
module knn_comb_BMR_W16_K3_N128 ( p_input, o );
  input [2063:0] p_input;
  output [47:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
         n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
         n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
         n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
         n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
         n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507,
         n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
         n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
         n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
         n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539,
         n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
         n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555,
         n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
         n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
         n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579,
         n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
         n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
         n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
         n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611,
         n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
         n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
         n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
         n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
         n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
         n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683,
         n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
         n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
         n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755,
         n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
         n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
         n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
         n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
         n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827,
         n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
         n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843,
         n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
         n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
         n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891,
         n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899,
         n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
         n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
         n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
         n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987,
         n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
         n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
         n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
         n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
         n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
         n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
         n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
         n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059,
         n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
         n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
         n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083,
         n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
         n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
         n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
         n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
         n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
         n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131,
         n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
         n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
         n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155,
         n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
         n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
         n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
         n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
         n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203,
         n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
         n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
         n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
         n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
         n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
         n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
         n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
         n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275,
         n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
         n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
         n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299,
         n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
         n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
         n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
         n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
         n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
         n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
         n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
         n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
         n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395,
         n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
         n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
         n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419,
         n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
         n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
         n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443,
         n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
         n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
         n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
         n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
         n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
         n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491,
         n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
         n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
         n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
         n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
         n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
         n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539,
         n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
         n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
         n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563,
         n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
         n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
         n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587,
         n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
         n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603,
         n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611,
         n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
         n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
         n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635,
         n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
         n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651,
         n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659,
         n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
         n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675,
         n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683,
         n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
         n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
         n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707,
         n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
         n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723,
         n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731,
         n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
         n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
         n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755,
         n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
         n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779,
         n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
         n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795,
         n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803,
         n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
         n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
         n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827,
         n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
         n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
         n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851,
         n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
         n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
         n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875,
         n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
         n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
         n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899,
         n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907,
         n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
         n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923,
         n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
         n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939,
         n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
         n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955,
         n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
         n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971,
         n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979,
         n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
         n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
         n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
         n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
         n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
         n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
         n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035,
         n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043,
         n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051,
         n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
         n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
         n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
         n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083,
         n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
         n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
         n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
         n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115,
         n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
         n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
         n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
         n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
         n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
         n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187,
         n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
         n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
         n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211,
         n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
         n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
         n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
         n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
         n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259,
         n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
         n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
         n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
         n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
         n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
         n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307,
         n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
         n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
         n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331,
         n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
         n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
         n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355,
         n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
         n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
         n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379,
         n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387,
         n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395,
         n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403,
         n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
         n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
         n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427,
         n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
         n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
         n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
         n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499,
         n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
         n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
         n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523,
         n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531,
         n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539,
         n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547,
         n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
         n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
         n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571,
         n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
         n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
         n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595,
         n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
         n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
         n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
         n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643,
         n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
         n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
         n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667,
         n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675,
         n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
         n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691,
         n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
         n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
         n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715,
         n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
         n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
         n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739,
         n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747,
         n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755,
         n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763,
         n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771,
         n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
         n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787,
         n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
         n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803,
         n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811,
         n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
         n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827,
         n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835,
         n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843,
         n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
         n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859,
         n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
         n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875,
         n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883,
         n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891,
         n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899,
         n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907,
         n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
         n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
         n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931,
         n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
         n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947,
         n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955,
         n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
         n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
         n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
         n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987,
         n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
         n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003,
         n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
         n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019,
         n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027,
         n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035,
         n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
         n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
         n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059,
         n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
         n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075,
         n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
         n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091,
         n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099,
         n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
         n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
         n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123,
         n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131,
         n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
         n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147,
         n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
         n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
         n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171,
         n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
         n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
         n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195,
         n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203,
         n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
         n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
         n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
         n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
         n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243,
         n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251,
         n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
         n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267,
         n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275,
         n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
         n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291,
         n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
         n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307,
         n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315,
         n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
         n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
         n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
         n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347,
         n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
         n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363,
         n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
         n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379,
         n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387,
         n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
         n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
         n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
         n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419,
         n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
         n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
         n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
         n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
         n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
         n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
         n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
         n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
         n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
         n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
         n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
         n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579,
         n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
         n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
         n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603,
         n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
         n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
         n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
         n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635,
         n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
         n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
         n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
         n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675,
         n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
         n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
         n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
         n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707,
         n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
         n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723,
         n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
         n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
         n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
         n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
         n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
         n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795,
         n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
         n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
         n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
         n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
         n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
         n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
         n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
         n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
         n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
         n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923,
         n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
         n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
         n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
         n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
         n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
         n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
         n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
         n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
         n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995,
         n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
         n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011,
         n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
         n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
         n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
         n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
         n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
         n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059,
         n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067,
         n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
         n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
         n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
         n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
         n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
         n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131,
         n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139,
         n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
         n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155,
         n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
         n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
         n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179,
         n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
         n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
         n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203,
         n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211,
         n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
         n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227,
         n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
         n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
         n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251,
         n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
         n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
         n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275,
         n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
         n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
         n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
         n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323,
         n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
         n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
         n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347,
         n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355,
         n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
         n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371,
         n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
         n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
         n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395,
         n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
         n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411,
         n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419,
         n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
         n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
         n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443,
         n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
         n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
         n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467,
         n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
         n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483,
         n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491,
         n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499,
         n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
         n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515,
         n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
         n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531,
         n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539,
         n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
         n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555,
         n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563,
         n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571,
         n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
         n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587,
         n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
         n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603,
         n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
         n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619,
         n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627,
         n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635,
         n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643,
         n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
         n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659,
         n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
         n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675,
         n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683,
         n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691,
         n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
         n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707,
         n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
         n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
         n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731,
         n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
         n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747,
         n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755,
         n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763,
         n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771,
         n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779,
         n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
         n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
         n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803,
         n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
         n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819,
         n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827,
         n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835,
         n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843,
         n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851,
         n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859,
         n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
         n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
         n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
         n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891,
         n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899,
         n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
         n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915,
         n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923,
         n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931,
         n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
         n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947,
         n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
         n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
         n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971,
         n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
         n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
         n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995,
         n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003,
         n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
         n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019,
         n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
         n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
         n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043,
         n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
         n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059,
         n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067,
         n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075,
         n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
         n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091,
         n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
         n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107,
         n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115,
         n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
         n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131,
         n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139,
         n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147,
         n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
         n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163,
         n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
         n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179,
         n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187,
         n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
         n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203,
         n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
         n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219,
         n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
         n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235,
         n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
         n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251,
         n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259,
         n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267,
         n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
         n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
         n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291,
         n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
         n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307,
         n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
         n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323,
         n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331,
         n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
         n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347,
         n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355,
         n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363,
         n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
         n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379,
         n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
         n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395,
         n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403,
         n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
         n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
         n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427,
         n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435,
         n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
         n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451,
         n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
         n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
         n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475,
         n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483,
         n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491,
         n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499,
         n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507,
         n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
         n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523,
         n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
         n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
         n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547,
         n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
         n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563,
         n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571,
         n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579,
         n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
         n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595,
         n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
         n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611,
         n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619,
         n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
         n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635,
         n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643,
         n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651,
         n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
         n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667,
         n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
         n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683,
         n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691,
         n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699,
         n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707,
         n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715,
         n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723,
         n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
         n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739,
         n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
         n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
         n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
         n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
         n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787,
         n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
         n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
         n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811,
         n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
         n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827,
         n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835,
         n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843,
         n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851,
         n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
         n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
         n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883,
         n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
         n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899,
         n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907,
         n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
         n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
         n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931,
         n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
         n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
         n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955,
         n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
         n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971,
         n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979,
         n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
         n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
         n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
         n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011,
         n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
         n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027,
         n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
         n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
         n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
         n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
         n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067,
         n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
         n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083,
         n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
         n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099,
         n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
         n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
         n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
         n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131,
         n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139,
         n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147,
         n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155,
         n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
         n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171,
         n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
         n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
         n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195,
         n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203,
         n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211,
         n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219,
         n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227,
         n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
         n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243,
         n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
         n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259,
         n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267,
         n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275,
         n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
         n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291,
         n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299,
         n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
         n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
         n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
         n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331,
         n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339,
         n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347,
         n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
         n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363,
         n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371,
         n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
         n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
         n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
         n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403,
         n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411,
         n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419,
         n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
         n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
         n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443,
         n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
         n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
         n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
         n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475,
         n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483,
         n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491,
         n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
         n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507,
         n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515,
         n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
         n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531,
         n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
         n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547,
         n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555,
         n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563,
         n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
         n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579,
         n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587,
         n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
         n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603,
         n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
         n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619,
         n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627,
         n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
         n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
         n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651,
         n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659,
         n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
         n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
         n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
         n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
         n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699,
         n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
         n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
         n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723,
         n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731,
         n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
         n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
         n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
         n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
         n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771,
         n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
         n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
         n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
         n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
         n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
         n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
         n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
         n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
         n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
         n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
         n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859,
         n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867,
         n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875,
         n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
         n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891,
         n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
         n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
         n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915,
         n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
         n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987,
         n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
         n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
         n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011,
         n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
         n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
         n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
         n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
         n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
         n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059,
         n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
         n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
         n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
         n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091,
         n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
         n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
         n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
         n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
         n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
         n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155,
         n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163,
         n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
         n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179,
         n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
         n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
         n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
         n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
         n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227,
         n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
         n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
         n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251,
         n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
         n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
         n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
         n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283,
         n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291,
         n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299,
         n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307,
         n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
         n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323,
         n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
         n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
         n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
         n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
         n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371,
         n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379,
         n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
         n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395,
         n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
         n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411,
         n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419,
         n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
         n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435,
         n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443,
         n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451,
         n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
         n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467,
         n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
         n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483,
         n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
         n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499,
         n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507,
         n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515,
         n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523,
         n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531,
         n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539,
         n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547,
         n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555,
         n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563,
         n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571,
         n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579,
         n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587,
         n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595,
         n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603,
         n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611,
         n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619,
         n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
         n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635,
         n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643,
         n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651,
         n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659,
         n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667,
         n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675,
         n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683,
         n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
         n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699,
         n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707,
         n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715,
         n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723,
         n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731,
         n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739,
         n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747,
         n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755,
         n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763,
         n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771,
         n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779,
         n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787,
         n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795,
         n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803,
         n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811,
         n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819,
         n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827,
         n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835,
         n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
         n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851,
         n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
         n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
         n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875,
         n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
         n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
         n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899,
         n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907,
         n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915,
         n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923,
         n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931,
         n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939,
         n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947,
         n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955,
         n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963,
         n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971,
         n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
         n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987,
         n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995,
         n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003,
         n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011,
         n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019,
         n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027,
         n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035,
         n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043,
         n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
         n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059,
         n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067,
         n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075,
         n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083,
         n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091,
         n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099,
         n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
         n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115,
         n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
         n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131,
         n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139,
         n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147,
         n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155,
         n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163,
         n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171,
         n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179,
         n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187,
         n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195,
         n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203,
         n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211,
         n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219,
         n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227,
         n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235,
         n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243,
         n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251,
         n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259,
         n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
         n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275,
         n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283,
         n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291,
         n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299,
         n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307,
         n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315,
         n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
         n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331,
         n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
         n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
         n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355,
         n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363,
         n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371,
         n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379,
         n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387,
         n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395,
         n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403,
         n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411,
         n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419,
         n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427,
         n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435,
         n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443,
         n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451,
         n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459,
         n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467,
         n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475,
         n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483,
         n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491,
         n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499,
         n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507,
         n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515,
         n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523,
         n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531,
         n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
         n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547,
         n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
         n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563,
         n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571,
         n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579,
         n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587,
         n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595,
         n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603,
         n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
         n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619,
         n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627,
         n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635,
         n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643,
         n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651,
         n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659,
         n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667,
         n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675,
         n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683,
         n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691,
         n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699,
         n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707,
         n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715,
         n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723,
         n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731,
         n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739,
         n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747,
         n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
         n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763,
         n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771,
         n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779,
         n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787,
         n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795,
         n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
         n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811,
         n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819,
         n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
         n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835,
         n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
         n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851,
         n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859,
         n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867,
         n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875,
         n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883,
         n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891,
         n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
         n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907,
         n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915,
         n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923,
         n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931,
         n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939,
         n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947,
         n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955,
         n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963,
         n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
         n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979,
         n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987,
         n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
         n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003,
         n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011,
         n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019,
         n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027,
         n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035,
         n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
         n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051,
         n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
         n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067,
         n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075,
         n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083,
         n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091,
         n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099,
         n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107,
         n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
         n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123,
         n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131,
         n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139,
         n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147,
         n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155,
         n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163,
         n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171,
         n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179,
         n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
         n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195,
         n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
         n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211,
         n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219,
         n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227,
         n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235,
         n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243,
         n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251,
         n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259,
         n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267,
         n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275,
         n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283,
         n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291,
         n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299,
         n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307,
         n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315,
         n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
         n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331,
         n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339,
         n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
         n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355,
         n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363,
         n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371,
         n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379,
         n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387,
         n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395,
         n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403,
         n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411,
         n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419,
         n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427,
         n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435,
         n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443,
         n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451,
         n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459,
         n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467,
         n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475,
         n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483,
         n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
         n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499,
         n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507,
         n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
         n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523,
         n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531,
         n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539,
         n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
         n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555,
         n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
         n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
         n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579,
         n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
         n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595,
         n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603,
         n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611,
         n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
         n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627,
         n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
         n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643,
         n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651,
         n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659,
         n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667,
         n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675,
         n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683,
         n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
         n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699,
         n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707,
         n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715,
         n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723,
         n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731,
         n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739,
         n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747,
         n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755,
         n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763,
         n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771,
         n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
         n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787,
         n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795,
         n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803,
         n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811,
         n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819,
         n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827,
         n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
         n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843,
         n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851,
         n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859,
         n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867,
         n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875,
         n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883,
         n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891,
         n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899,
         n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
         n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915,
         n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923,
         n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931,
         n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
         n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947,
         n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955,
         n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963,
         n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971,
         n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979,
         n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987,
         n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
         n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
         n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011,
         n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019,
         n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027,
         n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035,
         n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043,
         n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051,
         n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059,
         n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
         n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075,
         n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083,
         n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091,
         n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099,
         n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107,
         n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115,
         n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123,
         n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131,
         n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
         n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147,
         n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155,
         n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163,
         n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171,
         n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179,
         n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187,
         n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
         n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203,
         n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
         n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219,
         n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227,
         n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235,
         n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243,
         n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251,
         n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259,
         n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
         n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275,
         n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
         n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291,
         n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299,
         n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307,
         n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315,
         n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323,
         n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331,
         n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339,
         n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347,
         n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
         n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363,
         n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371,
         n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379,
         n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387,
         n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395,
         n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403,
         n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411,
         n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419,
         n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
         n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435,
         n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443,
         n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451,
         n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459,
         n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467,
         n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475,
         n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
         n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
         n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
         n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507,
         n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515,
         n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523,
         n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531,
         n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539,
         n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547,
         n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
         n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
         n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
         n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
         n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587,
         n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
         n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603,
         n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611,
         n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
         n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
         n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
         n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
         n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
         n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659,
         n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667,
         n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675,
         n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683,
         n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691,
         n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
         n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
         n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
         n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723,
         n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731,
         n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739,
         n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747,
         n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755,
         n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763,
         n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
         n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779,
         n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
         n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795,
         n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803,
         n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
         n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819,
         n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827,
         n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835,
         n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
         n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851,
         n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
         n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867,
         n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875,
         n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
         n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891,
         n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
         n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907,
         n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
         n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923,
         n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
         n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
         n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947,
         n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
         n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963,
         n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971,
         n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979,
         n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
         n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995,
         n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
         n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
         n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019,
         n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027,
         n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035,
         n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043,
         n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051,
         n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
         n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067,
         n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
         n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083,
         n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091,
         n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099,
         n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107,
         n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115,
         n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123,
         n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
         n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139,
         n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
         n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155,
         n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163,
         n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171,
         n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179,
         n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
         n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195,
         n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
         n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211,
         n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
         n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227,
         n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235,
         n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243,
         n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251,
         n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259,
         n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267,
         n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
         n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283,
         n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
         n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299,
         n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307,
         n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
         n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323,
         n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
         n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339,
         n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
         n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355,
         n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
         n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371,
         n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379,
         n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387,
         n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395,
         n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403,
         n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411,
         n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419,
         n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427,
         n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435,
         n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443,
         n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451,
         n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459,
         n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467,
         n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475,
         n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483,
         n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491,
         n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499,
         n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
         n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515,
         n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523,
         n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531,
         n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539,
         n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547,
         n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555,
         n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563,
         n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
         n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579,
         n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587,
         n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595,
         n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603,
         n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611,
         n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619,
         n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627,
         n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
         n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643,
         n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
         n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659,
         n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667,
         n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675,
         n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683,
         n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691,
         n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699,
         n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707,
         n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715,
         n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723,
         n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731,
         n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739,
         n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747,
         n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755,
         n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763,
         n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771,
         n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779,
         n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787,
         n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
         n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
         n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811,
         n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819,
         n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827,
         n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835,
         n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843,
         n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851,
         n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859,
         n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867,
         n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875,
         n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883,
         n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
         n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899,
         n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907,
         n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915,
         n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
         n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931,
         n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
         n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
         n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955,
         n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963,
         n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971,
         n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979,
         n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987,
         n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995,
         n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003,
         n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011,
         n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019,
         n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027,
         n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035,
         n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043,
         n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051,
         n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059,
         n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
         n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075,
         n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083,
         n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091,
         n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099,
         n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107,
         n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115,
         n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123,
         n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131,
         n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139,
         n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147,
         n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
         n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163,
         n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171,
         n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179,
         n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187,
         n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195,
         n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203,
         n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211,
         n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219,
         n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
         n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235,
         n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243,
         n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251,
         n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259,
         n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267,
         n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275,
         n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283,
         n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291,
         n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
         n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
         n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315,
         n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323,
         n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331,
         n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339,
         n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347,
         n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
         n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363,
         n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371,
         n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379,
         n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387,
         n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395,
         n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403,
         n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411,
         n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419,
         n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427,
         n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435,
         n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
         n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451,
         n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459,
         n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467,
         n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475,
         n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483,
         n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491,
         n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
         n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507,
         n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
         n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
         n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531,
         n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539,
         n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547,
         n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555,
         n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563,
         n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
         n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579,
         n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587,
         n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595,
         n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603,
         n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611,
         n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619,
         n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627,
         n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635,
         n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643,
         n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651,
         n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659,
         n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667,
         n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675,
         n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683,
         n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691,
         n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699,
         n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707,
         n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715,
         n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723,
         n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731,
         n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739,
         n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747,
         n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755,
         n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763,
         n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771,
         n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779,
         n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787,
         n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795,
         n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803,
         n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811,
         n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819,
         n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827,
         n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835,
         n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843,
         n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851,
         n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859,
         n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867,
         n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875,
         n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883,
         n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891,
         n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899,
         n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907,
         n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915,
         n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923,
         n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931,
         n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939,
         n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947,
         n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955,
         n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963,
         n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971,
         n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979,
         n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987,
         n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995,
         n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
         n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011,
         n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
         n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027,
         n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035,
         n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043,
         n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051,
         n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059,
         n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067,
         n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
         n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083,
         n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
         n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099,
         n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107,
         n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115,
         n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123,
         n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131,
         n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139,
         n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
         n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155,
         n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
         n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171,
         n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179,
         n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187,
         n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195,
         n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203,
         n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211,
         n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
         n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227,
         n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
         n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
         n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251,
         n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259,
         n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267,
         n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275,
         n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283,
         n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
         n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299,
         n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
         n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315,
         n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323,
         n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
         n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339,
         n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347,
         n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355,
         n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
         n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371,
         n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
         n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387,
         n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395,
         n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
         n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411,
         n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419,
         n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427,
         n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
         n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443,
         n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
         n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459,
         n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467,
         n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475,
         n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483,
         n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491,
         n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499,
         n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
         n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515,
         n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
         n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531,
         n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539,
         n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547,
         n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555,
         n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563,
         n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571,
         n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
         n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
         n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
         n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603,
         n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611,
         n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
         n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
         n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
         n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643,
         n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
         n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659,
         n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
         n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
         n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683,
         n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
         n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699,
         n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707,
         n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
         n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
         n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731,
         n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
         n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747,
         n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
         n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
         n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771,
         n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779,
         n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787,
         n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
         n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803,
         n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
         n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819,
         n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827,
         n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
         n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
         n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851,
         n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859,
         n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
         n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875,
         n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
         n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891,
         n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899,
         n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
         n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915,
         n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923,
         n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931,
         n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
         n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947,
         n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
         n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963,
         n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
         n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
         n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987,
         n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995,
         n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003,
         n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
         n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019,
         n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
         n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035,
         n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043,
         n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
         n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059,
         n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067,
         n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075,
         n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
         n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091,
         n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
         n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107,
         n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115,
         n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
         n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131,
         n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139,
         n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147,
         n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
         n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163,
         n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
         n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179,
         n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187,
         n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
         n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
         n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211,
         n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219,
         n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
         n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235,
         n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
         n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251,
         n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259,
         n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
         n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275,
         n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283,
         n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291,
         n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
         n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307,
         n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
         n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323,
         n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331,
         n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
         n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347,
         n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355,
         n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363,
         n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
         n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379,
         n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
         n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
         n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403,
         n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
         n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419,
         n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427,
         n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435,
         n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
         n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451,
         n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
         n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467,
         n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475,
         n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
         n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491,
         n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499,
         n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507,
         n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
         n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523,
         n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
         n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539,
         n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547,
         n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
         n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563,
         n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571,
         n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579,
         n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
         n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595,
         n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
         n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611,
         n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619,
         n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
         n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635,
         n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643,
         n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651,
         n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
         n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667,
         n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
         n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683,
         n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691,
         n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
         n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707,
         n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715,
         n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723,
         n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
         n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739,
         n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
         n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755,
         n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763,
         n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
         n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779,
         n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787,
         n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795,
         n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
         n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811,
         n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
         n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827,
         n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835,
         n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
         n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851,
         n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859,
         n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867,
         n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
         n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883,
         n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
         n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899,
         n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907,
         n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
         n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923,
         n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931,
         n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939,
         n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
         n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955,
         n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
         n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971,
         n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979,
         n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
         n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995,
         n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003,
         n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011,
         n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
         n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027,
         n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
         n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043,
         n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051,
         n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
         n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067,
         n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075,
         n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083,
         n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
         n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099,
         n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
         n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115,
         n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123,
         n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
         n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139,
         n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147,
         n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155,
         n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
         n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171,
         n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
         n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187,
         n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195,
         n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
         n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211,
         n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219,
         n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227,
         n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
         n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243,
         n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251,
         n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259,
         n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267,
         n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275,
         n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283,
         n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291,
         n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299,
         n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307,
         n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315,
         n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
         n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331,
         n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339,
         n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347,
         n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355,
         n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363,
         n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371,
         n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379,
         n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387,
         n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
         n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403,
         n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411,
         n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419,
         n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427,
         n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435,
         n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443,
         n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
         n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459,
         n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467,
         n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475,
         n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483,
         n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491,
         n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499,
         n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507,
         n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515,
         n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523,
         n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531,
         n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539,
         n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547,
         n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555,
         n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563,
         n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571,
         n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579,
         n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587,
         n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595,
         n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603,
         n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611,
         n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619,
         n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627,
         n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635,
         n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643,
         n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651,
         n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659,
         n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667,
         n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675,
         n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683,
         n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691,
         n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699,
         n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707,
         n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715,
         n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723,
         n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731,
         n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739,
         n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747,
         n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755,
         n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763,
         n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771,
         n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779,
         n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787,
         n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795,
         n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803,
         n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811,
         n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819,
         n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827,
         n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835,
         n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843,
         n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851,
         n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859,
         n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867,
         n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875,
         n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883,
         n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891,
         n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
         n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907,
         n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915,
         n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923,
         n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931,
         n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939,
         n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947,
         n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955,
         n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963,
         n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971,
         n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979,
         n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987,
         n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995,
         n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003,
         n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011,
         n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019,
         n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027,
         n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035,
         n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
         n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051,
         n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059,
         n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067,
         n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075,
         n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083,
         n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091,
         n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099,
         n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107,
         n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
         n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123,
         n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131,
         n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139,
         n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147,
         n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155,
         n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163,
         n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171,
         n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179,
         n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
         n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195,
         n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203,
         n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211,
         n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219,
         n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227,
         n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235,
         n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243,
         n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251,
         n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
         n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267,
         n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275,
         n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283,
         n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291,
         n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299,
         n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307,
         n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315,
         n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323,
         n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
         n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339,
         n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347,
         n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
         n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363,
         n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371,
         n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379,
         n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387,
         n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395,
         n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
         n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411,
         n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419,
         n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427,
         n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435,
         n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443,
         n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451,
         n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459,
         n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467,
         n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475,
         n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483,
         n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491,
         n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499,
         n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507,
         n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515,
         n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523,
         n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531,
         n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539,
         n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547,
         n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555,
         n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563,
         n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571,
         n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579,
         n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587,
         n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595,
         n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603,
         n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611,
         n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619,
         n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627,
         n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635,
         n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643,
         n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651,
         n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659,
         n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667,
         n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675,
         n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683,
         n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
         n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699,
         n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707,
         n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715,
         n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723,
         n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731,
         n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739,
         n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747,
         n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755,
         n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763,
         n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771,
         n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779,
         n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787,
         n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795,
         n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803,
         n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811,
         n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
         n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827,
         n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835,
         n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843,
         n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851,
         n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859,
         n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867,
         n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875,
         n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883,
         n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891,
         n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899,
         n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907,
         n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915,
         n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923,
         n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931,
         n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939,
         n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947,
         n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955,
         n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
         n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971,
         n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979,
         n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987,
         n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995,
         n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003,
         n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011,
         n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019,
         n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027,
         n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035,
         n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043,
         n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051,
         n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059,
         n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067,
         n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075,
         n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083,
         n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091,
         n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099,
         n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107,
         n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115,
         n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123,
         n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131,
         n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139,
         n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147,
         n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155,
         n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163,
         n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171,
         n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179,
         n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187,
         n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195,
         n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203,
         n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211,
         n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219,
         n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227,
         n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235,
         n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243,
         n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251,
         n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259,
         n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267,
         n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275,
         n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283,
         n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291,
         n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299,
         n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307,
         n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315,
         n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323,
         n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331,
         n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339,
         n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347,
         n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355,
         n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363,
         n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371,
         n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379,
         n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387,
         n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395,
         n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403,
         n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411,
         n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419,
         n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427,
         n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435,
         n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443,
         n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451,
         n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459,
         n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467,
         n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475,
         n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
         n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491,
         n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499,
         n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
         n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515,
         n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523,
         n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531,
         n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539,
         n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547,
         n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555,
         n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563,
         n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571,
         n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579,
         n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587,
         n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595,
         n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603,
         n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611,
         n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619,
         n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
         n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635,
         n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643,
         n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651,
         n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659,
         n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667,
         n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675,
         n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683,
         n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691,
         n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
         n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707,
         n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715,
         n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723,
         n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731,
         n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739,
         n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747,
         n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755,
         n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763,
         n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771,
         n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779,
         n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787,
         n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795,
         n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803,
         n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811,
         n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819,
         n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827,
         n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835,
         n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843,
         n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851,
         n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859,
         n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867,
         n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875,
         n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883,
         n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891,
         n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899,
         n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907,
         n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915,
         n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923,
         n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931,
         n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939,
         n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947,
         n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955,
         n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963,
         n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971,
         n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979,
         n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987,
         n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995,
         n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003,
         n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
         n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019,
         n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027,
         n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035,
         n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043,
         n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051,
         n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059,
         n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067,
         n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075,
         n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083,
         n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091,
         n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099,
         n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107,
         n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115,
         n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123,
         n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131,
         n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139,
         n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147,
         n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155,
         n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163,
         n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171,
         n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179,
         n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187,
         n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195,
         n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203,
         n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211,
         n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219,
         n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227,
         n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235,
         n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243,
         n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251,
         n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259,
         n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267,
         n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275,
         n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283,
         n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291,
         n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299,
         n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307,
         n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315,
         n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323,
         n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331,
         n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339,
         n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347,
         n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355,
         n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363,
         n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371,
         n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379,
         n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387,
         n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395,
         n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403,
         n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411,
         n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419,
         n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427,
         n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435,
         n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443,
         n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451,
         n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459,
         n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467,
         n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475,
         n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483,
         n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491,
         n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499,
         n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507,
         n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515,
         n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523,
         n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531,
         n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539,
         n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547,
         n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555,
         n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563,
         n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571,
         n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579,
         n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587,
         n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595,
         n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603,
         n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611,
         n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619,
         n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627,
         n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635,
         n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643,
         n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651,
         n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659,
         n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667,
         n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675,
         n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683,
         n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691,
         n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699,
         n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707,
         n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715,
         n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723,
         n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731,
         n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739,
         n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747,
         n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755,
         n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763,
         n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771,
         n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779,
         n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787,
         n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795,
         n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
         n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811,
         n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819,
         n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827,
         n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835,
         n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843,
         n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851,
         n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859,
         n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867,
         n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875,
         n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883,
         n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891,
         n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899,
         n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907,
         n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915,
         n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923,
         n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931,
         n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939,
         n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947,
         n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955,
         n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963,
         n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971,
         n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979,
         n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987,
         n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995,
         n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003,
         n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011,
         n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019,
         n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027,
         n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035,
         n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043,
         n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051,
         n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059,
         n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067,
         n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075,
         n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083,
         n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091,
         n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099,
         n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107,
         n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115,
         n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123,
         n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131,
         n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139,
         n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147,
         n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155,
         n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163,
         n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171,
         n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179,
         n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187,
         n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195,
         n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203,
         n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211,
         n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219,
         n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227,
         n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235,
         n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243,
         n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251,
         n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259,
         n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267,
         n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275,
         n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283,
         n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291,
         n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299,
         n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307,
         n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315,
         n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323,
         n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331,
         n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339,
         n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347,
         n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355,
         n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363,
         n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371,
         n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379,
         n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387,
         n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395,
         n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403,
         n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411,
         n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419,
         n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427,
         n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435,
         n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443,
         n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451,
         n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459,
         n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467,
         n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475,
         n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483,
         n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491,
         n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499,
         n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507,
         n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515,
         n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523,
         n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531,
         n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539,
         n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547,
         n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555,
         n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563,
         n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571,
         n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579,
         n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587,
         n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595,
         n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603,
         n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611,
         n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619,
         n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627,
         n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635,
         n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643,
         n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651,
         n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659,
         n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667,
         n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675,
         n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683,
         n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691,
         n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699,
         n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707,
         n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715,
         n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723,
         n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731,
         n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739,
         n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747,
         n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755,
         n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763,
         n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771,
         n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779,
         n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787,
         n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795,
         n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803,
         n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811,
         n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819,
         n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827,
         n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835,
         n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843,
         n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851,
         n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859,
         n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867,
         n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875,
         n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883,
         n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891,
         n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899,
         n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907,
         n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915,
         n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923,
         n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931,
         n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939,
         n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947,
         n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955,
         n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963,
         n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971,
         n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979,
         n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987,
         n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995,
         n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003,
         n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011,
         n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019,
         n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027,
         n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035,
         n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043,
         n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051,
         n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059,
         n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067,
         n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075,
         n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083,
         n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091,
         n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099,
         n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107,
         n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115,
         n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123,
         n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131,
         n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139,
         n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147,
         n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155,
         n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163,
         n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171,
         n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179,
         n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187,
         n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195,
         n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203,
         n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211,
         n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219,
         n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227,
         n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235,
         n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243,
         n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251,
         n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259,
         n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267,
         n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275,
         n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283,
         n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291,
         n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299,
         n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307,
         n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315,
         n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323,
         n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331,
         n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339,
         n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347,
         n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355,
         n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363,
         n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371,
         n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379,
         n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387,
         n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395,
         n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403,
         n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411,
         n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419,
         n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427,
         n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435,
         n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443,
         n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451,
         n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459,
         n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467,
         n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475,
         n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483,
         n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491,
         n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499,
         n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
         n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515,
         n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523,
         n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531,
         n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539,
         n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547,
         n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555,
         n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
         n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571,
         n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579,
         n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587,
         n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595,
         n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603,
         n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611,
         n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619,
         n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627,
         n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635,
         n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643,
         n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651,
         n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659,
         n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667,
         n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675,
         n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683,
         n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691,
         n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699,
         n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
         n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715,
         n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723,
         n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731,
         n50732, n50733, n50734, n50735, n50736, n50737, n50738, n50739,
         n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747,
         n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755,
         n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763,
         n50764, n50765, n50766, n50767, n50768, n50769, n50770, n50771,
         n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779,
         n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787,
         n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795,
         n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803,
         n50804, n50805, n50806, n50807, n50808, n50809, n50810, n50811,
         n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819,
         n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827,
         n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835,
         n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843,
         n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851,
         n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859,
         n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867,
         n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875,
         n50876, n50877, n50878, n50879, n50880, n50881, n50882, n50883,
         n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891,
         n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899,
         n50900, n50901, n50902, n50903, n50904, n50905, n50906, n50907,
         n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915,
         n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923,
         n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931,
         n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939,
         n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947,
         n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955,
         n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963,
         n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971,
         n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979,
         n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987,
         n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995,
         n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003,
         n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011,
         n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019,
         n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51027,
         n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035,
         n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043,
         n51044, n51045, n51046, n51047, n51048, n51049, n51050, n51051,
         n51052, n51053, n51054, n51055, n51056, n51057, n51058, n51059,
         n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067,
         n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075,
         n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083,
         n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091,
         n51092, n51093, n51094, n51095, n51096, n51097, n51098, n51099,
         n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107,
         n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115,
         n51116, n51117, n51118, n51119, n51120, n51121, n51122, n51123,
         n51124, n51125, n51126, n51127, n51128, n51129, n51130, n51131,
         n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139,
         n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147,
         n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155,
         n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163,
         n51164, n51165, n51166, n51167, n51168, n51169, n51170, n51171,
         n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179,
         n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187,
         n51188, n51189, n51190, n51191, n51192, n51193, n51194, n51195,
         n51196, n51197, n51198, n51199, n51200, n51201, n51202, n51203,
         n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211,
         n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219,
         n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227,
         n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235,
         n51236, n51237, n51238, n51239, n51240, n51241, n51242, n51243,
         n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251,
         n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259,
         n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267,
         n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275,
         n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283,
         n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291,
         n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299,
         n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307,
         n51308, n51309, n51310, n51311, n51312, n51313, n51314, n51315,
         n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323,
         n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331,
         n51332, n51333, n51334, n51335, n51336, n51337, n51338, n51339,
         n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347,
         n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355,
         n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363,
         n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371,
         n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379,
         n51380, n51381, n51382, n51383, n51384, n51385, n51386, n51387,
         n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395,
         n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403,
         n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411,
         n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419,
         n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427,
         n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435,
         n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443,
         n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451,
         n51452, n51453, n51454, n51455, n51456, n51457, n51458, n51459,
         n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467,
         n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475,
         n51476, n51477, n51478, n51479, n51480, n51481, n51482, n51483,
         n51484, n51485, n51486, n51487, n51488, n51489, n51490, n51491,
         n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499,
         n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507,
         n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515,
         n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523,
         n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531,
         n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539,
         n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547,
         n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555,
         n51556, n51557, n51558, n51559, n51560, n51561, n51562, n51563,
         n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571,
         n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579,
         n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587,
         n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595,
         n51596, n51597, n51598, n51599, n51600, n51601, n51602, n51603,
         n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611,
         n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619,
         n51620, n51621, n51622, n51623, n51624, n51625, n51626, n51627,
         n51628, n51629, n51630, n51631, n51632, n51633, n51634, n51635,
         n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643,
         n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651,
         n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659,
         n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667,
         n51668, n51669, n51670, n51671, n51672, n51673, n51674, n51675,
         n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683,
         n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691,
         n51692, n51693, n51694, n51695, n51696, n51697, n51698, n51699,
         n51700, n51701, n51702, n51703, n51704, n51705, n51706, n51707,
         n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715,
         n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723,
         n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731,
         n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739,
         n51740, n51741, n51742, n51743, n51744, n51745, n51746, n51747,
         n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755,
         n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763,
         n51764, n51765, n51766, n51767, n51768, n51769, n51770, n51771,
         n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779,
         n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787,
         n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795,
         n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803,
         n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811,
         n51812, n51813, n51814, n51815, n51816, n51817, n51818, n51819,
         n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827,
         n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835,
         n51836, n51837, n51838, n51839, n51840, n51841, n51842, n51843,
         n51844, n51845, n51846, n51847, n51848, n51849, n51850, n51851,
         n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859,
         n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867,
         n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875,
         n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883,
         n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51891,
         n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899,
         n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907,
         n51908, n51909, n51910, n51911, n51912, n51913, n51914, n51915,
         n51916, n51917, n51918, n51919, n51920, n51921, n51922, n51923,
         n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931,
         n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939,
         n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947,
         n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955,
         n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963,
         n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971,
         n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979,
         n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987,
         n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995,
         n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003,
         n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011,
         n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019,
         n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027,
         n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035,
         n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043,
         n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051,
         n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059,
         n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067,
         n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075,
         n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083,
         n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091,
         n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099,
         n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107,
         n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115,
         n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123,
         n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131,
         n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139,
         n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147,
         n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155,
         n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163,
         n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171,
         n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179,
         n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187,
         n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195,
         n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203,
         n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211,
         n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219,
         n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227,
         n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235,
         n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243,
         n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251,
         n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259,
         n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267,
         n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275,
         n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283,
         n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291,
         n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299,
         n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307,
         n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315,
         n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323,
         n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331,
         n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339,
         n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347,
         n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355,
         n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363,
         n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371,
         n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379,
         n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387,
         n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395,
         n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403,
         n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411,
         n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419,
         n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427,
         n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435,
         n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443,
         n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451,
         n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459,
         n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467,
         n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475,
         n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483,
         n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491,
         n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499,
         n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507,
         n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515,
         n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523,
         n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531,
         n52532, n52533, n52534, n52535, n52536, n52537, n52538, n52539,
         n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547,
         n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555,
         n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563,
         n52564, n52565, n52566, n52567, n52568, n52569, n52570, n52571,
         n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579,
         n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587,
         n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595,
         n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603,
         n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611,
         n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619,
         n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627,
         n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635,
         n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643,
         n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651,
         n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659,
         n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667,
         n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675,
         n52676, n52677, n52678, n52679, n52680, n52681, n52682, n52683,
         n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691,
         n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699,
         n52700, n52701, n52702, n52703, n52704, n52705, n52706, n52707,
         n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715,
         n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723,
         n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731,
         n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739,
         n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747,
         n52748, n52749, n52750, n52751, n52752, n52753, n52754, n52755,
         n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763,
         n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771,
         n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779,
         n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787,
         n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795,
         n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803,
         n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811,
         n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819,
         n52820, n52821, n52822, n52823, n52824, n52825, n52826, n52827,
         n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835,
         n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843,
         n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851,
         n52852, n52853, n52854, n52855, n52856, n52857, n52858, n52859,
         n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867,
         n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875,
         n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883,
         n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891,
         n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899,
         n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907,
         n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915,
         n52916, n52917, n52918, n52919, n52920, n52921, n52922, n52923,
         n52924, n52925, n52926, n52927, n52928, n52929, n52930, n52931,
         n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939,
         n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947,
         n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955,
         n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963,
         n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971,
         n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979,
         n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987,
         n52988, n52989, n52990, n52991, n52992, n52993, n52994, n52995,
         n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003,
         n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011,
         n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019,
         n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027,
         n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035,
         n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043,
         n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051,
         n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059,
         n53060, n53061, n53062, n53063, n53064, n53065, n53066, n53067,
         n53068, n53069, n53070, n53071, n53072, n53073, n53074, n53075,
         n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083,
         n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091,
         n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099,
         n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107,
         n53108, n53109, n53110, n53111, n53112, n53113, n53114, n53115,
         n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123,
         n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131,
         n53132, n53133, n53134, n53135, n53136, n53137, n53138, n53139,
         n53140, n53141, n53142, n53143, n53144, n53145, n53146, n53147,
         n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155,
         n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163,
         n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171,
         n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179,
         n53180, n53181, n53182, n53183, n53184, n53185, n53186, n53187,
         n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195,
         n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203,
         n53204, n53205, n53206, n53207, n53208, n53209, n53210, n53211,
         n53212, n53213, n53214, n53215, n53216, n53217, n53218, n53219,
         n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227,
         n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235,
         n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243,
         n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251,
         n53252, n53253, n53254, n53255, n53256, n53257, n53258, n53259,
         n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267,
         n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275,
         n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283,
         n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291,
         n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299,
         n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307,
         n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315,
         n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323,
         n53324, n53325, n53326, n53327, n53328, n53329, n53330, n53331,
         n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339,
         n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347,
         n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355,
         n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363,
         n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371,
         n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379,
         n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387,
         n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395,
         n53396, n53397, n53398, n53399, n53400, n53401, n53402, n53403,
         n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411,
         n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419,
         n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427,
         n53428, n53429, n53430, n53431, n53432, n53433, n53434, n53435,
         n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443,
         n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451,
         n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459,
         n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467,
         n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475,
         n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483,
         n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491,
         n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499,
         n53500, n53501, n53502, n53503, n53504, n53505, n53506, n53507,
         n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515,
         n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523,
         n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531,
         n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539,
         n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547,
         n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555,
         n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563,
         n53564, n53565, n53566, n53567, n53568, n53569, n53570, n53571,
         n53572, n53573, n53574, n53575, n53576, n53577, n53578, n53579,
         n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587,
         n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595,
         n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603,
         n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611,
         n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619,
         n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627,
         n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635,
         n53636, n53637, n53638, n53639, n53640, n53641, n53642, n53643,
         n53644, n53645, n53646, n53647, n53648, n53649, n53650, n53651,
         n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659,
         n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667,
         n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675,
         n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683,
         n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691,
         n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699,
         n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707,
         n53708, n53709, n53710, n53711, n53712, n53713, n53714, n53715,
         n53716, n53717, n53718, n53719, n53720, n53721, n53722, n53723,
         n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731,
         n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739,
         n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747,
         n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755,
         n53756, n53757, n53758, n53759, n53760, n53761, n53762, n53763,
         n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771,
         n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779,
         n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787,
         n53788, n53789, n53790, n53791, n53792, n53793, n53794, n53795,
         n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803,
         n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811,
         n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819,
         n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827,
         n53828, n53829, n53830, n53831, n53832, n53833, n53834, n53835,
         n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843,
         n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851,
         n53852, n53853, n53854, n53855, n53856, n53857, n53858, n53859,
         n53860, n53861, n53862, n53863, n53864, n53865, n53866, n53867,
         n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875,
         n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883,
         n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891,
         n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899,
         n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907,
         n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915,
         n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923,
         n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931,
         n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939,
         n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947,
         n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955,
         n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963,
         n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971,
         n53972, n53973, n53974, n53975, n53976, n53977, n53978, n53979,
         n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987,
         n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995,
         n53996, n53997, n53998, n53999, n54000, n54001, n54002, n54003,
         n54004, n54005, n54006, n54007, n54008, n54009, n54010, n54011,
         n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019,
         n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027,
         n54028, n54029, n54030, n54031, n54032, n54033, n54034, n54035,
         n54036, n54037, n54038, n54039, n54040, n54041, n54042, n54043,
         n54044, n54045, n54046, n54047, n54048, n54049, n54050, n54051,
         n54052, n54053, n54054, n54055, n54056, n54057, n54058, n54059,
         n54060, n54061, n54062, n54063, n54064, n54065, n54066, n54067,
         n54068, n54069, n54070, n54071, n54072, n54073, n54074, n54075,
         n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083,
         n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091,
         n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099,
         n54100, n54101, n54102, n54103, n54104, n54105, n54106, n54107,
         n54108, n54109, n54110, n54111, n54112, n54113, n54114, n54115,
         n54116, n54117, n54118, n54119, n54120, n54121, n54122, n54123,
         n54124, n54125, n54126, n54127, n54128, n54129, n54130, n54131,
         n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139,
         n54140, n54141, n54142, n54143, n54144, n54145, n54146, n54147,
         n54148, n54149, n54150, n54151, n54152, n54153, n54154, n54155,
         n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163,
         n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171,
         n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179,
         n54180, n54181, n54182, n54183, n54184, n54185, n54186, n54187,
         n54188, n54189, n54190, n54191, n54192, n54193, n54194, n54195,
         n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203,
         n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211,
         n54212, n54213, n54214, n54215, n54216, n54217, n54218, n54219,
         n54220, n54221, n54222, n54223, n54224, n54225, n54226, n54227,
         n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235,
         n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243,
         n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251,
         n54252, n54253, n54254, n54255, n54256, n54257, n54258, n54259,
         n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267,
         n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275,
         n54276, n54277, n54278, n54279, n54280, n54281, n54282, n54283,
         n54284, n54285, n54286, n54287, n54288, n54289, n54290, n54291,
         n54292, n54293, n54294, n54295, n54296, n54297, n54298, n54299,
         n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307,
         n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315,
         n54316, n54317, n54318, n54319, n54320, n54321, n54322, n54323,
         n54324, n54325, n54326, n54327, n54328, n54329, n54330, n54331,
         n54332, n54333, n54334, n54335, n54336, n54337, n54338, n54339,
         n54340, n54341, n54342, n54343, n54344, n54345, n54346, n54347,
         n54348, n54349, n54350, n54351, n54352, n54353, n54354, n54355,
         n54356, n54357, n54358, n54359, n54360, n54361, n54362, n54363,
         n54364, n54365, n54366, n54367, n54368, n54369, n54370, n54371,
         n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379,
         n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387,
         n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395,
         n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403,
         n54404, n54405, n54406, n54407, n54408, n54409, n54410, n54411,
         n54412, n54413, n54414, n54415, n54416, n54417, n54418, n54419,
         n54420, n54421, n54422, n54423, n54424, n54425, n54426, n54427,
         n54428, n54429, n54430, n54431, n54432, n54433, n54434, n54435,
         n54436, n54437, n54438, n54439, n54440, n54441, n54442, n54443,
         n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451,
         n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459,
         n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467,
         n54468, n54469, n54470, n54471, n54472, n54473, n54474, n54475,
         n54476, n54477, n54478, n54479, n54480, n54481, n54482, n54483,
         n54484, n54485, n54486, n54487, n54488, n54489, n54490, n54491,
         n54492, n54493, n54494, n54495, n54496, n54497, n54498, n54499,
         n54500, n54501, n54502, n54503, n54504, n54505, n54506, n54507,
         n54508, n54509, n54510, n54511, n54512, n54513, n54514, n54515,
         n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523,
         n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531,
         n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539,
         n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547,
         n54548, n54549, n54550, n54551, n54552, n54553, n54554, n54555,
         n54556, n54557, n54558, n54559, n54560, n54561, n54562, n54563,
         n54564, n54565, n54566, n54567, n54568, n54569, n54570, n54571,
         n54572, n54573, n54574, n54575, n54576, n54577, n54578, n54579,
         n54580, n54581, n54582, n54583, n54584, n54585, n54586, n54587,
         n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595,
         n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603,
         n54604, n54605, n54606, n54607, n54608, n54609, n54610, n54611,
         n54612, n54613, n54614, n54615, n54616, n54617, n54618, n54619,
         n54620, n54621, n54622, n54623, n54624, n54625, n54626, n54627,
         n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635,
         n54636, n54637, n54638, n54639, n54640, n54641, n54642, n54643,
         n54644, n54645, n54646, n54647, n54648, n54649, n54650, n54651,
         n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659,
         n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667,
         n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675,
         n54676, n54677, n54678, n54679, n54680, n54681, n54682, n54683,
         n54684, n54685, n54686, n54687, n54688, n54689, n54690, n54691,
         n54692, n54693, n54694, n54695, n54696, n54697, n54698, n54699,
         n54700, n54701, n54702, n54703, n54704, n54705, n54706, n54707,
         n54708, n54709, n54710, n54711, n54712, n54713, n54714, n54715,
         n54716, n54717, n54718, n54719, n54720, n54721, n54722, n54723,
         n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731,
         n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739,
         n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747,
         n54748, n54749, n54750, n54751, n54752, n54753, n54754, n54755,
         n54756, n54757, n54758, n54759, n54760, n54761, n54762, n54763,
         n54764, n54765, n54766, n54767, n54768, n54769, n54770, n54771,
         n54772, n54773, n54774, n54775, n54776, n54777, n54778, n54779,
         n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787,
         n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795,
         n54796, n54797, n54798, n54799, n54800, n54801, n54802, n54803,
         n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811,
         n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819,
         n54820, n54821, n54822, n54823, n54824, n54825, n54826, n54827,
         n54828, n54829, n54830, n54831, n54832, n54833, n54834, n54835,
         n54836, n54837, n54838, n54839, n54840, n54841, n54842, n54843,
         n54844, n54845, n54846, n54847, n54848, n54849, n54850, n54851,
         n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54859,
         n54860, n54861, n54862, n54863, n54864, n54865, n54866, n54867,
         n54868, n54869, n54870, n54871, n54872, n54873, n54874, n54875,
         n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883,
         n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891,
         n54892, n54893, n54894, n54895, n54896, n54897, n54898, n54899,
         n54900, n54901, n54902, n54903, n54904, n54905, n54906, n54907,
         n54908, n54909, n54910, n54911, n54912, n54913, n54914, n54915,
         n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923,
         n54924, n54925, n54926, n54927, n54928, n54929, n54930, n54931,
         n54932, n54933, n54934, n54935, n54936, n54937, n54938, n54939,
         n54940, n54941, n54942, n54943, n54944, n54945, n54946, n54947,
         n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955,
         n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963,
         n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971,
         n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979,
         n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987,
         n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995,
         n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003,
         n55004, n55005, n55006, n55007, n55008, n55009, n55010, n55011,
         n55012, n55013, n55014, n55015, n55016, n55017, n55018, n55019,
         n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027,
         n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035,
         n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043,
         n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051,
         n55052, n55053, n55054, n55055, n55056, n55057, n55058, n55059,
         n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067,
         n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075,
         n55076, n55077, n55078, n55079, n55080, n55081, n55082, n55083,
         n55084, n55085, n55086, n55087, n55088, n55089, n55090, n55091,
         n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099,
         n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107,
         n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115,
         n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123,
         n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131,
         n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139,
         n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147,
         n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155,
         n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163,
         n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171,
         n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179,
         n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187,
         n55188, n55189, n55190, n55191, n55192, n55193, n55194, n55195,
         n55196, n55197, n55198, n55199, n55200, n55201, n55202, n55203,
         n55204, n55205, n55206, n55207, n55208, n55209, n55210, n55211,
         n55212, n55213, n55214, n55215, n55216, n55217, n55218, n55219,
         n55220, n55221, n55222, n55223, n55224, n55225, n55226, n55227,
         n55228, n55229, n55230, n55231, n55232, n55233, n55234, n55235,
         n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243,
         n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251,
         n55252, n55253, n55254, n55255, n55256, n55257, n55258, n55259,
         n55260, n55261, n55262, n55263, n55264, n55265, n55266, n55267,
         n55268, n55269, n55270, n55271, n55272, n55273, n55274, n55275,
         n55276, n55277, n55278, n55279, n55280, n55281, n55282, n55283,
         n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291,
         n55292, n55293, n55294, n55295, n55296, n55297, n55298, n55299,
         n55300, n55301, n55302, n55303, n55304, n55305, n55306, n55307,
         n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315,
         n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323,
         n55324, n55325, n55326, n55327, n55328, n55329, n55330, n55331,
         n55332, n55333, n55334, n55335, n55336, n55337, n55338, n55339,
         n55340, n55341, n55342, n55343, n55344, n55345, n55346, n55347,
         n55348, n55349, n55350, n55351, n55352, n55353, n55354, n55355,
         n55356, n55357, n55358, n55359, n55360, n55361, n55362, n55363,
         n55364, n55365, n55366, n55367, n55368, n55369, n55370, n55371,
         n55372, n55373, n55374, n55375, n55376, n55377, n55378, n55379,
         n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387,
         n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395,
         n55396, n55397, n55398, n55399, n55400, n55401, n55402, n55403,
         n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411,
         n55412, n55413, n55414, n55415, n55416, n55417, n55418, n55419,
         n55420, n55421, n55422, n55423, n55424, n55425, n55426, n55427,
         n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435,
         n55436, n55437, n55438, n55439, n55440, n55441, n55442, n55443,
         n55444, n55445, n55446, n55447, n55448, n55449, n55450, n55451,
         n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459,
         n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467,
         n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475,
         n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483,
         n55484, n55485, n55486, n55487, n55488, n55489, n55490, n55491,
         n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499,
         n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507,
         n55508, n55509, n55510, n55511, n55512, n55513, n55514, n55515,
         n55516, n55517, n55518, n55519, n55520, n55521, n55522, n55523,
         n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531,
         n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539,
         n55540, n55541, n55542, n55543, n55544, n55545, n55546, n55547,
         n55548, n55549, n55550, n55551, n55552, n55553, n55554, n55555,
         n55556, n55557, n55558, n55559, n55560, n55561, n55562, n55563,
         n55564, n55565, n55566, n55567, n55568, n55569, n55570, n55571,
         n55572, n55573, n55574, n55575, n55576, n55577, n55578, n55579,
         n55580, n55581, n55582, n55583, n55584, n55585, n55586, n55587,
         n55588, n55589, n55590, n55591, n55592, n55593, n55594, n55595,
         n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603,
         n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611,
         n55612, n55613, n55614, n55615, n55616, n55617, n55618, n55619,
         n55620, n55621, n55622, n55623, n55624, n55625, n55626, n55627,
         n55628, n55629, n55630, n55631, n55632, n55633, n55634, n55635,
         n55636, n55637, n55638, n55639, n55640, n55641, n55642, n55643,
         n55644, n55645, n55646, n55647, n55648, n55649, n55650, n55651,
         n55652, n55653, n55654, n55655, n55656, n55657, n55658, n55659,
         n55660, n55661, n55662, n55663, n55664, n55665, n55666, n55667,
         n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675,
         n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683,
         n55684, n55685, n55686, n55687, n55688, n55689, n55690, n55691,
         n55692, n55693, n55694, n55695, n55696, n55697, n55698, n55699,
         n55700, n55701, n55702, n55703, n55704, n55705, n55706, n55707,
         n55708, n55709, n55710, n55711, n55712, n55713, n55714, n55715,
         n55716, n55717, n55718, n55719, n55720, n55721, n55722, n55723,
         n55724, n55725, n55726, n55727, n55728, n55729, n55730, n55731,
         n55732, n55733, n55734, n55735, n55736, n55737, n55738, n55739,
         n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747,
         n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755,
         n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763,
         n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771,
         n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779,
         n55780, n55781, n55782, n55783, n55784, n55785, n55786, n55787,
         n55788, n55789, n55790, n55791, n55792, n55793, n55794, n55795,
         n55796, n55797, n55798, n55799, n55800, n55801, n55802, n55803,
         n55804, n55805, n55806, n55807, n55808, n55809, n55810, n55811,
         n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819,
         n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827,
         n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835,
         n55836, n55837, n55838, n55839, n55840, n55841, n55842, n55843,
         n55844, n55845, n55846, n55847, n55848, n55849, n55850, n55851,
         n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859,
         n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867,
         n55868, n55869, n55870, n55871, n55872, n55873, n55874, n55875,
         n55876, n55877, n55878, n55879, n55880, n55881, n55882, n55883,
         n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891,
         n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899,
         n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55907,
         n55908, n55909, n55910, n55911, n55912, n55913, n55914, n55915,
         n55916, n55917, n55918, n55919, n55920, n55921, n55922, n55923,
         n55924, n55925, n55926, n55927, n55928, n55929, n55930, n55931,
         n55932, n55933, n55934, n55935, n55936, n55937, n55938, n55939,
         n55940, n55941, n55942, n55943, n55944, n55945, n55946, n55947,
         n55948, n55949, n55950, n55951, n55952, n55953, n55954, n55955,
         n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963,
         n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971,
         n55972, n55973, n55974, n55975, n55976, n55977, n55978, n55979,
         n55980, n55981, n55982, n55983, n55984, n55985, n55986, n55987,
         n55988, n55989, n55990, n55991, n55992, n55993, n55994, n55995,
         n55996, n55997, n55998, n55999, n56000, n56001, n56002, n56003,
         n56004, n56005, n56006, n56007, n56008, n56009, n56010, n56011,
         n56012, n56013, n56014, n56015, n56016, n56017, n56018, n56019,
         n56020, n56021, n56022, n56023, n56024, n56025, n56026, n56027,
         n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035,
         n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043,
         n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051,
         n56052, n56053, n56054, n56055, n56056, n56057, n56058, n56059,
         n56060, n56061, n56062, n56063, n56064, n56065, n56066, n56067,
         n56068, n56069, n56070, n56071, n56072, n56073, n56074, n56075,
         n56076, n56077, n56078, n56079, n56080, n56081, n56082, n56083,
         n56084, n56085, n56086, n56087, n56088, n56089, n56090, n56091,
         n56092, n56093, n56094, n56095, n56096, n56097, n56098, n56099,
         n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107,
         n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115,
         n56116, n56117, n56118, n56119, n56120, n56121, n56122, n56123,
         n56124, n56125, n56126, n56127, n56128, n56129, n56130, n56131,
         n56132, n56133, n56134, n56135, n56136, n56137, n56138, n56139,
         n56140, n56141, n56142, n56143, n56144, n56145, n56146, n56147,
         n56148, n56149, n56150, n56151, n56152, n56153, n56154, n56155,
         n56156, n56157, n56158, n56159, n56160, n56161, n56162, n56163,
         n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171,
         n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179,
         n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187,
         n56188, n56189, n56190, n56191, n56192, n56193, n56194, n56195,
         n56196, n56197, n56198, n56199, n56200, n56201, n56202, n56203,
         n56204, n56205, n56206, n56207, n56208, n56209, n56210, n56211,
         n56212, n56213, n56214, n56215, n56216, n56217, n56218, n56219,
         n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227,
         n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235,
         n56236, n56237, n56238, n56239, n56240, n56241, n56242, n56243,
         n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251,
         n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259,
         n56260, n56261, n56262, n56263, n56264, n56265, n56266, n56267,
         n56268, n56269, n56270, n56271, n56272, n56273, n56274, n56275,
         n56276, n56277, n56278, n56279, n56280, n56281, n56282, n56283,
         n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291,
         n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299,
         n56300, n56301, n56302, n56303, n56304, n56305, n56306, n56307,
         n56308, n56309, n56310, n56311, n56312, n56313, n56314, n56315,
         n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323,
         n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331,
         n56332, n56333, n56334, n56335, n56336, n56337, n56338, n56339,
         n56340, n56341, n56342, n56343, n56344, n56345, n56346, n56347,
         n56348, n56349, n56350, n56351, n56352, n56353, n56354, n56355,
         n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363,
         n56364, n56365, n56366, n56367, n56368, n56369, n56370, n56371,
         n56372, n56373, n56374, n56375, n56376, n56377, n56378, n56379,
         n56380, n56381, n56382, n56383, n56384, n56385, n56386, n56387,
         n56388, n56389, n56390, n56391, n56392, n56393, n56394, n56395,
         n56396, n56397, n56398, n56399, n56400, n56401, n56402, n56403,
         n56404, n56405, n56406, n56407, n56408, n56409, n56410, n56411,
         n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419,
         n56420, n56421, n56422, n56423, n56424, n56425, n56426, n56427,
         n56428, n56429, n56430, n56431, n56432, n56433, n56434, n56435,
         n56436, n56437, n56438, n56439, n56440, n56441, n56442, n56443,
         n56444, n56445, n56446, n56447, n56448, n56449, n56450, n56451,
         n56452, n56453, n56454, n56455, n56456, n56457, n56458, n56459,
         n56460, n56461, n56462, n56463, n56464, n56465, n56466, n56467,
         n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475,
         n56476, n56477, n56478, n56479, n56480, n56481, n56482, n56483,
         n56484, n56485, n56486, n56487, n56488, n56489, n56490, n56491,
         n56492, n56493, n56494, n56495, n56496, n56497, n56498, n56499,
         n56500, n56501, n56502, n56503, n56504, n56505, n56506, n56507,
         n56508, n56509, n56510, n56511, n56512, n56513, n56514, n56515,
         n56516, n56517, n56518, n56519, n56520, n56521, n56522, n56523,
         n56524, n56525, n56526, n56527, n56528, n56529, n56530, n56531,
         n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539,
         n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547,
         n56548, n56549, n56550, n56551, n56552, n56553, n56554, n56555,
         n56556, n56557, n56558, n56559, n56560, n56561, n56562, n56563,
         n56564, n56565, n56566, n56567, n56568, n56569, n56570, n56571,
         n56572, n56573, n56574, n56575, n56576, n56577, n56578, n56579,
         n56580, n56581, n56582, n56583, n56584, n56585, n56586, n56587,
         n56588, n56589, n56590, n56591, n56592, n56593, n56594, n56595,
         n56596, n56597, n56598, n56599, n56600, n56601, n56602, n56603,
         n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611,
         n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619,
         n56620, n56621, n56622, n56623, n56624, n56625, n56626, n56627,
         n56628, n56629, n56630, n56631, n56632, n56633, n56634, n56635,
         n56636, n56637, n56638, n56639, n56640, n56641, n56642, n56643,
         n56644, n56645, n56646, n56647, n56648, n56649, n56650, n56651,
         n56652, n56653, n56654, n56655, n56656, n56657, n56658, n56659,
         n56660, n56661, n56662, n56663, n56664, n56665, n56666, n56667,
         n56668, n56669, n56670, n56671, n56672, n56673, n56674, n56675,
         n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683,
         n56684, n56685, n56686, n56687, n56688, n56689, n56690, n56691,
         n56692, n56693, n56694, n56695, n56696, n56697, n56698, n56699,
         n56700, n56701, n56702, n56703, n56704, n56705, n56706, n56707,
         n56708, n56709, n56710, n56711, n56712, n56713, n56714, n56715,
         n56716, n56717, n56718, n56719, n56720, n56721, n56722, n56723,
         n56724, n56725, n56726, n56727, n56728, n56729, n56730, n56731,
         n56732, n56733, n56734, n56735, n56736, n56737, n56738, n56739,
         n56740, n56741, n56742, n56743, n56744, n56745, n56746, n56747,
         n56748, n56749, n56750, n56751, n56752, n56753, n56754, n56755,
         n56756, n56757, n56758, n56759, n56760, n56761, n56762, n56763,
         n56764, n56765, n56766, n56767, n56768, n56769, n56770, n56771,
         n56772, n56773, n56774, n56775, n56776, n56777, n56778, n56779,
         n56780, n56781, n56782, n56783, n56784, n56785, n56786, n56787,
         n56788, n56789, n56790, n56791, n56792, n56793, n56794, n56795,
         n56796, n56797, n56798, n56799, n56800, n56801, n56802, n56803,
         n56804, n56805, n56806, n56807, n56808, n56809, n56810, n56811,
         n56812, n56813, n56814, n56815, n56816, n56817, n56818, n56819,
         n56820, n56821, n56822, n56823, n56824, n56825, n56826, n56827,
         n56828, n56829, n56830, n56831, n56832, n56833, n56834, n56835,
         n56836, n56837, n56838, n56839, n56840, n56841, n56842, n56843,
         n56844, n56845, n56846, n56847, n56848, n56849, n56850, n56851,
         n56852, n56853, n56854, n56855, n56856, n56857, n56858, n56859,
         n56860, n56861, n56862, n56863, n56864, n56865, n56866, n56867,
         n56868, n56869, n56870, n56871, n56872, n56873, n56874, n56875,
         n56876, n56877, n56878, n56879, n56880, n56881, n56882, n56883,
         n56884, n56885, n56886, n56887, n56888, n56889, n56890, n56891,
         n56892, n56893, n56894, n56895, n56896, n56897, n56898, n56899,
         n56900, n56901, n56902, n56903, n56904, n56905, n56906, n56907,
         n56908, n56909, n56910, n56911, n56912, n56913, n56914, n56915,
         n56916, n56917, n56918, n56919, n56920, n56921, n56922, n56923,
         n56924, n56925, n56926, n56927, n56928, n56929, n56930, n56931,
         n56932, n56933, n56934, n56935, n56936, n56937, n56938, n56939,
         n56940, n56941, n56942, n56943, n56944, n56945, n56946, n56947,
         n56948, n56949, n56950, n56951, n56952, n56953, n56954, n56955,
         n56956, n56957, n56958, n56959, n56960, n56961, n56962, n56963,
         n56964, n56965, n56966, n56967, n56968, n56969, n56970, n56971,
         n56972, n56973, n56974, n56975, n56976, n56977, n56978, n56979,
         n56980, n56981, n56982, n56983, n56984, n56985, n56986, n56987,
         n56988, n56989, n56990, n56991, n56992, n56993, n56994, n56995,
         n56996, n56997, n56998, n56999, n57000, n57001, n57002, n57003,
         n57004, n57005, n57006, n57007, n57008, n57009, n57010, n57011,
         n57012, n57013, n57014, n57015, n57016, n57017, n57018, n57019,
         n57020, n57021, n57022, n57023, n57024, n57025, n57026, n57027,
         n57028, n57029, n57030, n57031, n57032, n57033, n57034, n57035,
         n57036, n57037, n57038, n57039, n57040, n57041, n57042, n57043,
         n57044, n57045, n57046, n57047, n57048, n57049, n57050, n57051,
         n57052, n57053, n57054, n57055, n57056, n57057, n57058, n57059,
         n57060, n57061, n57062, n57063, n57064, n57065, n57066, n57067,
         n57068, n57069, n57070, n57071, n57072, n57073, n57074, n57075,
         n57076, n57077, n57078, n57079, n57080, n57081, n57082, n57083,
         n57084, n57085, n57086, n57087, n57088, n57089, n57090, n57091,
         n57092, n57093, n57094, n57095, n57096, n57097, n57098, n57099,
         n57100, n57101, n57102, n57103, n57104, n57105, n57106, n57107,
         n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115,
         n57116, n57117, n57118, n57119, n57120, n57121, n57122, n57123,
         n57124, n57125, n57126, n57127, n57128, n57129, n57130, n57131,
         n57132, n57133, n57134, n57135, n57136, n57137, n57138, n57139,
         n57140, n57141, n57142, n57143, n57144, n57145, n57146, n57147,
         n57148, n57149, n57150, n57151, n57152, n57153, n57154, n57155,
         n57156, n57157, n57158, n57159, n57160, n57161, n57162, n57163,
         n57164, n57165, n57166, n57167, n57168, n57169, n57170, n57171,
         n57172, n57173, n57174, n57175, n57176, n57177, n57178, n57179,
         n57180, n57181, n57182, n57183, n57184, n57185, n57186, n57187,
         n57188, n57189, n57190, n57191, n57192, n57193, n57194, n57195,
         n57196, n57197, n57198, n57199, n57200, n57201, n57202, n57203,
         n57204, n57205, n57206, n57207, n57208, n57209, n57210, n57211,
         n57212, n57213, n57214, n57215, n57216, n57217, n57218, n57219,
         n57220, n57221, n57222, n57223, n57224, n57225, n57226, n57227,
         n57228, n57229, n57230, n57231, n57232, n57233, n57234, n57235,
         n57236, n57237, n57238, n57239, n57240, n57241, n57242, n57243,
         n57244, n57245, n57246, n57247, n57248, n57249, n57250, n57251,
         n57252, n57253, n57254, n57255, n57256, n57257, n57258, n57259,
         n57260, n57261, n57262, n57263, n57264, n57265, n57266, n57267,
         n57268, n57269, n57270, n57271, n57272, n57273, n57274, n57275,
         n57276, n57277, n57278, n57279, n57280, n57281, n57282, n57283,
         n57284, n57285, n57286, n57287, n57288, n57289, n57290, n57291,
         n57292, n57293, n57294, n57295, n57296, n57297, n57298, n57299,
         n57300, n57301, n57302, n57303, n57304, n57305, n57306, n57307,
         n57308, n57309, n57310, n57311, n57312, n57313, n57314, n57315,
         n57316, n57317, n57318, n57319, n57320, n57321, n57322, n57323,
         n57324, n57325, n57326, n57327, n57328, n57329, n57330, n57331,
         n57332, n57333, n57334, n57335, n57336, n57337, n57338, n57339,
         n57340, n57341, n57342, n57343, n57344, n57345, n57346, n57347,
         n57348, n57349, n57350, n57351, n57352, n57353, n57354, n57355,
         n57356, n57357, n57358, n57359, n57360, n57361, n57362, n57363,
         n57364, n57365, n57366, n57367, n57368, n57369, n57370, n57371,
         n57372, n57373, n57374, n57375, n57376, n57377, n57378, n57379,
         n57380, n57381, n57382, n57383, n57384, n57385, n57386, n57387,
         n57388, n57389, n57390, n57391, n57392, n57393, n57394, n57395,
         n57396, n57397, n57398, n57399, n57400, n57401, n57402, n57403,
         n57404, n57405, n57406, n57407, n57408, n57409, n57410, n57411,
         n57412, n57413, n57414, n57415, n57416, n57417, n57418, n57419,
         n57420, n57421, n57422, n57423, n57424, n57425, n57426, n57427,
         n57428, n57429, n57430, n57431, n57432, n57433, n57434, n57435,
         n57436, n57437, n57438, n57439, n57440, n57441, n57442, n57443,
         n57444, n57445, n57446, n57447, n57448, n57449, n57450, n57451,
         n57452, n57453, n57454, n57455, n57456, n57457, n57458, n57459,
         n57460, n57461, n57462, n57463, n57464, n57465, n57466, n57467,
         n57468, n57469, n57470, n57471, n57472, n57473, n57474, n57475,
         n57476, n57477, n57478, n57479, n57480, n57481, n57482, n57483,
         n57484, n57485, n57486, n57487, n57488, n57489, n57490, n57491,
         n57492, n57493, n57494, n57495, n57496, n57497, n57498, n57499,
         n57500, n57501, n57502, n57503, n57504, n57505, n57506, n57507,
         n57508, n57509, n57510, n57511, n57512, n57513, n57514, n57515,
         n57516, n57517, n57518, n57519, n57520, n57521, n57522, n57523,
         n57524, n57525, n57526, n57527, n57528, n57529, n57530, n57531,
         n57532, n57533, n57534, n57535, n57536, n57537, n57538, n57539,
         n57540, n57541, n57542, n57543, n57544, n57545, n57546, n57547,
         n57548, n57549, n57550, n57551, n57552, n57553, n57554, n57555,
         n57556, n57557, n57558, n57559, n57560, n57561, n57562, n57563,
         n57564, n57565, n57566, n57567, n57568, n57569, n57570, n57571,
         n57572, n57573;
  assign \knn_comb_/min_val_out[0][0]  = p_input[2032];
  assign \knn_comb_/min_val_out[0][1]  = p_input[2033];
  assign \knn_comb_/min_val_out[0][2]  = p_input[2034];
  assign \knn_comb_/min_val_out[0][3]  = p_input[2035];
  assign \knn_comb_/min_val_out[0][4]  = p_input[2036];
  assign \knn_comb_/min_val_out[0][5]  = p_input[2037];
  assign \knn_comb_/min_val_out[0][6]  = p_input[2038];
  assign \knn_comb_/min_val_out[0][7]  = p_input[2039];
  assign \knn_comb_/min_val_out[0][8]  = p_input[2040];
  assign \knn_comb_/min_val_out[0][9]  = p_input[2041];
  assign \knn_comb_/min_val_out[0][10]  = p_input[2042];
  assign \knn_comb_/min_val_out[0][11]  = p_input[2043];
  assign \knn_comb_/min_val_out[0][12]  = p_input[2044];
  assign \knn_comb_/min_val_out[0][13]  = p_input[2045];
  assign \knn_comb_/min_val_out[0][14]  = p_input[2046];
  assign \knn_comb_/min_val_out[0][15]  = p_input[2047];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[2000];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[2001];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[2002];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[2003];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[2004];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[2005];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[2006];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[2007];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[2008];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[2009];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[2010];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[2011];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[2012];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[2013];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[2014];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[2015];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[2016];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[2017];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[2018];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[2019];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[2020];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[2021];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[2022];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[2023];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[2024];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[2025];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[2026];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[2027];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[2028];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[2029];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[2030];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[2031];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[47]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[46]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[45]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[44]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[43]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[42]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[41]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[40]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[3]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[39]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[38]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[37]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[36]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[35]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[34]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[33]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[32]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[31]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[30]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[2]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[29]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[28]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[27]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[26]) );
  XOR U31 ( .A(n1), .B(n61), .Z(o[25]) );
  AND U32 ( .A(n62), .B(n63), .Z(n1) );
  XOR U33 ( .A(n2), .B(n61), .Z(n63) );
  XOR U34 ( .A(n64), .B(n25), .Z(n61) );
  AND U35 ( .A(n65), .B(n66), .Z(n25) );
  XNOR U36 ( .A(n67), .B(n26), .Z(n66) );
  XOR U37 ( .A(n68), .B(n69), .Z(n26) );
  AND U38 ( .A(n70), .B(n71), .Z(n69) );
  XOR U39 ( .A(p_input[9]), .B(n68), .Z(n71) );
  XOR U40 ( .A(n72), .B(n73), .Z(n68) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  IV U42 ( .A(n64), .Z(n67) );
  XOR U43 ( .A(n76), .B(n77), .Z(n64) );
  AND U44 ( .A(n78), .B(n79), .Z(n77) );
  XOR U45 ( .A(n80), .B(n81), .Z(n2) );
  AND U46 ( .A(n82), .B(n79), .Z(n81) );
  XNOR U47 ( .A(n83), .B(n76), .Z(n79) );
  XOR U48 ( .A(n84), .B(n85), .Z(n76) );
  AND U49 ( .A(n86), .B(n75), .Z(n85) );
  XNOR U50 ( .A(n87), .B(n72), .Z(n75) );
  XOR U51 ( .A(n88), .B(n89), .Z(n72) );
  AND U52 ( .A(n90), .B(n91), .Z(n89) );
  XOR U53 ( .A(p_input[25]), .B(n88), .Z(n91) );
  XOR U54 ( .A(n92), .B(n93), .Z(n88) );
  AND U55 ( .A(n94), .B(n95), .Z(n93) );
  IV U56 ( .A(n84), .Z(n87) );
  XOR U57 ( .A(n96), .B(n97), .Z(n84) );
  AND U58 ( .A(n98), .B(n99), .Z(n97) );
  IV U59 ( .A(n80), .Z(n83) );
  XNOR U60 ( .A(n100), .B(n101), .Z(n80) );
  AND U61 ( .A(n102), .B(n99), .Z(n101) );
  XNOR U62 ( .A(n100), .B(n96), .Z(n99) );
  XOR U63 ( .A(n103), .B(n104), .Z(n96) );
  AND U64 ( .A(n105), .B(n95), .Z(n104) );
  XNOR U65 ( .A(n106), .B(n92), .Z(n95) );
  XOR U66 ( .A(n107), .B(n108), .Z(n92) );
  AND U67 ( .A(n109), .B(n110), .Z(n108) );
  XOR U68 ( .A(p_input[41]), .B(n107), .Z(n110) );
  XOR U69 ( .A(n111), .B(n112), .Z(n107) );
  AND U70 ( .A(n113), .B(n114), .Z(n112) );
  IV U71 ( .A(n103), .Z(n106) );
  XOR U72 ( .A(n115), .B(n116), .Z(n103) );
  AND U73 ( .A(n117), .B(n118), .Z(n116) );
  XOR U74 ( .A(n119), .B(n120), .Z(n100) );
  AND U75 ( .A(n121), .B(n118), .Z(n120) );
  XNOR U76 ( .A(n119), .B(n115), .Z(n118) );
  XOR U77 ( .A(n122), .B(n123), .Z(n115) );
  AND U78 ( .A(n124), .B(n114), .Z(n123) );
  XNOR U79 ( .A(n125), .B(n111), .Z(n114) );
  XOR U80 ( .A(n126), .B(n127), .Z(n111) );
  AND U81 ( .A(n128), .B(n129), .Z(n127) );
  XOR U82 ( .A(p_input[57]), .B(n126), .Z(n129) );
  XOR U83 ( .A(n130), .B(n131), .Z(n126) );
  AND U84 ( .A(n132), .B(n133), .Z(n131) );
  IV U85 ( .A(n122), .Z(n125) );
  XOR U86 ( .A(n134), .B(n135), .Z(n122) );
  AND U87 ( .A(n136), .B(n137), .Z(n135) );
  XOR U88 ( .A(n138), .B(n139), .Z(n119) );
  AND U89 ( .A(n140), .B(n137), .Z(n139) );
  XNOR U90 ( .A(n138), .B(n134), .Z(n137) );
  XOR U91 ( .A(n141), .B(n142), .Z(n134) );
  AND U92 ( .A(n143), .B(n133), .Z(n142) );
  XNOR U93 ( .A(n144), .B(n130), .Z(n133) );
  XOR U94 ( .A(n145), .B(n146), .Z(n130) );
  AND U95 ( .A(n147), .B(n148), .Z(n146) );
  XOR U96 ( .A(p_input[73]), .B(n145), .Z(n148) );
  XOR U97 ( .A(n149), .B(n150), .Z(n145) );
  AND U98 ( .A(n151), .B(n152), .Z(n150) );
  IV U99 ( .A(n141), .Z(n144) );
  XOR U100 ( .A(n153), .B(n154), .Z(n141) );
  AND U101 ( .A(n155), .B(n156), .Z(n154) );
  XOR U102 ( .A(n157), .B(n158), .Z(n138) );
  AND U103 ( .A(n159), .B(n156), .Z(n158) );
  XNOR U104 ( .A(n157), .B(n153), .Z(n156) );
  XOR U105 ( .A(n160), .B(n161), .Z(n153) );
  AND U106 ( .A(n162), .B(n152), .Z(n161) );
  XNOR U107 ( .A(n163), .B(n149), .Z(n152) );
  XOR U108 ( .A(n164), .B(n165), .Z(n149) );
  AND U109 ( .A(n166), .B(n167), .Z(n165) );
  XOR U110 ( .A(p_input[89]), .B(n164), .Z(n167) );
  XOR U111 ( .A(n168), .B(n169), .Z(n164) );
  AND U112 ( .A(n170), .B(n171), .Z(n169) );
  IV U113 ( .A(n160), .Z(n163) );
  XOR U114 ( .A(n172), .B(n173), .Z(n160) );
  AND U115 ( .A(n174), .B(n175), .Z(n173) );
  XOR U116 ( .A(n176), .B(n177), .Z(n157) );
  AND U117 ( .A(n178), .B(n175), .Z(n177) );
  XNOR U118 ( .A(n176), .B(n172), .Z(n175) );
  XOR U119 ( .A(n179), .B(n180), .Z(n172) );
  AND U120 ( .A(n181), .B(n171), .Z(n180) );
  XNOR U121 ( .A(n182), .B(n168), .Z(n171) );
  XOR U122 ( .A(n183), .B(n184), .Z(n168) );
  AND U123 ( .A(n185), .B(n186), .Z(n184) );
  XOR U124 ( .A(p_input[105]), .B(n183), .Z(n186) );
  XOR U125 ( .A(n187), .B(n188), .Z(n183) );
  AND U126 ( .A(n189), .B(n190), .Z(n188) );
  IV U127 ( .A(n179), .Z(n182) );
  XOR U128 ( .A(n191), .B(n192), .Z(n179) );
  AND U129 ( .A(n193), .B(n194), .Z(n192) );
  XOR U130 ( .A(n195), .B(n196), .Z(n176) );
  AND U131 ( .A(n197), .B(n194), .Z(n196) );
  XNOR U132 ( .A(n195), .B(n191), .Z(n194) );
  XOR U133 ( .A(n198), .B(n199), .Z(n191) );
  AND U134 ( .A(n200), .B(n190), .Z(n199) );
  XNOR U135 ( .A(n201), .B(n187), .Z(n190) );
  XOR U136 ( .A(n202), .B(n203), .Z(n187) );
  AND U137 ( .A(n204), .B(n205), .Z(n203) );
  XOR U138 ( .A(p_input[121]), .B(n202), .Z(n205) );
  XOR U139 ( .A(n206), .B(n207), .Z(n202) );
  AND U140 ( .A(n208), .B(n209), .Z(n207) );
  IV U141 ( .A(n198), .Z(n201) );
  XOR U142 ( .A(n210), .B(n211), .Z(n198) );
  AND U143 ( .A(n212), .B(n213), .Z(n211) );
  XOR U144 ( .A(n214), .B(n215), .Z(n195) );
  AND U145 ( .A(n216), .B(n213), .Z(n215) );
  XNOR U146 ( .A(n214), .B(n210), .Z(n213) );
  XOR U147 ( .A(n217), .B(n218), .Z(n210) );
  AND U148 ( .A(n219), .B(n209), .Z(n218) );
  XNOR U149 ( .A(n220), .B(n206), .Z(n209) );
  XOR U150 ( .A(n221), .B(n222), .Z(n206) );
  AND U151 ( .A(n223), .B(n224), .Z(n222) );
  XOR U152 ( .A(p_input[137]), .B(n221), .Z(n224) );
  XOR U153 ( .A(n225), .B(n226), .Z(n221) );
  AND U154 ( .A(n227), .B(n228), .Z(n226) );
  IV U155 ( .A(n217), .Z(n220) );
  XOR U156 ( .A(n229), .B(n230), .Z(n217) );
  AND U157 ( .A(n231), .B(n232), .Z(n230) );
  XOR U158 ( .A(n233), .B(n234), .Z(n214) );
  AND U159 ( .A(n235), .B(n232), .Z(n234) );
  XNOR U160 ( .A(n233), .B(n229), .Z(n232) );
  XOR U161 ( .A(n236), .B(n237), .Z(n229) );
  AND U162 ( .A(n238), .B(n228), .Z(n237) );
  XNOR U163 ( .A(n239), .B(n225), .Z(n228) );
  XOR U164 ( .A(n240), .B(n241), .Z(n225) );
  AND U165 ( .A(n242), .B(n243), .Z(n241) );
  XOR U166 ( .A(p_input[153]), .B(n240), .Z(n243) );
  XOR U167 ( .A(n244), .B(n245), .Z(n240) );
  AND U168 ( .A(n246), .B(n247), .Z(n245) );
  IV U169 ( .A(n236), .Z(n239) );
  XOR U170 ( .A(n248), .B(n249), .Z(n236) );
  AND U171 ( .A(n250), .B(n251), .Z(n249) );
  XOR U172 ( .A(n252), .B(n253), .Z(n233) );
  AND U173 ( .A(n254), .B(n251), .Z(n253) );
  XNOR U174 ( .A(n252), .B(n248), .Z(n251) );
  XOR U175 ( .A(n255), .B(n256), .Z(n248) );
  AND U176 ( .A(n257), .B(n247), .Z(n256) );
  XNOR U177 ( .A(n258), .B(n244), .Z(n247) );
  XOR U178 ( .A(n259), .B(n260), .Z(n244) );
  AND U179 ( .A(n261), .B(n262), .Z(n260) );
  XOR U180 ( .A(p_input[169]), .B(n259), .Z(n262) );
  XOR U181 ( .A(n263), .B(n264), .Z(n259) );
  AND U182 ( .A(n265), .B(n266), .Z(n264) );
  IV U183 ( .A(n255), .Z(n258) );
  XOR U184 ( .A(n267), .B(n268), .Z(n255) );
  AND U185 ( .A(n269), .B(n270), .Z(n268) );
  XOR U186 ( .A(n271), .B(n272), .Z(n252) );
  AND U187 ( .A(n273), .B(n270), .Z(n272) );
  XNOR U188 ( .A(n271), .B(n267), .Z(n270) );
  XOR U189 ( .A(n274), .B(n275), .Z(n267) );
  AND U190 ( .A(n276), .B(n266), .Z(n275) );
  XNOR U191 ( .A(n277), .B(n263), .Z(n266) );
  XOR U192 ( .A(n278), .B(n279), .Z(n263) );
  AND U193 ( .A(n280), .B(n281), .Z(n279) );
  XOR U194 ( .A(p_input[185]), .B(n278), .Z(n281) );
  XOR U195 ( .A(n282), .B(n283), .Z(n278) );
  AND U196 ( .A(n284), .B(n285), .Z(n283) );
  IV U197 ( .A(n274), .Z(n277) );
  XOR U198 ( .A(n286), .B(n287), .Z(n274) );
  AND U199 ( .A(n288), .B(n289), .Z(n287) );
  XOR U200 ( .A(n290), .B(n291), .Z(n271) );
  AND U201 ( .A(n292), .B(n289), .Z(n291) );
  XNOR U202 ( .A(n290), .B(n286), .Z(n289) );
  XOR U203 ( .A(n293), .B(n294), .Z(n286) );
  AND U204 ( .A(n295), .B(n285), .Z(n294) );
  XNOR U205 ( .A(n296), .B(n282), .Z(n285) );
  XOR U206 ( .A(n297), .B(n298), .Z(n282) );
  AND U207 ( .A(n299), .B(n300), .Z(n298) );
  XOR U208 ( .A(p_input[201]), .B(n297), .Z(n300) );
  XOR U209 ( .A(n301), .B(n302), .Z(n297) );
  AND U210 ( .A(n303), .B(n304), .Z(n302) );
  IV U211 ( .A(n293), .Z(n296) );
  XOR U212 ( .A(n305), .B(n306), .Z(n293) );
  AND U213 ( .A(n307), .B(n308), .Z(n306) );
  XOR U214 ( .A(n309), .B(n310), .Z(n290) );
  AND U215 ( .A(n311), .B(n308), .Z(n310) );
  XNOR U216 ( .A(n309), .B(n305), .Z(n308) );
  XOR U217 ( .A(n312), .B(n313), .Z(n305) );
  AND U218 ( .A(n314), .B(n304), .Z(n313) );
  XNOR U219 ( .A(n315), .B(n301), .Z(n304) );
  XOR U220 ( .A(n316), .B(n317), .Z(n301) );
  AND U221 ( .A(n318), .B(n319), .Z(n317) );
  XOR U222 ( .A(p_input[217]), .B(n316), .Z(n319) );
  XOR U223 ( .A(n320), .B(n321), .Z(n316) );
  AND U224 ( .A(n322), .B(n323), .Z(n321) );
  IV U225 ( .A(n312), .Z(n315) );
  XOR U226 ( .A(n324), .B(n325), .Z(n312) );
  AND U227 ( .A(n326), .B(n327), .Z(n325) );
  XOR U228 ( .A(n328), .B(n329), .Z(n309) );
  AND U229 ( .A(n330), .B(n327), .Z(n329) );
  XNOR U230 ( .A(n328), .B(n324), .Z(n327) );
  XOR U231 ( .A(n331), .B(n332), .Z(n324) );
  AND U232 ( .A(n333), .B(n323), .Z(n332) );
  XNOR U233 ( .A(n334), .B(n320), .Z(n323) );
  XOR U234 ( .A(n335), .B(n336), .Z(n320) );
  AND U235 ( .A(n337), .B(n338), .Z(n336) );
  XOR U236 ( .A(p_input[233]), .B(n335), .Z(n338) );
  XOR U237 ( .A(n339), .B(n340), .Z(n335) );
  AND U238 ( .A(n341), .B(n342), .Z(n340) );
  IV U239 ( .A(n331), .Z(n334) );
  XOR U240 ( .A(n343), .B(n344), .Z(n331) );
  AND U241 ( .A(n345), .B(n346), .Z(n344) );
  XOR U242 ( .A(n347), .B(n348), .Z(n328) );
  AND U243 ( .A(n349), .B(n346), .Z(n348) );
  XNOR U244 ( .A(n347), .B(n343), .Z(n346) );
  XOR U245 ( .A(n350), .B(n351), .Z(n343) );
  AND U246 ( .A(n352), .B(n342), .Z(n351) );
  XNOR U247 ( .A(n353), .B(n339), .Z(n342) );
  XOR U248 ( .A(n354), .B(n355), .Z(n339) );
  AND U249 ( .A(n356), .B(n357), .Z(n355) );
  XOR U250 ( .A(p_input[249]), .B(n354), .Z(n357) );
  XOR U251 ( .A(n358), .B(n359), .Z(n354) );
  AND U252 ( .A(n360), .B(n361), .Z(n359) );
  IV U253 ( .A(n350), .Z(n353) );
  XOR U254 ( .A(n362), .B(n363), .Z(n350) );
  AND U255 ( .A(n364), .B(n365), .Z(n363) );
  XOR U256 ( .A(n366), .B(n367), .Z(n347) );
  AND U257 ( .A(n368), .B(n365), .Z(n367) );
  XNOR U258 ( .A(n366), .B(n362), .Z(n365) );
  XOR U259 ( .A(n369), .B(n370), .Z(n362) );
  AND U260 ( .A(n371), .B(n361), .Z(n370) );
  XNOR U261 ( .A(n372), .B(n358), .Z(n361) );
  XOR U262 ( .A(n373), .B(n374), .Z(n358) );
  AND U263 ( .A(n375), .B(n376), .Z(n374) );
  XOR U264 ( .A(p_input[265]), .B(n373), .Z(n376) );
  XOR U265 ( .A(n377), .B(n378), .Z(n373) );
  AND U266 ( .A(n379), .B(n380), .Z(n378) );
  IV U267 ( .A(n369), .Z(n372) );
  XOR U268 ( .A(n381), .B(n382), .Z(n369) );
  AND U269 ( .A(n383), .B(n384), .Z(n382) );
  XOR U270 ( .A(n385), .B(n386), .Z(n366) );
  AND U271 ( .A(n387), .B(n384), .Z(n386) );
  XNOR U272 ( .A(n385), .B(n381), .Z(n384) );
  XOR U273 ( .A(n388), .B(n389), .Z(n381) );
  AND U274 ( .A(n390), .B(n380), .Z(n389) );
  XNOR U275 ( .A(n391), .B(n377), .Z(n380) );
  XOR U276 ( .A(n392), .B(n393), .Z(n377) );
  AND U277 ( .A(n394), .B(n395), .Z(n393) );
  XOR U278 ( .A(p_input[281]), .B(n392), .Z(n395) );
  XOR U279 ( .A(n396), .B(n397), .Z(n392) );
  AND U280 ( .A(n398), .B(n399), .Z(n397) );
  IV U281 ( .A(n388), .Z(n391) );
  XOR U282 ( .A(n400), .B(n401), .Z(n388) );
  AND U283 ( .A(n402), .B(n403), .Z(n401) );
  XOR U284 ( .A(n404), .B(n405), .Z(n385) );
  AND U285 ( .A(n406), .B(n403), .Z(n405) );
  XNOR U286 ( .A(n404), .B(n400), .Z(n403) );
  XOR U287 ( .A(n407), .B(n408), .Z(n400) );
  AND U288 ( .A(n409), .B(n399), .Z(n408) );
  XNOR U289 ( .A(n410), .B(n396), .Z(n399) );
  XOR U290 ( .A(n411), .B(n412), .Z(n396) );
  AND U291 ( .A(n413), .B(n414), .Z(n412) );
  XOR U292 ( .A(p_input[297]), .B(n411), .Z(n414) );
  XOR U293 ( .A(n415), .B(n416), .Z(n411) );
  AND U294 ( .A(n417), .B(n418), .Z(n416) );
  IV U295 ( .A(n407), .Z(n410) );
  XOR U296 ( .A(n419), .B(n420), .Z(n407) );
  AND U297 ( .A(n421), .B(n422), .Z(n420) );
  XOR U298 ( .A(n423), .B(n424), .Z(n404) );
  AND U299 ( .A(n425), .B(n422), .Z(n424) );
  XNOR U300 ( .A(n423), .B(n419), .Z(n422) );
  XOR U301 ( .A(n426), .B(n427), .Z(n419) );
  AND U302 ( .A(n428), .B(n418), .Z(n427) );
  XNOR U303 ( .A(n429), .B(n415), .Z(n418) );
  XOR U304 ( .A(n430), .B(n431), .Z(n415) );
  AND U305 ( .A(n432), .B(n433), .Z(n431) );
  XOR U306 ( .A(p_input[313]), .B(n430), .Z(n433) );
  XOR U307 ( .A(n434), .B(n435), .Z(n430) );
  AND U308 ( .A(n436), .B(n437), .Z(n435) );
  IV U309 ( .A(n426), .Z(n429) );
  XOR U310 ( .A(n438), .B(n439), .Z(n426) );
  AND U311 ( .A(n440), .B(n441), .Z(n439) );
  XOR U312 ( .A(n442), .B(n443), .Z(n423) );
  AND U313 ( .A(n444), .B(n441), .Z(n443) );
  XNOR U314 ( .A(n442), .B(n438), .Z(n441) );
  XOR U315 ( .A(n445), .B(n446), .Z(n438) );
  AND U316 ( .A(n447), .B(n437), .Z(n446) );
  XNOR U317 ( .A(n448), .B(n434), .Z(n437) );
  XOR U318 ( .A(n449), .B(n450), .Z(n434) );
  AND U319 ( .A(n451), .B(n452), .Z(n450) );
  XOR U320 ( .A(p_input[329]), .B(n449), .Z(n452) );
  XOR U321 ( .A(n453), .B(n454), .Z(n449) );
  AND U322 ( .A(n455), .B(n456), .Z(n454) );
  IV U323 ( .A(n445), .Z(n448) );
  XOR U324 ( .A(n457), .B(n458), .Z(n445) );
  AND U325 ( .A(n459), .B(n460), .Z(n458) );
  XOR U326 ( .A(n461), .B(n462), .Z(n442) );
  AND U327 ( .A(n463), .B(n460), .Z(n462) );
  XNOR U328 ( .A(n461), .B(n457), .Z(n460) );
  XOR U329 ( .A(n464), .B(n465), .Z(n457) );
  AND U330 ( .A(n466), .B(n456), .Z(n465) );
  XNOR U331 ( .A(n467), .B(n453), .Z(n456) );
  XOR U332 ( .A(n468), .B(n469), .Z(n453) );
  AND U333 ( .A(n470), .B(n471), .Z(n469) );
  XOR U334 ( .A(p_input[345]), .B(n468), .Z(n471) );
  XOR U335 ( .A(n472), .B(n473), .Z(n468) );
  AND U336 ( .A(n474), .B(n475), .Z(n473) );
  IV U337 ( .A(n464), .Z(n467) );
  XOR U338 ( .A(n476), .B(n477), .Z(n464) );
  AND U339 ( .A(n478), .B(n479), .Z(n477) );
  XOR U340 ( .A(n480), .B(n481), .Z(n461) );
  AND U341 ( .A(n482), .B(n479), .Z(n481) );
  XNOR U342 ( .A(n480), .B(n476), .Z(n479) );
  XOR U343 ( .A(n483), .B(n484), .Z(n476) );
  AND U344 ( .A(n485), .B(n475), .Z(n484) );
  XNOR U345 ( .A(n486), .B(n472), .Z(n475) );
  XOR U346 ( .A(n487), .B(n488), .Z(n472) );
  AND U347 ( .A(n489), .B(n490), .Z(n488) );
  XOR U348 ( .A(p_input[361]), .B(n487), .Z(n490) );
  XOR U349 ( .A(n491), .B(n492), .Z(n487) );
  AND U350 ( .A(n493), .B(n494), .Z(n492) );
  IV U351 ( .A(n483), .Z(n486) );
  XOR U352 ( .A(n495), .B(n496), .Z(n483) );
  AND U353 ( .A(n497), .B(n498), .Z(n496) );
  XOR U354 ( .A(n499), .B(n500), .Z(n480) );
  AND U355 ( .A(n501), .B(n498), .Z(n500) );
  XNOR U356 ( .A(n499), .B(n495), .Z(n498) );
  XOR U357 ( .A(n502), .B(n503), .Z(n495) );
  AND U358 ( .A(n504), .B(n494), .Z(n503) );
  XNOR U359 ( .A(n505), .B(n491), .Z(n494) );
  XOR U360 ( .A(n506), .B(n507), .Z(n491) );
  AND U361 ( .A(n508), .B(n509), .Z(n507) );
  XOR U362 ( .A(p_input[377]), .B(n506), .Z(n509) );
  XOR U363 ( .A(n510), .B(n511), .Z(n506) );
  AND U364 ( .A(n512), .B(n513), .Z(n511) );
  IV U365 ( .A(n502), .Z(n505) );
  XOR U366 ( .A(n514), .B(n515), .Z(n502) );
  AND U367 ( .A(n516), .B(n517), .Z(n515) );
  XOR U368 ( .A(n518), .B(n519), .Z(n499) );
  AND U369 ( .A(n520), .B(n517), .Z(n519) );
  XNOR U370 ( .A(n518), .B(n514), .Z(n517) );
  XOR U371 ( .A(n521), .B(n522), .Z(n514) );
  AND U372 ( .A(n523), .B(n513), .Z(n522) );
  XNOR U373 ( .A(n524), .B(n510), .Z(n513) );
  XOR U374 ( .A(n525), .B(n526), .Z(n510) );
  AND U375 ( .A(n527), .B(n528), .Z(n526) );
  XOR U376 ( .A(p_input[393]), .B(n525), .Z(n528) );
  XOR U377 ( .A(n529), .B(n530), .Z(n525) );
  AND U378 ( .A(n531), .B(n532), .Z(n530) );
  IV U379 ( .A(n521), .Z(n524) );
  XOR U380 ( .A(n533), .B(n534), .Z(n521) );
  AND U381 ( .A(n535), .B(n536), .Z(n534) );
  XOR U382 ( .A(n537), .B(n538), .Z(n518) );
  AND U383 ( .A(n539), .B(n536), .Z(n538) );
  XNOR U384 ( .A(n537), .B(n533), .Z(n536) );
  XOR U385 ( .A(n540), .B(n541), .Z(n533) );
  AND U386 ( .A(n542), .B(n532), .Z(n541) );
  XNOR U387 ( .A(n543), .B(n529), .Z(n532) );
  XOR U388 ( .A(n544), .B(n545), .Z(n529) );
  AND U389 ( .A(n546), .B(n547), .Z(n545) );
  XOR U390 ( .A(p_input[409]), .B(n544), .Z(n547) );
  XOR U391 ( .A(n548), .B(n549), .Z(n544) );
  AND U392 ( .A(n550), .B(n551), .Z(n549) );
  IV U393 ( .A(n540), .Z(n543) );
  XOR U394 ( .A(n552), .B(n553), .Z(n540) );
  AND U395 ( .A(n554), .B(n555), .Z(n553) );
  XOR U396 ( .A(n556), .B(n557), .Z(n537) );
  AND U397 ( .A(n558), .B(n555), .Z(n557) );
  XNOR U398 ( .A(n556), .B(n552), .Z(n555) );
  XOR U399 ( .A(n559), .B(n560), .Z(n552) );
  AND U400 ( .A(n561), .B(n551), .Z(n560) );
  XNOR U401 ( .A(n562), .B(n548), .Z(n551) );
  XOR U402 ( .A(n563), .B(n564), .Z(n548) );
  AND U403 ( .A(n565), .B(n566), .Z(n564) );
  XOR U404 ( .A(p_input[425]), .B(n563), .Z(n566) );
  XOR U405 ( .A(n567), .B(n568), .Z(n563) );
  AND U406 ( .A(n569), .B(n570), .Z(n568) );
  IV U407 ( .A(n559), .Z(n562) );
  XOR U408 ( .A(n571), .B(n572), .Z(n559) );
  AND U409 ( .A(n573), .B(n574), .Z(n572) );
  XOR U410 ( .A(n575), .B(n576), .Z(n556) );
  AND U411 ( .A(n577), .B(n574), .Z(n576) );
  XNOR U412 ( .A(n575), .B(n571), .Z(n574) );
  XOR U413 ( .A(n578), .B(n579), .Z(n571) );
  AND U414 ( .A(n580), .B(n570), .Z(n579) );
  XNOR U415 ( .A(n581), .B(n567), .Z(n570) );
  XOR U416 ( .A(n582), .B(n583), .Z(n567) );
  AND U417 ( .A(n584), .B(n585), .Z(n583) );
  XOR U418 ( .A(p_input[441]), .B(n582), .Z(n585) );
  XOR U419 ( .A(n586), .B(n587), .Z(n582) );
  AND U420 ( .A(n588), .B(n589), .Z(n587) );
  IV U421 ( .A(n578), .Z(n581) );
  XOR U422 ( .A(n590), .B(n591), .Z(n578) );
  AND U423 ( .A(n592), .B(n593), .Z(n591) );
  XOR U424 ( .A(n594), .B(n595), .Z(n575) );
  AND U425 ( .A(n596), .B(n593), .Z(n595) );
  XNOR U426 ( .A(n594), .B(n590), .Z(n593) );
  XOR U427 ( .A(n597), .B(n598), .Z(n590) );
  AND U428 ( .A(n599), .B(n589), .Z(n598) );
  XNOR U429 ( .A(n600), .B(n586), .Z(n589) );
  XOR U430 ( .A(n601), .B(n602), .Z(n586) );
  AND U431 ( .A(n603), .B(n604), .Z(n602) );
  XOR U432 ( .A(p_input[457]), .B(n601), .Z(n604) );
  XOR U433 ( .A(n605), .B(n606), .Z(n601) );
  AND U434 ( .A(n607), .B(n608), .Z(n606) );
  IV U435 ( .A(n597), .Z(n600) );
  XOR U436 ( .A(n609), .B(n610), .Z(n597) );
  AND U437 ( .A(n611), .B(n612), .Z(n610) );
  XOR U438 ( .A(n613), .B(n614), .Z(n594) );
  AND U439 ( .A(n615), .B(n612), .Z(n614) );
  XNOR U440 ( .A(n613), .B(n609), .Z(n612) );
  XOR U441 ( .A(n616), .B(n617), .Z(n609) );
  AND U442 ( .A(n618), .B(n608), .Z(n617) );
  XNOR U443 ( .A(n619), .B(n605), .Z(n608) );
  XOR U444 ( .A(n620), .B(n621), .Z(n605) );
  AND U445 ( .A(n622), .B(n623), .Z(n621) );
  XOR U446 ( .A(p_input[473]), .B(n620), .Z(n623) );
  XOR U447 ( .A(n624), .B(n625), .Z(n620) );
  AND U448 ( .A(n626), .B(n627), .Z(n625) );
  IV U449 ( .A(n616), .Z(n619) );
  XOR U450 ( .A(n628), .B(n629), .Z(n616) );
  AND U451 ( .A(n630), .B(n631), .Z(n629) );
  XOR U452 ( .A(n632), .B(n633), .Z(n613) );
  AND U453 ( .A(n634), .B(n631), .Z(n633) );
  XNOR U454 ( .A(n632), .B(n628), .Z(n631) );
  XOR U455 ( .A(n635), .B(n636), .Z(n628) );
  AND U456 ( .A(n637), .B(n627), .Z(n636) );
  XNOR U457 ( .A(n638), .B(n624), .Z(n627) );
  XOR U458 ( .A(n639), .B(n640), .Z(n624) );
  AND U459 ( .A(n641), .B(n642), .Z(n640) );
  XOR U460 ( .A(p_input[489]), .B(n639), .Z(n642) );
  XOR U461 ( .A(n643), .B(n644), .Z(n639) );
  AND U462 ( .A(n645), .B(n646), .Z(n644) );
  IV U463 ( .A(n635), .Z(n638) );
  XOR U464 ( .A(n647), .B(n648), .Z(n635) );
  AND U465 ( .A(n649), .B(n650), .Z(n648) );
  XOR U466 ( .A(n651), .B(n652), .Z(n632) );
  AND U467 ( .A(n653), .B(n650), .Z(n652) );
  XNOR U468 ( .A(n651), .B(n647), .Z(n650) );
  XOR U469 ( .A(n654), .B(n655), .Z(n647) );
  AND U470 ( .A(n656), .B(n646), .Z(n655) );
  XNOR U471 ( .A(n657), .B(n643), .Z(n646) );
  XOR U472 ( .A(n658), .B(n659), .Z(n643) );
  AND U473 ( .A(n660), .B(n661), .Z(n659) );
  XOR U474 ( .A(p_input[505]), .B(n658), .Z(n661) );
  XOR U475 ( .A(n662), .B(n663), .Z(n658) );
  AND U476 ( .A(n664), .B(n665), .Z(n663) );
  IV U477 ( .A(n654), .Z(n657) );
  XOR U478 ( .A(n666), .B(n667), .Z(n654) );
  AND U479 ( .A(n668), .B(n669), .Z(n667) );
  XOR U480 ( .A(n670), .B(n671), .Z(n651) );
  AND U481 ( .A(n672), .B(n669), .Z(n671) );
  XNOR U482 ( .A(n670), .B(n666), .Z(n669) );
  XOR U483 ( .A(n673), .B(n674), .Z(n666) );
  AND U484 ( .A(n675), .B(n665), .Z(n674) );
  XNOR U485 ( .A(n676), .B(n662), .Z(n665) );
  XOR U486 ( .A(n677), .B(n678), .Z(n662) );
  AND U487 ( .A(n679), .B(n680), .Z(n678) );
  XOR U488 ( .A(p_input[521]), .B(n677), .Z(n680) );
  XOR U489 ( .A(n681), .B(n682), .Z(n677) );
  AND U490 ( .A(n683), .B(n684), .Z(n682) );
  IV U491 ( .A(n673), .Z(n676) );
  XOR U492 ( .A(n685), .B(n686), .Z(n673) );
  AND U493 ( .A(n687), .B(n688), .Z(n686) );
  XOR U494 ( .A(n689), .B(n690), .Z(n670) );
  AND U495 ( .A(n691), .B(n688), .Z(n690) );
  XNOR U496 ( .A(n689), .B(n685), .Z(n688) );
  XOR U497 ( .A(n692), .B(n693), .Z(n685) );
  AND U498 ( .A(n694), .B(n684), .Z(n693) );
  XNOR U499 ( .A(n695), .B(n681), .Z(n684) );
  XOR U500 ( .A(n696), .B(n697), .Z(n681) );
  AND U501 ( .A(n698), .B(n699), .Z(n697) );
  XOR U502 ( .A(p_input[537]), .B(n696), .Z(n699) );
  XOR U503 ( .A(n700), .B(n701), .Z(n696) );
  AND U504 ( .A(n702), .B(n703), .Z(n701) );
  IV U505 ( .A(n692), .Z(n695) );
  XOR U506 ( .A(n704), .B(n705), .Z(n692) );
  AND U507 ( .A(n706), .B(n707), .Z(n705) );
  XOR U508 ( .A(n708), .B(n709), .Z(n689) );
  AND U509 ( .A(n710), .B(n707), .Z(n709) );
  XNOR U510 ( .A(n708), .B(n704), .Z(n707) );
  XOR U511 ( .A(n711), .B(n712), .Z(n704) );
  AND U512 ( .A(n713), .B(n703), .Z(n712) );
  XNOR U513 ( .A(n714), .B(n700), .Z(n703) );
  XOR U514 ( .A(n715), .B(n716), .Z(n700) );
  AND U515 ( .A(n717), .B(n718), .Z(n716) );
  XOR U516 ( .A(p_input[553]), .B(n715), .Z(n718) );
  XOR U517 ( .A(n719), .B(n720), .Z(n715) );
  AND U518 ( .A(n721), .B(n722), .Z(n720) );
  IV U519 ( .A(n711), .Z(n714) );
  XOR U520 ( .A(n723), .B(n724), .Z(n711) );
  AND U521 ( .A(n725), .B(n726), .Z(n724) );
  XOR U522 ( .A(n727), .B(n728), .Z(n708) );
  AND U523 ( .A(n729), .B(n726), .Z(n728) );
  XNOR U524 ( .A(n727), .B(n723), .Z(n726) );
  XOR U525 ( .A(n730), .B(n731), .Z(n723) );
  AND U526 ( .A(n732), .B(n722), .Z(n731) );
  XNOR U527 ( .A(n733), .B(n719), .Z(n722) );
  XOR U528 ( .A(n734), .B(n735), .Z(n719) );
  AND U529 ( .A(n736), .B(n737), .Z(n735) );
  XOR U530 ( .A(p_input[569]), .B(n734), .Z(n737) );
  XOR U531 ( .A(n738), .B(n739), .Z(n734) );
  AND U532 ( .A(n740), .B(n741), .Z(n739) );
  IV U533 ( .A(n730), .Z(n733) );
  XOR U534 ( .A(n742), .B(n743), .Z(n730) );
  AND U535 ( .A(n744), .B(n745), .Z(n743) );
  XOR U536 ( .A(n746), .B(n747), .Z(n727) );
  AND U537 ( .A(n748), .B(n745), .Z(n747) );
  XNOR U538 ( .A(n746), .B(n742), .Z(n745) );
  XOR U539 ( .A(n749), .B(n750), .Z(n742) );
  AND U540 ( .A(n751), .B(n741), .Z(n750) );
  XNOR U541 ( .A(n752), .B(n738), .Z(n741) );
  XOR U542 ( .A(n753), .B(n754), .Z(n738) );
  AND U543 ( .A(n755), .B(n756), .Z(n754) );
  XOR U544 ( .A(p_input[585]), .B(n753), .Z(n756) );
  XOR U545 ( .A(n757), .B(n758), .Z(n753) );
  AND U546 ( .A(n759), .B(n760), .Z(n758) );
  IV U547 ( .A(n749), .Z(n752) );
  XOR U548 ( .A(n761), .B(n762), .Z(n749) );
  AND U549 ( .A(n763), .B(n764), .Z(n762) );
  XOR U550 ( .A(n765), .B(n766), .Z(n746) );
  AND U551 ( .A(n767), .B(n764), .Z(n766) );
  XNOR U552 ( .A(n765), .B(n761), .Z(n764) );
  XOR U553 ( .A(n768), .B(n769), .Z(n761) );
  AND U554 ( .A(n770), .B(n760), .Z(n769) );
  XNOR U555 ( .A(n771), .B(n757), .Z(n760) );
  XOR U556 ( .A(n772), .B(n773), .Z(n757) );
  AND U557 ( .A(n774), .B(n775), .Z(n773) );
  XOR U558 ( .A(p_input[601]), .B(n772), .Z(n775) );
  XOR U559 ( .A(n776), .B(n777), .Z(n772) );
  AND U560 ( .A(n778), .B(n779), .Z(n777) );
  IV U561 ( .A(n768), .Z(n771) );
  XOR U562 ( .A(n780), .B(n781), .Z(n768) );
  AND U563 ( .A(n782), .B(n783), .Z(n781) );
  XOR U564 ( .A(n784), .B(n785), .Z(n765) );
  AND U565 ( .A(n786), .B(n783), .Z(n785) );
  XNOR U566 ( .A(n784), .B(n780), .Z(n783) );
  XOR U567 ( .A(n787), .B(n788), .Z(n780) );
  AND U568 ( .A(n789), .B(n779), .Z(n788) );
  XNOR U569 ( .A(n790), .B(n776), .Z(n779) );
  XOR U570 ( .A(n791), .B(n792), .Z(n776) );
  AND U571 ( .A(n793), .B(n794), .Z(n792) );
  XOR U572 ( .A(p_input[617]), .B(n791), .Z(n794) );
  XOR U573 ( .A(n795), .B(n796), .Z(n791) );
  AND U574 ( .A(n797), .B(n798), .Z(n796) );
  IV U575 ( .A(n787), .Z(n790) );
  XOR U576 ( .A(n799), .B(n800), .Z(n787) );
  AND U577 ( .A(n801), .B(n802), .Z(n800) );
  XOR U578 ( .A(n803), .B(n804), .Z(n784) );
  AND U579 ( .A(n805), .B(n802), .Z(n804) );
  XNOR U580 ( .A(n803), .B(n799), .Z(n802) );
  XOR U581 ( .A(n806), .B(n807), .Z(n799) );
  AND U582 ( .A(n808), .B(n798), .Z(n807) );
  XNOR U583 ( .A(n809), .B(n795), .Z(n798) );
  XOR U584 ( .A(n810), .B(n811), .Z(n795) );
  AND U585 ( .A(n812), .B(n813), .Z(n811) );
  XOR U586 ( .A(p_input[633]), .B(n810), .Z(n813) );
  XOR U587 ( .A(n814), .B(n815), .Z(n810) );
  AND U588 ( .A(n816), .B(n817), .Z(n815) );
  IV U589 ( .A(n806), .Z(n809) );
  XOR U590 ( .A(n818), .B(n819), .Z(n806) );
  AND U591 ( .A(n820), .B(n821), .Z(n819) );
  XOR U592 ( .A(n822), .B(n823), .Z(n803) );
  AND U593 ( .A(n824), .B(n821), .Z(n823) );
  XNOR U594 ( .A(n822), .B(n818), .Z(n821) );
  XOR U595 ( .A(n825), .B(n826), .Z(n818) );
  AND U596 ( .A(n827), .B(n817), .Z(n826) );
  XNOR U597 ( .A(n828), .B(n814), .Z(n817) );
  XOR U598 ( .A(n829), .B(n830), .Z(n814) );
  AND U599 ( .A(n831), .B(n832), .Z(n830) );
  XOR U600 ( .A(p_input[649]), .B(n829), .Z(n832) );
  XOR U601 ( .A(n833), .B(n834), .Z(n829) );
  AND U602 ( .A(n835), .B(n836), .Z(n834) );
  IV U603 ( .A(n825), .Z(n828) );
  XOR U604 ( .A(n837), .B(n838), .Z(n825) );
  AND U605 ( .A(n839), .B(n840), .Z(n838) );
  XOR U606 ( .A(n841), .B(n842), .Z(n822) );
  AND U607 ( .A(n843), .B(n840), .Z(n842) );
  XNOR U608 ( .A(n841), .B(n837), .Z(n840) );
  XOR U609 ( .A(n844), .B(n845), .Z(n837) );
  AND U610 ( .A(n846), .B(n836), .Z(n845) );
  XNOR U611 ( .A(n847), .B(n833), .Z(n836) );
  XOR U612 ( .A(n848), .B(n849), .Z(n833) );
  AND U613 ( .A(n850), .B(n851), .Z(n849) );
  XOR U614 ( .A(p_input[665]), .B(n848), .Z(n851) );
  XOR U615 ( .A(n852), .B(n853), .Z(n848) );
  AND U616 ( .A(n854), .B(n855), .Z(n853) );
  IV U617 ( .A(n844), .Z(n847) );
  XOR U618 ( .A(n856), .B(n857), .Z(n844) );
  AND U619 ( .A(n858), .B(n859), .Z(n857) );
  XOR U620 ( .A(n860), .B(n861), .Z(n841) );
  AND U621 ( .A(n862), .B(n859), .Z(n861) );
  XNOR U622 ( .A(n860), .B(n856), .Z(n859) );
  XOR U623 ( .A(n863), .B(n864), .Z(n856) );
  AND U624 ( .A(n865), .B(n855), .Z(n864) );
  XNOR U625 ( .A(n866), .B(n852), .Z(n855) );
  XOR U626 ( .A(n867), .B(n868), .Z(n852) );
  AND U627 ( .A(n869), .B(n870), .Z(n868) );
  XOR U628 ( .A(p_input[681]), .B(n867), .Z(n870) );
  XOR U629 ( .A(n871), .B(n872), .Z(n867) );
  AND U630 ( .A(n873), .B(n874), .Z(n872) );
  IV U631 ( .A(n863), .Z(n866) );
  XOR U632 ( .A(n875), .B(n876), .Z(n863) );
  AND U633 ( .A(n877), .B(n878), .Z(n876) );
  XOR U634 ( .A(n879), .B(n880), .Z(n860) );
  AND U635 ( .A(n881), .B(n878), .Z(n880) );
  XNOR U636 ( .A(n879), .B(n875), .Z(n878) );
  XOR U637 ( .A(n882), .B(n883), .Z(n875) );
  AND U638 ( .A(n884), .B(n874), .Z(n883) );
  XNOR U639 ( .A(n885), .B(n871), .Z(n874) );
  XOR U640 ( .A(n886), .B(n887), .Z(n871) );
  AND U641 ( .A(n888), .B(n889), .Z(n887) );
  XOR U642 ( .A(p_input[697]), .B(n886), .Z(n889) );
  XOR U643 ( .A(n890), .B(n891), .Z(n886) );
  AND U644 ( .A(n892), .B(n893), .Z(n891) );
  IV U645 ( .A(n882), .Z(n885) );
  XOR U646 ( .A(n894), .B(n895), .Z(n882) );
  AND U647 ( .A(n896), .B(n897), .Z(n895) );
  XOR U648 ( .A(n898), .B(n899), .Z(n879) );
  AND U649 ( .A(n900), .B(n897), .Z(n899) );
  XNOR U650 ( .A(n898), .B(n894), .Z(n897) );
  XOR U651 ( .A(n901), .B(n902), .Z(n894) );
  AND U652 ( .A(n903), .B(n893), .Z(n902) );
  XNOR U653 ( .A(n904), .B(n890), .Z(n893) );
  XOR U654 ( .A(n905), .B(n906), .Z(n890) );
  AND U655 ( .A(n907), .B(n908), .Z(n906) );
  XOR U656 ( .A(p_input[713]), .B(n905), .Z(n908) );
  XOR U657 ( .A(n909), .B(n910), .Z(n905) );
  AND U658 ( .A(n911), .B(n912), .Z(n910) );
  IV U659 ( .A(n901), .Z(n904) );
  XOR U660 ( .A(n913), .B(n914), .Z(n901) );
  AND U661 ( .A(n915), .B(n916), .Z(n914) );
  XOR U662 ( .A(n917), .B(n918), .Z(n898) );
  AND U663 ( .A(n919), .B(n916), .Z(n918) );
  XNOR U664 ( .A(n917), .B(n913), .Z(n916) );
  XOR U665 ( .A(n920), .B(n921), .Z(n913) );
  AND U666 ( .A(n922), .B(n912), .Z(n921) );
  XNOR U667 ( .A(n923), .B(n909), .Z(n912) );
  XOR U668 ( .A(n924), .B(n925), .Z(n909) );
  AND U669 ( .A(n926), .B(n927), .Z(n925) );
  XOR U670 ( .A(p_input[729]), .B(n924), .Z(n927) );
  XOR U671 ( .A(n928), .B(n929), .Z(n924) );
  AND U672 ( .A(n930), .B(n931), .Z(n929) );
  IV U673 ( .A(n920), .Z(n923) );
  XOR U674 ( .A(n932), .B(n933), .Z(n920) );
  AND U675 ( .A(n934), .B(n935), .Z(n933) );
  XOR U676 ( .A(n936), .B(n937), .Z(n917) );
  AND U677 ( .A(n938), .B(n935), .Z(n937) );
  XNOR U678 ( .A(n936), .B(n932), .Z(n935) );
  XOR U679 ( .A(n939), .B(n940), .Z(n932) );
  AND U680 ( .A(n941), .B(n931), .Z(n940) );
  XNOR U681 ( .A(n942), .B(n928), .Z(n931) );
  XOR U682 ( .A(n943), .B(n944), .Z(n928) );
  AND U683 ( .A(n945), .B(n946), .Z(n944) );
  XOR U684 ( .A(p_input[745]), .B(n943), .Z(n946) );
  XOR U685 ( .A(n947), .B(n948), .Z(n943) );
  AND U686 ( .A(n949), .B(n950), .Z(n948) );
  IV U687 ( .A(n939), .Z(n942) );
  XOR U688 ( .A(n951), .B(n952), .Z(n939) );
  AND U689 ( .A(n953), .B(n954), .Z(n952) );
  XOR U690 ( .A(n955), .B(n956), .Z(n936) );
  AND U691 ( .A(n957), .B(n954), .Z(n956) );
  XNOR U692 ( .A(n955), .B(n951), .Z(n954) );
  XOR U693 ( .A(n958), .B(n959), .Z(n951) );
  AND U694 ( .A(n960), .B(n950), .Z(n959) );
  XNOR U695 ( .A(n961), .B(n947), .Z(n950) );
  XOR U696 ( .A(n962), .B(n963), .Z(n947) );
  AND U697 ( .A(n964), .B(n965), .Z(n963) );
  XOR U698 ( .A(p_input[761]), .B(n962), .Z(n965) );
  XOR U699 ( .A(n966), .B(n967), .Z(n962) );
  AND U700 ( .A(n968), .B(n969), .Z(n967) );
  IV U701 ( .A(n958), .Z(n961) );
  XOR U702 ( .A(n970), .B(n971), .Z(n958) );
  AND U703 ( .A(n972), .B(n973), .Z(n971) );
  XOR U704 ( .A(n974), .B(n975), .Z(n955) );
  AND U705 ( .A(n976), .B(n973), .Z(n975) );
  XNOR U706 ( .A(n974), .B(n970), .Z(n973) );
  XOR U707 ( .A(n977), .B(n978), .Z(n970) );
  AND U708 ( .A(n979), .B(n969), .Z(n978) );
  XNOR U709 ( .A(n980), .B(n966), .Z(n969) );
  XOR U710 ( .A(n981), .B(n982), .Z(n966) );
  AND U711 ( .A(n983), .B(n984), .Z(n982) );
  XOR U712 ( .A(p_input[777]), .B(n981), .Z(n984) );
  XOR U713 ( .A(n985), .B(n986), .Z(n981) );
  AND U714 ( .A(n987), .B(n988), .Z(n986) );
  IV U715 ( .A(n977), .Z(n980) );
  XOR U716 ( .A(n989), .B(n990), .Z(n977) );
  AND U717 ( .A(n991), .B(n992), .Z(n990) );
  XOR U718 ( .A(n993), .B(n994), .Z(n974) );
  AND U719 ( .A(n995), .B(n992), .Z(n994) );
  XNOR U720 ( .A(n993), .B(n989), .Z(n992) );
  XOR U721 ( .A(n996), .B(n997), .Z(n989) );
  AND U722 ( .A(n998), .B(n988), .Z(n997) );
  XNOR U723 ( .A(n999), .B(n985), .Z(n988) );
  XOR U724 ( .A(n1000), .B(n1001), .Z(n985) );
  AND U725 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U726 ( .A(p_input[793]), .B(n1000), .Z(n1003) );
  XOR U727 ( .A(n1004), .B(n1005), .Z(n1000) );
  AND U728 ( .A(n1006), .B(n1007), .Z(n1005) );
  IV U729 ( .A(n996), .Z(n999) );
  XOR U730 ( .A(n1008), .B(n1009), .Z(n996) );
  AND U731 ( .A(n1010), .B(n1011), .Z(n1009) );
  XOR U732 ( .A(n1012), .B(n1013), .Z(n993) );
  AND U733 ( .A(n1014), .B(n1011), .Z(n1013) );
  XNOR U734 ( .A(n1012), .B(n1008), .Z(n1011) );
  XOR U735 ( .A(n1015), .B(n1016), .Z(n1008) );
  AND U736 ( .A(n1017), .B(n1007), .Z(n1016) );
  XNOR U737 ( .A(n1018), .B(n1004), .Z(n1007) );
  XOR U738 ( .A(n1019), .B(n1020), .Z(n1004) );
  AND U739 ( .A(n1021), .B(n1022), .Z(n1020) );
  XOR U740 ( .A(p_input[809]), .B(n1019), .Z(n1022) );
  XOR U741 ( .A(n1023), .B(n1024), .Z(n1019) );
  AND U742 ( .A(n1025), .B(n1026), .Z(n1024) );
  IV U743 ( .A(n1015), .Z(n1018) );
  XOR U744 ( .A(n1027), .B(n1028), .Z(n1015) );
  AND U745 ( .A(n1029), .B(n1030), .Z(n1028) );
  XOR U746 ( .A(n1031), .B(n1032), .Z(n1012) );
  AND U747 ( .A(n1033), .B(n1030), .Z(n1032) );
  XNOR U748 ( .A(n1031), .B(n1027), .Z(n1030) );
  XOR U749 ( .A(n1034), .B(n1035), .Z(n1027) );
  AND U750 ( .A(n1036), .B(n1026), .Z(n1035) );
  XNOR U751 ( .A(n1037), .B(n1023), .Z(n1026) );
  XOR U752 ( .A(n1038), .B(n1039), .Z(n1023) );
  AND U753 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U754 ( .A(p_input[825]), .B(n1038), .Z(n1041) );
  XOR U755 ( .A(n1042), .B(n1043), .Z(n1038) );
  AND U756 ( .A(n1044), .B(n1045), .Z(n1043) );
  IV U757 ( .A(n1034), .Z(n1037) );
  XOR U758 ( .A(n1046), .B(n1047), .Z(n1034) );
  AND U759 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U760 ( .A(n1050), .B(n1051), .Z(n1031) );
  AND U761 ( .A(n1052), .B(n1049), .Z(n1051) );
  XNOR U762 ( .A(n1050), .B(n1046), .Z(n1049) );
  XOR U763 ( .A(n1053), .B(n1054), .Z(n1046) );
  AND U764 ( .A(n1055), .B(n1045), .Z(n1054) );
  XNOR U765 ( .A(n1056), .B(n1042), .Z(n1045) );
  XOR U766 ( .A(n1057), .B(n1058), .Z(n1042) );
  AND U767 ( .A(n1059), .B(n1060), .Z(n1058) );
  XOR U768 ( .A(p_input[841]), .B(n1057), .Z(n1060) );
  XOR U769 ( .A(n1061), .B(n1062), .Z(n1057) );
  AND U770 ( .A(n1063), .B(n1064), .Z(n1062) );
  IV U771 ( .A(n1053), .Z(n1056) );
  XOR U772 ( .A(n1065), .B(n1066), .Z(n1053) );
  AND U773 ( .A(n1067), .B(n1068), .Z(n1066) );
  XOR U774 ( .A(n1069), .B(n1070), .Z(n1050) );
  AND U775 ( .A(n1071), .B(n1068), .Z(n1070) );
  XNOR U776 ( .A(n1069), .B(n1065), .Z(n1068) );
  XOR U777 ( .A(n1072), .B(n1073), .Z(n1065) );
  AND U778 ( .A(n1074), .B(n1064), .Z(n1073) );
  XNOR U779 ( .A(n1075), .B(n1061), .Z(n1064) );
  XOR U780 ( .A(n1076), .B(n1077), .Z(n1061) );
  AND U781 ( .A(n1078), .B(n1079), .Z(n1077) );
  XOR U782 ( .A(p_input[857]), .B(n1076), .Z(n1079) );
  XOR U783 ( .A(n1080), .B(n1081), .Z(n1076) );
  AND U784 ( .A(n1082), .B(n1083), .Z(n1081) );
  IV U785 ( .A(n1072), .Z(n1075) );
  XOR U786 ( .A(n1084), .B(n1085), .Z(n1072) );
  AND U787 ( .A(n1086), .B(n1087), .Z(n1085) );
  XOR U788 ( .A(n1088), .B(n1089), .Z(n1069) );
  AND U789 ( .A(n1090), .B(n1087), .Z(n1089) );
  XNOR U790 ( .A(n1088), .B(n1084), .Z(n1087) );
  XOR U791 ( .A(n1091), .B(n1092), .Z(n1084) );
  AND U792 ( .A(n1093), .B(n1083), .Z(n1092) );
  XNOR U793 ( .A(n1094), .B(n1080), .Z(n1083) );
  XOR U794 ( .A(n1095), .B(n1096), .Z(n1080) );
  AND U795 ( .A(n1097), .B(n1098), .Z(n1096) );
  XOR U796 ( .A(p_input[873]), .B(n1095), .Z(n1098) );
  XOR U797 ( .A(n1099), .B(n1100), .Z(n1095) );
  AND U798 ( .A(n1101), .B(n1102), .Z(n1100) );
  IV U799 ( .A(n1091), .Z(n1094) );
  XOR U800 ( .A(n1103), .B(n1104), .Z(n1091) );
  AND U801 ( .A(n1105), .B(n1106), .Z(n1104) );
  XOR U802 ( .A(n1107), .B(n1108), .Z(n1088) );
  AND U803 ( .A(n1109), .B(n1106), .Z(n1108) );
  XNOR U804 ( .A(n1107), .B(n1103), .Z(n1106) );
  XOR U805 ( .A(n1110), .B(n1111), .Z(n1103) );
  AND U806 ( .A(n1112), .B(n1102), .Z(n1111) );
  XNOR U807 ( .A(n1113), .B(n1099), .Z(n1102) );
  XOR U808 ( .A(n1114), .B(n1115), .Z(n1099) );
  AND U809 ( .A(n1116), .B(n1117), .Z(n1115) );
  XOR U810 ( .A(p_input[889]), .B(n1114), .Z(n1117) );
  XOR U811 ( .A(n1118), .B(n1119), .Z(n1114) );
  AND U812 ( .A(n1120), .B(n1121), .Z(n1119) );
  IV U813 ( .A(n1110), .Z(n1113) );
  XOR U814 ( .A(n1122), .B(n1123), .Z(n1110) );
  AND U815 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U816 ( .A(n1126), .B(n1127), .Z(n1107) );
  AND U817 ( .A(n1128), .B(n1125), .Z(n1127) );
  XNOR U818 ( .A(n1126), .B(n1122), .Z(n1125) );
  XOR U819 ( .A(n1129), .B(n1130), .Z(n1122) );
  AND U820 ( .A(n1131), .B(n1121), .Z(n1130) );
  XNOR U821 ( .A(n1132), .B(n1118), .Z(n1121) );
  XOR U822 ( .A(n1133), .B(n1134), .Z(n1118) );
  AND U823 ( .A(n1135), .B(n1136), .Z(n1134) );
  XOR U824 ( .A(p_input[905]), .B(n1133), .Z(n1136) );
  XOR U825 ( .A(n1137), .B(n1138), .Z(n1133) );
  AND U826 ( .A(n1139), .B(n1140), .Z(n1138) );
  IV U827 ( .A(n1129), .Z(n1132) );
  XOR U828 ( .A(n1141), .B(n1142), .Z(n1129) );
  AND U829 ( .A(n1143), .B(n1144), .Z(n1142) );
  XOR U830 ( .A(n1145), .B(n1146), .Z(n1126) );
  AND U831 ( .A(n1147), .B(n1144), .Z(n1146) );
  XNOR U832 ( .A(n1145), .B(n1141), .Z(n1144) );
  XOR U833 ( .A(n1148), .B(n1149), .Z(n1141) );
  AND U834 ( .A(n1150), .B(n1140), .Z(n1149) );
  XNOR U835 ( .A(n1151), .B(n1137), .Z(n1140) );
  XOR U836 ( .A(n1152), .B(n1153), .Z(n1137) );
  AND U837 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U838 ( .A(p_input[921]), .B(n1152), .Z(n1155) );
  XOR U839 ( .A(n1156), .B(n1157), .Z(n1152) );
  AND U840 ( .A(n1158), .B(n1159), .Z(n1157) );
  IV U841 ( .A(n1148), .Z(n1151) );
  XOR U842 ( .A(n1160), .B(n1161), .Z(n1148) );
  AND U843 ( .A(n1162), .B(n1163), .Z(n1161) );
  XOR U844 ( .A(n1164), .B(n1165), .Z(n1145) );
  AND U845 ( .A(n1166), .B(n1163), .Z(n1165) );
  XNOR U846 ( .A(n1164), .B(n1160), .Z(n1163) );
  XOR U847 ( .A(n1167), .B(n1168), .Z(n1160) );
  AND U848 ( .A(n1169), .B(n1159), .Z(n1168) );
  XNOR U849 ( .A(n1170), .B(n1156), .Z(n1159) );
  XOR U850 ( .A(n1171), .B(n1172), .Z(n1156) );
  AND U851 ( .A(n1173), .B(n1174), .Z(n1172) );
  XOR U852 ( .A(p_input[937]), .B(n1171), .Z(n1174) );
  XOR U853 ( .A(n1175), .B(n1176), .Z(n1171) );
  AND U854 ( .A(n1177), .B(n1178), .Z(n1176) );
  IV U855 ( .A(n1167), .Z(n1170) );
  XOR U856 ( .A(n1179), .B(n1180), .Z(n1167) );
  AND U857 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U858 ( .A(n1183), .B(n1184), .Z(n1164) );
  AND U859 ( .A(n1185), .B(n1182), .Z(n1184) );
  XNOR U860 ( .A(n1183), .B(n1179), .Z(n1182) );
  XOR U861 ( .A(n1186), .B(n1187), .Z(n1179) );
  AND U862 ( .A(n1188), .B(n1178), .Z(n1187) );
  XNOR U863 ( .A(n1189), .B(n1175), .Z(n1178) );
  XOR U864 ( .A(n1190), .B(n1191), .Z(n1175) );
  AND U865 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U866 ( .A(p_input[953]), .B(n1190), .Z(n1193) );
  XOR U867 ( .A(n1194), .B(n1195), .Z(n1190) );
  AND U868 ( .A(n1196), .B(n1197), .Z(n1195) );
  IV U869 ( .A(n1186), .Z(n1189) );
  XOR U870 ( .A(n1198), .B(n1199), .Z(n1186) );
  AND U871 ( .A(n1200), .B(n1201), .Z(n1199) );
  XOR U872 ( .A(n1202), .B(n1203), .Z(n1183) );
  AND U873 ( .A(n1204), .B(n1201), .Z(n1203) );
  XNOR U874 ( .A(n1202), .B(n1198), .Z(n1201) );
  XOR U875 ( .A(n1205), .B(n1206), .Z(n1198) );
  AND U876 ( .A(n1207), .B(n1197), .Z(n1206) );
  XNOR U877 ( .A(n1208), .B(n1194), .Z(n1197) );
  XOR U878 ( .A(n1209), .B(n1210), .Z(n1194) );
  AND U879 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U880 ( .A(p_input[969]), .B(n1209), .Z(n1212) );
  XOR U881 ( .A(n1213), .B(n1214), .Z(n1209) );
  AND U882 ( .A(n1215), .B(n1216), .Z(n1214) );
  IV U883 ( .A(n1205), .Z(n1208) );
  XOR U884 ( .A(n1217), .B(n1218), .Z(n1205) );
  AND U885 ( .A(n1219), .B(n1220), .Z(n1218) );
  XOR U886 ( .A(n1221), .B(n1222), .Z(n1202) );
  AND U887 ( .A(n1223), .B(n1220), .Z(n1222) );
  XNOR U888 ( .A(n1221), .B(n1217), .Z(n1220) );
  XOR U889 ( .A(n1224), .B(n1225), .Z(n1217) );
  AND U890 ( .A(n1226), .B(n1216), .Z(n1225) );
  XNOR U891 ( .A(n1227), .B(n1213), .Z(n1216) );
  XOR U892 ( .A(n1228), .B(n1229), .Z(n1213) );
  AND U893 ( .A(n1230), .B(n1231), .Z(n1229) );
  XOR U894 ( .A(p_input[985]), .B(n1228), .Z(n1231) );
  XOR U895 ( .A(n1232), .B(n1233), .Z(n1228) );
  AND U896 ( .A(n1234), .B(n1235), .Z(n1233) );
  IV U897 ( .A(n1224), .Z(n1227) );
  XOR U898 ( .A(n1236), .B(n1237), .Z(n1224) );
  AND U899 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U900 ( .A(n1240), .B(n1241), .Z(n1221) );
  AND U901 ( .A(n1242), .B(n1239), .Z(n1241) );
  XNOR U902 ( .A(n1240), .B(n1236), .Z(n1239) );
  XOR U903 ( .A(n1243), .B(n1244), .Z(n1236) );
  AND U904 ( .A(n1245), .B(n1235), .Z(n1244) );
  XNOR U905 ( .A(n1246), .B(n1232), .Z(n1235) );
  XOR U906 ( .A(n1247), .B(n1248), .Z(n1232) );
  AND U907 ( .A(n1249), .B(n1250), .Z(n1248) );
  XOR U908 ( .A(p_input[1001]), .B(n1247), .Z(n1250) );
  XOR U909 ( .A(n1251), .B(n1252), .Z(n1247) );
  AND U910 ( .A(n1253), .B(n1254), .Z(n1252) );
  IV U911 ( .A(n1243), .Z(n1246) );
  XOR U912 ( .A(n1255), .B(n1256), .Z(n1243) );
  AND U913 ( .A(n1257), .B(n1258), .Z(n1256) );
  XOR U914 ( .A(n1259), .B(n1260), .Z(n1240) );
  AND U915 ( .A(n1261), .B(n1258), .Z(n1260) );
  XNOR U916 ( .A(n1259), .B(n1255), .Z(n1258) );
  XOR U917 ( .A(n1262), .B(n1263), .Z(n1255) );
  AND U918 ( .A(n1264), .B(n1254), .Z(n1263) );
  XNOR U919 ( .A(n1265), .B(n1251), .Z(n1254) );
  XOR U920 ( .A(n1266), .B(n1267), .Z(n1251) );
  AND U921 ( .A(n1268), .B(n1269), .Z(n1267) );
  XOR U922 ( .A(p_input[1017]), .B(n1266), .Z(n1269) );
  XOR U923 ( .A(n1270), .B(n1271), .Z(n1266) );
  AND U924 ( .A(n1272), .B(n1273), .Z(n1271) );
  IV U925 ( .A(n1262), .Z(n1265) );
  XOR U926 ( .A(n1274), .B(n1275), .Z(n1262) );
  AND U927 ( .A(n1276), .B(n1277), .Z(n1275) );
  XOR U928 ( .A(n1278), .B(n1279), .Z(n1259) );
  AND U929 ( .A(n1280), .B(n1277), .Z(n1279) );
  XNOR U930 ( .A(n1278), .B(n1274), .Z(n1277) );
  XOR U931 ( .A(n1281), .B(n1282), .Z(n1274) );
  AND U932 ( .A(n1283), .B(n1273), .Z(n1282) );
  XNOR U933 ( .A(n1284), .B(n1270), .Z(n1273) );
  XOR U934 ( .A(n1285), .B(n1286), .Z(n1270) );
  AND U935 ( .A(n1287), .B(n1288), .Z(n1286) );
  XOR U936 ( .A(p_input[1033]), .B(n1285), .Z(n1288) );
  XOR U937 ( .A(n1289), .B(n1290), .Z(n1285) );
  AND U938 ( .A(n1291), .B(n1292), .Z(n1290) );
  IV U939 ( .A(n1281), .Z(n1284) );
  XOR U940 ( .A(n1293), .B(n1294), .Z(n1281) );
  AND U941 ( .A(n1295), .B(n1296), .Z(n1294) );
  XOR U942 ( .A(n1297), .B(n1298), .Z(n1278) );
  AND U943 ( .A(n1299), .B(n1296), .Z(n1298) );
  XNOR U944 ( .A(n1297), .B(n1293), .Z(n1296) );
  XOR U945 ( .A(n1300), .B(n1301), .Z(n1293) );
  AND U946 ( .A(n1302), .B(n1292), .Z(n1301) );
  XNOR U947 ( .A(n1303), .B(n1289), .Z(n1292) );
  XOR U948 ( .A(n1304), .B(n1305), .Z(n1289) );
  AND U949 ( .A(n1306), .B(n1307), .Z(n1305) );
  XOR U950 ( .A(p_input[1049]), .B(n1304), .Z(n1307) );
  XOR U951 ( .A(n1308), .B(n1309), .Z(n1304) );
  AND U952 ( .A(n1310), .B(n1311), .Z(n1309) );
  IV U953 ( .A(n1300), .Z(n1303) );
  XOR U954 ( .A(n1312), .B(n1313), .Z(n1300) );
  AND U955 ( .A(n1314), .B(n1315), .Z(n1313) );
  XOR U956 ( .A(n1316), .B(n1317), .Z(n1297) );
  AND U957 ( .A(n1318), .B(n1315), .Z(n1317) );
  XNOR U958 ( .A(n1316), .B(n1312), .Z(n1315) );
  XOR U959 ( .A(n1319), .B(n1320), .Z(n1312) );
  AND U960 ( .A(n1321), .B(n1311), .Z(n1320) );
  XNOR U961 ( .A(n1322), .B(n1308), .Z(n1311) );
  XOR U962 ( .A(n1323), .B(n1324), .Z(n1308) );
  AND U963 ( .A(n1325), .B(n1326), .Z(n1324) );
  XOR U964 ( .A(p_input[1065]), .B(n1323), .Z(n1326) );
  XOR U965 ( .A(n1327), .B(n1328), .Z(n1323) );
  AND U966 ( .A(n1329), .B(n1330), .Z(n1328) );
  IV U967 ( .A(n1319), .Z(n1322) );
  XOR U968 ( .A(n1331), .B(n1332), .Z(n1319) );
  AND U969 ( .A(n1333), .B(n1334), .Z(n1332) );
  XOR U970 ( .A(n1335), .B(n1336), .Z(n1316) );
  AND U971 ( .A(n1337), .B(n1334), .Z(n1336) );
  XNOR U972 ( .A(n1335), .B(n1331), .Z(n1334) );
  XOR U973 ( .A(n1338), .B(n1339), .Z(n1331) );
  AND U974 ( .A(n1340), .B(n1330), .Z(n1339) );
  XNOR U975 ( .A(n1341), .B(n1327), .Z(n1330) );
  XOR U976 ( .A(n1342), .B(n1343), .Z(n1327) );
  AND U977 ( .A(n1344), .B(n1345), .Z(n1343) );
  XOR U978 ( .A(p_input[1081]), .B(n1342), .Z(n1345) );
  XOR U979 ( .A(n1346), .B(n1347), .Z(n1342) );
  AND U980 ( .A(n1348), .B(n1349), .Z(n1347) );
  IV U981 ( .A(n1338), .Z(n1341) );
  XOR U982 ( .A(n1350), .B(n1351), .Z(n1338) );
  AND U983 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR U984 ( .A(n1354), .B(n1355), .Z(n1335) );
  AND U985 ( .A(n1356), .B(n1353), .Z(n1355) );
  XNOR U986 ( .A(n1354), .B(n1350), .Z(n1353) );
  XOR U987 ( .A(n1357), .B(n1358), .Z(n1350) );
  AND U988 ( .A(n1359), .B(n1349), .Z(n1358) );
  XNOR U989 ( .A(n1360), .B(n1346), .Z(n1349) );
  XOR U990 ( .A(n1361), .B(n1362), .Z(n1346) );
  AND U991 ( .A(n1363), .B(n1364), .Z(n1362) );
  XOR U992 ( .A(p_input[1097]), .B(n1361), .Z(n1364) );
  XOR U993 ( .A(n1365), .B(n1366), .Z(n1361) );
  AND U994 ( .A(n1367), .B(n1368), .Z(n1366) );
  IV U995 ( .A(n1357), .Z(n1360) );
  XOR U996 ( .A(n1369), .B(n1370), .Z(n1357) );
  AND U997 ( .A(n1371), .B(n1372), .Z(n1370) );
  XOR U998 ( .A(n1373), .B(n1374), .Z(n1354) );
  AND U999 ( .A(n1375), .B(n1372), .Z(n1374) );
  XNOR U1000 ( .A(n1373), .B(n1369), .Z(n1372) );
  XOR U1001 ( .A(n1376), .B(n1377), .Z(n1369) );
  AND U1002 ( .A(n1378), .B(n1368), .Z(n1377) );
  XNOR U1003 ( .A(n1379), .B(n1365), .Z(n1368) );
  XOR U1004 ( .A(n1380), .B(n1381), .Z(n1365) );
  AND U1005 ( .A(n1382), .B(n1383), .Z(n1381) );
  XOR U1006 ( .A(p_input[1113]), .B(n1380), .Z(n1383) );
  XOR U1007 ( .A(n1384), .B(n1385), .Z(n1380) );
  AND U1008 ( .A(n1386), .B(n1387), .Z(n1385) );
  IV U1009 ( .A(n1376), .Z(n1379) );
  XOR U1010 ( .A(n1388), .B(n1389), .Z(n1376) );
  AND U1011 ( .A(n1390), .B(n1391), .Z(n1389) );
  XOR U1012 ( .A(n1392), .B(n1393), .Z(n1373) );
  AND U1013 ( .A(n1394), .B(n1391), .Z(n1393) );
  XNOR U1014 ( .A(n1392), .B(n1388), .Z(n1391) );
  XOR U1015 ( .A(n1395), .B(n1396), .Z(n1388) );
  AND U1016 ( .A(n1397), .B(n1387), .Z(n1396) );
  XNOR U1017 ( .A(n1398), .B(n1384), .Z(n1387) );
  XOR U1018 ( .A(n1399), .B(n1400), .Z(n1384) );
  AND U1019 ( .A(n1401), .B(n1402), .Z(n1400) );
  XOR U1020 ( .A(p_input[1129]), .B(n1399), .Z(n1402) );
  XOR U1021 ( .A(n1403), .B(n1404), .Z(n1399) );
  AND U1022 ( .A(n1405), .B(n1406), .Z(n1404) );
  IV U1023 ( .A(n1395), .Z(n1398) );
  XOR U1024 ( .A(n1407), .B(n1408), .Z(n1395) );
  AND U1025 ( .A(n1409), .B(n1410), .Z(n1408) );
  XOR U1026 ( .A(n1411), .B(n1412), .Z(n1392) );
  AND U1027 ( .A(n1413), .B(n1410), .Z(n1412) );
  XNOR U1028 ( .A(n1411), .B(n1407), .Z(n1410) );
  XOR U1029 ( .A(n1414), .B(n1415), .Z(n1407) );
  AND U1030 ( .A(n1416), .B(n1406), .Z(n1415) );
  XNOR U1031 ( .A(n1417), .B(n1403), .Z(n1406) );
  XOR U1032 ( .A(n1418), .B(n1419), .Z(n1403) );
  AND U1033 ( .A(n1420), .B(n1421), .Z(n1419) );
  XOR U1034 ( .A(p_input[1145]), .B(n1418), .Z(n1421) );
  XOR U1035 ( .A(n1422), .B(n1423), .Z(n1418) );
  AND U1036 ( .A(n1424), .B(n1425), .Z(n1423) );
  IV U1037 ( .A(n1414), .Z(n1417) );
  XOR U1038 ( .A(n1426), .B(n1427), .Z(n1414) );
  AND U1039 ( .A(n1428), .B(n1429), .Z(n1427) );
  XOR U1040 ( .A(n1430), .B(n1431), .Z(n1411) );
  AND U1041 ( .A(n1432), .B(n1429), .Z(n1431) );
  XNOR U1042 ( .A(n1430), .B(n1426), .Z(n1429) );
  XOR U1043 ( .A(n1433), .B(n1434), .Z(n1426) );
  AND U1044 ( .A(n1435), .B(n1425), .Z(n1434) );
  XNOR U1045 ( .A(n1436), .B(n1422), .Z(n1425) );
  XOR U1046 ( .A(n1437), .B(n1438), .Z(n1422) );
  AND U1047 ( .A(n1439), .B(n1440), .Z(n1438) );
  XOR U1048 ( .A(p_input[1161]), .B(n1437), .Z(n1440) );
  XOR U1049 ( .A(n1441), .B(n1442), .Z(n1437) );
  AND U1050 ( .A(n1443), .B(n1444), .Z(n1442) );
  IV U1051 ( .A(n1433), .Z(n1436) );
  XOR U1052 ( .A(n1445), .B(n1446), .Z(n1433) );
  AND U1053 ( .A(n1447), .B(n1448), .Z(n1446) );
  XOR U1054 ( .A(n1449), .B(n1450), .Z(n1430) );
  AND U1055 ( .A(n1451), .B(n1448), .Z(n1450) );
  XNOR U1056 ( .A(n1449), .B(n1445), .Z(n1448) );
  XOR U1057 ( .A(n1452), .B(n1453), .Z(n1445) );
  AND U1058 ( .A(n1454), .B(n1444), .Z(n1453) );
  XNOR U1059 ( .A(n1455), .B(n1441), .Z(n1444) );
  XOR U1060 ( .A(n1456), .B(n1457), .Z(n1441) );
  AND U1061 ( .A(n1458), .B(n1459), .Z(n1457) );
  XOR U1062 ( .A(p_input[1177]), .B(n1456), .Z(n1459) );
  XOR U1063 ( .A(n1460), .B(n1461), .Z(n1456) );
  AND U1064 ( .A(n1462), .B(n1463), .Z(n1461) );
  IV U1065 ( .A(n1452), .Z(n1455) );
  XOR U1066 ( .A(n1464), .B(n1465), .Z(n1452) );
  AND U1067 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U1068 ( .A(n1468), .B(n1469), .Z(n1449) );
  AND U1069 ( .A(n1470), .B(n1467), .Z(n1469) );
  XNOR U1070 ( .A(n1468), .B(n1464), .Z(n1467) );
  XOR U1071 ( .A(n1471), .B(n1472), .Z(n1464) );
  AND U1072 ( .A(n1473), .B(n1463), .Z(n1472) );
  XNOR U1073 ( .A(n1474), .B(n1460), .Z(n1463) );
  XOR U1074 ( .A(n1475), .B(n1476), .Z(n1460) );
  AND U1075 ( .A(n1477), .B(n1478), .Z(n1476) );
  XOR U1076 ( .A(p_input[1193]), .B(n1475), .Z(n1478) );
  XOR U1077 ( .A(n1479), .B(n1480), .Z(n1475) );
  AND U1078 ( .A(n1481), .B(n1482), .Z(n1480) );
  IV U1079 ( .A(n1471), .Z(n1474) );
  XOR U1080 ( .A(n1483), .B(n1484), .Z(n1471) );
  AND U1081 ( .A(n1485), .B(n1486), .Z(n1484) );
  XOR U1082 ( .A(n1487), .B(n1488), .Z(n1468) );
  AND U1083 ( .A(n1489), .B(n1486), .Z(n1488) );
  XNOR U1084 ( .A(n1487), .B(n1483), .Z(n1486) );
  XOR U1085 ( .A(n1490), .B(n1491), .Z(n1483) );
  AND U1086 ( .A(n1492), .B(n1482), .Z(n1491) );
  XNOR U1087 ( .A(n1493), .B(n1479), .Z(n1482) );
  XOR U1088 ( .A(n1494), .B(n1495), .Z(n1479) );
  AND U1089 ( .A(n1496), .B(n1497), .Z(n1495) );
  XOR U1090 ( .A(p_input[1209]), .B(n1494), .Z(n1497) );
  XOR U1091 ( .A(n1498), .B(n1499), .Z(n1494) );
  AND U1092 ( .A(n1500), .B(n1501), .Z(n1499) );
  IV U1093 ( .A(n1490), .Z(n1493) );
  XOR U1094 ( .A(n1502), .B(n1503), .Z(n1490) );
  AND U1095 ( .A(n1504), .B(n1505), .Z(n1503) );
  XOR U1096 ( .A(n1506), .B(n1507), .Z(n1487) );
  AND U1097 ( .A(n1508), .B(n1505), .Z(n1507) );
  XNOR U1098 ( .A(n1506), .B(n1502), .Z(n1505) );
  XOR U1099 ( .A(n1509), .B(n1510), .Z(n1502) );
  AND U1100 ( .A(n1511), .B(n1501), .Z(n1510) );
  XNOR U1101 ( .A(n1512), .B(n1498), .Z(n1501) );
  XOR U1102 ( .A(n1513), .B(n1514), .Z(n1498) );
  AND U1103 ( .A(n1515), .B(n1516), .Z(n1514) );
  XOR U1104 ( .A(p_input[1225]), .B(n1513), .Z(n1516) );
  XOR U1105 ( .A(n1517), .B(n1518), .Z(n1513) );
  AND U1106 ( .A(n1519), .B(n1520), .Z(n1518) );
  IV U1107 ( .A(n1509), .Z(n1512) );
  XOR U1108 ( .A(n1521), .B(n1522), .Z(n1509) );
  AND U1109 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U1110 ( .A(n1525), .B(n1526), .Z(n1506) );
  AND U1111 ( .A(n1527), .B(n1524), .Z(n1526) );
  XNOR U1112 ( .A(n1525), .B(n1521), .Z(n1524) );
  XOR U1113 ( .A(n1528), .B(n1529), .Z(n1521) );
  AND U1114 ( .A(n1530), .B(n1520), .Z(n1529) );
  XNOR U1115 ( .A(n1531), .B(n1517), .Z(n1520) );
  XOR U1116 ( .A(n1532), .B(n1533), .Z(n1517) );
  AND U1117 ( .A(n1534), .B(n1535), .Z(n1533) );
  XOR U1118 ( .A(p_input[1241]), .B(n1532), .Z(n1535) );
  XOR U1119 ( .A(n1536), .B(n1537), .Z(n1532) );
  AND U1120 ( .A(n1538), .B(n1539), .Z(n1537) );
  IV U1121 ( .A(n1528), .Z(n1531) );
  XOR U1122 ( .A(n1540), .B(n1541), .Z(n1528) );
  AND U1123 ( .A(n1542), .B(n1543), .Z(n1541) );
  XOR U1124 ( .A(n1544), .B(n1545), .Z(n1525) );
  AND U1125 ( .A(n1546), .B(n1543), .Z(n1545) );
  XNOR U1126 ( .A(n1544), .B(n1540), .Z(n1543) );
  XOR U1127 ( .A(n1547), .B(n1548), .Z(n1540) );
  AND U1128 ( .A(n1549), .B(n1539), .Z(n1548) );
  XNOR U1129 ( .A(n1550), .B(n1536), .Z(n1539) );
  XOR U1130 ( .A(n1551), .B(n1552), .Z(n1536) );
  AND U1131 ( .A(n1553), .B(n1554), .Z(n1552) );
  XOR U1132 ( .A(p_input[1257]), .B(n1551), .Z(n1554) );
  XOR U1133 ( .A(n1555), .B(n1556), .Z(n1551) );
  AND U1134 ( .A(n1557), .B(n1558), .Z(n1556) );
  IV U1135 ( .A(n1547), .Z(n1550) );
  XOR U1136 ( .A(n1559), .B(n1560), .Z(n1547) );
  AND U1137 ( .A(n1561), .B(n1562), .Z(n1560) );
  XOR U1138 ( .A(n1563), .B(n1564), .Z(n1544) );
  AND U1139 ( .A(n1565), .B(n1562), .Z(n1564) );
  XNOR U1140 ( .A(n1563), .B(n1559), .Z(n1562) );
  XOR U1141 ( .A(n1566), .B(n1567), .Z(n1559) );
  AND U1142 ( .A(n1568), .B(n1558), .Z(n1567) );
  XNOR U1143 ( .A(n1569), .B(n1555), .Z(n1558) );
  XOR U1144 ( .A(n1570), .B(n1571), .Z(n1555) );
  AND U1145 ( .A(n1572), .B(n1573), .Z(n1571) );
  XOR U1146 ( .A(p_input[1273]), .B(n1570), .Z(n1573) );
  XOR U1147 ( .A(n1574), .B(n1575), .Z(n1570) );
  AND U1148 ( .A(n1576), .B(n1577), .Z(n1575) );
  IV U1149 ( .A(n1566), .Z(n1569) );
  XOR U1150 ( .A(n1578), .B(n1579), .Z(n1566) );
  AND U1151 ( .A(n1580), .B(n1581), .Z(n1579) );
  XOR U1152 ( .A(n1582), .B(n1583), .Z(n1563) );
  AND U1153 ( .A(n1584), .B(n1581), .Z(n1583) );
  XNOR U1154 ( .A(n1582), .B(n1578), .Z(n1581) );
  XOR U1155 ( .A(n1585), .B(n1586), .Z(n1578) );
  AND U1156 ( .A(n1587), .B(n1577), .Z(n1586) );
  XNOR U1157 ( .A(n1588), .B(n1574), .Z(n1577) );
  XOR U1158 ( .A(n1589), .B(n1590), .Z(n1574) );
  AND U1159 ( .A(n1591), .B(n1592), .Z(n1590) );
  XOR U1160 ( .A(p_input[1289]), .B(n1589), .Z(n1592) );
  XOR U1161 ( .A(n1593), .B(n1594), .Z(n1589) );
  AND U1162 ( .A(n1595), .B(n1596), .Z(n1594) );
  IV U1163 ( .A(n1585), .Z(n1588) );
  XOR U1164 ( .A(n1597), .B(n1598), .Z(n1585) );
  AND U1165 ( .A(n1599), .B(n1600), .Z(n1598) );
  XOR U1166 ( .A(n1601), .B(n1602), .Z(n1582) );
  AND U1167 ( .A(n1603), .B(n1600), .Z(n1602) );
  XNOR U1168 ( .A(n1601), .B(n1597), .Z(n1600) );
  XOR U1169 ( .A(n1604), .B(n1605), .Z(n1597) );
  AND U1170 ( .A(n1606), .B(n1596), .Z(n1605) );
  XNOR U1171 ( .A(n1607), .B(n1593), .Z(n1596) );
  XOR U1172 ( .A(n1608), .B(n1609), .Z(n1593) );
  AND U1173 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U1174 ( .A(p_input[1305]), .B(n1608), .Z(n1611) );
  XOR U1175 ( .A(n1612), .B(n1613), .Z(n1608) );
  AND U1176 ( .A(n1614), .B(n1615), .Z(n1613) );
  IV U1177 ( .A(n1604), .Z(n1607) );
  XOR U1178 ( .A(n1616), .B(n1617), .Z(n1604) );
  AND U1179 ( .A(n1618), .B(n1619), .Z(n1617) );
  XOR U1180 ( .A(n1620), .B(n1621), .Z(n1601) );
  AND U1181 ( .A(n1622), .B(n1619), .Z(n1621) );
  XNOR U1182 ( .A(n1620), .B(n1616), .Z(n1619) );
  XOR U1183 ( .A(n1623), .B(n1624), .Z(n1616) );
  AND U1184 ( .A(n1625), .B(n1615), .Z(n1624) );
  XNOR U1185 ( .A(n1626), .B(n1612), .Z(n1615) );
  XOR U1186 ( .A(n1627), .B(n1628), .Z(n1612) );
  AND U1187 ( .A(n1629), .B(n1630), .Z(n1628) );
  XOR U1188 ( .A(p_input[1321]), .B(n1627), .Z(n1630) );
  XOR U1189 ( .A(n1631), .B(n1632), .Z(n1627) );
  AND U1190 ( .A(n1633), .B(n1634), .Z(n1632) );
  IV U1191 ( .A(n1623), .Z(n1626) );
  XOR U1192 ( .A(n1635), .B(n1636), .Z(n1623) );
  AND U1193 ( .A(n1637), .B(n1638), .Z(n1636) );
  XOR U1194 ( .A(n1639), .B(n1640), .Z(n1620) );
  AND U1195 ( .A(n1641), .B(n1638), .Z(n1640) );
  XNOR U1196 ( .A(n1639), .B(n1635), .Z(n1638) );
  XOR U1197 ( .A(n1642), .B(n1643), .Z(n1635) );
  AND U1198 ( .A(n1644), .B(n1634), .Z(n1643) );
  XNOR U1199 ( .A(n1645), .B(n1631), .Z(n1634) );
  XOR U1200 ( .A(n1646), .B(n1647), .Z(n1631) );
  AND U1201 ( .A(n1648), .B(n1649), .Z(n1647) );
  XOR U1202 ( .A(p_input[1337]), .B(n1646), .Z(n1649) );
  XOR U1203 ( .A(n1650), .B(n1651), .Z(n1646) );
  AND U1204 ( .A(n1652), .B(n1653), .Z(n1651) );
  IV U1205 ( .A(n1642), .Z(n1645) );
  XOR U1206 ( .A(n1654), .B(n1655), .Z(n1642) );
  AND U1207 ( .A(n1656), .B(n1657), .Z(n1655) );
  XOR U1208 ( .A(n1658), .B(n1659), .Z(n1639) );
  AND U1209 ( .A(n1660), .B(n1657), .Z(n1659) );
  XNOR U1210 ( .A(n1658), .B(n1654), .Z(n1657) );
  XOR U1211 ( .A(n1661), .B(n1662), .Z(n1654) );
  AND U1212 ( .A(n1663), .B(n1653), .Z(n1662) );
  XNOR U1213 ( .A(n1664), .B(n1650), .Z(n1653) );
  XOR U1214 ( .A(n1665), .B(n1666), .Z(n1650) );
  AND U1215 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U1216 ( .A(p_input[1353]), .B(n1665), .Z(n1668) );
  XOR U1217 ( .A(n1669), .B(n1670), .Z(n1665) );
  AND U1218 ( .A(n1671), .B(n1672), .Z(n1670) );
  IV U1219 ( .A(n1661), .Z(n1664) );
  XOR U1220 ( .A(n1673), .B(n1674), .Z(n1661) );
  AND U1221 ( .A(n1675), .B(n1676), .Z(n1674) );
  XOR U1222 ( .A(n1677), .B(n1678), .Z(n1658) );
  AND U1223 ( .A(n1679), .B(n1676), .Z(n1678) );
  XNOR U1224 ( .A(n1677), .B(n1673), .Z(n1676) );
  XOR U1225 ( .A(n1680), .B(n1681), .Z(n1673) );
  AND U1226 ( .A(n1682), .B(n1672), .Z(n1681) );
  XNOR U1227 ( .A(n1683), .B(n1669), .Z(n1672) );
  XOR U1228 ( .A(n1684), .B(n1685), .Z(n1669) );
  AND U1229 ( .A(n1686), .B(n1687), .Z(n1685) );
  XOR U1230 ( .A(p_input[1369]), .B(n1684), .Z(n1687) );
  XOR U1231 ( .A(n1688), .B(n1689), .Z(n1684) );
  AND U1232 ( .A(n1690), .B(n1691), .Z(n1689) );
  IV U1233 ( .A(n1680), .Z(n1683) );
  XOR U1234 ( .A(n1692), .B(n1693), .Z(n1680) );
  AND U1235 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U1236 ( .A(n1696), .B(n1697), .Z(n1677) );
  AND U1237 ( .A(n1698), .B(n1695), .Z(n1697) );
  XNOR U1238 ( .A(n1696), .B(n1692), .Z(n1695) );
  XOR U1239 ( .A(n1699), .B(n1700), .Z(n1692) );
  AND U1240 ( .A(n1701), .B(n1691), .Z(n1700) );
  XNOR U1241 ( .A(n1702), .B(n1688), .Z(n1691) );
  XOR U1242 ( .A(n1703), .B(n1704), .Z(n1688) );
  AND U1243 ( .A(n1705), .B(n1706), .Z(n1704) );
  XOR U1244 ( .A(p_input[1385]), .B(n1703), .Z(n1706) );
  XOR U1245 ( .A(n1707), .B(n1708), .Z(n1703) );
  AND U1246 ( .A(n1709), .B(n1710), .Z(n1708) );
  IV U1247 ( .A(n1699), .Z(n1702) );
  XOR U1248 ( .A(n1711), .B(n1712), .Z(n1699) );
  AND U1249 ( .A(n1713), .B(n1714), .Z(n1712) );
  XOR U1250 ( .A(n1715), .B(n1716), .Z(n1696) );
  AND U1251 ( .A(n1717), .B(n1714), .Z(n1716) );
  XNOR U1252 ( .A(n1715), .B(n1711), .Z(n1714) );
  XOR U1253 ( .A(n1718), .B(n1719), .Z(n1711) );
  AND U1254 ( .A(n1720), .B(n1710), .Z(n1719) );
  XNOR U1255 ( .A(n1721), .B(n1707), .Z(n1710) );
  XOR U1256 ( .A(n1722), .B(n1723), .Z(n1707) );
  AND U1257 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U1258 ( .A(p_input[1401]), .B(n1722), .Z(n1725) );
  XOR U1259 ( .A(n1726), .B(n1727), .Z(n1722) );
  AND U1260 ( .A(n1728), .B(n1729), .Z(n1727) );
  IV U1261 ( .A(n1718), .Z(n1721) );
  XOR U1262 ( .A(n1730), .B(n1731), .Z(n1718) );
  AND U1263 ( .A(n1732), .B(n1733), .Z(n1731) );
  XOR U1264 ( .A(n1734), .B(n1735), .Z(n1715) );
  AND U1265 ( .A(n1736), .B(n1733), .Z(n1735) );
  XNOR U1266 ( .A(n1734), .B(n1730), .Z(n1733) );
  XOR U1267 ( .A(n1737), .B(n1738), .Z(n1730) );
  AND U1268 ( .A(n1739), .B(n1729), .Z(n1738) );
  XNOR U1269 ( .A(n1740), .B(n1726), .Z(n1729) );
  XOR U1270 ( .A(n1741), .B(n1742), .Z(n1726) );
  AND U1271 ( .A(n1743), .B(n1744), .Z(n1742) );
  XOR U1272 ( .A(p_input[1417]), .B(n1741), .Z(n1744) );
  XOR U1273 ( .A(n1745), .B(n1746), .Z(n1741) );
  AND U1274 ( .A(n1747), .B(n1748), .Z(n1746) );
  IV U1275 ( .A(n1737), .Z(n1740) );
  XOR U1276 ( .A(n1749), .B(n1750), .Z(n1737) );
  AND U1277 ( .A(n1751), .B(n1752), .Z(n1750) );
  XOR U1278 ( .A(n1753), .B(n1754), .Z(n1734) );
  AND U1279 ( .A(n1755), .B(n1752), .Z(n1754) );
  XNOR U1280 ( .A(n1753), .B(n1749), .Z(n1752) );
  XOR U1281 ( .A(n1756), .B(n1757), .Z(n1749) );
  AND U1282 ( .A(n1758), .B(n1748), .Z(n1757) );
  XNOR U1283 ( .A(n1759), .B(n1745), .Z(n1748) );
  XOR U1284 ( .A(n1760), .B(n1761), .Z(n1745) );
  AND U1285 ( .A(n1762), .B(n1763), .Z(n1761) );
  XOR U1286 ( .A(p_input[1433]), .B(n1760), .Z(n1763) );
  XOR U1287 ( .A(n1764), .B(n1765), .Z(n1760) );
  AND U1288 ( .A(n1766), .B(n1767), .Z(n1765) );
  IV U1289 ( .A(n1756), .Z(n1759) );
  XOR U1290 ( .A(n1768), .B(n1769), .Z(n1756) );
  AND U1291 ( .A(n1770), .B(n1771), .Z(n1769) );
  XOR U1292 ( .A(n1772), .B(n1773), .Z(n1753) );
  AND U1293 ( .A(n1774), .B(n1771), .Z(n1773) );
  XNOR U1294 ( .A(n1772), .B(n1768), .Z(n1771) );
  XOR U1295 ( .A(n1775), .B(n1776), .Z(n1768) );
  AND U1296 ( .A(n1777), .B(n1767), .Z(n1776) );
  XNOR U1297 ( .A(n1778), .B(n1764), .Z(n1767) );
  XOR U1298 ( .A(n1779), .B(n1780), .Z(n1764) );
  AND U1299 ( .A(n1781), .B(n1782), .Z(n1780) );
  XOR U1300 ( .A(p_input[1449]), .B(n1779), .Z(n1782) );
  XOR U1301 ( .A(n1783), .B(n1784), .Z(n1779) );
  AND U1302 ( .A(n1785), .B(n1786), .Z(n1784) );
  IV U1303 ( .A(n1775), .Z(n1778) );
  XOR U1304 ( .A(n1787), .B(n1788), .Z(n1775) );
  AND U1305 ( .A(n1789), .B(n1790), .Z(n1788) );
  XOR U1306 ( .A(n1791), .B(n1792), .Z(n1772) );
  AND U1307 ( .A(n1793), .B(n1790), .Z(n1792) );
  XNOR U1308 ( .A(n1791), .B(n1787), .Z(n1790) );
  XOR U1309 ( .A(n1794), .B(n1795), .Z(n1787) );
  AND U1310 ( .A(n1796), .B(n1786), .Z(n1795) );
  XNOR U1311 ( .A(n1797), .B(n1783), .Z(n1786) );
  XOR U1312 ( .A(n1798), .B(n1799), .Z(n1783) );
  AND U1313 ( .A(n1800), .B(n1801), .Z(n1799) );
  XOR U1314 ( .A(p_input[1465]), .B(n1798), .Z(n1801) );
  XOR U1315 ( .A(n1802), .B(n1803), .Z(n1798) );
  AND U1316 ( .A(n1804), .B(n1805), .Z(n1803) );
  IV U1317 ( .A(n1794), .Z(n1797) );
  XOR U1318 ( .A(n1806), .B(n1807), .Z(n1794) );
  AND U1319 ( .A(n1808), .B(n1809), .Z(n1807) );
  XOR U1320 ( .A(n1810), .B(n1811), .Z(n1791) );
  AND U1321 ( .A(n1812), .B(n1809), .Z(n1811) );
  XNOR U1322 ( .A(n1810), .B(n1806), .Z(n1809) );
  XOR U1323 ( .A(n1813), .B(n1814), .Z(n1806) );
  AND U1324 ( .A(n1815), .B(n1805), .Z(n1814) );
  XNOR U1325 ( .A(n1816), .B(n1802), .Z(n1805) );
  XOR U1326 ( .A(n1817), .B(n1818), .Z(n1802) );
  AND U1327 ( .A(n1819), .B(n1820), .Z(n1818) );
  XOR U1328 ( .A(p_input[1481]), .B(n1817), .Z(n1820) );
  XOR U1329 ( .A(n1821), .B(n1822), .Z(n1817) );
  AND U1330 ( .A(n1823), .B(n1824), .Z(n1822) );
  IV U1331 ( .A(n1813), .Z(n1816) );
  XOR U1332 ( .A(n1825), .B(n1826), .Z(n1813) );
  AND U1333 ( .A(n1827), .B(n1828), .Z(n1826) );
  XOR U1334 ( .A(n1829), .B(n1830), .Z(n1810) );
  AND U1335 ( .A(n1831), .B(n1828), .Z(n1830) );
  XNOR U1336 ( .A(n1829), .B(n1825), .Z(n1828) );
  XOR U1337 ( .A(n1832), .B(n1833), .Z(n1825) );
  AND U1338 ( .A(n1834), .B(n1824), .Z(n1833) );
  XNOR U1339 ( .A(n1835), .B(n1821), .Z(n1824) );
  XOR U1340 ( .A(n1836), .B(n1837), .Z(n1821) );
  AND U1341 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U1342 ( .A(p_input[1497]), .B(n1836), .Z(n1839) );
  XOR U1343 ( .A(n1840), .B(n1841), .Z(n1836) );
  AND U1344 ( .A(n1842), .B(n1843), .Z(n1841) );
  IV U1345 ( .A(n1832), .Z(n1835) );
  XOR U1346 ( .A(n1844), .B(n1845), .Z(n1832) );
  AND U1347 ( .A(n1846), .B(n1847), .Z(n1845) );
  XOR U1348 ( .A(n1848), .B(n1849), .Z(n1829) );
  AND U1349 ( .A(n1850), .B(n1847), .Z(n1849) );
  XNOR U1350 ( .A(n1848), .B(n1844), .Z(n1847) );
  XOR U1351 ( .A(n1851), .B(n1852), .Z(n1844) );
  AND U1352 ( .A(n1853), .B(n1843), .Z(n1852) );
  XNOR U1353 ( .A(n1854), .B(n1840), .Z(n1843) );
  XOR U1354 ( .A(n1855), .B(n1856), .Z(n1840) );
  AND U1355 ( .A(n1857), .B(n1858), .Z(n1856) );
  XOR U1356 ( .A(p_input[1513]), .B(n1855), .Z(n1858) );
  XOR U1357 ( .A(n1859), .B(n1860), .Z(n1855) );
  AND U1358 ( .A(n1861), .B(n1862), .Z(n1860) );
  IV U1359 ( .A(n1851), .Z(n1854) );
  XOR U1360 ( .A(n1863), .B(n1864), .Z(n1851) );
  AND U1361 ( .A(n1865), .B(n1866), .Z(n1864) );
  XOR U1362 ( .A(n1867), .B(n1868), .Z(n1848) );
  AND U1363 ( .A(n1869), .B(n1866), .Z(n1868) );
  XNOR U1364 ( .A(n1867), .B(n1863), .Z(n1866) );
  XOR U1365 ( .A(n1870), .B(n1871), .Z(n1863) );
  AND U1366 ( .A(n1872), .B(n1862), .Z(n1871) );
  XNOR U1367 ( .A(n1873), .B(n1859), .Z(n1862) );
  XOR U1368 ( .A(n1874), .B(n1875), .Z(n1859) );
  AND U1369 ( .A(n1876), .B(n1877), .Z(n1875) );
  XOR U1370 ( .A(p_input[1529]), .B(n1874), .Z(n1877) );
  XOR U1371 ( .A(n1878), .B(n1879), .Z(n1874) );
  AND U1372 ( .A(n1880), .B(n1881), .Z(n1879) );
  IV U1373 ( .A(n1870), .Z(n1873) );
  XOR U1374 ( .A(n1882), .B(n1883), .Z(n1870) );
  AND U1375 ( .A(n1884), .B(n1885), .Z(n1883) );
  XOR U1376 ( .A(n1886), .B(n1887), .Z(n1867) );
  AND U1377 ( .A(n1888), .B(n1885), .Z(n1887) );
  XNOR U1378 ( .A(n1886), .B(n1882), .Z(n1885) );
  XOR U1379 ( .A(n1889), .B(n1890), .Z(n1882) );
  AND U1380 ( .A(n1891), .B(n1881), .Z(n1890) );
  XNOR U1381 ( .A(n1892), .B(n1878), .Z(n1881) );
  XOR U1382 ( .A(n1893), .B(n1894), .Z(n1878) );
  AND U1383 ( .A(n1895), .B(n1896), .Z(n1894) );
  XOR U1384 ( .A(p_input[1545]), .B(n1893), .Z(n1896) );
  XOR U1385 ( .A(n1897), .B(n1898), .Z(n1893) );
  AND U1386 ( .A(n1899), .B(n1900), .Z(n1898) );
  IV U1387 ( .A(n1889), .Z(n1892) );
  XOR U1388 ( .A(n1901), .B(n1902), .Z(n1889) );
  AND U1389 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U1390 ( .A(n1905), .B(n1906), .Z(n1886) );
  AND U1391 ( .A(n1907), .B(n1904), .Z(n1906) );
  XNOR U1392 ( .A(n1905), .B(n1901), .Z(n1904) );
  XOR U1393 ( .A(n1908), .B(n1909), .Z(n1901) );
  AND U1394 ( .A(n1910), .B(n1900), .Z(n1909) );
  XNOR U1395 ( .A(n1911), .B(n1897), .Z(n1900) );
  XOR U1396 ( .A(n1912), .B(n1913), .Z(n1897) );
  AND U1397 ( .A(n1914), .B(n1915), .Z(n1913) );
  XOR U1398 ( .A(p_input[1561]), .B(n1912), .Z(n1915) );
  XOR U1399 ( .A(n1916), .B(n1917), .Z(n1912) );
  AND U1400 ( .A(n1918), .B(n1919), .Z(n1917) );
  IV U1401 ( .A(n1908), .Z(n1911) );
  XOR U1402 ( .A(n1920), .B(n1921), .Z(n1908) );
  AND U1403 ( .A(n1922), .B(n1923), .Z(n1921) );
  XOR U1404 ( .A(n1924), .B(n1925), .Z(n1905) );
  AND U1405 ( .A(n1926), .B(n1923), .Z(n1925) );
  XNOR U1406 ( .A(n1924), .B(n1920), .Z(n1923) );
  XOR U1407 ( .A(n1927), .B(n1928), .Z(n1920) );
  AND U1408 ( .A(n1929), .B(n1919), .Z(n1928) );
  XNOR U1409 ( .A(n1930), .B(n1916), .Z(n1919) );
  XOR U1410 ( .A(n1931), .B(n1932), .Z(n1916) );
  AND U1411 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U1412 ( .A(p_input[1577]), .B(n1931), .Z(n1934) );
  XOR U1413 ( .A(n1935), .B(n1936), .Z(n1931) );
  AND U1414 ( .A(n1937), .B(n1938), .Z(n1936) );
  IV U1415 ( .A(n1927), .Z(n1930) );
  XOR U1416 ( .A(n1939), .B(n1940), .Z(n1927) );
  AND U1417 ( .A(n1941), .B(n1942), .Z(n1940) );
  XOR U1418 ( .A(n1943), .B(n1944), .Z(n1924) );
  AND U1419 ( .A(n1945), .B(n1942), .Z(n1944) );
  XNOR U1420 ( .A(n1943), .B(n1939), .Z(n1942) );
  XOR U1421 ( .A(n1946), .B(n1947), .Z(n1939) );
  AND U1422 ( .A(n1948), .B(n1938), .Z(n1947) );
  XNOR U1423 ( .A(n1949), .B(n1935), .Z(n1938) );
  XOR U1424 ( .A(n1950), .B(n1951), .Z(n1935) );
  AND U1425 ( .A(n1952), .B(n1953), .Z(n1951) );
  XOR U1426 ( .A(p_input[1593]), .B(n1950), .Z(n1953) );
  XOR U1427 ( .A(n1954), .B(n1955), .Z(n1950) );
  AND U1428 ( .A(n1956), .B(n1957), .Z(n1955) );
  IV U1429 ( .A(n1946), .Z(n1949) );
  XOR U1430 ( .A(n1958), .B(n1959), .Z(n1946) );
  AND U1431 ( .A(n1960), .B(n1961), .Z(n1959) );
  XOR U1432 ( .A(n1962), .B(n1963), .Z(n1943) );
  AND U1433 ( .A(n1964), .B(n1961), .Z(n1963) );
  XNOR U1434 ( .A(n1962), .B(n1958), .Z(n1961) );
  XOR U1435 ( .A(n1965), .B(n1966), .Z(n1958) );
  AND U1436 ( .A(n1967), .B(n1957), .Z(n1966) );
  XNOR U1437 ( .A(n1968), .B(n1954), .Z(n1957) );
  XOR U1438 ( .A(n1969), .B(n1970), .Z(n1954) );
  AND U1439 ( .A(n1971), .B(n1972), .Z(n1970) );
  XOR U1440 ( .A(p_input[1609]), .B(n1969), .Z(n1972) );
  XOR U1441 ( .A(n1973), .B(n1974), .Z(n1969) );
  AND U1442 ( .A(n1975), .B(n1976), .Z(n1974) );
  IV U1443 ( .A(n1965), .Z(n1968) );
  XOR U1444 ( .A(n1977), .B(n1978), .Z(n1965) );
  AND U1445 ( .A(n1979), .B(n1980), .Z(n1978) );
  XOR U1446 ( .A(n1981), .B(n1982), .Z(n1962) );
  AND U1447 ( .A(n1983), .B(n1980), .Z(n1982) );
  XNOR U1448 ( .A(n1981), .B(n1977), .Z(n1980) );
  XOR U1449 ( .A(n1984), .B(n1985), .Z(n1977) );
  AND U1450 ( .A(n1986), .B(n1976), .Z(n1985) );
  XNOR U1451 ( .A(n1987), .B(n1973), .Z(n1976) );
  XOR U1452 ( .A(n1988), .B(n1989), .Z(n1973) );
  AND U1453 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U1454 ( .A(p_input[1625]), .B(n1988), .Z(n1991) );
  XOR U1455 ( .A(n1992), .B(n1993), .Z(n1988) );
  AND U1456 ( .A(n1994), .B(n1995), .Z(n1993) );
  IV U1457 ( .A(n1984), .Z(n1987) );
  XOR U1458 ( .A(n1996), .B(n1997), .Z(n1984) );
  AND U1459 ( .A(n1998), .B(n1999), .Z(n1997) );
  XOR U1460 ( .A(n2000), .B(n2001), .Z(n1981) );
  AND U1461 ( .A(n2002), .B(n1999), .Z(n2001) );
  XNOR U1462 ( .A(n2000), .B(n1996), .Z(n1999) );
  XOR U1463 ( .A(n2003), .B(n2004), .Z(n1996) );
  AND U1464 ( .A(n2005), .B(n1995), .Z(n2004) );
  XNOR U1465 ( .A(n2006), .B(n1992), .Z(n1995) );
  XOR U1466 ( .A(n2007), .B(n2008), .Z(n1992) );
  AND U1467 ( .A(n2009), .B(n2010), .Z(n2008) );
  XOR U1468 ( .A(p_input[1641]), .B(n2007), .Z(n2010) );
  XOR U1469 ( .A(n2011), .B(n2012), .Z(n2007) );
  AND U1470 ( .A(n2013), .B(n2014), .Z(n2012) );
  IV U1471 ( .A(n2003), .Z(n2006) );
  XOR U1472 ( .A(n2015), .B(n2016), .Z(n2003) );
  AND U1473 ( .A(n2017), .B(n2018), .Z(n2016) );
  XOR U1474 ( .A(n2019), .B(n2020), .Z(n2000) );
  AND U1475 ( .A(n2021), .B(n2018), .Z(n2020) );
  XNOR U1476 ( .A(n2019), .B(n2015), .Z(n2018) );
  XOR U1477 ( .A(n2022), .B(n2023), .Z(n2015) );
  AND U1478 ( .A(n2024), .B(n2014), .Z(n2023) );
  XNOR U1479 ( .A(n2025), .B(n2011), .Z(n2014) );
  XOR U1480 ( .A(n2026), .B(n2027), .Z(n2011) );
  AND U1481 ( .A(n2028), .B(n2029), .Z(n2027) );
  XOR U1482 ( .A(p_input[1657]), .B(n2026), .Z(n2029) );
  XOR U1483 ( .A(n2030), .B(n2031), .Z(n2026) );
  AND U1484 ( .A(n2032), .B(n2033), .Z(n2031) );
  IV U1485 ( .A(n2022), .Z(n2025) );
  XOR U1486 ( .A(n2034), .B(n2035), .Z(n2022) );
  AND U1487 ( .A(n2036), .B(n2037), .Z(n2035) );
  XOR U1488 ( .A(n2038), .B(n2039), .Z(n2019) );
  AND U1489 ( .A(n2040), .B(n2037), .Z(n2039) );
  XNOR U1490 ( .A(n2038), .B(n2034), .Z(n2037) );
  XOR U1491 ( .A(n2041), .B(n2042), .Z(n2034) );
  AND U1492 ( .A(n2043), .B(n2033), .Z(n2042) );
  XNOR U1493 ( .A(n2044), .B(n2030), .Z(n2033) );
  XOR U1494 ( .A(n2045), .B(n2046), .Z(n2030) );
  AND U1495 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U1496 ( .A(p_input[1673]), .B(n2045), .Z(n2048) );
  XOR U1497 ( .A(n2049), .B(n2050), .Z(n2045) );
  AND U1498 ( .A(n2051), .B(n2052), .Z(n2050) );
  IV U1499 ( .A(n2041), .Z(n2044) );
  XOR U1500 ( .A(n2053), .B(n2054), .Z(n2041) );
  AND U1501 ( .A(n2055), .B(n2056), .Z(n2054) );
  XOR U1502 ( .A(n2057), .B(n2058), .Z(n2038) );
  AND U1503 ( .A(n2059), .B(n2056), .Z(n2058) );
  XNOR U1504 ( .A(n2057), .B(n2053), .Z(n2056) );
  XOR U1505 ( .A(n2060), .B(n2061), .Z(n2053) );
  AND U1506 ( .A(n2062), .B(n2052), .Z(n2061) );
  XNOR U1507 ( .A(n2063), .B(n2049), .Z(n2052) );
  XOR U1508 ( .A(n2064), .B(n2065), .Z(n2049) );
  AND U1509 ( .A(n2066), .B(n2067), .Z(n2065) );
  XOR U1510 ( .A(p_input[1689]), .B(n2064), .Z(n2067) );
  XOR U1511 ( .A(n2068), .B(n2069), .Z(n2064) );
  AND U1512 ( .A(n2070), .B(n2071), .Z(n2069) );
  IV U1513 ( .A(n2060), .Z(n2063) );
  XOR U1514 ( .A(n2072), .B(n2073), .Z(n2060) );
  AND U1515 ( .A(n2074), .B(n2075), .Z(n2073) );
  XOR U1516 ( .A(n2076), .B(n2077), .Z(n2057) );
  AND U1517 ( .A(n2078), .B(n2075), .Z(n2077) );
  XNOR U1518 ( .A(n2076), .B(n2072), .Z(n2075) );
  XOR U1519 ( .A(n2079), .B(n2080), .Z(n2072) );
  AND U1520 ( .A(n2081), .B(n2071), .Z(n2080) );
  XNOR U1521 ( .A(n2082), .B(n2068), .Z(n2071) );
  XOR U1522 ( .A(n2083), .B(n2084), .Z(n2068) );
  AND U1523 ( .A(n2085), .B(n2086), .Z(n2084) );
  XOR U1524 ( .A(p_input[1705]), .B(n2083), .Z(n2086) );
  XOR U1525 ( .A(n2087), .B(n2088), .Z(n2083) );
  AND U1526 ( .A(n2089), .B(n2090), .Z(n2088) );
  IV U1527 ( .A(n2079), .Z(n2082) );
  XOR U1528 ( .A(n2091), .B(n2092), .Z(n2079) );
  AND U1529 ( .A(n2093), .B(n2094), .Z(n2092) );
  XOR U1530 ( .A(n2095), .B(n2096), .Z(n2076) );
  AND U1531 ( .A(n2097), .B(n2094), .Z(n2096) );
  XNOR U1532 ( .A(n2095), .B(n2091), .Z(n2094) );
  XOR U1533 ( .A(n2098), .B(n2099), .Z(n2091) );
  AND U1534 ( .A(n2100), .B(n2090), .Z(n2099) );
  XNOR U1535 ( .A(n2101), .B(n2087), .Z(n2090) );
  XOR U1536 ( .A(n2102), .B(n2103), .Z(n2087) );
  AND U1537 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR U1538 ( .A(p_input[1721]), .B(n2102), .Z(n2105) );
  XOR U1539 ( .A(n2106), .B(n2107), .Z(n2102) );
  AND U1540 ( .A(n2108), .B(n2109), .Z(n2107) );
  IV U1541 ( .A(n2098), .Z(n2101) );
  XOR U1542 ( .A(n2110), .B(n2111), .Z(n2098) );
  AND U1543 ( .A(n2112), .B(n2113), .Z(n2111) );
  XOR U1544 ( .A(n2114), .B(n2115), .Z(n2095) );
  AND U1545 ( .A(n2116), .B(n2113), .Z(n2115) );
  XNOR U1546 ( .A(n2114), .B(n2110), .Z(n2113) );
  XOR U1547 ( .A(n2117), .B(n2118), .Z(n2110) );
  AND U1548 ( .A(n2119), .B(n2109), .Z(n2118) );
  XNOR U1549 ( .A(n2120), .B(n2106), .Z(n2109) );
  XOR U1550 ( .A(n2121), .B(n2122), .Z(n2106) );
  AND U1551 ( .A(n2123), .B(n2124), .Z(n2122) );
  XOR U1552 ( .A(p_input[1737]), .B(n2121), .Z(n2124) );
  XOR U1553 ( .A(n2125), .B(n2126), .Z(n2121) );
  AND U1554 ( .A(n2127), .B(n2128), .Z(n2126) );
  IV U1555 ( .A(n2117), .Z(n2120) );
  XOR U1556 ( .A(n2129), .B(n2130), .Z(n2117) );
  AND U1557 ( .A(n2131), .B(n2132), .Z(n2130) );
  XOR U1558 ( .A(n2133), .B(n2134), .Z(n2114) );
  AND U1559 ( .A(n2135), .B(n2132), .Z(n2134) );
  XNOR U1560 ( .A(n2133), .B(n2129), .Z(n2132) );
  XOR U1561 ( .A(n2136), .B(n2137), .Z(n2129) );
  AND U1562 ( .A(n2138), .B(n2128), .Z(n2137) );
  XNOR U1563 ( .A(n2139), .B(n2125), .Z(n2128) );
  XOR U1564 ( .A(n2140), .B(n2141), .Z(n2125) );
  AND U1565 ( .A(n2142), .B(n2143), .Z(n2141) );
  XOR U1566 ( .A(p_input[1753]), .B(n2140), .Z(n2143) );
  XOR U1567 ( .A(n2144), .B(n2145), .Z(n2140) );
  AND U1568 ( .A(n2146), .B(n2147), .Z(n2145) );
  IV U1569 ( .A(n2136), .Z(n2139) );
  XOR U1570 ( .A(n2148), .B(n2149), .Z(n2136) );
  AND U1571 ( .A(n2150), .B(n2151), .Z(n2149) );
  XOR U1572 ( .A(n2152), .B(n2153), .Z(n2133) );
  AND U1573 ( .A(n2154), .B(n2151), .Z(n2153) );
  XNOR U1574 ( .A(n2152), .B(n2148), .Z(n2151) );
  XOR U1575 ( .A(n2155), .B(n2156), .Z(n2148) );
  AND U1576 ( .A(n2157), .B(n2147), .Z(n2156) );
  XNOR U1577 ( .A(n2158), .B(n2144), .Z(n2147) );
  XOR U1578 ( .A(n2159), .B(n2160), .Z(n2144) );
  AND U1579 ( .A(n2161), .B(n2162), .Z(n2160) );
  XOR U1580 ( .A(p_input[1769]), .B(n2159), .Z(n2162) );
  XOR U1581 ( .A(n2163), .B(n2164), .Z(n2159) );
  AND U1582 ( .A(n2165), .B(n2166), .Z(n2164) );
  IV U1583 ( .A(n2155), .Z(n2158) );
  XOR U1584 ( .A(n2167), .B(n2168), .Z(n2155) );
  AND U1585 ( .A(n2169), .B(n2170), .Z(n2168) );
  XOR U1586 ( .A(n2171), .B(n2172), .Z(n2152) );
  AND U1587 ( .A(n2173), .B(n2170), .Z(n2172) );
  XNOR U1588 ( .A(n2171), .B(n2167), .Z(n2170) );
  XOR U1589 ( .A(n2174), .B(n2175), .Z(n2167) );
  AND U1590 ( .A(n2176), .B(n2166), .Z(n2175) );
  XNOR U1591 ( .A(n2177), .B(n2163), .Z(n2166) );
  XOR U1592 ( .A(n2178), .B(n2179), .Z(n2163) );
  AND U1593 ( .A(n2180), .B(n2181), .Z(n2179) );
  XOR U1594 ( .A(p_input[1785]), .B(n2178), .Z(n2181) );
  XOR U1595 ( .A(n2182), .B(n2183), .Z(n2178) );
  AND U1596 ( .A(n2184), .B(n2185), .Z(n2183) );
  IV U1597 ( .A(n2174), .Z(n2177) );
  XOR U1598 ( .A(n2186), .B(n2187), .Z(n2174) );
  AND U1599 ( .A(n2188), .B(n2189), .Z(n2187) );
  XOR U1600 ( .A(n2190), .B(n2191), .Z(n2171) );
  AND U1601 ( .A(n2192), .B(n2189), .Z(n2191) );
  XNOR U1602 ( .A(n2190), .B(n2186), .Z(n2189) );
  XOR U1603 ( .A(n2193), .B(n2194), .Z(n2186) );
  AND U1604 ( .A(n2195), .B(n2185), .Z(n2194) );
  XNOR U1605 ( .A(n2196), .B(n2182), .Z(n2185) );
  XOR U1606 ( .A(n2197), .B(n2198), .Z(n2182) );
  AND U1607 ( .A(n2199), .B(n2200), .Z(n2198) );
  XOR U1608 ( .A(p_input[1801]), .B(n2197), .Z(n2200) );
  XOR U1609 ( .A(n2201), .B(n2202), .Z(n2197) );
  AND U1610 ( .A(n2203), .B(n2204), .Z(n2202) );
  IV U1611 ( .A(n2193), .Z(n2196) );
  XOR U1612 ( .A(n2205), .B(n2206), .Z(n2193) );
  AND U1613 ( .A(n2207), .B(n2208), .Z(n2206) );
  XOR U1614 ( .A(n2209), .B(n2210), .Z(n2190) );
  AND U1615 ( .A(n2211), .B(n2208), .Z(n2210) );
  XNOR U1616 ( .A(n2209), .B(n2205), .Z(n2208) );
  XOR U1617 ( .A(n2212), .B(n2213), .Z(n2205) );
  AND U1618 ( .A(n2214), .B(n2204), .Z(n2213) );
  XNOR U1619 ( .A(n2215), .B(n2201), .Z(n2204) );
  XOR U1620 ( .A(n2216), .B(n2217), .Z(n2201) );
  AND U1621 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U1622 ( .A(p_input[1817]), .B(n2216), .Z(n2219) );
  XOR U1623 ( .A(n2220), .B(n2221), .Z(n2216) );
  AND U1624 ( .A(n2222), .B(n2223), .Z(n2221) );
  IV U1625 ( .A(n2212), .Z(n2215) );
  XOR U1626 ( .A(n2224), .B(n2225), .Z(n2212) );
  AND U1627 ( .A(n2226), .B(n2227), .Z(n2225) );
  XOR U1628 ( .A(n2228), .B(n2229), .Z(n2209) );
  AND U1629 ( .A(n2230), .B(n2227), .Z(n2229) );
  XNOR U1630 ( .A(n2228), .B(n2224), .Z(n2227) );
  XOR U1631 ( .A(n2231), .B(n2232), .Z(n2224) );
  AND U1632 ( .A(n2233), .B(n2223), .Z(n2232) );
  XNOR U1633 ( .A(n2234), .B(n2220), .Z(n2223) );
  XOR U1634 ( .A(n2235), .B(n2236), .Z(n2220) );
  AND U1635 ( .A(n2237), .B(n2238), .Z(n2236) );
  XOR U1636 ( .A(p_input[1833]), .B(n2235), .Z(n2238) );
  XOR U1637 ( .A(n2239), .B(n2240), .Z(n2235) );
  AND U1638 ( .A(n2241), .B(n2242), .Z(n2240) );
  IV U1639 ( .A(n2231), .Z(n2234) );
  XOR U1640 ( .A(n2243), .B(n2244), .Z(n2231) );
  AND U1641 ( .A(n2245), .B(n2246), .Z(n2244) );
  XOR U1642 ( .A(n2247), .B(n2248), .Z(n2228) );
  AND U1643 ( .A(n2249), .B(n2246), .Z(n2248) );
  XNOR U1644 ( .A(n2247), .B(n2243), .Z(n2246) );
  XOR U1645 ( .A(n2250), .B(n2251), .Z(n2243) );
  AND U1646 ( .A(n2252), .B(n2242), .Z(n2251) );
  XNOR U1647 ( .A(n2253), .B(n2239), .Z(n2242) );
  XOR U1648 ( .A(n2254), .B(n2255), .Z(n2239) );
  AND U1649 ( .A(n2256), .B(n2257), .Z(n2255) );
  XOR U1650 ( .A(p_input[1849]), .B(n2254), .Z(n2257) );
  XOR U1651 ( .A(n2258), .B(n2259), .Z(n2254) );
  AND U1652 ( .A(n2260), .B(n2261), .Z(n2259) );
  IV U1653 ( .A(n2250), .Z(n2253) );
  XOR U1654 ( .A(n2262), .B(n2263), .Z(n2250) );
  AND U1655 ( .A(n2264), .B(n2265), .Z(n2263) );
  XOR U1656 ( .A(n2266), .B(n2267), .Z(n2247) );
  AND U1657 ( .A(n2268), .B(n2265), .Z(n2267) );
  XNOR U1658 ( .A(n2266), .B(n2262), .Z(n2265) );
  XOR U1659 ( .A(n2269), .B(n2270), .Z(n2262) );
  AND U1660 ( .A(n2271), .B(n2261), .Z(n2270) );
  XNOR U1661 ( .A(n2272), .B(n2258), .Z(n2261) );
  XOR U1662 ( .A(n2273), .B(n2274), .Z(n2258) );
  AND U1663 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U1664 ( .A(p_input[1865]), .B(n2273), .Z(n2276) );
  XOR U1665 ( .A(n2277), .B(n2278), .Z(n2273) );
  AND U1666 ( .A(n2279), .B(n2280), .Z(n2278) );
  IV U1667 ( .A(n2269), .Z(n2272) );
  XOR U1668 ( .A(n2281), .B(n2282), .Z(n2269) );
  AND U1669 ( .A(n2283), .B(n2284), .Z(n2282) );
  XOR U1670 ( .A(n2285), .B(n2286), .Z(n2266) );
  AND U1671 ( .A(n2287), .B(n2284), .Z(n2286) );
  XNOR U1672 ( .A(n2285), .B(n2281), .Z(n2284) );
  XOR U1673 ( .A(n2288), .B(n2289), .Z(n2281) );
  AND U1674 ( .A(n2290), .B(n2280), .Z(n2289) );
  XNOR U1675 ( .A(n2291), .B(n2277), .Z(n2280) );
  XOR U1676 ( .A(n2292), .B(n2293), .Z(n2277) );
  AND U1677 ( .A(n2294), .B(n2295), .Z(n2293) );
  XOR U1678 ( .A(p_input[1881]), .B(n2292), .Z(n2295) );
  XOR U1679 ( .A(n2296), .B(n2297), .Z(n2292) );
  AND U1680 ( .A(n2298), .B(n2299), .Z(n2297) );
  IV U1681 ( .A(n2288), .Z(n2291) );
  XOR U1682 ( .A(n2300), .B(n2301), .Z(n2288) );
  AND U1683 ( .A(n2302), .B(n2303), .Z(n2301) );
  XOR U1684 ( .A(n2304), .B(n2305), .Z(n2285) );
  AND U1685 ( .A(n2306), .B(n2303), .Z(n2305) );
  XNOR U1686 ( .A(n2304), .B(n2300), .Z(n2303) );
  XOR U1687 ( .A(n2307), .B(n2308), .Z(n2300) );
  AND U1688 ( .A(n2309), .B(n2299), .Z(n2308) );
  XNOR U1689 ( .A(n2310), .B(n2296), .Z(n2299) );
  XOR U1690 ( .A(n2311), .B(n2312), .Z(n2296) );
  AND U1691 ( .A(n2313), .B(n2314), .Z(n2312) );
  XOR U1692 ( .A(p_input[1897]), .B(n2311), .Z(n2314) );
  XOR U1693 ( .A(n2315), .B(n2316), .Z(n2311) );
  AND U1694 ( .A(n2317), .B(n2318), .Z(n2316) );
  IV U1695 ( .A(n2307), .Z(n2310) );
  XOR U1696 ( .A(n2319), .B(n2320), .Z(n2307) );
  AND U1697 ( .A(n2321), .B(n2322), .Z(n2320) );
  XOR U1698 ( .A(n2323), .B(n2324), .Z(n2304) );
  AND U1699 ( .A(n2325), .B(n2322), .Z(n2324) );
  XNOR U1700 ( .A(n2323), .B(n2319), .Z(n2322) );
  XOR U1701 ( .A(n2326), .B(n2327), .Z(n2319) );
  AND U1702 ( .A(n2328), .B(n2318), .Z(n2327) );
  XNOR U1703 ( .A(n2329), .B(n2315), .Z(n2318) );
  XOR U1704 ( .A(n2330), .B(n2331), .Z(n2315) );
  AND U1705 ( .A(n2332), .B(n2333), .Z(n2331) );
  XOR U1706 ( .A(p_input[1913]), .B(n2330), .Z(n2333) );
  XOR U1707 ( .A(n2334), .B(n2335), .Z(n2330) );
  AND U1708 ( .A(n2336), .B(n2337), .Z(n2335) );
  IV U1709 ( .A(n2326), .Z(n2329) );
  XOR U1710 ( .A(n2338), .B(n2339), .Z(n2326) );
  AND U1711 ( .A(n2340), .B(n2341), .Z(n2339) );
  XOR U1712 ( .A(n2342), .B(n2343), .Z(n2323) );
  AND U1713 ( .A(n2344), .B(n2341), .Z(n2343) );
  XNOR U1714 ( .A(n2342), .B(n2338), .Z(n2341) );
  XOR U1715 ( .A(n2345), .B(n2346), .Z(n2338) );
  AND U1716 ( .A(n2347), .B(n2337), .Z(n2346) );
  XNOR U1717 ( .A(n2348), .B(n2334), .Z(n2337) );
  XOR U1718 ( .A(n2349), .B(n2350), .Z(n2334) );
  AND U1719 ( .A(n2351), .B(n2352), .Z(n2350) );
  XOR U1720 ( .A(p_input[1929]), .B(n2349), .Z(n2352) );
  XOR U1721 ( .A(n2353), .B(n2354), .Z(n2349) );
  AND U1722 ( .A(n2355), .B(n2356), .Z(n2354) );
  IV U1723 ( .A(n2345), .Z(n2348) );
  XOR U1724 ( .A(n2357), .B(n2358), .Z(n2345) );
  AND U1725 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U1726 ( .A(n2361), .B(n2362), .Z(n2342) );
  AND U1727 ( .A(n2363), .B(n2360), .Z(n2362) );
  XNOR U1728 ( .A(n2361), .B(n2357), .Z(n2360) );
  XOR U1729 ( .A(n2364), .B(n2365), .Z(n2357) );
  AND U1730 ( .A(n2366), .B(n2356), .Z(n2365) );
  XNOR U1731 ( .A(n2367), .B(n2353), .Z(n2356) );
  XOR U1732 ( .A(n2368), .B(n2369), .Z(n2353) );
  AND U1733 ( .A(n2370), .B(n2371), .Z(n2369) );
  XOR U1734 ( .A(p_input[1945]), .B(n2368), .Z(n2371) );
  XOR U1735 ( .A(n2372), .B(n2373), .Z(n2368) );
  AND U1736 ( .A(n2374), .B(n2375), .Z(n2373) );
  IV U1737 ( .A(n2364), .Z(n2367) );
  XOR U1738 ( .A(n2376), .B(n2377), .Z(n2364) );
  AND U1739 ( .A(n2378), .B(n2379), .Z(n2377) );
  XOR U1740 ( .A(n2380), .B(n2381), .Z(n2361) );
  AND U1741 ( .A(n2382), .B(n2379), .Z(n2381) );
  XNOR U1742 ( .A(n2380), .B(n2376), .Z(n2379) );
  XOR U1743 ( .A(n2383), .B(n2384), .Z(n2376) );
  AND U1744 ( .A(n2385), .B(n2375), .Z(n2384) );
  XNOR U1745 ( .A(n2386), .B(n2372), .Z(n2375) );
  XOR U1746 ( .A(n2387), .B(n2388), .Z(n2372) );
  AND U1747 ( .A(n2389), .B(n2390), .Z(n2388) );
  XOR U1748 ( .A(p_input[1961]), .B(n2387), .Z(n2390) );
  XOR U1749 ( .A(n2391), .B(n2392), .Z(n2387) );
  AND U1750 ( .A(n2393), .B(n2394), .Z(n2392) );
  IV U1751 ( .A(n2383), .Z(n2386) );
  XOR U1752 ( .A(n2395), .B(n2396), .Z(n2383) );
  AND U1753 ( .A(n2397), .B(n2398), .Z(n2396) );
  XOR U1754 ( .A(n2399), .B(n2400), .Z(n2380) );
  AND U1755 ( .A(n2401), .B(n2398), .Z(n2400) );
  XNOR U1756 ( .A(n2399), .B(n2395), .Z(n2398) );
  XOR U1757 ( .A(n2402), .B(n2403), .Z(n2395) );
  AND U1758 ( .A(n2404), .B(n2394), .Z(n2403) );
  XNOR U1759 ( .A(n2405), .B(n2391), .Z(n2394) );
  XOR U1760 ( .A(n2406), .B(n2407), .Z(n2391) );
  AND U1761 ( .A(n2408), .B(n2409), .Z(n2407) );
  XOR U1762 ( .A(p_input[1977]), .B(n2406), .Z(n2409) );
  XOR U1763 ( .A(n2410), .B(n2411), .Z(n2406) );
  AND U1764 ( .A(n2412), .B(n2413), .Z(n2411) );
  IV U1765 ( .A(n2402), .Z(n2405) );
  XOR U1766 ( .A(n2414), .B(n2415), .Z(n2402) );
  AND U1767 ( .A(n2416), .B(n2417), .Z(n2415) );
  XOR U1768 ( .A(n2418), .B(n2419), .Z(n2399) );
  AND U1769 ( .A(n2420), .B(n2417), .Z(n2419) );
  XNOR U1770 ( .A(n2418), .B(n2414), .Z(n2417) );
  XOR U1771 ( .A(n2421), .B(n2422), .Z(n2414) );
  AND U1772 ( .A(n2423), .B(n2413), .Z(n2422) );
  XNOR U1773 ( .A(n2424), .B(n2410), .Z(n2413) );
  XOR U1774 ( .A(n2425), .B(n2426), .Z(n2410) );
  AND U1775 ( .A(n2427), .B(n2428), .Z(n2426) );
  XOR U1776 ( .A(p_input[1993]), .B(n2425), .Z(n2428) );
  XOR U1777 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n2429), 
        .Z(n2425) );
  AND U1778 ( .A(n2430), .B(n2431), .Z(n2429) );
  IV U1779 ( .A(n2421), .Z(n2424) );
  XOR U1780 ( .A(n2432), .B(n2433), .Z(n2421) );
  AND U1781 ( .A(n2434), .B(n2435), .Z(n2433) );
  XOR U1782 ( .A(n2436), .B(n2437), .Z(n2418) );
  AND U1783 ( .A(n2438), .B(n2435), .Z(n2437) );
  XNOR U1784 ( .A(n2436), .B(n2432), .Z(n2435) );
  XNOR U1785 ( .A(n2439), .B(n2440), .Z(n2432) );
  AND U1786 ( .A(n2441), .B(n2431), .Z(n2440) );
  XNOR U1787 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n2439), 
        .Z(n2431) );
  XNOR U1788 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n2442), 
        .Z(n2439) );
  AND U1789 ( .A(n2443), .B(n2444), .Z(n2442) );
  XNOR U1790 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n2445), .Z(n2436) );
  AND U1791 ( .A(n2446), .B(n2444), .Z(n2445) );
  XOR U1792 ( .A(n2447), .B(n2448), .Z(n2444) );
  XOR U1793 ( .A(n3), .B(n2449), .Z(o[24]) );
  AND U1794 ( .A(n62), .B(n2450), .Z(n3) );
  XOR U1795 ( .A(n4), .B(n2449), .Z(n2450) );
  XOR U1796 ( .A(n2451), .B(n27), .Z(n2449) );
  AND U1797 ( .A(n65), .B(n2452), .Z(n27) );
  XNOR U1798 ( .A(n2453), .B(n28), .Z(n2452) );
  XOR U1799 ( .A(n2454), .B(n2455), .Z(n28) );
  AND U1800 ( .A(n70), .B(n2456), .Z(n2455) );
  XOR U1801 ( .A(p_input[8]), .B(n2454), .Z(n2456) );
  XOR U1802 ( .A(n2457), .B(n2458), .Z(n2454) );
  AND U1803 ( .A(n74), .B(n2459), .Z(n2458) );
  IV U1804 ( .A(n2451), .Z(n2453) );
  XOR U1805 ( .A(n2460), .B(n2461), .Z(n2451) );
  AND U1806 ( .A(n78), .B(n2462), .Z(n2461) );
  XOR U1807 ( .A(n2463), .B(n2464), .Z(n4) );
  AND U1808 ( .A(n82), .B(n2462), .Z(n2464) );
  XNOR U1809 ( .A(n2465), .B(n2460), .Z(n2462) );
  XOR U1810 ( .A(n2466), .B(n2467), .Z(n2460) );
  AND U1811 ( .A(n86), .B(n2459), .Z(n2467) );
  XNOR U1812 ( .A(n2468), .B(n2457), .Z(n2459) );
  XOR U1813 ( .A(n2469), .B(n2470), .Z(n2457) );
  AND U1814 ( .A(n90), .B(n2471), .Z(n2470) );
  XOR U1815 ( .A(p_input[24]), .B(n2469), .Z(n2471) );
  XOR U1816 ( .A(n2472), .B(n2473), .Z(n2469) );
  AND U1817 ( .A(n94), .B(n2474), .Z(n2473) );
  IV U1818 ( .A(n2466), .Z(n2468) );
  XOR U1819 ( .A(n2475), .B(n2476), .Z(n2466) );
  AND U1820 ( .A(n98), .B(n2477), .Z(n2476) );
  IV U1821 ( .A(n2463), .Z(n2465) );
  XNOR U1822 ( .A(n2478), .B(n2479), .Z(n2463) );
  AND U1823 ( .A(n102), .B(n2477), .Z(n2479) );
  XNOR U1824 ( .A(n2478), .B(n2475), .Z(n2477) );
  XOR U1825 ( .A(n2480), .B(n2481), .Z(n2475) );
  AND U1826 ( .A(n105), .B(n2474), .Z(n2481) );
  XNOR U1827 ( .A(n2482), .B(n2472), .Z(n2474) );
  XOR U1828 ( .A(n2483), .B(n2484), .Z(n2472) );
  AND U1829 ( .A(n109), .B(n2485), .Z(n2484) );
  XOR U1830 ( .A(p_input[40]), .B(n2483), .Z(n2485) );
  XOR U1831 ( .A(n2486), .B(n2487), .Z(n2483) );
  AND U1832 ( .A(n113), .B(n2488), .Z(n2487) );
  IV U1833 ( .A(n2480), .Z(n2482) );
  XOR U1834 ( .A(n2489), .B(n2490), .Z(n2480) );
  AND U1835 ( .A(n117), .B(n2491), .Z(n2490) );
  XOR U1836 ( .A(n2492), .B(n2493), .Z(n2478) );
  AND U1837 ( .A(n121), .B(n2491), .Z(n2493) );
  XNOR U1838 ( .A(n2492), .B(n2489), .Z(n2491) );
  XOR U1839 ( .A(n2494), .B(n2495), .Z(n2489) );
  AND U1840 ( .A(n124), .B(n2488), .Z(n2495) );
  XNOR U1841 ( .A(n2496), .B(n2486), .Z(n2488) );
  XOR U1842 ( .A(n2497), .B(n2498), .Z(n2486) );
  AND U1843 ( .A(n128), .B(n2499), .Z(n2498) );
  XOR U1844 ( .A(p_input[56]), .B(n2497), .Z(n2499) );
  XOR U1845 ( .A(n2500), .B(n2501), .Z(n2497) );
  AND U1846 ( .A(n132), .B(n2502), .Z(n2501) );
  IV U1847 ( .A(n2494), .Z(n2496) );
  XOR U1848 ( .A(n2503), .B(n2504), .Z(n2494) );
  AND U1849 ( .A(n136), .B(n2505), .Z(n2504) );
  XOR U1850 ( .A(n2506), .B(n2507), .Z(n2492) );
  AND U1851 ( .A(n140), .B(n2505), .Z(n2507) );
  XNOR U1852 ( .A(n2506), .B(n2503), .Z(n2505) );
  XOR U1853 ( .A(n2508), .B(n2509), .Z(n2503) );
  AND U1854 ( .A(n143), .B(n2502), .Z(n2509) );
  XNOR U1855 ( .A(n2510), .B(n2500), .Z(n2502) );
  XOR U1856 ( .A(n2511), .B(n2512), .Z(n2500) );
  AND U1857 ( .A(n147), .B(n2513), .Z(n2512) );
  XOR U1858 ( .A(p_input[72]), .B(n2511), .Z(n2513) );
  XOR U1859 ( .A(n2514), .B(n2515), .Z(n2511) );
  AND U1860 ( .A(n151), .B(n2516), .Z(n2515) );
  IV U1861 ( .A(n2508), .Z(n2510) );
  XOR U1862 ( .A(n2517), .B(n2518), .Z(n2508) );
  AND U1863 ( .A(n155), .B(n2519), .Z(n2518) );
  XOR U1864 ( .A(n2520), .B(n2521), .Z(n2506) );
  AND U1865 ( .A(n159), .B(n2519), .Z(n2521) );
  XNOR U1866 ( .A(n2520), .B(n2517), .Z(n2519) );
  XOR U1867 ( .A(n2522), .B(n2523), .Z(n2517) );
  AND U1868 ( .A(n162), .B(n2516), .Z(n2523) );
  XNOR U1869 ( .A(n2524), .B(n2514), .Z(n2516) );
  XOR U1870 ( .A(n2525), .B(n2526), .Z(n2514) );
  AND U1871 ( .A(n166), .B(n2527), .Z(n2526) );
  XOR U1872 ( .A(p_input[88]), .B(n2525), .Z(n2527) );
  XOR U1873 ( .A(n2528), .B(n2529), .Z(n2525) );
  AND U1874 ( .A(n170), .B(n2530), .Z(n2529) );
  IV U1875 ( .A(n2522), .Z(n2524) );
  XOR U1876 ( .A(n2531), .B(n2532), .Z(n2522) );
  AND U1877 ( .A(n174), .B(n2533), .Z(n2532) );
  XOR U1878 ( .A(n2534), .B(n2535), .Z(n2520) );
  AND U1879 ( .A(n178), .B(n2533), .Z(n2535) );
  XNOR U1880 ( .A(n2534), .B(n2531), .Z(n2533) );
  XOR U1881 ( .A(n2536), .B(n2537), .Z(n2531) );
  AND U1882 ( .A(n181), .B(n2530), .Z(n2537) );
  XNOR U1883 ( .A(n2538), .B(n2528), .Z(n2530) );
  XOR U1884 ( .A(n2539), .B(n2540), .Z(n2528) );
  AND U1885 ( .A(n185), .B(n2541), .Z(n2540) );
  XOR U1886 ( .A(p_input[104]), .B(n2539), .Z(n2541) );
  XOR U1887 ( .A(n2542), .B(n2543), .Z(n2539) );
  AND U1888 ( .A(n189), .B(n2544), .Z(n2543) );
  IV U1889 ( .A(n2536), .Z(n2538) );
  XOR U1890 ( .A(n2545), .B(n2546), .Z(n2536) );
  AND U1891 ( .A(n193), .B(n2547), .Z(n2546) );
  XOR U1892 ( .A(n2548), .B(n2549), .Z(n2534) );
  AND U1893 ( .A(n197), .B(n2547), .Z(n2549) );
  XNOR U1894 ( .A(n2548), .B(n2545), .Z(n2547) );
  XOR U1895 ( .A(n2550), .B(n2551), .Z(n2545) );
  AND U1896 ( .A(n200), .B(n2544), .Z(n2551) );
  XNOR U1897 ( .A(n2552), .B(n2542), .Z(n2544) );
  XOR U1898 ( .A(n2553), .B(n2554), .Z(n2542) );
  AND U1899 ( .A(n204), .B(n2555), .Z(n2554) );
  XOR U1900 ( .A(p_input[120]), .B(n2553), .Z(n2555) );
  XOR U1901 ( .A(n2556), .B(n2557), .Z(n2553) );
  AND U1902 ( .A(n208), .B(n2558), .Z(n2557) );
  IV U1903 ( .A(n2550), .Z(n2552) );
  XOR U1904 ( .A(n2559), .B(n2560), .Z(n2550) );
  AND U1905 ( .A(n212), .B(n2561), .Z(n2560) );
  XOR U1906 ( .A(n2562), .B(n2563), .Z(n2548) );
  AND U1907 ( .A(n216), .B(n2561), .Z(n2563) );
  XNOR U1908 ( .A(n2562), .B(n2559), .Z(n2561) );
  XOR U1909 ( .A(n2564), .B(n2565), .Z(n2559) );
  AND U1910 ( .A(n219), .B(n2558), .Z(n2565) );
  XNOR U1911 ( .A(n2566), .B(n2556), .Z(n2558) );
  XOR U1912 ( .A(n2567), .B(n2568), .Z(n2556) );
  AND U1913 ( .A(n223), .B(n2569), .Z(n2568) );
  XOR U1914 ( .A(p_input[136]), .B(n2567), .Z(n2569) );
  XOR U1915 ( .A(n2570), .B(n2571), .Z(n2567) );
  AND U1916 ( .A(n227), .B(n2572), .Z(n2571) );
  IV U1917 ( .A(n2564), .Z(n2566) );
  XOR U1918 ( .A(n2573), .B(n2574), .Z(n2564) );
  AND U1919 ( .A(n231), .B(n2575), .Z(n2574) );
  XOR U1920 ( .A(n2576), .B(n2577), .Z(n2562) );
  AND U1921 ( .A(n235), .B(n2575), .Z(n2577) );
  XNOR U1922 ( .A(n2576), .B(n2573), .Z(n2575) );
  XOR U1923 ( .A(n2578), .B(n2579), .Z(n2573) );
  AND U1924 ( .A(n238), .B(n2572), .Z(n2579) );
  XNOR U1925 ( .A(n2580), .B(n2570), .Z(n2572) );
  XOR U1926 ( .A(n2581), .B(n2582), .Z(n2570) );
  AND U1927 ( .A(n242), .B(n2583), .Z(n2582) );
  XOR U1928 ( .A(p_input[152]), .B(n2581), .Z(n2583) );
  XOR U1929 ( .A(n2584), .B(n2585), .Z(n2581) );
  AND U1930 ( .A(n246), .B(n2586), .Z(n2585) );
  IV U1931 ( .A(n2578), .Z(n2580) );
  XOR U1932 ( .A(n2587), .B(n2588), .Z(n2578) );
  AND U1933 ( .A(n250), .B(n2589), .Z(n2588) );
  XOR U1934 ( .A(n2590), .B(n2591), .Z(n2576) );
  AND U1935 ( .A(n254), .B(n2589), .Z(n2591) );
  XNOR U1936 ( .A(n2590), .B(n2587), .Z(n2589) );
  XOR U1937 ( .A(n2592), .B(n2593), .Z(n2587) );
  AND U1938 ( .A(n257), .B(n2586), .Z(n2593) );
  XNOR U1939 ( .A(n2594), .B(n2584), .Z(n2586) );
  XOR U1940 ( .A(n2595), .B(n2596), .Z(n2584) );
  AND U1941 ( .A(n261), .B(n2597), .Z(n2596) );
  XOR U1942 ( .A(p_input[168]), .B(n2595), .Z(n2597) );
  XOR U1943 ( .A(n2598), .B(n2599), .Z(n2595) );
  AND U1944 ( .A(n265), .B(n2600), .Z(n2599) );
  IV U1945 ( .A(n2592), .Z(n2594) );
  XOR U1946 ( .A(n2601), .B(n2602), .Z(n2592) );
  AND U1947 ( .A(n269), .B(n2603), .Z(n2602) );
  XOR U1948 ( .A(n2604), .B(n2605), .Z(n2590) );
  AND U1949 ( .A(n273), .B(n2603), .Z(n2605) );
  XNOR U1950 ( .A(n2604), .B(n2601), .Z(n2603) );
  XOR U1951 ( .A(n2606), .B(n2607), .Z(n2601) );
  AND U1952 ( .A(n276), .B(n2600), .Z(n2607) );
  XNOR U1953 ( .A(n2608), .B(n2598), .Z(n2600) );
  XOR U1954 ( .A(n2609), .B(n2610), .Z(n2598) );
  AND U1955 ( .A(n280), .B(n2611), .Z(n2610) );
  XOR U1956 ( .A(p_input[184]), .B(n2609), .Z(n2611) );
  XOR U1957 ( .A(n2612), .B(n2613), .Z(n2609) );
  AND U1958 ( .A(n284), .B(n2614), .Z(n2613) );
  IV U1959 ( .A(n2606), .Z(n2608) );
  XOR U1960 ( .A(n2615), .B(n2616), .Z(n2606) );
  AND U1961 ( .A(n288), .B(n2617), .Z(n2616) );
  XOR U1962 ( .A(n2618), .B(n2619), .Z(n2604) );
  AND U1963 ( .A(n292), .B(n2617), .Z(n2619) );
  XNOR U1964 ( .A(n2618), .B(n2615), .Z(n2617) );
  XOR U1965 ( .A(n2620), .B(n2621), .Z(n2615) );
  AND U1966 ( .A(n295), .B(n2614), .Z(n2621) );
  XNOR U1967 ( .A(n2622), .B(n2612), .Z(n2614) );
  XOR U1968 ( .A(n2623), .B(n2624), .Z(n2612) );
  AND U1969 ( .A(n299), .B(n2625), .Z(n2624) );
  XOR U1970 ( .A(p_input[200]), .B(n2623), .Z(n2625) );
  XOR U1971 ( .A(n2626), .B(n2627), .Z(n2623) );
  AND U1972 ( .A(n303), .B(n2628), .Z(n2627) );
  IV U1973 ( .A(n2620), .Z(n2622) );
  XOR U1974 ( .A(n2629), .B(n2630), .Z(n2620) );
  AND U1975 ( .A(n307), .B(n2631), .Z(n2630) );
  XOR U1976 ( .A(n2632), .B(n2633), .Z(n2618) );
  AND U1977 ( .A(n311), .B(n2631), .Z(n2633) );
  XNOR U1978 ( .A(n2632), .B(n2629), .Z(n2631) );
  XOR U1979 ( .A(n2634), .B(n2635), .Z(n2629) );
  AND U1980 ( .A(n314), .B(n2628), .Z(n2635) );
  XNOR U1981 ( .A(n2636), .B(n2626), .Z(n2628) );
  XOR U1982 ( .A(n2637), .B(n2638), .Z(n2626) );
  AND U1983 ( .A(n318), .B(n2639), .Z(n2638) );
  XOR U1984 ( .A(p_input[216]), .B(n2637), .Z(n2639) );
  XOR U1985 ( .A(n2640), .B(n2641), .Z(n2637) );
  AND U1986 ( .A(n322), .B(n2642), .Z(n2641) );
  IV U1987 ( .A(n2634), .Z(n2636) );
  XOR U1988 ( .A(n2643), .B(n2644), .Z(n2634) );
  AND U1989 ( .A(n326), .B(n2645), .Z(n2644) );
  XOR U1990 ( .A(n2646), .B(n2647), .Z(n2632) );
  AND U1991 ( .A(n330), .B(n2645), .Z(n2647) );
  XNOR U1992 ( .A(n2646), .B(n2643), .Z(n2645) );
  XOR U1993 ( .A(n2648), .B(n2649), .Z(n2643) );
  AND U1994 ( .A(n333), .B(n2642), .Z(n2649) );
  XNOR U1995 ( .A(n2650), .B(n2640), .Z(n2642) );
  XOR U1996 ( .A(n2651), .B(n2652), .Z(n2640) );
  AND U1997 ( .A(n337), .B(n2653), .Z(n2652) );
  XOR U1998 ( .A(p_input[232]), .B(n2651), .Z(n2653) );
  XOR U1999 ( .A(n2654), .B(n2655), .Z(n2651) );
  AND U2000 ( .A(n341), .B(n2656), .Z(n2655) );
  IV U2001 ( .A(n2648), .Z(n2650) );
  XOR U2002 ( .A(n2657), .B(n2658), .Z(n2648) );
  AND U2003 ( .A(n345), .B(n2659), .Z(n2658) );
  XOR U2004 ( .A(n2660), .B(n2661), .Z(n2646) );
  AND U2005 ( .A(n349), .B(n2659), .Z(n2661) );
  XNOR U2006 ( .A(n2660), .B(n2657), .Z(n2659) );
  XOR U2007 ( .A(n2662), .B(n2663), .Z(n2657) );
  AND U2008 ( .A(n352), .B(n2656), .Z(n2663) );
  XNOR U2009 ( .A(n2664), .B(n2654), .Z(n2656) );
  XOR U2010 ( .A(n2665), .B(n2666), .Z(n2654) );
  AND U2011 ( .A(n356), .B(n2667), .Z(n2666) );
  XOR U2012 ( .A(p_input[248]), .B(n2665), .Z(n2667) );
  XOR U2013 ( .A(n2668), .B(n2669), .Z(n2665) );
  AND U2014 ( .A(n360), .B(n2670), .Z(n2669) );
  IV U2015 ( .A(n2662), .Z(n2664) );
  XOR U2016 ( .A(n2671), .B(n2672), .Z(n2662) );
  AND U2017 ( .A(n364), .B(n2673), .Z(n2672) );
  XOR U2018 ( .A(n2674), .B(n2675), .Z(n2660) );
  AND U2019 ( .A(n368), .B(n2673), .Z(n2675) );
  XNOR U2020 ( .A(n2674), .B(n2671), .Z(n2673) );
  XOR U2021 ( .A(n2676), .B(n2677), .Z(n2671) );
  AND U2022 ( .A(n371), .B(n2670), .Z(n2677) );
  XNOR U2023 ( .A(n2678), .B(n2668), .Z(n2670) );
  XOR U2024 ( .A(n2679), .B(n2680), .Z(n2668) );
  AND U2025 ( .A(n375), .B(n2681), .Z(n2680) );
  XOR U2026 ( .A(p_input[264]), .B(n2679), .Z(n2681) );
  XOR U2027 ( .A(n2682), .B(n2683), .Z(n2679) );
  AND U2028 ( .A(n379), .B(n2684), .Z(n2683) );
  IV U2029 ( .A(n2676), .Z(n2678) );
  XOR U2030 ( .A(n2685), .B(n2686), .Z(n2676) );
  AND U2031 ( .A(n383), .B(n2687), .Z(n2686) );
  XOR U2032 ( .A(n2688), .B(n2689), .Z(n2674) );
  AND U2033 ( .A(n387), .B(n2687), .Z(n2689) );
  XNOR U2034 ( .A(n2688), .B(n2685), .Z(n2687) );
  XOR U2035 ( .A(n2690), .B(n2691), .Z(n2685) );
  AND U2036 ( .A(n390), .B(n2684), .Z(n2691) );
  XNOR U2037 ( .A(n2692), .B(n2682), .Z(n2684) );
  XOR U2038 ( .A(n2693), .B(n2694), .Z(n2682) );
  AND U2039 ( .A(n394), .B(n2695), .Z(n2694) );
  XOR U2040 ( .A(p_input[280]), .B(n2693), .Z(n2695) );
  XOR U2041 ( .A(n2696), .B(n2697), .Z(n2693) );
  AND U2042 ( .A(n398), .B(n2698), .Z(n2697) );
  IV U2043 ( .A(n2690), .Z(n2692) );
  XOR U2044 ( .A(n2699), .B(n2700), .Z(n2690) );
  AND U2045 ( .A(n402), .B(n2701), .Z(n2700) );
  XOR U2046 ( .A(n2702), .B(n2703), .Z(n2688) );
  AND U2047 ( .A(n406), .B(n2701), .Z(n2703) );
  XNOR U2048 ( .A(n2702), .B(n2699), .Z(n2701) );
  XOR U2049 ( .A(n2704), .B(n2705), .Z(n2699) );
  AND U2050 ( .A(n409), .B(n2698), .Z(n2705) );
  XNOR U2051 ( .A(n2706), .B(n2696), .Z(n2698) );
  XOR U2052 ( .A(n2707), .B(n2708), .Z(n2696) );
  AND U2053 ( .A(n413), .B(n2709), .Z(n2708) );
  XOR U2054 ( .A(p_input[296]), .B(n2707), .Z(n2709) );
  XOR U2055 ( .A(n2710), .B(n2711), .Z(n2707) );
  AND U2056 ( .A(n417), .B(n2712), .Z(n2711) );
  IV U2057 ( .A(n2704), .Z(n2706) );
  XOR U2058 ( .A(n2713), .B(n2714), .Z(n2704) );
  AND U2059 ( .A(n421), .B(n2715), .Z(n2714) );
  XOR U2060 ( .A(n2716), .B(n2717), .Z(n2702) );
  AND U2061 ( .A(n425), .B(n2715), .Z(n2717) );
  XNOR U2062 ( .A(n2716), .B(n2713), .Z(n2715) );
  XOR U2063 ( .A(n2718), .B(n2719), .Z(n2713) );
  AND U2064 ( .A(n428), .B(n2712), .Z(n2719) );
  XNOR U2065 ( .A(n2720), .B(n2710), .Z(n2712) );
  XOR U2066 ( .A(n2721), .B(n2722), .Z(n2710) );
  AND U2067 ( .A(n432), .B(n2723), .Z(n2722) );
  XOR U2068 ( .A(p_input[312]), .B(n2721), .Z(n2723) );
  XOR U2069 ( .A(n2724), .B(n2725), .Z(n2721) );
  AND U2070 ( .A(n436), .B(n2726), .Z(n2725) );
  IV U2071 ( .A(n2718), .Z(n2720) );
  XOR U2072 ( .A(n2727), .B(n2728), .Z(n2718) );
  AND U2073 ( .A(n440), .B(n2729), .Z(n2728) );
  XOR U2074 ( .A(n2730), .B(n2731), .Z(n2716) );
  AND U2075 ( .A(n444), .B(n2729), .Z(n2731) );
  XNOR U2076 ( .A(n2730), .B(n2727), .Z(n2729) );
  XOR U2077 ( .A(n2732), .B(n2733), .Z(n2727) );
  AND U2078 ( .A(n447), .B(n2726), .Z(n2733) );
  XNOR U2079 ( .A(n2734), .B(n2724), .Z(n2726) );
  XOR U2080 ( .A(n2735), .B(n2736), .Z(n2724) );
  AND U2081 ( .A(n451), .B(n2737), .Z(n2736) );
  XOR U2082 ( .A(p_input[328]), .B(n2735), .Z(n2737) );
  XOR U2083 ( .A(n2738), .B(n2739), .Z(n2735) );
  AND U2084 ( .A(n455), .B(n2740), .Z(n2739) );
  IV U2085 ( .A(n2732), .Z(n2734) );
  XOR U2086 ( .A(n2741), .B(n2742), .Z(n2732) );
  AND U2087 ( .A(n459), .B(n2743), .Z(n2742) );
  XOR U2088 ( .A(n2744), .B(n2745), .Z(n2730) );
  AND U2089 ( .A(n463), .B(n2743), .Z(n2745) );
  XNOR U2090 ( .A(n2744), .B(n2741), .Z(n2743) );
  XOR U2091 ( .A(n2746), .B(n2747), .Z(n2741) );
  AND U2092 ( .A(n466), .B(n2740), .Z(n2747) );
  XNOR U2093 ( .A(n2748), .B(n2738), .Z(n2740) );
  XOR U2094 ( .A(n2749), .B(n2750), .Z(n2738) );
  AND U2095 ( .A(n470), .B(n2751), .Z(n2750) );
  XOR U2096 ( .A(p_input[344]), .B(n2749), .Z(n2751) );
  XOR U2097 ( .A(n2752), .B(n2753), .Z(n2749) );
  AND U2098 ( .A(n474), .B(n2754), .Z(n2753) );
  IV U2099 ( .A(n2746), .Z(n2748) );
  XOR U2100 ( .A(n2755), .B(n2756), .Z(n2746) );
  AND U2101 ( .A(n478), .B(n2757), .Z(n2756) );
  XOR U2102 ( .A(n2758), .B(n2759), .Z(n2744) );
  AND U2103 ( .A(n482), .B(n2757), .Z(n2759) );
  XNOR U2104 ( .A(n2758), .B(n2755), .Z(n2757) );
  XOR U2105 ( .A(n2760), .B(n2761), .Z(n2755) );
  AND U2106 ( .A(n485), .B(n2754), .Z(n2761) );
  XNOR U2107 ( .A(n2762), .B(n2752), .Z(n2754) );
  XOR U2108 ( .A(n2763), .B(n2764), .Z(n2752) );
  AND U2109 ( .A(n489), .B(n2765), .Z(n2764) );
  XOR U2110 ( .A(p_input[360]), .B(n2763), .Z(n2765) );
  XOR U2111 ( .A(n2766), .B(n2767), .Z(n2763) );
  AND U2112 ( .A(n493), .B(n2768), .Z(n2767) );
  IV U2113 ( .A(n2760), .Z(n2762) );
  XOR U2114 ( .A(n2769), .B(n2770), .Z(n2760) );
  AND U2115 ( .A(n497), .B(n2771), .Z(n2770) );
  XOR U2116 ( .A(n2772), .B(n2773), .Z(n2758) );
  AND U2117 ( .A(n501), .B(n2771), .Z(n2773) );
  XNOR U2118 ( .A(n2772), .B(n2769), .Z(n2771) );
  XOR U2119 ( .A(n2774), .B(n2775), .Z(n2769) );
  AND U2120 ( .A(n504), .B(n2768), .Z(n2775) );
  XNOR U2121 ( .A(n2776), .B(n2766), .Z(n2768) );
  XOR U2122 ( .A(n2777), .B(n2778), .Z(n2766) );
  AND U2123 ( .A(n508), .B(n2779), .Z(n2778) );
  XOR U2124 ( .A(p_input[376]), .B(n2777), .Z(n2779) );
  XOR U2125 ( .A(n2780), .B(n2781), .Z(n2777) );
  AND U2126 ( .A(n512), .B(n2782), .Z(n2781) );
  IV U2127 ( .A(n2774), .Z(n2776) );
  XOR U2128 ( .A(n2783), .B(n2784), .Z(n2774) );
  AND U2129 ( .A(n516), .B(n2785), .Z(n2784) );
  XOR U2130 ( .A(n2786), .B(n2787), .Z(n2772) );
  AND U2131 ( .A(n520), .B(n2785), .Z(n2787) );
  XNOR U2132 ( .A(n2786), .B(n2783), .Z(n2785) );
  XOR U2133 ( .A(n2788), .B(n2789), .Z(n2783) );
  AND U2134 ( .A(n523), .B(n2782), .Z(n2789) );
  XNOR U2135 ( .A(n2790), .B(n2780), .Z(n2782) );
  XOR U2136 ( .A(n2791), .B(n2792), .Z(n2780) );
  AND U2137 ( .A(n527), .B(n2793), .Z(n2792) );
  XOR U2138 ( .A(p_input[392]), .B(n2791), .Z(n2793) );
  XOR U2139 ( .A(n2794), .B(n2795), .Z(n2791) );
  AND U2140 ( .A(n531), .B(n2796), .Z(n2795) );
  IV U2141 ( .A(n2788), .Z(n2790) );
  XOR U2142 ( .A(n2797), .B(n2798), .Z(n2788) );
  AND U2143 ( .A(n535), .B(n2799), .Z(n2798) );
  XOR U2144 ( .A(n2800), .B(n2801), .Z(n2786) );
  AND U2145 ( .A(n539), .B(n2799), .Z(n2801) );
  XNOR U2146 ( .A(n2800), .B(n2797), .Z(n2799) );
  XOR U2147 ( .A(n2802), .B(n2803), .Z(n2797) );
  AND U2148 ( .A(n542), .B(n2796), .Z(n2803) );
  XNOR U2149 ( .A(n2804), .B(n2794), .Z(n2796) );
  XOR U2150 ( .A(n2805), .B(n2806), .Z(n2794) );
  AND U2151 ( .A(n546), .B(n2807), .Z(n2806) );
  XOR U2152 ( .A(p_input[408]), .B(n2805), .Z(n2807) );
  XOR U2153 ( .A(n2808), .B(n2809), .Z(n2805) );
  AND U2154 ( .A(n550), .B(n2810), .Z(n2809) );
  IV U2155 ( .A(n2802), .Z(n2804) );
  XOR U2156 ( .A(n2811), .B(n2812), .Z(n2802) );
  AND U2157 ( .A(n554), .B(n2813), .Z(n2812) );
  XOR U2158 ( .A(n2814), .B(n2815), .Z(n2800) );
  AND U2159 ( .A(n558), .B(n2813), .Z(n2815) );
  XNOR U2160 ( .A(n2814), .B(n2811), .Z(n2813) );
  XOR U2161 ( .A(n2816), .B(n2817), .Z(n2811) );
  AND U2162 ( .A(n561), .B(n2810), .Z(n2817) );
  XNOR U2163 ( .A(n2818), .B(n2808), .Z(n2810) );
  XOR U2164 ( .A(n2819), .B(n2820), .Z(n2808) );
  AND U2165 ( .A(n565), .B(n2821), .Z(n2820) );
  XOR U2166 ( .A(p_input[424]), .B(n2819), .Z(n2821) );
  XOR U2167 ( .A(n2822), .B(n2823), .Z(n2819) );
  AND U2168 ( .A(n569), .B(n2824), .Z(n2823) );
  IV U2169 ( .A(n2816), .Z(n2818) );
  XOR U2170 ( .A(n2825), .B(n2826), .Z(n2816) );
  AND U2171 ( .A(n573), .B(n2827), .Z(n2826) );
  XOR U2172 ( .A(n2828), .B(n2829), .Z(n2814) );
  AND U2173 ( .A(n577), .B(n2827), .Z(n2829) );
  XNOR U2174 ( .A(n2828), .B(n2825), .Z(n2827) );
  XOR U2175 ( .A(n2830), .B(n2831), .Z(n2825) );
  AND U2176 ( .A(n580), .B(n2824), .Z(n2831) );
  XNOR U2177 ( .A(n2832), .B(n2822), .Z(n2824) );
  XOR U2178 ( .A(n2833), .B(n2834), .Z(n2822) );
  AND U2179 ( .A(n584), .B(n2835), .Z(n2834) );
  XOR U2180 ( .A(p_input[440]), .B(n2833), .Z(n2835) );
  XOR U2181 ( .A(n2836), .B(n2837), .Z(n2833) );
  AND U2182 ( .A(n588), .B(n2838), .Z(n2837) );
  IV U2183 ( .A(n2830), .Z(n2832) );
  XOR U2184 ( .A(n2839), .B(n2840), .Z(n2830) );
  AND U2185 ( .A(n592), .B(n2841), .Z(n2840) );
  XOR U2186 ( .A(n2842), .B(n2843), .Z(n2828) );
  AND U2187 ( .A(n596), .B(n2841), .Z(n2843) );
  XNOR U2188 ( .A(n2842), .B(n2839), .Z(n2841) );
  XOR U2189 ( .A(n2844), .B(n2845), .Z(n2839) );
  AND U2190 ( .A(n599), .B(n2838), .Z(n2845) );
  XNOR U2191 ( .A(n2846), .B(n2836), .Z(n2838) );
  XOR U2192 ( .A(n2847), .B(n2848), .Z(n2836) );
  AND U2193 ( .A(n603), .B(n2849), .Z(n2848) );
  XOR U2194 ( .A(p_input[456]), .B(n2847), .Z(n2849) );
  XOR U2195 ( .A(n2850), .B(n2851), .Z(n2847) );
  AND U2196 ( .A(n607), .B(n2852), .Z(n2851) );
  IV U2197 ( .A(n2844), .Z(n2846) );
  XOR U2198 ( .A(n2853), .B(n2854), .Z(n2844) );
  AND U2199 ( .A(n611), .B(n2855), .Z(n2854) );
  XOR U2200 ( .A(n2856), .B(n2857), .Z(n2842) );
  AND U2201 ( .A(n615), .B(n2855), .Z(n2857) );
  XNOR U2202 ( .A(n2856), .B(n2853), .Z(n2855) );
  XOR U2203 ( .A(n2858), .B(n2859), .Z(n2853) );
  AND U2204 ( .A(n618), .B(n2852), .Z(n2859) );
  XNOR U2205 ( .A(n2860), .B(n2850), .Z(n2852) );
  XOR U2206 ( .A(n2861), .B(n2862), .Z(n2850) );
  AND U2207 ( .A(n622), .B(n2863), .Z(n2862) );
  XOR U2208 ( .A(p_input[472]), .B(n2861), .Z(n2863) );
  XOR U2209 ( .A(n2864), .B(n2865), .Z(n2861) );
  AND U2210 ( .A(n626), .B(n2866), .Z(n2865) );
  IV U2211 ( .A(n2858), .Z(n2860) );
  XOR U2212 ( .A(n2867), .B(n2868), .Z(n2858) );
  AND U2213 ( .A(n630), .B(n2869), .Z(n2868) );
  XOR U2214 ( .A(n2870), .B(n2871), .Z(n2856) );
  AND U2215 ( .A(n634), .B(n2869), .Z(n2871) );
  XNOR U2216 ( .A(n2870), .B(n2867), .Z(n2869) );
  XOR U2217 ( .A(n2872), .B(n2873), .Z(n2867) );
  AND U2218 ( .A(n637), .B(n2866), .Z(n2873) );
  XNOR U2219 ( .A(n2874), .B(n2864), .Z(n2866) );
  XOR U2220 ( .A(n2875), .B(n2876), .Z(n2864) );
  AND U2221 ( .A(n641), .B(n2877), .Z(n2876) );
  XOR U2222 ( .A(p_input[488]), .B(n2875), .Z(n2877) );
  XOR U2223 ( .A(n2878), .B(n2879), .Z(n2875) );
  AND U2224 ( .A(n645), .B(n2880), .Z(n2879) );
  IV U2225 ( .A(n2872), .Z(n2874) );
  XOR U2226 ( .A(n2881), .B(n2882), .Z(n2872) );
  AND U2227 ( .A(n649), .B(n2883), .Z(n2882) );
  XOR U2228 ( .A(n2884), .B(n2885), .Z(n2870) );
  AND U2229 ( .A(n653), .B(n2883), .Z(n2885) );
  XNOR U2230 ( .A(n2884), .B(n2881), .Z(n2883) );
  XOR U2231 ( .A(n2886), .B(n2887), .Z(n2881) );
  AND U2232 ( .A(n656), .B(n2880), .Z(n2887) );
  XNOR U2233 ( .A(n2888), .B(n2878), .Z(n2880) );
  XOR U2234 ( .A(n2889), .B(n2890), .Z(n2878) );
  AND U2235 ( .A(n660), .B(n2891), .Z(n2890) );
  XOR U2236 ( .A(p_input[504]), .B(n2889), .Z(n2891) );
  XOR U2237 ( .A(n2892), .B(n2893), .Z(n2889) );
  AND U2238 ( .A(n664), .B(n2894), .Z(n2893) );
  IV U2239 ( .A(n2886), .Z(n2888) );
  XOR U2240 ( .A(n2895), .B(n2896), .Z(n2886) );
  AND U2241 ( .A(n668), .B(n2897), .Z(n2896) );
  XOR U2242 ( .A(n2898), .B(n2899), .Z(n2884) );
  AND U2243 ( .A(n672), .B(n2897), .Z(n2899) );
  XNOR U2244 ( .A(n2898), .B(n2895), .Z(n2897) );
  XOR U2245 ( .A(n2900), .B(n2901), .Z(n2895) );
  AND U2246 ( .A(n675), .B(n2894), .Z(n2901) );
  XNOR U2247 ( .A(n2902), .B(n2892), .Z(n2894) );
  XOR U2248 ( .A(n2903), .B(n2904), .Z(n2892) );
  AND U2249 ( .A(n679), .B(n2905), .Z(n2904) );
  XOR U2250 ( .A(p_input[520]), .B(n2903), .Z(n2905) );
  XOR U2251 ( .A(n2906), .B(n2907), .Z(n2903) );
  AND U2252 ( .A(n683), .B(n2908), .Z(n2907) );
  IV U2253 ( .A(n2900), .Z(n2902) );
  XOR U2254 ( .A(n2909), .B(n2910), .Z(n2900) );
  AND U2255 ( .A(n687), .B(n2911), .Z(n2910) );
  XOR U2256 ( .A(n2912), .B(n2913), .Z(n2898) );
  AND U2257 ( .A(n691), .B(n2911), .Z(n2913) );
  XNOR U2258 ( .A(n2912), .B(n2909), .Z(n2911) );
  XOR U2259 ( .A(n2914), .B(n2915), .Z(n2909) );
  AND U2260 ( .A(n694), .B(n2908), .Z(n2915) );
  XNOR U2261 ( .A(n2916), .B(n2906), .Z(n2908) );
  XOR U2262 ( .A(n2917), .B(n2918), .Z(n2906) );
  AND U2263 ( .A(n698), .B(n2919), .Z(n2918) );
  XOR U2264 ( .A(p_input[536]), .B(n2917), .Z(n2919) );
  XOR U2265 ( .A(n2920), .B(n2921), .Z(n2917) );
  AND U2266 ( .A(n702), .B(n2922), .Z(n2921) );
  IV U2267 ( .A(n2914), .Z(n2916) );
  XOR U2268 ( .A(n2923), .B(n2924), .Z(n2914) );
  AND U2269 ( .A(n706), .B(n2925), .Z(n2924) );
  XOR U2270 ( .A(n2926), .B(n2927), .Z(n2912) );
  AND U2271 ( .A(n710), .B(n2925), .Z(n2927) );
  XNOR U2272 ( .A(n2926), .B(n2923), .Z(n2925) );
  XOR U2273 ( .A(n2928), .B(n2929), .Z(n2923) );
  AND U2274 ( .A(n713), .B(n2922), .Z(n2929) );
  XNOR U2275 ( .A(n2930), .B(n2920), .Z(n2922) );
  XOR U2276 ( .A(n2931), .B(n2932), .Z(n2920) );
  AND U2277 ( .A(n717), .B(n2933), .Z(n2932) );
  XOR U2278 ( .A(p_input[552]), .B(n2931), .Z(n2933) );
  XOR U2279 ( .A(n2934), .B(n2935), .Z(n2931) );
  AND U2280 ( .A(n721), .B(n2936), .Z(n2935) );
  IV U2281 ( .A(n2928), .Z(n2930) );
  XOR U2282 ( .A(n2937), .B(n2938), .Z(n2928) );
  AND U2283 ( .A(n725), .B(n2939), .Z(n2938) );
  XOR U2284 ( .A(n2940), .B(n2941), .Z(n2926) );
  AND U2285 ( .A(n729), .B(n2939), .Z(n2941) );
  XNOR U2286 ( .A(n2940), .B(n2937), .Z(n2939) );
  XOR U2287 ( .A(n2942), .B(n2943), .Z(n2937) );
  AND U2288 ( .A(n732), .B(n2936), .Z(n2943) );
  XNOR U2289 ( .A(n2944), .B(n2934), .Z(n2936) );
  XOR U2290 ( .A(n2945), .B(n2946), .Z(n2934) );
  AND U2291 ( .A(n736), .B(n2947), .Z(n2946) );
  XOR U2292 ( .A(p_input[568]), .B(n2945), .Z(n2947) );
  XOR U2293 ( .A(n2948), .B(n2949), .Z(n2945) );
  AND U2294 ( .A(n740), .B(n2950), .Z(n2949) );
  IV U2295 ( .A(n2942), .Z(n2944) );
  XOR U2296 ( .A(n2951), .B(n2952), .Z(n2942) );
  AND U2297 ( .A(n744), .B(n2953), .Z(n2952) );
  XOR U2298 ( .A(n2954), .B(n2955), .Z(n2940) );
  AND U2299 ( .A(n748), .B(n2953), .Z(n2955) );
  XNOR U2300 ( .A(n2954), .B(n2951), .Z(n2953) );
  XOR U2301 ( .A(n2956), .B(n2957), .Z(n2951) );
  AND U2302 ( .A(n751), .B(n2950), .Z(n2957) );
  XNOR U2303 ( .A(n2958), .B(n2948), .Z(n2950) );
  XOR U2304 ( .A(n2959), .B(n2960), .Z(n2948) );
  AND U2305 ( .A(n755), .B(n2961), .Z(n2960) );
  XOR U2306 ( .A(p_input[584]), .B(n2959), .Z(n2961) );
  XOR U2307 ( .A(n2962), .B(n2963), .Z(n2959) );
  AND U2308 ( .A(n759), .B(n2964), .Z(n2963) );
  IV U2309 ( .A(n2956), .Z(n2958) );
  XOR U2310 ( .A(n2965), .B(n2966), .Z(n2956) );
  AND U2311 ( .A(n763), .B(n2967), .Z(n2966) );
  XOR U2312 ( .A(n2968), .B(n2969), .Z(n2954) );
  AND U2313 ( .A(n767), .B(n2967), .Z(n2969) );
  XNOR U2314 ( .A(n2968), .B(n2965), .Z(n2967) );
  XOR U2315 ( .A(n2970), .B(n2971), .Z(n2965) );
  AND U2316 ( .A(n770), .B(n2964), .Z(n2971) );
  XNOR U2317 ( .A(n2972), .B(n2962), .Z(n2964) );
  XOR U2318 ( .A(n2973), .B(n2974), .Z(n2962) );
  AND U2319 ( .A(n774), .B(n2975), .Z(n2974) );
  XOR U2320 ( .A(p_input[600]), .B(n2973), .Z(n2975) );
  XOR U2321 ( .A(n2976), .B(n2977), .Z(n2973) );
  AND U2322 ( .A(n778), .B(n2978), .Z(n2977) );
  IV U2323 ( .A(n2970), .Z(n2972) );
  XOR U2324 ( .A(n2979), .B(n2980), .Z(n2970) );
  AND U2325 ( .A(n782), .B(n2981), .Z(n2980) );
  XOR U2326 ( .A(n2982), .B(n2983), .Z(n2968) );
  AND U2327 ( .A(n786), .B(n2981), .Z(n2983) );
  XNOR U2328 ( .A(n2982), .B(n2979), .Z(n2981) );
  XOR U2329 ( .A(n2984), .B(n2985), .Z(n2979) );
  AND U2330 ( .A(n789), .B(n2978), .Z(n2985) );
  XNOR U2331 ( .A(n2986), .B(n2976), .Z(n2978) );
  XOR U2332 ( .A(n2987), .B(n2988), .Z(n2976) );
  AND U2333 ( .A(n793), .B(n2989), .Z(n2988) );
  XOR U2334 ( .A(p_input[616]), .B(n2987), .Z(n2989) );
  XOR U2335 ( .A(n2990), .B(n2991), .Z(n2987) );
  AND U2336 ( .A(n797), .B(n2992), .Z(n2991) );
  IV U2337 ( .A(n2984), .Z(n2986) );
  XOR U2338 ( .A(n2993), .B(n2994), .Z(n2984) );
  AND U2339 ( .A(n801), .B(n2995), .Z(n2994) );
  XOR U2340 ( .A(n2996), .B(n2997), .Z(n2982) );
  AND U2341 ( .A(n805), .B(n2995), .Z(n2997) );
  XNOR U2342 ( .A(n2996), .B(n2993), .Z(n2995) );
  XOR U2343 ( .A(n2998), .B(n2999), .Z(n2993) );
  AND U2344 ( .A(n808), .B(n2992), .Z(n2999) );
  XNOR U2345 ( .A(n3000), .B(n2990), .Z(n2992) );
  XOR U2346 ( .A(n3001), .B(n3002), .Z(n2990) );
  AND U2347 ( .A(n812), .B(n3003), .Z(n3002) );
  XOR U2348 ( .A(p_input[632]), .B(n3001), .Z(n3003) );
  XOR U2349 ( .A(n3004), .B(n3005), .Z(n3001) );
  AND U2350 ( .A(n816), .B(n3006), .Z(n3005) );
  IV U2351 ( .A(n2998), .Z(n3000) );
  XOR U2352 ( .A(n3007), .B(n3008), .Z(n2998) );
  AND U2353 ( .A(n820), .B(n3009), .Z(n3008) );
  XOR U2354 ( .A(n3010), .B(n3011), .Z(n2996) );
  AND U2355 ( .A(n824), .B(n3009), .Z(n3011) );
  XNOR U2356 ( .A(n3010), .B(n3007), .Z(n3009) );
  XOR U2357 ( .A(n3012), .B(n3013), .Z(n3007) );
  AND U2358 ( .A(n827), .B(n3006), .Z(n3013) );
  XNOR U2359 ( .A(n3014), .B(n3004), .Z(n3006) );
  XOR U2360 ( .A(n3015), .B(n3016), .Z(n3004) );
  AND U2361 ( .A(n831), .B(n3017), .Z(n3016) );
  XOR U2362 ( .A(p_input[648]), .B(n3015), .Z(n3017) );
  XOR U2363 ( .A(n3018), .B(n3019), .Z(n3015) );
  AND U2364 ( .A(n835), .B(n3020), .Z(n3019) );
  IV U2365 ( .A(n3012), .Z(n3014) );
  XOR U2366 ( .A(n3021), .B(n3022), .Z(n3012) );
  AND U2367 ( .A(n839), .B(n3023), .Z(n3022) );
  XOR U2368 ( .A(n3024), .B(n3025), .Z(n3010) );
  AND U2369 ( .A(n843), .B(n3023), .Z(n3025) );
  XNOR U2370 ( .A(n3024), .B(n3021), .Z(n3023) );
  XOR U2371 ( .A(n3026), .B(n3027), .Z(n3021) );
  AND U2372 ( .A(n846), .B(n3020), .Z(n3027) );
  XNOR U2373 ( .A(n3028), .B(n3018), .Z(n3020) );
  XOR U2374 ( .A(n3029), .B(n3030), .Z(n3018) );
  AND U2375 ( .A(n850), .B(n3031), .Z(n3030) );
  XOR U2376 ( .A(p_input[664]), .B(n3029), .Z(n3031) );
  XOR U2377 ( .A(n3032), .B(n3033), .Z(n3029) );
  AND U2378 ( .A(n854), .B(n3034), .Z(n3033) );
  IV U2379 ( .A(n3026), .Z(n3028) );
  XOR U2380 ( .A(n3035), .B(n3036), .Z(n3026) );
  AND U2381 ( .A(n858), .B(n3037), .Z(n3036) );
  XOR U2382 ( .A(n3038), .B(n3039), .Z(n3024) );
  AND U2383 ( .A(n862), .B(n3037), .Z(n3039) );
  XNOR U2384 ( .A(n3038), .B(n3035), .Z(n3037) );
  XOR U2385 ( .A(n3040), .B(n3041), .Z(n3035) );
  AND U2386 ( .A(n865), .B(n3034), .Z(n3041) );
  XNOR U2387 ( .A(n3042), .B(n3032), .Z(n3034) );
  XOR U2388 ( .A(n3043), .B(n3044), .Z(n3032) );
  AND U2389 ( .A(n869), .B(n3045), .Z(n3044) );
  XOR U2390 ( .A(p_input[680]), .B(n3043), .Z(n3045) );
  XOR U2391 ( .A(n3046), .B(n3047), .Z(n3043) );
  AND U2392 ( .A(n873), .B(n3048), .Z(n3047) );
  IV U2393 ( .A(n3040), .Z(n3042) );
  XOR U2394 ( .A(n3049), .B(n3050), .Z(n3040) );
  AND U2395 ( .A(n877), .B(n3051), .Z(n3050) );
  XOR U2396 ( .A(n3052), .B(n3053), .Z(n3038) );
  AND U2397 ( .A(n881), .B(n3051), .Z(n3053) );
  XNOR U2398 ( .A(n3052), .B(n3049), .Z(n3051) );
  XOR U2399 ( .A(n3054), .B(n3055), .Z(n3049) );
  AND U2400 ( .A(n884), .B(n3048), .Z(n3055) );
  XNOR U2401 ( .A(n3056), .B(n3046), .Z(n3048) );
  XOR U2402 ( .A(n3057), .B(n3058), .Z(n3046) );
  AND U2403 ( .A(n888), .B(n3059), .Z(n3058) );
  XOR U2404 ( .A(p_input[696]), .B(n3057), .Z(n3059) );
  XOR U2405 ( .A(n3060), .B(n3061), .Z(n3057) );
  AND U2406 ( .A(n892), .B(n3062), .Z(n3061) );
  IV U2407 ( .A(n3054), .Z(n3056) );
  XOR U2408 ( .A(n3063), .B(n3064), .Z(n3054) );
  AND U2409 ( .A(n896), .B(n3065), .Z(n3064) );
  XOR U2410 ( .A(n3066), .B(n3067), .Z(n3052) );
  AND U2411 ( .A(n900), .B(n3065), .Z(n3067) );
  XNOR U2412 ( .A(n3066), .B(n3063), .Z(n3065) );
  XOR U2413 ( .A(n3068), .B(n3069), .Z(n3063) );
  AND U2414 ( .A(n903), .B(n3062), .Z(n3069) );
  XNOR U2415 ( .A(n3070), .B(n3060), .Z(n3062) );
  XOR U2416 ( .A(n3071), .B(n3072), .Z(n3060) );
  AND U2417 ( .A(n907), .B(n3073), .Z(n3072) );
  XOR U2418 ( .A(p_input[712]), .B(n3071), .Z(n3073) );
  XOR U2419 ( .A(n3074), .B(n3075), .Z(n3071) );
  AND U2420 ( .A(n911), .B(n3076), .Z(n3075) );
  IV U2421 ( .A(n3068), .Z(n3070) );
  XOR U2422 ( .A(n3077), .B(n3078), .Z(n3068) );
  AND U2423 ( .A(n915), .B(n3079), .Z(n3078) );
  XOR U2424 ( .A(n3080), .B(n3081), .Z(n3066) );
  AND U2425 ( .A(n919), .B(n3079), .Z(n3081) );
  XNOR U2426 ( .A(n3080), .B(n3077), .Z(n3079) );
  XOR U2427 ( .A(n3082), .B(n3083), .Z(n3077) );
  AND U2428 ( .A(n922), .B(n3076), .Z(n3083) );
  XNOR U2429 ( .A(n3084), .B(n3074), .Z(n3076) );
  XOR U2430 ( .A(n3085), .B(n3086), .Z(n3074) );
  AND U2431 ( .A(n926), .B(n3087), .Z(n3086) );
  XOR U2432 ( .A(p_input[728]), .B(n3085), .Z(n3087) );
  XOR U2433 ( .A(n3088), .B(n3089), .Z(n3085) );
  AND U2434 ( .A(n930), .B(n3090), .Z(n3089) );
  IV U2435 ( .A(n3082), .Z(n3084) );
  XOR U2436 ( .A(n3091), .B(n3092), .Z(n3082) );
  AND U2437 ( .A(n934), .B(n3093), .Z(n3092) );
  XOR U2438 ( .A(n3094), .B(n3095), .Z(n3080) );
  AND U2439 ( .A(n938), .B(n3093), .Z(n3095) );
  XNOR U2440 ( .A(n3094), .B(n3091), .Z(n3093) );
  XOR U2441 ( .A(n3096), .B(n3097), .Z(n3091) );
  AND U2442 ( .A(n941), .B(n3090), .Z(n3097) );
  XNOR U2443 ( .A(n3098), .B(n3088), .Z(n3090) );
  XOR U2444 ( .A(n3099), .B(n3100), .Z(n3088) );
  AND U2445 ( .A(n945), .B(n3101), .Z(n3100) );
  XOR U2446 ( .A(p_input[744]), .B(n3099), .Z(n3101) );
  XOR U2447 ( .A(n3102), .B(n3103), .Z(n3099) );
  AND U2448 ( .A(n949), .B(n3104), .Z(n3103) );
  IV U2449 ( .A(n3096), .Z(n3098) );
  XOR U2450 ( .A(n3105), .B(n3106), .Z(n3096) );
  AND U2451 ( .A(n953), .B(n3107), .Z(n3106) );
  XOR U2452 ( .A(n3108), .B(n3109), .Z(n3094) );
  AND U2453 ( .A(n957), .B(n3107), .Z(n3109) );
  XNOR U2454 ( .A(n3108), .B(n3105), .Z(n3107) );
  XOR U2455 ( .A(n3110), .B(n3111), .Z(n3105) );
  AND U2456 ( .A(n960), .B(n3104), .Z(n3111) );
  XNOR U2457 ( .A(n3112), .B(n3102), .Z(n3104) );
  XOR U2458 ( .A(n3113), .B(n3114), .Z(n3102) );
  AND U2459 ( .A(n964), .B(n3115), .Z(n3114) );
  XOR U2460 ( .A(p_input[760]), .B(n3113), .Z(n3115) );
  XOR U2461 ( .A(n3116), .B(n3117), .Z(n3113) );
  AND U2462 ( .A(n968), .B(n3118), .Z(n3117) );
  IV U2463 ( .A(n3110), .Z(n3112) );
  XOR U2464 ( .A(n3119), .B(n3120), .Z(n3110) );
  AND U2465 ( .A(n972), .B(n3121), .Z(n3120) );
  XOR U2466 ( .A(n3122), .B(n3123), .Z(n3108) );
  AND U2467 ( .A(n976), .B(n3121), .Z(n3123) );
  XNOR U2468 ( .A(n3122), .B(n3119), .Z(n3121) );
  XOR U2469 ( .A(n3124), .B(n3125), .Z(n3119) );
  AND U2470 ( .A(n979), .B(n3118), .Z(n3125) );
  XNOR U2471 ( .A(n3126), .B(n3116), .Z(n3118) );
  XOR U2472 ( .A(n3127), .B(n3128), .Z(n3116) );
  AND U2473 ( .A(n983), .B(n3129), .Z(n3128) );
  XOR U2474 ( .A(p_input[776]), .B(n3127), .Z(n3129) );
  XOR U2475 ( .A(n3130), .B(n3131), .Z(n3127) );
  AND U2476 ( .A(n987), .B(n3132), .Z(n3131) );
  IV U2477 ( .A(n3124), .Z(n3126) );
  XOR U2478 ( .A(n3133), .B(n3134), .Z(n3124) );
  AND U2479 ( .A(n991), .B(n3135), .Z(n3134) );
  XOR U2480 ( .A(n3136), .B(n3137), .Z(n3122) );
  AND U2481 ( .A(n995), .B(n3135), .Z(n3137) );
  XNOR U2482 ( .A(n3136), .B(n3133), .Z(n3135) );
  XOR U2483 ( .A(n3138), .B(n3139), .Z(n3133) );
  AND U2484 ( .A(n998), .B(n3132), .Z(n3139) );
  XNOR U2485 ( .A(n3140), .B(n3130), .Z(n3132) );
  XOR U2486 ( .A(n3141), .B(n3142), .Z(n3130) );
  AND U2487 ( .A(n1002), .B(n3143), .Z(n3142) );
  XOR U2488 ( .A(p_input[792]), .B(n3141), .Z(n3143) );
  XOR U2489 ( .A(n3144), .B(n3145), .Z(n3141) );
  AND U2490 ( .A(n1006), .B(n3146), .Z(n3145) );
  IV U2491 ( .A(n3138), .Z(n3140) );
  XOR U2492 ( .A(n3147), .B(n3148), .Z(n3138) );
  AND U2493 ( .A(n1010), .B(n3149), .Z(n3148) );
  XOR U2494 ( .A(n3150), .B(n3151), .Z(n3136) );
  AND U2495 ( .A(n1014), .B(n3149), .Z(n3151) );
  XNOR U2496 ( .A(n3150), .B(n3147), .Z(n3149) );
  XOR U2497 ( .A(n3152), .B(n3153), .Z(n3147) );
  AND U2498 ( .A(n1017), .B(n3146), .Z(n3153) );
  XNOR U2499 ( .A(n3154), .B(n3144), .Z(n3146) );
  XOR U2500 ( .A(n3155), .B(n3156), .Z(n3144) );
  AND U2501 ( .A(n1021), .B(n3157), .Z(n3156) );
  XOR U2502 ( .A(p_input[808]), .B(n3155), .Z(n3157) );
  XOR U2503 ( .A(n3158), .B(n3159), .Z(n3155) );
  AND U2504 ( .A(n1025), .B(n3160), .Z(n3159) );
  IV U2505 ( .A(n3152), .Z(n3154) );
  XOR U2506 ( .A(n3161), .B(n3162), .Z(n3152) );
  AND U2507 ( .A(n1029), .B(n3163), .Z(n3162) );
  XOR U2508 ( .A(n3164), .B(n3165), .Z(n3150) );
  AND U2509 ( .A(n1033), .B(n3163), .Z(n3165) );
  XNOR U2510 ( .A(n3164), .B(n3161), .Z(n3163) );
  XOR U2511 ( .A(n3166), .B(n3167), .Z(n3161) );
  AND U2512 ( .A(n1036), .B(n3160), .Z(n3167) );
  XNOR U2513 ( .A(n3168), .B(n3158), .Z(n3160) );
  XOR U2514 ( .A(n3169), .B(n3170), .Z(n3158) );
  AND U2515 ( .A(n1040), .B(n3171), .Z(n3170) );
  XOR U2516 ( .A(p_input[824]), .B(n3169), .Z(n3171) );
  XOR U2517 ( .A(n3172), .B(n3173), .Z(n3169) );
  AND U2518 ( .A(n1044), .B(n3174), .Z(n3173) );
  IV U2519 ( .A(n3166), .Z(n3168) );
  XOR U2520 ( .A(n3175), .B(n3176), .Z(n3166) );
  AND U2521 ( .A(n1048), .B(n3177), .Z(n3176) );
  XOR U2522 ( .A(n3178), .B(n3179), .Z(n3164) );
  AND U2523 ( .A(n1052), .B(n3177), .Z(n3179) );
  XNOR U2524 ( .A(n3178), .B(n3175), .Z(n3177) );
  XOR U2525 ( .A(n3180), .B(n3181), .Z(n3175) );
  AND U2526 ( .A(n1055), .B(n3174), .Z(n3181) );
  XNOR U2527 ( .A(n3182), .B(n3172), .Z(n3174) );
  XOR U2528 ( .A(n3183), .B(n3184), .Z(n3172) );
  AND U2529 ( .A(n1059), .B(n3185), .Z(n3184) );
  XOR U2530 ( .A(p_input[840]), .B(n3183), .Z(n3185) );
  XOR U2531 ( .A(n3186), .B(n3187), .Z(n3183) );
  AND U2532 ( .A(n1063), .B(n3188), .Z(n3187) );
  IV U2533 ( .A(n3180), .Z(n3182) );
  XOR U2534 ( .A(n3189), .B(n3190), .Z(n3180) );
  AND U2535 ( .A(n1067), .B(n3191), .Z(n3190) );
  XOR U2536 ( .A(n3192), .B(n3193), .Z(n3178) );
  AND U2537 ( .A(n1071), .B(n3191), .Z(n3193) );
  XNOR U2538 ( .A(n3192), .B(n3189), .Z(n3191) );
  XOR U2539 ( .A(n3194), .B(n3195), .Z(n3189) );
  AND U2540 ( .A(n1074), .B(n3188), .Z(n3195) );
  XNOR U2541 ( .A(n3196), .B(n3186), .Z(n3188) );
  XOR U2542 ( .A(n3197), .B(n3198), .Z(n3186) );
  AND U2543 ( .A(n1078), .B(n3199), .Z(n3198) );
  XOR U2544 ( .A(p_input[856]), .B(n3197), .Z(n3199) );
  XOR U2545 ( .A(n3200), .B(n3201), .Z(n3197) );
  AND U2546 ( .A(n1082), .B(n3202), .Z(n3201) );
  IV U2547 ( .A(n3194), .Z(n3196) );
  XOR U2548 ( .A(n3203), .B(n3204), .Z(n3194) );
  AND U2549 ( .A(n1086), .B(n3205), .Z(n3204) );
  XOR U2550 ( .A(n3206), .B(n3207), .Z(n3192) );
  AND U2551 ( .A(n1090), .B(n3205), .Z(n3207) );
  XNOR U2552 ( .A(n3206), .B(n3203), .Z(n3205) );
  XOR U2553 ( .A(n3208), .B(n3209), .Z(n3203) );
  AND U2554 ( .A(n1093), .B(n3202), .Z(n3209) );
  XNOR U2555 ( .A(n3210), .B(n3200), .Z(n3202) );
  XOR U2556 ( .A(n3211), .B(n3212), .Z(n3200) );
  AND U2557 ( .A(n1097), .B(n3213), .Z(n3212) );
  XOR U2558 ( .A(p_input[872]), .B(n3211), .Z(n3213) );
  XOR U2559 ( .A(n3214), .B(n3215), .Z(n3211) );
  AND U2560 ( .A(n1101), .B(n3216), .Z(n3215) );
  IV U2561 ( .A(n3208), .Z(n3210) );
  XOR U2562 ( .A(n3217), .B(n3218), .Z(n3208) );
  AND U2563 ( .A(n1105), .B(n3219), .Z(n3218) );
  XOR U2564 ( .A(n3220), .B(n3221), .Z(n3206) );
  AND U2565 ( .A(n1109), .B(n3219), .Z(n3221) );
  XNOR U2566 ( .A(n3220), .B(n3217), .Z(n3219) );
  XOR U2567 ( .A(n3222), .B(n3223), .Z(n3217) );
  AND U2568 ( .A(n1112), .B(n3216), .Z(n3223) );
  XNOR U2569 ( .A(n3224), .B(n3214), .Z(n3216) );
  XOR U2570 ( .A(n3225), .B(n3226), .Z(n3214) );
  AND U2571 ( .A(n1116), .B(n3227), .Z(n3226) );
  XOR U2572 ( .A(p_input[888]), .B(n3225), .Z(n3227) );
  XOR U2573 ( .A(n3228), .B(n3229), .Z(n3225) );
  AND U2574 ( .A(n1120), .B(n3230), .Z(n3229) );
  IV U2575 ( .A(n3222), .Z(n3224) );
  XOR U2576 ( .A(n3231), .B(n3232), .Z(n3222) );
  AND U2577 ( .A(n1124), .B(n3233), .Z(n3232) );
  XOR U2578 ( .A(n3234), .B(n3235), .Z(n3220) );
  AND U2579 ( .A(n1128), .B(n3233), .Z(n3235) );
  XNOR U2580 ( .A(n3234), .B(n3231), .Z(n3233) );
  XOR U2581 ( .A(n3236), .B(n3237), .Z(n3231) );
  AND U2582 ( .A(n1131), .B(n3230), .Z(n3237) );
  XNOR U2583 ( .A(n3238), .B(n3228), .Z(n3230) );
  XOR U2584 ( .A(n3239), .B(n3240), .Z(n3228) );
  AND U2585 ( .A(n1135), .B(n3241), .Z(n3240) );
  XOR U2586 ( .A(p_input[904]), .B(n3239), .Z(n3241) );
  XOR U2587 ( .A(n3242), .B(n3243), .Z(n3239) );
  AND U2588 ( .A(n1139), .B(n3244), .Z(n3243) );
  IV U2589 ( .A(n3236), .Z(n3238) );
  XOR U2590 ( .A(n3245), .B(n3246), .Z(n3236) );
  AND U2591 ( .A(n1143), .B(n3247), .Z(n3246) );
  XOR U2592 ( .A(n3248), .B(n3249), .Z(n3234) );
  AND U2593 ( .A(n1147), .B(n3247), .Z(n3249) );
  XNOR U2594 ( .A(n3248), .B(n3245), .Z(n3247) );
  XOR U2595 ( .A(n3250), .B(n3251), .Z(n3245) );
  AND U2596 ( .A(n1150), .B(n3244), .Z(n3251) );
  XNOR U2597 ( .A(n3252), .B(n3242), .Z(n3244) );
  XOR U2598 ( .A(n3253), .B(n3254), .Z(n3242) );
  AND U2599 ( .A(n1154), .B(n3255), .Z(n3254) );
  XOR U2600 ( .A(p_input[920]), .B(n3253), .Z(n3255) );
  XOR U2601 ( .A(n3256), .B(n3257), .Z(n3253) );
  AND U2602 ( .A(n1158), .B(n3258), .Z(n3257) );
  IV U2603 ( .A(n3250), .Z(n3252) );
  XOR U2604 ( .A(n3259), .B(n3260), .Z(n3250) );
  AND U2605 ( .A(n1162), .B(n3261), .Z(n3260) );
  XOR U2606 ( .A(n3262), .B(n3263), .Z(n3248) );
  AND U2607 ( .A(n1166), .B(n3261), .Z(n3263) );
  XNOR U2608 ( .A(n3262), .B(n3259), .Z(n3261) );
  XOR U2609 ( .A(n3264), .B(n3265), .Z(n3259) );
  AND U2610 ( .A(n1169), .B(n3258), .Z(n3265) );
  XNOR U2611 ( .A(n3266), .B(n3256), .Z(n3258) );
  XOR U2612 ( .A(n3267), .B(n3268), .Z(n3256) );
  AND U2613 ( .A(n1173), .B(n3269), .Z(n3268) );
  XOR U2614 ( .A(p_input[936]), .B(n3267), .Z(n3269) );
  XOR U2615 ( .A(n3270), .B(n3271), .Z(n3267) );
  AND U2616 ( .A(n1177), .B(n3272), .Z(n3271) );
  IV U2617 ( .A(n3264), .Z(n3266) );
  XOR U2618 ( .A(n3273), .B(n3274), .Z(n3264) );
  AND U2619 ( .A(n1181), .B(n3275), .Z(n3274) );
  XOR U2620 ( .A(n3276), .B(n3277), .Z(n3262) );
  AND U2621 ( .A(n1185), .B(n3275), .Z(n3277) );
  XNOR U2622 ( .A(n3276), .B(n3273), .Z(n3275) );
  XOR U2623 ( .A(n3278), .B(n3279), .Z(n3273) );
  AND U2624 ( .A(n1188), .B(n3272), .Z(n3279) );
  XNOR U2625 ( .A(n3280), .B(n3270), .Z(n3272) );
  XOR U2626 ( .A(n3281), .B(n3282), .Z(n3270) );
  AND U2627 ( .A(n1192), .B(n3283), .Z(n3282) );
  XOR U2628 ( .A(p_input[952]), .B(n3281), .Z(n3283) );
  XOR U2629 ( .A(n3284), .B(n3285), .Z(n3281) );
  AND U2630 ( .A(n1196), .B(n3286), .Z(n3285) );
  IV U2631 ( .A(n3278), .Z(n3280) );
  XOR U2632 ( .A(n3287), .B(n3288), .Z(n3278) );
  AND U2633 ( .A(n1200), .B(n3289), .Z(n3288) );
  XOR U2634 ( .A(n3290), .B(n3291), .Z(n3276) );
  AND U2635 ( .A(n1204), .B(n3289), .Z(n3291) );
  XNOR U2636 ( .A(n3290), .B(n3287), .Z(n3289) );
  XOR U2637 ( .A(n3292), .B(n3293), .Z(n3287) );
  AND U2638 ( .A(n1207), .B(n3286), .Z(n3293) );
  XNOR U2639 ( .A(n3294), .B(n3284), .Z(n3286) );
  XOR U2640 ( .A(n3295), .B(n3296), .Z(n3284) );
  AND U2641 ( .A(n1211), .B(n3297), .Z(n3296) );
  XOR U2642 ( .A(p_input[968]), .B(n3295), .Z(n3297) );
  XOR U2643 ( .A(n3298), .B(n3299), .Z(n3295) );
  AND U2644 ( .A(n1215), .B(n3300), .Z(n3299) );
  IV U2645 ( .A(n3292), .Z(n3294) );
  XOR U2646 ( .A(n3301), .B(n3302), .Z(n3292) );
  AND U2647 ( .A(n1219), .B(n3303), .Z(n3302) );
  XOR U2648 ( .A(n3304), .B(n3305), .Z(n3290) );
  AND U2649 ( .A(n1223), .B(n3303), .Z(n3305) );
  XNOR U2650 ( .A(n3304), .B(n3301), .Z(n3303) );
  XOR U2651 ( .A(n3306), .B(n3307), .Z(n3301) );
  AND U2652 ( .A(n1226), .B(n3300), .Z(n3307) );
  XNOR U2653 ( .A(n3308), .B(n3298), .Z(n3300) );
  XOR U2654 ( .A(n3309), .B(n3310), .Z(n3298) );
  AND U2655 ( .A(n1230), .B(n3311), .Z(n3310) );
  XOR U2656 ( .A(p_input[984]), .B(n3309), .Z(n3311) );
  XOR U2657 ( .A(n3312), .B(n3313), .Z(n3309) );
  AND U2658 ( .A(n1234), .B(n3314), .Z(n3313) );
  IV U2659 ( .A(n3306), .Z(n3308) );
  XOR U2660 ( .A(n3315), .B(n3316), .Z(n3306) );
  AND U2661 ( .A(n1238), .B(n3317), .Z(n3316) );
  XOR U2662 ( .A(n3318), .B(n3319), .Z(n3304) );
  AND U2663 ( .A(n1242), .B(n3317), .Z(n3319) );
  XNOR U2664 ( .A(n3318), .B(n3315), .Z(n3317) );
  XOR U2665 ( .A(n3320), .B(n3321), .Z(n3315) );
  AND U2666 ( .A(n1245), .B(n3314), .Z(n3321) );
  XNOR U2667 ( .A(n3322), .B(n3312), .Z(n3314) );
  XOR U2668 ( .A(n3323), .B(n3324), .Z(n3312) );
  AND U2669 ( .A(n1249), .B(n3325), .Z(n3324) );
  XOR U2670 ( .A(p_input[1000]), .B(n3323), .Z(n3325) );
  XOR U2671 ( .A(n3326), .B(n3327), .Z(n3323) );
  AND U2672 ( .A(n1253), .B(n3328), .Z(n3327) );
  IV U2673 ( .A(n3320), .Z(n3322) );
  XOR U2674 ( .A(n3329), .B(n3330), .Z(n3320) );
  AND U2675 ( .A(n1257), .B(n3331), .Z(n3330) );
  XOR U2676 ( .A(n3332), .B(n3333), .Z(n3318) );
  AND U2677 ( .A(n1261), .B(n3331), .Z(n3333) );
  XNOR U2678 ( .A(n3332), .B(n3329), .Z(n3331) );
  XOR U2679 ( .A(n3334), .B(n3335), .Z(n3329) );
  AND U2680 ( .A(n1264), .B(n3328), .Z(n3335) );
  XNOR U2681 ( .A(n3336), .B(n3326), .Z(n3328) );
  XOR U2682 ( .A(n3337), .B(n3338), .Z(n3326) );
  AND U2683 ( .A(n1268), .B(n3339), .Z(n3338) );
  XOR U2684 ( .A(p_input[1016]), .B(n3337), .Z(n3339) );
  XOR U2685 ( .A(n3340), .B(n3341), .Z(n3337) );
  AND U2686 ( .A(n1272), .B(n3342), .Z(n3341) );
  IV U2687 ( .A(n3334), .Z(n3336) );
  XOR U2688 ( .A(n3343), .B(n3344), .Z(n3334) );
  AND U2689 ( .A(n1276), .B(n3345), .Z(n3344) );
  XOR U2690 ( .A(n3346), .B(n3347), .Z(n3332) );
  AND U2691 ( .A(n1280), .B(n3345), .Z(n3347) );
  XNOR U2692 ( .A(n3346), .B(n3343), .Z(n3345) );
  XOR U2693 ( .A(n3348), .B(n3349), .Z(n3343) );
  AND U2694 ( .A(n1283), .B(n3342), .Z(n3349) );
  XNOR U2695 ( .A(n3350), .B(n3340), .Z(n3342) );
  XOR U2696 ( .A(n3351), .B(n3352), .Z(n3340) );
  AND U2697 ( .A(n1287), .B(n3353), .Z(n3352) );
  XOR U2698 ( .A(p_input[1032]), .B(n3351), .Z(n3353) );
  XOR U2699 ( .A(n3354), .B(n3355), .Z(n3351) );
  AND U2700 ( .A(n1291), .B(n3356), .Z(n3355) );
  IV U2701 ( .A(n3348), .Z(n3350) );
  XOR U2702 ( .A(n3357), .B(n3358), .Z(n3348) );
  AND U2703 ( .A(n1295), .B(n3359), .Z(n3358) );
  XOR U2704 ( .A(n3360), .B(n3361), .Z(n3346) );
  AND U2705 ( .A(n1299), .B(n3359), .Z(n3361) );
  XNOR U2706 ( .A(n3360), .B(n3357), .Z(n3359) );
  XOR U2707 ( .A(n3362), .B(n3363), .Z(n3357) );
  AND U2708 ( .A(n1302), .B(n3356), .Z(n3363) );
  XNOR U2709 ( .A(n3364), .B(n3354), .Z(n3356) );
  XOR U2710 ( .A(n3365), .B(n3366), .Z(n3354) );
  AND U2711 ( .A(n1306), .B(n3367), .Z(n3366) );
  XOR U2712 ( .A(p_input[1048]), .B(n3365), .Z(n3367) );
  XOR U2713 ( .A(n3368), .B(n3369), .Z(n3365) );
  AND U2714 ( .A(n1310), .B(n3370), .Z(n3369) );
  IV U2715 ( .A(n3362), .Z(n3364) );
  XOR U2716 ( .A(n3371), .B(n3372), .Z(n3362) );
  AND U2717 ( .A(n1314), .B(n3373), .Z(n3372) );
  XOR U2718 ( .A(n3374), .B(n3375), .Z(n3360) );
  AND U2719 ( .A(n1318), .B(n3373), .Z(n3375) );
  XNOR U2720 ( .A(n3374), .B(n3371), .Z(n3373) );
  XOR U2721 ( .A(n3376), .B(n3377), .Z(n3371) );
  AND U2722 ( .A(n1321), .B(n3370), .Z(n3377) );
  XNOR U2723 ( .A(n3378), .B(n3368), .Z(n3370) );
  XOR U2724 ( .A(n3379), .B(n3380), .Z(n3368) );
  AND U2725 ( .A(n1325), .B(n3381), .Z(n3380) );
  XOR U2726 ( .A(p_input[1064]), .B(n3379), .Z(n3381) );
  XOR U2727 ( .A(n3382), .B(n3383), .Z(n3379) );
  AND U2728 ( .A(n1329), .B(n3384), .Z(n3383) );
  IV U2729 ( .A(n3376), .Z(n3378) );
  XOR U2730 ( .A(n3385), .B(n3386), .Z(n3376) );
  AND U2731 ( .A(n1333), .B(n3387), .Z(n3386) );
  XOR U2732 ( .A(n3388), .B(n3389), .Z(n3374) );
  AND U2733 ( .A(n1337), .B(n3387), .Z(n3389) );
  XNOR U2734 ( .A(n3388), .B(n3385), .Z(n3387) );
  XOR U2735 ( .A(n3390), .B(n3391), .Z(n3385) );
  AND U2736 ( .A(n1340), .B(n3384), .Z(n3391) );
  XNOR U2737 ( .A(n3392), .B(n3382), .Z(n3384) );
  XOR U2738 ( .A(n3393), .B(n3394), .Z(n3382) );
  AND U2739 ( .A(n1344), .B(n3395), .Z(n3394) );
  XOR U2740 ( .A(p_input[1080]), .B(n3393), .Z(n3395) );
  XOR U2741 ( .A(n3396), .B(n3397), .Z(n3393) );
  AND U2742 ( .A(n1348), .B(n3398), .Z(n3397) );
  IV U2743 ( .A(n3390), .Z(n3392) );
  XOR U2744 ( .A(n3399), .B(n3400), .Z(n3390) );
  AND U2745 ( .A(n1352), .B(n3401), .Z(n3400) );
  XOR U2746 ( .A(n3402), .B(n3403), .Z(n3388) );
  AND U2747 ( .A(n1356), .B(n3401), .Z(n3403) );
  XNOR U2748 ( .A(n3402), .B(n3399), .Z(n3401) );
  XOR U2749 ( .A(n3404), .B(n3405), .Z(n3399) );
  AND U2750 ( .A(n1359), .B(n3398), .Z(n3405) );
  XNOR U2751 ( .A(n3406), .B(n3396), .Z(n3398) );
  XOR U2752 ( .A(n3407), .B(n3408), .Z(n3396) );
  AND U2753 ( .A(n1363), .B(n3409), .Z(n3408) );
  XOR U2754 ( .A(p_input[1096]), .B(n3407), .Z(n3409) );
  XOR U2755 ( .A(n3410), .B(n3411), .Z(n3407) );
  AND U2756 ( .A(n1367), .B(n3412), .Z(n3411) );
  IV U2757 ( .A(n3404), .Z(n3406) );
  XOR U2758 ( .A(n3413), .B(n3414), .Z(n3404) );
  AND U2759 ( .A(n1371), .B(n3415), .Z(n3414) );
  XOR U2760 ( .A(n3416), .B(n3417), .Z(n3402) );
  AND U2761 ( .A(n1375), .B(n3415), .Z(n3417) );
  XNOR U2762 ( .A(n3416), .B(n3413), .Z(n3415) );
  XOR U2763 ( .A(n3418), .B(n3419), .Z(n3413) );
  AND U2764 ( .A(n1378), .B(n3412), .Z(n3419) );
  XNOR U2765 ( .A(n3420), .B(n3410), .Z(n3412) );
  XOR U2766 ( .A(n3421), .B(n3422), .Z(n3410) );
  AND U2767 ( .A(n1382), .B(n3423), .Z(n3422) );
  XOR U2768 ( .A(p_input[1112]), .B(n3421), .Z(n3423) );
  XOR U2769 ( .A(n3424), .B(n3425), .Z(n3421) );
  AND U2770 ( .A(n1386), .B(n3426), .Z(n3425) );
  IV U2771 ( .A(n3418), .Z(n3420) );
  XOR U2772 ( .A(n3427), .B(n3428), .Z(n3418) );
  AND U2773 ( .A(n1390), .B(n3429), .Z(n3428) );
  XOR U2774 ( .A(n3430), .B(n3431), .Z(n3416) );
  AND U2775 ( .A(n1394), .B(n3429), .Z(n3431) );
  XNOR U2776 ( .A(n3430), .B(n3427), .Z(n3429) );
  XOR U2777 ( .A(n3432), .B(n3433), .Z(n3427) );
  AND U2778 ( .A(n1397), .B(n3426), .Z(n3433) );
  XNOR U2779 ( .A(n3434), .B(n3424), .Z(n3426) );
  XOR U2780 ( .A(n3435), .B(n3436), .Z(n3424) );
  AND U2781 ( .A(n1401), .B(n3437), .Z(n3436) );
  XOR U2782 ( .A(p_input[1128]), .B(n3435), .Z(n3437) );
  XOR U2783 ( .A(n3438), .B(n3439), .Z(n3435) );
  AND U2784 ( .A(n1405), .B(n3440), .Z(n3439) );
  IV U2785 ( .A(n3432), .Z(n3434) );
  XOR U2786 ( .A(n3441), .B(n3442), .Z(n3432) );
  AND U2787 ( .A(n1409), .B(n3443), .Z(n3442) );
  XOR U2788 ( .A(n3444), .B(n3445), .Z(n3430) );
  AND U2789 ( .A(n1413), .B(n3443), .Z(n3445) );
  XNOR U2790 ( .A(n3444), .B(n3441), .Z(n3443) );
  XOR U2791 ( .A(n3446), .B(n3447), .Z(n3441) );
  AND U2792 ( .A(n1416), .B(n3440), .Z(n3447) );
  XNOR U2793 ( .A(n3448), .B(n3438), .Z(n3440) );
  XOR U2794 ( .A(n3449), .B(n3450), .Z(n3438) );
  AND U2795 ( .A(n1420), .B(n3451), .Z(n3450) );
  XOR U2796 ( .A(p_input[1144]), .B(n3449), .Z(n3451) );
  XOR U2797 ( .A(n3452), .B(n3453), .Z(n3449) );
  AND U2798 ( .A(n1424), .B(n3454), .Z(n3453) );
  IV U2799 ( .A(n3446), .Z(n3448) );
  XOR U2800 ( .A(n3455), .B(n3456), .Z(n3446) );
  AND U2801 ( .A(n1428), .B(n3457), .Z(n3456) );
  XOR U2802 ( .A(n3458), .B(n3459), .Z(n3444) );
  AND U2803 ( .A(n1432), .B(n3457), .Z(n3459) );
  XNOR U2804 ( .A(n3458), .B(n3455), .Z(n3457) );
  XOR U2805 ( .A(n3460), .B(n3461), .Z(n3455) );
  AND U2806 ( .A(n1435), .B(n3454), .Z(n3461) );
  XNOR U2807 ( .A(n3462), .B(n3452), .Z(n3454) );
  XOR U2808 ( .A(n3463), .B(n3464), .Z(n3452) );
  AND U2809 ( .A(n1439), .B(n3465), .Z(n3464) );
  XOR U2810 ( .A(p_input[1160]), .B(n3463), .Z(n3465) );
  XOR U2811 ( .A(n3466), .B(n3467), .Z(n3463) );
  AND U2812 ( .A(n1443), .B(n3468), .Z(n3467) );
  IV U2813 ( .A(n3460), .Z(n3462) );
  XOR U2814 ( .A(n3469), .B(n3470), .Z(n3460) );
  AND U2815 ( .A(n1447), .B(n3471), .Z(n3470) );
  XOR U2816 ( .A(n3472), .B(n3473), .Z(n3458) );
  AND U2817 ( .A(n1451), .B(n3471), .Z(n3473) );
  XNOR U2818 ( .A(n3472), .B(n3469), .Z(n3471) );
  XOR U2819 ( .A(n3474), .B(n3475), .Z(n3469) );
  AND U2820 ( .A(n1454), .B(n3468), .Z(n3475) );
  XNOR U2821 ( .A(n3476), .B(n3466), .Z(n3468) );
  XOR U2822 ( .A(n3477), .B(n3478), .Z(n3466) );
  AND U2823 ( .A(n1458), .B(n3479), .Z(n3478) );
  XOR U2824 ( .A(p_input[1176]), .B(n3477), .Z(n3479) );
  XOR U2825 ( .A(n3480), .B(n3481), .Z(n3477) );
  AND U2826 ( .A(n1462), .B(n3482), .Z(n3481) );
  IV U2827 ( .A(n3474), .Z(n3476) );
  XOR U2828 ( .A(n3483), .B(n3484), .Z(n3474) );
  AND U2829 ( .A(n1466), .B(n3485), .Z(n3484) );
  XOR U2830 ( .A(n3486), .B(n3487), .Z(n3472) );
  AND U2831 ( .A(n1470), .B(n3485), .Z(n3487) );
  XNOR U2832 ( .A(n3486), .B(n3483), .Z(n3485) );
  XOR U2833 ( .A(n3488), .B(n3489), .Z(n3483) );
  AND U2834 ( .A(n1473), .B(n3482), .Z(n3489) );
  XNOR U2835 ( .A(n3490), .B(n3480), .Z(n3482) );
  XOR U2836 ( .A(n3491), .B(n3492), .Z(n3480) );
  AND U2837 ( .A(n1477), .B(n3493), .Z(n3492) );
  XOR U2838 ( .A(p_input[1192]), .B(n3491), .Z(n3493) );
  XOR U2839 ( .A(n3494), .B(n3495), .Z(n3491) );
  AND U2840 ( .A(n1481), .B(n3496), .Z(n3495) );
  IV U2841 ( .A(n3488), .Z(n3490) );
  XOR U2842 ( .A(n3497), .B(n3498), .Z(n3488) );
  AND U2843 ( .A(n1485), .B(n3499), .Z(n3498) );
  XOR U2844 ( .A(n3500), .B(n3501), .Z(n3486) );
  AND U2845 ( .A(n1489), .B(n3499), .Z(n3501) );
  XNOR U2846 ( .A(n3500), .B(n3497), .Z(n3499) );
  XOR U2847 ( .A(n3502), .B(n3503), .Z(n3497) );
  AND U2848 ( .A(n1492), .B(n3496), .Z(n3503) );
  XNOR U2849 ( .A(n3504), .B(n3494), .Z(n3496) );
  XOR U2850 ( .A(n3505), .B(n3506), .Z(n3494) );
  AND U2851 ( .A(n1496), .B(n3507), .Z(n3506) );
  XOR U2852 ( .A(p_input[1208]), .B(n3505), .Z(n3507) );
  XOR U2853 ( .A(n3508), .B(n3509), .Z(n3505) );
  AND U2854 ( .A(n1500), .B(n3510), .Z(n3509) );
  IV U2855 ( .A(n3502), .Z(n3504) );
  XOR U2856 ( .A(n3511), .B(n3512), .Z(n3502) );
  AND U2857 ( .A(n1504), .B(n3513), .Z(n3512) );
  XOR U2858 ( .A(n3514), .B(n3515), .Z(n3500) );
  AND U2859 ( .A(n1508), .B(n3513), .Z(n3515) );
  XNOR U2860 ( .A(n3514), .B(n3511), .Z(n3513) );
  XOR U2861 ( .A(n3516), .B(n3517), .Z(n3511) );
  AND U2862 ( .A(n1511), .B(n3510), .Z(n3517) );
  XNOR U2863 ( .A(n3518), .B(n3508), .Z(n3510) );
  XOR U2864 ( .A(n3519), .B(n3520), .Z(n3508) );
  AND U2865 ( .A(n1515), .B(n3521), .Z(n3520) );
  XOR U2866 ( .A(p_input[1224]), .B(n3519), .Z(n3521) );
  XOR U2867 ( .A(n3522), .B(n3523), .Z(n3519) );
  AND U2868 ( .A(n1519), .B(n3524), .Z(n3523) );
  IV U2869 ( .A(n3516), .Z(n3518) );
  XOR U2870 ( .A(n3525), .B(n3526), .Z(n3516) );
  AND U2871 ( .A(n1523), .B(n3527), .Z(n3526) );
  XOR U2872 ( .A(n3528), .B(n3529), .Z(n3514) );
  AND U2873 ( .A(n1527), .B(n3527), .Z(n3529) );
  XNOR U2874 ( .A(n3528), .B(n3525), .Z(n3527) );
  XOR U2875 ( .A(n3530), .B(n3531), .Z(n3525) );
  AND U2876 ( .A(n1530), .B(n3524), .Z(n3531) );
  XNOR U2877 ( .A(n3532), .B(n3522), .Z(n3524) );
  XOR U2878 ( .A(n3533), .B(n3534), .Z(n3522) );
  AND U2879 ( .A(n1534), .B(n3535), .Z(n3534) );
  XOR U2880 ( .A(p_input[1240]), .B(n3533), .Z(n3535) );
  XOR U2881 ( .A(n3536), .B(n3537), .Z(n3533) );
  AND U2882 ( .A(n1538), .B(n3538), .Z(n3537) );
  IV U2883 ( .A(n3530), .Z(n3532) );
  XOR U2884 ( .A(n3539), .B(n3540), .Z(n3530) );
  AND U2885 ( .A(n1542), .B(n3541), .Z(n3540) );
  XOR U2886 ( .A(n3542), .B(n3543), .Z(n3528) );
  AND U2887 ( .A(n1546), .B(n3541), .Z(n3543) );
  XNOR U2888 ( .A(n3542), .B(n3539), .Z(n3541) );
  XOR U2889 ( .A(n3544), .B(n3545), .Z(n3539) );
  AND U2890 ( .A(n1549), .B(n3538), .Z(n3545) );
  XNOR U2891 ( .A(n3546), .B(n3536), .Z(n3538) );
  XOR U2892 ( .A(n3547), .B(n3548), .Z(n3536) );
  AND U2893 ( .A(n1553), .B(n3549), .Z(n3548) );
  XOR U2894 ( .A(p_input[1256]), .B(n3547), .Z(n3549) );
  XOR U2895 ( .A(n3550), .B(n3551), .Z(n3547) );
  AND U2896 ( .A(n1557), .B(n3552), .Z(n3551) );
  IV U2897 ( .A(n3544), .Z(n3546) );
  XOR U2898 ( .A(n3553), .B(n3554), .Z(n3544) );
  AND U2899 ( .A(n1561), .B(n3555), .Z(n3554) );
  XOR U2900 ( .A(n3556), .B(n3557), .Z(n3542) );
  AND U2901 ( .A(n1565), .B(n3555), .Z(n3557) );
  XNOR U2902 ( .A(n3556), .B(n3553), .Z(n3555) );
  XOR U2903 ( .A(n3558), .B(n3559), .Z(n3553) );
  AND U2904 ( .A(n1568), .B(n3552), .Z(n3559) );
  XNOR U2905 ( .A(n3560), .B(n3550), .Z(n3552) );
  XOR U2906 ( .A(n3561), .B(n3562), .Z(n3550) );
  AND U2907 ( .A(n1572), .B(n3563), .Z(n3562) );
  XOR U2908 ( .A(p_input[1272]), .B(n3561), .Z(n3563) );
  XOR U2909 ( .A(n3564), .B(n3565), .Z(n3561) );
  AND U2910 ( .A(n1576), .B(n3566), .Z(n3565) );
  IV U2911 ( .A(n3558), .Z(n3560) );
  XOR U2912 ( .A(n3567), .B(n3568), .Z(n3558) );
  AND U2913 ( .A(n1580), .B(n3569), .Z(n3568) );
  XOR U2914 ( .A(n3570), .B(n3571), .Z(n3556) );
  AND U2915 ( .A(n1584), .B(n3569), .Z(n3571) );
  XNOR U2916 ( .A(n3570), .B(n3567), .Z(n3569) );
  XOR U2917 ( .A(n3572), .B(n3573), .Z(n3567) );
  AND U2918 ( .A(n1587), .B(n3566), .Z(n3573) );
  XNOR U2919 ( .A(n3574), .B(n3564), .Z(n3566) );
  XOR U2920 ( .A(n3575), .B(n3576), .Z(n3564) );
  AND U2921 ( .A(n1591), .B(n3577), .Z(n3576) );
  XOR U2922 ( .A(p_input[1288]), .B(n3575), .Z(n3577) );
  XOR U2923 ( .A(n3578), .B(n3579), .Z(n3575) );
  AND U2924 ( .A(n1595), .B(n3580), .Z(n3579) );
  IV U2925 ( .A(n3572), .Z(n3574) );
  XOR U2926 ( .A(n3581), .B(n3582), .Z(n3572) );
  AND U2927 ( .A(n1599), .B(n3583), .Z(n3582) );
  XOR U2928 ( .A(n3584), .B(n3585), .Z(n3570) );
  AND U2929 ( .A(n1603), .B(n3583), .Z(n3585) );
  XNOR U2930 ( .A(n3584), .B(n3581), .Z(n3583) );
  XOR U2931 ( .A(n3586), .B(n3587), .Z(n3581) );
  AND U2932 ( .A(n1606), .B(n3580), .Z(n3587) );
  XNOR U2933 ( .A(n3588), .B(n3578), .Z(n3580) );
  XOR U2934 ( .A(n3589), .B(n3590), .Z(n3578) );
  AND U2935 ( .A(n1610), .B(n3591), .Z(n3590) );
  XOR U2936 ( .A(p_input[1304]), .B(n3589), .Z(n3591) );
  XOR U2937 ( .A(n3592), .B(n3593), .Z(n3589) );
  AND U2938 ( .A(n1614), .B(n3594), .Z(n3593) );
  IV U2939 ( .A(n3586), .Z(n3588) );
  XOR U2940 ( .A(n3595), .B(n3596), .Z(n3586) );
  AND U2941 ( .A(n1618), .B(n3597), .Z(n3596) );
  XOR U2942 ( .A(n3598), .B(n3599), .Z(n3584) );
  AND U2943 ( .A(n1622), .B(n3597), .Z(n3599) );
  XNOR U2944 ( .A(n3598), .B(n3595), .Z(n3597) );
  XOR U2945 ( .A(n3600), .B(n3601), .Z(n3595) );
  AND U2946 ( .A(n1625), .B(n3594), .Z(n3601) );
  XNOR U2947 ( .A(n3602), .B(n3592), .Z(n3594) );
  XOR U2948 ( .A(n3603), .B(n3604), .Z(n3592) );
  AND U2949 ( .A(n1629), .B(n3605), .Z(n3604) );
  XOR U2950 ( .A(p_input[1320]), .B(n3603), .Z(n3605) );
  XOR U2951 ( .A(n3606), .B(n3607), .Z(n3603) );
  AND U2952 ( .A(n1633), .B(n3608), .Z(n3607) );
  IV U2953 ( .A(n3600), .Z(n3602) );
  XOR U2954 ( .A(n3609), .B(n3610), .Z(n3600) );
  AND U2955 ( .A(n1637), .B(n3611), .Z(n3610) );
  XOR U2956 ( .A(n3612), .B(n3613), .Z(n3598) );
  AND U2957 ( .A(n1641), .B(n3611), .Z(n3613) );
  XNOR U2958 ( .A(n3612), .B(n3609), .Z(n3611) );
  XOR U2959 ( .A(n3614), .B(n3615), .Z(n3609) );
  AND U2960 ( .A(n1644), .B(n3608), .Z(n3615) );
  XNOR U2961 ( .A(n3616), .B(n3606), .Z(n3608) );
  XOR U2962 ( .A(n3617), .B(n3618), .Z(n3606) );
  AND U2963 ( .A(n1648), .B(n3619), .Z(n3618) );
  XOR U2964 ( .A(p_input[1336]), .B(n3617), .Z(n3619) );
  XOR U2965 ( .A(n3620), .B(n3621), .Z(n3617) );
  AND U2966 ( .A(n1652), .B(n3622), .Z(n3621) );
  IV U2967 ( .A(n3614), .Z(n3616) );
  XOR U2968 ( .A(n3623), .B(n3624), .Z(n3614) );
  AND U2969 ( .A(n1656), .B(n3625), .Z(n3624) );
  XOR U2970 ( .A(n3626), .B(n3627), .Z(n3612) );
  AND U2971 ( .A(n1660), .B(n3625), .Z(n3627) );
  XNOR U2972 ( .A(n3626), .B(n3623), .Z(n3625) );
  XOR U2973 ( .A(n3628), .B(n3629), .Z(n3623) );
  AND U2974 ( .A(n1663), .B(n3622), .Z(n3629) );
  XNOR U2975 ( .A(n3630), .B(n3620), .Z(n3622) );
  XOR U2976 ( .A(n3631), .B(n3632), .Z(n3620) );
  AND U2977 ( .A(n1667), .B(n3633), .Z(n3632) );
  XOR U2978 ( .A(p_input[1352]), .B(n3631), .Z(n3633) );
  XOR U2979 ( .A(n3634), .B(n3635), .Z(n3631) );
  AND U2980 ( .A(n1671), .B(n3636), .Z(n3635) );
  IV U2981 ( .A(n3628), .Z(n3630) );
  XOR U2982 ( .A(n3637), .B(n3638), .Z(n3628) );
  AND U2983 ( .A(n1675), .B(n3639), .Z(n3638) );
  XOR U2984 ( .A(n3640), .B(n3641), .Z(n3626) );
  AND U2985 ( .A(n1679), .B(n3639), .Z(n3641) );
  XNOR U2986 ( .A(n3640), .B(n3637), .Z(n3639) );
  XOR U2987 ( .A(n3642), .B(n3643), .Z(n3637) );
  AND U2988 ( .A(n1682), .B(n3636), .Z(n3643) );
  XNOR U2989 ( .A(n3644), .B(n3634), .Z(n3636) );
  XOR U2990 ( .A(n3645), .B(n3646), .Z(n3634) );
  AND U2991 ( .A(n1686), .B(n3647), .Z(n3646) );
  XOR U2992 ( .A(p_input[1368]), .B(n3645), .Z(n3647) );
  XOR U2993 ( .A(n3648), .B(n3649), .Z(n3645) );
  AND U2994 ( .A(n1690), .B(n3650), .Z(n3649) );
  IV U2995 ( .A(n3642), .Z(n3644) );
  XOR U2996 ( .A(n3651), .B(n3652), .Z(n3642) );
  AND U2997 ( .A(n1694), .B(n3653), .Z(n3652) );
  XOR U2998 ( .A(n3654), .B(n3655), .Z(n3640) );
  AND U2999 ( .A(n1698), .B(n3653), .Z(n3655) );
  XNOR U3000 ( .A(n3654), .B(n3651), .Z(n3653) );
  XOR U3001 ( .A(n3656), .B(n3657), .Z(n3651) );
  AND U3002 ( .A(n1701), .B(n3650), .Z(n3657) );
  XNOR U3003 ( .A(n3658), .B(n3648), .Z(n3650) );
  XOR U3004 ( .A(n3659), .B(n3660), .Z(n3648) );
  AND U3005 ( .A(n1705), .B(n3661), .Z(n3660) );
  XOR U3006 ( .A(p_input[1384]), .B(n3659), .Z(n3661) );
  XOR U3007 ( .A(n3662), .B(n3663), .Z(n3659) );
  AND U3008 ( .A(n1709), .B(n3664), .Z(n3663) );
  IV U3009 ( .A(n3656), .Z(n3658) );
  XOR U3010 ( .A(n3665), .B(n3666), .Z(n3656) );
  AND U3011 ( .A(n1713), .B(n3667), .Z(n3666) );
  XOR U3012 ( .A(n3668), .B(n3669), .Z(n3654) );
  AND U3013 ( .A(n1717), .B(n3667), .Z(n3669) );
  XNOR U3014 ( .A(n3668), .B(n3665), .Z(n3667) );
  XOR U3015 ( .A(n3670), .B(n3671), .Z(n3665) );
  AND U3016 ( .A(n1720), .B(n3664), .Z(n3671) );
  XNOR U3017 ( .A(n3672), .B(n3662), .Z(n3664) );
  XOR U3018 ( .A(n3673), .B(n3674), .Z(n3662) );
  AND U3019 ( .A(n1724), .B(n3675), .Z(n3674) );
  XOR U3020 ( .A(p_input[1400]), .B(n3673), .Z(n3675) );
  XOR U3021 ( .A(n3676), .B(n3677), .Z(n3673) );
  AND U3022 ( .A(n1728), .B(n3678), .Z(n3677) );
  IV U3023 ( .A(n3670), .Z(n3672) );
  XOR U3024 ( .A(n3679), .B(n3680), .Z(n3670) );
  AND U3025 ( .A(n1732), .B(n3681), .Z(n3680) );
  XOR U3026 ( .A(n3682), .B(n3683), .Z(n3668) );
  AND U3027 ( .A(n1736), .B(n3681), .Z(n3683) );
  XNOR U3028 ( .A(n3682), .B(n3679), .Z(n3681) );
  XOR U3029 ( .A(n3684), .B(n3685), .Z(n3679) );
  AND U3030 ( .A(n1739), .B(n3678), .Z(n3685) );
  XNOR U3031 ( .A(n3686), .B(n3676), .Z(n3678) );
  XOR U3032 ( .A(n3687), .B(n3688), .Z(n3676) );
  AND U3033 ( .A(n1743), .B(n3689), .Z(n3688) );
  XOR U3034 ( .A(p_input[1416]), .B(n3687), .Z(n3689) );
  XOR U3035 ( .A(n3690), .B(n3691), .Z(n3687) );
  AND U3036 ( .A(n1747), .B(n3692), .Z(n3691) );
  IV U3037 ( .A(n3684), .Z(n3686) );
  XOR U3038 ( .A(n3693), .B(n3694), .Z(n3684) );
  AND U3039 ( .A(n1751), .B(n3695), .Z(n3694) );
  XOR U3040 ( .A(n3696), .B(n3697), .Z(n3682) );
  AND U3041 ( .A(n1755), .B(n3695), .Z(n3697) );
  XNOR U3042 ( .A(n3696), .B(n3693), .Z(n3695) );
  XOR U3043 ( .A(n3698), .B(n3699), .Z(n3693) );
  AND U3044 ( .A(n1758), .B(n3692), .Z(n3699) );
  XNOR U3045 ( .A(n3700), .B(n3690), .Z(n3692) );
  XOR U3046 ( .A(n3701), .B(n3702), .Z(n3690) );
  AND U3047 ( .A(n1762), .B(n3703), .Z(n3702) );
  XOR U3048 ( .A(p_input[1432]), .B(n3701), .Z(n3703) );
  XOR U3049 ( .A(n3704), .B(n3705), .Z(n3701) );
  AND U3050 ( .A(n1766), .B(n3706), .Z(n3705) );
  IV U3051 ( .A(n3698), .Z(n3700) );
  XOR U3052 ( .A(n3707), .B(n3708), .Z(n3698) );
  AND U3053 ( .A(n1770), .B(n3709), .Z(n3708) );
  XOR U3054 ( .A(n3710), .B(n3711), .Z(n3696) );
  AND U3055 ( .A(n1774), .B(n3709), .Z(n3711) );
  XNOR U3056 ( .A(n3710), .B(n3707), .Z(n3709) );
  XOR U3057 ( .A(n3712), .B(n3713), .Z(n3707) );
  AND U3058 ( .A(n1777), .B(n3706), .Z(n3713) );
  XNOR U3059 ( .A(n3714), .B(n3704), .Z(n3706) );
  XOR U3060 ( .A(n3715), .B(n3716), .Z(n3704) );
  AND U3061 ( .A(n1781), .B(n3717), .Z(n3716) );
  XOR U3062 ( .A(p_input[1448]), .B(n3715), .Z(n3717) );
  XOR U3063 ( .A(n3718), .B(n3719), .Z(n3715) );
  AND U3064 ( .A(n1785), .B(n3720), .Z(n3719) );
  IV U3065 ( .A(n3712), .Z(n3714) );
  XOR U3066 ( .A(n3721), .B(n3722), .Z(n3712) );
  AND U3067 ( .A(n1789), .B(n3723), .Z(n3722) );
  XOR U3068 ( .A(n3724), .B(n3725), .Z(n3710) );
  AND U3069 ( .A(n1793), .B(n3723), .Z(n3725) );
  XNOR U3070 ( .A(n3724), .B(n3721), .Z(n3723) );
  XOR U3071 ( .A(n3726), .B(n3727), .Z(n3721) );
  AND U3072 ( .A(n1796), .B(n3720), .Z(n3727) );
  XNOR U3073 ( .A(n3728), .B(n3718), .Z(n3720) );
  XOR U3074 ( .A(n3729), .B(n3730), .Z(n3718) );
  AND U3075 ( .A(n1800), .B(n3731), .Z(n3730) );
  XOR U3076 ( .A(p_input[1464]), .B(n3729), .Z(n3731) );
  XOR U3077 ( .A(n3732), .B(n3733), .Z(n3729) );
  AND U3078 ( .A(n1804), .B(n3734), .Z(n3733) );
  IV U3079 ( .A(n3726), .Z(n3728) );
  XOR U3080 ( .A(n3735), .B(n3736), .Z(n3726) );
  AND U3081 ( .A(n1808), .B(n3737), .Z(n3736) );
  XOR U3082 ( .A(n3738), .B(n3739), .Z(n3724) );
  AND U3083 ( .A(n1812), .B(n3737), .Z(n3739) );
  XNOR U3084 ( .A(n3738), .B(n3735), .Z(n3737) );
  XOR U3085 ( .A(n3740), .B(n3741), .Z(n3735) );
  AND U3086 ( .A(n1815), .B(n3734), .Z(n3741) );
  XNOR U3087 ( .A(n3742), .B(n3732), .Z(n3734) );
  XOR U3088 ( .A(n3743), .B(n3744), .Z(n3732) );
  AND U3089 ( .A(n1819), .B(n3745), .Z(n3744) );
  XOR U3090 ( .A(p_input[1480]), .B(n3743), .Z(n3745) );
  XOR U3091 ( .A(n3746), .B(n3747), .Z(n3743) );
  AND U3092 ( .A(n1823), .B(n3748), .Z(n3747) );
  IV U3093 ( .A(n3740), .Z(n3742) );
  XOR U3094 ( .A(n3749), .B(n3750), .Z(n3740) );
  AND U3095 ( .A(n1827), .B(n3751), .Z(n3750) );
  XOR U3096 ( .A(n3752), .B(n3753), .Z(n3738) );
  AND U3097 ( .A(n1831), .B(n3751), .Z(n3753) );
  XNOR U3098 ( .A(n3752), .B(n3749), .Z(n3751) );
  XOR U3099 ( .A(n3754), .B(n3755), .Z(n3749) );
  AND U3100 ( .A(n1834), .B(n3748), .Z(n3755) );
  XNOR U3101 ( .A(n3756), .B(n3746), .Z(n3748) );
  XOR U3102 ( .A(n3757), .B(n3758), .Z(n3746) );
  AND U3103 ( .A(n1838), .B(n3759), .Z(n3758) );
  XOR U3104 ( .A(p_input[1496]), .B(n3757), .Z(n3759) );
  XOR U3105 ( .A(n3760), .B(n3761), .Z(n3757) );
  AND U3106 ( .A(n1842), .B(n3762), .Z(n3761) );
  IV U3107 ( .A(n3754), .Z(n3756) );
  XOR U3108 ( .A(n3763), .B(n3764), .Z(n3754) );
  AND U3109 ( .A(n1846), .B(n3765), .Z(n3764) );
  XOR U3110 ( .A(n3766), .B(n3767), .Z(n3752) );
  AND U3111 ( .A(n1850), .B(n3765), .Z(n3767) );
  XNOR U3112 ( .A(n3766), .B(n3763), .Z(n3765) );
  XOR U3113 ( .A(n3768), .B(n3769), .Z(n3763) );
  AND U3114 ( .A(n1853), .B(n3762), .Z(n3769) );
  XNOR U3115 ( .A(n3770), .B(n3760), .Z(n3762) );
  XOR U3116 ( .A(n3771), .B(n3772), .Z(n3760) );
  AND U3117 ( .A(n1857), .B(n3773), .Z(n3772) );
  XOR U3118 ( .A(p_input[1512]), .B(n3771), .Z(n3773) );
  XOR U3119 ( .A(n3774), .B(n3775), .Z(n3771) );
  AND U3120 ( .A(n1861), .B(n3776), .Z(n3775) );
  IV U3121 ( .A(n3768), .Z(n3770) );
  XOR U3122 ( .A(n3777), .B(n3778), .Z(n3768) );
  AND U3123 ( .A(n1865), .B(n3779), .Z(n3778) );
  XOR U3124 ( .A(n3780), .B(n3781), .Z(n3766) );
  AND U3125 ( .A(n1869), .B(n3779), .Z(n3781) );
  XNOR U3126 ( .A(n3780), .B(n3777), .Z(n3779) );
  XOR U3127 ( .A(n3782), .B(n3783), .Z(n3777) );
  AND U3128 ( .A(n1872), .B(n3776), .Z(n3783) );
  XNOR U3129 ( .A(n3784), .B(n3774), .Z(n3776) );
  XOR U3130 ( .A(n3785), .B(n3786), .Z(n3774) );
  AND U3131 ( .A(n1876), .B(n3787), .Z(n3786) );
  XOR U3132 ( .A(p_input[1528]), .B(n3785), .Z(n3787) );
  XOR U3133 ( .A(n3788), .B(n3789), .Z(n3785) );
  AND U3134 ( .A(n1880), .B(n3790), .Z(n3789) );
  IV U3135 ( .A(n3782), .Z(n3784) );
  XOR U3136 ( .A(n3791), .B(n3792), .Z(n3782) );
  AND U3137 ( .A(n1884), .B(n3793), .Z(n3792) );
  XOR U3138 ( .A(n3794), .B(n3795), .Z(n3780) );
  AND U3139 ( .A(n1888), .B(n3793), .Z(n3795) );
  XNOR U3140 ( .A(n3794), .B(n3791), .Z(n3793) );
  XOR U3141 ( .A(n3796), .B(n3797), .Z(n3791) );
  AND U3142 ( .A(n1891), .B(n3790), .Z(n3797) );
  XNOR U3143 ( .A(n3798), .B(n3788), .Z(n3790) );
  XOR U3144 ( .A(n3799), .B(n3800), .Z(n3788) );
  AND U3145 ( .A(n1895), .B(n3801), .Z(n3800) );
  XOR U3146 ( .A(p_input[1544]), .B(n3799), .Z(n3801) );
  XOR U3147 ( .A(n3802), .B(n3803), .Z(n3799) );
  AND U3148 ( .A(n1899), .B(n3804), .Z(n3803) );
  IV U3149 ( .A(n3796), .Z(n3798) );
  XOR U3150 ( .A(n3805), .B(n3806), .Z(n3796) );
  AND U3151 ( .A(n1903), .B(n3807), .Z(n3806) );
  XOR U3152 ( .A(n3808), .B(n3809), .Z(n3794) );
  AND U3153 ( .A(n1907), .B(n3807), .Z(n3809) );
  XNOR U3154 ( .A(n3808), .B(n3805), .Z(n3807) );
  XOR U3155 ( .A(n3810), .B(n3811), .Z(n3805) );
  AND U3156 ( .A(n1910), .B(n3804), .Z(n3811) );
  XNOR U3157 ( .A(n3812), .B(n3802), .Z(n3804) );
  XOR U3158 ( .A(n3813), .B(n3814), .Z(n3802) );
  AND U3159 ( .A(n1914), .B(n3815), .Z(n3814) );
  XOR U3160 ( .A(p_input[1560]), .B(n3813), .Z(n3815) );
  XOR U3161 ( .A(n3816), .B(n3817), .Z(n3813) );
  AND U3162 ( .A(n1918), .B(n3818), .Z(n3817) );
  IV U3163 ( .A(n3810), .Z(n3812) );
  XOR U3164 ( .A(n3819), .B(n3820), .Z(n3810) );
  AND U3165 ( .A(n1922), .B(n3821), .Z(n3820) );
  XOR U3166 ( .A(n3822), .B(n3823), .Z(n3808) );
  AND U3167 ( .A(n1926), .B(n3821), .Z(n3823) );
  XNOR U3168 ( .A(n3822), .B(n3819), .Z(n3821) );
  XOR U3169 ( .A(n3824), .B(n3825), .Z(n3819) );
  AND U3170 ( .A(n1929), .B(n3818), .Z(n3825) );
  XNOR U3171 ( .A(n3826), .B(n3816), .Z(n3818) );
  XOR U3172 ( .A(n3827), .B(n3828), .Z(n3816) );
  AND U3173 ( .A(n1933), .B(n3829), .Z(n3828) );
  XOR U3174 ( .A(p_input[1576]), .B(n3827), .Z(n3829) );
  XOR U3175 ( .A(n3830), .B(n3831), .Z(n3827) );
  AND U3176 ( .A(n1937), .B(n3832), .Z(n3831) );
  IV U3177 ( .A(n3824), .Z(n3826) );
  XOR U3178 ( .A(n3833), .B(n3834), .Z(n3824) );
  AND U3179 ( .A(n1941), .B(n3835), .Z(n3834) );
  XOR U3180 ( .A(n3836), .B(n3837), .Z(n3822) );
  AND U3181 ( .A(n1945), .B(n3835), .Z(n3837) );
  XNOR U3182 ( .A(n3836), .B(n3833), .Z(n3835) );
  XOR U3183 ( .A(n3838), .B(n3839), .Z(n3833) );
  AND U3184 ( .A(n1948), .B(n3832), .Z(n3839) );
  XNOR U3185 ( .A(n3840), .B(n3830), .Z(n3832) );
  XOR U3186 ( .A(n3841), .B(n3842), .Z(n3830) );
  AND U3187 ( .A(n1952), .B(n3843), .Z(n3842) );
  XOR U3188 ( .A(p_input[1592]), .B(n3841), .Z(n3843) );
  XOR U3189 ( .A(n3844), .B(n3845), .Z(n3841) );
  AND U3190 ( .A(n1956), .B(n3846), .Z(n3845) );
  IV U3191 ( .A(n3838), .Z(n3840) );
  XOR U3192 ( .A(n3847), .B(n3848), .Z(n3838) );
  AND U3193 ( .A(n1960), .B(n3849), .Z(n3848) );
  XOR U3194 ( .A(n3850), .B(n3851), .Z(n3836) );
  AND U3195 ( .A(n1964), .B(n3849), .Z(n3851) );
  XNOR U3196 ( .A(n3850), .B(n3847), .Z(n3849) );
  XOR U3197 ( .A(n3852), .B(n3853), .Z(n3847) );
  AND U3198 ( .A(n1967), .B(n3846), .Z(n3853) );
  XNOR U3199 ( .A(n3854), .B(n3844), .Z(n3846) );
  XOR U3200 ( .A(n3855), .B(n3856), .Z(n3844) );
  AND U3201 ( .A(n1971), .B(n3857), .Z(n3856) );
  XOR U3202 ( .A(p_input[1608]), .B(n3855), .Z(n3857) );
  XOR U3203 ( .A(n3858), .B(n3859), .Z(n3855) );
  AND U3204 ( .A(n1975), .B(n3860), .Z(n3859) );
  IV U3205 ( .A(n3852), .Z(n3854) );
  XOR U3206 ( .A(n3861), .B(n3862), .Z(n3852) );
  AND U3207 ( .A(n1979), .B(n3863), .Z(n3862) );
  XOR U3208 ( .A(n3864), .B(n3865), .Z(n3850) );
  AND U3209 ( .A(n1983), .B(n3863), .Z(n3865) );
  XNOR U3210 ( .A(n3864), .B(n3861), .Z(n3863) );
  XOR U3211 ( .A(n3866), .B(n3867), .Z(n3861) );
  AND U3212 ( .A(n1986), .B(n3860), .Z(n3867) );
  XNOR U3213 ( .A(n3868), .B(n3858), .Z(n3860) );
  XOR U3214 ( .A(n3869), .B(n3870), .Z(n3858) );
  AND U3215 ( .A(n1990), .B(n3871), .Z(n3870) );
  XOR U3216 ( .A(p_input[1624]), .B(n3869), .Z(n3871) );
  XOR U3217 ( .A(n3872), .B(n3873), .Z(n3869) );
  AND U3218 ( .A(n1994), .B(n3874), .Z(n3873) );
  IV U3219 ( .A(n3866), .Z(n3868) );
  XOR U3220 ( .A(n3875), .B(n3876), .Z(n3866) );
  AND U3221 ( .A(n1998), .B(n3877), .Z(n3876) );
  XOR U3222 ( .A(n3878), .B(n3879), .Z(n3864) );
  AND U3223 ( .A(n2002), .B(n3877), .Z(n3879) );
  XNOR U3224 ( .A(n3878), .B(n3875), .Z(n3877) );
  XOR U3225 ( .A(n3880), .B(n3881), .Z(n3875) );
  AND U3226 ( .A(n2005), .B(n3874), .Z(n3881) );
  XNOR U3227 ( .A(n3882), .B(n3872), .Z(n3874) );
  XOR U3228 ( .A(n3883), .B(n3884), .Z(n3872) );
  AND U3229 ( .A(n2009), .B(n3885), .Z(n3884) );
  XOR U3230 ( .A(p_input[1640]), .B(n3883), .Z(n3885) );
  XOR U3231 ( .A(n3886), .B(n3887), .Z(n3883) );
  AND U3232 ( .A(n2013), .B(n3888), .Z(n3887) );
  IV U3233 ( .A(n3880), .Z(n3882) );
  XOR U3234 ( .A(n3889), .B(n3890), .Z(n3880) );
  AND U3235 ( .A(n2017), .B(n3891), .Z(n3890) );
  XOR U3236 ( .A(n3892), .B(n3893), .Z(n3878) );
  AND U3237 ( .A(n2021), .B(n3891), .Z(n3893) );
  XNOR U3238 ( .A(n3892), .B(n3889), .Z(n3891) );
  XOR U3239 ( .A(n3894), .B(n3895), .Z(n3889) );
  AND U3240 ( .A(n2024), .B(n3888), .Z(n3895) );
  XNOR U3241 ( .A(n3896), .B(n3886), .Z(n3888) );
  XOR U3242 ( .A(n3897), .B(n3898), .Z(n3886) );
  AND U3243 ( .A(n2028), .B(n3899), .Z(n3898) );
  XOR U3244 ( .A(p_input[1656]), .B(n3897), .Z(n3899) );
  XOR U3245 ( .A(n3900), .B(n3901), .Z(n3897) );
  AND U3246 ( .A(n2032), .B(n3902), .Z(n3901) );
  IV U3247 ( .A(n3894), .Z(n3896) );
  XOR U3248 ( .A(n3903), .B(n3904), .Z(n3894) );
  AND U3249 ( .A(n2036), .B(n3905), .Z(n3904) );
  XOR U3250 ( .A(n3906), .B(n3907), .Z(n3892) );
  AND U3251 ( .A(n2040), .B(n3905), .Z(n3907) );
  XNOR U3252 ( .A(n3906), .B(n3903), .Z(n3905) );
  XOR U3253 ( .A(n3908), .B(n3909), .Z(n3903) );
  AND U3254 ( .A(n2043), .B(n3902), .Z(n3909) );
  XNOR U3255 ( .A(n3910), .B(n3900), .Z(n3902) );
  XOR U3256 ( .A(n3911), .B(n3912), .Z(n3900) );
  AND U3257 ( .A(n2047), .B(n3913), .Z(n3912) );
  XOR U3258 ( .A(p_input[1672]), .B(n3911), .Z(n3913) );
  XOR U3259 ( .A(n3914), .B(n3915), .Z(n3911) );
  AND U3260 ( .A(n2051), .B(n3916), .Z(n3915) );
  IV U3261 ( .A(n3908), .Z(n3910) );
  XOR U3262 ( .A(n3917), .B(n3918), .Z(n3908) );
  AND U3263 ( .A(n2055), .B(n3919), .Z(n3918) );
  XOR U3264 ( .A(n3920), .B(n3921), .Z(n3906) );
  AND U3265 ( .A(n2059), .B(n3919), .Z(n3921) );
  XNOR U3266 ( .A(n3920), .B(n3917), .Z(n3919) );
  XOR U3267 ( .A(n3922), .B(n3923), .Z(n3917) );
  AND U3268 ( .A(n2062), .B(n3916), .Z(n3923) );
  XNOR U3269 ( .A(n3924), .B(n3914), .Z(n3916) );
  XOR U3270 ( .A(n3925), .B(n3926), .Z(n3914) );
  AND U3271 ( .A(n2066), .B(n3927), .Z(n3926) );
  XOR U3272 ( .A(p_input[1688]), .B(n3925), .Z(n3927) );
  XOR U3273 ( .A(n3928), .B(n3929), .Z(n3925) );
  AND U3274 ( .A(n2070), .B(n3930), .Z(n3929) );
  IV U3275 ( .A(n3922), .Z(n3924) );
  XOR U3276 ( .A(n3931), .B(n3932), .Z(n3922) );
  AND U3277 ( .A(n2074), .B(n3933), .Z(n3932) );
  XOR U3278 ( .A(n3934), .B(n3935), .Z(n3920) );
  AND U3279 ( .A(n2078), .B(n3933), .Z(n3935) );
  XNOR U3280 ( .A(n3934), .B(n3931), .Z(n3933) );
  XOR U3281 ( .A(n3936), .B(n3937), .Z(n3931) );
  AND U3282 ( .A(n2081), .B(n3930), .Z(n3937) );
  XNOR U3283 ( .A(n3938), .B(n3928), .Z(n3930) );
  XOR U3284 ( .A(n3939), .B(n3940), .Z(n3928) );
  AND U3285 ( .A(n2085), .B(n3941), .Z(n3940) );
  XOR U3286 ( .A(p_input[1704]), .B(n3939), .Z(n3941) );
  XOR U3287 ( .A(n3942), .B(n3943), .Z(n3939) );
  AND U3288 ( .A(n2089), .B(n3944), .Z(n3943) );
  IV U3289 ( .A(n3936), .Z(n3938) );
  XOR U3290 ( .A(n3945), .B(n3946), .Z(n3936) );
  AND U3291 ( .A(n2093), .B(n3947), .Z(n3946) );
  XOR U3292 ( .A(n3948), .B(n3949), .Z(n3934) );
  AND U3293 ( .A(n2097), .B(n3947), .Z(n3949) );
  XNOR U3294 ( .A(n3948), .B(n3945), .Z(n3947) );
  XOR U3295 ( .A(n3950), .B(n3951), .Z(n3945) );
  AND U3296 ( .A(n2100), .B(n3944), .Z(n3951) );
  XNOR U3297 ( .A(n3952), .B(n3942), .Z(n3944) );
  XOR U3298 ( .A(n3953), .B(n3954), .Z(n3942) );
  AND U3299 ( .A(n2104), .B(n3955), .Z(n3954) );
  XOR U3300 ( .A(p_input[1720]), .B(n3953), .Z(n3955) );
  XOR U3301 ( .A(n3956), .B(n3957), .Z(n3953) );
  AND U3302 ( .A(n2108), .B(n3958), .Z(n3957) );
  IV U3303 ( .A(n3950), .Z(n3952) );
  XOR U3304 ( .A(n3959), .B(n3960), .Z(n3950) );
  AND U3305 ( .A(n2112), .B(n3961), .Z(n3960) );
  XOR U3306 ( .A(n3962), .B(n3963), .Z(n3948) );
  AND U3307 ( .A(n2116), .B(n3961), .Z(n3963) );
  XNOR U3308 ( .A(n3962), .B(n3959), .Z(n3961) );
  XOR U3309 ( .A(n3964), .B(n3965), .Z(n3959) );
  AND U3310 ( .A(n2119), .B(n3958), .Z(n3965) );
  XNOR U3311 ( .A(n3966), .B(n3956), .Z(n3958) );
  XOR U3312 ( .A(n3967), .B(n3968), .Z(n3956) );
  AND U3313 ( .A(n2123), .B(n3969), .Z(n3968) );
  XOR U3314 ( .A(p_input[1736]), .B(n3967), .Z(n3969) );
  XOR U3315 ( .A(n3970), .B(n3971), .Z(n3967) );
  AND U3316 ( .A(n2127), .B(n3972), .Z(n3971) );
  IV U3317 ( .A(n3964), .Z(n3966) );
  XOR U3318 ( .A(n3973), .B(n3974), .Z(n3964) );
  AND U3319 ( .A(n2131), .B(n3975), .Z(n3974) );
  XOR U3320 ( .A(n3976), .B(n3977), .Z(n3962) );
  AND U3321 ( .A(n2135), .B(n3975), .Z(n3977) );
  XNOR U3322 ( .A(n3976), .B(n3973), .Z(n3975) );
  XOR U3323 ( .A(n3978), .B(n3979), .Z(n3973) );
  AND U3324 ( .A(n2138), .B(n3972), .Z(n3979) );
  XNOR U3325 ( .A(n3980), .B(n3970), .Z(n3972) );
  XOR U3326 ( .A(n3981), .B(n3982), .Z(n3970) );
  AND U3327 ( .A(n2142), .B(n3983), .Z(n3982) );
  XOR U3328 ( .A(p_input[1752]), .B(n3981), .Z(n3983) );
  XOR U3329 ( .A(n3984), .B(n3985), .Z(n3981) );
  AND U3330 ( .A(n2146), .B(n3986), .Z(n3985) );
  IV U3331 ( .A(n3978), .Z(n3980) );
  XOR U3332 ( .A(n3987), .B(n3988), .Z(n3978) );
  AND U3333 ( .A(n2150), .B(n3989), .Z(n3988) );
  XOR U3334 ( .A(n3990), .B(n3991), .Z(n3976) );
  AND U3335 ( .A(n2154), .B(n3989), .Z(n3991) );
  XNOR U3336 ( .A(n3990), .B(n3987), .Z(n3989) );
  XOR U3337 ( .A(n3992), .B(n3993), .Z(n3987) );
  AND U3338 ( .A(n2157), .B(n3986), .Z(n3993) );
  XNOR U3339 ( .A(n3994), .B(n3984), .Z(n3986) );
  XOR U3340 ( .A(n3995), .B(n3996), .Z(n3984) );
  AND U3341 ( .A(n2161), .B(n3997), .Z(n3996) );
  XOR U3342 ( .A(p_input[1768]), .B(n3995), .Z(n3997) );
  XOR U3343 ( .A(n3998), .B(n3999), .Z(n3995) );
  AND U3344 ( .A(n2165), .B(n4000), .Z(n3999) );
  IV U3345 ( .A(n3992), .Z(n3994) );
  XOR U3346 ( .A(n4001), .B(n4002), .Z(n3992) );
  AND U3347 ( .A(n2169), .B(n4003), .Z(n4002) );
  XOR U3348 ( .A(n4004), .B(n4005), .Z(n3990) );
  AND U3349 ( .A(n2173), .B(n4003), .Z(n4005) );
  XNOR U3350 ( .A(n4004), .B(n4001), .Z(n4003) );
  XOR U3351 ( .A(n4006), .B(n4007), .Z(n4001) );
  AND U3352 ( .A(n2176), .B(n4000), .Z(n4007) );
  XNOR U3353 ( .A(n4008), .B(n3998), .Z(n4000) );
  XOR U3354 ( .A(n4009), .B(n4010), .Z(n3998) );
  AND U3355 ( .A(n2180), .B(n4011), .Z(n4010) );
  XOR U3356 ( .A(p_input[1784]), .B(n4009), .Z(n4011) );
  XOR U3357 ( .A(n4012), .B(n4013), .Z(n4009) );
  AND U3358 ( .A(n2184), .B(n4014), .Z(n4013) );
  IV U3359 ( .A(n4006), .Z(n4008) );
  XOR U3360 ( .A(n4015), .B(n4016), .Z(n4006) );
  AND U3361 ( .A(n2188), .B(n4017), .Z(n4016) );
  XOR U3362 ( .A(n4018), .B(n4019), .Z(n4004) );
  AND U3363 ( .A(n2192), .B(n4017), .Z(n4019) );
  XNOR U3364 ( .A(n4018), .B(n4015), .Z(n4017) );
  XOR U3365 ( .A(n4020), .B(n4021), .Z(n4015) );
  AND U3366 ( .A(n2195), .B(n4014), .Z(n4021) );
  XNOR U3367 ( .A(n4022), .B(n4012), .Z(n4014) );
  XOR U3368 ( .A(n4023), .B(n4024), .Z(n4012) );
  AND U3369 ( .A(n2199), .B(n4025), .Z(n4024) );
  XOR U3370 ( .A(p_input[1800]), .B(n4023), .Z(n4025) );
  XOR U3371 ( .A(n4026), .B(n4027), .Z(n4023) );
  AND U3372 ( .A(n2203), .B(n4028), .Z(n4027) );
  IV U3373 ( .A(n4020), .Z(n4022) );
  XOR U3374 ( .A(n4029), .B(n4030), .Z(n4020) );
  AND U3375 ( .A(n2207), .B(n4031), .Z(n4030) );
  XOR U3376 ( .A(n4032), .B(n4033), .Z(n4018) );
  AND U3377 ( .A(n2211), .B(n4031), .Z(n4033) );
  XNOR U3378 ( .A(n4032), .B(n4029), .Z(n4031) );
  XOR U3379 ( .A(n4034), .B(n4035), .Z(n4029) );
  AND U3380 ( .A(n2214), .B(n4028), .Z(n4035) );
  XNOR U3381 ( .A(n4036), .B(n4026), .Z(n4028) );
  XOR U3382 ( .A(n4037), .B(n4038), .Z(n4026) );
  AND U3383 ( .A(n2218), .B(n4039), .Z(n4038) );
  XOR U3384 ( .A(p_input[1816]), .B(n4037), .Z(n4039) );
  XOR U3385 ( .A(n4040), .B(n4041), .Z(n4037) );
  AND U3386 ( .A(n2222), .B(n4042), .Z(n4041) );
  IV U3387 ( .A(n4034), .Z(n4036) );
  XOR U3388 ( .A(n4043), .B(n4044), .Z(n4034) );
  AND U3389 ( .A(n2226), .B(n4045), .Z(n4044) );
  XOR U3390 ( .A(n4046), .B(n4047), .Z(n4032) );
  AND U3391 ( .A(n2230), .B(n4045), .Z(n4047) );
  XNOR U3392 ( .A(n4046), .B(n4043), .Z(n4045) );
  XOR U3393 ( .A(n4048), .B(n4049), .Z(n4043) );
  AND U3394 ( .A(n2233), .B(n4042), .Z(n4049) );
  XNOR U3395 ( .A(n4050), .B(n4040), .Z(n4042) );
  XOR U3396 ( .A(n4051), .B(n4052), .Z(n4040) );
  AND U3397 ( .A(n2237), .B(n4053), .Z(n4052) );
  XOR U3398 ( .A(p_input[1832]), .B(n4051), .Z(n4053) );
  XOR U3399 ( .A(n4054), .B(n4055), .Z(n4051) );
  AND U3400 ( .A(n2241), .B(n4056), .Z(n4055) );
  IV U3401 ( .A(n4048), .Z(n4050) );
  XOR U3402 ( .A(n4057), .B(n4058), .Z(n4048) );
  AND U3403 ( .A(n2245), .B(n4059), .Z(n4058) );
  XOR U3404 ( .A(n4060), .B(n4061), .Z(n4046) );
  AND U3405 ( .A(n2249), .B(n4059), .Z(n4061) );
  XNOR U3406 ( .A(n4060), .B(n4057), .Z(n4059) );
  XOR U3407 ( .A(n4062), .B(n4063), .Z(n4057) );
  AND U3408 ( .A(n2252), .B(n4056), .Z(n4063) );
  XNOR U3409 ( .A(n4064), .B(n4054), .Z(n4056) );
  XOR U3410 ( .A(n4065), .B(n4066), .Z(n4054) );
  AND U3411 ( .A(n2256), .B(n4067), .Z(n4066) );
  XOR U3412 ( .A(p_input[1848]), .B(n4065), .Z(n4067) );
  XOR U3413 ( .A(n4068), .B(n4069), .Z(n4065) );
  AND U3414 ( .A(n2260), .B(n4070), .Z(n4069) );
  IV U3415 ( .A(n4062), .Z(n4064) );
  XOR U3416 ( .A(n4071), .B(n4072), .Z(n4062) );
  AND U3417 ( .A(n2264), .B(n4073), .Z(n4072) );
  XOR U3418 ( .A(n4074), .B(n4075), .Z(n4060) );
  AND U3419 ( .A(n2268), .B(n4073), .Z(n4075) );
  XNOR U3420 ( .A(n4074), .B(n4071), .Z(n4073) );
  XOR U3421 ( .A(n4076), .B(n4077), .Z(n4071) );
  AND U3422 ( .A(n2271), .B(n4070), .Z(n4077) );
  XNOR U3423 ( .A(n4078), .B(n4068), .Z(n4070) );
  XOR U3424 ( .A(n4079), .B(n4080), .Z(n4068) );
  AND U3425 ( .A(n2275), .B(n4081), .Z(n4080) );
  XOR U3426 ( .A(p_input[1864]), .B(n4079), .Z(n4081) );
  XOR U3427 ( .A(n4082), .B(n4083), .Z(n4079) );
  AND U3428 ( .A(n2279), .B(n4084), .Z(n4083) );
  IV U3429 ( .A(n4076), .Z(n4078) );
  XOR U3430 ( .A(n4085), .B(n4086), .Z(n4076) );
  AND U3431 ( .A(n2283), .B(n4087), .Z(n4086) );
  XOR U3432 ( .A(n4088), .B(n4089), .Z(n4074) );
  AND U3433 ( .A(n2287), .B(n4087), .Z(n4089) );
  XNOR U3434 ( .A(n4088), .B(n4085), .Z(n4087) );
  XOR U3435 ( .A(n4090), .B(n4091), .Z(n4085) );
  AND U3436 ( .A(n2290), .B(n4084), .Z(n4091) );
  XNOR U3437 ( .A(n4092), .B(n4082), .Z(n4084) );
  XOR U3438 ( .A(n4093), .B(n4094), .Z(n4082) );
  AND U3439 ( .A(n2294), .B(n4095), .Z(n4094) );
  XOR U3440 ( .A(p_input[1880]), .B(n4093), .Z(n4095) );
  XOR U3441 ( .A(n4096), .B(n4097), .Z(n4093) );
  AND U3442 ( .A(n2298), .B(n4098), .Z(n4097) );
  IV U3443 ( .A(n4090), .Z(n4092) );
  XOR U3444 ( .A(n4099), .B(n4100), .Z(n4090) );
  AND U3445 ( .A(n2302), .B(n4101), .Z(n4100) );
  XOR U3446 ( .A(n4102), .B(n4103), .Z(n4088) );
  AND U3447 ( .A(n2306), .B(n4101), .Z(n4103) );
  XNOR U3448 ( .A(n4102), .B(n4099), .Z(n4101) );
  XOR U3449 ( .A(n4104), .B(n4105), .Z(n4099) );
  AND U3450 ( .A(n2309), .B(n4098), .Z(n4105) );
  XNOR U3451 ( .A(n4106), .B(n4096), .Z(n4098) );
  XOR U3452 ( .A(n4107), .B(n4108), .Z(n4096) );
  AND U3453 ( .A(n2313), .B(n4109), .Z(n4108) );
  XOR U3454 ( .A(p_input[1896]), .B(n4107), .Z(n4109) );
  XOR U3455 ( .A(n4110), .B(n4111), .Z(n4107) );
  AND U3456 ( .A(n2317), .B(n4112), .Z(n4111) );
  IV U3457 ( .A(n4104), .Z(n4106) );
  XOR U3458 ( .A(n4113), .B(n4114), .Z(n4104) );
  AND U3459 ( .A(n2321), .B(n4115), .Z(n4114) );
  XOR U3460 ( .A(n4116), .B(n4117), .Z(n4102) );
  AND U3461 ( .A(n2325), .B(n4115), .Z(n4117) );
  XNOR U3462 ( .A(n4116), .B(n4113), .Z(n4115) );
  XOR U3463 ( .A(n4118), .B(n4119), .Z(n4113) );
  AND U3464 ( .A(n2328), .B(n4112), .Z(n4119) );
  XNOR U3465 ( .A(n4120), .B(n4110), .Z(n4112) );
  XOR U3466 ( .A(n4121), .B(n4122), .Z(n4110) );
  AND U3467 ( .A(n2332), .B(n4123), .Z(n4122) );
  XOR U3468 ( .A(p_input[1912]), .B(n4121), .Z(n4123) );
  XOR U3469 ( .A(n4124), .B(n4125), .Z(n4121) );
  AND U3470 ( .A(n2336), .B(n4126), .Z(n4125) );
  IV U3471 ( .A(n4118), .Z(n4120) );
  XOR U3472 ( .A(n4127), .B(n4128), .Z(n4118) );
  AND U3473 ( .A(n2340), .B(n4129), .Z(n4128) );
  XOR U3474 ( .A(n4130), .B(n4131), .Z(n4116) );
  AND U3475 ( .A(n2344), .B(n4129), .Z(n4131) );
  XNOR U3476 ( .A(n4130), .B(n4127), .Z(n4129) );
  XOR U3477 ( .A(n4132), .B(n4133), .Z(n4127) );
  AND U3478 ( .A(n2347), .B(n4126), .Z(n4133) );
  XNOR U3479 ( .A(n4134), .B(n4124), .Z(n4126) );
  XOR U3480 ( .A(n4135), .B(n4136), .Z(n4124) );
  AND U3481 ( .A(n2351), .B(n4137), .Z(n4136) );
  XOR U3482 ( .A(p_input[1928]), .B(n4135), .Z(n4137) );
  XOR U3483 ( .A(n4138), .B(n4139), .Z(n4135) );
  AND U3484 ( .A(n2355), .B(n4140), .Z(n4139) );
  IV U3485 ( .A(n4132), .Z(n4134) );
  XOR U3486 ( .A(n4141), .B(n4142), .Z(n4132) );
  AND U3487 ( .A(n2359), .B(n4143), .Z(n4142) );
  XOR U3488 ( .A(n4144), .B(n4145), .Z(n4130) );
  AND U3489 ( .A(n2363), .B(n4143), .Z(n4145) );
  XNOR U3490 ( .A(n4144), .B(n4141), .Z(n4143) );
  XOR U3491 ( .A(n4146), .B(n4147), .Z(n4141) );
  AND U3492 ( .A(n2366), .B(n4140), .Z(n4147) );
  XNOR U3493 ( .A(n4148), .B(n4138), .Z(n4140) );
  XOR U3494 ( .A(n4149), .B(n4150), .Z(n4138) );
  AND U3495 ( .A(n2370), .B(n4151), .Z(n4150) );
  XOR U3496 ( .A(p_input[1944]), .B(n4149), .Z(n4151) );
  XOR U3497 ( .A(n4152), .B(n4153), .Z(n4149) );
  AND U3498 ( .A(n2374), .B(n4154), .Z(n4153) );
  IV U3499 ( .A(n4146), .Z(n4148) );
  XOR U3500 ( .A(n4155), .B(n4156), .Z(n4146) );
  AND U3501 ( .A(n2378), .B(n4157), .Z(n4156) );
  XOR U3502 ( .A(n4158), .B(n4159), .Z(n4144) );
  AND U3503 ( .A(n2382), .B(n4157), .Z(n4159) );
  XNOR U3504 ( .A(n4158), .B(n4155), .Z(n4157) );
  XOR U3505 ( .A(n4160), .B(n4161), .Z(n4155) );
  AND U3506 ( .A(n2385), .B(n4154), .Z(n4161) );
  XNOR U3507 ( .A(n4162), .B(n4152), .Z(n4154) );
  XOR U3508 ( .A(n4163), .B(n4164), .Z(n4152) );
  AND U3509 ( .A(n2389), .B(n4165), .Z(n4164) );
  XOR U3510 ( .A(p_input[1960]), .B(n4163), .Z(n4165) );
  XOR U3511 ( .A(n4166), .B(n4167), .Z(n4163) );
  AND U3512 ( .A(n2393), .B(n4168), .Z(n4167) );
  IV U3513 ( .A(n4160), .Z(n4162) );
  XOR U3514 ( .A(n4169), .B(n4170), .Z(n4160) );
  AND U3515 ( .A(n2397), .B(n4171), .Z(n4170) );
  XOR U3516 ( .A(n4172), .B(n4173), .Z(n4158) );
  AND U3517 ( .A(n2401), .B(n4171), .Z(n4173) );
  XNOR U3518 ( .A(n4172), .B(n4169), .Z(n4171) );
  XOR U3519 ( .A(n4174), .B(n4175), .Z(n4169) );
  AND U3520 ( .A(n2404), .B(n4168), .Z(n4175) );
  XNOR U3521 ( .A(n4176), .B(n4166), .Z(n4168) );
  XOR U3522 ( .A(n4177), .B(n4178), .Z(n4166) );
  AND U3523 ( .A(n2408), .B(n4179), .Z(n4178) );
  XOR U3524 ( .A(p_input[1976]), .B(n4177), .Z(n4179) );
  XOR U3525 ( .A(n4180), .B(n4181), .Z(n4177) );
  AND U3526 ( .A(n2412), .B(n4182), .Z(n4181) );
  IV U3527 ( .A(n4174), .Z(n4176) );
  XOR U3528 ( .A(n4183), .B(n4184), .Z(n4174) );
  AND U3529 ( .A(n2416), .B(n4185), .Z(n4184) );
  XOR U3530 ( .A(n4186), .B(n4187), .Z(n4172) );
  AND U3531 ( .A(n2420), .B(n4185), .Z(n4187) );
  XNOR U3532 ( .A(n4186), .B(n4183), .Z(n4185) );
  XOR U3533 ( .A(n4188), .B(n4189), .Z(n4183) );
  AND U3534 ( .A(n2423), .B(n4182), .Z(n4189) );
  XNOR U3535 ( .A(n4190), .B(n4180), .Z(n4182) );
  XOR U3536 ( .A(n4191), .B(n4192), .Z(n4180) );
  AND U3537 ( .A(n2427), .B(n4193), .Z(n4192) );
  XOR U3538 ( .A(p_input[1992]), .B(n4191), .Z(n4193) );
  XOR U3539 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n4194), 
        .Z(n4191) );
  AND U3540 ( .A(n2430), .B(n4195), .Z(n4194) );
  IV U3541 ( .A(n4188), .Z(n4190) );
  XOR U3542 ( .A(n4196), .B(n4197), .Z(n4188) );
  AND U3543 ( .A(n2434), .B(n4198), .Z(n4197) );
  XOR U3544 ( .A(n4199), .B(n4200), .Z(n4186) );
  AND U3545 ( .A(n2438), .B(n4198), .Z(n4200) );
  XNOR U3546 ( .A(n4199), .B(n4196), .Z(n4198) );
  XNOR U3547 ( .A(n4201), .B(n4202), .Z(n4196) );
  AND U3548 ( .A(n2441), .B(n4195), .Z(n4202) );
  XNOR U3549 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n4201), 
        .Z(n4195) );
  XNOR U3550 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n4203), 
        .Z(n4201) );
  AND U3551 ( .A(n2443), .B(n4204), .Z(n4203) );
  XNOR U3552 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n4205), .Z(n4199) );
  AND U3553 ( .A(n2446), .B(n4204), .Z(n4205) );
  XOR U3554 ( .A(n4206), .B(n4207), .Z(n4204) );
  XOR U3555 ( .A(n5), .B(n4208), .Z(o[23]) );
  AND U3556 ( .A(n62), .B(n4209), .Z(n5) );
  XOR U3557 ( .A(n6), .B(n4208), .Z(n4209) );
  XOR U3558 ( .A(n4210), .B(n31), .Z(n4208) );
  AND U3559 ( .A(n65), .B(n4211), .Z(n31) );
  XNOR U3560 ( .A(n4212), .B(n32), .Z(n4211) );
  XOR U3561 ( .A(n4213), .B(n4214), .Z(n32) );
  AND U3562 ( .A(n70), .B(n4215), .Z(n4214) );
  XOR U3563 ( .A(p_input[7]), .B(n4213), .Z(n4215) );
  XOR U3564 ( .A(n4216), .B(n4217), .Z(n4213) );
  AND U3565 ( .A(n74), .B(n4218), .Z(n4217) );
  IV U3566 ( .A(n4210), .Z(n4212) );
  XOR U3567 ( .A(n4219), .B(n4220), .Z(n4210) );
  AND U3568 ( .A(n78), .B(n4221), .Z(n4220) );
  XOR U3569 ( .A(n4222), .B(n4223), .Z(n6) );
  AND U3570 ( .A(n82), .B(n4221), .Z(n4223) );
  XNOR U3571 ( .A(n4224), .B(n4219), .Z(n4221) );
  XOR U3572 ( .A(n4225), .B(n4226), .Z(n4219) );
  AND U3573 ( .A(n86), .B(n4218), .Z(n4226) );
  XNOR U3574 ( .A(n4227), .B(n4216), .Z(n4218) );
  XOR U3575 ( .A(n4228), .B(n4229), .Z(n4216) );
  AND U3576 ( .A(n90), .B(n4230), .Z(n4229) );
  XOR U3577 ( .A(p_input[23]), .B(n4228), .Z(n4230) );
  XOR U3578 ( .A(n4231), .B(n4232), .Z(n4228) );
  AND U3579 ( .A(n94), .B(n4233), .Z(n4232) );
  IV U3580 ( .A(n4225), .Z(n4227) );
  XOR U3581 ( .A(n4234), .B(n4235), .Z(n4225) );
  AND U3582 ( .A(n98), .B(n4236), .Z(n4235) );
  IV U3583 ( .A(n4222), .Z(n4224) );
  XNOR U3584 ( .A(n4237), .B(n4238), .Z(n4222) );
  AND U3585 ( .A(n102), .B(n4236), .Z(n4238) );
  XNOR U3586 ( .A(n4237), .B(n4234), .Z(n4236) );
  XOR U3587 ( .A(n4239), .B(n4240), .Z(n4234) );
  AND U3588 ( .A(n105), .B(n4233), .Z(n4240) );
  XNOR U3589 ( .A(n4241), .B(n4231), .Z(n4233) );
  XOR U3590 ( .A(n4242), .B(n4243), .Z(n4231) );
  AND U3591 ( .A(n109), .B(n4244), .Z(n4243) );
  XOR U3592 ( .A(p_input[39]), .B(n4242), .Z(n4244) );
  XOR U3593 ( .A(n4245), .B(n4246), .Z(n4242) );
  AND U3594 ( .A(n113), .B(n4247), .Z(n4246) );
  IV U3595 ( .A(n4239), .Z(n4241) );
  XOR U3596 ( .A(n4248), .B(n4249), .Z(n4239) );
  AND U3597 ( .A(n117), .B(n4250), .Z(n4249) );
  XOR U3598 ( .A(n4251), .B(n4252), .Z(n4237) );
  AND U3599 ( .A(n121), .B(n4250), .Z(n4252) );
  XNOR U3600 ( .A(n4251), .B(n4248), .Z(n4250) );
  XOR U3601 ( .A(n4253), .B(n4254), .Z(n4248) );
  AND U3602 ( .A(n124), .B(n4247), .Z(n4254) );
  XNOR U3603 ( .A(n4255), .B(n4245), .Z(n4247) );
  XOR U3604 ( .A(n4256), .B(n4257), .Z(n4245) );
  AND U3605 ( .A(n128), .B(n4258), .Z(n4257) );
  XOR U3606 ( .A(p_input[55]), .B(n4256), .Z(n4258) );
  XOR U3607 ( .A(n4259), .B(n4260), .Z(n4256) );
  AND U3608 ( .A(n132), .B(n4261), .Z(n4260) );
  IV U3609 ( .A(n4253), .Z(n4255) );
  XOR U3610 ( .A(n4262), .B(n4263), .Z(n4253) );
  AND U3611 ( .A(n136), .B(n4264), .Z(n4263) );
  XOR U3612 ( .A(n4265), .B(n4266), .Z(n4251) );
  AND U3613 ( .A(n140), .B(n4264), .Z(n4266) );
  XNOR U3614 ( .A(n4265), .B(n4262), .Z(n4264) );
  XOR U3615 ( .A(n4267), .B(n4268), .Z(n4262) );
  AND U3616 ( .A(n143), .B(n4261), .Z(n4268) );
  XNOR U3617 ( .A(n4269), .B(n4259), .Z(n4261) );
  XOR U3618 ( .A(n4270), .B(n4271), .Z(n4259) );
  AND U3619 ( .A(n147), .B(n4272), .Z(n4271) );
  XOR U3620 ( .A(p_input[71]), .B(n4270), .Z(n4272) );
  XOR U3621 ( .A(n4273), .B(n4274), .Z(n4270) );
  AND U3622 ( .A(n151), .B(n4275), .Z(n4274) );
  IV U3623 ( .A(n4267), .Z(n4269) );
  XOR U3624 ( .A(n4276), .B(n4277), .Z(n4267) );
  AND U3625 ( .A(n155), .B(n4278), .Z(n4277) );
  XOR U3626 ( .A(n4279), .B(n4280), .Z(n4265) );
  AND U3627 ( .A(n159), .B(n4278), .Z(n4280) );
  XNOR U3628 ( .A(n4279), .B(n4276), .Z(n4278) );
  XOR U3629 ( .A(n4281), .B(n4282), .Z(n4276) );
  AND U3630 ( .A(n162), .B(n4275), .Z(n4282) );
  XNOR U3631 ( .A(n4283), .B(n4273), .Z(n4275) );
  XOR U3632 ( .A(n4284), .B(n4285), .Z(n4273) );
  AND U3633 ( .A(n166), .B(n4286), .Z(n4285) );
  XOR U3634 ( .A(p_input[87]), .B(n4284), .Z(n4286) );
  XOR U3635 ( .A(n4287), .B(n4288), .Z(n4284) );
  AND U3636 ( .A(n170), .B(n4289), .Z(n4288) );
  IV U3637 ( .A(n4281), .Z(n4283) );
  XOR U3638 ( .A(n4290), .B(n4291), .Z(n4281) );
  AND U3639 ( .A(n174), .B(n4292), .Z(n4291) );
  XOR U3640 ( .A(n4293), .B(n4294), .Z(n4279) );
  AND U3641 ( .A(n178), .B(n4292), .Z(n4294) );
  XNOR U3642 ( .A(n4293), .B(n4290), .Z(n4292) );
  XOR U3643 ( .A(n4295), .B(n4296), .Z(n4290) );
  AND U3644 ( .A(n181), .B(n4289), .Z(n4296) );
  XNOR U3645 ( .A(n4297), .B(n4287), .Z(n4289) );
  XOR U3646 ( .A(n4298), .B(n4299), .Z(n4287) );
  AND U3647 ( .A(n185), .B(n4300), .Z(n4299) );
  XOR U3648 ( .A(p_input[103]), .B(n4298), .Z(n4300) );
  XOR U3649 ( .A(n4301), .B(n4302), .Z(n4298) );
  AND U3650 ( .A(n189), .B(n4303), .Z(n4302) );
  IV U3651 ( .A(n4295), .Z(n4297) );
  XOR U3652 ( .A(n4304), .B(n4305), .Z(n4295) );
  AND U3653 ( .A(n193), .B(n4306), .Z(n4305) );
  XOR U3654 ( .A(n4307), .B(n4308), .Z(n4293) );
  AND U3655 ( .A(n197), .B(n4306), .Z(n4308) );
  XNOR U3656 ( .A(n4307), .B(n4304), .Z(n4306) );
  XOR U3657 ( .A(n4309), .B(n4310), .Z(n4304) );
  AND U3658 ( .A(n200), .B(n4303), .Z(n4310) );
  XNOR U3659 ( .A(n4311), .B(n4301), .Z(n4303) );
  XOR U3660 ( .A(n4312), .B(n4313), .Z(n4301) );
  AND U3661 ( .A(n204), .B(n4314), .Z(n4313) );
  XOR U3662 ( .A(p_input[119]), .B(n4312), .Z(n4314) );
  XOR U3663 ( .A(n4315), .B(n4316), .Z(n4312) );
  AND U3664 ( .A(n208), .B(n4317), .Z(n4316) );
  IV U3665 ( .A(n4309), .Z(n4311) );
  XOR U3666 ( .A(n4318), .B(n4319), .Z(n4309) );
  AND U3667 ( .A(n212), .B(n4320), .Z(n4319) );
  XOR U3668 ( .A(n4321), .B(n4322), .Z(n4307) );
  AND U3669 ( .A(n216), .B(n4320), .Z(n4322) );
  XNOR U3670 ( .A(n4321), .B(n4318), .Z(n4320) );
  XOR U3671 ( .A(n4323), .B(n4324), .Z(n4318) );
  AND U3672 ( .A(n219), .B(n4317), .Z(n4324) );
  XNOR U3673 ( .A(n4325), .B(n4315), .Z(n4317) );
  XOR U3674 ( .A(n4326), .B(n4327), .Z(n4315) );
  AND U3675 ( .A(n223), .B(n4328), .Z(n4327) );
  XOR U3676 ( .A(p_input[135]), .B(n4326), .Z(n4328) );
  XOR U3677 ( .A(n4329), .B(n4330), .Z(n4326) );
  AND U3678 ( .A(n227), .B(n4331), .Z(n4330) );
  IV U3679 ( .A(n4323), .Z(n4325) );
  XOR U3680 ( .A(n4332), .B(n4333), .Z(n4323) );
  AND U3681 ( .A(n231), .B(n4334), .Z(n4333) );
  XOR U3682 ( .A(n4335), .B(n4336), .Z(n4321) );
  AND U3683 ( .A(n235), .B(n4334), .Z(n4336) );
  XNOR U3684 ( .A(n4335), .B(n4332), .Z(n4334) );
  XOR U3685 ( .A(n4337), .B(n4338), .Z(n4332) );
  AND U3686 ( .A(n238), .B(n4331), .Z(n4338) );
  XNOR U3687 ( .A(n4339), .B(n4329), .Z(n4331) );
  XOR U3688 ( .A(n4340), .B(n4341), .Z(n4329) );
  AND U3689 ( .A(n242), .B(n4342), .Z(n4341) );
  XOR U3690 ( .A(p_input[151]), .B(n4340), .Z(n4342) );
  XOR U3691 ( .A(n4343), .B(n4344), .Z(n4340) );
  AND U3692 ( .A(n246), .B(n4345), .Z(n4344) );
  IV U3693 ( .A(n4337), .Z(n4339) );
  XOR U3694 ( .A(n4346), .B(n4347), .Z(n4337) );
  AND U3695 ( .A(n250), .B(n4348), .Z(n4347) );
  XOR U3696 ( .A(n4349), .B(n4350), .Z(n4335) );
  AND U3697 ( .A(n254), .B(n4348), .Z(n4350) );
  XNOR U3698 ( .A(n4349), .B(n4346), .Z(n4348) );
  XOR U3699 ( .A(n4351), .B(n4352), .Z(n4346) );
  AND U3700 ( .A(n257), .B(n4345), .Z(n4352) );
  XNOR U3701 ( .A(n4353), .B(n4343), .Z(n4345) );
  XOR U3702 ( .A(n4354), .B(n4355), .Z(n4343) );
  AND U3703 ( .A(n261), .B(n4356), .Z(n4355) );
  XOR U3704 ( .A(p_input[167]), .B(n4354), .Z(n4356) );
  XOR U3705 ( .A(n4357), .B(n4358), .Z(n4354) );
  AND U3706 ( .A(n265), .B(n4359), .Z(n4358) );
  IV U3707 ( .A(n4351), .Z(n4353) );
  XOR U3708 ( .A(n4360), .B(n4361), .Z(n4351) );
  AND U3709 ( .A(n269), .B(n4362), .Z(n4361) );
  XOR U3710 ( .A(n4363), .B(n4364), .Z(n4349) );
  AND U3711 ( .A(n273), .B(n4362), .Z(n4364) );
  XNOR U3712 ( .A(n4363), .B(n4360), .Z(n4362) );
  XOR U3713 ( .A(n4365), .B(n4366), .Z(n4360) );
  AND U3714 ( .A(n276), .B(n4359), .Z(n4366) );
  XNOR U3715 ( .A(n4367), .B(n4357), .Z(n4359) );
  XOR U3716 ( .A(n4368), .B(n4369), .Z(n4357) );
  AND U3717 ( .A(n280), .B(n4370), .Z(n4369) );
  XOR U3718 ( .A(p_input[183]), .B(n4368), .Z(n4370) );
  XOR U3719 ( .A(n4371), .B(n4372), .Z(n4368) );
  AND U3720 ( .A(n284), .B(n4373), .Z(n4372) );
  IV U3721 ( .A(n4365), .Z(n4367) );
  XOR U3722 ( .A(n4374), .B(n4375), .Z(n4365) );
  AND U3723 ( .A(n288), .B(n4376), .Z(n4375) );
  XOR U3724 ( .A(n4377), .B(n4378), .Z(n4363) );
  AND U3725 ( .A(n292), .B(n4376), .Z(n4378) );
  XNOR U3726 ( .A(n4377), .B(n4374), .Z(n4376) );
  XOR U3727 ( .A(n4379), .B(n4380), .Z(n4374) );
  AND U3728 ( .A(n295), .B(n4373), .Z(n4380) );
  XNOR U3729 ( .A(n4381), .B(n4371), .Z(n4373) );
  XOR U3730 ( .A(n4382), .B(n4383), .Z(n4371) );
  AND U3731 ( .A(n299), .B(n4384), .Z(n4383) );
  XOR U3732 ( .A(p_input[199]), .B(n4382), .Z(n4384) );
  XOR U3733 ( .A(n4385), .B(n4386), .Z(n4382) );
  AND U3734 ( .A(n303), .B(n4387), .Z(n4386) );
  IV U3735 ( .A(n4379), .Z(n4381) );
  XOR U3736 ( .A(n4388), .B(n4389), .Z(n4379) );
  AND U3737 ( .A(n307), .B(n4390), .Z(n4389) );
  XOR U3738 ( .A(n4391), .B(n4392), .Z(n4377) );
  AND U3739 ( .A(n311), .B(n4390), .Z(n4392) );
  XNOR U3740 ( .A(n4391), .B(n4388), .Z(n4390) );
  XOR U3741 ( .A(n4393), .B(n4394), .Z(n4388) );
  AND U3742 ( .A(n314), .B(n4387), .Z(n4394) );
  XNOR U3743 ( .A(n4395), .B(n4385), .Z(n4387) );
  XOR U3744 ( .A(n4396), .B(n4397), .Z(n4385) );
  AND U3745 ( .A(n318), .B(n4398), .Z(n4397) );
  XOR U3746 ( .A(p_input[215]), .B(n4396), .Z(n4398) );
  XOR U3747 ( .A(n4399), .B(n4400), .Z(n4396) );
  AND U3748 ( .A(n322), .B(n4401), .Z(n4400) );
  IV U3749 ( .A(n4393), .Z(n4395) );
  XOR U3750 ( .A(n4402), .B(n4403), .Z(n4393) );
  AND U3751 ( .A(n326), .B(n4404), .Z(n4403) );
  XOR U3752 ( .A(n4405), .B(n4406), .Z(n4391) );
  AND U3753 ( .A(n330), .B(n4404), .Z(n4406) );
  XNOR U3754 ( .A(n4405), .B(n4402), .Z(n4404) );
  XOR U3755 ( .A(n4407), .B(n4408), .Z(n4402) );
  AND U3756 ( .A(n333), .B(n4401), .Z(n4408) );
  XNOR U3757 ( .A(n4409), .B(n4399), .Z(n4401) );
  XOR U3758 ( .A(n4410), .B(n4411), .Z(n4399) );
  AND U3759 ( .A(n337), .B(n4412), .Z(n4411) );
  XOR U3760 ( .A(p_input[231]), .B(n4410), .Z(n4412) );
  XOR U3761 ( .A(n4413), .B(n4414), .Z(n4410) );
  AND U3762 ( .A(n341), .B(n4415), .Z(n4414) );
  IV U3763 ( .A(n4407), .Z(n4409) );
  XOR U3764 ( .A(n4416), .B(n4417), .Z(n4407) );
  AND U3765 ( .A(n345), .B(n4418), .Z(n4417) );
  XOR U3766 ( .A(n4419), .B(n4420), .Z(n4405) );
  AND U3767 ( .A(n349), .B(n4418), .Z(n4420) );
  XNOR U3768 ( .A(n4419), .B(n4416), .Z(n4418) );
  XOR U3769 ( .A(n4421), .B(n4422), .Z(n4416) );
  AND U3770 ( .A(n352), .B(n4415), .Z(n4422) );
  XNOR U3771 ( .A(n4423), .B(n4413), .Z(n4415) );
  XOR U3772 ( .A(n4424), .B(n4425), .Z(n4413) );
  AND U3773 ( .A(n356), .B(n4426), .Z(n4425) );
  XOR U3774 ( .A(p_input[247]), .B(n4424), .Z(n4426) );
  XOR U3775 ( .A(n4427), .B(n4428), .Z(n4424) );
  AND U3776 ( .A(n360), .B(n4429), .Z(n4428) );
  IV U3777 ( .A(n4421), .Z(n4423) );
  XOR U3778 ( .A(n4430), .B(n4431), .Z(n4421) );
  AND U3779 ( .A(n364), .B(n4432), .Z(n4431) );
  XOR U3780 ( .A(n4433), .B(n4434), .Z(n4419) );
  AND U3781 ( .A(n368), .B(n4432), .Z(n4434) );
  XNOR U3782 ( .A(n4433), .B(n4430), .Z(n4432) );
  XOR U3783 ( .A(n4435), .B(n4436), .Z(n4430) );
  AND U3784 ( .A(n371), .B(n4429), .Z(n4436) );
  XNOR U3785 ( .A(n4437), .B(n4427), .Z(n4429) );
  XOR U3786 ( .A(n4438), .B(n4439), .Z(n4427) );
  AND U3787 ( .A(n375), .B(n4440), .Z(n4439) );
  XOR U3788 ( .A(p_input[263]), .B(n4438), .Z(n4440) );
  XOR U3789 ( .A(n4441), .B(n4442), .Z(n4438) );
  AND U3790 ( .A(n379), .B(n4443), .Z(n4442) );
  IV U3791 ( .A(n4435), .Z(n4437) );
  XOR U3792 ( .A(n4444), .B(n4445), .Z(n4435) );
  AND U3793 ( .A(n383), .B(n4446), .Z(n4445) );
  XOR U3794 ( .A(n4447), .B(n4448), .Z(n4433) );
  AND U3795 ( .A(n387), .B(n4446), .Z(n4448) );
  XNOR U3796 ( .A(n4447), .B(n4444), .Z(n4446) );
  XOR U3797 ( .A(n4449), .B(n4450), .Z(n4444) );
  AND U3798 ( .A(n390), .B(n4443), .Z(n4450) );
  XNOR U3799 ( .A(n4451), .B(n4441), .Z(n4443) );
  XOR U3800 ( .A(n4452), .B(n4453), .Z(n4441) );
  AND U3801 ( .A(n394), .B(n4454), .Z(n4453) );
  XOR U3802 ( .A(p_input[279]), .B(n4452), .Z(n4454) );
  XOR U3803 ( .A(n4455), .B(n4456), .Z(n4452) );
  AND U3804 ( .A(n398), .B(n4457), .Z(n4456) );
  IV U3805 ( .A(n4449), .Z(n4451) );
  XOR U3806 ( .A(n4458), .B(n4459), .Z(n4449) );
  AND U3807 ( .A(n402), .B(n4460), .Z(n4459) );
  XOR U3808 ( .A(n4461), .B(n4462), .Z(n4447) );
  AND U3809 ( .A(n406), .B(n4460), .Z(n4462) );
  XNOR U3810 ( .A(n4461), .B(n4458), .Z(n4460) );
  XOR U3811 ( .A(n4463), .B(n4464), .Z(n4458) );
  AND U3812 ( .A(n409), .B(n4457), .Z(n4464) );
  XNOR U3813 ( .A(n4465), .B(n4455), .Z(n4457) );
  XOR U3814 ( .A(n4466), .B(n4467), .Z(n4455) );
  AND U3815 ( .A(n413), .B(n4468), .Z(n4467) );
  XOR U3816 ( .A(p_input[295]), .B(n4466), .Z(n4468) );
  XOR U3817 ( .A(n4469), .B(n4470), .Z(n4466) );
  AND U3818 ( .A(n417), .B(n4471), .Z(n4470) );
  IV U3819 ( .A(n4463), .Z(n4465) );
  XOR U3820 ( .A(n4472), .B(n4473), .Z(n4463) );
  AND U3821 ( .A(n421), .B(n4474), .Z(n4473) );
  XOR U3822 ( .A(n4475), .B(n4476), .Z(n4461) );
  AND U3823 ( .A(n425), .B(n4474), .Z(n4476) );
  XNOR U3824 ( .A(n4475), .B(n4472), .Z(n4474) );
  XOR U3825 ( .A(n4477), .B(n4478), .Z(n4472) );
  AND U3826 ( .A(n428), .B(n4471), .Z(n4478) );
  XNOR U3827 ( .A(n4479), .B(n4469), .Z(n4471) );
  XOR U3828 ( .A(n4480), .B(n4481), .Z(n4469) );
  AND U3829 ( .A(n432), .B(n4482), .Z(n4481) );
  XOR U3830 ( .A(p_input[311]), .B(n4480), .Z(n4482) );
  XOR U3831 ( .A(n4483), .B(n4484), .Z(n4480) );
  AND U3832 ( .A(n436), .B(n4485), .Z(n4484) );
  IV U3833 ( .A(n4477), .Z(n4479) );
  XOR U3834 ( .A(n4486), .B(n4487), .Z(n4477) );
  AND U3835 ( .A(n440), .B(n4488), .Z(n4487) );
  XOR U3836 ( .A(n4489), .B(n4490), .Z(n4475) );
  AND U3837 ( .A(n444), .B(n4488), .Z(n4490) );
  XNOR U3838 ( .A(n4489), .B(n4486), .Z(n4488) );
  XOR U3839 ( .A(n4491), .B(n4492), .Z(n4486) );
  AND U3840 ( .A(n447), .B(n4485), .Z(n4492) );
  XNOR U3841 ( .A(n4493), .B(n4483), .Z(n4485) );
  XOR U3842 ( .A(n4494), .B(n4495), .Z(n4483) );
  AND U3843 ( .A(n451), .B(n4496), .Z(n4495) );
  XOR U3844 ( .A(p_input[327]), .B(n4494), .Z(n4496) );
  XOR U3845 ( .A(n4497), .B(n4498), .Z(n4494) );
  AND U3846 ( .A(n455), .B(n4499), .Z(n4498) );
  IV U3847 ( .A(n4491), .Z(n4493) );
  XOR U3848 ( .A(n4500), .B(n4501), .Z(n4491) );
  AND U3849 ( .A(n459), .B(n4502), .Z(n4501) );
  XOR U3850 ( .A(n4503), .B(n4504), .Z(n4489) );
  AND U3851 ( .A(n463), .B(n4502), .Z(n4504) );
  XNOR U3852 ( .A(n4503), .B(n4500), .Z(n4502) );
  XOR U3853 ( .A(n4505), .B(n4506), .Z(n4500) );
  AND U3854 ( .A(n466), .B(n4499), .Z(n4506) );
  XNOR U3855 ( .A(n4507), .B(n4497), .Z(n4499) );
  XOR U3856 ( .A(n4508), .B(n4509), .Z(n4497) );
  AND U3857 ( .A(n470), .B(n4510), .Z(n4509) );
  XOR U3858 ( .A(p_input[343]), .B(n4508), .Z(n4510) );
  XOR U3859 ( .A(n4511), .B(n4512), .Z(n4508) );
  AND U3860 ( .A(n474), .B(n4513), .Z(n4512) );
  IV U3861 ( .A(n4505), .Z(n4507) );
  XOR U3862 ( .A(n4514), .B(n4515), .Z(n4505) );
  AND U3863 ( .A(n478), .B(n4516), .Z(n4515) );
  XOR U3864 ( .A(n4517), .B(n4518), .Z(n4503) );
  AND U3865 ( .A(n482), .B(n4516), .Z(n4518) );
  XNOR U3866 ( .A(n4517), .B(n4514), .Z(n4516) );
  XOR U3867 ( .A(n4519), .B(n4520), .Z(n4514) );
  AND U3868 ( .A(n485), .B(n4513), .Z(n4520) );
  XNOR U3869 ( .A(n4521), .B(n4511), .Z(n4513) );
  XOR U3870 ( .A(n4522), .B(n4523), .Z(n4511) );
  AND U3871 ( .A(n489), .B(n4524), .Z(n4523) );
  XOR U3872 ( .A(p_input[359]), .B(n4522), .Z(n4524) );
  XOR U3873 ( .A(n4525), .B(n4526), .Z(n4522) );
  AND U3874 ( .A(n493), .B(n4527), .Z(n4526) );
  IV U3875 ( .A(n4519), .Z(n4521) );
  XOR U3876 ( .A(n4528), .B(n4529), .Z(n4519) );
  AND U3877 ( .A(n497), .B(n4530), .Z(n4529) );
  XOR U3878 ( .A(n4531), .B(n4532), .Z(n4517) );
  AND U3879 ( .A(n501), .B(n4530), .Z(n4532) );
  XNOR U3880 ( .A(n4531), .B(n4528), .Z(n4530) );
  XOR U3881 ( .A(n4533), .B(n4534), .Z(n4528) );
  AND U3882 ( .A(n504), .B(n4527), .Z(n4534) );
  XNOR U3883 ( .A(n4535), .B(n4525), .Z(n4527) );
  XOR U3884 ( .A(n4536), .B(n4537), .Z(n4525) );
  AND U3885 ( .A(n508), .B(n4538), .Z(n4537) );
  XOR U3886 ( .A(p_input[375]), .B(n4536), .Z(n4538) );
  XOR U3887 ( .A(n4539), .B(n4540), .Z(n4536) );
  AND U3888 ( .A(n512), .B(n4541), .Z(n4540) );
  IV U3889 ( .A(n4533), .Z(n4535) );
  XOR U3890 ( .A(n4542), .B(n4543), .Z(n4533) );
  AND U3891 ( .A(n516), .B(n4544), .Z(n4543) );
  XOR U3892 ( .A(n4545), .B(n4546), .Z(n4531) );
  AND U3893 ( .A(n520), .B(n4544), .Z(n4546) );
  XNOR U3894 ( .A(n4545), .B(n4542), .Z(n4544) );
  XOR U3895 ( .A(n4547), .B(n4548), .Z(n4542) );
  AND U3896 ( .A(n523), .B(n4541), .Z(n4548) );
  XNOR U3897 ( .A(n4549), .B(n4539), .Z(n4541) );
  XOR U3898 ( .A(n4550), .B(n4551), .Z(n4539) );
  AND U3899 ( .A(n527), .B(n4552), .Z(n4551) );
  XOR U3900 ( .A(p_input[391]), .B(n4550), .Z(n4552) );
  XOR U3901 ( .A(n4553), .B(n4554), .Z(n4550) );
  AND U3902 ( .A(n531), .B(n4555), .Z(n4554) );
  IV U3903 ( .A(n4547), .Z(n4549) );
  XOR U3904 ( .A(n4556), .B(n4557), .Z(n4547) );
  AND U3905 ( .A(n535), .B(n4558), .Z(n4557) );
  XOR U3906 ( .A(n4559), .B(n4560), .Z(n4545) );
  AND U3907 ( .A(n539), .B(n4558), .Z(n4560) );
  XNOR U3908 ( .A(n4559), .B(n4556), .Z(n4558) );
  XOR U3909 ( .A(n4561), .B(n4562), .Z(n4556) );
  AND U3910 ( .A(n542), .B(n4555), .Z(n4562) );
  XNOR U3911 ( .A(n4563), .B(n4553), .Z(n4555) );
  XOR U3912 ( .A(n4564), .B(n4565), .Z(n4553) );
  AND U3913 ( .A(n546), .B(n4566), .Z(n4565) );
  XOR U3914 ( .A(p_input[407]), .B(n4564), .Z(n4566) );
  XOR U3915 ( .A(n4567), .B(n4568), .Z(n4564) );
  AND U3916 ( .A(n550), .B(n4569), .Z(n4568) );
  IV U3917 ( .A(n4561), .Z(n4563) );
  XOR U3918 ( .A(n4570), .B(n4571), .Z(n4561) );
  AND U3919 ( .A(n554), .B(n4572), .Z(n4571) );
  XOR U3920 ( .A(n4573), .B(n4574), .Z(n4559) );
  AND U3921 ( .A(n558), .B(n4572), .Z(n4574) );
  XNOR U3922 ( .A(n4573), .B(n4570), .Z(n4572) );
  XOR U3923 ( .A(n4575), .B(n4576), .Z(n4570) );
  AND U3924 ( .A(n561), .B(n4569), .Z(n4576) );
  XNOR U3925 ( .A(n4577), .B(n4567), .Z(n4569) );
  XOR U3926 ( .A(n4578), .B(n4579), .Z(n4567) );
  AND U3927 ( .A(n565), .B(n4580), .Z(n4579) );
  XOR U3928 ( .A(p_input[423]), .B(n4578), .Z(n4580) );
  XOR U3929 ( .A(n4581), .B(n4582), .Z(n4578) );
  AND U3930 ( .A(n569), .B(n4583), .Z(n4582) );
  IV U3931 ( .A(n4575), .Z(n4577) );
  XOR U3932 ( .A(n4584), .B(n4585), .Z(n4575) );
  AND U3933 ( .A(n573), .B(n4586), .Z(n4585) );
  XOR U3934 ( .A(n4587), .B(n4588), .Z(n4573) );
  AND U3935 ( .A(n577), .B(n4586), .Z(n4588) );
  XNOR U3936 ( .A(n4587), .B(n4584), .Z(n4586) );
  XOR U3937 ( .A(n4589), .B(n4590), .Z(n4584) );
  AND U3938 ( .A(n580), .B(n4583), .Z(n4590) );
  XNOR U3939 ( .A(n4591), .B(n4581), .Z(n4583) );
  XOR U3940 ( .A(n4592), .B(n4593), .Z(n4581) );
  AND U3941 ( .A(n584), .B(n4594), .Z(n4593) );
  XOR U3942 ( .A(p_input[439]), .B(n4592), .Z(n4594) );
  XOR U3943 ( .A(n4595), .B(n4596), .Z(n4592) );
  AND U3944 ( .A(n588), .B(n4597), .Z(n4596) );
  IV U3945 ( .A(n4589), .Z(n4591) );
  XOR U3946 ( .A(n4598), .B(n4599), .Z(n4589) );
  AND U3947 ( .A(n592), .B(n4600), .Z(n4599) );
  XOR U3948 ( .A(n4601), .B(n4602), .Z(n4587) );
  AND U3949 ( .A(n596), .B(n4600), .Z(n4602) );
  XNOR U3950 ( .A(n4601), .B(n4598), .Z(n4600) );
  XOR U3951 ( .A(n4603), .B(n4604), .Z(n4598) );
  AND U3952 ( .A(n599), .B(n4597), .Z(n4604) );
  XNOR U3953 ( .A(n4605), .B(n4595), .Z(n4597) );
  XOR U3954 ( .A(n4606), .B(n4607), .Z(n4595) );
  AND U3955 ( .A(n603), .B(n4608), .Z(n4607) );
  XOR U3956 ( .A(p_input[455]), .B(n4606), .Z(n4608) );
  XOR U3957 ( .A(n4609), .B(n4610), .Z(n4606) );
  AND U3958 ( .A(n607), .B(n4611), .Z(n4610) );
  IV U3959 ( .A(n4603), .Z(n4605) );
  XOR U3960 ( .A(n4612), .B(n4613), .Z(n4603) );
  AND U3961 ( .A(n611), .B(n4614), .Z(n4613) );
  XOR U3962 ( .A(n4615), .B(n4616), .Z(n4601) );
  AND U3963 ( .A(n615), .B(n4614), .Z(n4616) );
  XNOR U3964 ( .A(n4615), .B(n4612), .Z(n4614) );
  XOR U3965 ( .A(n4617), .B(n4618), .Z(n4612) );
  AND U3966 ( .A(n618), .B(n4611), .Z(n4618) );
  XNOR U3967 ( .A(n4619), .B(n4609), .Z(n4611) );
  XOR U3968 ( .A(n4620), .B(n4621), .Z(n4609) );
  AND U3969 ( .A(n622), .B(n4622), .Z(n4621) );
  XOR U3970 ( .A(p_input[471]), .B(n4620), .Z(n4622) );
  XOR U3971 ( .A(n4623), .B(n4624), .Z(n4620) );
  AND U3972 ( .A(n626), .B(n4625), .Z(n4624) );
  IV U3973 ( .A(n4617), .Z(n4619) );
  XOR U3974 ( .A(n4626), .B(n4627), .Z(n4617) );
  AND U3975 ( .A(n630), .B(n4628), .Z(n4627) );
  XOR U3976 ( .A(n4629), .B(n4630), .Z(n4615) );
  AND U3977 ( .A(n634), .B(n4628), .Z(n4630) );
  XNOR U3978 ( .A(n4629), .B(n4626), .Z(n4628) );
  XOR U3979 ( .A(n4631), .B(n4632), .Z(n4626) );
  AND U3980 ( .A(n637), .B(n4625), .Z(n4632) );
  XNOR U3981 ( .A(n4633), .B(n4623), .Z(n4625) );
  XOR U3982 ( .A(n4634), .B(n4635), .Z(n4623) );
  AND U3983 ( .A(n641), .B(n4636), .Z(n4635) );
  XOR U3984 ( .A(p_input[487]), .B(n4634), .Z(n4636) );
  XOR U3985 ( .A(n4637), .B(n4638), .Z(n4634) );
  AND U3986 ( .A(n645), .B(n4639), .Z(n4638) );
  IV U3987 ( .A(n4631), .Z(n4633) );
  XOR U3988 ( .A(n4640), .B(n4641), .Z(n4631) );
  AND U3989 ( .A(n649), .B(n4642), .Z(n4641) );
  XOR U3990 ( .A(n4643), .B(n4644), .Z(n4629) );
  AND U3991 ( .A(n653), .B(n4642), .Z(n4644) );
  XNOR U3992 ( .A(n4643), .B(n4640), .Z(n4642) );
  XOR U3993 ( .A(n4645), .B(n4646), .Z(n4640) );
  AND U3994 ( .A(n656), .B(n4639), .Z(n4646) );
  XNOR U3995 ( .A(n4647), .B(n4637), .Z(n4639) );
  XOR U3996 ( .A(n4648), .B(n4649), .Z(n4637) );
  AND U3997 ( .A(n660), .B(n4650), .Z(n4649) );
  XOR U3998 ( .A(p_input[503]), .B(n4648), .Z(n4650) );
  XOR U3999 ( .A(n4651), .B(n4652), .Z(n4648) );
  AND U4000 ( .A(n664), .B(n4653), .Z(n4652) );
  IV U4001 ( .A(n4645), .Z(n4647) );
  XOR U4002 ( .A(n4654), .B(n4655), .Z(n4645) );
  AND U4003 ( .A(n668), .B(n4656), .Z(n4655) );
  XOR U4004 ( .A(n4657), .B(n4658), .Z(n4643) );
  AND U4005 ( .A(n672), .B(n4656), .Z(n4658) );
  XNOR U4006 ( .A(n4657), .B(n4654), .Z(n4656) );
  XOR U4007 ( .A(n4659), .B(n4660), .Z(n4654) );
  AND U4008 ( .A(n675), .B(n4653), .Z(n4660) );
  XNOR U4009 ( .A(n4661), .B(n4651), .Z(n4653) );
  XOR U4010 ( .A(n4662), .B(n4663), .Z(n4651) );
  AND U4011 ( .A(n679), .B(n4664), .Z(n4663) );
  XOR U4012 ( .A(p_input[519]), .B(n4662), .Z(n4664) );
  XOR U4013 ( .A(n4665), .B(n4666), .Z(n4662) );
  AND U4014 ( .A(n683), .B(n4667), .Z(n4666) );
  IV U4015 ( .A(n4659), .Z(n4661) );
  XOR U4016 ( .A(n4668), .B(n4669), .Z(n4659) );
  AND U4017 ( .A(n687), .B(n4670), .Z(n4669) );
  XOR U4018 ( .A(n4671), .B(n4672), .Z(n4657) );
  AND U4019 ( .A(n691), .B(n4670), .Z(n4672) );
  XNOR U4020 ( .A(n4671), .B(n4668), .Z(n4670) );
  XOR U4021 ( .A(n4673), .B(n4674), .Z(n4668) );
  AND U4022 ( .A(n694), .B(n4667), .Z(n4674) );
  XNOR U4023 ( .A(n4675), .B(n4665), .Z(n4667) );
  XOR U4024 ( .A(n4676), .B(n4677), .Z(n4665) );
  AND U4025 ( .A(n698), .B(n4678), .Z(n4677) );
  XOR U4026 ( .A(p_input[535]), .B(n4676), .Z(n4678) );
  XOR U4027 ( .A(n4679), .B(n4680), .Z(n4676) );
  AND U4028 ( .A(n702), .B(n4681), .Z(n4680) );
  IV U4029 ( .A(n4673), .Z(n4675) );
  XOR U4030 ( .A(n4682), .B(n4683), .Z(n4673) );
  AND U4031 ( .A(n706), .B(n4684), .Z(n4683) );
  XOR U4032 ( .A(n4685), .B(n4686), .Z(n4671) );
  AND U4033 ( .A(n710), .B(n4684), .Z(n4686) );
  XNOR U4034 ( .A(n4685), .B(n4682), .Z(n4684) );
  XOR U4035 ( .A(n4687), .B(n4688), .Z(n4682) );
  AND U4036 ( .A(n713), .B(n4681), .Z(n4688) );
  XNOR U4037 ( .A(n4689), .B(n4679), .Z(n4681) );
  XOR U4038 ( .A(n4690), .B(n4691), .Z(n4679) );
  AND U4039 ( .A(n717), .B(n4692), .Z(n4691) );
  XOR U4040 ( .A(p_input[551]), .B(n4690), .Z(n4692) );
  XOR U4041 ( .A(n4693), .B(n4694), .Z(n4690) );
  AND U4042 ( .A(n721), .B(n4695), .Z(n4694) );
  IV U4043 ( .A(n4687), .Z(n4689) );
  XOR U4044 ( .A(n4696), .B(n4697), .Z(n4687) );
  AND U4045 ( .A(n725), .B(n4698), .Z(n4697) );
  XOR U4046 ( .A(n4699), .B(n4700), .Z(n4685) );
  AND U4047 ( .A(n729), .B(n4698), .Z(n4700) );
  XNOR U4048 ( .A(n4699), .B(n4696), .Z(n4698) );
  XOR U4049 ( .A(n4701), .B(n4702), .Z(n4696) );
  AND U4050 ( .A(n732), .B(n4695), .Z(n4702) );
  XNOR U4051 ( .A(n4703), .B(n4693), .Z(n4695) );
  XOR U4052 ( .A(n4704), .B(n4705), .Z(n4693) );
  AND U4053 ( .A(n736), .B(n4706), .Z(n4705) );
  XOR U4054 ( .A(p_input[567]), .B(n4704), .Z(n4706) );
  XOR U4055 ( .A(n4707), .B(n4708), .Z(n4704) );
  AND U4056 ( .A(n740), .B(n4709), .Z(n4708) );
  IV U4057 ( .A(n4701), .Z(n4703) );
  XOR U4058 ( .A(n4710), .B(n4711), .Z(n4701) );
  AND U4059 ( .A(n744), .B(n4712), .Z(n4711) );
  XOR U4060 ( .A(n4713), .B(n4714), .Z(n4699) );
  AND U4061 ( .A(n748), .B(n4712), .Z(n4714) );
  XNOR U4062 ( .A(n4713), .B(n4710), .Z(n4712) );
  XOR U4063 ( .A(n4715), .B(n4716), .Z(n4710) );
  AND U4064 ( .A(n751), .B(n4709), .Z(n4716) );
  XNOR U4065 ( .A(n4717), .B(n4707), .Z(n4709) );
  XOR U4066 ( .A(n4718), .B(n4719), .Z(n4707) );
  AND U4067 ( .A(n755), .B(n4720), .Z(n4719) );
  XOR U4068 ( .A(p_input[583]), .B(n4718), .Z(n4720) );
  XOR U4069 ( .A(n4721), .B(n4722), .Z(n4718) );
  AND U4070 ( .A(n759), .B(n4723), .Z(n4722) );
  IV U4071 ( .A(n4715), .Z(n4717) );
  XOR U4072 ( .A(n4724), .B(n4725), .Z(n4715) );
  AND U4073 ( .A(n763), .B(n4726), .Z(n4725) );
  XOR U4074 ( .A(n4727), .B(n4728), .Z(n4713) );
  AND U4075 ( .A(n767), .B(n4726), .Z(n4728) );
  XNOR U4076 ( .A(n4727), .B(n4724), .Z(n4726) );
  XOR U4077 ( .A(n4729), .B(n4730), .Z(n4724) );
  AND U4078 ( .A(n770), .B(n4723), .Z(n4730) );
  XNOR U4079 ( .A(n4731), .B(n4721), .Z(n4723) );
  XOR U4080 ( .A(n4732), .B(n4733), .Z(n4721) );
  AND U4081 ( .A(n774), .B(n4734), .Z(n4733) );
  XOR U4082 ( .A(p_input[599]), .B(n4732), .Z(n4734) );
  XOR U4083 ( .A(n4735), .B(n4736), .Z(n4732) );
  AND U4084 ( .A(n778), .B(n4737), .Z(n4736) );
  IV U4085 ( .A(n4729), .Z(n4731) );
  XOR U4086 ( .A(n4738), .B(n4739), .Z(n4729) );
  AND U4087 ( .A(n782), .B(n4740), .Z(n4739) );
  XOR U4088 ( .A(n4741), .B(n4742), .Z(n4727) );
  AND U4089 ( .A(n786), .B(n4740), .Z(n4742) );
  XNOR U4090 ( .A(n4741), .B(n4738), .Z(n4740) );
  XOR U4091 ( .A(n4743), .B(n4744), .Z(n4738) );
  AND U4092 ( .A(n789), .B(n4737), .Z(n4744) );
  XNOR U4093 ( .A(n4745), .B(n4735), .Z(n4737) );
  XOR U4094 ( .A(n4746), .B(n4747), .Z(n4735) );
  AND U4095 ( .A(n793), .B(n4748), .Z(n4747) );
  XOR U4096 ( .A(p_input[615]), .B(n4746), .Z(n4748) );
  XOR U4097 ( .A(n4749), .B(n4750), .Z(n4746) );
  AND U4098 ( .A(n797), .B(n4751), .Z(n4750) );
  IV U4099 ( .A(n4743), .Z(n4745) );
  XOR U4100 ( .A(n4752), .B(n4753), .Z(n4743) );
  AND U4101 ( .A(n801), .B(n4754), .Z(n4753) );
  XOR U4102 ( .A(n4755), .B(n4756), .Z(n4741) );
  AND U4103 ( .A(n805), .B(n4754), .Z(n4756) );
  XNOR U4104 ( .A(n4755), .B(n4752), .Z(n4754) );
  XOR U4105 ( .A(n4757), .B(n4758), .Z(n4752) );
  AND U4106 ( .A(n808), .B(n4751), .Z(n4758) );
  XNOR U4107 ( .A(n4759), .B(n4749), .Z(n4751) );
  XOR U4108 ( .A(n4760), .B(n4761), .Z(n4749) );
  AND U4109 ( .A(n812), .B(n4762), .Z(n4761) );
  XOR U4110 ( .A(p_input[631]), .B(n4760), .Z(n4762) );
  XOR U4111 ( .A(n4763), .B(n4764), .Z(n4760) );
  AND U4112 ( .A(n816), .B(n4765), .Z(n4764) );
  IV U4113 ( .A(n4757), .Z(n4759) );
  XOR U4114 ( .A(n4766), .B(n4767), .Z(n4757) );
  AND U4115 ( .A(n820), .B(n4768), .Z(n4767) );
  XOR U4116 ( .A(n4769), .B(n4770), .Z(n4755) );
  AND U4117 ( .A(n824), .B(n4768), .Z(n4770) );
  XNOR U4118 ( .A(n4769), .B(n4766), .Z(n4768) );
  XOR U4119 ( .A(n4771), .B(n4772), .Z(n4766) );
  AND U4120 ( .A(n827), .B(n4765), .Z(n4772) );
  XNOR U4121 ( .A(n4773), .B(n4763), .Z(n4765) );
  XOR U4122 ( .A(n4774), .B(n4775), .Z(n4763) );
  AND U4123 ( .A(n831), .B(n4776), .Z(n4775) );
  XOR U4124 ( .A(p_input[647]), .B(n4774), .Z(n4776) );
  XOR U4125 ( .A(n4777), .B(n4778), .Z(n4774) );
  AND U4126 ( .A(n835), .B(n4779), .Z(n4778) );
  IV U4127 ( .A(n4771), .Z(n4773) );
  XOR U4128 ( .A(n4780), .B(n4781), .Z(n4771) );
  AND U4129 ( .A(n839), .B(n4782), .Z(n4781) );
  XOR U4130 ( .A(n4783), .B(n4784), .Z(n4769) );
  AND U4131 ( .A(n843), .B(n4782), .Z(n4784) );
  XNOR U4132 ( .A(n4783), .B(n4780), .Z(n4782) );
  XOR U4133 ( .A(n4785), .B(n4786), .Z(n4780) );
  AND U4134 ( .A(n846), .B(n4779), .Z(n4786) );
  XNOR U4135 ( .A(n4787), .B(n4777), .Z(n4779) );
  XOR U4136 ( .A(n4788), .B(n4789), .Z(n4777) );
  AND U4137 ( .A(n850), .B(n4790), .Z(n4789) );
  XOR U4138 ( .A(p_input[663]), .B(n4788), .Z(n4790) );
  XOR U4139 ( .A(n4791), .B(n4792), .Z(n4788) );
  AND U4140 ( .A(n854), .B(n4793), .Z(n4792) );
  IV U4141 ( .A(n4785), .Z(n4787) );
  XOR U4142 ( .A(n4794), .B(n4795), .Z(n4785) );
  AND U4143 ( .A(n858), .B(n4796), .Z(n4795) );
  XOR U4144 ( .A(n4797), .B(n4798), .Z(n4783) );
  AND U4145 ( .A(n862), .B(n4796), .Z(n4798) );
  XNOR U4146 ( .A(n4797), .B(n4794), .Z(n4796) );
  XOR U4147 ( .A(n4799), .B(n4800), .Z(n4794) );
  AND U4148 ( .A(n865), .B(n4793), .Z(n4800) );
  XNOR U4149 ( .A(n4801), .B(n4791), .Z(n4793) );
  XOR U4150 ( .A(n4802), .B(n4803), .Z(n4791) );
  AND U4151 ( .A(n869), .B(n4804), .Z(n4803) );
  XOR U4152 ( .A(p_input[679]), .B(n4802), .Z(n4804) );
  XOR U4153 ( .A(n4805), .B(n4806), .Z(n4802) );
  AND U4154 ( .A(n873), .B(n4807), .Z(n4806) );
  IV U4155 ( .A(n4799), .Z(n4801) );
  XOR U4156 ( .A(n4808), .B(n4809), .Z(n4799) );
  AND U4157 ( .A(n877), .B(n4810), .Z(n4809) );
  XOR U4158 ( .A(n4811), .B(n4812), .Z(n4797) );
  AND U4159 ( .A(n881), .B(n4810), .Z(n4812) );
  XNOR U4160 ( .A(n4811), .B(n4808), .Z(n4810) );
  XOR U4161 ( .A(n4813), .B(n4814), .Z(n4808) );
  AND U4162 ( .A(n884), .B(n4807), .Z(n4814) );
  XNOR U4163 ( .A(n4815), .B(n4805), .Z(n4807) );
  XOR U4164 ( .A(n4816), .B(n4817), .Z(n4805) );
  AND U4165 ( .A(n888), .B(n4818), .Z(n4817) );
  XOR U4166 ( .A(p_input[695]), .B(n4816), .Z(n4818) );
  XOR U4167 ( .A(n4819), .B(n4820), .Z(n4816) );
  AND U4168 ( .A(n892), .B(n4821), .Z(n4820) );
  IV U4169 ( .A(n4813), .Z(n4815) );
  XOR U4170 ( .A(n4822), .B(n4823), .Z(n4813) );
  AND U4171 ( .A(n896), .B(n4824), .Z(n4823) );
  XOR U4172 ( .A(n4825), .B(n4826), .Z(n4811) );
  AND U4173 ( .A(n900), .B(n4824), .Z(n4826) );
  XNOR U4174 ( .A(n4825), .B(n4822), .Z(n4824) );
  XOR U4175 ( .A(n4827), .B(n4828), .Z(n4822) );
  AND U4176 ( .A(n903), .B(n4821), .Z(n4828) );
  XNOR U4177 ( .A(n4829), .B(n4819), .Z(n4821) );
  XOR U4178 ( .A(n4830), .B(n4831), .Z(n4819) );
  AND U4179 ( .A(n907), .B(n4832), .Z(n4831) );
  XOR U4180 ( .A(p_input[711]), .B(n4830), .Z(n4832) );
  XOR U4181 ( .A(n4833), .B(n4834), .Z(n4830) );
  AND U4182 ( .A(n911), .B(n4835), .Z(n4834) );
  IV U4183 ( .A(n4827), .Z(n4829) );
  XOR U4184 ( .A(n4836), .B(n4837), .Z(n4827) );
  AND U4185 ( .A(n915), .B(n4838), .Z(n4837) );
  XOR U4186 ( .A(n4839), .B(n4840), .Z(n4825) );
  AND U4187 ( .A(n919), .B(n4838), .Z(n4840) );
  XNOR U4188 ( .A(n4839), .B(n4836), .Z(n4838) );
  XOR U4189 ( .A(n4841), .B(n4842), .Z(n4836) );
  AND U4190 ( .A(n922), .B(n4835), .Z(n4842) );
  XNOR U4191 ( .A(n4843), .B(n4833), .Z(n4835) );
  XOR U4192 ( .A(n4844), .B(n4845), .Z(n4833) );
  AND U4193 ( .A(n926), .B(n4846), .Z(n4845) );
  XOR U4194 ( .A(p_input[727]), .B(n4844), .Z(n4846) );
  XOR U4195 ( .A(n4847), .B(n4848), .Z(n4844) );
  AND U4196 ( .A(n930), .B(n4849), .Z(n4848) );
  IV U4197 ( .A(n4841), .Z(n4843) );
  XOR U4198 ( .A(n4850), .B(n4851), .Z(n4841) );
  AND U4199 ( .A(n934), .B(n4852), .Z(n4851) );
  XOR U4200 ( .A(n4853), .B(n4854), .Z(n4839) );
  AND U4201 ( .A(n938), .B(n4852), .Z(n4854) );
  XNOR U4202 ( .A(n4853), .B(n4850), .Z(n4852) );
  XOR U4203 ( .A(n4855), .B(n4856), .Z(n4850) );
  AND U4204 ( .A(n941), .B(n4849), .Z(n4856) );
  XNOR U4205 ( .A(n4857), .B(n4847), .Z(n4849) );
  XOR U4206 ( .A(n4858), .B(n4859), .Z(n4847) );
  AND U4207 ( .A(n945), .B(n4860), .Z(n4859) );
  XOR U4208 ( .A(p_input[743]), .B(n4858), .Z(n4860) );
  XOR U4209 ( .A(n4861), .B(n4862), .Z(n4858) );
  AND U4210 ( .A(n949), .B(n4863), .Z(n4862) );
  IV U4211 ( .A(n4855), .Z(n4857) );
  XOR U4212 ( .A(n4864), .B(n4865), .Z(n4855) );
  AND U4213 ( .A(n953), .B(n4866), .Z(n4865) );
  XOR U4214 ( .A(n4867), .B(n4868), .Z(n4853) );
  AND U4215 ( .A(n957), .B(n4866), .Z(n4868) );
  XNOR U4216 ( .A(n4867), .B(n4864), .Z(n4866) );
  XOR U4217 ( .A(n4869), .B(n4870), .Z(n4864) );
  AND U4218 ( .A(n960), .B(n4863), .Z(n4870) );
  XNOR U4219 ( .A(n4871), .B(n4861), .Z(n4863) );
  XOR U4220 ( .A(n4872), .B(n4873), .Z(n4861) );
  AND U4221 ( .A(n964), .B(n4874), .Z(n4873) );
  XOR U4222 ( .A(p_input[759]), .B(n4872), .Z(n4874) );
  XOR U4223 ( .A(n4875), .B(n4876), .Z(n4872) );
  AND U4224 ( .A(n968), .B(n4877), .Z(n4876) );
  IV U4225 ( .A(n4869), .Z(n4871) );
  XOR U4226 ( .A(n4878), .B(n4879), .Z(n4869) );
  AND U4227 ( .A(n972), .B(n4880), .Z(n4879) );
  XOR U4228 ( .A(n4881), .B(n4882), .Z(n4867) );
  AND U4229 ( .A(n976), .B(n4880), .Z(n4882) );
  XNOR U4230 ( .A(n4881), .B(n4878), .Z(n4880) );
  XOR U4231 ( .A(n4883), .B(n4884), .Z(n4878) );
  AND U4232 ( .A(n979), .B(n4877), .Z(n4884) );
  XNOR U4233 ( .A(n4885), .B(n4875), .Z(n4877) );
  XOR U4234 ( .A(n4886), .B(n4887), .Z(n4875) );
  AND U4235 ( .A(n983), .B(n4888), .Z(n4887) );
  XOR U4236 ( .A(p_input[775]), .B(n4886), .Z(n4888) );
  XOR U4237 ( .A(n4889), .B(n4890), .Z(n4886) );
  AND U4238 ( .A(n987), .B(n4891), .Z(n4890) );
  IV U4239 ( .A(n4883), .Z(n4885) );
  XOR U4240 ( .A(n4892), .B(n4893), .Z(n4883) );
  AND U4241 ( .A(n991), .B(n4894), .Z(n4893) );
  XOR U4242 ( .A(n4895), .B(n4896), .Z(n4881) );
  AND U4243 ( .A(n995), .B(n4894), .Z(n4896) );
  XNOR U4244 ( .A(n4895), .B(n4892), .Z(n4894) );
  XOR U4245 ( .A(n4897), .B(n4898), .Z(n4892) );
  AND U4246 ( .A(n998), .B(n4891), .Z(n4898) );
  XNOR U4247 ( .A(n4899), .B(n4889), .Z(n4891) );
  XOR U4248 ( .A(n4900), .B(n4901), .Z(n4889) );
  AND U4249 ( .A(n1002), .B(n4902), .Z(n4901) );
  XOR U4250 ( .A(p_input[791]), .B(n4900), .Z(n4902) );
  XOR U4251 ( .A(n4903), .B(n4904), .Z(n4900) );
  AND U4252 ( .A(n1006), .B(n4905), .Z(n4904) );
  IV U4253 ( .A(n4897), .Z(n4899) );
  XOR U4254 ( .A(n4906), .B(n4907), .Z(n4897) );
  AND U4255 ( .A(n1010), .B(n4908), .Z(n4907) );
  XOR U4256 ( .A(n4909), .B(n4910), .Z(n4895) );
  AND U4257 ( .A(n1014), .B(n4908), .Z(n4910) );
  XNOR U4258 ( .A(n4909), .B(n4906), .Z(n4908) );
  XOR U4259 ( .A(n4911), .B(n4912), .Z(n4906) );
  AND U4260 ( .A(n1017), .B(n4905), .Z(n4912) );
  XNOR U4261 ( .A(n4913), .B(n4903), .Z(n4905) );
  XOR U4262 ( .A(n4914), .B(n4915), .Z(n4903) );
  AND U4263 ( .A(n1021), .B(n4916), .Z(n4915) );
  XOR U4264 ( .A(p_input[807]), .B(n4914), .Z(n4916) );
  XOR U4265 ( .A(n4917), .B(n4918), .Z(n4914) );
  AND U4266 ( .A(n1025), .B(n4919), .Z(n4918) );
  IV U4267 ( .A(n4911), .Z(n4913) );
  XOR U4268 ( .A(n4920), .B(n4921), .Z(n4911) );
  AND U4269 ( .A(n1029), .B(n4922), .Z(n4921) );
  XOR U4270 ( .A(n4923), .B(n4924), .Z(n4909) );
  AND U4271 ( .A(n1033), .B(n4922), .Z(n4924) );
  XNOR U4272 ( .A(n4923), .B(n4920), .Z(n4922) );
  XOR U4273 ( .A(n4925), .B(n4926), .Z(n4920) );
  AND U4274 ( .A(n1036), .B(n4919), .Z(n4926) );
  XNOR U4275 ( .A(n4927), .B(n4917), .Z(n4919) );
  XOR U4276 ( .A(n4928), .B(n4929), .Z(n4917) );
  AND U4277 ( .A(n1040), .B(n4930), .Z(n4929) );
  XOR U4278 ( .A(p_input[823]), .B(n4928), .Z(n4930) );
  XOR U4279 ( .A(n4931), .B(n4932), .Z(n4928) );
  AND U4280 ( .A(n1044), .B(n4933), .Z(n4932) );
  IV U4281 ( .A(n4925), .Z(n4927) );
  XOR U4282 ( .A(n4934), .B(n4935), .Z(n4925) );
  AND U4283 ( .A(n1048), .B(n4936), .Z(n4935) );
  XOR U4284 ( .A(n4937), .B(n4938), .Z(n4923) );
  AND U4285 ( .A(n1052), .B(n4936), .Z(n4938) );
  XNOR U4286 ( .A(n4937), .B(n4934), .Z(n4936) );
  XOR U4287 ( .A(n4939), .B(n4940), .Z(n4934) );
  AND U4288 ( .A(n1055), .B(n4933), .Z(n4940) );
  XNOR U4289 ( .A(n4941), .B(n4931), .Z(n4933) );
  XOR U4290 ( .A(n4942), .B(n4943), .Z(n4931) );
  AND U4291 ( .A(n1059), .B(n4944), .Z(n4943) );
  XOR U4292 ( .A(p_input[839]), .B(n4942), .Z(n4944) );
  XOR U4293 ( .A(n4945), .B(n4946), .Z(n4942) );
  AND U4294 ( .A(n1063), .B(n4947), .Z(n4946) );
  IV U4295 ( .A(n4939), .Z(n4941) );
  XOR U4296 ( .A(n4948), .B(n4949), .Z(n4939) );
  AND U4297 ( .A(n1067), .B(n4950), .Z(n4949) );
  XOR U4298 ( .A(n4951), .B(n4952), .Z(n4937) );
  AND U4299 ( .A(n1071), .B(n4950), .Z(n4952) );
  XNOR U4300 ( .A(n4951), .B(n4948), .Z(n4950) );
  XOR U4301 ( .A(n4953), .B(n4954), .Z(n4948) );
  AND U4302 ( .A(n1074), .B(n4947), .Z(n4954) );
  XNOR U4303 ( .A(n4955), .B(n4945), .Z(n4947) );
  XOR U4304 ( .A(n4956), .B(n4957), .Z(n4945) );
  AND U4305 ( .A(n1078), .B(n4958), .Z(n4957) );
  XOR U4306 ( .A(p_input[855]), .B(n4956), .Z(n4958) );
  XOR U4307 ( .A(n4959), .B(n4960), .Z(n4956) );
  AND U4308 ( .A(n1082), .B(n4961), .Z(n4960) );
  IV U4309 ( .A(n4953), .Z(n4955) );
  XOR U4310 ( .A(n4962), .B(n4963), .Z(n4953) );
  AND U4311 ( .A(n1086), .B(n4964), .Z(n4963) );
  XOR U4312 ( .A(n4965), .B(n4966), .Z(n4951) );
  AND U4313 ( .A(n1090), .B(n4964), .Z(n4966) );
  XNOR U4314 ( .A(n4965), .B(n4962), .Z(n4964) );
  XOR U4315 ( .A(n4967), .B(n4968), .Z(n4962) );
  AND U4316 ( .A(n1093), .B(n4961), .Z(n4968) );
  XNOR U4317 ( .A(n4969), .B(n4959), .Z(n4961) );
  XOR U4318 ( .A(n4970), .B(n4971), .Z(n4959) );
  AND U4319 ( .A(n1097), .B(n4972), .Z(n4971) );
  XOR U4320 ( .A(p_input[871]), .B(n4970), .Z(n4972) );
  XOR U4321 ( .A(n4973), .B(n4974), .Z(n4970) );
  AND U4322 ( .A(n1101), .B(n4975), .Z(n4974) );
  IV U4323 ( .A(n4967), .Z(n4969) );
  XOR U4324 ( .A(n4976), .B(n4977), .Z(n4967) );
  AND U4325 ( .A(n1105), .B(n4978), .Z(n4977) );
  XOR U4326 ( .A(n4979), .B(n4980), .Z(n4965) );
  AND U4327 ( .A(n1109), .B(n4978), .Z(n4980) );
  XNOR U4328 ( .A(n4979), .B(n4976), .Z(n4978) );
  XOR U4329 ( .A(n4981), .B(n4982), .Z(n4976) );
  AND U4330 ( .A(n1112), .B(n4975), .Z(n4982) );
  XNOR U4331 ( .A(n4983), .B(n4973), .Z(n4975) );
  XOR U4332 ( .A(n4984), .B(n4985), .Z(n4973) );
  AND U4333 ( .A(n1116), .B(n4986), .Z(n4985) );
  XOR U4334 ( .A(p_input[887]), .B(n4984), .Z(n4986) );
  XOR U4335 ( .A(n4987), .B(n4988), .Z(n4984) );
  AND U4336 ( .A(n1120), .B(n4989), .Z(n4988) );
  IV U4337 ( .A(n4981), .Z(n4983) );
  XOR U4338 ( .A(n4990), .B(n4991), .Z(n4981) );
  AND U4339 ( .A(n1124), .B(n4992), .Z(n4991) );
  XOR U4340 ( .A(n4993), .B(n4994), .Z(n4979) );
  AND U4341 ( .A(n1128), .B(n4992), .Z(n4994) );
  XNOR U4342 ( .A(n4993), .B(n4990), .Z(n4992) );
  XOR U4343 ( .A(n4995), .B(n4996), .Z(n4990) );
  AND U4344 ( .A(n1131), .B(n4989), .Z(n4996) );
  XNOR U4345 ( .A(n4997), .B(n4987), .Z(n4989) );
  XOR U4346 ( .A(n4998), .B(n4999), .Z(n4987) );
  AND U4347 ( .A(n1135), .B(n5000), .Z(n4999) );
  XOR U4348 ( .A(p_input[903]), .B(n4998), .Z(n5000) );
  XOR U4349 ( .A(n5001), .B(n5002), .Z(n4998) );
  AND U4350 ( .A(n1139), .B(n5003), .Z(n5002) );
  IV U4351 ( .A(n4995), .Z(n4997) );
  XOR U4352 ( .A(n5004), .B(n5005), .Z(n4995) );
  AND U4353 ( .A(n1143), .B(n5006), .Z(n5005) );
  XOR U4354 ( .A(n5007), .B(n5008), .Z(n4993) );
  AND U4355 ( .A(n1147), .B(n5006), .Z(n5008) );
  XNOR U4356 ( .A(n5007), .B(n5004), .Z(n5006) );
  XOR U4357 ( .A(n5009), .B(n5010), .Z(n5004) );
  AND U4358 ( .A(n1150), .B(n5003), .Z(n5010) );
  XNOR U4359 ( .A(n5011), .B(n5001), .Z(n5003) );
  XOR U4360 ( .A(n5012), .B(n5013), .Z(n5001) );
  AND U4361 ( .A(n1154), .B(n5014), .Z(n5013) );
  XOR U4362 ( .A(p_input[919]), .B(n5012), .Z(n5014) );
  XOR U4363 ( .A(n5015), .B(n5016), .Z(n5012) );
  AND U4364 ( .A(n1158), .B(n5017), .Z(n5016) );
  IV U4365 ( .A(n5009), .Z(n5011) );
  XOR U4366 ( .A(n5018), .B(n5019), .Z(n5009) );
  AND U4367 ( .A(n1162), .B(n5020), .Z(n5019) );
  XOR U4368 ( .A(n5021), .B(n5022), .Z(n5007) );
  AND U4369 ( .A(n1166), .B(n5020), .Z(n5022) );
  XNOR U4370 ( .A(n5021), .B(n5018), .Z(n5020) );
  XOR U4371 ( .A(n5023), .B(n5024), .Z(n5018) );
  AND U4372 ( .A(n1169), .B(n5017), .Z(n5024) );
  XNOR U4373 ( .A(n5025), .B(n5015), .Z(n5017) );
  XOR U4374 ( .A(n5026), .B(n5027), .Z(n5015) );
  AND U4375 ( .A(n1173), .B(n5028), .Z(n5027) );
  XOR U4376 ( .A(p_input[935]), .B(n5026), .Z(n5028) );
  XOR U4377 ( .A(n5029), .B(n5030), .Z(n5026) );
  AND U4378 ( .A(n1177), .B(n5031), .Z(n5030) );
  IV U4379 ( .A(n5023), .Z(n5025) );
  XOR U4380 ( .A(n5032), .B(n5033), .Z(n5023) );
  AND U4381 ( .A(n1181), .B(n5034), .Z(n5033) );
  XOR U4382 ( .A(n5035), .B(n5036), .Z(n5021) );
  AND U4383 ( .A(n1185), .B(n5034), .Z(n5036) );
  XNOR U4384 ( .A(n5035), .B(n5032), .Z(n5034) );
  XOR U4385 ( .A(n5037), .B(n5038), .Z(n5032) );
  AND U4386 ( .A(n1188), .B(n5031), .Z(n5038) );
  XNOR U4387 ( .A(n5039), .B(n5029), .Z(n5031) );
  XOR U4388 ( .A(n5040), .B(n5041), .Z(n5029) );
  AND U4389 ( .A(n1192), .B(n5042), .Z(n5041) );
  XOR U4390 ( .A(p_input[951]), .B(n5040), .Z(n5042) );
  XOR U4391 ( .A(n5043), .B(n5044), .Z(n5040) );
  AND U4392 ( .A(n1196), .B(n5045), .Z(n5044) );
  IV U4393 ( .A(n5037), .Z(n5039) );
  XOR U4394 ( .A(n5046), .B(n5047), .Z(n5037) );
  AND U4395 ( .A(n1200), .B(n5048), .Z(n5047) );
  XOR U4396 ( .A(n5049), .B(n5050), .Z(n5035) );
  AND U4397 ( .A(n1204), .B(n5048), .Z(n5050) );
  XNOR U4398 ( .A(n5049), .B(n5046), .Z(n5048) );
  XOR U4399 ( .A(n5051), .B(n5052), .Z(n5046) );
  AND U4400 ( .A(n1207), .B(n5045), .Z(n5052) );
  XNOR U4401 ( .A(n5053), .B(n5043), .Z(n5045) );
  XOR U4402 ( .A(n5054), .B(n5055), .Z(n5043) );
  AND U4403 ( .A(n1211), .B(n5056), .Z(n5055) );
  XOR U4404 ( .A(p_input[967]), .B(n5054), .Z(n5056) );
  XOR U4405 ( .A(n5057), .B(n5058), .Z(n5054) );
  AND U4406 ( .A(n1215), .B(n5059), .Z(n5058) );
  IV U4407 ( .A(n5051), .Z(n5053) );
  XOR U4408 ( .A(n5060), .B(n5061), .Z(n5051) );
  AND U4409 ( .A(n1219), .B(n5062), .Z(n5061) );
  XOR U4410 ( .A(n5063), .B(n5064), .Z(n5049) );
  AND U4411 ( .A(n1223), .B(n5062), .Z(n5064) );
  XNOR U4412 ( .A(n5063), .B(n5060), .Z(n5062) );
  XOR U4413 ( .A(n5065), .B(n5066), .Z(n5060) );
  AND U4414 ( .A(n1226), .B(n5059), .Z(n5066) );
  XNOR U4415 ( .A(n5067), .B(n5057), .Z(n5059) );
  XOR U4416 ( .A(n5068), .B(n5069), .Z(n5057) );
  AND U4417 ( .A(n1230), .B(n5070), .Z(n5069) );
  XOR U4418 ( .A(p_input[983]), .B(n5068), .Z(n5070) );
  XOR U4419 ( .A(n5071), .B(n5072), .Z(n5068) );
  AND U4420 ( .A(n1234), .B(n5073), .Z(n5072) );
  IV U4421 ( .A(n5065), .Z(n5067) );
  XOR U4422 ( .A(n5074), .B(n5075), .Z(n5065) );
  AND U4423 ( .A(n1238), .B(n5076), .Z(n5075) );
  XOR U4424 ( .A(n5077), .B(n5078), .Z(n5063) );
  AND U4425 ( .A(n1242), .B(n5076), .Z(n5078) );
  XNOR U4426 ( .A(n5077), .B(n5074), .Z(n5076) );
  XOR U4427 ( .A(n5079), .B(n5080), .Z(n5074) );
  AND U4428 ( .A(n1245), .B(n5073), .Z(n5080) );
  XNOR U4429 ( .A(n5081), .B(n5071), .Z(n5073) );
  XOR U4430 ( .A(n5082), .B(n5083), .Z(n5071) );
  AND U4431 ( .A(n1249), .B(n5084), .Z(n5083) );
  XOR U4432 ( .A(p_input[999]), .B(n5082), .Z(n5084) );
  XOR U4433 ( .A(n5085), .B(n5086), .Z(n5082) );
  AND U4434 ( .A(n1253), .B(n5087), .Z(n5086) );
  IV U4435 ( .A(n5079), .Z(n5081) );
  XOR U4436 ( .A(n5088), .B(n5089), .Z(n5079) );
  AND U4437 ( .A(n1257), .B(n5090), .Z(n5089) );
  XOR U4438 ( .A(n5091), .B(n5092), .Z(n5077) );
  AND U4439 ( .A(n1261), .B(n5090), .Z(n5092) );
  XNOR U4440 ( .A(n5091), .B(n5088), .Z(n5090) );
  XOR U4441 ( .A(n5093), .B(n5094), .Z(n5088) );
  AND U4442 ( .A(n1264), .B(n5087), .Z(n5094) );
  XNOR U4443 ( .A(n5095), .B(n5085), .Z(n5087) );
  XOR U4444 ( .A(n5096), .B(n5097), .Z(n5085) );
  AND U4445 ( .A(n1268), .B(n5098), .Z(n5097) );
  XOR U4446 ( .A(p_input[1015]), .B(n5096), .Z(n5098) );
  XOR U4447 ( .A(n5099), .B(n5100), .Z(n5096) );
  AND U4448 ( .A(n1272), .B(n5101), .Z(n5100) );
  IV U4449 ( .A(n5093), .Z(n5095) );
  XOR U4450 ( .A(n5102), .B(n5103), .Z(n5093) );
  AND U4451 ( .A(n1276), .B(n5104), .Z(n5103) );
  XOR U4452 ( .A(n5105), .B(n5106), .Z(n5091) );
  AND U4453 ( .A(n1280), .B(n5104), .Z(n5106) );
  XNOR U4454 ( .A(n5105), .B(n5102), .Z(n5104) );
  XOR U4455 ( .A(n5107), .B(n5108), .Z(n5102) );
  AND U4456 ( .A(n1283), .B(n5101), .Z(n5108) );
  XNOR U4457 ( .A(n5109), .B(n5099), .Z(n5101) );
  XOR U4458 ( .A(n5110), .B(n5111), .Z(n5099) );
  AND U4459 ( .A(n1287), .B(n5112), .Z(n5111) );
  XOR U4460 ( .A(p_input[1031]), .B(n5110), .Z(n5112) );
  XOR U4461 ( .A(n5113), .B(n5114), .Z(n5110) );
  AND U4462 ( .A(n1291), .B(n5115), .Z(n5114) );
  IV U4463 ( .A(n5107), .Z(n5109) );
  XOR U4464 ( .A(n5116), .B(n5117), .Z(n5107) );
  AND U4465 ( .A(n1295), .B(n5118), .Z(n5117) );
  XOR U4466 ( .A(n5119), .B(n5120), .Z(n5105) );
  AND U4467 ( .A(n1299), .B(n5118), .Z(n5120) );
  XNOR U4468 ( .A(n5119), .B(n5116), .Z(n5118) );
  XOR U4469 ( .A(n5121), .B(n5122), .Z(n5116) );
  AND U4470 ( .A(n1302), .B(n5115), .Z(n5122) );
  XNOR U4471 ( .A(n5123), .B(n5113), .Z(n5115) );
  XOR U4472 ( .A(n5124), .B(n5125), .Z(n5113) );
  AND U4473 ( .A(n1306), .B(n5126), .Z(n5125) );
  XOR U4474 ( .A(p_input[1047]), .B(n5124), .Z(n5126) );
  XOR U4475 ( .A(n5127), .B(n5128), .Z(n5124) );
  AND U4476 ( .A(n1310), .B(n5129), .Z(n5128) );
  IV U4477 ( .A(n5121), .Z(n5123) );
  XOR U4478 ( .A(n5130), .B(n5131), .Z(n5121) );
  AND U4479 ( .A(n1314), .B(n5132), .Z(n5131) );
  XOR U4480 ( .A(n5133), .B(n5134), .Z(n5119) );
  AND U4481 ( .A(n1318), .B(n5132), .Z(n5134) );
  XNOR U4482 ( .A(n5133), .B(n5130), .Z(n5132) );
  XOR U4483 ( .A(n5135), .B(n5136), .Z(n5130) );
  AND U4484 ( .A(n1321), .B(n5129), .Z(n5136) );
  XNOR U4485 ( .A(n5137), .B(n5127), .Z(n5129) );
  XOR U4486 ( .A(n5138), .B(n5139), .Z(n5127) );
  AND U4487 ( .A(n1325), .B(n5140), .Z(n5139) );
  XOR U4488 ( .A(p_input[1063]), .B(n5138), .Z(n5140) );
  XOR U4489 ( .A(n5141), .B(n5142), .Z(n5138) );
  AND U4490 ( .A(n1329), .B(n5143), .Z(n5142) );
  IV U4491 ( .A(n5135), .Z(n5137) );
  XOR U4492 ( .A(n5144), .B(n5145), .Z(n5135) );
  AND U4493 ( .A(n1333), .B(n5146), .Z(n5145) );
  XOR U4494 ( .A(n5147), .B(n5148), .Z(n5133) );
  AND U4495 ( .A(n1337), .B(n5146), .Z(n5148) );
  XNOR U4496 ( .A(n5147), .B(n5144), .Z(n5146) );
  XOR U4497 ( .A(n5149), .B(n5150), .Z(n5144) );
  AND U4498 ( .A(n1340), .B(n5143), .Z(n5150) );
  XNOR U4499 ( .A(n5151), .B(n5141), .Z(n5143) );
  XOR U4500 ( .A(n5152), .B(n5153), .Z(n5141) );
  AND U4501 ( .A(n1344), .B(n5154), .Z(n5153) );
  XOR U4502 ( .A(p_input[1079]), .B(n5152), .Z(n5154) );
  XOR U4503 ( .A(n5155), .B(n5156), .Z(n5152) );
  AND U4504 ( .A(n1348), .B(n5157), .Z(n5156) );
  IV U4505 ( .A(n5149), .Z(n5151) );
  XOR U4506 ( .A(n5158), .B(n5159), .Z(n5149) );
  AND U4507 ( .A(n1352), .B(n5160), .Z(n5159) );
  XOR U4508 ( .A(n5161), .B(n5162), .Z(n5147) );
  AND U4509 ( .A(n1356), .B(n5160), .Z(n5162) );
  XNOR U4510 ( .A(n5161), .B(n5158), .Z(n5160) );
  XOR U4511 ( .A(n5163), .B(n5164), .Z(n5158) );
  AND U4512 ( .A(n1359), .B(n5157), .Z(n5164) );
  XNOR U4513 ( .A(n5165), .B(n5155), .Z(n5157) );
  XOR U4514 ( .A(n5166), .B(n5167), .Z(n5155) );
  AND U4515 ( .A(n1363), .B(n5168), .Z(n5167) );
  XOR U4516 ( .A(p_input[1095]), .B(n5166), .Z(n5168) );
  XOR U4517 ( .A(n5169), .B(n5170), .Z(n5166) );
  AND U4518 ( .A(n1367), .B(n5171), .Z(n5170) );
  IV U4519 ( .A(n5163), .Z(n5165) );
  XOR U4520 ( .A(n5172), .B(n5173), .Z(n5163) );
  AND U4521 ( .A(n1371), .B(n5174), .Z(n5173) );
  XOR U4522 ( .A(n5175), .B(n5176), .Z(n5161) );
  AND U4523 ( .A(n1375), .B(n5174), .Z(n5176) );
  XNOR U4524 ( .A(n5175), .B(n5172), .Z(n5174) );
  XOR U4525 ( .A(n5177), .B(n5178), .Z(n5172) );
  AND U4526 ( .A(n1378), .B(n5171), .Z(n5178) );
  XNOR U4527 ( .A(n5179), .B(n5169), .Z(n5171) );
  XOR U4528 ( .A(n5180), .B(n5181), .Z(n5169) );
  AND U4529 ( .A(n1382), .B(n5182), .Z(n5181) );
  XOR U4530 ( .A(p_input[1111]), .B(n5180), .Z(n5182) );
  XOR U4531 ( .A(n5183), .B(n5184), .Z(n5180) );
  AND U4532 ( .A(n1386), .B(n5185), .Z(n5184) );
  IV U4533 ( .A(n5177), .Z(n5179) );
  XOR U4534 ( .A(n5186), .B(n5187), .Z(n5177) );
  AND U4535 ( .A(n1390), .B(n5188), .Z(n5187) );
  XOR U4536 ( .A(n5189), .B(n5190), .Z(n5175) );
  AND U4537 ( .A(n1394), .B(n5188), .Z(n5190) );
  XNOR U4538 ( .A(n5189), .B(n5186), .Z(n5188) );
  XOR U4539 ( .A(n5191), .B(n5192), .Z(n5186) );
  AND U4540 ( .A(n1397), .B(n5185), .Z(n5192) );
  XNOR U4541 ( .A(n5193), .B(n5183), .Z(n5185) );
  XOR U4542 ( .A(n5194), .B(n5195), .Z(n5183) );
  AND U4543 ( .A(n1401), .B(n5196), .Z(n5195) );
  XOR U4544 ( .A(p_input[1127]), .B(n5194), .Z(n5196) );
  XOR U4545 ( .A(n5197), .B(n5198), .Z(n5194) );
  AND U4546 ( .A(n1405), .B(n5199), .Z(n5198) );
  IV U4547 ( .A(n5191), .Z(n5193) );
  XOR U4548 ( .A(n5200), .B(n5201), .Z(n5191) );
  AND U4549 ( .A(n1409), .B(n5202), .Z(n5201) );
  XOR U4550 ( .A(n5203), .B(n5204), .Z(n5189) );
  AND U4551 ( .A(n1413), .B(n5202), .Z(n5204) );
  XNOR U4552 ( .A(n5203), .B(n5200), .Z(n5202) );
  XOR U4553 ( .A(n5205), .B(n5206), .Z(n5200) );
  AND U4554 ( .A(n1416), .B(n5199), .Z(n5206) );
  XNOR U4555 ( .A(n5207), .B(n5197), .Z(n5199) );
  XOR U4556 ( .A(n5208), .B(n5209), .Z(n5197) );
  AND U4557 ( .A(n1420), .B(n5210), .Z(n5209) );
  XOR U4558 ( .A(p_input[1143]), .B(n5208), .Z(n5210) );
  XOR U4559 ( .A(n5211), .B(n5212), .Z(n5208) );
  AND U4560 ( .A(n1424), .B(n5213), .Z(n5212) );
  IV U4561 ( .A(n5205), .Z(n5207) );
  XOR U4562 ( .A(n5214), .B(n5215), .Z(n5205) );
  AND U4563 ( .A(n1428), .B(n5216), .Z(n5215) );
  XOR U4564 ( .A(n5217), .B(n5218), .Z(n5203) );
  AND U4565 ( .A(n1432), .B(n5216), .Z(n5218) );
  XNOR U4566 ( .A(n5217), .B(n5214), .Z(n5216) );
  XOR U4567 ( .A(n5219), .B(n5220), .Z(n5214) );
  AND U4568 ( .A(n1435), .B(n5213), .Z(n5220) );
  XNOR U4569 ( .A(n5221), .B(n5211), .Z(n5213) );
  XOR U4570 ( .A(n5222), .B(n5223), .Z(n5211) );
  AND U4571 ( .A(n1439), .B(n5224), .Z(n5223) );
  XOR U4572 ( .A(p_input[1159]), .B(n5222), .Z(n5224) );
  XOR U4573 ( .A(n5225), .B(n5226), .Z(n5222) );
  AND U4574 ( .A(n1443), .B(n5227), .Z(n5226) );
  IV U4575 ( .A(n5219), .Z(n5221) );
  XOR U4576 ( .A(n5228), .B(n5229), .Z(n5219) );
  AND U4577 ( .A(n1447), .B(n5230), .Z(n5229) );
  XOR U4578 ( .A(n5231), .B(n5232), .Z(n5217) );
  AND U4579 ( .A(n1451), .B(n5230), .Z(n5232) );
  XNOR U4580 ( .A(n5231), .B(n5228), .Z(n5230) );
  XOR U4581 ( .A(n5233), .B(n5234), .Z(n5228) );
  AND U4582 ( .A(n1454), .B(n5227), .Z(n5234) );
  XNOR U4583 ( .A(n5235), .B(n5225), .Z(n5227) );
  XOR U4584 ( .A(n5236), .B(n5237), .Z(n5225) );
  AND U4585 ( .A(n1458), .B(n5238), .Z(n5237) );
  XOR U4586 ( .A(p_input[1175]), .B(n5236), .Z(n5238) );
  XOR U4587 ( .A(n5239), .B(n5240), .Z(n5236) );
  AND U4588 ( .A(n1462), .B(n5241), .Z(n5240) );
  IV U4589 ( .A(n5233), .Z(n5235) );
  XOR U4590 ( .A(n5242), .B(n5243), .Z(n5233) );
  AND U4591 ( .A(n1466), .B(n5244), .Z(n5243) );
  XOR U4592 ( .A(n5245), .B(n5246), .Z(n5231) );
  AND U4593 ( .A(n1470), .B(n5244), .Z(n5246) );
  XNOR U4594 ( .A(n5245), .B(n5242), .Z(n5244) );
  XOR U4595 ( .A(n5247), .B(n5248), .Z(n5242) );
  AND U4596 ( .A(n1473), .B(n5241), .Z(n5248) );
  XNOR U4597 ( .A(n5249), .B(n5239), .Z(n5241) );
  XOR U4598 ( .A(n5250), .B(n5251), .Z(n5239) );
  AND U4599 ( .A(n1477), .B(n5252), .Z(n5251) );
  XOR U4600 ( .A(p_input[1191]), .B(n5250), .Z(n5252) );
  XOR U4601 ( .A(n5253), .B(n5254), .Z(n5250) );
  AND U4602 ( .A(n1481), .B(n5255), .Z(n5254) );
  IV U4603 ( .A(n5247), .Z(n5249) );
  XOR U4604 ( .A(n5256), .B(n5257), .Z(n5247) );
  AND U4605 ( .A(n1485), .B(n5258), .Z(n5257) );
  XOR U4606 ( .A(n5259), .B(n5260), .Z(n5245) );
  AND U4607 ( .A(n1489), .B(n5258), .Z(n5260) );
  XNOR U4608 ( .A(n5259), .B(n5256), .Z(n5258) );
  XOR U4609 ( .A(n5261), .B(n5262), .Z(n5256) );
  AND U4610 ( .A(n1492), .B(n5255), .Z(n5262) );
  XNOR U4611 ( .A(n5263), .B(n5253), .Z(n5255) );
  XOR U4612 ( .A(n5264), .B(n5265), .Z(n5253) );
  AND U4613 ( .A(n1496), .B(n5266), .Z(n5265) );
  XOR U4614 ( .A(p_input[1207]), .B(n5264), .Z(n5266) );
  XOR U4615 ( .A(n5267), .B(n5268), .Z(n5264) );
  AND U4616 ( .A(n1500), .B(n5269), .Z(n5268) );
  IV U4617 ( .A(n5261), .Z(n5263) );
  XOR U4618 ( .A(n5270), .B(n5271), .Z(n5261) );
  AND U4619 ( .A(n1504), .B(n5272), .Z(n5271) );
  XOR U4620 ( .A(n5273), .B(n5274), .Z(n5259) );
  AND U4621 ( .A(n1508), .B(n5272), .Z(n5274) );
  XNOR U4622 ( .A(n5273), .B(n5270), .Z(n5272) );
  XOR U4623 ( .A(n5275), .B(n5276), .Z(n5270) );
  AND U4624 ( .A(n1511), .B(n5269), .Z(n5276) );
  XNOR U4625 ( .A(n5277), .B(n5267), .Z(n5269) );
  XOR U4626 ( .A(n5278), .B(n5279), .Z(n5267) );
  AND U4627 ( .A(n1515), .B(n5280), .Z(n5279) );
  XOR U4628 ( .A(p_input[1223]), .B(n5278), .Z(n5280) );
  XOR U4629 ( .A(n5281), .B(n5282), .Z(n5278) );
  AND U4630 ( .A(n1519), .B(n5283), .Z(n5282) );
  IV U4631 ( .A(n5275), .Z(n5277) );
  XOR U4632 ( .A(n5284), .B(n5285), .Z(n5275) );
  AND U4633 ( .A(n1523), .B(n5286), .Z(n5285) );
  XOR U4634 ( .A(n5287), .B(n5288), .Z(n5273) );
  AND U4635 ( .A(n1527), .B(n5286), .Z(n5288) );
  XNOR U4636 ( .A(n5287), .B(n5284), .Z(n5286) );
  XOR U4637 ( .A(n5289), .B(n5290), .Z(n5284) );
  AND U4638 ( .A(n1530), .B(n5283), .Z(n5290) );
  XNOR U4639 ( .A(n5291), .B(n5281), .Z(n5283) );
  XOR U4640 ( .A(n5292), .B(n5293), .Z(n5281) );
  AND U4641 ( .A(n1534), .B(n5294), .Z(n5293) );
  XOR U4642 ( .A(p_input[1239]), .B(n5292), .Z(n5294) );
  XOR U4643 ( .A(n5295), .B(n5296), .Z(n5292) );
  AND U4644 ( .A(n1538), .B(n5297), .Z(n5296) );
  IV U4645 ( .A(n5289), .Z(n5291) );
  XOR U4646 ( .A(n5298), .B(n5299), .Z(n5289) );
  AND U4647 ( .A(n1542), .B(n5300), .Z(n5299) );
  XOR U4648 ( .A(n5301), .B(n5302), .Z(n5287) );
  AND U4649 ( .A(n1546), .B(n5300), .Z(n5302) );
  XNOR U4650 ( .A(n5301), .B(n5298), .Z(n5300) );
  XOR U4651 ( .A(n5303), .B(n5304), .Z(n5298) );
  AND U4652 ( .A(n1549), .B(n5297), .Z(n5304) );
  XNOR U4653 ( .A(n5305), .B(n5295), .Z(n5297) );
  XOR U4654 ( .A(n5306), .B(n5307), .Z(n5295) );
  AND U4655 ( .A(n1553), .B(n5308), .Z(n5307) );
  XOR U4656 ( .A(p_input[1255]), .B(n5306), .Z(n5308) );
  XOR U4657 ( .A(n5309), .B(n5310), .Z(n5306) );
  AND U4658 ( .A(n1557), .B(n5311), .Z(n5310) );
  IV U4659 ( .A(n5303), .Z(n5305) );
  XOR U4660 ( .A(n5312), .B(n5313), .Z(n5303) );
  AND U4661 ( .A(n1561), .B(n5314), .Z(n5313) );
  XOR U4662 ( .A(n5315), .B(n5316), .Z(n5301) );
  AND U4663 ( .A(n1565), .B(n5314), .Z(n5316) );
  XNOR U4664 ( .A(n5315), .B(n5312), .Z(n5314) );
  XOR U4665 ( .A(n5317), .B(n5318), .Z(n5312) );
  AND U4666 ( .A(n1568), .B(n5311), .Z(n5318) );
  XNOR U4667 ( .A(n5319), .B(n5309), .Z(n5311) );
  XOR U4668 ( .A(n5320), .B(n5321), .Z(n5309) );
  AND U4669 ( .A(n1572), .B(n5322), .Z(n5321) );
  XOR U4670 ( .A(p_input[1271]), .B(n5320), .Z(n5322) );
  XOR U4671 ( .A(n5323), .B(n5324), .Z(n5320) );
  AND U4672 ( .A(n1576), .B(n5325), .Z(n5324) );
  IV U4673 ( .A(n5317), .Z(n5319) );
  XOR U4674 ( .A(n5326), .B(n5327), .Z(n5317) );
  AND U4675 ( .A(n1580), .B(n5328), .Z(n5327) );
  XOR U4676 ( .A(n5329), .B(n5330), .Z(n5315) );
  AND U4677 ( .A(n1584), .B(n5328), .Z(n5330) );
  XNOR U4678 ( .A(n5329), .B(n5326), .Z(n5328) );
  XOR U4679 ( .A(n5331), .B(n5332), .Z(n5326) );
  AND U4680 ( .A(n1587), .B(n5325), .Z(n5332) );
  XNOR U4681 ( .A(n5333), .B(n5323), .Z(n5325) );
  XOR U4682 ( .A(n5334), .B(n5335), .Z(n5323) );
  AND U4683 ( .A(n1591), .B(n5336), .Z(n5335) );
  XOR U4684 ( .A(p_input[1287]), .B(n5334), .Z(n5336) );
  XOR U4685 ( .A(n5337), .B(n5338), .Z(n5334) );
  AND U4686 ( .A(n1595), .B(n5339), .Z(n5338) );
  IV U4687 ( .A(n5331), .Z(n5333) );
  XOR U4688 ( .A(n5340), .B(n5341), .Z(n5331) );
  AND U4689 ( .A(n1599), .B(n5342), .Z(n5341) );
  XOR U4690 ( .A(n5343), .B(n5344), .Z(n5329) );
  AND U4691 ( .A(n1603), .B(n5342), .Z(n5344) );
  XNOR U4692 ( .A(n5343), .B(n5340), .Z(n5342) );
  XOR U4693 ( .A(n5345), .B(n5346), .Z(n5340) );
  AND U4694 ( .A(n1606), .B(n5339), .Z(n5346) );
  XNOR U4695 ( .A(n5347), .B(n5337), .Z(n5339) );
  XOR U4696 ( .A(n5348), .B(n5349), .Z(n5337) );
  AND U4697 ( .A(n1610), .B(n5350), .Z(n5349) );
  XOR U4698 ( .A(p_input[1303]), .B(n5348), .Z(n5350) );
  XOR U4699 ( .A(n5351), .B(n5352), .Z(n5348) );
  AND U4700 ( .A(n1614), .B(n5353), .Z(n5352) );
  IV U4701 ( .A(n5345), .Z(n5347) );
  XOR U4702 ( .A(n5354), .B(n5355), .Z(n5345) );
  AND U4703 ( .A(n1618), .B(n5356), .Z(n5355) );
  XOR U4704 ( .A(n5357), .B(n5358), .Z(n5343) );
  AND U4705 ( .A(n1622), .B(n5356), .Z(n5358) );
  XNOR U4706 ( .A(n5357), .B(n5354), .Z(n5356) );
  XOR U4707 ( .A(n5359), .B(n5360), .Z(n5354) );
  AND U4708 ( .A(n1625), .B(n5353), .Z(n5360) );
  XNOR U4709 ( .A(n5361), .B(n5351), .Z(n5353) );
  XOR U4710 ( .A(n5362), .B(n5363), .Z(n5351) );
  AND U4711 ( .A(n1629), .B(n5364), .Z(n5363) );
  XOR U4712 ( .A(p_input[1319]), .B(n5362), .Z(n5364) );
  XOR U4713 ( .A(n5365), .B(n5366), .Z(n5362) );
  AND U4714 ( .A(n1633), .B(n5367), .Z(n5366) );
  IV U4715 ( .A(n5359), .Z(n5361) );
  XOR U4716 ( .A(n5368), .B(n5369), .Z(n5359) );
  AND U4717 ( .A(n1637), .B(n5370), .Z(n5369) );
  XOR U4718 ( .A(n5371), .B(n5372), .Z(n5357) );
  AND U4719 ( .A(n1641), .B(n5370), .Z(n5372) );
  XNOR U4720 ( .A(n5371), .B(n5368), .Z(n5370) );
  XOR U4721 ( .A(n5373), .B(n5374), .Z(n5368) );
  AND U4722 ( .A(n1644), .B(n5367), .Z(n5374) );
  XNOR U4723 ( .A(n5375), .B(n5365), .Z(n5367) );
  XOR U4724 ( .A(n5376), .B(n5377), .Z(n5365) );
  AND U4725 ( .A(n1648), .B(n5378), .Z(n5377) );
  XOR U4726 ( .A(p_input[1335]), .B(n5376), .Z(n5378) );
  XOR U4727 ( .A(n5379), .B(n5380), .Z(n5376) );
  AND U4728 ( .A(n1652), .B(n5381), .Z(n5380) );
  IV U4729 ( .A(n5373), .Z(n5375) );
  XOR U4730 ( .A(n5382), .B(n5383), .Z(n5373) );
  AND U4731 ( .A(n1656), .B(n5384), .Z(n5383) );
  XOR U4732 ( .A(n5385), .B(n5386), .Z(n5371) );
  AND U4733 ( .A(n1660), .B(n5384), .Z(n5386) );
  XNOR U4734 ( .A(n5385), .B(n5382), .Z(n5384) );
  XOR U4735 ( .A(n5387), .B(n5388), .Z(n5382) );
  AND U4736 ( .A(n1663), .B(n5381), .Z(n5388) );
  XNOR U4737 ( .A(n5389), .B(n5379), .Z(n5381) );
  XOR U4738 ( .A(n5390), .B(n5391), .Z(n5379) );
  AND U4739 ( .A(n1667), .B(n5392), .Z(n5391) );
  XOR U4740 ( .A(p_input[1351]), .B(n5390), .Z(n5392) );
  XOR U4741 ( .A(n5393), .B(n5394), .Z(n5390) );
  AND U4742 ( .A(n1671), .B(n5395), .Z(n5394) );
  IV U4743 ( .A(n5387), .Z(n5389) );
  XOR U4744 ( .A(n5396), .B(n5397), .Z(n5387) );
  AND U4745 ( .A(n1675), .B(n5398), .Z(n5397) );
  XOR U4746 ( .A(n5399), .B(n5400), .Z(n5385) );
  AND U4747 ( .A(n1679), .B(n5398), .Z(n5400) );
  XNOR U4748 ( .A(n5399), .B(n5396), .Z(n5398) );
  XOR U4749 ( .A(n5401), .B(n5402), .Z(n5396) );
  AND U4750 ( .A(n1682), .B(n5395), .Z(n5402) );
  XNOR U4751 ( .A(n5403), .B(n5393), .Z(n5395) );
  XOR U4752 ( .A(n5404), .B(n5405), .Z(n5393) );
  AND U4753 ( .A(n1686), .B(n5406), .Z(n5405) );
  XOR U4754 ( .A(p_input[1367]), .B(n5404), .Z(n5406) );
  XOR U4755 ( .A(n5407), .B(n5408), .Z(n5404) );
  AND U4756 ( .A(n1690), .B(n5409), .Z(n5408) );
  IV U4757 ( .A(n5401), .Z(n5403) );
  XOR U4758 ( .A(n5410), .B(n5411), .Z(n5401) );
  AND U4759 ( .A(n1694), .B(n5412), .Z(n5411) );
  XOR U4760 ( .A(n5413), .B(n5414), .Z(n5399) );
  AND U4761 ( .A(n1698), .B(n5412), .Z(n5414) );
  XNOR U4762 ( .A(n5413), .B(n5410), .Z(n5412) );
  XOR U4763 ( .A(n5415), .B(n5416), .Z(n5410) );
  AND U4764 ( .A(n1701), .B(n5409), .Z(n5416) );
  XNOR U4765 ( .A(n5417), .B(n5407), .Z(n5409) );
  XOR U4766 ( .A(n5418), .B(n5419), .Z(n5407) );
  AND U4767 ( .A(n1705), .B(n5420), .Z(n5419) );
  XOR U4768 ( .A(p_input[1383]), .B(n5418), .Z(n5420) );
  XOR U4769 ( .A(n5421), .B(n5422), .Z(n5418) );
  AND U4770 ( .A(n1709), .B(n5423), .Z(n5422) );
  IV U4771 ( .A(n5415), .Z(n5417) );
  XOR U4772 ( .A(n5424), .B(n5425), .Z(n5415) );
  AND U4773 ( .A(n1713), .B(n5426), .Z(n5425) );
  XOR U4774 ( .A(n5427), .B(n5428), .Z(n5413) );
  AND U4775 ( .A(n1717), .B(n5426), .Z(n5428) );
  XNOR U4776 ( .A(n5427), .B(n5424), .Z(n5426) );
  XOR U4777 ( .A(n5429), .B(n5430), .Z(n5424) );
  AND U4778 ( .A(n1720), .B(n5423), .Z(n5430) );
  XNOR U4779 ( .A(n5431), .B(n5421), .Z(n5423) );
  XOR U4780 ( .A(n5432), .B(n5433), .Z(n5421) );
  AND U4781 ( .A(n1724), .B(n5434), .Z(n5433) );
  XOR U4782 ( .A(p_input[1399]), .B(n5432), .Z(n5434) );
  XOR U4783 ( .A(n5435), .B(n5436), .Z(n5432) );
  AND U4784 ( .A(n1728), .B(n5437), .Z(n5436) );
  IV U4785 ( .A(n5429), .Z(n5431) );
  XOR U4786 ( .A(n5438), .B(n5439), .Z(n5429) );
  AND U4787 ( .A(n1732), .B(n5440), .Z(n5439) );
  XOR U4788 ( .A(n5441), .B(n5442), .Z(n5427) );
  AND U4789 ( .A(n1736), .B(n5440), .Z(n5442) );
  XNOR U4790 ( .A(n5441), .B(n5438), .Z(n5440) );
  XOR U4791 ( .A(n5443), .B(n5444), .Z(n5438) );
  AND U4792 ( .A(n1739), .B(n5437), .Z(n5444) );
  XNOR U4793 ( .A(n5445), .B(n5435), .Z(n5437) );
  XOR U4794 ( .A(n5446), .B(n5447), .Z(n5435) );
  AND U4795 ( .A(n1743), .B(n5448), .Z(n5447) );
  XOR U4796 ( .A(p_input[1415]), .B(n5446), .Z(n5448) );
  XOR U4797 ( .A(n5449), .B(n5450), .Z(n5446) );
  AND U4798 ( .A(n1747), .B(n5451), .Z(n5450) );
  IV U4799 ( .A(n5443), .Z(n5445) );
  XOR U4800 ( .A(n5452), .B(n5453), .Z(n5443) );
  AND U4801 ( .A(n1751), .B(n5454), .Z(n5453) );
  XOR U4802 ( .A(n5455), .B(n5456), .Z(n5441) );
  AND U4803 ( .A(n1755), .B(n5454), .Z(n5456) );
  XNOR U4804 ( .A(n5455), .B(n5452), .Z(n5454) );
  XOR U4805 ( .A(n5457), .B(n5458), .Z(n5452) );
  AND U4806 ( .A(n1758), .B(n5451), .Z(n5458) );
  XNOR U4807 ( .A(n5459), .B(n5449), .Z(n5451) );
  XOR U4808 ( .A(n5460), .B(n5461), .Z(n5449) );
  AND U4809 ( .A(n1762), .B(n5462), .Z(n5461) );
  XOR U4810 ( .A(p_input[1431]), .B(n5460), .Z(n5462) );
  XOR U4811 ( .A(n5463), .B(n5464), .Z(n5460) );
  AND U4812 ( .A(n1766), .B(n5465), .Z(n5464) );
  IV U4813 ( .A(n5457), .Z(n5459) );
  XOR U4814 ( .A(n5466), .B(n5467), .Z(n5457) );
  AND U4815 ( .A(n1770), .B(n5468), .Z(n5467) );
  XOR U4816 ( .A(n5469), .B(n5470), .Z(n5455) );
  AND U4817 ( .A(n1774), .B(n5468), .Z(n5470) );
  XNOR U4818 ( .A(n5469), .B(n5466), .Z(n5468) );
  XOR U4819 ( .A(n5471), .B(n5472), .Z(n5466) );
  AND U4820 ( .A(n1777), .B(n5465), .Z(n5472) );
  XNOR U4821 ( .A(n5473), .B(n5463), .Z(n5465) );
  XOR U4822 ( .A(n5474), .B(n5475), .Z(n5463) );
  AND U4823 ( .A(n1781), .B(n5476), .Z(n5475) );
  XOR U4824 ( .A(p_input[1447]), .B(n5474), .Z(n5476) );
  XOR U4825 ( .A(n5477), .B(n5478), .Z(n5474) );
  AND U4826 ( .A(n1785), .B(n5479), .Z(n5478) );
  IV U4827 ( .A(n5471), .Z(n5473) );
  XOR U4828 ( .A(n5480), .B(n5481), .Z(n5471) );
  AND U4829 ( .A(n1789), .B(n5482), .Z(n5481) );
  XOR U4830 ( .A(n5483), .B(n5484), .Z(n5469) );
  AND U4831 ( .A(n1793), .B(n5482), .Z(n5484) );
  XNOR U4832 ( .A(n5483), .B(n5480), .Z(n5482) );
  XOR U4833 ( .A(n5485), .B(n5486), .Z(n5480) );
  AND U4834 ( .A(n1796), .B(n5479), .Z(n5486) );
  XNOR U4835 ( .A(n5487), .B(n5477), .Z(n5479) );
  XOR U4836 ( .A(n5488), .B(n5489), .Z(n5477) );
  AND U4837 ( .A(n1800), .B(n5490), .Z(n5489) );
  XOR U4838 ( .A(p_input[1463]), .B(n5488), .Z(n5490) );
  XOR U4839 ( .A(n5491), .B(n5492), .Z(n5488) );
  AND U4840 ( .A(n1804), .B(n5493), .Z(n5492) );
  IV U4841 ( .A(n5485), .Z(n5487) );
  XOR U4842 ( .A(n5494), .B(n5495), .Z(n5485) );
  AND U4843 ( .A(n1808), .B(n5496), .Z(n5495) );
  XOR U4844 ( .A(n5497), .B(n5498), .Z(n5483) );
  AND U4845 ( .A(n1812), .B(n5496), .Z(n5498) );
  XNOR U4846 ( .A(n5497), .B(n5494), .Z(n5496) );
  XOR U4847 ( .A(n5499), .B(n5500), .Z(n5494) );
  AND U4848 ( .A(n1815), .B(n5493), .Z(n5500) );
  XNOR U4849 ( .A(n5501), .B(n5491), .Z(n5493) );
  XOR U4850 ( .A(n5502), .B(n5503), .Z(n5491) );
  AND U4851 ( .A(n1819), .B(n5504), .Z(n5503) );
  XOR U4852 ( .A(p_input[1479]), .B(n5502), .Z(n5504) );
  XOR U4853 ( .A(n5505), .B(n5506), .Z(n5502) );
  AND U4854 ( .A(n1823), .B(n5507), .Z(n5506) );
  IV U4855 ( .A(n5499), .Z(n5501) );
  XOR U4856 ( .A(n5508), .B(n5509), .Z(n5499) );
  AND U4857 ( .A(n1827), .B(n5510), .Z(n5509) );
  XOR U4858 ( .A(n5511), .B(n5512), .Z(n5497) );
  AND U4859 ( .A(n1831), .B(n5510), .Z(n5512) );
  XNOR U4860 ( .A(n5511), .B(n5508), .Z(n5510) );
  XOR U4861 ( .A(n5513), .B(n5514), .Z(n5508) );
  AND U4862 ( .A(n1834), .B(n5507), .Z(n5514) );
  XNOR U4863 ( .A(n5515), .B(n5505), .Z(n5507) );
  XOR U4864 ( .A(n5516), .B(n5517), .Z(n5505) );
  AND U4865 ( .A(n1838), .B(n5518), .Z(n5517) );
  XOR U4866 ( .A(p_input[1495]), .B(n5516), .Z(n5518) );
  XOR U4867 ( .A(n5519), .B(n5520), .Z(n5516) );
  AND U4868 ( .A(n1842), .B(n5521), .Z(n5520) );
  IV U4869 ( .A(n5513), .Z(n5515) );
  XOR U4870 ( .A(n5522), .B(n5523), .Z(n5513) );
  AND U4871 ( .A(n1846), .B(n5524), .Z(n5523) );
  XOR U4872 ( .A(n5525), .B(n5526), .Z(n5511) );
  AND U4873 ( .A(n1850), .B(n5524), .Z(n5526) );
  XNOR U4874 ( .A(n5525), .B(n5522), .Z(n5524) );
  XOR U4875 ( .A(n5527), .B(n5528), .Z(n5522) );
  AND U4876 ( .A(n1853), .B(n5521), .Z(n5528) );
  XNOR U4877 ( .A(n5529), .B(n5519), .Z(n5521) );
  XOR U4878 ( .A(n5530), .B(n5531), .Z(n5519) );
  AND U4879 ( .A(n1857), .B(n5532), .Z(n5531) );
  XOR U4880 ( .A(p_input[1511]), .B(n5530), .Z(n5532) );
  XOR U4881 ( .A(n5533), .B(n5534), .Z(n5530) );
  AND U4882 ( .A(n1861), .B(n5535), .Z(n5534) );
  IV U4883 ( .A(n5527), .Z(n5529) );
  XOR U4884 ( .A(n5536), .B(n5537), .Z(n5527) );
  AND U4885 ( .A(n1865), .B(n5538), .Z(n5537) );
  XOR U4886 ( .A(n5539), .B(n5540), .Z(n5525) );
  AND U4887 ( .A(n1869), .B(n5538), .Z(n5540) );
  XNOR U4888 ( .A(n5539), .B(n5536), .Z(n5538) );
  XOR U4889 ( .A(n5541), .B(n5542), .Z(n5536) );
  AND U4890 ( .A(n1872), .B(n5535), .Z(n5542) );
  XNOR U4891 ( .A(n5543), .B(n5533), .Z(n5535) );
  XOR U4892 ( .A(n5544), .B(n5545), .Z(n5533) );
  AND U4893 ( .A(n1876), .B(n5546), .Z(n5545) );
  XOR U4894 ( .A(p_input[1527]), .B(n5544), .Z(n5546) );
  XOR U4895 ( .A(n5547), .B(n5548), .Z(n5544) );
  AND U4896 ( .A(n1880), .B(n5549), .Z(n5548) );
  IV U4897 ( .A(n5541), .Z(n5543) );
  XOR U4898 ( .A(n5550), .B(n5551), .Z(n5541) );
  AND U4899 ( .A(n1884), .B(n5552), .Z(n5551) );
  XOR U4900 ( .A(n5553), .B(n5554), .Z(n5539) );
  AND U4901 ( .A(n1888), .B(n5552), .Z(n5554) );
  XNOR U4902 ( .A(n5553), .B(n5550), .Z(n5552) );
  XOR U4903 ( .A(n5555), .B(n5556), .Z(n5550) );
  AND U4904 ( .A(n1891), .B(n5549), .Z(n5556) );
  XNOR U4905 ( .A(n5557), .B(n5547), .Z(n5549) );
  XOR U4906 ( .A(n5558), .B(n5559), .Z(n5547) );
  AND U4907 ( .A(n1895), .B(n5560), .Z(n5559) );
  XOR U4908 ( .A(p_input[1543]), .B(n5558), .Z(n5560) );
  XOR U4909 ( .A(n5561), .B(n5562), .Z(n5558) );
  AND U4910 ( .A(n1899), .B(n5563), .Z(n5562) );
  IV U4911 ( .A(n5555), .Z(n5557) );
  XOR U4912 ( .A(n5564), .B(n5565), .Z(n5555) );
  AND U4913 ( .A(n1903), .B(n5566), .Z(n5565) );
  XOR U4914 ( .A(n5567), .B(n5568), .Z(n5553) );
  AND U4915 ( .A(n1907), .B(n5566), .Z(n5568) );
  XNOR U4916 ( .A(n5567), .B(n5564), .Z(n5566) );
  XOR U4917 ( .A(n5569), .B(n5570), .Z(n5564) );
  AND U4918 ( .A(n1910), .B(n5563), .Z(n5570) );
  XNOR U4919 ( .A(n5571), .B(n5561), .Z(n5563) );
  XOR U4920 ( .A(n5572), .B(n5573), .Z(n5561) );
  AND U4921 ( .A(n1914), .B(n5574), .Z(n5573) );
  XOR U4922 ( .A(p_input[1559]), .B(n5572), .Z(n5574) );
  XOR U4923 ( .A(n5575), .B(n5576), .Z(n5572) );
  AND U4924 ( .A(n1918), .B(n5577), .Z(n5576) );
  IV U4925 ( .A(n5569), .Z(n5571) );
  XOR U4926 ( .A(n5578), .B(n5579), .Z(n5569) );
  AND U4927 ( .A(n1922), .B(n5580), .Z(n5579) );
  XOR U4928 ( .A(n5581), .B(n5582), .Z(n5567) );
  AND U4929 ( .A(n1926), .B(n5580), .Z(n5582) );
  XNOR U4930 ( .A(n5581), .B(n5578), .Z(n5580) );
  XOR U4931 ( .A(n5583), .B(n5584), .Z(n5578) );
  AND U4932 ( .A(n1929), .B(n5577), .Z(n5584) );
  XNOR U4933 ( .A(n5585), .B(n5575), .Z(n5577) );
  XOR U4934 ( .A(n5586), .B(n5587), .Z(n5575) );
  AND U4935 ( .A(n1933), .B(n5588), .Z(n5587) );
  XOR U4936 ( .A(p_input[1575]), .B(n5586), .Z(n5588) );
  XOR U4937 ( .A(n5589), .B(n5590), .Z(n5586) );
  AND U4938 ( .A(n1937), .B(n5591), .Z(n5590) );
  IV U4939 ( .A(n5583), .Z(n5585) );
  XOR U4940 ( .A(n5592), .B(n5593), .Z(n5583) );
  AND U4941 ( .A(n1941), .B(n5594), .Z(n5593) );
  XOR U4942 ( .A(n5595), .B(n5596), .Z(n5581) );
  AND U4943 ( .A(n1945), .B(n5594), .Z(n5596) );
  XNOR U4944 ( .A(n5595), .B(n5592), .Z(n5594) );
  XOR U4945 ( .A(n5597), .B(n5598), .Z(n5592) );
  AND U4946 ( .A(n1948), .B(n5591), .Z(n5598) );
  XNOR U4947 ( .A(n5599), .B(n5589), .Z(n5591) );
  XOR U4948 ( .A(n5600), .B(n5601), .Z(n5589) );
  AND U4949 ( .A(n1952), .B(n5602), .Z(n5601) );
  XOR U4950 ( .A(p_input[1591]), .B(n5600), .Z(n5602) );
  XOR U4951 ( .A(n5603), .B(n5604), .Z(n5600) );
  AND U4952 ( .A(n1956), .B(n5605), .Z(n5604) );
  IV U4953 ( .A(n5597), .Z(n5599) );
  XOR U4954 ( .A(n5606), .B(n5607), .Z(n5597) );
  AND U4955 ( .A(n1960), .B(n5608), .Z(n5607) );
  XOR U4956 ( .A(n5609), .B(n5610), .Z(n5595) );
  AND U4957 ( .A(n1964), .B(n5608), .Z(n5610) );
  XNOR U4958 ( .A(n5609), .B(n5606), .Z(n5608) );
  XOR U4959 ( .A(n5611), .B(n5612), .Z(n5606) );
  AND U4960 ( .A(n1967), .B(n5605), .Z(n5612) );
  XNOR U4961 ( .A(n5613), .B(n5603), .Z(n5605) );
  XOR U4962 ( .A(n5614), .B(n5615), .Z(n5603) );
  AND U4963 ( .A(n1971), .B(n5616), .Z(n5615) );
  XOR U4964 ( .A(p_input[1607]), .B(n5614), .Z(n5616) );
  XOR U4965 ( .A(n5617), .B(n5618), .Z(n5614) );
  AND U4966 ( .A(n1975), .B(n5619), .Z(n5618) );
  IV U4967 ( .A(n5611), .Z(n5613) );
  XOR U4968 ( .A(n5620), .B(n5621), .Z(n5611) );
  AND U4969 ( .A(n1979), .B(n5622), .Z(n5621) );
  XOR U4970 ( .A(n5623), .B(n5624), .Z(n5609) );
  AND U4971 ( .A(n1983), .B(n5622), .Z(n5624) );
  XNOR U4972 ( .A(n5623), .B(n5620), .Z(n5622) );
  XOR U4973 ( .A(n5625), .B(n5626), .Z(n5620) );
  AND U4974 ( .A(n1986), .B(n5619), .Z(n5626) );
  XNOR U4975 ( .A(n5627), .B(n5617), .Z(n5619) );
  XOR U4976 ( .A(n5628), .B(n5629), .Z(n5617) );
  AND U4977 ( .A(n1990), .B(n5630), .Z(n5629) );
  XOR U4978 ( .A(p_input[1623]), .B(n5628), .Z(n5630) );
  XOR U4979 ( .A(n5631), .B(n5632), .Z(n5628) );
  AND U4980 ( .A(n1994), .B(n5633), .Z(n5632) );
  IV U4981 ( .A(n5625), .Z(n5627) );
  XOR U4982 ( .A(n5634), .B(n5635), .Z(n5625) );
  AND U4983 ( .A(n1998), .B(n5636), .Z(n5635) );
  XOR U4984 ( .A(n5637), .B(n5638), .Z(n5623) );
  AND U4985 ( .A(n2002), .B(n5636), .Z(n5638) );
  XNOR U4986 ( .A(n5637), .B(n5634), .Z(n5636) );
  XOR U4987 ( .A(n5639), .B(n5640), .Z(n5634) );
  AND U4988 ( .A(n2005), .B(n5633), .Z(n5640) );
  XNOR U4989 ( .A(n5641), .B(n5631), .Z(n5633) );
  XOR U4990 ( .A(n5642), .B(n5643), .Z(n5631) );
  AND U4991 ( .A(n2009), .B(n5644), .Z(n5643) );
  XOR U4992 ( .A(p_input[1639]), .B(n5642), .Z(n5644) );
  XOR U4993 ( .A(n5645), .B(n5646), .Z(n5642) );
  AND U4994 ( .A(n2013), .B(n5647), .Z(n5646) );
  IV U4995 ( .A(n5639), .Z(n5641) );
  XOR U4996 ( .A(n5648), .B(n5649), .Z(n5639) );
  AND U4997 ( .A(n2017), .B(n5650), .Z(n5649) );
  XOR U4998 ( .A(n5651), .B(n5652), .Z(n5637) );
  AND U4999 ( .A(n2021), .B(n5650), .Z(n5652) );
  XNOR U5000 ( .A(n5651), .B(n5648), .Z(n5650) );
  XOR U5001 ( .A(n5653), .B(n5654), .Z(n5648) );
  AND U5002 ( .A(n2024), .B(n5647), .Z(n5654) );
  XNOR U5003 ( .A(n5655), .B(n5645), .Z(n5647) );
  XOR U5004 ( .A(n5656), .B(n5657), .Z(n5645) );
  AND U5005 ( .A(n2028), .B(n5658), .Z(n5657) );
  XOR U5006 ( .A(p_input[1655]), .B(n5656), .Z(n5658) );
  XOR U5007 ( .A(n5659), .B(n5660), .Z(n5656) );
  AND U5008 ( .A(n2032), .B(n5661), .Z(n5660) );
  IV U5009 ( .A(n5653), .Z(n5655) );
  XOR U5010 ( .A(n5662), .B(n5663), .Z(n5653) );
  AND U5011 ( .A(n2036), .B(n5664), .Z(n5663) );
  XOR U5012 ( .A(n5665), .B(n5666), .Z(n5651) );
  AND U5013 ( .A(n2040), .B(n5664), .Z(n5666) );
  XNOR U5014 ( .A(n5665), .B(n5662), .Z(n5664) );
  XOR U5015 ( .A(n5667), .B(n5668), .Z(n5662) );
  AND U5016 ( .A(n2043), .B(n5661), .Z(n5668) );
  XNOR U5017 ( .A(n5669), .B(n5659), .Z(n5661) );
  XOR U5018 ( .A(n5670), .B(n5671), .Z(n5659) );
  AND U5019 ( .A(n2047), .B(n5672), .Z(n5671) );
  XOR U5020 ( .A(p_input[1671]), .B(n5670), .Z(n5672) );
  XOR U5021 ( .A(n5673), .B(n5674), .Z(n5670) );
  AND U5022 ( .A(n2051), .B(n5675), .Z(n5674) );
  IV U5023 ( .A(n5667), .Z(n5669) );
  XOR U5024 ( .A(n5676), .B(n5677), .Z(n5667) );
  AND U5025 ( .A(n2055), .B(n5678), .Z(n5677) );
  XOR U5026 ( .A(n5679), .B(n5680), .Z(n5665) );
  AND U5027 ( .A(n2059), .B(n5678), .Z(n5680) );
  XNOR U5028 ( .A(n5679), .B(n5676), .Z(n5678) );
  XOR U5029 ( .A(n5681), .B(n5682), .Z(n5676) );
  AND U5030 ( .A(n2062), .B(n5675), .Z(n5682) );
  XNOR U5031 ( .A(n5683), .B(n5673), .Z(n5675) );
  XOR U5032 ( .A(n5684), .B(n5685), .Z(n5673) );
  AND U5033 ( .A(n2066), .B(n5686), .Z(n5685) );
  XOR U5034 ( .A(p_input[1687]), .B(n5684), .Z(n5686) );
  XOR U5035 ( .A(n5687), .B(n5688), .Z(n5684) );
  AND U5036 ( .A(n2070), .B(n5689), .Z(n5688) );
  IV U5037 ( .A(n5681), .Z(n5683) );
  XOR U5038 ( .A(n5690), .B(n5691), .Z(n5681) );
  AND U5039 ( .A(n2074), .B(n5692), .Z(n5691) );
  XOR U5040 ( .A(n5693), .B(n5694), .Z(n5679) );
  AND U5041 ( .A(n2078), .B(n5692), .Z(n5694) );
  XNOR U5042 ( .A(n5693), .B(n5690), .Z(n5692) );
  XOR U5043 ( .A(n5695), .B(n5696), .Z(n5690) );
  AND U5044 ( .A(n2081), .B(n5689), .Z(n5696) );
  XNOR U5045 ( .A(n5697), .B(n5687), .Z(n5689) );
  XOR U5046 ( .A(n5698), .B(n5699), .Z(n5687) );
  AND U5047 ( .A(n2085), .B(n5700), .Z(n5699) );
  XOR U5048 ( .A(p_input[1703]), .B(n5698), .Z(n5700) );
  XOR U5049 ( .A(n5701), .B(n5702), .Z(n5698) );
  AND U5050 ( .A(n2089), .B(n5703), .Z(n5702) );
  IV U5051 ( .A(n5695), .Z(n5697) );
  XOR U5052 ( .A(n5704), .B(n5705), .Z(n5695) );
  AND U5053 ( .A(n2093), .B(n5706), .Z(n5705) );
  XOR U5054 ( .A(n5707), .B(n5708), .Z(n5693) );
  AND U5055 ( .A(n2097), .B(n5706), .Z(n5708) );
  XNOR U5056 ( .A(n5707), .B(n5704), .Z(n5706) );
  XOR U5057 ( .A(n5709), .B(n5710), .Z(n5704) );
  AND U5058 ( .A(n2100), .B(n5703), .Z(n5710) );
  XNOR U5059 ( .A(n5711), .B(n5701), .Z(n5703) );
  XOR U5060 ( .A(n5712), .B(n5713), .Z(n5701) );
  AND U5061 ( .A(n2104), .B(n5714), .Z(n5713) );
  XOR U5062 ( .A(p_input[1719]), .B(n5712), .Z(n5714) );
  XOR U5063 ( .A(n5715), .B(n5716), .Z(n5712) );
  AND U5064 ( .A(n2108), .B(n5717), .Z(n5716) );
  IV U5065 ( .A(n5709), .Z(n5711) );
  XOR U5066 ( .A(n5718), .B(n5719), .Z(n5709) );
  AND U5067 ( .A(n2112), .B(n5720), .Z(n5719) );
  XOR U5068 ( .A(n5721), .B(n5722), .Z(n5707) );
  AND U5069 ( .A(n2116), .B(n5720), .Z(n5722) );
  XNOR U5070 ( .A(n5721), .B(n5718), .Z(n5720) );
  XOR U5071 ( .A(n5723), .B(n5724), .Z(n5718) );
  AND U5072 ( .A(n2119), .B(n5717), .Z(n5724) );
  XNOR U5073 ( .A(n5725), .B(n5715), .Z(n5717) );
  XOR U5074 ( .A(n5726), .B(n5727), .Z(n5715) );
  AND U5075 ( .A(n2123), .B(n5728), .Z(n5727) );
  XOR U5076 ( .A(p_input[1735]), .B(n5726), .Z(n5728) );
  XOR U5077 ( .A(n5729), .B(n5730), .Z(n5726) );
  AND U5078 ( .A(n2127), .B(n5731), .Z(n5730) );
  IV U5079 ( .A(n5723), .Z(n5725) );
  XOR U5080 ( .A(n5732), .B(n5733), .Z(n5723) );
  AND U5081 ( .A(n2131), .B(n5734), .Z(n5733) );
  XOR U5082 ( .A(n5735), .B(n5736), .Z(n5721) );
  AND U5083 ( .A(n2135), .B(n5734), .Z(n5736) );
  XNOR U5084 ( .A(n5735), .B(n5732), .Z(n5734) );
  XOR U5085 ( .A(n5737), .B(n5738), .Z(n5732) );
  AND U5086 ( .A(n2138), .B(n5731), .Z(n5738) );
  XNOR U5087 ( .A(n5739), .B(n5729), .Z(n5731) );
  XOR U5088 ( .A(n5740), .B(n5741), .Z(n5729) );
  AND U5089 ( .A(n2142), .B(n5742), .Z(n5741) );
  XOR U5090 ( .A(p_input[1751]), .B(n5740), .Z(n5742) );
  XOR U5091 ( .A(n5743), .B(n5744), .Z(n5740) );
  AND U5092 ( .A(n2146), .B(n5745), .Z(n5744) );
  IV U5093 ( .A(n5737), .Z(n5739) );
  XOR U5094 ( .A(n5746), .B(n5747), .Z(n5737) );
  AND U5095 ( .A(n2150), .B(n5748), .Z(n5747) );
  XOR U5096 ( .A(n5749), .B(n5750), .Z(n5735) );
  AND U5097 ( .A(n2154), .B(n5748), .Z(n5750) );
  XNOR U5098 ( .A(n5749), .B(n5746), .Z(n5748) );
  XOR U5099 ( .A(n5751), .B(n5752), .Z(n5746) );
  AND U5100 ( .A(n2157), .B(n5745), .Z(n5752) );
  XNOR U5101 ( .A(n5753), .B(n5743), .Z(n5745) );
  XOR U5102 ( .A(n5754), .B(n5755), .Z(n5743) );
  AND U5103 ( .A(n2161), .B(n5756), .Z(n5755) );
  XOR U5104 ( .A(p_input[1767]), .B(n5754), .Z(n5756) );
  XOR U5105 ( .A(n5757), .B(n5758), .Z(n5754) );
  AND U5106 ( .A(n2165), .B(n5759), .Z(n5758) );
  IV U5107 ( .A(n5751), .Z(n5753) );
  XOR U5108 ( .A(n5760), .B(n5761), .Z(n5751) );
  AND U5109 ( .A(n2169), .B(n5762), .Z(n5761) );
  XOR U5110 ( .A(n5763), .B(n5764), .Z(n5749) );
  AND U5111 ( .A(n2173), .B(n5762), .Z(n5764) );
  XNOR U5112 ( .A(n5763), .B(n5760), .Z(n5762) );
  XOR U5113 ( .A(n5765), .B(n5766), .Z(n5760) );
  AND U5114 ( .A(n2176), .B(n5759), .Z(n5766) );
  XNOR U5115 ( .A(n5767), .B(n5757), .Z(n5759) );
  XOR U5116 ( .A(n5768), .B(n5769), .Z(n5757) );
  AND U5117 ( .A(n2180), .B(n5770), .Z(n5769) );
  XOR U5118 ( .A(p_input[1783]), .B(n5768), .Z(n5770) );
  XOR U5119 ( .A(n5771), .B(n5772), .Z(n5768) );
  AND U5120 ( .A(n2184), .B(n5773), .Z(n5772) );
  IV U5121 ( .A(n5765), .Z(n5767) );
  XOR U5122 ( .A(n5774), .B(n5775), .Z(n5765) );
  AND U5123 ( .A(n2188), .B(n5776), .Z(n5775) );
  XOR U5124 ( .A(n5777), .B(n5778), .Z(n5763) );
  AND U5125 ( .A(n2192), .B(n5776), .Z(n5778) );
  XNOR U5126 ( .A(n5777), .B(n5774), .Z(n5776) );
  XOR U5127 ( .A(n5779), .B(n5780), .Z(n5774) );
  AND U5128 ( .A(n2195), .B(n5773), .Z(n5780) );
  XNOR U5129 ( .A(n5781), .B(n5771), .Z(n5773) );
  XOR U5130 ( .A(n5782), .B(n5783), .Z(n5771) );
  AND U5131 ( .A(n2199), .B(n5784), .Z(n5783) );
  XOR U5132 ( .A(p_input[1799]), .B(n5782), .Z(n5784) );
  XOR U5133 ( .A(n5785), .B(n5786), .Z(n5782) );
  AND U5134 ( .A(n2203), .B(n5787), .Z(n5786) );
  IV U5135 ( .A(n5779), .Z(n5781) );
  XOR U5136 ( .A(n5788), .B(n5789), .Z(n5779) );
  AND U5137 ( .A(n2207), .B(n5790), .Z(n5789) );
  XOR U5138 ( .A(n5791), .B(n5792), .Z(n5777) );
  AND U5139 ( .A(n2211), .B(n5790), .Z(n5792) );
  XNOR U5140 ( .A(n5791), .B(n5788), .Z(n5790) );
  XOR U5141 ( .A(n5793), .B(n5794), .Z(n5788) );
  AND U5142 ( .A(n2214), .B(n5787), .Z(n5794) );
  XNOR U5143 ( .A(n5795), .B(n5785), .Z(n5787) );
  XOR U5144 ( .A(n5796), .B(n5797), .Z(n5785) );
  AND U5145 ( .A(n2218), .B(n5798), .Z(n5797) );
  XOR U5146 ( .A(p_input[1815]), .B(n5796), .Z(n5798) );
  XOR U5147 ( .A(n5799), .B(n5800), .Z(n5796) );
  AND U5148 ( .A(n2222), .B(n5801), .Z(n5800) );
  IV U5149 ( .A(n5793), .Z(n5795) );
  XOR U5150 ( .A(n5802), .B(n5803), .Z(n5793) );
  AND U5151 ( .A(n2226), .B(n5804), .Z(n5803) );
  XOR U5152 ( .A(n5805), .B(n5806), .Z(n5791) );
  AND U5153 ( .A(n2230), .B(n5804), .Z(n5806) );
  XNOR U5154 ( .A(n5805), .B(n5802), .Z(n5804) );
  XOR U5155 ( .A(n5807), .B(n5808), .Z(n5802) );
  AND U5156 ( .A(n2233), .B(n5801), .Z(n5808) );
  XNOR U5157 ( .A(n5809), .B(n5799), .Z(n5801) );
  XOR U5158 ( .A(n5810), .B(n5811), .Z(n5799) );
  AND U5159 ( .A(n2237), .B(n5812), .Z(n5811) );
  XOR U5160 ( .A(p_input[1831]), .B(n5810), .Z(n5812) );
  XOR U5161 ( .A(n5813), .B(n5814), .Z(n5810) );
  AND U5162 ( .A(n2241), .B(n5815), .Z(n5814) );
  IV U5163 ( .A(n5807), .Z(n5809) );
  XOR U5164 ( .A(n5816), .B(n5817), .Z(n5807) );
  AND U5165 ( .A(n2245), .B(n5818), .Z(n5817) );
  XOR U5166 ( .A(n5819), .B(n5820), .Z(n5805) );
  AND U5167 ( .A(n2249), .B(n5818), .Z(n5820) );
  XNOR U5168 ( .A(n5819), .B(n5816), .Z(n5818) );
  XOR U5169 ( .A(n5821), .B(n5822), .Z(n5816) );
  AND U5170 ( .A(n2252), .B(n5815), .Z(n5822) );
  XNOR U5171 ( .A(n5823), .B(n5813), .Z(n5815) );
  XOR U5172 ( .A(n5824), .B(n5825), .Z(n5813) );
  AND U5173 ( .A(n2256), .B(n5826), .Z(n5825) );
  XOR U5174 ( .A(p_input[1847]), .B(n5824), .Z(n5826) );
  XOR U5175 ( .A(n5827), .B(n5828), .Z(n5824) );
  AND U5176 ( .A(n2260), .B(n5829), .Z(n5828) );
  IV U5177 ( .A(n5821), .Z(n5823) );
  XOR U5178 ( .A(n5830), .B(n5831), .Z(n5821) );
  AND U5179 ( .A(n2264), .B(n5832), .Z(n5831) );
  XOR U5180 ( .A(n5833), .B(n5834), .Z(n5819) );
  AND U5181 ( .A(n2268), .B(n5832), .Z(n5834) );
  XNOR U5182 ( .A(n5833), .B(n5830), .Z(n5832) );
  XOR U5183 ( .A(n5835), .B(n5836), .Z(n5830) );
  AND U5184 ( .A(n2271), .B(n5829), .Z(n5836) );
  XNOR U5185 ( .A(n5837), .B(n5827), .Z(n5829) );
  XOR U5186 ( .A(n5838), .B(n5839), .Z(n5827) );
  AND U5187 ( .A(n2275), .B(n5840), .Z(n5839) );
  XOR U5188 ( .A(p_input[1863]), .B(n5838), .Z(n5840) );
  XOR U5189 ( .A(n5841), .B(n5842), .Z(n5838) );
  AND U5190 ( .A(n2279), .B(n5843), .Z(n5842) );
  IV U5191 ( .A(n5835), .Z(n5837) );
  XOR U5192 ( .A(n5844), .B(n5845), .Z(n5835) );
  AND U5193 ( .A(n2283), .B(n5846), .Z(n5845) );
  XOR U5194 ( .A(n5847), .B(n5848), .Z(n5833) );
  AND U5195 ( .A(n2287), .B(n5846), .Z(n5848) );
  XNOR U5196 ( .A(n5847), .B(n5844), .Z(n5846) );
  XOR U5197 ( .A(n5849), .B(n5850), .Z(n5844) );
  AND U5198 ( .A(n2290), .B(n5843), .Z(n5850) );
  XNOR U5199 ( .A(n5851), .B(n5841), .Z(n5843) );
  XOR U5200 ( .A(n5852), .B(n5853), .Z(n5841) );
  AND U5201 ( .A(n2294), .B(n5854), .Z(n5853) );
  XOR U5202 ( .A(p_input[1879]), .B(n5852), .Z(n5854) );
  XOR U5203 ( .A(n5855), .B(n5856), .Z(n5852) );
  AND U5204 ( .A(n2298), .B(n5857), .Z(n5856) );
  IV U5205 ( .A(n5849), .Z(n5851) );
  XOR U5206 ( .A(n5858), .B(n5859), .Z(n5849) );
  AND U5207 ( .A(n2302), .B(n5860), .Z(n5859) );
  XOR U5208 ( .A(n5861), .B(n5862), .Z(n5847) );
  AND U5209 ( .A(n2306), .B(n5860), .Z(n5862) );
  XNOR U5210 ( .A(n5861), .B(n5858), .Z(n5860) );
  XOR U5211 ( .A(n5863), .B(n5864), .Z(n5858) );
  AND U5212 ( .A(n2309), .B(n5857), .Z(n5864) );
  XNOR U5213 ( .A(n5865), .B(n5855), .Z(n5857) );
  XOR U5214 ( .A(n5866), .B(n5867), .Z(n5855) );
  AND U5215 ( .A(n2313), .B(n5868), .Z(n5867) );
  XOR U5216 ( .A(p_input[1895]), .B(n5866), .Z(n5868) );
  XOR U5217 ( .A(n5869), .B(n5870), .Z(n5866) );
  AND U5218 ( .A(n2317), .B(n5871), .Z(n5870) );
  IV U5219 ( .A(n5863), .Z(n5865) );
  XOR U5220 ( .A(n5872), .B(n5873), .Z(n5863) );
  AND U5221 ( .A(n2321), .B(n5874), .Z(n5873) );
  XOR U5222 ( .A(n5875), .B(n5876), .Z(n5861) );
  AND U5223 ( .A(n2325), .B(n5874), .Z(n5876) );
  XNOR U5224 ( .A(n5875), .B(n5872), .Z(n5874) );
  XOR U5225 ( .A(n5877), .B(n5878), .Z(n5872) );
  AND U5226 ( .A(n2328), .B(n5871), .Z(n5878) );
  XNOR U5227 ( .A(n5879), .B(n5869), .Z(n5871) );
  XOR U5228 ( .A(n5880), .B(n5881), .Z(n5869) );
  AND U5229 ( .A(n2332), .B(n5882), .Z(n5881) );
  XOR U5230 ( .A(p_input[1911]), .B(n5880), .Z(n5882) );
  XOR U5231 ( .A(n5883), .B(n5884), .Z(n5880) );
  AND U5232 ( .A(n2336), .B(n5885), .Z(n5884) );
  IV U5233 ( .A(n5877), .Z(n5879) );
  XOR U5234 ( .A(n5886), .B(n5887), .Z(n5877) );
  AND U5235 ( .A(n2340), .B(n5888), .Z(n5887) );
  XOR U5236 ( .A(n5889), .B(n5890), .Z(n5875) );
  AND U5237 ( .A(n2344), .B(n5888), .Z(n5890) );
  XNOR U5238 ( .A(n5889), .B(n5886), .Z(n5888) );
  XOR U5239 ( .A(n5891), .B(n5892), .Z(n5886) );
  AND U5240 ( .A(n2347), .B(n5885), .Z(n5892) );
  XNOR U5241 ( .A(n5893), .B(n5883), .Z(n5885) );
  XOR U5242 ( .A(n5894), .B(n5895), .Z(n5883) );
  AND U5243 ( .A(n2351), .B(n5896), .Z(n5895) );
  XOR U5244 ( .A(p_input[1927]), .B(n5894), .Z(n5896) );
  XOR U5245 ( .A(n5897), .B(n5898), .Z(n5894) );
  AND U5246 ( .A(n2355), .B(n5899), .Z(n5898) );
  IV U5247 ( .A(n5891), .Z(n5893) );
  XOR U5248 ( .A(n5900), .B(n5901), .Z(n5891) );
  AND U5249 ( .A(n2359), .B(n5902), .Z(n5901) );
  XOR U5250 ( .A(n5903), .B(n5904), .Z(n5889) );
  AND U5251 ( .A(n2363), .B(n5902), .Z(n5904) );
  XNOR U5252 ( .A(n5903), .B(n5900), .Z(n5902) );
  XOR U5253 ( .A(n5905), .B(n5906), .Z(n5900) );
  AND U5254 ( .A(n2366), .B(n5899), .Z(n5906) );
  XNOR U5255 ( .A(n5907), .B(n5897), .Z(n5899) );
  XOR U5256 ( .A(n5908), .B(n5909), .Z(n5897) );
  AND U5257 ( .A(n2370), .B(n5910), .Z(n5909) );
  XOR U5258 ( .A(p_input[1943]), .B(n5908), .Z(n5910) );
  XOR U5259 ( .A(n5911), .B(n5912), .Z(n5908) );
  AND U5260 ( .A(n2374), .B(n5913), .Z(n5912) );
  IV U5261 ( .A(n5905), .Z(n5907) );
  XOR U5262 ( .A(n5914), .B(n5915), .Z(n5905) );
  AND U5263 ( .A(n2378), .B(n5916), .Z(n5915) );
  XOR U5264 ( .A(n5917), .B(n5918), .Z(n5903) );
  AND U5265 ( .A(n2382), .B(n5916), .Z(n5918) );
  XNOR U5266 ( .A(n5917), .B(n5914), .Z(n5916) );
  XOR U5267 ( .A(n5919), .B(n5920), .Z(n5914) );
  AND U5268 ( .A(n2385), .B(n5913), .Z(n5920) );
  XNOR U5269 ( .A(n5921), .B(n5911), .Z(n5913) );
  XOR U5270 ( .A(n5922), .B(n5923), .Z(n5911) );
  AND U5271 ( .A(n2389), .B(n5924), .Z(n5923) );
  XOR U5272 ( .A(p_input[1959]), .B(n5922), .Z(n5924) );
  XOR U5273 ( .A(n5925), .B(n5926), .Z(n5922) );
  AND U5274 ( .A(n2393), .B(n5927), .Z(n5926) );
  IV U5275 ( .A(n5919), .Z(n5921) );
  XOR U5276 ( .A(n5928), .B(n5929), .Z(n5919) );
  AND U5277 ( .A(n2397), .B(n5930), .Z(n5929) );
  XOR U5278 ( .A(n5931), .B(n5932), .Z(n5917) );
  AND U5279 ( .A(n2401), .B(n5930), .Z(n5932) );
  XNOR U5280 ( .A(n5931), .B(n5928), .Z(n5930) );
  XOR U5281 ( .A(n5933), .B(n5934), .Z(n5928) );
  AND U5282 ( .A(n2404), .B(n5927), .Z(n5934) );
  XNOR U5283 ( .A(n5935), .B(n5925), .Z(n5927) );
  XOR U5284 ( .A(n5936), .B(n5937), .Z(n5925) );
  AND U5285 ( .A(n2408), .B(n5938), .Z(n5937) );
  XOR U5286 ( .A(p_input[1975]), .B(n5936), .Z(n5938) );
  XOR U5287 ( .A(n5939), .B(n5940), .Z(n5936) );
  AND U5288 ( .A(n2412), .B(n5941), .Z(n5940) );
  IV U5289 ( .A(n5933), .Z(n5935) );
  XOR U5290 ( .A(n5942), .B(n5943), .Z(n5933) );
  AND U5291 ( .A(n2416), .B(n5944), .Z(n5943) );
  XOR U5292 ( .A(n5945), .B(n5946), .Z(n5931) );
  AND U5293 ( .A(n2420), .B(n5944), .Z(n5946) );
  XNOR U5294 ( .A(n5945), .B(n5942), .Z(n5944) );
  XOR U5295 ( .A(n5947), .B(n5948), .Z(n5942) );
  AND U5296 ( .A(n2423), .B(n5941), .Z(n5948) );
  XNOR U5297 ( .A(n5949), .B(n5939), .Z(n5941) );
  XOR U5298 ( .A(n5950), .B(n5951), .Z(n5939) );
  AND U5299 ( .A(n2427), .B(n5952), .Z(n5951) );
  XOR U5300 ( .A(p_input[1991]), .B(n5950), .Z(n5952) );
  XOR U5301 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n5953), 
        .Z(n5950) );
  AND U5302 ( .A(n2430), .B(n5954), .Z(n5953) );
  IV U5303 ( .A(n5947), .Z(n5949) );
  XOR U5304 ( .A(n5955), .B(n5956), .Z(n5947) );
  AND U5305 ( .A(n2434), .B(n5957), .Z(n5956) );
  XOR U5306 ( .A(n5958), .B(n5959), .Z(n5945) );
  AND U5307 ( .A(n2438), .B(n5957), .Z(n5959) );
  XNOR U5308 ( .A(n5958), .B(n5955), .Z(n5957) );
  XNOR U5309 ( .A(n5960), .B(n5961), .Z(n5955) );
  AND U5310 ( .A(n2441), .B(n5954), .Z(n5961) );
  XNOR U5311 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n5960), 
        .Z(n5954) );
  XNOR U5312 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n5962), 
        .Z(n5960) );
  AND U5313 ( .A(n2443), .B(n5963), .Z(n5962) );
  XNOR U5314 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n5964), .Z(n5958) );
  AND U5315 ( .A(n2446), .B(n5963), .Z(n5964) );
  XOR U5316 ( .A(n5965), .B(n5966), .Z(n5963) );
  IV U5317 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n5966) );
  IV U5318 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n5965) );
  XOR U5319 ( .A(n7), .B(n5967), .Z(o[22]) );
  AND U5320 ( .A(n62), .B(n5968), .Z(n7) );
  XOR U5321 ( .A(n8), .B(n5967), .Z(n5968) );
  XOR U5322 ( .A(n5969), .B(n33), .Z(n5967) );
  AND U5323 ( .A(n65), .B(n5970), .Z(n33) );
  XNOR U5324 ( .A(n5971), .B(n34), .Z(n5970) );
  XOR U5325 ( .A(n5972), .B(n5973), .Z(n34) );
  AND U5326 ( .A(n70), .B(n5974), .Z(n5973) );
  XOR U5327 ( .A(p_input[6]), .B(n5972), .Z(n5974) );
  XOR U5328 ( .A(n5975), .B(n5976), .Z(n5972) );
  AND U5329 ( .A(n74), .B(n5977), .Z(n5976) );
  IV U5330 ( .A(n5969), .Z(n5971) );
  XOR U5331 ( .A(n5978), .B(n5979), .Z(n5969) );
  AND U5332 ( .A(n78), .B(n5980), .Z(n5979) );
  XOR U5333 ( .A(n5981), .B(n5982), .Z(n8) );
  AND U5334 ( .A(n82), .B(n5980), .Z(n5982) );
  XNOR U5335 ( .A(n5983), .B(n5978), .Z(n5980) );
  XOR U5336 ( .A(n5984), .B(n5985), .Z(n5978) );
  AND U5337 ( .A(n86), .B(n5977), .Z(n5985) );
  XNOR U5338 ( .A(n5986), .B(n5975), .Z(n5977) );
  XOR U5339 ( .A(n5987), .B(n5988), .Z(n5975) );
  AND U5340 ( .A(n90), .B(n5989), .Z(n5988) );
  XOR U5341 ( .A(p_input[22]), .B(n5987), .Z(n5989) );
  XOR U5342 ( .A(n5990), .B(n5991), .Z(n5987) );
  AND U5343 ( .A(n94), .B(n5992), .Z(n5991) );
  IV U5344 ( .A(n5984), .Z(n5986) );
  XOR U5345 ( .A(n5993), .B(n5994), .Z(n5984) );
  AND U5346 ( .A(n98), .B(n5995), .Z(n5994) );
  IV U5347 ( .A(n5981), .Z(n5983) );
  XNOR U5348 ( .A(n5996), .B(n5997), .Z(n5981) );
  AND U5349 ( .A(n102), .B(n5995), .Z(n5997) );
  XNOR U5350 ( .A(n5996), .B(n5993), .Z(n5995) );
  XOR U5351 ( .A(n5998), .B(n5999), .Z(n5993) );
  AND U5352 ( .A(n105), .B(n5992), .Z(n5999) );
  XNOR U5353 ( .A(n6000), .B(n5990), .Z(n5992) );
  XOR U5354 ( .A(n6001), .B(n6002), .Z(n5990) );
  AND U5355 ( .A(n109), .B(n6003), .Z(n6002) );
  XOR U5356 ( .A(p_input[38]), .B(n6001), .Z(n6003) );
  XOR U5357 ( .A(n6004), .B(n6005), .Z(n6001) );
  AND U5358 ( .A(n113), .B(n6006), .Z(n6005) );
  IV U5359 ( .A(n5998), .Z(n6000) );
  XOR U5360 ( .A(n6007), .B(n6008), .Z(n5998) );
  AND U5361 ( .A(n117), .B(n6009), .Z(n6008) );
  XOR U5362 ( .A(n6010), .B(n6011), .Z(n5996) );
  AND U5363 ( .A(n121), .B(n6009), .Z(n6011) );
  XNOR U5364 ( .A(n6010), .B(n6007), .Z(n6009) );
  XOR U5365 ( .A(n6012), .B(n6013), .Z(n6007) );
  AND U5366 ( .A(n124), .B(n6006), .Z(n6013) );
  XNOR U5367 ( .A(n6014), .B(n6004), .Z(n6006) );
  XOR U5368 ( .A(n6015), .B(n6016), .Z(n6004) );
  AND U5369 ( .A(n128), .B(n6017), .Z(n6016) );
  XOR U5370 ( .A(p_input[54]), .B(n6015), .Z(n6017) );
  XOR U5371 ( .A(n6018), .B(n6019), .Z(n6015) );
  AND U5372 ( .A(n132), .B(n6020), .Z(n6019) );
  IV U5373 ( .A(n6012), .Z(n6014) );
  XOR U5374 ( .A(n6021), .B(n6022), .Z(n6012) );
  AND U5375 ( .A(n136), .B(n6023), .Z(n6022) );
  XOR U5376 ( .A(n6024), .B(n6025), .Z(n6010) );
  AND U5377 ( .A(n140), .B(n6023), .Z(n6025) );
  XNOR U5378 ( .A(n6024), .B(n6021), .Z(n6023) );
  XOR U5379 ( .A(n6026), .B(n6027), .Z(n6021) );
  AND U5380 ( .A(n143), .B(n6020), .Z(n6027) );
  XNOR U5381 ( .A(n6028), .B(n6018), .Z(n6020) );
  XOR U5382 ( .A(n6029), .B(n6030), .Z(n6018) );
  AND U5383 ( .A(n147), .B(n6031), .Z(n6030) );
  XOR U5384 ( .A(p_input[70]), .B(n6029), .Z(n6031) );
  XOR U5385 ( .A(n6032), .B(n6033), .Z(n6029) );
  AND U5386 ( .A(n151), .B(n6034), .Z(n6033) );
  IV U5387 ( .A(n6026), .Z(n6028) );
  XOR U5388 ( .A(n6035), .B(n6036), .Z(n6026) );
  AND U5389 ( .A(n155), .B(n6037), .Z(n6036) );
  XOR U5390 ( .A(n6038), .B(n6039), .Z(n6024) );
  AND U5391 ( .A(n159), .B(n6037), .Z(n6039) );
  XNOR U5392 ( .A(n6038), .B(n6035), .Z(n6037) );
  XOR U5393 ( .A(n6040), .B(n6041), .Z(n6035) );
  AND U5394 ( .A(n162), .B(n6034), .Z(n6041) );
  XNOR U5395 ( .A(n6042), .B(n6032), .Z(n6034) );
  XOR U5396 ( .A(n6043), .B(n6044), .Z(n6032) );
  AND U5397 ( .A(n166), .B(n6045), .Z(n6044) );
  XOR U5398 ( .A(p_input[86]), .B(n6043), .Z(n6045) );
  XOR U5399 ( .A(n6046), .B(n6047), .Z(n6043) );
  AND U5400 ( .A(n170), .B(n6048), .Z(n6047) );
  IV U5401 ( .A(n6040), .Z(n6042) );
  XOR U5402 ( .A(n6049), .B(n6050), .Z(n6040) );
  AND U5403 ( .A(n174), .B(n6051), .Z(n6050) );
  XOR U5404 ( .A(n6052), .B(n6053), .Z(n6038) );
  AND U5405 ( .A(n178), .B(n6051), .Z(n6053) );
  XNOR U5406 ( .A(n6052), .B(n6049), .Z(n6051) );
  XOR U5407 ( .A(n6054), .B(n6055), .Z(n6049) );
  AND U5408 ( .A(n181), .B(n6048), .Z(n6055) );
  XNOR U5409 ( .A(n6056), .B(n6046), .Z(n6048) );
  XOR U5410 ( .A(n6057), .B(n6058), .Z(n6046) );
  AND U5411 ( .A(n185), .B(n6059), .Z(n6058) );
  XOR U5412 ( .A(p_input[102]), .B(n6057), .Z(n6059) );
  XOR U5413 ( .A(n6060), .B(n6061), .Z(n6057) );
  AND U5414 ( .A(n189), .B(n6062), .Z(n6061) );
  IV U5415 ( .A(n6054), .Z(n6056) );
  XOR U5416 ( .A(n6063), .B(n6064), .Z(n6054) );
  AND U5417 ( .A(n193), .B(n6065), .Z(n6064) );
  XOR U5418 ( .A(n6066), .B(n6067), .Z(n6052) );
  AND U5419 ( .A(n197), .B(n6065), .Z(n6067) );
  XNOR U5420 ( .A(n6066), .B(n6063), .Z(n6065) );
  XOR U5421 ( .A(n6068), .B(n6069), .Z(n6063) );
  AND U5422 ( .A(n200), .B(n6062), .Z(n6069) );
  XNOR U5423 ( .A(n6070), .B(n6060), .Z(n6062) );
  XOR U5424 ( .A(n6071), .B(n6072), .Z(n6060) );
  AND U5425 ( .A(n204), .B(n6073), .Z(n6072) );
  XOR U5426 ( .A(p_input[118]), .B(n6071), .Z(n6073) );
  XOR U5427 ( .A(n6074), .B(n6075), .Z(n6071) );
  AND U5428 ( .A(n208), .B(n6076), .Z(n6075) );
  IV U5429 ( .A(n6068), .Z(n6070) );
  XOR U5430 ( .A(n6077), .B(n6078), .Z(n6068) );
  AND U5431 ( .A(n212), .B(n6079), .Z(n6078) );
  XOR U5432 ( .A(n6080), .B(n6081), .Z(n6066) );
  AND U5433 ( .A(n216), .B(n6079), .Z(n6081) );
  XNOR U5434 ( .A(n6080), .B(n6077), .Z(n6079) );
  XOR U5435 ( .A(n6082), .B(n6083), .Z(n6077) );
  AND U5436 ( .A(n219), .B(n6076), .Z(n6083) );
  XNOR U5437 ( .A(n6084), .B(n6074), .Z(n6076) );
  XOR U5438 ( .A(n6085), .B(n6086), .Z(n6074) );
  AND U5439 ( .A(n223), .B(n6087), .Z(n6086) );
  XOR U5440 ( .A(p_input[134]), .B(n6085), .Z(n6087) );
  XOR U5441 ( .A(n6088), .B(n6089), .Z(n6085) );
  AND U5442 ( .A(n227), .B(n6090), .Z(n6089) );
  IV U5443 ( .A(n6082), .Z(n6084) );
  XOR U5444 ( .A(n6091), .B(n6092), .Z(n6082) );
  AND U5445 ( .A(n231), .B(n6093), .Z(n6092) );
  XOR U5446 ( .A(n6094), .B(n6095), .Z(n6080) );
  AND U5447 ( .A(n235), .B(n6093), .Z(n6095) );
  XNOR U5448 ( .A(n6094), .B(n6091), .Z(n6093) );
  XOR U5449 ( .A(n6096), .B(n6097), .Z(n6091) );
  AND U5450 ( .A(n238), .B(n6090), .Z(n6097) );
  XNOR U5451 ( .A(n6098), .B(n6088), .Z(n6090) );
  XOR U5452 ( .A(n6099), .B(n6100), .Z(n6088) );
  AND U5453 ( .A(n242), .B(n6101), .Z(n6100) );
  XOR U5454 ( .A(p_input[150]), .B(n6099), .Z(n6101) );
  XOR U5455 ( .A(n6102), .B(n6103), .Z(n6099) );
  AND U5456 ( .A(n246), .B(n6104), .Z(n6103) );
  IV U5457 ( .A(n6096), .Z(n6098) );
  XOR U5458 ( .A(n6105), .B(n6106), .Z(n6096) );
  AND U5459 ( .A(n250), .B(n6107), .Z(n6106) );
  XOR U5460 ( .A(n6108), .B(n6109), .Z(n6094) );
  AND U5461 ( .A(n254), .B(n6107), .Z(n6109) );
  XNOR U5462 ( .A(n6108), .B(n6105), .Z(n6107) );
  XOR U5463 ( .A(n6110), .B(n6111), .Z(n6105) );
  AND U5464 ( .A(n257), .B(n6104), .Z(n6111) );
  XNOR U5465 ( .A(n6112), .B(n6102), .Z(n6104) );
  XOR U5466 ( .A(n6113), .B(n6114), .Z(n6102) );
  AND U5467 ( .A(n261), .B(n6115), .Z(n6114) );
  XOR U5468 ( .A(p_input[166]), .B(n6113), .Z(n6115) );
  XOR U5469 ( .A(n6116), .B(n6117), .Z(n6113) );
  AND U5470 ( .A(n265), .B(n6118), .Z(n6117) );
  IV U5471 ( .A(n6110), .Z(n6112) );
  XOR U5472 ( .A(n6119), .B(n6120), .Z(n6110) );
  AND U5473 ( .A(n269), .B(n6121), .Z(n6120) );
  XOR U5474 ( .A(n6122), .B(n6123), .Z(n6108) );
  AND U5475 ( .A(n273), .B(n6121), .Z(n6123) );
  XNOR U5476 ( .A(n6122), .B(n6119), .Z(n6121) );
  XOR U5477 ( .A(n6124), .B(n6125), .Z(n6119) );
  AND U5478 ( .A(n276), .B(n6118), .Z(n6125) );
  XNOR U5479 ( .A(n6126), .B(n6116), .Z(n6118) );
  XOR U5480 ( .A(n6127), .B(n6128), .Z(n6116) );
  AND U5481 ( .A(n280), .B(n6129), .Z(n6128) );
  XOR U5482 ( .A(p_input[182]), .B(n6127), .Z(n6129) );
  XOR U5483 ( .A(n6130), .B(n6131), .Z(n6127) );
  AND U5484 ( .A(n284), .B(n6132), .Z(n6131) );
  IV U5485 ( .A(n6124), .Z(n6126) );
  XOR U5486 ( .A(n6133), .B(n6134), .Z(n6124) );
  AND U5487 ( .A(n288), .B(n6135), .Z(n6134) );
  XOR U5488 ( .A(n6136), .B(n6137), .Z(n6122) );
  AND U5489 ( .A(n292), .B(n6135), .Z(n6137) );
  XNOR U5490 ( .A(n6136), .B(n6133), .Z(n6135) );
  XOR U5491 ( .A(n6138), .B(n6139), .Z(n6133) );
  AND U5492 ( .A(n295), .B(n6132), .Z(n6139) );
  XNOR U5493 ( .A(n6140), .B(n6130), .Z(n6132) );
  XOR U5494 ( .A(n6141), .B(n6142), .Z(n6130) );
  AND U5495 ( .A(n299), .B(n6143), .Z(n6142) );
  XOR U5496 ( .A(p_input[198]), .B(n6141), .Z(n6143) );
  XOR U5497 ( .A(n6144), .B(n6145), .Z(n6141) );
  AND U5498 ( .A(n303), .B(n6146), .Z(n6145) );
  IV U5499 ( .A(n6138), .Z(n6140) );
  XOR U5500 ( .A(n6147), .B(n6148), .Z(n6138) );
  AND U5501 ( .A(n307), .B(n6149), .Z(n6148) );
  XOR U5502 ( .A(n6150), .B(n6151), .Z(n6136) );
  AND U5503 ( .A(n311), .B(n6149), .Z(n6151) );
  XNOR U5504 ( .A(n6150), .B(n6147), .Z(n6149) );
  XOR U5505 ( .A(n6152), .B(n6153), .Z(n6147) );
  AND U5506 ( .A(n314), .B(n6146), .Z(n6153) );
  XNOR U5507 ( .A(n6154), .B(n6144), .Z(n6146) );
  XOR U5508 ( .A(n6155), .B(n6156), .Z(n6144) );
  AND U5509 ( .A(n318), .B(n6157), .Z(n6156) );
  XOR U5510 ( .A(p_input[214]), .B(n6155), .Z(n6157) );
  XOR U5511 ( .A(n6158), .B(n6159), .Z(n6155) );
  AND U5512 ( .A(n322), .B(n6160), .Z(n6159) );
  IV U5513 ( .A(n6152), .Z(n6154) );
  XOR U5514 ( .A(n6161), .B(n6162), .Z(n6152) );
  AND U5515 ( .A(n326), .B(n6163), .Z(n6162) );
  XOR U5516 ( .A(n6164), .B(n6165), .Z(n6150) );
  AND U5517 ( .A(n330), .B(n6163), .Z(n6165) );
  XNOR U5518 ( .A(n6164), .B(n6161), .Z(n6163) );
  XOR U5519 ( .A(n6166), .B(n6167), .Z(n6161) );
  AND U5520 ( .A(n333), .B(n6160), .Z(n6167) );
  XNOR U5521 ( .A(n6168), .B(n6158), .Z(n6160) );
  XOR U5522 ( .A(n6169), .B(n6170), .Z(n6158) );
  AND U5523 ( .A(n337), .B(n6171), .Z(n6170) );
  XOR U5524 ( .A(p_input[230]), .B(n6169), .Z(n6171) );
  XOR U5525 ( .A(n6172), .B(n6173), .Z(n6169) );
  AND U5526 ( .A(n341), .B(n6174), .Z(n6173) );
  IV U5527 ( .A(n6166), .Z(n6168) );
  XOR U5528 ( .A(n6175), .B(n6176), .Z(n6166) );
  AND U5529 ( .A(n345), .B(n6177), .Z(n6176) );
  XOR U5530 ( .A(n6178), .B(n6179), .Z(n6164) );
  AND U5531 ( .A(n349), .B(n6177), .Z(n6179) );
  XNOR U5532 ( .A(n6178), .B(n6175), .Z(n6177) );
  XOR U5533 ( .A(n6180), .B(n6181), .Z(n6175) );
  AND U5534 ( .A(n352), .B(n6174), .Z(n6181) );
  XNOR U5535 ( .A(n6182), .B(n6172), .Z(n6174) );
  XOR U5536 ( .A(n6183), .B(n6184), .Z(n6172) );
  AND U5537 ( .A(n356), .B(n6185), .Z(n6184) );
  XOR U5538 ( .A(p_input[246]), .B(n6183), .Z(n6185) );
  XOR U5539 ( .A(n6186), .B(n6187), .Z(n6183) );
  AND U5540 ( .A(n360), .B(n6188), .Z(n6187) );
  IV U5541 ( .A(n6180), .Z(n6182) );
  XOR U5542 ( .A(n6189), .B(n6190), .Z(n6180) );
  AND U5543 ( .A(n364), .B(n6191), .Z(n6190) );
  XOR U5544 ( .A(n6192), .B(n6193), .Z(n6178) );
  AND U5545 ( .A(n368), .B(n6191), .Z(n6193) );
  XNOR U5546 ( .A(n6192), .B(n6189), .Z(n6191) );
  XOR U5547 ( .A(n6194), .B(n6195), .Z(n6189) );
  AND U5548 ( .A(n371), .B(n6188), .Z(n6195) );
  XNOR U5549 ( .A(n6196), .B(n6186), .Z(n6188) );
  XOR U5550 ( .A(n6197), .B(n6198), .Z(n6186) );
  AND U5551 ( .A(n375), .B(n6199), .Z(n6198) );
  XOR U5552 ( .A(p_input[262]), .B(n6197), .Z(n6199) );
  XOR U5553 ( .A(n6200), .B(n6201), .Z(n6197) );
  AND U5554 ( .A(n379), .B(n6202), .Z(n6201) );
  IV U5555 ( .A(n6194), .Z(n6196) );
  XOR U5556 ( .A(n6203), .B(n6204), .Z(n6194) );
  AND U5557 ( .A(n383), .B(n6205), .Z(n6204) );
  XOR U5558 ( .A(n6206), .B(n6207), .Z(n6192) );
  AND U5559 ( .A(n387), .B(n6205), .Z(n6207) );
  XNOR U5560 ( .A(n6206), .B(n6203), .Z(n6205) );
  XOR U5561 ( .A(n6208), .B(n6209), .Z(n6203) );
  AND U5562 ( .A(n390), .B(n6202), .Z(n6209) );
  XNOR U5563 ( .A(n6210), .B(n6200), .Z(n6202) );
  XOR U5564 ( .A(n6211), .B(n6212), .Z(n6200) );
  AND U5565 ( .A(n394), .B(n6213), .Z(n6212) );
  XOR U5566 ( .A(p_input[278]), .B(n6211), .Z(n6213) );
  XOR U5567 ( .A(n6214), .B(n6215), .Z(n6211) );
  AND U5568 ( .A(n398), .B(n6216), .Z(n6215) );
  IV U5569 ( .A(n6208), .Z(n6210) );
  XOR U5570 ( .A(n6217), .B(n6218), .Z(n6208) );
  AND U5571 ( .A(n402), .B(n6219), .Z(n6218) );
  XOR U5572 ( .A(n6220), .B(n6221), .Z(n6206) );
  AND U5573 ( .A(n406), .B(n6219), .Z(n6221) );
  XNOR U5574 ( .A(n6220), .B(n6217), .Z(n6219) );
  XOR U5575 ( .A(n6222), .B(n6223), .Z(n6217) );
  AND U5576 ( .A(n409), .B(n6216), .Z(n6223) );
  XNOR U5577 ( .A(n6224), .B(n6214), .Z(n6216) );
  XOR U5578 ( .A(n6225), .B(n6226), .Z(n6214) );
  AND U5579 ( .A(n413), .B(n6227), .Z(n6226) );
  XOR U5580 ( .A(p_input[294]), .B(n6225), .Z(n6227) );
  XOR U5581 ( .A(n6228), .B(n6229), .Z(n6225) );
  AND U5582 ( .A(n417), .B(n6230), .Z(n6229) );
  IV U5583 ( .A(n6222), .Z(n6224) );
  XOR U5584 ( .A(n6231), .B(n6232), .Z(n6222) );
  AND U5585 ( .A(n421), .B(n6233), .Z(n6232) );
  XOR U5586 ( .A(n6234), .B(n6235), .Z(n6220) );
  AND U5587 ( .A(n425), .B(n6233), .Z(n6235) );
  XNOR U5588 ( .A(n6234), .B(n6231), .Z(n6233) );
  XOR U5589 ( .A(n6236), .B(n6237), .Z(n6231) );
  AND U5590 ( .A(n428), .B(n6230), .Z(n6237) );
  XNOR U5591 ( .A(n6238), .B(n6228), .Z(n6230) );
  XOR U5592 ( .A(n6239), .B(n6240), .Z(n6228) );
  AND U5593 ( .A(n432), .B(n6241), .Z(n6240) );
  XOR U5594 ( .A(p_input[310]), .B(n6239), .Z(n6241) );
  XOR U5595 ( .A(n6242), .B(n6243), .Z(n6239) );
  AND U5596 ( .A(n436), .B(n6244), .Z(n6243) );
  IV U5597 ( .A(n6236), .Z(n6238) );
  XOR U5598 ( .A(n6245), .B(n6246), .Z(n6236) );
  AND U5599 ( .A(n440), .B(n6247), .Z(n6246) );
  XOR U5600 ( .A(n6248), .B(n6249), .Z(n6234) );
  AND U5601 ( .A(n444), .B(n6247), .Z(n6249) );
  XNOR U5602 ( .A(n6248), .B(n6245), .Z(n6247) );
  XOR U5603 ( .A(n6250), .B(n6251), .Z(n6245) );
  AND U5604 ( .A(n447), .B(n6244), .Z(n6251) );
  XNOR U5605 ( .A(n6252), .B(n6242), .Z(n6244) );
  XOR U5606 ( .A(n6253), .B(n6254), .Z(n6242) );
  AND U5607 ( .A(n451), .B(n6255), .Z(n6254) );
  XOR U5608 ( .A(p_input[326]), .B(n6253), .Z(n6255) );
  XOR U5609 ( .A(n6256), .B(n6257), .Z(n6253) );
  AND U5610 ( .A(n455), .B(n6258), .Z(n6257) );
  IV U5611 ( .A(n6250), .Z(n6252) );
  XOR U5612 ( .A(n6259), .B(n6260), .Z(n6250) );
  AND U5613 ( .A(n459), .B(n6261), .Z(n6260) );
  XOR U5614 ( .A(n6262), .B(n6263), .Z(n6248) );
  AND U5615 ( .A(n463), .B(n6261), .Z(n6263) );
  XNOR U5616 ( .A(n6262), .B(n6259), .Z(n6261) );
  XOR U5617 ( .A(n6264), .B(n6265), .Z(n6259) );
  AND U5618 ( .A(n466), .B(n6258), .Z(n6265) );
  XNOR U5619 ( .A(n6266), .B(n6256), .Z(n6258) );
  XOR U5620 ( .A(n6267), .B(n6268), .Z(n6256) );
  AND U5621 ( .A(n470), .B(n6269), .Z(n6268) );
  XOR U5622 ( .A(p_input[342]), .B(n6267), .Z(n6269) );
  XOR U5623 ( .A(n6270), .B(n6271), .Z(n6267) );
  AND U5624 ( .A(n474), .B(n6272), .Z(n6271) );
  IV U5625 ( .A(n6264), .Z(n6266) );
  XOR U5626 ( .A(n6273), .B(n6274), .Z(n6264) );
  AND U5627 ( .A(n478), .B(n6275), .Z(n6274) );
  XOR U5628 ( .A(n6276), .B(n6277), .Z(n6262) );
  AND U5629 ( .A(n482), .B(n6275), .Z(n6277) );
  XNOR U5630 ( .A(n6276), .B(n6273), .Z(n6275) );
  XOR U5631 ( .A(n6278), .B(n6279), .Z(n6273) );
  AND U5632 ( .A(n485), .B(n6272), .Z(n6279) );
  XNOR U5633 ( .A(n6280), .B(n6270), .Z(n6272) );
  XOR U5634 ( .A(n6281), .B(n6282), .Z(n6270) );
  AND U5635 ( .A(n489), .B(n6283), .Z(n6282) );
  XOR U5636 ( .A(p_input[358]), .B(n6281), .Z(n6283) );
  XOR U5637 ( .A(n6284), .B(n6285), .Z(n6281) );
  AND U5638 ( .A(n493), .B(n6286), .Z(n6285) );
  IV U5639 ( .A(n6278), .Z(n6280) );
  XOR U5640 ( .A(n6287), .B(n6288), .Z(n6278) );
  AND U5641 ( .A(n497), .B(n6289), .Z(n6288) );
  XOR U5642 ( .A(n6290), .B(n6291), .Z(n6276) );
  AND U5643 ( .A(n501), .B(n6289), .Z(n6291) );
  XNOR U5644 ( .A(n6290), .B(n6287), .Z(n6289) );
  XOR U5645 ( .A(n6292), .B(n6293), .Z(n6287) );
  AND U5646 ( .A(n504), .B(n6286), .Z(n6293) );
  XNOR U5647 ( .A(n6294), .B(n6284), .Z(n6286) );
  XOR U5648 ( .A(n6295), .B(n6296), .Z(n6284) );
  AND U5649 ( .A(n508), .B(n6297), .Z(n6296) );
  XOR U5650 ( .A(p_input[374]), .B(n6295), .Z(n6297) );
  XOR U5651 ( .A(n6298), .B(n6299), .Z(n6295) );
  AND U5652 ( .A(n512), .B(n6300), .Z(n6299) );
  IV U5653 ( .A(n6292), .Z(n6294) );
  XOR U5654 ( .A(n6301), .B(n6302), .Z(n6292) );
  AND U5655 ( .A(n516), .B(n6303), .Z(n6302) );
  XOR U5656 ( .A(n6304), .B(n6305), .Z(n6290) );
  AND U5657 ( .A(n520), .B(n6303), .Z(n6305) );
  XNOR U5658 ( .A(n6304), .B(n6301), .Z(n6303) );
  XOR U5659 ( .A(n6306), .B(n6307), .Z(n6301) );
  AND U5660 ( .A(n523), .B(n6300), .Z(n6307) );
  XNOR U5661 ( .A(n6308), .B(n6298), .Z(n6300) );
  XOR U5662 ( .A(n6309), .B(n6310), .Z(n6298) );
  AND U5663 ( .A(n527), .B(n6311), .Z(n6310) );
  XOR U5664 ( .A(p_input[390]), .B(n6309), .Z(n6311) );
  XOR U5665 ( .A(n6312), .B(n6313), .Z(n6309) );
  AND U5666 ( .A(n531), .B(n6314), .Z(n6313) );
  IV U5667 ( .A(n6306), .Z(n6308) );
  XOR U5668 ( .A(n6315), .B(n6316), .Z(n6306) );
  AND U5669 ( .A(n535), .B(n6317), .Z(n6316) );
  XOR U5670 ( .A(n6318), .B(n6319), .Z(n6304) );
  AND U5671 ( .A(n539), .B(n6317), .Z(n6319) );
  XNOR U5672 ( .A(n6318), .B(n6315), .Z(n6317) );
  XOR U5673 ( .A(n6320), .B(n6321), .Z(n6315) );
  AND U5674 ( .A(n542), .B(n6314), .Z(n6321) );
  XNOR U5675 ( .A(n6322), .B(n6312), .Z(n6314) );
  XOR U5676 ( .A(n6323), .B(n6324), .Z(n6312) );
  AND U5677 ( .A(n546), .B(n6325), .Z(n6324) );
  XOR U5678 ( .A(p_input[406]), .B(n6323), .Z(n6325) );
  XOR U5679 ( .A(n6326), .B(n6327), .Z(n6323) );
  AND U5680 ( .A(n550), .B(n6328), .Z(n6327) );
  IV U5681 ( .A(n6320), .Z(n6322) );
  XOR U5682 ( .A(n6329), .B(n6330), .Z(n6320) );
  AND U5683 ( .A(n554), .B(n6331), .Z(n6330) );
  XOR U5684 ( .A(n6332), .B(n6333), .Z(n6318) );
  AND U5685 ( .A(n558), .B(n6331), .Z(n6333) );
  XNOR U5686 ( .A(n6332), .B(n6329), .Z(n6331) );
  XOR U5687 ( .A(n6334), .B(n6335), .Z(n6329) );
  AND U5688 ( .A(n561), .B(n6328), .Z(n6335) );
  XNOR U5689 ( .A(n6336), .B(n6326), .Z(n6328) );
  XOR U5690 ( .A(n6337), .B(n6338), .Z(n6326) );
  AND U5691 ( .A(n565), .B(n6339), .Z(n6338) );
  XOR U5692 ( .A(p_input[422]), .B(n6337), .Z(n6339) );
  XOR U5693 ( .A(n6340), .B(n6341), .Z(n6337) );
  AND U5694 ( .A(n569), .B(n6342), .Z(n6341) );
  IV U5695 ( .A(n6334), .Z(n6336) );
  XOR U5696 ( .A(n6343), .B(n6344), .Z(n6334) );
  AND U5697 ( .A(n573), .B(n6345), .Z(n6344) );
  XOR U5698 ( .A(n6346), .B(n6347), .Z(n6332) );
  AND U5699 ( .A(n577), .B(n6345), .Z(n6347) );
  XNOR U5700 ( .A(n6346), .B(n6343), .Z(n6345) );
  XOR U5701 ( .A(n6348), .B(n6349), .Z(n6343) );
  AND U5702 ( .A(n580), .B(n6342), .Z(n6349) );
  XNOR U5703 ( .A(n6350), .B(n6340), .Z(n6342) );
  XOR U5704 ( .A(n6351), .B(n6352), .Z(n6340) );
  AND U5705 ( .A(n584), .B(n6353), .Z(n6352) );
  XOR U5706 ( .A(p_input[438]), .B(n6351), .Z(n6353) );
  XOR U5707 ( .A(n6354), .B(n6355), .Z(n6351) );
  AND U5708 ( .A(n588), .B(n6356), .Z(n6355) );
  IV U5709 ( .A(n6348), .Z(n6350) );
  XOR U5710 ( .A(n6357), .B(n6358), .Z(n6348) );
  AND U5711 ( .A(n592), .B(n6359), .Z(n6358) );
  XOR U5712 ( .A(n6360), .B(n6361), .Z(n6346) );
  AND U5713 ( .A(n596), .B(n6359), .Z(n6361) );
  XNOR U5714 ( .A(n6360), .B(n6357), .Z(n6359) );
  XOR U5715 ( .A(n6362), .B(n6363), .Z(n6357) );
  AND U5716 ( .A(n599), .B(n6356), .Z(n6363) );
  XNOR U5717 ( .A(n6364), .B(n6354), .Z(n6356) );
  XOR U5718 ( .A(n6365), .B(n6366), .Z(n6354) );
  AND U5719 ( .A(n603), .B(n6367), .Z(n6366) );
  XOR U5720 ( .A(p_input[454]), .B(n6365), .Z(n6367) );
  XOR U5721 ( .A(n6368), .B(n6369), .Z(n6365) );
  AND U5722 ( .A(n607), .B(n6370), .Z(n6369) );
  IV U5723 ( .A(n6362), .Z(n6364) );
  XOR U5724 ( .A(n6371), .B(n6372), .Z(n6362) );
  AND U5725 ( .A(n611), .B(n6373), .Z(n6372) );
  XOR U5726 ( .A(n6374), .B(n6375), .Z(n6360) );
  AND U5727 ( .A(n615), .B(n6373), .Z(n6375) );
  XNOR U5728 ( .A(n6374), .B(n6371), .Z(n6373) );
  XOR U5729 ( .A(n6376), .B(n6377), .Z(n6371) );
  AND U5730 ( .A(n618), .B(n6370), .Z(n6377) );
  XNOR U5731 ( .A(n6378), .B(n6368), .Z(n6370) );
  XOR U5732 ( .A(n6379), .B(n6380), .Z(n6368) );
  AND U5733 ( .A(n622), .B(n6381), .Z(n6380) );
  XOR U5734 ( .A(p_input[470]), .B(n6379), .Z(n6381) );
  XOR U5735 ( .A(n6382), .B(n6383), .Z(n6379) );
  AND U5736 ( .A(n626), .B(n6384), .Z(n6383) );
  IV U5737 ( .A(n6376), .Z(n6378) );
  XOR U5738 ( .A(n6385), .B(n6386), .Z(n6376) );
  AND U5739 ( .A(n630), .B(n6387), .Z(n6386) );
  XOR U5740 ( .A(n6388), .B(n6389), .Z(n6374) );
  AND U5741 ( .A(n634), .B(n6387), .Z(n6389) );
  XNOR U5742 ( .A(n6388), .B(n6385), .Z(n6387) );
  XOR U5743 ( .A(n6390), .B(n6391), .Z(n6385) );
  AND U5744 ( .A(n637), .B(n6384), .Z(n6391) );
  XNOR U5745 ( .A(n6392), .B(n6382), .Z(n6384) );
  XOR U5746 ( .A(n6393), .B(n6394), .Z(n6382) );
  AND U5747 ( .A(n641), .B(n6395), .Z(n6394) );
  XOR U5748 ( .A(p_input[486]), .B(n6393), .Z(n6395) );
  XOR U5749 ( .A(n6396), .B(n6397), .Z(n6393) );
  AND U5750 ( .A(n645), .B(n6398), .Z(n6397) );
  IV U5751 ( .A(n6390), .Z(n6392) );
  XOR U5752 ( .A(n6399), .B(n6400), .Z(n6390) );
  AND U5753 ( .A(n649), .B(n6401), .Z(n6400) );
  XOR U5754 ( .A(n6402), .B(n6403), .Z(n6388) );
  AND U5755 ( .A(n653), .B(n6401), .Z(n6403) );
  XNOR U5756 ( .A(n6402), .B(n6399), .Z(n6401) );
  XOR U5757 ( .A(n6404), .B(n6405), .Z(n6399) );
  AND U5758 ( .A(n656), .B(n6398), .Z(n6405) );
  XNOR U5759 ( .A(n6406), .B(n6396), .Z(n6398) );
  XOR U5760 ( .A(n6407), .B(n6408), .Z(n6396) );
  AND U5761 ( .A(n660), .B(n6409), .Z(n6408) );
  XOR U5762 ( .A(p_input[502]), .B(n6407), .Z(n6409) );
  XOR U5763 ( .A(n6410), .B(n6411), .Z(n6407) );
  AND U5764 ( .A(n664), .B(n6412), .Z(n6411) );
  IV U5765 ( .A(n6404), .Z(n6406) );
  XOR U5766 ( .A(n6413), .B(n6414), .Z(n6404) );
  AND U5767 ( .A(n668), .B(n6415), .Z(n6414) );
  XOR U5768 ( .A(n6416), .B(n6417), .Z(n6402) );
  AND U5769 ( .A(n672), .B(n6415), .Z(n6417) );
  XNOR U5770 ( .A(n6416), .B(n6413), .Z(n6415) );
  XOR U5771 ( .A(n6418), .B(n6419), .Z(n6413) );
  AND U5772 ( .A(n675), .B(n6412), .Z(n6419) );
  XNOR U5773 ( .A(n6420), .B(n6410), .Z(n6412) );
  XOR U5774 ( .A(n6421), .B(n6422), .Z(n6410) );
  AND U5775 ( .A(n679), .B(n6423), .Z(n6422) );
  XOR U5776 ( .A(p_input[518]), .B(n6421), .Z(n6423) );
  XOR U5777 ( .A(n6424), .B(n6425), .Z(n6421) );
  AND U5778 ( .A(n683), .B(n6426), .Z(n6425) );
  IV U5779 ( .A(n6418), .Z(n6420) );
  XOR U5780 ( .A(n6427), .B(n6428), .Z(n6418) );
  AND U5781 ( .A(n687), .B(n6429), .Z(n6428) );
  XOR U5782 ( .A(n6430), .B(n6431), .Z(n6416) );
  AND U5783 ( .A(n691), .B(n6429), .Z(n6431) );
  XNOR U5784 ( .A(n6430), .B(n6427), .Z(n6429) );
  XOR U5785 ( .A(n6432), .B(n6433), .Z(n6427) );
  AND U5786 ( .A(n694), .B(n6426), .Z(n6433) );
  XNOR U5787 ( .A(n6434), .B(n6424), .Z(n6426) );
  XOR U5788 ( .A(n6435), .B(n6436), .Z(n6424) );
  AND U5789 ( .A(n698), .B(n6437), .Z(n6436) );
  XOR U5790 ( .A(p_input[534]), .B(n6435), .Z(n6437) );
  XOR U5791 ( .A(n6438), .B(n6439), .Z(n6435) );
  AND U5792 ( .A(n702), .B(n6440), .Z(n6439) );
  IV U5793 ( .A(n6432), .Z(n6434) );
  XOR U5794 ( .A(n6441), .B(n6442), .Z(n6432) );
  AND U5795 ( .A(n706), .B(n6443), .Z(n6442) );
  XOR U5796 ( .A(n6444), .B(n6445), .Z(n6430) );
  AND U5797 ( .A(n710), .B(n6443), .Z(n6445) );
  XNOR U5798 ( .A(n6444), .B(n6441), .Z(n6443) );
  XOR U5799 ( .A(n6446), .B(n6447), .Z(n6441) );
  AND U5800 ( .A(n713), .B(n6440), .Z(n6447) );
  XNOR U5801 ( .A(n6448), .B(n6438), .Z(n6440) );
  XOR U5802 ( .A(n6449), .B(n6450), .Z(n6438) );
  AND U5803 ( .A(n717), .B(n6451), .Z(n6450) );
  XOR U5804 ( .A(p_input[550]), .B(n6449), .Z(n6451) );
  XOR U5805 ( .A(n6452), .B(n6453), .Z(n6449) );
  AND U5806 ( .A(n721), .B(n6454), .Z(n6453) );
  IV U5807 ( .A(n6446), .Z(n6448) );
  XOR U5808 ( .A(n6455), .B(n6456), .Z(n6446) );
  AND U5809 ( .A(n725), .B(n6457), .Z(n6456) );
  XOR U5810 ( .A(n6458), .B(n6459), .Z(n6444) );
  AND U5811 ( .A(n729), .B(n6457), .Z(n6459) );
  XNOR U5812 ( .A(n6458), .B(n6455), .Z(n6457) );
  XOR U5813 ( .A(n6460), .B(n6461), .Z(n6455) );
  AND U5814 ( .A(n732), .B(n6454), .Z(n6461) );
  XNOR U5815 ( .A(n6462), .B(n6452), .Z(n6454) );
  XOR U5816 ( .A(n6463), .B(n6464), .Z(n6452) );
  AND U5817 ( .A(n736), .B(n6465), .Z(n6464) );
  XOR U5818 ( .A(p_input[566]), .B(n6463), .Z(n6465) );
  XOR U5819 ( .A(n6466), .B(n6467), .Z(n6463) );
  AND U5820 ( .A(n740), .B(n6468), .Z(n6467) );
  IV U5821 ( .A(n6460), .Z(n6462) );
  XOR U5822 ( .A(n6469), .B(n6470), .Z(n6460) );
  AND U5823 ( .A(n744), .B(n6471), .Z(n6470) );
  XOR U5824 ( .A(n6472), .B(n6473), .Z(n6458) );
  AND U5825 ( .A(n748), .B(n6471), .Z(n6473) );
  XNOR U5826 ( .A(n6472), .B(n6469), .Z(n6471) );
  XOR U5827 ( .A(n6474), .B(n6475), .Z(n6469) );
  AND U5828 ( .A(n751), .B(n6468), .Z(n6475) );
  XNOR U5829 ( .A(n6476), .B(n6466), .Z(n6468) );
  XOR U5830 ( .A(n6477), .B(n6478), .Z(n6466) );
  AND U5831 ( .A(n755), .B(n6479), .Z(n6478) );
  XOR U5832 ( .A(p_input[582]), .B(n6477), .Z(n6479) );
  XOR U5833 ( .A(n6480), .B(n6481), .Z(n6477) );
  AND U5834 ( .A(n759), .B(n6482), .Z(n6481) );
  IV U5835 ( .A(n6474), .Z(n6476) );
  XOR U5836 ( .A(n6483), .B(n6484), .Z(n6474) );
  AND U5837 ( .A(n763), .B(n6485), .Z(n6484) );
  XOR U5838 ( .A(n6486), .B(n6487), .Z(n6472) );
  AND U5839 ( .A(n767), .B(n6485), .Z(n6487) );
  XNOR U5840 ( .A(n6486), .B(n6483), .Z(n6485) );
  XOR U5841 ( .A(n6488), .B(n6489), .Z(n6483) );
  AND U5842 ( .A(n770), .B(n6482), .Z(n6489) );
  XNOR U5843 ( .A(n6490), .B(n6480), .Z(n6482) );
  XOR U5844 ( .A(n6491), .B(n6492), .Z(n6480) );
  AND U5845 ( .A(n774), .B(n6493), .Z(n6492) );
  XOR U5846 ( .A(p_input[598]), .B(n6491), .Z(n6493) );
  XOR U5847 ( .A(n6494), .B(n6495), .Z(n6491) );
  AND U5848 ( .A(n778), .B(n6496), .Z(n6495) );
  IV U5849 ( .A(n6488), .Z(n6490) );
  XOR U5850 ( .A(n6497), .B(n6498), .Z(n6488) );
  AND U5851 ( .A(n782), .B(n6499), .Z(n6498) );
  XOR U5852 ( .A(n6500), .B(n6501), .Z(n6486) );
  AND U5853 ( .A(n786), .B(n6499), .Z(n6501) );
  XNOR U5854 ( .A(n6500), .B(n6497), .Z(n6499) );
  XOR U5855 ( .A(n6502), .B(n6503), .Z(n6497) );
  AND U5856 ( .A(n789), .B(n6496), .Z(n6503) );
  XNOR U5857 ( .A(n6504), .B(n6494), .Z(n6496) );
  XOR U5858 ( .A(n6505), .B(n6506), .Z(n6494) );
  AND U5859 ( .A(n793), .B(n6507), .Z(n6506) );
  XOR U5860 ( .A(p_input[614]), .B(n6505), .Z(n6507) );
  XOR U5861 ( .A(n6508), .B(n6509), .Z(n6505) );
  AND U5862 ( .A(n797), .B(n6510), .Z(n6509) );
  IV U5863 ( .A(n6502), .Z(n6504) );
  XOR U5864 ( .A(n6511), .B(n6512), .Z(n6502) );
  AND U5865 ( .A(n801), .B(n6513), .Z(n6512) );
  XOR U5866 ( .A(n6514), .B(n6515), .Z(n6500) );
  AND U5867 ( .A(n805), .B(n6513), .Z(n6515) );
  XNOR U5868 ( .A(n6514), .B(n6511), .Z(n6513) );
  XOR U5869 ( .A(n6516), .B(n6517), .Z(n6511) );
  AND U5870 ( .A(n808), .B(n6510), .Z(n6517) );
  XNOR U5871 ( .A(n6518), .B(n6508), .Z(n6510) );
  XOR U5872 ( .A(n6519), .B(n6520), .Z(n6508) );
  AND U5873 ( .A(n812), .B(n6521), .Z(n6520) );
  XOR U5874 ( .A(p_input[630]), .B(n6519), .Z(n6521) );
  XOR U5875 ( .A(n6522), .B(n6523), .Z(n6519) );
  AND U5876 ( .A(n816), .B(n6524), .Z(n6523) );
  IV U5877 ( .A(n6516), .Z(n6518) );
  XOR U5878 ( .A(n6525), .B(n6526), .Z(n6516) );
  AND U5879 ( .A(n820), .B(n6527), .Z(n6526) );
  XOR U5880 ( .A(n6528), .B(n6529), .Z(n6514) );
  AND U5881 ( .A(n824), .B(n6527), .Z(n6529) );
  XNOR U5882 ( .A(n6528), .B(n6525), .Z(n6527) );
  XOR U5883 ( .A(n6530), .B(n6531), .Z(n6525) );
  AND U5884 ( .A(n827), .B(n6524), .Z(n6531) );
  XNOR U5885 ( .A(n6532), .B(n6522), .Z(n6524) );
  XOR U5886 ( .A(n6533), .B(n6534), .Z(n6522) );
  AND U5887 ( .A(n831), .B(n6535), .Z(n6534) );
  XOR U5888 ( .A(p_input[646]), .B(n6533), .Z(n6535) );
  XOR U5889 ( .A(n6536), .B(n6537), .Z(n6533) );
  AND U5890 ( .A(n835), .B(n6538), .Z(n6537) );
  IV U5891 ( .A(n6530), .Z(n6532) );
  XOR U5892 ( .A(n6539), .B(n6540), .Z(n6530) );
  AND U5893 ( .A(n839), .B(n6541), .Z(n6540) );
  XOR U5894 ( .A(n6542), .B(n6543), .Z(n6528) );
  AND U5895 ( .A(n843), .B(n6541), .Z(n6543) );
  XNOR U5896 ( .A(n6542), .B(n6539), .Z(n6541) );
  XOR U5897 ( .A(n6544), .B(n6545), .Z(n6539) );
  AND U5898 ( .A(n846), .B(n6538), .Z(n6545) );
  XNOR U5899 ( .A(n6546), .B(n6536), .Z(n6538) );
  XOR U5900 ( .A(n6547), .B(n6548), .Z(n6536) );
  AND U5901 ( .A(n850), .B(n6549), .Z(n6548) );
  XOR U5902 ( .A(p_input[662]), .B(n6547), .Z(n6549) );
  XOR U5903 ( .A(n6550), .B(n6551), .Z(n6547) );
  AND U5904 ( .A(n854), .B(n6552), .Z(n6551) );
  IV U5905 ( .A(n6544), .Z(n6546) );
  XOR U5906 ( .A(n6553), .B(n6554), .Z(n6544) );
  AND U5907 ( .A(n858), .B(n6555), .Z(n6554) );
  XOR U5908 ( .A(n6556), .B(n6557), .Z(n6542) );
  AND U5909 ( .A(n862), .B(n6555), .Z(n6557) );
  XNOR U5910 ( .A(n6556), .B(n6553), .Z(n6555) );
  XOR U5911 ( .A(n6558), .B(n6559), .Z(n6553) );
  AND U5912 ( .A(n865), .B(n6552), .Z(n6559) );
  XNOR U5913 ( .A(n6560), .B(n6550), .Z(n6552) );
  XOR U5914 ( .A(n6561), .B(n6562), .Z(n6550) );
  AND U5915 ( .A(n869), .B(n6563), .Z(n6562) );
  XOR U5916 ( .A(p_input[678]), .B(n6561), .Z(n6563) );
  XOR U5917 ( .A(n6564), .B(n6565), .Z(n6561) );
  AND U5918 ( .A(n873), .B(n6566), .Z(n6565) );
  IV U5919 ( .A(n6558), .Z(n6560) );
  XOR U5920 ( .A(n6567), .B(n6568), .Z(n6558) );
  AND U5921 ( .A(n877), .B(n6569), .Z(n6568) );
  XOR U5922 ( .A(n6570), .B(n6571), .Z(n6556) );
  AND U5923 ( .A(n881), .B(n6569), .Z(n6571) );
  XNOR U5924 ( .A(n6570), .B(n6567), .Z(n6569) );
  XOR U5925 ( .A(n6572), .B(n6573), .Z(n6567) );
  AND U5926 ( .A(n884), .B(n6566), .Z(n6573) );
  XNOR U5927 ( .A(n6574), .B(n6564), .Z(n6566) );
  XOR U5928 ( .A(n6575), .B(n6576), .Z(n6564) );
  AND U5929 ( .A(n888), .B(n6577), .Z(n6576) );
  XOR U5930 ( .A(p_input[694]), .B(n6575), .Z(n6577) );
  XOR U5931 ( .A(n6578), .B(n6579), .Z(n6575) );
  AND U5932 ( .A(n892), .B(n6580), .Z(n6579) );
  IV U5933 ( .A(n6572), .Z(n6574) );
  XOR U5934 ( .A(n6581), .B(n6582), .Z(n6572) );
  AND U5935 ( .A(n896), .B(n6583), .Z(n6582) );
  XOR U5936 ( .A(n6584), .B(n6585), .Z(n6570) );
  AND U5937 ( .A(n900), .B(n6583), .Z(n6585) );
  XNOR U5938 ( .A(n6584), .B(n6581), .Z(n6583) );
  XOR U5939 ( .A(n6586), .B(n6587), .Z(n6581) );
  AND U5940 ( .A(n903), .B(n6580), .Z(n6587) );
  XNOR U5941 ( .A(n6588), .B(n6578), .Z(n6580) );
  XOR U5942 ( .A(n6589), .B(n6590), .Z(n6578) );
  AND U5943 ( .A(n907), .B(n6591), .Z(n6590) );
  XOR U5944 ( .A(p_input[710]), .B(n6589), .Z(n6591) );
  XOR U5945 ( .A(n6592), .B(n6593), .Z(n6589) );
  AND U5946 ( .A(n911), .B(n6594), .Z(n6593) );
  IV U5947 ( .A(n6586), .Z(n6588) );
  XOR U5948 ( .A(n6595), .B(n6596), .Z(n6586) );
  AND U5949 ( .A(n915), .B(n6597), .Z(n6596) );
  XOR U5950 ( .A(n6598), .B(n6599), .Z(n6584) );
  AND U5951 ( .A(n919), .B(n6597), .Z(n6599) );
  XNOR U5952 ( .A(n6598), .B(n6595), .Z(n6597) );
  XOR U5953 ( .A(n6600), .B(n6601), .Z(n6595) );
  AND U5954 ( .A(n922), .B(n6594), .Z(n6601) );
  XNOR U5955 ( .A(n6602), .B(n6592), .Z(n6594) );
  XOR U5956 ( .A(n6603), .B(n6604), .Z(n6592) );
  AND U5957 ( .A(n926), .B(n6605), .Z(n6604) );
  XOR U5958 ( .A(p_input[726]), .B(n6603), .Z(n6605) );
  XOR U5959 ( .A(n6606), .B(n6607), .Z(n6603) );
  AND U5960 ( .A(n930), .B(n6608), .Z(n6607) );
  IV U5961 ( .A(n6600), .Z(n6602) );
  XOR U5962 ( .A(n6609), .B(n6610), .Z(n6600) );
  AND U5963 ( .A(n934), .B(n6611), .Z(n6610) );
  XOR U5964 ( .A(n6612), .B(n6613), .Z(n6598) );
  AND U5965 ( .A(n938), .B(n6611), .Z(n6613) );
  XNOR U5966 ( .A(n6612), .B(n6609), .Z(n6611) );
  XOR U5967 ( .A(n6614), .B(n6615), .Z(n6609) );
  AND U5968 ( .A(n941), .B(n6608), .Z(n6615) );
  XNOR U5969 ( .A(n6616), .B(n6606), .Z(n6608) );
  XOR U5970 ( .A(n6617), .B(n6618), .Z(n6606) );
  AND U5971 ( .A(n945), .B(n6619), .Z(n6618) );
  XOR U5972 ( .A(p_input[742]), .B(n6617), .Z(n6619) );
  XOR U5973 ( .A(n6620), .B(n6621), .Z(n6617) );
  AND U5974 ( .A(n949), .B(n6622), .Z(n6621) );
  IV U5975 ( .A(n6614), .Z(n6616) );
  XOR U5976 ( .A(n6623), .B(n6624), .Z(n6614) );
  AND U5977 ( .A(n953), .B(n6625), .Z(n6624) );
  XOR U5978 ( .A(n6626), .B(n6627), .Z(n6612) );
  AND U5979 ( .A(n957), .B(n6625), .Z(n6627) );
  XNOR U5980 ( .A(n6626), .B(n6623), .Z(n6625) );
  XOR U5981 ( .A(n6628), .B(n6629), .Z(n6623) );
  AND U5982 ( .A(n960), .B(n6622), .Z(n6629) );
  XNOR U5983 ( .A(n6630), .B(n6620), .Z(n6622) );
  XOR U5984 ( .A(n6631), .B(n6632), .Z(n6620) );
  AND U5985 ( .A(n964), .B(n6633), .Z(n6632) );
  XOR U5986 ( .A(p_input[758]), .B(n6631), .Z(n6633) );
  XOR U5987 ( .A(n6634), .B(n6635), .Z(n6631) );
  AND U5988 ( .A(n968), .B(n6636), .Z(n6635) );
  IV U5989 ( .A(n6628), .Z(n6630) );
  XOR U5990 ( .A(n6637), .B(n6638), .Z(n6628) );
  AND U5991 ( .A(n972), .B(n6639), .Z(n6638) );
  XOR U5992 ( .A(n6640), .B(n6641), .Z(n6626) );
  AND U5993 ( .A(n976), .B(n6639), .Z(n6641) );
  XNOR U5994 ( .A(n6640), .B(n6637), .Z(n6639) );
  XOR U5995 ( .A(n6642), .B(n6643), .Z(n6637) );
  AND U5996 ( .A(n979), .B(n6636), .Z(n6643) );
  XNOR U5997 ( .A(n6644), .B(n6634), .Z(n6636) );
  XOR U5998 ( .A(n6645), .B(n6646), .Z(n6634) );
  AND U5999 ( .A(n983), .B(n6647), .Z(n6646) );
  XOR U6000 ( .A(p_input[774]), .B(n6645), .Z(n6647) );
  XOR U6001 ( .A(n6648), .B(n6649), .Z(n6645) );
  AND U6002 ( .A(n987), .B(n6650), .Z(n6649) );
  IV U6003 ( .A(n6642), .Z(n6644) );
  XOR U6004 ( .A(n6651), .B(n6652), .Z(n6642) );
  AND U6005 ( .A(n991), .B(n6653), .Z(n6652) );
  XOR U6006 ( .A(n6654), .B(n6655), .Z(n6640) );
  AND U6007 ( .A(n995), .B(n6653), .Z(n6655) );
  XNOR U6008 ( .A(n6654), .B(n6651), .Z(n6653) );
  XOR U6009 ( .A(n6656), .B(n6657), .Z(n6651) );
  AND U6010 ( .A(n998), .B(n6650), .Z(n6657) );
  XNOR U6011 ( .A(n6658), .B(n6648), .Z(n6650) );
  XOR U6012 ( .A(n6659), .B(n6660), .Z(n6648) );
  AND U6013 ( .A(n1002), .B(n6661), .Z(n6660) );
  XOR U6014 ( .A(p_input[790]), .B(n6659), .Z(n6661) );
  XOR U6015 ( .A(n6662), .B(n6663), .Z(n6659) );
  AND U6016 ( .A(n1006), .B(n6664), .Z(n6663) );
  IV U6017 ( .A(n6656), .Z(n6658) );
  XOR U6018 ( .A(n6665), .B(n6666), .Z(n6656) );
  AND U6019 ( .A(n1010), .B(n6667), .Z(n6666) );
  XOR U6020 ( .A(n6668), .B(n6669), .Z(n6654) );
  AND U6021 ( .A(n1014), .B(n6667), .Z(n6669) );
  XNOR U6022 ( .A(n6668), .B(n6665), .Z(n6667) );
  XOR U6023 ( .A(n6670), .B(n6671), .Z(n6665) );
  AND U6024 ( .A(n1017), .B(n6664), .Z(n6671) );
  XNOR U6025 ( .A(n6672), .B(n6662), .Z(n6664) );
  XOR U6026 ( .A(n6673), .B(n6674), .Z(n6662) );
  AND U6027 ( .A(n1021), .B(n6675), .Z(n6674) );
  XOR U6028 ( .A(p_input[806]), .B(n6673), .Z(n6675) );
  XOR U6029 ( .A(n6676), .B(n6677), .Z(n6673) );
  AND U6030 ( .A(n1025), .B(n6678), .Z(n6677) );
  IV U6031 ( .A(n6670), .Z(n6672) );
  XOR U6032 ( .A(n6679), .B(n6680), .Z(n6670) );
  AND U6033 ( .A(n1029), .B(n6681), .Z(n6680) );
  XOR U6034 ( .A(n6682), .B(n6683), .Z(n6668) );
  AND U6035 ( .A(n1033), .B(n6681), .Z(n6683) );
  XNOR U6036 ( .A(n6682), .B(n6679), .Z(n6681) );
  XOR U6037 ( .A(n6684), .B(n6685), .Z(n6679) );
  AND U6038 ( .A(n1036), .B(n6678), .Z(n6685) );
  XNOR U6039 ( .A(n6686), .B(n6676), .Z(n6678) );
  XOR U6040 ( .A(n6687), .B(n6688), .Z(n6676) );
  AND U6041 ( .A(n1040), .B(n6689), .Z(n6688) );
  XOR U6042 ( .A(p_input[822]), .B(n6687), .Z(n6689) );
  XOR U6043 ( .A(n6690), .B(n6691), .Z(n6687) );
  AND U6044 ( .A(n1044), .B(n6692), .Z(n6691) );
  IV U6045 ( .A(n6684), .Z(n6686) );
  XOR U6046 ( .A(n6693), .B(n6694), .Z(n6684) );
  AND U6047 ( .A(n1048), .B(n6695), .Z(n6694) );
  XOR U6048 ( .A(n6696), .B(n6697), .Z(n6682) );
  AND U6049 ( .A(n1052), .B(n6695), .Z(n6697) );
  XNOR U6050 ( .A(n6696), .B(n6693), .Z(n6695) );
  XOR U6051 ( .A(n6698), .B(n6699), .Z(n6693) );
  AND U6052 ( .A(n1055), .B(n6692), .Z(n6699) );
  XNOR U6053 ( .A(n6700), .B(n6690), .Z(n6692) );
  XOR U6054 ( .A(n6701), .B(n6702), .Z(n6690) );
  AND U6055 ( .A(n1059), .B(n6703), .Z(n6702) );
  XOR U6056 ( .A(p_input[838]), .B(n6701), .Z(n6703) );
  XOR U6057 ( .A(n6704), .B(n6705), .Z(n6701) );
  AND U6058 ( .A(n1063), .B(n6706), .Z(n6705) );
  IV U6059 ( .A(n6698), .Z(n6700) );
  XOR U6060 ( .A(n6707), .B(n6708), .Z(n6698) );
  AND U6061 ( .A(n1067), .B(n6709), .Z(n6708) );
  XOR U6062 ( .A(n6710), .B(n6711), .Z(n6696) );
  AND U6063 ( .A(n1071), .B(n6709), .Z(n6711) );
  XNOR U6064 ( .A(n6710), .B(n6707), .Z(n6709) );
  XOR U6065 ( .A(n6712), .B(n6713), .Z(n6707) );
  AND U6066 ( .A(n1074), .B(n6706), .Z(n6713) );
  XNOR U6067 ( .A(n6714), .B(n6704), .Z(n6706) );
  XOR U6068 ( .A(n6715), .B(n6716), .Z(n6704) );
  AND U6069 ( .A(n1078), .B(n6717), .Z(n6716) );
  XOR U6070 ( .A(p_input[854]), .B(n6715), .Z(n6717) );
  XOR U6071 ( .A(n6718), .B(n6719), .Z(n6715) );
  AND U6072 ( .A(n1082), .B(n6720), .Z(n6719) );
  IV U6073 ( .A(n6712), .Z(n6714) );
  XOR U6074 ( .A(n6721), .B(n6722), .Z(n6712) );
  AND U6075 ( .A(n1086), .B(n6723), .Z(n6722) );
  XOR U6076 ( .A(n6724), .B(n6725), .Z(n6710) );
  AND U6077 ( .A(n1090), .B(n6723), .Z(n6725) );
  XNOR U6078 ( .A(n6724), .B(n6721), .Z(n6723) );
  XOR U6079 ( .A(n6726), .B(n6727), .Z(n6721) );
  AND U6080 ( .A(n1093), .B(n6720), .Z(n6727) );
  XNOR U6081 ( .A(n6728), .B(n6718), .Z(n6720) );
  XOR U6082 ( .A(n6729), .B(n6730), .Z(n6718) );
  AND U6083 ( .A(n1097), .B(n6731), .Z(n6730) );
  XOR U6084 ( .A(p_input[870]), .B(n6729), .Z(n6731) );
  XOR U6085 ( .A(n6732), .B(n6733), .Z(n6729) );
  AND U6086 ( .A(n1101), .B(n6734), .Z(n6733) );
  IV U6087 ( .A(n6726), .Z(n6728) );
  XOR U6088 ( .A(n6735), .B(n6736), .Z(n6726) );
  AND U6089 ( .A(n1105), .B(n6737), .Z(n6736) );
  XOR U6090 ( .A(n6738), .B(n6739), .Z(n6724) );
  AND U6091 ( .A(n1109), .B(n6737), .Z(n6739) );
  XNOR U6092 ( .A(n6738), .B(n6735), .Z(n6737) );
  XOR U6093 ( .A(n6740), .B(n6741), .Z(n6735) );
  AND U6094 ( .A(n1112), .B(n6734), .Z(n6741) );
  XNOR U6095 ( .A(n6742), .B(n6732), .Z(n6734) );
  XOR U6096 ( .A(n6743), .B(n6744), .Z(n6732) );
  AND U6097 ( .A(n1116), .B(n6745), .Z(n6744) );
  XOR U6098 ( .A(p_input[886]), .B(n6743), .Z(n6745) );
  XOR U6099 ( .A(n6746), .B(n6747), .Z(n6743) );
  AND U6100 ( .A(n1120), .B(n6748), .Z(n6747) );
  IV U6101 ( .A(n6740), .Z(n6742) );
  XOR U6102 ( .A(n6749), .B(n6750), .Z(n6740) );
  AND U6103 ( .A(n1124), .B(n6751), .Z(n6750) );
  XOR U6104 ( .A(n6752), .B(n6753), .Z(n6738) );
  AND U6105 ( .A(n1128), .B(n6751), .Z(n6753) );
  XNOR U6106 ( .A(n6752), .B(n6749), .Z(n6751) );
  XOR U6107 ( .A(n6754), .B(n6755), .Z(n6749) );
  AND U6108 ( .A(n1131), .B(n6748), .Z(n6755) );
  XNOR U6109 ( .A(n6756), .B(n6746), .Z(n6748) );
  XOR U6110 ( .A(n6757), .B(n6758), .Z(n6746) );
  AND U6111 ( .A(n1135), .B(n6759), .Z(n6758) );
  XOR U6112 ( .A(p_input[902]), .B(n6757), .Z(n6759) );
  XOR U6113 ( .A(n6760), .B(n6761), .Z(n6757) );
  AND U6114 ( .A(n1139), .B(n6762), .Z(n6761) );
  IV U6115 ( .A(n6754), .Z(n6756) );
  XOR U6116 ( .A(n6763), .B(n6764), .Z(n6754) );
  AND U6117 ( .A(n1143), .B(n6765), .Z(n6764) );
  XOR U6118 ( .A(n6766), .B(n6767), .Z(n6752) );
  AND U6119 ( .A(n1147), .B(n6765), .Z(n6767) );
  XNOR U6120 ( .A(n6766), .B(n6763), .Z(n6765) );
  XOR U6121 ( .A(n6768), .B(n6769), .Z(n6763) );
  AND U6122 ( .A(n1150), .B(n6762), .Z(n6769) );
  XNOR U6123 ( .A(n6770), .B(n6760), .Z(n6762) );
  XOR U6124 ( .A(n6771), .B(n6772), .Z(n6760) );
  AND U6125 ( .A(n1154), .B(n6773), .Z(n6772) );
  XOR U6126 ( .A(p_input[918]), .B(n6771), .Z(n6773) );
  XOR U6127 ( .A(n6774), .B(n6775), .Z(n6771) );
  AND U6128 ( .A(n1158), .B(n6776), .Z(n6775) );
  IV U6129 ( .A(n6768), .Z(n6770) );
  XOR U6130 ( .A(n6777), .B(n6778), .Z(n6768) );
  AND U6131 ( .A(n1162), .B(n6779), .Z(n6778) );
  XOR U6132 ( .A(n6780), .B(n6781), .Z(n6766) );
  AND U6133 ( .A(n1166), .B(n6779), .Z(n6781) );
  XNOR U6134 ( .A(n6780), .B(n6777), .Z(n6779) );
  XOR U6135 ( .A(n6782), .B(n6783), .Z(n6777) );
  AND U6136 ( .A(n1169), .B(n6776), .Z(n6783) );
  XNOR U6137 ( .A(n6784), .B(n6774), .Z(n6776) );
  XOR U6138 ( .A(n6785), .B(n6786), .Z(n6774) );
  AND U6139 ( .A(n1173), .B(n6787), .Z(n6786) );
  XOR U6140 ( .A(p_input[934]), .B(n6785), .Z(n6787) );
  XOR U6141 ( .A(n6788), .B(n6789), .Z(n6785) );
  AND U6142 ( .A(n1177), .B(n6790), .Z(n6789) );
  IV U6143 ( .A(n6782), .Z(n6784) );
  XOR U6144 ( .A(n6791), .B(n6792), .Z(n6782) );
  AND U6145 ( .A(n1181), .B(n6793), .Z(n6792) );
  XOR U6146 ( .A(n6794), .B(n6795), .Z(n6780) );
  AND U6147 ( .A(n1185), .B(n6793), .Z(n6795) );
  XNOR U6148 ( .A(n6794), .B(n6791), .Z(n6793) );
  XOR U6149 ( .A(n6796), .B(n6797), .Z(n6791) );
  AND U6150 ( .A(n1188), .B(n6790), .Z(n6797) );
  XNOR U6151 ( .A(n6798), .B(n6788), .Z(n6790) );
  XOR U6152 ( .A(n6799), .B(n6800), .Z(n6788) );
  AND U6153 ( .A(n1192), .B(n6801), .Z(n6800) );
  XOR U6154 ( .A(p_input[950]), .B(n6799), .Z(n6801) );
  XOR U6155 ( .A(n6802), .B(n6803), .Z(n6799) );
  AND U6156 ( .A(n1196), .B(n6804), .Z(n6803) );
  IV U6157 ( .A(n6796), .Z(n6798) );
  XOR U6158 ( .A(n6805), .B(n6806), .Z(n6796) );
  AND U6159 ( .A(n1200), .B(n6807), .Z(n6806) );
  XOR U6160 ( .A(n6808), .B(n6809), .Z(n6794) );
  AND U6161 ( .A(n1204), .B(n6807), .Z(n6809) );
  XNOR U6162 ( .A(n6808), .B(n6805), .Z(n6807) );
  XOR U6163 ( .A(n6810), .B(n6811), .Z(n6805) );
  AND U6164 ( .A(n1207), .B(n6804), .Z(n6811) );
  XNOR U6165 ( .A(n6812), .B(n6802), .Z(n6804) );
  XOR U6166 ( .A(n6813), .B(n6814), .Z(n6802) );
  AND U6167 ( .A(n1211), .B(n6815), .Z(n6814) );
  XOR U6168 ( .A(p_input[966]), .B(n6813), .Z(n6815) );
  XOR U6169 ( .A(n6816), .B(n6817), .Z(n6813) );
  AND U6170 ( .A(n1215), .B(n6818), .Z(n6817) );
  IV U6171 ( .A(n6810), .Z(n6812) );
  XOR U6172 ( .A(n6819), .B(n6820), .Z(n6810) );
  AND U6173 ( .A(n1219), .B(n6821), .Z(n6820) );
  XOR U6174 ( .A(n6822), .B(n6823), .Z(n6808) );
  AND U6175 ( .A(n1223), .B(n6821), .Z(n6823) );
  XNOR U6176 ( .A(n6822), .B(n6819), .Z(n6821) );
  XOR U6177 ( .A(n6824), .B(n6825), .Z(n6819) );
  AND U6178 ( .A(n1226), .B(n6818), .Z(n6825) );
  XNOR U6179 ( .A(n6826), .B(n6816), .Z(n6818) );
  XOR U6180 ( .A(n6827), .B(n6828), .Z(n6816) );
  AND U6181 ( .A(n1230), .B(n6829), .Z(n6828) );
  XOR U6182 ( .A(p_input[982]), .B(n6827), .Z(n6829) );
  XOR U6183 ( .A(n6830), .B(n6831), .Z(n6827) );
  AND U6184 ( .A(n1234), .B(n6832), .Z(n6831) );
  IV U6185 ( .A(n6824), .Z(n6826) );
  XOR U6186 ( .A(n6833), .B(n6834), .Z(n6824) );
  AND U6187 ( .A(n1238), .B(n6835), .Z(n6834) );
  XOR U6188 ( .A(n6836), .B(n6837), .Z(n6822) );
  AND U6189 ( .A(n1242), .B(n6835), .Z(n6837) );
  XNOR U6190 ( .A(n6836), .B(n6833), .Z(n6835) );
  XOR U6191 ( .A(n6838), .B(n6839), .Z(n6833) );
  AND U6192 ( .A(n1245), .B(n6832), .Z(n6839) );
  XNOR U6193 ( .A(n6840), .B(n6830), .Z(n6832) );
  XOR U6194 ( .A(n6841), .B(n6842), .Z(n6830) );
  AND U6195 ( .A(n1249), .B(n6843), .Z(n6842) );
  XOR U6196 ( .A(p_input[998]), .B(n6841), .Z(n6843) );
  XOR U6197 ( .A(n6844), .B(n6845), .Z(n6841) );
  AND U6198 ( .A(n1253), .B(n6846), .Z(n6845) );
  IV U6199 ( .A(n6838), .Z(n6840) );
  XOR U6200 ( .A(n6847), .B(n6848), .Z(n6838) );
  AND U6201 ( .A(n1257), .B(n6849), .Z(n6848) );
  XOR U6202 ( .A(n6850), .B(n6851), .Z(n6836) );
  AND U6203 ( .A(n1261), .B(n6849), .Z(n6851) );
  XNOR U6204 ( .A(n6850), .B(n6847), .Z(n6849) );
  XOR U6205 ( .A(n6852), .B(n6853), .Z(n6847) );
  AND U6206 ( .A(n1264), .B(n6846), .Z(n6853) );
  XNOR U6207 ( .A(n6854), .B(n6844), .Z(n6846) );
  XOR U6208 ( .A(n6855), .B(n6856), .Z(n6844) );
  AND U6209 ( .A(n1268), .B(n6857), .Z(n6856) );
  XOR U6210 ( .A(p_input[1014]), .B(n6855), .Z(n6857) );
  XOR U6211 ( .A(n6858), .B(n6859), .Z(n6855) );
  AND U6212 ( .A(n1272), .B(n6860), .Z(n6859) );
  IV U6213 ( .A(n6852), .Z(n6854) );
  XOR U6214 ( .A(n6861), .B(n6862), .Z(n6852) );
  AND U6215 ( .A(n1276), .B(n6863), .Z(n6862) );
  XOR U6216 ( .A(n6864), .B(n6865), .Z(n6850) );
  AND U6217 ( .A(n1280), .B(n6863), .Z(n6865) );
  XNOR U6218 ( .A(n6864), .B(n6861), .Z(n6863) );
  XOR U6219 ( .A(n6866), .B(n6867), .Z(n6861) );
  AND U6220 ( .A(n1283), .B(n6860), .Z(n6867) );
  XNOR U6221 ( .A(n6868), .B(n6858), .Z(n6860) );
  XOR U6222 ( .A(n6869), .B(n6870), .Z(n6858) );
  AND U6223 ( .A(n1287), .B(n6871), .Z(n6870) );
  XOR U6224 ( .A(p_input[1030]), .B(n6869), .Z(n6871) );
  XOR U6225 ( .A(n6872), .B(n6873), .Z(n6869) );
  AND U6226 ( .A(n1291), .B(n6874), .Z(n6873) );
  IV U6227 ( .A(n6866), .Z(n6868) );
  XOR U6228 ( .A(n6875), .B(n6876), .Z(n6866) );
  AND U6229 ( .A(n1295), .B(n6877), .Z(n6876) );
  XOR U6230 ( .A(n6878), .B(n6879), .Z(n6864) );
  AND U6231 ( .A(n1299), .B(n6877), .Z(n6879) );
  XNOR U6232 ( .A(n6878), .B(n6875), .Z(n6877) );
  XOR U6233 ( .A(n6880), .B(n6881), .Z(n6875) );
  AND U6234 ( .A(n1302), .B(n6874), .Z(n6881) );
  XNOR U6235 ( .A(n6882), .B(n6872), .Z(n6874) );
  XOR U6236 ( .A(n6883), .B(n6884), .Z(n6872) );
  AND U6237 ( .A(n1306), .B(n6885), .Z(n6884) );
  XOR U6238 ( .A(p_input[1046]), .B(n6883), .Z(n6885) );
  XOR U6239 ( .A(n6886), .B(n6887), .Z(n6883) );
  AND U6240 ( .A(n1310), .B(n6888), .Z(n6887) );
  IV U6241 ( .A(n6880), .Z(n6882) );
  XOR U6242 ( .A(n6889), .B(n6890), .Z(n6880) );
  AND U6243 ( .A(n1314), .B(n6891), .Z(n6890) );
  XOR U6244 ( .A(n6892), .B(n6893), .Z(n6878) );
  AND U6245 ( .A(n1318), .B(n6891), .Z(n6893) );
  XNOR U6246 ( .A(n6892), .B(n6889), .Z(n6891) );
  XOR U6247 ( .A(n6894), .B(n6895), .Z(n6889) );
  AND U6248 ( .A(n1321), .B(n6888), .Z(n6895) );
  XNOR U6249 ( .A(n6896), .B(n6886), .Z(n6888) );
  XOR U6250 ( .A(n6897), .B(n6898), .Z(n6886) );
  AND U6251 ( .A(n1325), .B(n6899), .Z(n6898) );
  XOR U6252 ( .A(p_input[1062]), .B(n6897), .Z(n6899) );
  XOR U6253 ( .A(n6900), .B(n6901), .Z(n6897) );
  AND U6254 ( .A(n1329), .B(n6902), .Z(n6901) );
  IV U6255 ( .A(n6894), .Z(n6896) );
  XOR U6256 ( .A(n6903), .B(n6904), .Z(n6894) );
  AND U6257 ( .A(n1333), .B(n6905), .Z(n6904) );
  XOR U6258 ( .A(n6906), .B(n6907), .Z(n6892) );
  AND U6259 ( .A(n1337), .B(n6905), .Z(n6907) );
  XNOR U6260 ( .A(n6906), .B(n6903), .Z(n6905) );
  XOR U6261 ( .A(n6908), .B(n6909), .Z(n6903) );
  AND U6262 ( .A(n1340), .B(n6902), .Z(n6909) );
  XNOR U6263 ( .A(n6910), .B(n6900), .Z(n6902) );
  XOR U6264 ( .A(n6911), .B(n6912), .Z(n6900) );
  AND U6265 ( .A(n1344), .B(n6913), .Z(n6912) );
  XOR U6266 ( .A(p_input[1078]), .B(n6911), .Z(n6913) );
  XOR U6267 ( .A(n6914), .B(n6915), .Z(n6911) );
  AND U6268 ( .A(n1348), .B(n6916), .Z(n6915) );
  IV U6269 ( .A(n6908), .Z(n6910) );
  XOR U6270 ( .A(n6917), .B(n6918), .Z(n6908) );
  AND U6271 ( .A(n1352), .B(n6919), .Z(n6918) );
  XOR U6272 ( .A(n6920), .B(n6921), .Z(n6906) );
  AND U6273 ( .A(n1356), .B(n6919), .Z(n6921) );
  XNOR U6274 ( .A(n6920), .B(n6917), .Z(n6919) );
  XOR U6275 ( .A(n6922), .B(n6923), .Z(n6917) );
  AND U6276 ( .A(n1359), .B(n6916), .Z(n6923) );
  XNOR U6277 ( .A(n6924), .B(n6914), .Z(n6916) );
  XOR U6278 ( .A(n6925), .B(n6926), .Z(n6914) );
  AND U6279 ( .A(n1363), .B(n6927), .Z(n6926) );
  XOR U6280 ( .A(p_input[1094]), .B(n6925), .Z(n6927) );
  XOR U6281 ( .A(n6928), .B(n6929), .Z(n6925) );
  AND U6282 ( .A(n1367), .B(n6930), .Z(n6929) );
  IV U6283 ( .A(n6922), .Z(n6924) );
  XOR U6284 ( .A(n6931), .B(n6932), .Z(n6922) );
  AND U6285 ( .A(n1371), .B(n6933), .Z(n6932) );
  XOR U6286 ( .A(n6934), .B(n6935), .Z(n6920) );
  AND U6287 ( .A(n1375), .B(n6933), .Z(n6935) );
  XNOR U6288 ( .A(n6934), .B(n6931), .Z(n6933) );
  XOR U6289 ( .A(n6936), .B(n6937), .Z(n6931) );
  AND U6290 ( .A(n1378), .B(n6930), .Z(n6937) );
  XNOR U6291 ( .A(n6938), .B(n6928), .Z(n6930) );
  XOR U6292 ( .A(n6939), .B(n6940), .Z(n6928) );
  AND U6293 ( .A(n1382), .B(n6941), .Z(n6940) );
  XOR U6294 ( .A(p_input[1110]), .B(n6939), .Z(n6941) );
  XOR U6295 ( .A(n6942), .B(n6943), .Z(n6939) );
  AND U6296 ( .A(n1386), .B(n6944), .Z(n6943) );
  IV U6297 ( .A(n6936), .Z(n6938) );
  XOR U6298 ( .A(n6945), .B(n6946), .Z(n6936) );
  AND U6299 ( .A(n1390), .B(n6947), .Z(n6946) );
  XOR U6300 ( .A(n6948), .B(n6949), .Z(n6934) );
  AND U6301 ( .A(n1394), .B(n6947), .Z(n6949) );
  XNOR U6302 ( .A(n6948), .B(n6945), .Z(n6947) );
  XOR U6303 ( .A(n6950), .B(n6951), .Z(n6945) );
  AND U6304 ( .A(n1397), .B(n6944), .Z(n6951) );
  XNOR U6305 ( .A(n6952), .B(n6942), .Z(n6944) );
  XOR U6306 ( .A(n6953), .B(n6954), .Z(n6942) );
  AND U6307 ( .A(n1401), .B(n6955), .Z(n6954) );
  XOR U6308 ( .A(p_input[1126]), .B(n6953), .Z(n6955) );
  XOR U6309 ( .A(n6956), .B(n6957), .Z(n6953) );
  AND U6310 ( .A(n1405), .B(n6958), .Z(n6957) );
  IV U6311 ( .A(n6950), .Z(n6952) );
  XOR U6312 ( .A(n6959), .B(n6960), .Z(n6950) );
  AND U6313 ( .A(n1409), .B(n6961), .Z(n6960) );
  XOR U6314 ( .A(n6962), .B(n6963), .Z(n6948) );
  AND U6315 ( .A(n1413), .B(n6961), .Z(n6963) );
  XNOR U6316 ( .A(n6962), .B(n6959), .Z(n6961) );
  XOR U6317 ( .A(n6964), .B(n6965), .Z(n6959) );
  AND U6318 ( .A(n1416), .B(n6958), .Z(n6965) );
  XNOR U6319 ( .A(n6966), .B(n6956), .Z(n6958) );
  XOR U6320 ( .A(n6967), .B(n6968), .Z(n6956) );
  AND U6321 ( .A(n1420), .B(n6969), .Z(n6968) );
  XOR U6322 ( .A(p_input[1142]), .B(n6967), .Z(n6969) );
  XOR U6323 ( .A(n6970), .B(n6971), .Z(n6967) );
  AND U6324 ( .A(n1424), .B(n6972), .Z(n6971) );
  IV U6325 ( .A(n6964), .Z(n6966) );
  XOR U6326 ( .A(n6973), .B(n6974), .Z(n6964) );
  AND U6327 ( .A(n1428), .B(n6975), .Z(n6974) );
  XOR U6328 ( .A(n6976), .B(n6977), .Z(n6962) );
  AND U6329 ( .A(n1432), .B(n6975), .Z(n6977) );
  XNOR U6330 ( .A(n6976), .B(n6973), .Z(n6975) );
  XOR U6331 ( .A(n6978), .B(n6979), .Z(n6973) );
  AND U6332 ( .A(n1435), .B(n6972), .Z(n6979) );
  XNOR U6333 ( .A(n6980), .B(n6970), .Z(n6972) );
  XOR U6334 ( .A(n6981), .B(n6982), .Z(n6970) );
  AND U6335 ( .A(n1439), .B(n6983), .Z(n6982) );
  XOR U6336 ( .A(p_input[1158]), .B(n6981), .Z(n6983) );
  XOR U6337 ( .A(n6984), .B(n6985), .Z(n6981) );
  AND U6338 ( .A(n1443), .B(n6986), .Z(n6985) );
  IV U6339 ( .A(n6978), .Z(n6980) );
  XOR U6340 ( .A(n6987), .B(n6988), .Z(n6978) );
  AND U6341 ( .A(n1447), .B(n6989), .Z(n6988) );
  XOR U6342 ( .A(n6990), .B(n6991), .Z(n6976) );
  AND U6343 ( .A(n1451), .B(n6989), .Z(n6991) );
  XNOR U6344 ( .A(n6990), .B(n6987), .Z(n6989) );
  XOR U6345 ( .A(n6992), .B(n6993), .Z(n6987) );
  AND U6346 ( .A(n1454), .B(n6986), .Z(n6993) );
  XNOR U6347 ( .A(n6994), .B(n6984), .Z(n6986) );
  XOR U6348 ( .A(n6995), .B(n6996), .Z(n6984) );
  AND U6349 ( .A(n1458), .B(n6997), .Z(n6996) );
  XOR U6350 ( .A(p_input[1174]), .B(n6995), .Z(n6997) );
  XOR U6351 ( .A(n6998), .B(n6999), .Z(n6995) );
  AND U6352 ( .A(n1462), .B(n7000), .Z(n6999) );
  IV U6353 ( .A(n6992), .Z(n6994) );
  XOR U6354 ( .A(n7001), .B(n7002), .Z(n6992) );
  AND U6355 ( .A(n1466), .B(n7003), .Z(n7002) );
  XOR U6356 ( .A(n7004), .B(n7005), .Z(n6990) );
  AND U6357 ( .A(n1470), .B(n7003), .Z(n7005) );
  XNOR U6358 ( .A(n7004), .B(n7001), .Z(n7003) );
  XOR U6359 ( .A(n7006), .B(n7007), .Z(n7001) );
  AND U6360 ( .A(n1473), .B(n7000), .Z(n7007) );
  XNOR U6361 ( .A(n7008), .B(n6998), .Z(n7000) );
  XOR U6362 ( .A(n7009), .B(n7010), .Z(n6998) );
  AND U6363 ( .A(n1477), .B(n7011), .Z(n7010) );
  XOR U6364 ( .A(p_input[1190]), .B(n7009), .Z(n7011) );
  XOR U6365 ( .A(n7012), .B(n7013), .Z(n7009) );
  AND U6366 ( .A(n1481), .B(n7014), .Z(n7013) );
  IV U6367 ( .A(n7006), .Z(n7008) );
  XOR U6368 ( .A(n7015), .B(n7016), .Z(n7006) );
  AND U6369 ( .A(n1485), .B(n7017), .Z(n7016) );
  XOR U6370 ( .A(n7018), .B(n7019), .Z(n7004) );
  AND U6371 ( .A(n1489), .B(n7017), .Z(n7019) );
  XNOR U6372 ( .A(n7018), .B(n7015), .Z(n7017) );
  XOR U6373 ( .A(n7020), .B(n7021), .Z(n7015) );
  AND U6374 ( .A(n1492), .B(n7014), .Z(n7021) );
  XNOR U6375 ( .A(n7022), .B(n7012), .Z(n7014) );
  XOR U6376 ( .A(n7023), .B(n7024), .Z(n7012) );
  AND U6377 ( .A(n1496), .B(n7025), .Z(n7024) );
  XOR U6378 ( .A(p_input[1206]), .B(n7023), .Z(n7025) );
  XOR U6379 ( .A(n7026), .B(n7027), .Z(n7023) );
  AND U6380 ( .A(n1500), .B(n7028), .Z(n7027) );
  IV U6381 ( .A(n7020), .Z(n7022) );
  XOR U6382 ( .A(n7029), .B(n7030), .Z(n7020) );
  AND U6383 ( .A(n1504), .B(n7031), .Z(n7030) );
  XOR U6384 ( .A(n7032), .B(n7033), .Z(n7018) );
  AND U6385 ( .A(n1508), .B(n7031), .Z(n7033) );
  XNOR U6386 ( .A(n7032), .B(n7029), .Z(n7031) );
  XOR U6387 ( .A(n7034), .B(n7035), .Z(n7029) );
  AND U6388 ( .A(n1511), .B(n7028), .Z(n7035) );
  XNOR U6389 ( .A(n7036), .B(n7026), .Z(n7028) );
  XOR U6390 ( .A(n7037), .B(n7038), .Z(n7026) );
  AND U6391 ( .A(n1515), .B(n7039), .Z(n7038) );
  XOR U6392 ( .A(p_input[1222]), .B(n7037), .Z(n7039) );
  XOR U6393 ( .A(n7040), .B(n7041), .Z(n7037) );
  AND U6394 ( .A(n1519), .B(n7042), .Z(n7041) );
  IV U6395 ( .A(n7034), .Z(n7036) );
  XOR U6396 ( .A(n7043), .B(n7044), .Z(n7034) );
  AND U6397 ( .A(n1523), .B(n7045), .Z(n7044) );
  XOR U6398 ( .A(n7046), .B(n7047), .Z(n7032) );
  AND U6399 ( .A(n1527), .B(n7045), .Z(n7047) );
  XNOR U6400 ( .A(n7046), .B(n7043), .Z(n7045) );
  XOR U6401 ( .A(n7048), .B(n7049), .Z(n7043) );
  AND U6402 ( .A(n1530), .B(n7042), .Z(n7049) );
  XNOR U6403 ( .A(n7050), .B(n7040), .Z(n7042) );
  XOR U6404 ( .A(n7051), .B(n7052), .Z(n7040) );
  AND U6405 ( .A(n1534), .B(n7053), .Z(n7052) );
  XOR U6406 ( .A(p_input[1238]), .B(n7051), .Z(n7053) );
  XOR U6407 ( .A(n7054), .B(n7055), .Z(n7051) );
  AND U6408 ( .A(n1538), .B(n7056), .Z(n7055) );
  IV U6409 ( .A(n7048), .Z(n7050) );
  XOR U6410 ( .A(n7057), .B(n7058), .Z(n7048) );
  AND U6411 ( .A(n1542), .B(n7059), .Z(n7058) );
  XOR U6412 ( .A(n7060), .B(n7061), .Z(n7046) );
  AND U6413 ( .A(n1546), .B(n7059), .Z(n7061) );
  XNOR U6414 ( .A(n7060), .B(n7057), .Z(n7059) );
  XOR U6415 ( .A(n7062), .B(n7063), .Z(n7057) );
  AND U6416 ( .A(n1549), .B(n7056), .Z(n7063) );
  XNOR U6417 ( .A(n7064), .B(n7054), .Z(n7056) );
  XOR U6418 ( .A(n7065), .B(n7066), .Z(n7054) );
  AND U6419 ( .A(n1553), .B(n7067), .Z(n7066) );
  XOR U6420 ( .A(p_input[1254]), .B(n7065), .Z(n7067) );
  XOR U6421 ( .A(n7068), .B(n7069), .Z(n7065) );
  AND U6422 ( .A(n1557), .B(n7070), .Z(n7069) );
  IV U6423 ( .A(n7062), .Z(n7064) );
  XOR U6424 ( .A(n7071), .B(n7072), .Z(n7062) );
  AND U6425 ( .A(n1561), .B(n7073), .Z(n7072) );
  XOR U6426 ( .A(n7074), .B(n7075), .Z(n7060) );
  AND U6427 ( .A(n1565), .B(n7073), .Z(n7075) );
  XNOR U6428 ( .A(n7074), .B(n7071), .Z(n7073) );
  XOR U6429 ( .A(n7076), .B(n7077), .Z(n7071) );
  AND U6430 ( .A(n1568), .B(n7070), .Z(n7077) );
  XNOR U6431 ( .A(n7078), .B(n7068), .Z(n7070) );
  XOR U6432 ( .A(n7079), .B(n7080), .Z(n7068) );
  AND U6433 ( .A(n1572), .B(n7081), .Z(n7080) );
  XOR U6434 ( .A(p_input[1270]), .B(n7079), .Z(n7081) );
  XOR U6435 ( .A(n7082), .B(n7083), .Z(n7079) );
  AND U6436 ( .A(n1576), .B(n7084), .Z(n7083) );
  IV U6437 ( .A(n7076), .Z(n7078) );
  XOR U6438 ( .A(n7085), .B(n7086), .Z(n7076) );
  AND U6439 ( .A(n1580), .B(n7087), .Z(n7086) );
  XOR U6440 ( .A(n7088), .B(n7089), .Z(n7074) );
  AND U6441 ( .A(n1584), .B(n7087), .Z(n7089) );
  XNOR U6442 ( .A(n7088), .B(n7085), .Z(n7087) );
  XOR U6443 ( .A(n7090), .B(n7091), .Z(n7085) );
  AND U6444 ( .A(n1587), .B(n7084), .Z(n7091) );
  XNOR U6445 ( .A(n7092), .B(n7082), .Z(n7084) );
  XOR U6446 ( .A(n7093), .B(n7094), .Z(n7082) );
  AND U6447 ( .A(n1591), .B(n7095), .Z(n7094) );
  XOR U6448 ( .A(p_input[1286]), .B(n7093), .Z(n7095) );
  XOR U6449 ( .A(n7096), .B(n7097), .Z(n7093) );
  AND U6450 ( .A(n1595), .B(n7098), .Z(n7097) );
  IV U6451 ( .A(n7090), .Z(n7092) );
  XOR U6452 ( .A(n7099), .B(n7100), .Z(n7090) );
  AND U6453 ( .A(n1599), .B(n7101), .Z(n7100) );
  XOR U6454 ( .A(n7102), .B(n7103), .Z(n7088) );
  AND U6455 ( .A(n1603), .B(n7101), .Z(n7103) );
  XNOR U6456 ( .A(n7102), .B(n7099), .Z(n7101) );
  XOR U6457 ( .A(n7104), .B(n7105), .Z(n7099) );
  AND U6458 ( .A(n1606), .B(n7098), .Z(n7105) );
  XNOR U6459 ( .A(n7106), .B(n7096), .Z(n7098) );
  XOR U6460 ( .A(n7107), .B(n7108), .Z(n7096) );
  AND U6461 ( .A(n1610), .B(n7109), .Z(n7108) );
  XOR U6462 ( .A(p_input[1302]), .B(n7107), .Z(n7109) );
  XOR U6463 ( .A(n7110), .B(n7111), .Z(n7107) );
  AND U6464 ( .A(n1614), .B(n7112), .Z(n7111) );
  IV U6465 ( .A(n7104), .Z(n7106) );
  XOR U6466 ( .A(n7113), .B(n7114), .Z(n7104) );
  AND U6467 ( .A(n1618), .B(n7115), .Z(n7114) );
  XOR U6468 ( .A(n7116), .B(n7117), .Z(n7102) );
  AND U6469 ( .A(n1622), .B(n7115), .Z(n7117) );
  XNOR U6470 ( .A(n7116), .B(n7113), .Z(n7115) );
  XOR U6471 ( .A(n7118), .B(n7119), .Z(n7113) );
  AND U6472 ( .A(n1625), .B(n7112), .Z(n7119) );
  XNOR U6473 ( .A(n7120), .B(n7110), .Z(n7112) );
  XOR U6474 ( .A(n7121), .B(n7122), .Z(n7110) );
  AND U6475 ( .A(n1629), .B(n7123), .Z(n7122) );
  XOR U6476 ( .A(p_input[1318]), .B(n7121), .Z(n7123) );
  XOR U6477 ( .A(n7124), .B(n7125), .Z(n7121) );
  AND U6478 ( .A(n1633), .B(n7126), .Z(n7125) );
  IV U6479 ( .A(n7118), .Z(n7120) );
  XOR U6480 ( .A(n7127), .B(n7128), .Z(n7118) );
  AND U6481 ( .A(n1637), .B(n7129), .Z(n7128) );
  XOR U6482 ( .A(n7130), .B(n7131), .Z(n7116) );
  AND U6483 ( .A(n1641), .B(n7129), .Z(n7131) );
  XNOR U6484 ( .A(n7130), .B(n7127), .Z(n7129) );
  XOR U6485 ( .A(n7132), .B(n7133), .Z(n7127) );
  AND U6486 ( .A(n1644), .B(n7126), .Z(n7133) );
  XNOR U6487 ( .A(n7134), .B(n7124), .Z(n7126) );
  XOR U6488 ( .A(n7135), .B(n7136), .Z(n7124) );
  AND U6489 ( .A(n1648), .B(n7137), .Z(n7136) );
  XOR U6490 ( .A(p_input[1334]), .B(n7135), .Z(n7137) );
  XOR U6491 ( .A(n7138), .B(n7139), .Z(n7135) );
  AND U6492 ( .A(n1652), .B(n7140), .Z(n7139) );
  IV U6493 ( .A(n7132), .Z(n7134) );
  XOR U6494 ( .A(n7141), .B(n7142), .Z(n7132) );
  AND U6495 ( .A(n1656), .B(n7143), .Z(n7142) );
  XOR U6496 ( .A(n7144), .B(n7145), .Z(n7130) );
  AND U6497 ( .A(n1660), .B(n7143), .Z(n7145) );
  XNOR U6498 ( .A(n7144), .B(n7141), .Z(n7143) );
  XOR U6499 ( .A(n7146), .B(n7147), .Z(n7141) );
  AND U6500 ( .A(n1663), .B(n7140), .Z(n7147) );
  XNOR U6501 ( .A(n7148), .B(n7138), .Z(n7140) );
  XOR U6502 ( .A(n7149), .B(n7150), .Z(n7138) );
  AND U6503 ( .A(n1667), .B(n7151), .Z(n7150) );
  XOR U6504 ( .A(p_input[1350]), .B(n7149), .Z(n7151) );
  XOR U6505 ( .A(n7152), .B(n7153), .Z(n7149) );
  AND U6506 ( .A(n1671), .B(n7154), .Z(n7153) );
  IV U6507 ( .A(n7146), .Z(n7148) );
  XOR U6508 ( .A(n7155), .B(n7156), .Z(n7146) );
  AND U6509 ( .A(n1675), .B(n7157), .Z(n7156) );
  XOR U6510 ( .A(n7158), .B(n7159), .Z(n7144) );
  AND U6511 ( .A(n1679), .B(n7157), .Z(n7159) );
  XNOR U6512 ( .A(n7158), .B(n7155), .Z(n7157) );
  XOR U6513 ( .A(n7160), .B(n7161), .Z(n7155) );
  AND U6514 ( .A(n1682), .B(n7154), .Z(n7161) );
  XNOR U6515 ( .A(n7162), .B(n7152), .Z(n7154) );
  XOR U6516 ( .A(n7163), .B(n7164), .Z(n7152) );
  AND U6517 ( .A(n1686), .B(n7165), .Z(n7164) );
  XOR U6518 ( .A(p_input[1366]), .B(n7163), .Z(n7165) );
  XOR U6519 ( .A(n7166), .B(n7167), .Z(n7163) );
  AND U6520 ( .A(n1690), .B(n7168), .Z(n7167) );
  IV U6521 ( .A(n7160), .Z(n7162) );
  XOR U6522 ( .A(n7169), .B(n7170), .Z(n7160) );
  AND U6523 ( .A(n1694), .B(n7171), .Z(n7170) );
  XOR U6524 ( .A(n7172), .B(n7173), .Z(n7158) );
  AND U6525 ( .A(n1698), .B(n7171), .Z(n7173) );
  XNOR U6526 ( .A(n7172), .B(n7169), .Z(n7171) );
  XOR U6527 ( .A(n7174), .B(n7175), .Z(n7169) );
  AND U6528 ( .A(n1701), .B(n7168), .Z(n7175) );
  XNOR U6529 ( .A(n7176), .B(n7166), .Z(n7168) );
  XOR U6530 ( .A(n7177), .B(n7178), .Z(n7166) );
  AND U6531 ( .A(n1705), .B(n7179), .Z(n7178) );
  XOR U6532 ( .A(p_input[1382]), .B(n7177), .Z(n7179) );
  XOR U6533 ( .A(n7180), .B(n7181), .Z(n7177) );
  AND U6534 ( .A(n1709), .B(n7182), .Z(n7181) );
  IV U6535 ( .A(n7174), .Z(n7176) );
  XOR U6536 ( .A(n7183), .B(n7184), .Z(n7174) );
  AND U6537 ( .A(n1713), .B(n7185), .Z(n7184) );
  XOR U6538 ( .A(n7186), .B(n7187), .Z(n7172) );
  AND U6539 ( .A(n1717), .B(n7185), .Z(n7187) );
  XNOR U6540 ( .A(n7186), .B(n7183), .Z(n7185) );
  XOR U6541 ( .A(n7188), .B(n7189), .Z(n7183) );
  AND U6542 ( .A(n1720), .B(n7182), .Z(n7189) );
  XNOR U6543 ( .A(n7190), .B(n7180), .Z(n7182) );
  XOR U6544 ( .A(n7191), .B(n7192), .Z(n7180) );
  AND U6545 ( .A(n1724), .B(n7193), .Z(n7192) );
  XOR U6546 ( .A(p_input[1398]), .B(n7191), .Z(n7193) );
  XOR U6547 ( .A(n7194), .B(n7195), .Z(n7191) );
  AND U6548 ( .A(n1728), .B(n7196), .Z(n7195) );
  IV U6549 ( .A(n7188), .Z(n7190) );
  XOR U6550 ( .A(n7197), .B(n7198), .Z(n7188) );
  AND U6551 ( .A(n1732), .B(n7199), .Z(n7198) );
  XOR U6552 ( .A(n7200), .B(n7201), .Z(n7186) );
  AND U6553 ( .A(n1736), .B(n7199), .Z(n7201) );
  XNOR U6554 ( .A(n7200), .B(n7197), .Z(n7199) );
  XOR U6555 ( .A(n7202), .B(n7203), .Z(n7197) );
  AND U6556 ( .A(n1739), .B(n7196), .Z(n7203) );
  XNOR U6557 ( .A(n7204), .B(n7194), .Z(n7196) );
  XOR U6558 ( .A(n7205), .B(n7206), .Z(n7194) );
  AND U6559 ( .A(n1743), .B(n7207), .Z(n7206) );
  XOR U6560 ( .A(p_input[1414]), .B(n7205), .Z(n7207) );
  XOR U6561 ( .A(n7208), .B(n7209), .Z(n7205) );
  AND U6562 ( .A(n1747), .B(n7210), .Z(n7209) );
  IV U6563 ( .A(n7202), .Z(n7204) );
  XOR U6564 ( .A(n7211), .B(n7212), .Z(n7202) );
  AND U6565 ( .A(n1751), .B(n7213), .Z(n7212) );
  XOR U6566 ( .A(n7214), .B(n7215), .Z(n7200) );
  AND U6567 ( .A(n1755), .B(n7213), .Z(n7215) );
  XNOR U6568 ( .A(n7214), .B(n7211), .Z(n7213) );
  XOR U6569 ( .A(n7216), .B(n7217), .Z(n7211) );
  AND U6570 ( .A(n1758), .B(n7210), .Z(n7217) );
  XNOR U6571 ( .A(n7218), .B(n7208), .Z(n7210) );
  XOR U6572 ( .A(n7219), .B(n7220), .Z(n7208) );
  AND U6573 ( .A(n1762), .B(n7221), .Z(n7220) );
  XOR U6574 ( .A(p_input[1430]), .B(n7219), .Z(n7221) );
  XOR U6575 ( .A(n7222), .B(n7223), .Z(n7219) );
  AND U6576 ( .A(n1766), .B(n7224), .Z(n7223) );
  IV U6577 ( .A(n7216), .Z(n7218) );
  XOR U6578 ( .A(n7225), .B(n7226), .Z(n7216) );
  AND U6579 ( .A(n1770), .B(n7227), .Z(n7226) );
  XOR U6580 ( .A(n7228), .B(n7229), .Z(n7214) );
  AND U6581 ( .A(n1774), .B(n7227), .Z(n7229) );
  XNOR U6582 ( .A(n7228), .B(n7225), .Z(n7227) );
  XOR U6583 ( .A(n7230), .B(n7231), .Z(n7225) );
  AND U6584 ( .A(n1777), .B(n7224), .Z(n7231) );
  XNOR U6585 ( .A(n7232), .B(n7222), .Z(n7224) );
  XOR U6586 ( .A(n7233), .B(n7234), .Z(n7222) );
  AND U6587 ( .A(n1781), .B(n7235), .Z(n7234) );
  XOR U6588 ( .A(p_input[1446]), .B(n7233), .Z(n7235) );
  XOR U6589 ( .A(n7236), .B(n7237), .Z(n7233) );
  AND U6590 ( .A(n1785), .B(n7238), .Z(n7237) );
  IV U6591 ( .A(n7230), .Z(n7232) );
  XOR U6592 ( .A(n7239), .B(n7240), .Z(n7230) );
  AND U6593 ( .A(n1789), .B(n7241), .Z(n7240) );
  XOR U6594 ( .A(n7242), .B(n7243), .Z(n7228) );
  AND U6595 ( .A(n1793), .B(n7241), .Z(n7243) );
  XNOR U6596 ( .A(n7242), .B(n7239), .Z(n7241) );
  XOR U6597 ( .A(n7244), .B(n7245), .Z(n7239) );
  AND U6598 ( .A(n1796), .B(n7238), .Z(n7245) );
  XNOR U6599 ( .A(n7246), .B(n7236), .Z(n7238) );
  XOR U6600 ( .A(n7247), .B(n7248), .Z(n7236) );
  AND U6601 ( .A(n1800), .B(n7249), .Z(n7248) );
  XOR U6602 ( .A(p_input[1462]), .B(n7247), .Z(n7249) );
  XOR U6603 ( .A(n7250), .B(n7251), .Z(n7247) );
  AND U6604 ( .A(n1804), .B(n7252), .Z(n7251) );
  IV U6605 ( .A(n7244), .Z(n7246) );
  XOR U6606 ( .A(n7253), .B(n7254), .Z(n7244) );
  AND U6607 ( .A(n1808), .B(n7255), .Z(n7254) );
  XOR U6608 ( .A(n7256), .B(n7257), .Z(n7242) );
  AND U6609 ( .A(n1812), .B(n7255), .Z(n7257) );
  XNOR U6610 ( .A(n7256), .B(n7253), .Z(n7255) );
  XOR U6611 ( .A(n7258), .B(n7259), .Z(n7253) );
  AND U6612 ( .A(n1815), .B(n7252), .Z(n7259) );
  XNOR U6613 ( .A(n7260), .B(n7250), .Z(n7252) );
  XOR U6614 ( .A(n7261), .B(n7262), .Z(n7250) );
  AND U6615 ( .A(n1819), .B(n7263), .Z(n7262) );
  XOR U6616 ( .A(p_input[1478]), .B(n7261), .Z(n7263) );
  XOR U6617 ( .A(n7264), .B(n7265), .Z(n7261) );
  AND U6618 ( .A(n1823), .B(n7266), .Z(n7265) );
  IV U6619 ( .A(n7258), .Z(n7260) );
  XOR U6620 ( .A(n7267), .B(n7268), .Z(n7258) );
  AND U6621 ( .A(n1827), .B(n7269), .Z(n7268) );
  XOR U6622 ( .A(n7270), .B(n7271), .Z(n7256) );
  AND U6623 ( .A(n1831), .B(n7269), .Z(n7271) );
  XNOR U6624 ( .A(n7270), .B(n7267), .Z(n7269) );
  XOR U6625 ( .A(n7272), .B(n7273), .Z(n7267) );
  AND U6626 ( .A(n1834), .B(n7266), .Z(n7273) );
  XNOR U6627 ( .A(n7274), .B(n7264), .Z(n7266) );
  XOR U6628 ( .A(n7275), .B(n7276), .Z(n7264) );
  AND U6629 ( .A(n1838), .B(n7277), .Z(n7276) );
  XOR U6630 ( .A(p_input[1494]), .B(n7275), .Z(n7277) );
  XOR U6631 ( .A(n7278), .B(n7279), .Z(n7275) );
  AND U6632 ( .A(n1842), .B(n7280), .Z(n7279) );
  IV U6633 ( .A(n7272), .Z(n7274) );
  XOR U6634 ( .A(n7281), .B(n7282), .Z(n7272) );
  AND U6635 ( .A(n1846), .B(n7283), .Z(n7282) );
  XOR U6636 ( .A(n7284), .B(n7285), .Z(n7270) );
  AND U6637 ( .A(n1850), .B(n7283), .Z(n7285) );
  XNOR U6638 ( .A(n7284), .B(n7281), .Z(n7283) );
  XOR U6639 ( .A(n7286), .B(n7287), .Z(n7281) );
  AND U6640 ( .A(n1853), .B(n7280), .Z(n7287) );
  XNOR U6641 ( .A(n7288), .B(n7278), .Z(n7280) );
  XOR U6642 ( .A(n7289), .B(n7290), .Z(n7278) );
  AND U6643 ( .A(n1857), .B(n7291), .Z(n7290) );
  XOR U6644 ( .A(p_input[1510]), .B(n7289), .Z(n7291) );
  XOR U6645 ( .A(n7292), .B(n7293), .Z(n7289) );
  AND U6646 ( .A(n1861), .B(n7294), .Z(n7293) );
  IV U6647 ( .A(n7286), .Z(n7288) );
  XOR U6648 ( .A(n7295), .B(n7296), .Z(n7286) );
  AND U6649 ( .A(n1865), .B(n7297), .Z(n7296) );
  XOR U6650 ( .A(n7298), .B(n7299), .Z(n7284) );
  AND U6651 ( .A(n1869), .B(n7297), .Z(n7299) );
  XNOR U6652 ( .A(n7298), .B(n7295), .Z(n7297) );
  XOR U6653 ( .A(n7300), .B(n7301), .Z(n7295) );
  AND U6654 ( .A(n1872), .B(n7294), .Z(n7301) );
  XNOR U6655 ( .A(n7302), .B(n7292), .Z(n7294) );
  XOR U6656 ( .A(n7303), .B(n7304), .Z(n7292) );
  AND U6657 ( .A(n1876), .B(n7305), .Z(n7304) );
  XOR U6658 ( .A(p_input[1526]), .B(n7303), .Z(n7305) );
  XOR U6659 ( .A(n7306), .B(n7307), .Z(n7303) );
  AND U6660 ( .A(n1880), .B(n7308), .Z(n7307) );
  IV U6661 ( .A(n7300), .Z(n7302) );
  XOR U6662 ( .A(n7309), .B(n7310), .Z(n7300) );
  AND U6663 ( .A(n1884), .B(n7311), .Z(n7310) );
  XOR U6664 ( .A(n7312), .B(n7313), .Z(n7298) );
  AND U6665 ( .A(n1888), .B(n7311), .Z(n7313) );
  XNOR U6666 ( .A(n7312), .B(n7309), .Z(n7311) );
  XOR U6667 ( .A(n7314), .B(n7315), .Z(n7309) );
  AND U6668 ( .A(n1891), .B(n7308), .Z(n7315) );
  XNOR U6669 ( .A(n7316), .B(n7306), .Z(n7308) );
  XOR U6670 ( .A(n7317), .B(n7318), .Z(n7306) );
  AND U6671 ( .A(n1895), .B(n7319), .Z(n7318) );
  XOR U6672 ( .A(p_input[1542]), .B(n7317), .Z(n7319) );
  XOR U6673 ( .A(n7320), .B(n7321), .Z(n7317) );
  AND U6674 ( .A(n1899), .B(n7322), .Z(n7321) );
  IV U6675 ( .A(n7314), .Z(n7316) );
  XOR U6676 ( .A(n7323), .B(n7324), .Z(n7314) );
  AND U6677 ( .A(n1903), .B(n7325), .Z(n7324) );
  XOR U6678 ( .A(n7326), .B(n7327), .Z(n7312) );
  AND U6679 ( .A(n1907), .B(n7325), .Z(n7327) );
  XNOR U6680 ( .A(n7326), .B(n7323), .Z(n7325) );
  XOR U6681 ( .A(n7328), .B(n7329), .Z(n7323) );
  AND U6682 ( .A(n1910), .B(n7322), .Z(n7329) );
  XNOR U6683 ( .A(n7330), .B(n7320), .Z(n7322) );
  XOR U6684 ( .A(n7331), .B(n7332), .Z(n7320) );
  AND U6685 ( .A(n1914), .B(n7333), .Z(n7332) );
  XOR U6686 ( .A(p_input[1558]), .B(n7331), .Z(n7333) );
  XOR U6687 ( .A(n7334), .B(n7335), .Z(n7331) );
  AND U6688 ( .A(n1918), .B(n7336), .Z(n7335) );
  IV U6689 ( .A(n7328), .Z(n7330) );
  XOR U6690 ( .A(n7337), .B(n7338), .Z(n7328) );
  AND U6691 ( .A(n1922), .B(n7339), .Z(n7338) );
  XOR U6692 ( .A(n7340), .B(n7341), .Z(n7326) );
  AND U6693 ( .A(n1926), .B(n7339), .Z(n7341) );
  XNOR U6694 ( .A(n7340), .B(n7337), .Z(n7339) );
  XOR U6695 ( .A(n7342), .B(n7343), .Z(n7337) );
  AND U6696 ( .A(n1929), .B(n7336), .Z(n7343) );
  XNOR U6697 ( .A(n7344), .B(n7334), .Z(n7336) );
  XOR U6698 ( .A(n7345), .B(n7346), .Z(n7334) );
  AND U6699 ( .A(n1933), .B(n7347), .Z(n7346) );
  XOR U6700 ( .A(p_input[1574]), .B(n7345), .Z(n7347) );
  XOR U6701 ( .A(n7348), .B(n7349), .Z(n7345) );
  AND U6702 ( .A(n1937), .B(n7350), .Z(n7349) );
  IV U6703 ( .A(n7342), .Z(n7344) );
  XOR U6704 ( .A(n7351), .B(n7352), .Z(n7342) );
  AND U6705 ( .A(n1941), .B(n7353), .Z(n7352) );
  XOR U6706 ( .A(n7354), .B(n7355), .Z(n7340) );
  AND U6707 ( .A(n1945), .B(n7353), .Z(n7355) );
  XNOR U6708 ( .A(n7354), .B(n7351), .Z(n7353) );
  XOR U6709 ( .A(n7356), .B(n7357), .Z(n7351) );
  AND U6710 ( .A(n1948), .B(n7350), .Z(n7357) );
  XNOR U6711 ( .A(n7358), .B(n7348), .Z(n7350) );
  XOR U6712 ( .A(n7359), .B(n7360), .Z(n7348) );
  AND U6713 ( .A(n1952), .B(n7361), .Z(n7360) );
  XOR U6714 ( .A(p_input[1590]), .B(n7359), .Z(n7361) );
  XOR U6715 ( .A(n7362), .B(n7363), .Z(n7359) );
  AND U6716 ( .A(n1956), .B(n7364), .Z(n7363) );
  IV U6717 ( .A(n7356), .Z(n7358) );
  XOR U6718 ( .A(n7365), .B(n7366), .Z(n7356) );
  AND U6719 ( .A(n1960), .B(n7367), .Z(n7366) );
  XOR U6720 ( .A(n7368), .B(n7369), .Z(n7354) );
  AND U6721 ( .A(n1964), .B(n7367), .Z(n7369) );
  XNOR U6722 ( .A(n7368), .B(n7365), .Z(n7367) );
  XOR U6723 ( .A(n7370), .B(n7371), .Z(n7365) );
  AND U6724 ( .A(n1967), .B(n7364), .Z(n7371) );
  XNOR U6725 ( .A(n7372), .B(n7362), .Z(n7364) );
  XOR U6726 ( .A(n7373), .B(n7374), .Z(n7362) );
  AND U6727 ( .A(n1971), .B(n7375), .Z(n7374) );
  XOR U6728 ( .A(p_input[1606]), .B(n7373), .Z(n7375) );
  XOR U6729 ( .A(n7376), .B(n7377), .Z(n7373) );
  AND U6730 ( .A(n1975), .B(n7378), .Z(n7377) );
  IV U6731 ( .A(n7370), .Z(n7372) );
  XOR U6732 ( .A(n7379), .B(n7380), .Z(n7370) );
  AND U6733 ( .A(n1979), .B(n7381), .Z(n7380) );
  XOR U6734 ( .A(n7382), .B(n7383), .Z(n7368) );
  AND U6735 ( .A(n1983), .B(n7381), .Z(n7383) );
  XNOR U6736 ( .A(n7382), .B(n7379), .Z(n7381) );
  XOR U6737 ( .A(n7384), .B(n7385), .Z(n7379) );
  AND U6738 ( .A(n1986), .B(n7378), .Z(n7385) );
  XNOR U6739 ( .A(n7386), .B(n7376), .Z(n7378) );
  XOR U6740 ( .A(n7387), .B(n7388), .Z(n7376) );
  AND U6741 ( .A(n1990), .B(n7389), .Z(n7388) );
  XOR U6742 ( .A(p_input[1622]), .B(n7387), .Z(n7389) );
  XOR U6743 ( .A(n7390), .B(n7391), .Z(n7387) );
  AND U6744 ( .A(n1994), .B(n7392), .Z(n7391) );
  IV U6745 ( .A(n7384), .Z(n7386) );
  XOR U6746 ( .A(n7393), .B(n7394), .Z(n7384) );
  AND U6747 ( .A(n1998), .B(n7395), .Z(n7394) );
  XOR U6748 ( .A(n7396), .B(n7397), .Z(n7382) );
  AND U6749 ( .A(n2002), .B(n7395), .Z(n7397) );
  XNOR U6750 ( .A(n7396), .B(n7393), .Z(n7395) );
  XOR U6751 ( .A(n7398), .B(n7399), .Z(n7393) );
  AND U6752 ( .A(n2005), .B(n7392), .Z(n7399) );
  XNOR U6753 ( .A(n7400), .B(n7390), .Z(n7392) );
  XOR U6754 ( .A(n7401), .B(n7402), .Z(n7390) );
  AND U6755 ( .A(n2009), .B(n7403), .Z(n7402) );
  XOR U6756 ( .A(p_input[1638]), .B(n7401), .Z(n7403) );
  XOR U6757 ( .A(n7404), .B(n7405), .Z(n7401) );
  AND U6758 ( .A(n2013), .B(n7406), .Z(n7405) );
  IV U6759 ( .A(n7398), .Z(n7400) );
  XOR U6760 ( .A(n7407), .B(n7408), .Z(n7398) );
  AND U6761 ( .A(n2017), .B(n7409), .Z(n7408) );
  XOR U6762 ( .A(n7410), .B(n7411), .Z(n7396) );
  AND U6763 ( .A(n2021), .B(n7409), .Z(n7411) );
  XNOR U6764 ( .A(n7410), .B(n7407), .Z(n7409) );
  XOR U6765 ( .A(n7412), .B(n7413), .Z(n7407) );
  AND U6766 ( .A(n2024), .B(n7406), .Z(n7413) );
  XNOR U6767 ( .A(n7414), .B(n7404), .Z(n7406) );
  XOR U6768 ( .A(n7415), .B(n7416), .Z(n7404) );
  AND U6769 ( .A(n2028), .B(n7417), .Z(n7416) );
  XOR U6770 ( .A(p_input[1654]), .B(n7415), .Z(n7417) );
  XOR U6771 ( .A(n7418), .B(n7419), .Z(n7415) );
  AND U6772 ( .A(n2032), .B(n7420), .Z(n7419) );
  IV U6773 ( .A(n7412), .Z(n7414) );
  XOR U6774 ( .A(n7421), .B(n7422), .Z(n7412) );
  AND U6775 ( .A(n2036), .B(n7423), .Z(n7422) );
  XOR U6776 ( .A(n7424), .B(n7425), .Z(n7410) );
  AND U6777 ( .A(n2040), .B(n7423), .Z(n7425) );
  XNOR U6778 ( .A(n7424), .B(n7421), .Z(n7423) );
  XOR U6779 ( .A(n7426), .B(n7427), .Z(n7421) );
  AND U6780 ( .A(n2043), .B(n7420), .Z(n7427) );
  XNOR U6781 ( .A(n7428), .B(n7418), .Z(n7420) );
  XOR U6782 ( .A(n7429), .B(n7430), .Z(n7418) );
  AND U6783 ( .A(n2047), .B(n7431), .Z(n7430) );
  XOR U6784 ( .A(p_input[1670]), .B(n7429), .Z(n7431) );
  XOR U6785 ( .A(n7432), .B(n7433), .Z(n7429) );
  AND U6786 ( .A(n2051), .B(n7434), .Z(n7433) );
  IV U6787 ( .A(n7426), .Z(n7428) );
  XOR U6788 ( .A(n7435), .B(n7436), .Z(n7426) );
  AND U6789 ( .A(n2055), .B(n7437), .Z(n7436) );
  XOR U6790 ( .A(n7438), .B(n7439), .Z(n7424) );
  AND U6791 ( .A(n2059), .B(n7437), .Z(n7439) );
  XNOR U6792 ( .A(n7438), .B(n7435), .Z(n7437) );
  XOR U6793 ( .A(n7440), .B(n7441), .Z(n7435) );
  AND U6794 ( .A(n2062), .B(n7434), .Z(n7441) );
  XNOR U6795 ( .A(n7442), .B(n7432), .Z(n7434) );
  XOR U6796 ( .A(n7443), .B(n7444), .Z(n7432) );
  AND U6797 ( .A(n2066), .B(n7445), .Z(n7444) );
  XOR U6798 ( .A(p_input[1686]), .B(n7443), .Z(n7445) );
  XOR U6799 ( .A(n7446), .B(n7447), .Z(n7443) );
  AND U6800 ( .A(n2070), .B(n7448), .Z(n7447) );
  IV U6801 ( .A(n7440), .Z(n7442) );
  XOR U6802 ( .A(n7449), .B(n7450), .Z(n7440) );
  AND U6803 ( .A(n2074), .B(n7451), .Z(n7450) );
  XOR U6804 ( .A(n7452), .B(n7453), .Z(n7438) );
  AND U6805 ( .A(n2078), .B(n7451), .Z(n7453) );
  XNOR U6806 ( .A(n7452), .B(n7449), .Z(n7451) );
  XOR U6807 ( .A(n7454), .B(n7455), .Z(n7449) );
  AND U6808 ( .A(n2081), .B(n7448), .Z(n7455) );
  XNOR U6809 ( .A(n7456), .B(n7446), .Z(n7448) );
  XOR U6810 ( .A(n7457), .B(n7458), .Z(n7446) );
  AND U6811 ( .A(n2085), .B(n7459), .Z(n7458) );
  XOR U6812 ( .A(p_input[1702]), .B(n7457), .Z(n7459) );
  XOR U6813 ( .A(n7460), .B(n7461), .Z(n7457) );
  AND U6814 ( .A(n2089), .B(n7462), .Z(n7461) );
  IV U6815 ( .A(n7454), .Z(n7456) );
  XOR U6816 ( .A(n7463), .B(n7464), .Z(n7454) );
  AND U6817 ( .A(n2093), .B(n7465), .Z(n7464) );
  XOR U6818 ( .A(n7466), .B(n7467), .Z(n7452) );
  AND U6819 ( .A(n2097), .B(n7465), .Z(n7467) );
  XNOR U6820 ( .A(n7466), .B(n7463), .Z(n7465) );
  XOR U6821 ( .A(n7468), .B(n7469), .Z(n7463) );
  AND U6822 ( .A(n2100), .B(n7462), .Z(n7469) );
  XNOR U6823 ( .A(n7470), .B(n7460), .Z(n7462) );
  XOR U6824 ( .A(n7471), .B(n7472), .Z(n7460) );
  AND U6825 ( .A(n2104), .B(n7473), .Z(n7472) );
  XOR U6826 ( .A(p_input[1718]), .B(n7471), .Z(n7473) );
  XOR U6827 ( .A(n7474), .B(n7475), .Z(n7471) );
  AND U6828 ( .A(n2108), .B(n7476), .Z(n7475) );
  IV U6829 ( .A(n7468), .Z(n7470) );
  XOR U6830 ( .A(n7477), .B(n7478), .Z(n7468) );
  AND U6831 ( .A(n2112), .B(n7479), .Z(n7478) );
  XOR U6832 ( .A(n7480), .B(n7481), .Z(n7466) );
  AND U6833 ( .A(n2116), .B(n7479), .Z(n7481) );
  XNOR U6834 ( .A(n7480), .B(n7477), .Z(n7479) );
  XOR U6835 ( .A(n7482), .B(n7483), .Z(n7477) );
  AND U6836 ( .A(n2119), .B(n7476), .Z(n7483) );
  XNOR U6837 ( .A(n7484), .B(n7474), .Z(n7476) );
  XOR U6838 ( .A(n7485), .B(n7486), .Z(n7474) );
  AND U6839 ( .A(n2123), .B(n7487), .Z(n7486) );
  XOR U6840 ( .A(p_input[1734]), .B(n7485), .Z(n7487) );
  XOR U6841 ( .A(n7488), .B(n7489), .Z(n7485) );
  AND U6842 ( .A(n2127), .B(n7490), .Z(n7489) );
  IV U6843 ( .A(n7482), .Z(n7484) );
  XOR U6844 ( .A(n7491), .B(n7492), .Z(n7482) );
  AND U6845 ( .A(n2131), .B(n7493), .Z(n7492) );
  XOR U6846 ( .A(n7494), .B(n7495), .Z(n7480) );
  AND U6847 ( .A(n2135), .B(n7493), .Z(n7495) );
  XNOR U6848 ( .A(n7494), .B(n7491), .Z(n7493) );
  XOR U6849 ( .A(n7496), .B(n7497), .Z(n7491) );
  AND U6850 ( .A(n2138), .B(n7490), .Z(n7497) );
  XNOR U6851 ( .A(n7498), .B(n7488), .Z(n7490) );
  XOR U6852 ( .A(n7499), .B(n7500), .Z(n7488) );
  AND U6853 ( .A(n2142), .B(n7501), .Z(n7500) );
  XOR U6854 ( .A(p_input[1750]), .B(n7499), .Z(n7501) );
  XOR U6855 ( .A(n7502), .B(n7503), .Z(n7499) );
  AND U6856 ( .A(n2146), .B(n7504), .Z(n7503) );
  IV U6857 ( .A(n7496), .Z(n7498) );
  XOR U6858 ( .A(n7505), .B(n7506), .Z(n7496) );
  AND U6859 ( .A(n2150), .B(n7507), .Z(n7506) );
  XOR U6860 ( .A(n7508), .B(n7509), .Z(n7494) );
  AND U6861 ( .A(n2154), .B(n7507), .Z(n7509) );
  XNOR U6862 ( .A(n7508), .B(n7505), .Z(n7507) );
  XOR U6863 ( .A(n7510), .B(n7511), .Z(n7505) );
  AND U6864 ( .A(n2157), .B(n7504), .Z(n7511) );
  XNOR U6865 ( .A(n7512), .B(n7502), .Z(n7504) );
  XOR U6866 ( .A(n7513), .B(n7514), .Z(n7502) );
  AND U6867 ( .A(n2161), .B(n7515), .Z(n7514) );
  XOR U6868 ( .A(p_input[1766]), .B(n7513), .Z(n7515) );
  XOR U6869 ( .A(n7516), .B(n7517), .Z(n7513) );
  AND U6870 ( .A(n2165), .B(n7518), .Z(n7517) );
  IV U6871 ( .A(n7510), .Z(n7512) );
  XOR U6872 ( .A(n7519), .B(n7520), .Z(n7510) );
  AND U6873 ( .A(n2169), .B(n7521), .Z(n7520) );
  XOR U6874 ( .A(n7522), .B(n7523), .Z(n7508) );
  AND U6875 ( .A(n2173), .B(n7521), .Z(n7523) );
  XNOR U6876 ( .A(n7522), .B(n7519), .Z(n7521) );
  XOR U6877 ( .A(n7524), .B(n7525), .Z(n7519) );
  AND U6878 ( .A(n2176), .B(n7518), .Z(n7525) );
  XNOR U6879 ( .A(n7526), .B(n7516), .Z(n7518) );
  XOR U6880 ( .A(n7527), .B(n7528), .Z(n7516) );
  AND U6881 ( .A(n2180), .B(n7529), .Z(n7528) );
  XOR U6882 ( .A(p_input[1782]), .B(n7527), .Z(n7529) );
  XOR U6883 ( .A(n7530), .B(n7531), .Z(n7527) );
  AND U6884 ( .A(n2184), .B(n7532), .Z(n7531) );
  IV U6885 ( .A(n7524), .Z(n7526) );
  XOR U6886 ( .A(n7533), .B(n7534), .Z(n7524) );
  AND U6887 ( .A(n2188), .B(n7535), .Z(n7534) );
  XOR U6888 ( .A(n7536), .B(n7537), .Z(n7522) );
  AND U6889 ( .A(n2192), .B(n7535), .Z(n7537) );
  XNOR U6890 ( .A(n7536), .B(n7533), .Z(n7535) );
  XOR U6891 ( .A(n7538), .B(n7539), .Z(n7533) );
  AND U6892 ( .A(n2195), .B(n7532), .Z(n7539) );
  XNOR U6893 ( .A(n7540), .B(n7530), .Z(n7532) );
  XOR U6894 ( .A(n7541), .B(n7542), .Z(n7530) );
  AND U6895 ( .A(n2199), .B(n7543), .Z(n7542) );
  XOR U6896 ( .A(p_input[1798]), .B(n7541), .Z(n7543) );
  XOR U6897 ( .A(n7544), .B(n7545), .Z(n7541) );
  AND U6898 ( .A(n2203), .B(n7546), .Z(n7545) );
  IV U6899 ( .A(n7538), .Z(n7540) );
  XOR U6900 ( .A(n7547), .B(n7548), .Z(n7538) );
  AND U6901 ( .A(n2207), .B(n7549), .Z(n7548) );
  XOR U6902 ( .A(n7550), .B(n7551), .Z(n7536) );
  AND U6903 ( .A(n2211), .B(n7549), .Z(n7551) );
  XNOR U6904 ( .A(n7550), .B(n7547), .Z(n7549) );
  XOR U6905 ( .A(n7552), .B(n7553), .Z(n7547) );
  AND U6906 ( .A(n2214), .B(n7546), .Z(n7553) );
  XNOR U6907 ( .A(n7554), .B(n7544), .Z(n7546) );
  XOR U6908 ( .A(n7555), .B(n7556), .Z(n7544) );
  AND U6909 ( .A(n2218), .B(n7557), .Z(n7556) );
  XOR U6910 ( .A(p_input[1814]), .B(n7555), .Z(n7557) );
  XOR U6911 ( .A(n7558), .B(n7559), .Z(n7555) );
  AND U6912 ( .A(n2222), .B(n7560), .Z(n7559) );
  IV U6913 ( .A(n7552), .Z(n7554) );
  XOR U6914 ( .A(n7561), .B(n7562), .Z(n7552) );
  AND U6915 ( .A(n2226), .B(n7563), .Z(n7562) );
  XOR U6916 ( .A(n7564), .B(n7565), .Z(n7550) );
  AND U6917 ( .A(n2230), .B(n7563), .Z(n7565) );
  XNOR U6918 ( .A(n7564), .B(n7561), .Z(n7563) );
  XOR U6919 ( .A(n7566), .B(n7567), .Z(n7561) );
  AND U6920 ( .A(n2233), .B(n7560), .Z(n7567) );
  XNOR U6921 ( .A(n7568), .B(n7558), .Z(n7560) );
  XOR U6922 ( .A(n7569), .B(n7570), .Z(n7558) );
  AND U6923 ( .A(n2237), .B(n7571), .Z(n7570) );
  XOR U6924 ( .A(p_input[1830]), .B(n7569), .Z(n7571) );
  XOR U6925 ( .A(n7572), .B(n7573), .Z(n7569) );
  AND U6926 ( .A(n2241), .B(n7574), .Z(n7573) );
  IV U6927 ( .A(n7566), .Z(n7568) );
  XOR U6928 ( .A(n7575), .B(n7576), .Z(n7566) );
  AND U6929 ( .A(n2245), .B(n7577), .Z(n7576) );
  XOR U6930 ( .A(n7578), .B(n7579), .Z(n7564) );
  AND U6931 ( .A(n2249), .B(n7577), .Z(n7579) );
  XNOR U6932 ( .A(n7578), .B(n7575), .Z(n7577) );
  XOR U6933 ( .A(n7580), .B(n7581), .Z(n7575) );
  AND U6934 ( .A(n2252), .B(n7574), .Z(n7581) );
  XNOR U6935 ( .A(n7582), .B(n7572), .Z(n7574) );
  XOR U6936 ( .A(n7583), .B(n7584), .Z(n7572) );
  AND U6937 ( .A(n2256), .B(n7585), .Z(n7584) );
  XOR U6938 ( .A(p_input[1846]), .B(n7583), .Z(n7585) );
  XOR U6939 ( .A(n7586), .B(n7587), .Z(n7583) );
  AND U6940 ( .A(n2260), .B(n7588), .Z(n7587) );
  IV U6941 ( .A(n7580), .Z(n7582) );
  XOR U6942 ( .A(n7589), .B(n7590), .Z(n7580) );
  AND U6943 ( .A(n2264), .B(n7591), .Z(n7590) );
  XOR U6944 ( .A(n7592), .B(n7593), .Z(n7578) );
  AND U6945 ( .A(n2268), .B(n7591), .Z(n7593) );
  XNOR U6946 ( .A(n7592), .B(n7589), .Z(n7591) );
  XOR U6947 ( .A(n7594), .B(n7595), .Z(n7589) );
  AND U6948 ( .A(n2271), .B(n7588), .Z(n7595) );
  XNOR U6949 ( .A(n7596), .B(n7586), .Z(n7588) );
  XOR U6950 ( .A(n7597), .B(n7598), .Z(n7586) );
  AND U6951 ( .A(n2275), .B(n7599), .Z(n7598) );
  XOR U6952 ( .A(p_input[1862]), .B(n7597), .Z(n7599) );
  XOR U6953 ( .A(n7600), .B(n7601), .Z(n7597) );
  AND U6954 ( .A(n2279), .B(n7602), .Z(n7601) );
  IV U6955 ( .A(n7594), .Z(n7596) );
  XOR U6956 ( .A(n7603), .B(n7604), .Z(n7594) );
  AND U6957 ( .A(n2283), .B(n7605), .Z(n7604) );
  XOR U6958 ( .A(n7606), .B(n7607), .Z(n7592) );
  AND U6959 ( .A(n2287), .B(n7605), .Z(n7607) );
  XNOR U6960 ( .A(n7606), .B(n7603), .Z(n7605) );
  XOR U6961 ( .A(n7608), .B(n7609), .Z(n7603) );
  AND U6962 ( .A(n2290), .B(n7602), .Z(n7609) );
  XNOR U6963 ( .A(n7610), .B(n7600), .Z(n7602) );
  XOR U6964 ( .A(n7611), .B(n7612), .Z(n7600) );
  AND U6965 ( .A(n2294), .B(n7613), .Z(n7612) );
  XOR U6966 ( .A(p_input[1878]), .B(n7611), .Z(n7613) );
  XOR U6967 ( .A(n7614), .B(n7615), .Z(n7611) );
  AND U6968 ( .A(n2298), .B(n7616), .Z(n7615) );
  IV U6969 ( .A(n7608), .Z(n7610) );
  XOR U6970 ( .A(n7617), .B(n7618), .Z(n7608) );
  AND U6971 ( .A(n2302), .B(n7619), .Z(n7618) );
  XOR U6972 ( .A(n7620), .B(n7621), .Z(n7606) );
  AND U6973 ( .A(n2306), .B(n7619), .Z(n7621) );
  XNOR U6974 ( .A(n7620), .B(n7617), .Z(n7619) );
  XOR U6975 ( .A(n7622), .B(n7623), .Z(n7617) );
  AND U6976 ( .A(n2309), .B(n7616), .Z(n7623) );
  XNOR U6977 ( .A(n7624), .B(n7614), .Z(n7616) );
  XOR U6978 ( .A(n7625), .B(n7626), .Z(n7614) );
  AND U6979 ( .A(n2313), .B(n7627), .Z(n7626) );
  XOR U6980 ( .A(p_input[1894]), .B(n7625), .Z(n7627) );
  XOR U6981 ( .A(n7628), .B(n7629), .Z(n7625) );
  AND U6982 ( .A(n2317), .B(n7630), .Z(n7629) );
  IV U6983 ( .A(n7622), .Z(n7624) );
  XOR U6984 ( .A(n7631), .B(n7632), .Z(n7622) );
  AND U6985 ( .A(n2321), .B(n7633), .Z(n7632) );
  XOR U6986 ( .A(n7634), .B(n7635), .Z(n7620) );
  AND U6987 ( .A(n2325), .B(n7633), .Z(n7635) );
  XNOR U6988 ( .A(n7634), .B(n7631), .Z(n7633) );
  XOR U6989 ( .A(n7636), .B(n7637), .Z(n7631) );
  AND U6990 ( .A(n2328), .B(n7630), .Z(n7637) );
  XNOR U6991 ( .A(n7638), .B(n7628), .Z(n7630) );
  XOR U6992 ( .A(n7639), .B(n7640), .Z(n7628) );
  AND U6993 ( .A(n2332), .B(n7641), .Z(n7640) );
  XOR U6994 ( .A(p_input[1910]), .B(n7639), .Z(n7641) );
  XOR U6995 ( .A(n7642), .B(n7643), .Z(n7639) );
  AND U6996 ( .A(n2336), .B(n7644), .Z(n7643) );
  IV U6997 ( .A(n7636), .Z(n7638) );
  XOR U6998 ( .A(n7645), .B(n7646), .Z(n7636) );
  AND U6999 ( .A(n2340), .B(n7647), .Z(n7646) );
  XOR U7000 ( .A(n7648), .B(n7649), .Z(n7634) );
  AND U7001 ( .A(n2344), .B(n7647), .Z(n7649) );
  XNOR U7002 ( .A(n7648), .B(n7645), .Z(n7647) );
  XOR U7003 ( .A(n7650), .B(n7651), .Z(n7645) );
  AND U7004 ( .A(n2347), .B(n7644), .Z(n7651) );
  XNOR U7005 ( .A(n7652), .B(n7642), .Z(n7644) );
  XOR U7006 ( .A(n7653), .B(n7654), .Z(n7642) );
  AND U7007 ( .A(n2351), .B(n7655), .Z(n7654) );
  XOR U7008 ( .A(p_input[1926]), .B(n7653), .Z(n7655) );
  XOR U7009 ( .A(n7656), .B(n7657), .Z(n7653) );
  AND U7010 ( .A(n2355), .B(n7658), .Z(n7657) );
  IV U7011 ( .A(n7650), .Z(n7652) );
  XOR U7012 ( .A(n7659), .B(n7660), .Z(n7650) );
  AND U7013 ( .A(n2359), .B(n7661), .Z(n7660) );
  XOR U7014 ( .A(n7662), .B(n7663), .Z(n7648) );
  AND U7015 ( .A(n2363), .B(n7661), .Z(n7663) );
  XNOR U7016 ( .A(n7662), .B(n7659), .Z(n7661) );
  XOR U7017 ( .A(n7664), .B(n7665), .Z(n7659) );
  AND U7018 ( .A(n2366), .B(n7658), .Z(n7665) );
  XNOR U7019 ( .A(n7666), .B(n7656), .Z(n7658) );
  XOR U7020 ( .A(n7667), .B(n7668), .Z(n7656) );
  AND U7021 ( .A(n2370), .B(n7669), .Z(n7668) );
  XOR U7022 ( .A(p_input[1942]), .B(n7667), .Z(n7669) );
  XOR U7023 ( .A(n7670), .B(n7671), .Z(n7667) );
  AND U7024 ( .A(n2374), .B(n7672), .Z(n7671) );
  IV U7025 ( .A(n7664), .Z(n7666) );
  XOR U7026 ( .A(n7673), .B(n7674), .Z(n7664) );
  AND U7027 ( .A(n2378), .B(n7675), .Z(n7674) );
  XOR U7028 ( .A(n7676), .B(n7677), .Z(n7662) );
  AND U7029 ( .A(n2382), .B(n7675), .Z(n7677) );
  XNOR U7030 ( .A(n7676), .B(n7673), .Z(n7675) );
  XOR U7031 ( .A(n7678), .B(n7679), .Z(n7673) );
  AND U7032 ( .A(n2385), .B(n7672), .Z(n7679) );
  XNOR U7033 ( .A(n7680), .B(n7670), .Z(n7672) );
  XOR U7034 ( .A(n7681), .B(n7682), .Z(n7670) );
  AND U7035 ( .A(n2389), .B(n7683), .Z(n7682) );
  XOR U7036 ( .A(p_input[1958]), .B(n7681), .Z(n7683) );
  XOR U7037 ( .A(n7684), .B(n7685), .Z(n7681) );
  AND U7038 ( .A(n2393), .B(n7686), .Z(n7685) );
  IV U7039 ( .A(n7678), .Z(n7680) );
  XOR U7040 ( .A(n7687), .B(n7688), .Z(n7678) );
  AND U7041 ( .A(n2397), .B(n7689), .Z(n7688) );
  XOR U7042 ( .A(n7690), .B(n7691), .Z(n7676) );
  AND U7043 ( .A(n2401), .B(n7689), .Z(n7691) );
  XNOR U7044 ( .A(n7690), .B(n7687), .Z(n7689) );
  XOR U7045 ( .A(n7692), .B(n7693), .Z(n7687) );
  AND U7046 ( .A(n2404), .B(n7686), .Z(n7693) );
  XNOR U7047 ( .A(n7694), .B(n7684), .Z(n7686) );
  XOR U7048 ( .A(n7695), .B(n7696), .Z(n7684) );
  AND U7049 ( .A(n2408), .B(n7697), .Z(n7696) );
  XOR U7050 ( .A(p_input[1974]), .B(n7695), .Z(n7697) );
  XOR U7051 ( .A(n7698), .B(n7699), .Z(n7695) );
  AND U7052 ( .A(n2412), .B(n7700), .Z(n7699) );
  IV U7053 ( .A(n7692), .Z(n7694) );
  XOR U7054 ( .A(n7701), .B(n7702), .Z(n7692) );
  AND U7055 ( .A(n2416), .B(n7703), .Z(n7702) );
  XOR U7056 ( .A(n7704), .B(n7705), .Z(n7690) );
  AND U7057 ( .A(n2420), .B(n7703), .Z(n7705) );
  XNOR U7058 ( .A(n7704), .B(n7701), .Z(n7703) );
  XOR U7059 ( .A(n7706), .B(n7707), .Z(n7701) );
  AND U7060 ( .A(n2423), .B(n7700), .Z(n7707) );
  XNOR U7061 ( .A(n7708), .B(n7698), .Z(n7700) );
  XOR U7062 ( .A(n7709), .B(n7710), .Z(n7698) );
  AND U7063 ( .A(n2427), .B(n7711), .Z(n7710) );
  XOR U7064 ( .A(p_input[1990]), .B(n7709), .Z(n7711) );
  XOR U7065 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n7712), 
        .Z(n7709) );
  AND U7066 ( .A(n2430), .B(n7713), .Z(n7712) );
  IV U7067 ( .A(n7706), .Z(n7708) );
  XOR U7068 ( .A(n7714), .B(n7715), .Z(n7706) );
  AND U7069 ( .A(n2434), .B(n7716), .Z(n7715) );
  XOR U7070 ( .A(n7717), .B(n7718), .Z(n7704) );
  AND U7071 ( .A(n2438), .B(n7716), .Z(n7718) );
  XNOR U7072 ( .A(n7717), .B(n7714), .Z(n7716) );
  XNOR U7073 ( .A(n7719), .B(n7720), .Z(n7714) );
  AND U7074 ( .A(n2441), .B(n7713), .Z(n7720) );
  XNOR U7075 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n7719), 
        .Z(n7713) );
  XNOR U7076 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n7721), 
        .Z(n7719) );
  AND U7077 ( .A(n2443), .B(n7722), .Z(n7721) );
  XNOR U7078 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n7723), .Z(n7717) );
  AND U7079 ( .A(n2446), .B(n7722), .Z(n7723) );
  XOR U7080 ( .A(n7724), .B(n7725), .Z(n7722) );
  XOR U7081 ( .A(n9), .B(n7726), .Z(o[21]) );
  AND U7082 ( .A(n62), .B(n7727), .Z(n9) );
  XOR U7083 ( .A(n10), .B(n7726), .Z(n7727) );
  XOR U7084 ( .A(n7728), .B(n35), .Z(n7726) );
  AND U7085 ( .A(n65), .B(n7729), .Z(n35) );
  XNOR U7086 ( .A(n7730), .B(n36), .Z(n7729) );
  XOR U7087 ( .A(n7731), .B(n7732), .Z(n36) );
  AND U7088 ( .A(n70), .B(n7733), .Z(n7732) );
  XOR U7089 ( .A(p_input[5]), .B(n7731), .Z(n7733) );
  XOR U7090 ( .A(n7734), .B(n7735), .Z(n7731) );
  AND U7091 ( .A(n74), .B(n7736), .Z(n7735) );
  IV U7092 ( .A(n7728), .Z(n7730) );
  XOR U7093 ( .A(n7737), .B(n7738), .Z(n7728) );
  AND U7094 ( .A(n78), .B(n7739), .Z(n7738) );
  XOR U7095 ( .A(n7740), .B(n7741), .Z(n10) );
  AND U7096 ( .A(n82), .B(n7739), .Z(n7741) );
  XNOR U7097 ( .A(n7742), .B(n7737), .Z(n7739) );
  XOR U7098 ( .A(n7743), .B(n7744), .Z(n7737) );
  AND U7099 ( .A(n86), .B(n7736), .Z(n7744) );
  XNOR U7100 ( .A(n7745), .B(n7734), .Z(n7736) );
  XOR U7101 ( .A(n7746), .B(n7747), .Z(n7734) );
  AND U7102 ( .A(n90), .B(n7748), .Z(n7747) );
  XOR U7103 ( .A(p_input[21]), .B(n7746), .Z(n7748) );
  XOR U7104 ( .A(n7749), .B(n7750), .Z(n7746) );
  AND U7105 ( .A(n94), .B(n7751), .Z(n7750) );
  IV U7106 ( .A(n7743), .Z(n7745) );
  XOR U7107 ( .A(n7752), .B(n7753), .Z(n7743) );
  AND U7108 ( .A(n98), .B(n7754), .Z(n7753) );
  IV U7109 ( .A(n7740), .Z(n7742) );
  XNOR U7110 ( .A(n7755), .B(n7756), .Z(n7740) );
  AND U7111 ( .A(n102), .B(n7754), .Z(n7756) );
  XNOR U7112 ( .A(n7755), .B(n7752), .Z(n7754) );
  XOR U7113 ( .A(n7757), .B(n7758), .Z(n7752) );
  AND U7114 ( .A(n105), .B(n7751), .Z(n7758) );
  XNOR U7115 ( .A(n7759), .B(n7749), .Z(n7751) );
  XOR U7116 ( .A(n7760), .B(n7761), .Z(n7749) );
  AND U7117 ( .A(n109), .B(n7762), .Z(n7761) );
  XOR U7118 ( .A(p_input[37]), .B(n7760), .Z(n7762) );
  XOR U7119 ( .A(n7763), .B(n7764), .Z(n7760) );
  AND U7120 ( .A(n113), .B(n7765), .Z(n7764) );
  IV U7121 ( .A(n7757), .Z(n7759) );
  XOR U7122 ( .A(n7766), .B(n7767), .Z(n7757) );
  AND U7123 ( .A(n117), .B(n7768), .Z(n7767) );
  XOR U7124 ( .A(n7769), .B(n7770), .Z(n7755) );
  AND U7125 ( .A(n121), .B(n7768), .Z(n7770) );
  XNOR U7126 ( .A(n7769), .B(n7766), .Z(n7768) );
  XOR U7127 ( .A(n7771), .B(n7772), .Z(n7766) );
  AND U7128 ( .A(n124), .B(n7765), .Z(n7772) );
  XNOR U7129 ( .A(n7773), .B(n7763), .Z(n7765) );
  XOR U7130 ( .A(n7774), .B(n7775), .Z(n7763) );
  AND U7131 ( .A(n128), .B(n7776), .Z(n7775) );
  XOR U7132 ( .A(p_input[53]), .B(n7774), .Z(n7776) );
  XOR U7133 ( .A(n7777), .B(n7778), .Z(n7774) );
  AND U7134 ( .A(n132), .B(n7779), .Z(n7778) );
  IV U7135 ( .A(n7771), .Z(n7773) );
  XOR U7136 ( .A(n7780), .B(n7781), .Z(n7771) );
  AND U7137 ( .A(n136), .B(n7782), .Z(n7781) );
  XOR U7138 ( .A(n7783), .B(n7784), .Z(n7769) );
  AND U7139 ( .A(n140), .B(n7782), .Z(n7784) );
  XNOR U7140 ( .A(n7783), .B(n7780), .Z(n7782) );
  XOR U7141 ( .A(n7785), .B(n7786), .Z(n7780) );
  AND U7142 ( .A(n143), .B(n7779), .Z(n7786) );
  XNOR U7143 ( .A(n7787), .B(n7777), .Z(n7779) );
  XOR U7144 ( .A(n7788), .B(n7789), .Z(n7777) );
  AND U7145 ( .A(n147), .B(n7790), .Z(n7789) );
  XOR U7146 ( .A(p_input[69]), .B(n7788), .Z(n7790) );
  XOR U7147 ( .A(n7791), .B(n7792), .Z(n7788) );
  AND U7148 ( .A(n151), .B(n7793), .Z(n7792) );
  IV U7149 ( .A(n7785), .Z(n7787) );
  XOR U7150 ( .A(n7794), .B(n7795), .Z(n7785) );
  AND U7151 ( .A(n155), .B(n7796), .Z(n7795) );
  XOR U7152 ( .A(n7797), .B(n7798), .Z(n7783) );
  AND U7153 ( .A(n159), .B(n7796), .Z(n7798) );
  XNOR U7154 ( .A(n7797), .B(n7794), .Z(n7796) );
  XOR U7155 ( .A(n7799), .B(n7800), .Z(n7794) );
  AND U7156 ( .A(n162), .B(n7793), .Z(n7800) );
  XNOR U7157 ( .A(n7801), .B(n7791), .Z(n7793) );
  XOR U7158 ( .A(n7802), .B(n7803), .Z(n7791) );
  AND U7159 ( .A(n166), .B(n7804), .Z(n7803) );
  XOR U7160 ( .A(p_input[85]), .B(n7802), .Z(n7804) );
  XOR U7161 ( .A(n7805), .B(n7806), .Z(n7802) );
  AND U7162 ( .A(n170), .B(n7807), .Z(n7806) );
  IV U7163 ( .A(n7799), .Z(n7801) );
  XOR U7164 ( .A(n7808), .B(n7809), .Z(n7799) );
  AND U7165 ( .A(n174), .B(n7810), .Z(n7809) );
  XOR U7166 ( .A(n7811), .B(n7812), .Z(n7797) );
  AND U7167 ( .A(n178), .B(n7810), .Z(n7812) );
  XNOR U7168 ( .A(n7811), .B(n7808), .Z(n7810) );
  XOR U7169 ( .A(n7813), .B(n7814), .Z(n7808) );
  AND U7170 ( .A(n181), .B(n7807), .Z(n7814) );
  XNOR U7171 ( .A(n7815), .B(n7805), .Z(n7807) );
  XOR U7172 ( .A(n7816), .B(n7817), .Z(n7805) );
  AND U7173 ( .A(n185), .B(n7818), .Z(n7817) );
  XOR U7174 ( .A(p_input[101]), .B(n7816), .Z(n7818) );
  XOR U7175 ( .A(n7819), .B(n7820), .Z(n7816) );
  AND U7176 ( .A(n189), .B(n7821), .Z(n7820) );
  IV U7177 ( .A(n7813), .Z(n7815) );
  XOR U7178 ( .A(n7822), .B(n7823), .Z(n7813) );
  AND U7179 ( .A(n193), .B(n7824), .Z(n7823) );
  XOR U7180 ( .A(n7825), .B(n7826), .Z(n7811) );
  AND U7181 ( .A(n197), .B(n7824), .Z(n7826) );
  XNOR U7182 ( .A(n7825), .B(n7822), .Z(n7824) );
  XOR U7183 ( .A(n7827), .B(n7828), .Z(n7822) );
  AND U7184 ( .A(n200), .B(n7821), .Z(n7828) );
  XNOR U7185 ( .A(n7829), .B(n7819), .Z(n7821) );
  XOR U7186 ( .A(n7830), .B(n7831), .Z(n7819) );
  AND U7187 ( .A(n204), .B(n7832), .Z(n7831) );
  XOR U7188 ( .A(p_input[117]), .B(n7830), .Z(n7832) );
  XOR U7189 ( .A(n7833), .B(n7834), .Z(n7830) );
  AND U7190 ( .A(n208), .B(n7835), .Z(n7834) );
  IV U7191 ( .A(n7827), .Z(n7829) );
  XOR U7192 ( .A(n7836), .B(n7837), .Z(n7827) );
  AND U7193 ( .A(n212), .B(n7838), .Z(n7837) );
  XOR U7194 ( .A(n7839), .B(n7840), .Z(n7825) );
  AND U7195 ( .A(n216), .B(n7838), .Z(n7840) );
  XNOR U7196 ( .A(n7839), .B(n7836), .Z(n7838) );
  XOR U7197 ( .A(n7841), .B(n7842), .Z(n7836) );
  AND U7198 ( .A(n219), .B(n7835), .Z(n7842) );
  XNOR U7199 ( .A(n7843), .B(n7833), .Z(n7835) );
  XOR U7200 ( .A(n7844), .B(n7845), .Z(n7833) );
  AND U7201 ( .A(n223), .B(n7846), .Z(n7845) );
  XOR U7202 ( .A(p_input[133]), .B(n7844), .Z(n7846) );
  XOR U7203 ( .A(n7847), .B(n7848), .Z(n7844) );
  AND U7204 ( .A(n227), .B(n7849), .Z(n7848) );
  IV U7205 ( .A(n7841), .Z(n7843) );
  XOR U7206 ( .A(n7850), .B(n7851), .Z(n7841) );
  AND U7207 ( .A(n231), .B(n7852), .Z(n7851) );
  XOR U7208 ( .A(n7853), .B(n7854), .Z(n7839) );
  AND U7209 ( .A(n235), .B(n7852), .Z(n7854) );
  XNOR U7210 ( .A(n7853), .B(n7850), .Z(n7852) );
  XOR U7211 ( .A(n7855), .B(n7856), .Z(n7850) );
  AND U7212 ( .A(n238), .B(n7849), .Z(n7856) );
  XNOR U7213 ( .A(n7857), .B(n7847), .Z(n7849) );
  XOR U7214 ( .A(n7858), .B(n7859), .Z(n7847) );
  AND U7215 ( .A(n242), .B(n7860), .Z(n7859) );
  XOR U7216 ( .A(p_input[149]), .B(n7858), .Z(n7860) );
  XOR U7217 ( .A(n7861), .B(n7862), .Z(n7858) );
  AND U7218 ( .A(n246), .B(n7863), .Z(n7862) );
  IV U7219 ( .A(n7855), .Z(n7857) );
  XOR U7220 ( .A(n7864), .B(n7865), .Z(n7855) );
  AND U7221 ( .A(n250), .B(n7866), .Z(n7865) );
  XOR U7222 ( .A(n7867), .B(n7868), .Z(n7853) );
  AND U7223 ( .A(n254), .B(n7866), .Z(n7868) );
  XNOR U7224 ( .A(n7867), .B(n7864), .Z(n7866) );
  XOR U7225 ( .A(n7869), .B(n7870), .Z(n7864) );
  AND U7226 ( .A(n257), .B(n7863), .Z(n7870) );
  XNOR U7227 ( .A(n7871), .B(n7861), .Z(n7863) );
  XOR U7228 ( .A(n7872), .B(n7873), .Z(n7861) );
  AND U7229 ( .A(n261), .B(n7874), .Z(n7873) );
  XOR U7230 ( .A(p_input[165]), .B(n7872), .Z(n7874) );
  XOR U7231 ( .A(n7875), .B(n7876), .Z(n7872) );
  AND U7232 ( .A(n265), .B(n7877), .Z(n7876) );
  IV U7233 ( .A(n7869), .Z(n7871) );
  XOR U7234 ( .A(n7878), .B(n7879), .Z(n7869) );
  AND U7235 ( .A(n269), .B(n7880), .Z(n7879) );
  XOR U7236 ( .A(n7881), .B(n7882), .Z(n7867) );
  AND U7237 ( .A(n273), .B(n7880), .Z(n7882) );
  XNOR U7238 ( .A(n7881), .B(n7878), .Z(n7880) );
  XOR U7239 ( .A(n7883), .B(n7884), .Z(n7878) );
  AND U7240 ( .A(n276), .B(n7877), .Z(n7884) );
  XNOR U7241 ( .A(n7885), .B(n7875), .Z(n7877) );
  XOR U7242 ( .A(n7886), .B(n7887), .Z(n7875) );
  AND U7243 ( .A(n280), .B(n7888), .Z(n7887) );
  XOR U7244 ( .A(p_input[181]), .B(n7886), .Z(n7888) );
  XOR U7245 ( .A(n7889), .B(n7890), .Z(n7886) );
  AND U7246 ( .A(n284), .B(n7891), .Z(n7890) );
  IV U7247 ( .A(n7883), .Z(n7885) );
  XOR U7248 ( .A(n7892), .B(n7893), .Z(n7883) );
  AND U7249 ( .A(n288), .B(n7894), .Z(n7893) );
  XOR U7250 ( .A(n7895), .B(n7896), .Z(n7881) );
  AND U7251 ( .A(n292), .B(n7894), .Z(n7896) );
  XNOR U7252 ( .A(n7895), .B(n7892), .Z(n7894) );
  XOR U7253 ( .A(n7897), .B(n7898), .Z(n7892) );
  AND U7254 ( .A(n295), .B(n7891), .Z(n7898) );
  XNOR U7255 ( .A(n7899), .B(n7889), .Z(n7891) );
  XOR U7256 ( .A(n7900), .B(n7901), .Z(n7889) );
  AND U7257 ( .A(n299), .B(n7902), .Z(n7901) );
  XOR U7258 ( .A(p_input[197]), .B(n7900), .Z(n7902) );
  XOR U7259 ( .A(n7903), .B(n7904), .Z(n7900) );
  AND U7260 ( .A(n303), .B(n7905), .Z(n7904) );
  IV U7261 ( .A(n7897), .Z(n7899) );
  XOR U7262 ( .A(n7906), .B(n7907), .Z(n7897) );
  AND U7263 ( .A(n307), .B(n7908), .Z(n7907) );
  XOR U7264 ( .A(n7909), .B(n7910), .Z(n7895) );
  AND U7265 ( .A(n311), .B(n7908), .Z(n7910) );
  XNOR U7266 ( .A(n7909), .B(n7906), .Z(n7908) );
  XOR U7267 ( .A(n7911), .B(n7912), .Z(n7906) );
  AND U7268 ( .A(n314), .B(n7905), .Z(n7912) );
  XNOR U7269 ( .A(n7913), .B(n7903), .Z(n7905) );
  XOR U7270 ( .A(n7914), .B(n7915), .Z(n7903) );
  AND U7271 ( .A(n318), .B(n7916), .Z(n7915) );
  XOR U7272 ( .A(p_input[213]), .B(n7914), .Z(n7916) );
  XOR U7273 ( .A(n7917), .B(n7918), .Z(n7914) );
  AND U7274 ( .A(n322), .B(n7919), .Z(n7918) );
  IV U7275 ( .A(n7911), .Z(n7913) );
  XOR U7276 ( .A(n7920), .B(n7921), .Z(n7911) );
  AND U7277 ( .A(n326), .B(n7922), .Z(n7921) );
  XOR U7278 ( .A(n7923), .B(n7924), .Z(n7909) );
  AND U7279 ( .A(n330), .B(n7922), .Z(n7924) );
  XNOR U7280 ( .A(n7923), .B(n7920), .Z(n7922) );
  XOR U7281 ( .A(n7925), .B(n7926), .Z(n7920) );
  AND U7282 ( .A(n333), .B(n7919), .Z(n7926) );
  XNOR U7283 ( .A(n7927), .B(n7917), .Z(n7919) );
  XOR U7284 ( .A(n7928), .B(n7929), .Z(n7917) );
  AND U7285 ( .A(n337), .B(n7930), .Z(n7929) );
  XOR U7286 ( .A(p_input[229]), .B(n7928), .Z(n7930) );
  XOR U7287 ( .A(n7931), .B(n7932), .Z(n7928) );
  AND U7288 ( .A(n341), .B(n7933), .Z(n7932) );
  IV U7289 ( .A(n7925), .Z(n7927) );
  XOR U7290 ( .A(n7934), .B(n7935), .Z(n7925) );
  AND U7291 ( .A(n345), .B(n7936), .Z(n7935) );
  XOR U7292 ( .A(n7937), .B(n7938), .Z(n7923) );
  AND U7293 ( .A(n349), .B(n7936), .Z(n7938) );
  XNOR U7294 ( .A(n7937), .B(n7934), .Z(n7936) );
  XOR U7295 ( .A(n7939), .B(n7940), .Z(n7934) );
  AND U7296 ( .A(n352), .B(n7933), .Z(n7940) );
  XNOR U7297 ( .A(n7941), .B(n7931), .Z(n7933) );
  XOR U7298 ( .A(n7942), .B(n7943), .Z(n7931) );
  AND U7299 ( .A(n356), .B(n7944), .Z(n7943) );
  XOR U7300 ( .A(p_input[245]), .B(n7942), .Z(n7944) );
  XOR U7301 ( .A(n7945), .B(n7946), .Z(n7942) );
  AND U7302 ( .A(n360), .B(n7947), .Z(n7946) );
  IV U7303 ( .A(n7939), .Z(n7941) );
  XOR U7304 ( .A(n7948), .B(n7949), .Z(n7939) );
  AND U7305 ( .A(n364), .B(n7950), .Z(n7949) );
  XOR U7306 ( .A(n7951), .B(n7952), .Z(n7937) );
  AND U7307 ( .A(n368), .B(n7950), .Z(n7952) );
  XNOR U7308 ( .A(n7951), .B(n7948), .Z(n7950) );
  XOR U7309 ( .A(n7953), .B(n7954), .Z(n7948) );
  AND U7310 ( .A(n371), .B(n7947), .Z(n7954) );
  XNOR U7311 ( .A(n7955), .B(n7945), .Z(n7947) );
  XOR U7312 ( .A(n7956), .B(n7957), .Z(n7945) );
  AND U7313 ( .A(n375), .B(n7958), .Z(n7957) );
  XOR U7314 ( .A(p_input[261]), .B(n7956), .Z(n7958) );
  XOR U7315 ( .A(n7959), .B(n7960), .Z(n7956) );
  AND U7316 ( .A(n379), .B(n7961), .Z(n7960) );
  IV U7317 ( .A(n7953), .Z(n7955) );
  XOR U7318 ( .A(n7962), .B(n7963), .Z(n7953) );
  AND U7319 ( .A(n383), .B(n7964), .Z(n7963) );
  XOR U7320 ( .A(n7965), .B(n7966), .Z(n7951) );
  AND U7321 ( .A(n387), .B(n7964), .Z(n7966) );
  XNOR U7322 ( .A(n7965), .B(n7962), .Z(n7964) );
  XOR U7323 ( .A(n7967), .B(n7968), .Z(n7962) );
  AND U7324 ( .A(n390), .B(n7961), .Z(n7968) );
  XNOR U7325 ( .A(n7969), .B(n7959), .Z(n7961) );
  XOR U7326 ( .A(n7970), .B(n7971), .Z(n7959) );
  AND U7327 ( .A(n394), .B(n7972), .Z(n7971) );
  XOR U7328 ( .A(p_input[277]), .B(n7970), .Z(n7972) );
  XOR U7329 ( .A(n7973), .B(n7974), .Z(n7970) );
  AND U7330 ( .A(n398), .B(n7975), .Z(n7974) );
  IV U7331 ( .A(n7967), .Z(n7969) );
  XOR U7332 ( .A(n7976), .B(n7977), .Z(n7967) );
  AND U7333 ( .A(n402), .B(n7978), .Z(n7977) );
  XOR U7334 ( .A(n7979), .B(n7980), .Z(n7965) );
  AND U7335 ( .A(n406), .B(n7978), .Z(n7980) );
  XNOR U7336 ( .A(n7979), .B(n7976), .Z(n7978) );
  XOR U7337 ( .A(n7981), .B(n7982), .Z(n7976) );
  AND U7338 ( .A(n409), .B(n7975), .Z(n7982) );
  XNOR U7339 ( .A(n7983), .B(n7973), .Z(n7975) );
  XOR U7340 ( .A(n7984), .B(n7985), .Z(n7973) );
  AND U7341 ( .A(n413), .B(n7986), .Z(n7985) );
  XOR U7342 ( .A(p_input[293]), .B(n7984), .Z(n7986) );
  XOR U7343 ( .A(n7987), .B(n7988), .Z(n7984) );
  AND U7344 ( .A(n417), .B(n7989), .Z(n7988) );
  IV U7345 ( .A(n7981), .Z(n7983) );
  XOR U7346 ( .A(n7990), .B(n7991), .Z(n7981) );
  AND U7347 ( .A(n421), .B(n7992), .Z(n7991) );
  XOR U7348 ( .A(n7993), .B(n7994), .Z(n7979) );
  AND U7349 ( .A(n425), .B(n7992), .Z(n7994) );
  XNOR U7350 ( .A(n7993), .B(n7990), .Z(n7992) );
  XOR U7351 ( .A(n7995), .B(n7996), .Z(n7990) );
  AND U7352 ( .A(n428), .B(n7989), .Z(n7996) );
  XNOR U7353 ( .A(n7997), .B(n7987), .Z(n7989) );
  XOR U7354 ( .A(n7998), .B(n7999), .Z(n7987) );
  AND U7355 ( .A(n432), .B(n8000), .Z(n7999) );
  XOR U7356 ( .A(p_input[309]), .B(n7998), .Z(n8000) );
  XOR U7357 ( .A(n8001), .B(n8002), .Z(n7998) );
  AND U7358 ( .A(n436), .B(n8003), .Z(n8002) );
  IV U7359 ( .A(n7995), .Z(n7997) );
  XOR U7360 ( .A(n8004), .B(n8005), .Z(n7995) );
  AND U7361 ( .A(n440), .B(n8006), .Z(n8005) );
  XOR U7362 ( .A(n8007), .B(n8008), .Z(n7993) );
  AND U7363 ( .A(n444), .B(n8006), .Z(n8008) );
  XNOR U7364 ( .A(n8007), .B(n8004), .Z(n8006) );
  XOR U7365 ( .A(n8009), .B(n8010), .Z(n8004) );
  AND U7366 ( .A(n447), .B(n8003), .Z(n8010) );
  XNOR U7367 ( .A(n8011), .B(n8001), .Z(n8003) );
  XOR U7368 ( .A(n8012), .B(n8013), .Z(n8001) );
  AND U7369 ( .A(n451), .B(n8014), .Z(n8013) );
  XOR U7370 ( .A(p_input[325]), .B(n8012), .Z(n8014) );
  XOR U7371 ( .A(n8015), .B(n8016), .Z(n8012) );
  AND U7372 ( .A(n455), .B(n8017), .Z(n8016) );
  IV U7373 ( .A(n8009), .Z(n8011) );
  XOR U7374 ( .A(n8018), .B(n8019), .Z(n8009) );
  AND U7375 ( .A(n459), .B(n8020), .Z(n8019) );
  XOR U7376 ( .A(n8021), .B(n8022), .Z(n8007) );
  AND U7377 ( .A(n463), .B(n8020), .Z(n8022) );
  XNOR U7378 ( .A(n8021), .B(n8018), .Z(n8020) );
  XOR U7379 ( .A(n8023), .B(n8024), .Z(n8018) );
  AND U7380 ( .A(n466), .B(n8017), .Z(n8024) );
  XNOR U7381 ( .A(n8025), .B(n8015), .Z(n8017) );
  XOR U7382 ( .A(n8026), .B(n8027), .Z(n8015) );
  AND U7383 ( .A(n470), .B(n8028), .Z(n8027) );
  XOR U7384 ( .A(p_input[341]), .B(n8026), .Z(n8028) );
  XOR U7385 ( .A(n8029), .B(n8030), .Z(n8026) );
  AND U7386 ( .A(n474), .B(n8031), .Z(n8030) );
  IV U7387 ( .A(n8023), .Z(n8025) );
  XOR U7388 ( .A(n8032), .B(n8033), .Z(n8023) );
  AND U7389 ( .A(n478), .B(n8034), .Z(n8033) );
  XOR U7390 ( .A(n8035), .B(n8036), .Z(n8021) );
  AND U7391 ( .A(n482), .B(n8034), .Z(n8036) );
  XNOR U7392 ( .A(n8035), .B(n8032), .Z(n8034) );
  XOR U7393 ( .A(n8037), .B(n8038), .Z(n8032) );
  AND U7394 ( .A(n485), .B(n8031), .Z(n8038) );
  XNOR U7395 ( .A(n8039), .B(n8029), .Z(n8031) );
  XOR U7396 ( .A(n8040), .B(n8041), .Z(n8029) );
  AND U7397 ( .A(n489), .B(n8042), .Z(n8041) );
  XOR U7398 ( .A(p_input[357]), .B(n8040), .Z(n8042) );
  XOR U7399 ( .A(n8043), .B(n8044), .Z(n8040) );
  AND U7400 ( .A(n493), .B(n8045), .Z(n8044) );
  IV U7401 ( .A(n8037), .Z(n8039) );
  XOR U7402 ( .A(n8046), .B(n8047), .Z(n8037) );
  AND U7403 ( .A(n497), .B(n8048), .Z(n8047) );
  XOR U7404 ( .A(n8049), .B(n8050), .Z(n8035) );
  AND U7405 ( .A(n501), .B(n8048), .Z(n8050) );
  XNOR U7406 ( .A(n8049), .B(n8046), .Z(n8048) );
  XOR U7407 ( .A(n8051), .B(n8052), .Z(n8046) );
  AND U7408 ( .A(n504), .B(n8045), .Z(n8052) );
  XNOR U7409 ( .A(n8053), .B(n8043), .Z(n8045) );
  XOR U7410 ( .A(n8054), .B(n8055), .Z(n8043) );
  AND U7411 ( .A(n508), .B(n8056), .Z(n8055) );
  XOR U7412 ( .A(p_input[373]), .B(n8054), .Z(n8056) );
  XOR U7413 ( .A(n8057), .B(n8058), .Z(n8054) );
  AND U7414 ( .A(n512), .B(n8059), .Z(n8058) );
  IV U7415 ( .A(n8051), .Z(n8053) );
  XOR U7416 ( .A(n8060), .B(n8061), .Z(n8051) );
  AND U7417 ( .A(n516), .B(n8062), .Z(n8061) );
  XOR U7418 ( .A(n8063), .B(n8064), .Z(n8049) );
  AND U7419 ( .A(n520), .B(n8062), .Z(n8064) );
  XNOR U7420 ( .A(n8063), .B(n8060), .Z(n8062) );
  XOR U7421 ( .A(n8065), .B(n8066), .Z(n8060) );
  AND U7422 ( .A(n523), .B(n8059), .Z(n8066) );
  XNOR U7423 ( .A(n8067), .B(n8057), .Z(n8059) );
  XOR U7424 ( .A(n8068), .B(n8069), .Z(n8057) );
  AND U7425 ( .A(n527), .B(n8070), .Z(n8069) );
  XOR U7426 ( .A(p_input[389]), .B(n8068), .Z(n8070) );
  XOR U7427 ( .A(n8071), .B(n8072), .Z(n8068) );
  AND U7428 ( .A(n531), .B(n8073), .Z(n8072) );
  IV U7429 ( .A(n8065), .Z(n8067) );
  XOR U7430 ( .A(n8074), .B(n8075), .Z(n8065) );
  AND U7431 ( .A(n535), .B(n8076), .Z(n8075) );
  XOR U7432 ( .A(n8077), .B(n8078), .Z(n8063) );
  AND U7433 ( .A(n539), .B(n8076), .Z(n8078) );
  XNOR U7434 ( .A(n8077), .B(n8074), .Z(n8076) );
  XOR U7435 ( .A(n8079), .B(n8080), .Z(n8074) );
  AND U7436 ( .A(n542), .B(n8073), .Z(n8080) );
  XNOR U7437 ( .A(n8081), .B(n8071), .Z(n8073) );
  XOR U7438 ( .A(n8082), .B(n8083), .Z(n8071) );
  AND U7439 ( .A(n546), .B(n8084), .Z(n8083) );
  XOR U7440 ( .A(p_input[405]), .B(n8082), .Z(n8084) );
  XOR U7441 ( .A(n8085), .B(n8086), .Z(n8082) );
  AND U7442 ( .A(n550), .B(n8087), .Z(n8086) );
  IV U7443 ( .A(n8079), .Z(n8081) );
  XOR U7444 ( .A(n8088), .B(n8089), .Z(n8079) );
  AND U7445 ( .A(n554), .B(n8090), .Z(n8089) );
  XOR U7446 ( .A(n8091), .B(n8092), .Z(n8077) );
  AND U7447 ( .A(n558), .B(n8090), .Z(n8092) );
  XNOR U7448 ( .A(n8091), .B(n8088), .Z(n8090) );
  XOR U7449 ( .A(n8093), .B(n8094), .Z(n8088) );
  AND U7450 ( .A(n561), .B(n8087), .Z(n8094) );
  XNOR U7451 ( .A(n8095), .B(n8085), .Z(n8087) );
  XOR U7452 ( .A(n8096), .B(n8097), .Z(n8085) );
  AND U7453 ( .A(n565), .B(n8098), .Z(n8097) );
  XOR U7454 ( .A(p_input[421]), .B(n8096), .Z(n8098) );
  XOR U7455 ( .A(n8099), .B(n8100), .Z(n8096) );
  AND U7456 ( .A(n569), .B(n8101), .Z(n8100) );
  IV U7457 ( .A(n8093), .Z(n8095) );
  XOR U7458 ( .A(n8102), .B(n8103), .Z(n8093) );
  AND U7459 ( .A(n573), .B(n8104), .Z(n8103) );
  XOR U7460 ( .A(n8105), .B(n8106), .Z(n8091) );
  AND U7461 ( .A(n577), .B(n8104), .Z(n8106) );
  XNOR U7462 ( .A(n8105), .B(n8102), .Z(n8104) );
  XOR U7463 ( .A(n8107), .B(n8108), .Z(n8102) );
  AND U7464 ( .A(n580), .B(n8101), .Z(n8108) );
  XNOR U7465 ( .A(n8109), .B(n8099), .Z(n8101) );
  XOR U7466 ( .A(n8110), .B(n8111), .Z(n8099) );
  AND U7467 ( .A(n584), .B(n8112), .Z(n8111) );
  XOR U7468 ( .A(p_input[437]), .B(n8110), .Z(n8112) );
  XOR U7469 ( .A(n8113), .B(n8114), .Z(n8110) );
  AND U7470 ( .A(n588), .B(n8115), .Z(n8114) );
  IV U7471 ( .A(n8107), .Z(n8109) );
  XOR U7472 ( .A(n8116), .B(n8117), .Z(n8107) );
  AND U7473 ( .A(n592), .B(n8118), .Z(n8117) );
  XOR U7474 ( .A(n8119), .B(n8120), .Z(n8105) );
  AND U7475 ( .A(n596), .B(n8118), .Z(n8120) );
  XNOR U7476 ( .A(n8119), .B(n8116), .Z(n8118) );
  XOR U7477 ( .A(n8121), .B(n8122), .Z(n8116) );
  AND U7478 ( .A(n599), .B(n8115), .Z(n8122) );
  XNOR U7479 ( .A(n8123), .B(n8113), .Z(n8115) );
  XOR U7480 ( .A(n8124), .B(n8125), .Z(n8113) );
  AND U7481 ( .A(n603), .B(n8126), .Z(n8125) );
  XOR U7482 ( .A(p_input[453]), .B(n8124), .Z(n8126) );
  XOR U7483 ( .A(n8127), .B(n8128), .Z(n8124) );
  AND U7484 ( .A(n607), .B(n8129), .Z(n8128) );
  IV U7485 ( .A(n8121), .Z(n8123) );
  XOR U7486 ( .A(n8130), .B(n8131), .Z(n8121) );
  AND U7487 ( .A(n611), .B(n8132), .Z(n8131) );
  XOR U7488 ( .A(n8133), .B(n8134), .Z(n8119) );
  AND U7489 ( .A(n615), .B(n8132), .Z(n8134) );
  XNOR U7490 ( .A(n8133), .B(n8130), .Z(n8132) );
  XOR U7491 ( .A(n8135), .B(n8136), .Z(n8130) );
  AND U7492 ( .A(n618), .B(n8129), .Z(n8136) );
  XNOR U7493 ( .A(n8137), .B(n8127), .Z(n8129) );
  XOR U7494 ( .A(n8138), .B(n8139), .Z(n8127) );
  AND U7495 ( .A(n622), .B(n8140), .Z(n8139) );
  XOR U7496 ( .A(p_input[469]), .B(n8138), .Z(n8140) );
  XOR U7497 ( .A(n8141), .B(n8142), .Z(n8138) );
  AND U7498 ( .A(n626), .B(n8143), .Z(n8142) );
  IV U7499 ( .A(n8135), .Z(n8137) );
  XOR U7500 ( .A(n8144), .B(n8145), .Z(n8135) );
  AND U7501 ( .A(n630), .B(n8146), .Z(n8145) );
  XOR U7502 ( .A(n8147), .B(n8148), .Z(n8133) );
  AND U7503 ( .A(n634), .B(n8146), .Z(n8148) );
  XNOR U7504 ( .A(n8147), .B(n8144), .Z(n8146) );
  XOR U7505 ( .A(n8149), .B(n8150), .Z(n8144) );
  AND U7506 ( .A(n637), .B(n8143), .Z(n8150) );
  XNOR U7507 ( .A(n8151), .B(n8141), .Z(n8143) );
  XOR U7508 ( .A(n8152), .B(n8153), .Z(n8141) );
  AND U7509 ( .A(n641), .B(n8154), .Z(n8153) );
  XOR U7510 ( .A(p_input[485]), .B(n8152), .Z(n8154) );
  XOR U7511 ( .A(n8155), .B(n8156), .Z(n8152) );
  AND U7512 ( .A(n645), .B(n8157), .Z(n8156) );
  IV U7513 ( .A(n8149), .Z(n8151) );
  XOR U7514 ( .A(n8158), .B(n8159), .Z(n8149) );
  AND U7515 ( .A(n649), .B(n8160), .Z(n8159) );
  XOR U7516 ( .A(n8161), .B(n8162), .Z(n8147) );
  AND U7517 ( .A(n653), .B(n8160), .Z(n8162) );
  XNOR U7518 ( .A(n8161), .B(n8158), .Z(n8160) );
  XOR U7519 ( .A(n8163), .B(n8164), .Z(n8158) );
  AND U7520 ( .A(n656), .B(n8157), .Z(n8164) );
  XNOR U7521 ( .A(n8165), .B(n8155), .Z(n8157) );
  XOR U7522 ( .A(n8166), .B(n8167), .Z(n8155) );
  AND U7523 ( .A(n660), .B(n8168), .Z(n8167) );
  XOR U7524 ( .A(p_input[501]), .B(n8166), .Z(n8168) );
  XOR U7525 ( .A(n8169), .B(n8170), .Z(n8166) );
  AND U7526 ( .A(n664), .B(n8171), .Z(n8170) );
  IV U7527 ( .A(n8163), .Z(n8165) );
  XOR U7528 ( .A(n8172), .B(n8173), .Z(n8163) );
  AND U7529 ( .A(n668), .B(n8174), .Z(n8173) );
  XOR U7530 ( .A(n8175), .B(n8176), .Z(n8161) );
  AND U7531 ( .A(n672), .B(n8174), .Z(n8176) );
  XNOR U7532 ( .A(n8175), .B(n8172), .Z(n8174) );
  XOR U7533 ( .A(n8177), .B(n8178), .Z(n8172) );
  AND U7534 ( .A(n675), .B(n8171), .Z(n8178) );
  XNOR U7535 ( .A(n8179), .B(n8169), .Z(n8171) );
  XOR U7536 ( .A(n8180), .B(n8181), .Z(n8169) );
  AND U7537 ( .A(n679), .B(n8182), .Z(n8181) );
  XOR U7538 ( .A(p_input[517]), .B(n8180), .Z(n8182) );
  XOR U7539 ( .A(n8183), .B(n8184), .Z(n8180) );
  AND U7540 ( .A(n683), .B(n8185), .Z(n8184) );
  IV U7541 ( .A(n8177), .Z(n8179) );
  XOR U7542 ( .A(n8186), .B(n8187), .Z(n8177) );
  AND U7543 ( .A(n687), .B(n8188), .Z(n8187) );
  XOR U7544 ( .A(n8189), .B(n8190), .Z(n8175) );
  AND U7545 ( .A(n691), .B(n8188), .Z(n8190) );
  XNOR U7546 ( .A(n8189), .B(n8186), .Z(n8188) );
  XOR U7547 ( .A(n8191), .B(n8192), .Z(n8186) );
  AND U7548 ( .A(n694), .B(n8185), .Z(n8192) );
  XNOR U7549 ( .A(n8193), .B(n8183), .Z(n8185) );
  XOR U7550 ( .A(n8194), .B(n8195), .Z(n8183) );
  AND U7551 ( .A(n698), .B(n8196), .Z(n8195) );
  XOR U7552 ( .A(p_input[533]), .B(n8194), .Z(n8196) );
  XOR U7553 ( .A(n8197), .B(n8198), .Z(n8194) );
  AND U7554 ( .A(n702), .B(n8199), .Z(n8198) );
  IV U7555 ( .A(n8191), .Z(n8193) );
  XOR U7556 ( .A(n8200), .B(n8201), .Z(n8191) );
  AND U7557 ( .A(n706), .B(n8202), .Z(n8201) );
  XOR U7558 ( .A(n8203), .B(n8204), .Z(n8189) );
  AND U7559 ( .A(n710), .B(n8202), .Z(n8204) );
  XNOR U7560 ( .A(n8203), .B(n8200), .Z(n8202) );
  XOR U7561 ( .A(n8205), .B(n8206), .Z(n8200) );
  AND U7562 ( .A(n713), .B(n8199), .Z(n8206) );
  XNOR U7563 ( .A(n8207), .B(n8197), .Z(n8199) );
  XOR U7564 ( .A(n8208), .B(n8209), .Z(n8197) );
  AND U7565 ( .A(n717), .B(n8210), .Z(n8209) );
  XOR U7566 ( .A(p_input[549]), .B(n8208), .Z(n8210) );
  XOR U7567 ( .A(n8211), .B(n8212), .Z(n8208) );
  AND U7568 ( .A(n721), .B(n8213), .Z(n8212) );
  IV U7569 ( .A(n8205), .Z(n8207) );
  XOR U7570 ( .A(n8214), .B(n8215), .Z(n8205) );
  AND U7571 ( .A(n725), .B(n8216), .Z(n8215) );
  XOR U7572 ( .A(n8217), .B(n8218), .Z(n8203) );
  AND U7573 ( .A(n729), .B(n8216), .Z(n8218) );
  XNOR U7574 ( .A(n8217), .B(n8214), .Z(n8216) );
  XOR U7575 ( .A(n8219), .B(n8220), .Z(n8214) );
  AND U7576 ( .A(n732), .B(n8213), .Z(n8220) );
  XNOR U7577 ( .A(n8221), .B(n8211), .Z(n8213) );
  XOR U7578 ( .A(n8222), .B(n8223), .Z(n8211) );
  AND U7579 ( .A(n736), .B(n8224), .Z(n8223) );
  XOR U7580 ( .A(p_input[565]), .B(n8222), .Z(n8224) );
  XOR U7581 ( .A(n8225), .B(n8226), .Z(n8222) );
  AND U7582 ( .A(n740), .B(n8227), .Z(n8226) );
  IV U7583 ( .A(n8219), .Z(n8221) );
  XOR U7584 ( .A(n8228), .B(n8229), .Z(n8219) );
  AND U7585 ( .A(n744), .B(n8230), .Z(n8229) );
  XOR U7586 ( .A(n8231), .B(n8232), .Z(n8217) );
  AND U7587 ( .A(n748), .B(n8230), .Z(n8232) );
  XNOR U7588 ( .A(n8231), .B(n8228), .Z(n8230) );
  XOR U7589 ( .A(n8233), .B(n8234), .Z(n8228) );
  AND U7590 ( .A(n751), .B(n8227), .Z(n8234) );
  XNOR U7591 ( .A(n8235), .B(n8225), .Z(n8227) );
  XOR U7592 ( .A(n8236), .B(n8237), .Z(n8225) );
  AND U7593 ( .A(n755), .B(n8238), .Z(n8237) );
  XOR U7594 ( .A(p_input[581]), .B(n8236), .Z(n8238) );
  XOR U7595 ( .A(n8239), .B(n8240), .Z(n8236) );
  AND U7596 ( .A(n759), .B(n8241), .Z(n8240) );
  IV U7597 ( .A(n8233), .Z(n8235) );
  XOR U7598 ( .A(n8242), .B(n8243), .Z(n8233) );
  AND U7599 ( .A(n763), .B(n8244), .Z(n8243) );
  XOR U7600 ( .A(n8245), .B(n8246), .Z(n8231) );
  AND U7601 ( .A(n767), .B(n8244), .Z(n8246) );
  XNOR U7602 ( .A(n8245), .B(n8242), .Z(n8244) );
  XOR U7603 ( .A(n8247), .B(n8248), .Z(n8242) );
  AND U7604 ( .A(n770), .B(n8241), .Z(n8248) );
  XNOR U7605 ( .A(n8249), .B(n8239), .Z(n8241) );
  XOR U7606 ( .A(n8250), .B(n8251), .Z(n8239) );
  AND U7607 ( .A(n774), .B(n8252), .Z(n8251) );
  XOR U7608 ( .A(p_input[597]), .B(n8250), .Z(n8252) );
  XOR U7609 ( .A(n8253), .B(n8254), .Z(n8250) );
  AND U7610 ( .A(n778), .B(n8255), .Z(n8254) );
  IV U7611 ( .A(n8247), .Z(n8249) );
  XOR U7612 ( .A(n8256), .B(n8257), .Z(n8247) );
  AND U7613 ( .A(n782), .B(n8258), .Z(n8257) );
  XOR U7614 ( .A(n8259), .B(n8260), .Z(n8245) );
  AND U7615 ( .A(n786), .B(n8258), .Z(n8260) );
  XNOR U7616 ( .A(n8259), .B(n8256), .Z(n8258) );
  XOR U7617 ( .A(n8261), .B(n8262), .Z(n8256) );
  AND U7618 ( .A(n789), .B(n8255), .Z(n8262) );
  XNOR U7619 ( .A(n8263), .B(n8253), .Z(n8255) );
  XOR U7620 ( .A(n8264), .B(n8265), .Z(n8253) );
  AND U7621 ( .A(n793), .B(n8266), .Z(n8265) );
  XOR U7622 ( .A(p_input[613]), .B(n8264), .Z(n8266) );
  XOR U7623 ( .A(n8267), .B(n8268), .Z(n8264) );
  AND U7624 ( .A(n797), .B(n8269), .Z(n8268) );
  IV U7625 ( .A(n8261), .Z(n8263) );
  XOR U7626 ( .A(n8270), .B(n8271), .Z(n8261) );
  AND U7627 ( .A(n801), .B(n8272), .Z(n8271) );
  XOR U7628 ( .A(n8273), .B(n8274), .Z(n8259) );
  AND U7629 ( .A(n805), .B(n8272), .Z(n8274) );
  XNOR U7630 ( .A(n8273), .B(n8270), .Z(n8272) );
  XOR U7631 ( .A(n8275), .B(n8276), .Z(n8270) );
  AND U7632 ( .A(n808), .B(n8269), .Z(n8276) );
  XNOR U7633 ( .A(n8277), .B(n8267), .Z(n8269) );
  XOR U7634 ( .A(n8278), .B(n8279), .Z(n8267) );
  AND U7635 ( .A(n812), .B(n8280), .Z(n8279) );
  XOR U7636 ( .A(p_input[629]), .B(n8278), .Z(n8280) );
  XOR U7637 ( .A(n8281), .B(n8282), .Z(n8278) );
  AND U7638 ( .A(n816), .B(n8283), .Z(n8282) );
  IV U7639 ( .A(n8275), .Z(n8277) );
  XOR U7640 ( .A(n8284), .B(n8285), .Z(n8275) );
  AND U7641 ( .A(n820), .B(n8286), .Z(n8285) );
  XOR U7642 ( .A(n8287), .B(n8288), .Z(n8273) );
  AND U7643 ( .A(n824), .B(n8286), .Z(n8288) );
  XNOR U7644 ( .A(n8287), .B(n8284), .Z(n8286) );
  XOR U7645 ( .A(n8289), .B(n8290), .Z(n8284) );
  AND U7646 ( .A(n827), .B(n8283), .Z(n8290) );
  XNOR U7647 ( .A(n8291), .B(n8281), .Z(n8283) );
  XOR U7648 ( .A(n8292), .B(n8293), .Z(n8281) );
  AND U7649 ( .A(n831), .B(n8294), .Z(n8293) );
  XOR U7650 ( .A(p_input[645]), .B(n8292), .Z(n8294) );
  XOR U7651 ( .A(n8295), .B(n8296), .Z(n8292) );
  AND U7652 ( .A(n835), .B(n8297), .Z(n8296) );
  IV U7653 ( .A(n8289), .Z(n8291) );
  XOR U7654 ( .A(n8298), .B(n8299), .Z(n8289) );
  AND U7655 ( .A(n839), .B(n8300), .Z(n8299) );
  XOR U7656 ( .A(n8301), .B(n8302), .Z(n8287) );
  AND U7657 ( .A(n843), .B(n8300), .Z(n8302) );
  XNOR U7658 ( .A(n8301), .B(n8298), .Z(n8300) );
  XOR U7659 ( .A(n8303), .B(n8304), .Z(n8298) );
  AND U7660 ( .A(n846), .B(n8297), .Z(n8304) );
  XNOR U7661 ( .A(n8305), .B(n8295), .Z(n8297) );
  XOR U7662 ( .A(n8306), .B(n8307), .Z(n8295) );
  AND U7663 ( .A(n850), .B(n8308), .Z(n8307) );
  XOR U7664 ( .A(p_input[661]), .B(n8306), .Z(n8308) );
  XOR U7665 ( .A(n8309), .B(n8310), .Z(n8306) );
  AND U7666 ( .A(n854), .B(n8311), .Z(n8310) );
  IV U7667 ( .A(n8303), .Z(n8305) );
  XOR U7668 ( .A(n8312), .B(n8313), .Z(n8303) );
  AND U7669 ( .A(n858), .B(n8314), .Z(n8313) );
  XOR U7670 ( .A(n8315), .B(n8316), .Z(n8301) );
  AND U7671 ( .A(n862), .B(n8314), .Z(n8316) );
  XNOR U7672 ( .A(n8315), .B(n8312), .Z(n8314) );
  XOR U7673 ( .A(n8317), .B(n8318), .Z(n8312) );
  AND U7674 ( .A(n865), .B(n8311), .Z(n8318) );
  XNOR U7675 ( .A(n8319), .B(n8309), .Z(n8311) );
  XOR U7676 ( .A(n8320), .B(n8321), .Z(n8309) );
  AND U7677 ( .A(n869), .B(n8322), .Z(n8321) );
  XOR U7678 ( .A(p_input[677]), .B(n8320), .Z(n8322) );
  XOR U7679 ( .A(n8323), .B(n8324), .Z(n8320) );
  AND U7680 ( .A(n873), .B(n8325), .Z(n8324) );
  IV U7681 ( .A(n8317), .Z(n8319) );
  XOR U7682 ( .A(n8326), .B(n8327), .Z(n8317) );
  AND U7683 ( .A(n877), .B(n8328), .Z(n8327) );
  XOR U7684 ( .A(n8329), .B(n8330), .Z(n8315) );
  AND U7685 ( .A(n881), .B(n8328), .Z(n8330) );
  XNOR U7686 ( .A(n8329), .B(n8326), .Z(n8328) );
  XOR U7687 ( .A(n8331), .B(n8332), .Z(n8326) );
  AND U7688 ( .A(n884), .B(n8325), .Z(n8332) );
  XNOR U7689 ( .A(n8333), .B(n8323), .Z(n8325) );
  XOR U7690 ( .A(n8334), .B(n8335), .Z(n8323) );
  AND U7691 ( .A(n888), .B(n8336), .Z(n8335) );
  XOR U7692 ( .A(p_input[693]), .B(n8334), .Z(n8336) );
  XOR U7693 ( .A(n8337), .B(n8338), .Z(n8334) );
  AND U7694 ( .A(n892), .B(n8339), .Z(n8338) );
  IV U7695 ( .A(n8331), .Z(n8333) );
  XOR U7696 ( .A(n8340), .B(n8341), .Z(n8331) );
  AND U7697 ( .A(n896), .B(n8342), .Z(n8341) );
  XOR U7698 ( .A(n8343), .B(n8344), .Z(n8329) );
  AND U7699 ( .A(n900), .B(n8342), .Z(n8344) );
  XNOR U7700 ( .A(n8343), .B(n8340), .Z(n8342) );
  XOR U7701 ( .A(n8345), .B(n8346), .Z(n8340) );
  AND U7702 ( .A(n903), .B(n8339), .Z(n8346) );
  XNOR U7703 ( .A(n8347), .B(n8337), .Z(n8339) );
  XOR U7704 ( .A(n8348), .B(n8349), .Z(n8337) );
  AND U7705 ( .A(n907), .B(n8350), .Z(n8349) );
  XOR U7706 ( .A(p_input[709]), .B(n8348), .Z(n8350) );
  XOR U7707 ( .A(n8351), .B(n8352), .Z(n8348) );
  AND U7708 ( .A(n911), .B(n8353), .Z(n8352) );
  IV U7709 ( .A(n8345), .Z(n8347) );
  XOR U7710 ( .A(n8354), .B(n8355), .Z(n8345) );
  AND U7711 ( .A(n915), .B(n8356), .Z(n8355) );
  XOR U7712 ( .A(n8357), .B(n8358), .Z(n8343) );
  AND U7713 ( .A(n919), .B(n8356), .Z(n8358) );
  XNOR U7714 ( .A(n8357), .B(n8354), .Z(n8356) );
  XOR U7715 ( .A(n8359), .B(n8360), .Z(n8354) );
  AND U7716 ( .A(n922), .B(n8353), .Z(n8360) );
  XNOR U7717 ( .A(n8361), .B(n8351), .Z(n8353) );
  XOR U7718 ( .A(n8362), .B(n8363), .Z(n8351) );
  AND U7719 ( .A(n926), .B(n8364), .Z(n8363) );
  XOR U7720 ( .A(p_input[725]), .B(n8362), .Z(n8364) );
  XOR U7721 ( .A(n8365), .B(n8366), .Z(n8362) );
  AND U7722 ( .A(n930), .B(n8367), .Z(n8366) );
  IV U7723 ( .A(n8359), .Z(n8361) );
  XOR U7724 ( .A(n8368), .B(n8369), .Z(n8359) );
  AND U7725 ( .A(n934), .B(n8370), .Z(n8369) );
  XOR U7726 ( .A(n8371), .B(n8372), .Z(n8357) );
  AND U7727 ( .A(n938), .B(n8370), .Z(n8372) );
  XNOR U7728 ( .A(n8371), .B(n8368), .Z(n8370) );
  XOR U7729 ( .A(n8373), .B(n8374), .Z(n8368) );
  AND U7730 ( .A(n941), .B(n8367), .Z(n8374) );
  XNOR U7731 ( .A(n8375), .B(n8365), .Z(n8367) );
  XOR U7732 ( .A(n8376), .B(n8377), .Z(n8365) );
  AND U7733 ( .A(n945), .B(n8378), .Z(n8377) );
  XOR U7734 ( .A(p_input[741]), .B(n8376), .Z(n8378) );
  XOR U7735 ( .A(n8379), .B(n8380), .Z(n8376) );
  AND U7736 ( .A(n949), .B(n8381), .Z(n8380) );
  IV U7737 ( .A(n8373), .Z(n8375) );
  XOR U7738 ( .A(n8382), .B(n8383), .Z(n8373) );
  AND U7739 ( .A(n953), .B(n8384), .Z(n8383) );
  XOR U7740 ( .A(n8385), .B(n8386), .Z(n8371) );
  AND U7741 ( .A(n957), .B(n8384), .Z(n8386) );
  XNOR U7742 ( .A(n8385), .B(n8382), .Z(n8384) );
  XOR U7743 ( .A(n8387), .B(n8388), .Z(n8382) );
  AND U7744 ( .A(n960), .B(n8381), .Z(n8388) );
  XNOR U7745 ( .A(n8389), .B(n8379), .Z(n8381) );
  XOR U7746 ( .A(n8390), .B(n8391), .Z(n8379) );
  AND U7747 ( .A(n964), .B(n8392), .Z(n8391) );
  XOR U7748 ( .A(p_input[757]), .B(n8390), .Z(n8392) );
  XOR U7749 ( .A(n8393), .B(n8394), .Z(n8390) );
  AND U7750 ( .A(n968), .B(n8395), .Z(n8394) );
  IV U7751 ( .A(n8387), .Z(n8389) );
  XOR U7752 ( .A(n8396), .B(n8397), .Z(n8387) );
  AND U7753 ( .A(n972), .B(n8398), .Z(n8397) );
  XOR U7754 ( .A(n8399), .B(n8400), .Z(n8385) );
  AND U7755 ( .A(n976), .B(n8398), .Z(n8400) );
  XNOR U7756 ( .A(n8399), .B(n8396), .Z(n8398) );
  XOR U7757 ( .A(n8401), .B(n8402), .Z(n8396) );
  AND U7758 ( .A(n979), .B(n8395), .Z(n8402) );
  XNOR U7759 ( .A(n8403), .B(n8393), .Z(n8395) );
  XOR U7760 ( .A(n8404), .B(n8405), .Z(n8393) );
  AND U7761 ( .A(n983), .B(n8406), .Z(n8405) );
  XOR U7762 ( .A(p_input[773]), .B(n8404), .Z(n8406) );
  XOR U7763 ( .A(n8407), .B(n8408), .Z(n8404) );
  AND U7764 ( .A(n987), .B(n8409), .Z(n8408) );
  IV U7765 ( .A(n8401), .Z(n8403) );
  XOR U7766 ( .A(n8410), .B(n8411), .Z(n8401) );
  AND U7767 ( .A(n991), .B(n8412), .Z(n8411) );
  XOR U7768 ( .A(n8413), .B(n8414), .Z(n8399) );
  AND U7769 ( .A(n995), .B(n8412), .Z(n8414) );
  XNOR U7770 ( .A(n8413), .B(n8410), .Z(n8412) );
  XOR U7771 ( .A(n8415), .B(n8416), .Z(n8410) );
  AND U7772 ( .A(n998), .B(n8409), .Z(n8416) );
  XNOR U7773 ( .A(n8417), .B(n8407), .Z(n8409) );
  XOR U7774 ( .A(n8418), .B(n8419), .Z(n8407) );
  AND U7775 ( .A(n1002), .B(n8420), .Z(n8419) );
  XOR U7776 ( .A(p_input[789]), .B(n8418), .Z(n8420) );
  XOR U7777 ( .A(n8421), .B(n8422), .Z(n8418) );
  AND U7778 ( .A(n1006), .B(n8423), .Z(n8422) );
  IV U7779 ( .A(n8415), .Z(n8417) );
  XOR U7780 ( .A(n8424), .B(n8425), .Z(n8415) );
  AND U7781 ( .A(n1010), .B(n8426), .Z(n8425) );
  XOR U7782 ( .A(n8427), .B(n8428), .Z(n8413) );
  AND U7783 ( .A(n1014), .B(n8426), .Z(n8428) );
  XNOR U7784 ( .A(n8427), .B(n8424), .Z(n8426) );
  XOR U7785 ( .A(n8429), .B(n8430), .Z(n8424) );
  AND U7786 ( .A(n1017), .B(n8423), .Z(n8430) );
  XNOR U7787 ( .A(n8431), .B(n8421), .Z(n8423) );
  XOR U7788 ( .A(n8432), .B(n8433), .Z(n8421) );
  AND U7789 ( .A(n1021), .B(n8434), .Z(n8433) );
  XOR U7790 ( .A(p_input[805]), .B(n8432), .Z(n8434) );
  XOR U7791 ( .A(n8435), .B(n8436), .Z(n8432) );
  AND U7792 ( .A(n1025), .B(n8437), .Z(n8436) );
  IV U7793 ( .A(n8429), .Z(n8431) );
  XOR U7794 ( .A(n8438), .B(n8439), .Z(n8429) );
  AND U7795 ( .A(n1029), .B(n8440), .Z(n8439) );
  XOR U7796 ( .A(n8441), .B(n8442), .Z(n8427) );
  AND U7797 ( .A(n1033), .B(n8440), .Z(n8442) );
  XNOR U7798 ( .A(n8441), .B(n8438), .Z(n8440) );
  XOR U7799 ( .A(n8443), .B(n8444), .Z(n8438) );
  AND U7800 ( .A(n1036), .B(n8437), .Z(n8444) );
  XNOR U7801 ( .A(n8445), .B(n8435), .Z(n8437) );
  XOR U7802 ( .A(n8446), .B(n8447), .Z(n8435) );
  AND U7803 ( .A(n1040), .B(n8448), .Z(n8447) );
  XOR U7804 ( .A(p_input[821]), .B(n8446), .Z(n8448) );
  XOR U7805 ( .A(n8449), .B(n8450), .Z(n8446) );
  AND U7806 ( .A(n1044), .B(n8451), .Z(n8450) );
  IV U7807 ( .A(n8443), .Z(n8445) );
  XOR U7808 ( .A(n8452), .B(n8453), .Z(n8443) );
  AND U7809 ( .A(n1048), .B(n8454), .Z(n8453) );
  XOR U7810 ( .A(n8455), .B(n8456), .Z(n8441) );
  AND U7811 ( .A(n1052), .B(n8454), .Z(n8456) );
  XNOR U7812 ( .A(n8455), .B(n8452), .Z(n8454) );
  XOR U7813 ( .A(n8457), .B(n8458), .Z(n8452) );
  AND U7814 ( .A(n1055), .B(n8451), .Z(n8458) );
  XNOR U7815 ( .A(n8459), .B(n8449), .Z(n8451) );
  XOR U7816 ( .A(n8460), .B(n8461), .Z(n8449) );
  AND U7817 ( .A(n1059), .B(n8462), .Z(n8461) );
  XOR U7818 ( .A(p_input[837]), .B(n8460), .Z(n8462) );
  XOR U7819 ( .A(n8463), .B(n8464), .Z(n8460) );
  AND U7820 ( .A(n1063), .B(n8465), .Z(n8464) );
  IV U7821 ( .A(n8457), .Z(n8459) );
  XOR U7822 ( .A(n8466), .B(n8467), .Z(n8457) );
  AND U7823 ( .A(n1067), .B(n8468), .Z(n8467) );
  XOR U7824 ( .A(n8469), .B(n8470), .Z(n8455) );
  AND U7825 ( .A(n1071), .B(n8468), .Z(n8470) );
  XNOR U7826 ( .A(n8469), .B(n8466), .Z(n8468) );
  XOR U7827 ( .A(n8471), .B(n8472), .Z(n8466) );
  AND U7828 ( .A(n1074), .B(n8465), .Z(n8472) );
  XNOR U7829 ( .A(n8473), .B(n8463), .Z(n8465) );
  XOR U7830 ( .A(n8474), .B(n8475), .Z(n8463) );
  AND U7831 ( .A(n1078), .B(n8476), .Z(n8475) );
  XOR U7832 ( .A(p_input[853]), .B(n8474), .Z(n8476) );
  XOR U7833 ( .A(n8477), .B(n8478), .Z(n8474) );
  AND U7834 ( .A(n1082), .B(n8479), .Z(n8478) );
  IV U7835 ( .A(n8471), .Z(n8473) );
  XOR U7836 ( .A(n8480), .B(n8481), .Z(n8471) );
  AND U7837 ( .A(n1086), .B(n8482), .Z(n8481) );
  XOR U7838 ( .A(n8483), .B(n8484), .Z(n8469) );
  AND U7839 ( .A(n1090), .B(n8482), .Z(n8484) );
  XNOR U7840 ( .A(n8483), .B(n8480), .Z(n8482) );
  XOR U7841 ( .A(n8485), .B(n8486), .Z(n8480) );
  AND U7842 ( .A(n1093), .B(n8479), .Z(n8486) );
  XNOR U7843 ( .A(n8487), .B(n8477), .Z(n8479) );
  XOR U7844 ( .A(n8488), .B(n8489), .Z(n8477) );
  AND U7845 ( .A(n1097), .B(n8490), .Z(n8489) );
  XOR U7846 ( .A(p_input[869]), .B(n8488), .Z(n8490) );
  XOR U7847 ( .A(n8491), .B(n8492), .Z(n8488) );
  AND U7848 ( .A(n1101), .B(n8493), .Z(n8492) );
  IV U7849 ( .A(n8485), .Z(n8487) );
  XOR U7850 ( .A(n8494), .B(n8495), .Z(n8485) );
  AND U7851 ( .A(n1105), .B(n8496), .Z(n8495) );
  XOR U7852 ( .A(n8497), .B(n8498), .Z(n8483) );
  AND U7853 ( .A(n1109), .B(n8496), .Z(n8498) );
  XNOR U7854 ( .A(n8497), .B(n8494), .Z(n8496) );
  XOR U7855 ( .A(n8499), .B(n8500), .Z(n8494) );
  AND U7856 ( .A(n1112), .B(n8493), .Z(n8500) );
  XNOR U7857 ( .A(n8501), .B(n8491), .Z(n8493) );
  XOR U7858 ( .A(n8502), .B(n8503), .Z(n8491) );
  AND U7859 ( .A(n1116), .B(n8504), .Z(n8503) );
  XOR U7860 ( .A(p_input[885]), .B(n8502), .Z(n8504) );
  XOR U7861 ( .A(n8505), .B(n8506), .Z(n8502) );
  AND U7862 ( .A(n1120), .B(n8507), .Z(n8506) );
  IV U7863 ( .A(n8499), .Z(n8501) );
  XOR U7864 ( .A(n8508), .B(n8509), .Z(n8499) );
  AND U7865 ( .A(n1124), .B(n8510), .Z(n8509) );
  XOR U7866 ( .A(n8511), .B(n8512), .Z(n8497) );
  AND U7867 ( .A(n1128), .B(n8510), .Z(n8512) );
  XNOR U7868 ( .A(n8511), .B(n8508), .Z(n8510) );
  XOR U7869 ( .A(n8513), .B(n8514), .Z(n8508) );
  AND U7870 ( .A(n1131), .B(n8507), .Z(n8514) );
  XNOR U7871 ( .A(n8515), .B(n8505), .Z(n8507) );
  XOR U7872 ( .A(n8516), .B(n8517), .Z(n8505) );
  AND U7873 ( .A(n1135), .B(n8518), .Z(n8517) );
  XOR U7874 ( .A(p_input[901]), .B(n8516), .Z(n8518) );
  XOR U7875 ( .A(n8519), .B(n8520), .Z(n8516) );
  AND U7876 ( .A(n1139), .B(n8521), .Z(n8520) );
  IV U7877 ( .A(n8513), .Z(n8515) );
  XOR U7878 ( .A(n8522), .B(n8523), .Z(n8513) );
  AND U7879 ( .A(n1143), .B(n8524), .Z(n8523) );
  XOR U7880 ( .A(n8525), .B(n8526), .Z(n8511) );
  AND U7881 ( .A(n1147), .B(n8524), .Z(n8526) );
  XNOR U7882 ( .A(n8525), .B(n8522), .Z(n8524) );
  XOR U7883 ( .A(n8527), .B(n8528), .Z(n8522) );
  AND U7884 ( .A(n1150), .B(n8521), .Z(n8528) );
  XNOR U7885 ( .A(n8529), .B(n8519), .Z(n8521) );
  XOR U7886 ( .A(n8530), .B(n8531), .Z(n8519) );
  AND U7887 ( .A(n1154), .B(n8532), .Z(n8531) );
  XOR U7888 ( .A(p_input[917]), .B(n8530), .Z(n8532) );
  XOR U7889 ( .A(n8533), .B(n8534), .Z(n8530) );
  AND U7890 ( .A(n1158), .B(n8535), .Z(n8534) );
  IV U7891 ( .A(n8527), .Z(n8529) );
  XOR U7892 ( .A(n8536), .B(n8537), .Z(n8527) );
  AND U7893 ( .A(n1162), .B(n8538), .Z(n8537) );
  XOR U7894 ( .A(n8539), .B(n8540), .Z(n8525) );
  AND U7895 ( .A(n1166), .B(n8538), .Z(n8540) );
  XNOR U7896 ( .A(n8539), .B(n8536), .Z(n8538) );
  XOR U7897 ( .A(n8541), .B(n8542), .Z(n8536) );
  AND U7898 ( .A(n1169), .B(n8535), .Z(n8542) );
  XNOR U7899 ( .A(n8543), .B(n8533), .Z(n8535) );
  XOR U7900 ( .A(n8544), .B(n8545), .Z(n8533) );
  AND U7901 ( .A(n1173), .B(n8546), .Z(n8545) );
  XOR U7902 ( .A(p_input[933]), .B(n8544), .Z(n8546) );
  XOR U7903 ( .A(n8547), .B(n8548), .Z(n8544) );
  AND U7904 ( .A(n1177), .B(n8549), .Z(n8548) );
  IV U7905 ( .A(n8541), .Z(n8543) );
  XOR U7906 ( .A(n8550), .B(n8551), .Z(n8541) );
  AND U7907 ( .A(n1181), .B(n8552), .Z(n8551) );
  XOR U7908 ( .A(n8553), .B(n8554), .Z(n8539) );
  AND U7909 ( .A(n1185), .B(n8552), .Z(n8554) );
  XNOR U7910 ( .A(n8553), .B(n8550), .Z(n8552) );
  XOR U7911 ( .A(n8555), .B(n8556), .Z(n8550) );
  AND U7912 ( .A(n1188), .B(n8549), .Z(n8556) );
  XNOR U7913 ( .A(n8557), .B(n8547), .Z(n8549) );
  XOR U7914 ( .A(n8558), .B(n8559), .Z(n8547) );
  AND U7915 ( .A(n1192), .B(n8560), .Z(n8559) );
  XOR U7916 ( .A(p_input[949]), .B(n8558), .Z(n8560) );
  XOR U7917 ( .A(n8561), .B(n8562), .Z(n8558) );
  AND U7918 ( .A(n1196), .B(n8563), .Z(n8562) );
  IV U7919 ( .A(n8555), .Z(n8557) );
  XOR U7920 ( .A(n8564), .B(n8565), .Z(n8555) );
  AND U7921 ( .A(n1200), .B(n8566), .Z(n8565) );
  XOR U7922 ( .A(n8567), .B(n8568), .Z(n8553) );
  AND U7923 ( .A(n1204), .B(n8566), .Z(n8568) );
  XNOR U7924 ( .A(n8567), .B(n8564), .Z(n8566) );
  XOR U7925 ( .A(n8569), .B(n8570), .Z(n8564) );
  AND U7926 ( .A(n1207), .B(n8563), .Z(n8570) );
  XNOR U7927 ( .A(n8571), .B(n8561), .Z(n8563) );
  XOR U7928 ( .A(n8572), .B(n8573), .Z(n8561) );
  AND U7929 ( .A(n1211), .B(n8574), .Z(n8573) );
  XOR U7930 ( .A(p_input[965]), .B(n8572), .Z(n8574) );
  XOR U7931 ( .A(n8575), .B(n8576), .Z(n8572) );
  AND U7932 ( .A(n1215), .B(n8577), .Z(n8576) );
  IV U7933 ( .A(n8569), .Z(n8571) );
  XOR U7934 ( .A(n8578), .B(n8579), .Z(n8569) );
  AND U7935 ( .A(n1219), .B(n8580), .Z(n8579) );
  XOR U7936 ( .A(n8581), .B(n8582), .Z(n8567) );
  AND U7937 ( .A(n1223), .B(n8580), .Z(n8582) );
  XNOR U7938 ( .A(n8581), .B(n8578), .Z(n8580) );
  XOR U7939 ( .A(n8583), .B(n8584), .Z(n8578) );
  AND U7940 ( .A(n1226), .B(n8577), .Z(n8584) );
  XNOR U7941 ( .A(n8585), .B(n8575), .Z(n8577) );
  XOR U7942 ( .A(n8586), .B(n8587), .Z(n8575) );
  AND U7943 ( .A(n1230), .B(n8588), .Z(n8587) );
  XOR U7944 ( .A(p_input[981]), .B(n8586), .Z(n8588) );
  XOR U7945 ( .A(n8589), .B(n8590), .Z(n8586) );
  AND U7946 ( .A(n1234), .B(n8591), .Z(n8590) );
  IV U7947 ( .A(n8583), .Z(n8585) );
  XOR U7948 ( .A(n8592), .B(n8593), .Z(n8583) );
  AND U7949 ( .A(n1238), .B(n8594), .Z(n8593) );
  XOR U7950 ( .A(n8595), .B(n8596), .Z(n8581) );
  AND U7951 ( .A(n1242), .B(n8594), .Z(n8596) );
  XNOR U7952 ( .A(n8595), .B(n8592), .Z(n8594) );
  XOR U7953 ( .A(n8597), .B(n8598), .Z(n8592) );
  AND U7954 ( .A(n1245), .B(n8591), .Z(n8598) );
  XNOR U7955 ( .A(n8599), .B(n8589), .Z(n8591) );
  XOR U7956 ( .A(n8600), .B(n8601), .Z(n8589) );
  AND U7957 ( .A(n1249), .B(n8602), .Z(n8601) );
  XOR U7958 ( .A(p_input[997]), .B(n8600), .Z(n8602) );
  XOR U7959 ( .A(n8603), .B(n8604), .Z(n8600) );
  AND U7960 ( .A(n1253), .B(n8605), .Z(n8604) );
  IV U7961 ( .A(n8597), .Z(n8599) );
  XOR U7962 ( .A(n8606), .B(n8607), .Z(n8597) );
  AND U7963 ( .A(n1257), .B(n8608), .Z(n8607) );
  XOR U7964 ( .A(n8609), .B(n8610), .Z(n8595) );
  AND U7965 ( .A(n1261), .B(n8608), .Z(n8610) );
  XNOR U7966 ( .A(n8609), .B(n8606), .Z(n8608) );
  XOR U7967 ( .A(n8611), .B(n8612), .Z(n8606) );
  AND U7968 ( .A(n1264), .B(n8605), .Z(n8612) );
  XNOR U7969 ( .A(n8613), .B(n8603), .Z(n8605) );
  XOR U7970 ( .A(n8614), .B(n8615), .Z(n8603) );
  AND U7971 ( .A(n1268), .B(n8616), .Z(n8615) );
  XOR U7972 ( .A(p_input[1013]), .B(n8614), .Z(n8616) );
  XOR U7973 ( .A(n8617), .B(n8618), .Z(n8614) );
  AND U7974 ( .A(n1272), .B(n8619), .Z(n8618) );
  IV U7975 ( .A(n8611), .Z(n8613) );
  XOR U7976 ( .A(n8620), .B(n8621), .Z(n8611) );
  AND U7977 ( .A(n1276), .B(n8622), .Z(n8621) );
  XOR U7978 ( .A(n8623), .B(n8624), .Z(n8609) );
  AND U7979 ( .A(n1280), .B(n8622), .Z(n8624) );
  XNOR U7980 ( .A(n8623), .B(n8620), .Z(n8622) );
  XOR U7981 ( .A(n8625), .B(n8626), .Z(n8620) );
  AND U7982 ( .A(n1283), .B(n8619), .Z(n8626) );
  XNOR U7983 ( .A(n8627), .B(n8617), .Z(n8619) );
  XOR U7984 ( .A(n8628), .B(n8629), .Z(n8617) );
  AND U7985 ( .A(n1287), .B(n8630), .Z(n8629) );
  XOR U7986 ( .A(p_input[1029]), .B(n8628), .Z(n8630) );
  XOR U7987 ( .A(n8631), .B(n8632), .Z(n8628) );
  AND U7988 ( .A(n1291), .B(n8633), .Z(n8632) );
  IV U7989 ( .A(n8625), .Z(n8627) );
  XOR U7990 ( .A(n8634), .B(n8635), .Z(n8625) );
  AND U7991 ( .A(n1295), .B(n8636), .Z(n8635) );
  XOR U7992 ( .A(n8637), .B(n8638), .Z(n8623) );
  AND U7993 ( .A(n1299), .B(n8636), .Z(n8638) );
  XNOR U7994 ( .A(n8637), .B(n8634), .Z(n8636) );
  XOR U7995 ( .A(n8639), .B(n8640), .Z(n8634) );
  AND U7996 ( .A(n1302), .B(n8633), .Z(n8640) );
  XNOR U7997 ( .A(n8641), .B(n8631), .Z(n8633) );
  XOR U7998 ( .A(n8642), .B(n8643), .Z(n8631) );
  AND U7999 ( .A(n1306), .B(n8644), .Z(n8643) );
  XOR U8000 ( .A(p_input[1045]), .B(n8642), .Z(n8644) );
  XOR U8001 ( .A(n8645), .B(n8646), .Z(n8642) );
  AND U8002 ( .A(n1310), .B(n8647), .Z(n8646) );
  IV U8003 ( .A(n8639), .Z(n8641) );
  XOR U8004 ( .A(n8648), .B(n8649), .Z(n8639) );
  AND U8005 ( .A(n1314), .B(n8650), .Z(n8649) );
  XOR U8006 ( .A(n8651), .B(n8652), .Z(n8637) );
  AND U8007 ( .A(n1318), .B(n8650), .Z(n8652) );
  XNOR U8008 ( .A(n8651), .B(n8648), .Z(n8650) );
  XOR U8009 ( .A(n8653), .B(n8654), .Z(n8648) );
  AND U8010 ( .A(n1321), .B(n8647), .Z(n8654) );
  XNOR U8011 ( .A(n8655), .B(n8645), .Z(n8647) );
  XOR U8012 ( .A(n8656), .B(n8657), .Z(n8645) );
  AND U8013 ( .A(n1325), .B(n8658), .Z(n8657) );
  XOR U8014 ( .A(p_input[1061]), .B(n8656), .Z(n8658) );
  XOR U8015 ( .A(n8659), .B(n8660), .Z(n8656) );
  AND U8016 ( .A(n1329), .B(n8661), .Z(n8660) );
  IV U8017 ( .A(n8653), .Z(n8655) );
  XOR U8018 ( .A(n8662), .B(n8663), .Z(n8653) );
  AND U8019 ( .A(n1333), .B(n8664), .Z(n8663) );
  XOR U8020 ( .A(n8665), .B(n8666), .Z(n8651) );
  AND U8021 ( .A(n1337), .B(n8664), .Z(n8666) );
  XNOR U8022 ( .A(n8665), .B(n8662), .Z(n8664) );
  XOR U8023 ( .A(n8667), .B(n8668), .Z(n8662) );
  AND U8024 ( .A(n1340), .B(n8661), .Z(n8668) );
  XNOR U8025 ( .A(n8669), .B(n8659), .Z(n8661) );
  XOR U8026 ( .A(n8670), .B(n8671), .Z(n8659) );
  AND U8027 ( .A(n1344), .B(n8672), .Z(n8671) );
  XOR U8028 ( .A(p_input[1077]), .B(n8670), .Z(n8672) );
  XOR U8029 ( .A(n8673), .B(n8674), .Z(n8670) );
  AND U8030 ( .A(n1348), .B(n8675), .Z(n8674) );
  IV U8031 ( .A(n8667), .Z(n8669) );
  XOR U8032 ( .A(n8676), .B(n8677), .Z(n8667) );
  AND U8033 ( .A(n1352), .B(n8678), .Z(n8677) );
  XOR U8034 ( .A(n8679), .B(n8680), .Z(n8665) );
  AND U8035 ( .A(n1356), .B(n8678), .Z(n8680) );
  XNOR U8036 ( .A(n8679), .B(n8676), .Z(n8678) );
  XOR U8037 ( .A(n8681), .B(n8682), .Z(n8676) );
  AND U8038 ( .A(n1359), .B(n8675), .Z(n8682) );
  XNOR U8039 ( .A(n8683), .B(n8673), .Z(n8675) );
  XOR U8040 ( .A(n8684), .B(n8685), .Z(n8673) );
  AND U8041 ( .A(n1363), .B(n8686), .Z(n8685) );
  XOR U8042 ( .A(p_input[1093]), .B(n8684), .Z(n8686) );
  XOR U8043 ( .A(n8687), .B(n8688), .Z(n8684) );
  AND U8044 ( .A(n1367), .B(n8689), .Z(n8688) );
  IV U8045 ( .A(n8681), .Z(n8683) );
  XOR U8046 ( .A(n8690), .B(n8691), .Z(n8681) );
  AND U8047 ( .A(n1371), .B(n8692), .Z(n8691) );
  XOR U8048 ( .A(n8693), .B(n8694), .Z(n8679) );
  AND U8049 ( .A(n1375), .B(n8692), .Z(n8694) );
  XNOR U8050 ( .A(n8693), .B(n8690), .Z(n8692) );
  XOR U8051 ( .A(n8695), .B(n8696), .Z(n8690) );
  AND U8052 ( .A(n1378), .B(n8689), .Z(n8696) );
  XNOR U8053 ( .A(n8697), .B(n8687), .Z(n8689) );
  XOR U8054 ( .A(n8698), .B(n8699), .Z(n8687) );
  AND U8055 ( .A(n1382), .B(n8700), .Z(n8699) );
  XOR U8056 ( .A(p_input[1109]), .B(n8698), .Z(n8700) );
  XOR U8057 ( .A(n8701), .B(n8702), .Z(n8698) );
  AND U8058 ( .A(n1386), .B(n8703), .Z(n8702) );
  IV U8059 ( .A(n8695), .Z(n8697) );
  XOR U8060 ( .A(n8704), .B(n8705), .Z(n8695) );
  AND U8061 ( .A(n1390), .B(n8706), .Z(n8705) );
  XOR U8062 ( .A(n8707), .B(n8708), .Z(n8693) );
  AND U8063 ( .A(n1394), .B(n8706), .Z(n8708) );
  XNOR U8064 ( .A(n8707), .B(n8704), .Z(n8706) );
  XOR U8065 ( .A(n8709), .B(n8710), .Z(n8704) );
  AND U8066 ( .A(n1397), .B(n8703), .Z(n8710) );
  XNOR U8067 ( .A(n8711), .B(n8701), .Z(n8703) );
  XOR U8068 ( .A(n8712), .B(n8713), .Z(n8701) );
  AND U8069 ( .A(n1401), .B(n8714), .Z(n8713) );
  XOR U8070 ( .A(p_input[1125]), .B(n8712), .Z(n8714) );
  XOR U8071 ( .A(n8715), .B(n8716), .Z(n8712) );
  AND U8072 ( .A(n1405), .B(n8717), .Z(n8716) );
  IV U8073 ( .A(n8709), .Z(n8711) );
  XOR U8074 ( .A(n8718), .B(n8719), .Z(n8709) );
  AND U8075 ( .A(n1409), .B(n8720), .Z(n8719) );
  XOR U8076 ( .A(n8721), .B(n8722), .Z(n8707) );
  AND U8077 ( .A(n1413), .B(n8720), .Z(n8722) );
  XNOR U8078 ( .A(n8721), .B(n8718), .Z(n8720) );
  XOR U8079 ( .A(n8723), .B(n8724), .Z(n8718) );
  AND U8080 ( .A(n1416), .B(n8717), .Z(n8724) );
  XNOR U8081 ( .A(n8725), .B(n8715), .Z(n8717) );
  XOR U8082 ( .A(n8726), .B(n8727), .Z(n8715) );
  AND U8083 ( .A(n1420), .B(n8728), .Z(n8727) );
  XOR U8084 ( .A(p_input[1141]), .B(n8726), .Z(n8728) );
  XOR U8085 ( .A(n8729), .B(n8730), .Z(n8726) );
  AND U8086 ( .A(n1424), .B(n8731), .Z(n8730) );
  IV U8087 ( .A(n8723), .Z(n8725) );
  XOR U8088 ( .A(n8732), .B(n8733), .Z(n8723) );
  AND U8089 ( .A(n1428), .B(n8734), .Z(n8733) );
  XOR U8090 ( .A(n8735), .B(n8736), .Z(n8721) );
  AND U8091 ( .A(n1432), .B(n8734), .Z(n8736) );
  XNOR U8092 ( .A(n8735), .B(n8732), .Z(n8734) );
  XOR U8093 ( .A(n8737), .B(n8738), .Z(n8732) );
  AND U8094 ( .A(n1435), .B(n8731), .Z(n8738) );
  XNOR U8095 ( .A(n8739), .B(n8729), .Z(n8731) );
  XOR U8096 ( .A(n8740), .B(n8741), .Z(n8729) );
  AND U8097 ( .A(n1439), .B(n8742), .Z(n8741) );
  XOR U8098 ( .A(p_input[1157]), .B(n8740), .Z(n8742) );
  XOR U8099 ( .A(n8743), .B(n8744), .Z(n8740) );
  AND U8100 ( .A(n1443), .B(n8745), .Z(n8744) );
  IV U8101 ( .A(n8737), .Z(n8739) );
  XOR U8102 ( .A(n8746), .B(n8747), .Z(n8737) );
  AND U8103 ( .A(n1447), .B(n8748), .Z(n8747) );
  XOR U8104 ( .A(n8749), .B(n8750), .Z(n8735) );
  AND U8105 ( .A(n1451), .B(n8748), .Z(n8750) );
  XNOR U8106 ( .A(n8749), .B(n8746), .Z(n8748) );
  XOR U8107 ( .A(n8751), .B(n8752), .Z(n8746) );
  AND U8108 ( .A(n1454), .B(n8745), .Z(n8752) );
  XNOR U8109 ( .A(n8753), .B(n8743), .Z(n8745) );
  XOR U8110 ( .A(n8754), .B(n8755), .Z(n8743) );
  AND U8111 ( .A(n1458), .B(n8756), .Z(n8755) );
  XOR U8112 ( .A(p_input[1173]), .B(n8754), .Z(n8756) );
  XOR U8113 ( .A(n8757), .B(n8758), .Z(n8754) );
  AND U8114 ( .A(n1462), .B(n8759), .Z(n8758) );
  IV U8115 ( .A(n8751), .Z(n8753) );
  XOR U8116 ( .A(n8760), .B(n8761), .Z(n8751) );
  AND U8117 ( .A(n1466), .B(n8762), .Z(n8761) );
  XOR U8118 ( .A(n8763), .B(n8764), .Z(n8749) );
  AND U8119 ( .A(n1470), .B(n8762), .Z(n8764) );
  XNOR U8120 ( .A(n8763), .B(n8760), .Z(n8762) );
  XOR U8121 ( .A(n8765), .B(n8766), .Z(n8760) );
  AND U8122 ( .A(n1473), .B(n8759), .Z(n8766) );
  XNOR U8123 ( .A(n8767), .B(n8757), .Z(n8759) );
  XOR U8124 ( .A(n8768), .B(n8769), .Z(n8757) );
  AND U8125 ( .A(n1477), .B(n8770), .Z(n8769) );
  XOR U8126 ( .A(p_input[1189]), .B(n8768), .Z(n8770) );
  XOR U8127 ( .A(n8771), .B(n8772), .Z(n8768) );
  AND U8128 ( .A(n1481), .B(n8773), .Z(n8772) );
  IV U8129 ( .A(n8765), .Z(n8767) );
  XOR U8130 ( .A(n8774), .B(n8775), .Z(n8765) );
  AND U8131 ( .A(n1485), .B(n8776), .Z(n8775) );
  XOR U8132 ( .A(n8777), .B(n8778), .Z(n8763) );
  AND U8133 ( .A(n1489), .B(n8776), .Z(n8778) );
  XNOR U8134 ( .A(n8777), .B(n8774), .Z(n8776) );
  XOR U8135 ( .A(n8779), .B(n8780), .Z(n8774) );
  AND U8136 ( .A(n1492), .B(n8773), .Z(n8780) );
  XNOR U8137 ( .A(n8781), .B(n8771), .Z(n8773) );
  XOR U8138 ( .A(n8782), .B(n8783), .Z(n8771) );
  AND U8139 ( .A(n1496), .B(n8784), .Z(n8783) );
  XOR U8140 ( .A(p_input[1205]), .B(n8782), .Z(n8784) );
  XOR U8141 ( .A(n8785), .B(n8786), .Z(n8782) );
  AND U8142 ( .A(n1500), .B(n8787), .Z(n8786) );
  IV U8143 ( .A(n8779), .Z(n8781) );
  XOR U8144 ( .A(n8788), .B(n8789), .Z(n8779) );
  AND U8145 ( .A(n1504), .B(n8790), .Z(n8789) );
  XOR U8146 ( .A(n8791), .B(n8792), .Z(n8777) );
  AND U8147 ( .A(n1508), .B(n8790), .Z(n8792) );
  XNOR U8148 ( .A(n8791), .B(n8788), .Z(n8790) );
  XOR U8149 ( .A(n8793), .B(n8794), .Z(n8788) );
  AND U8150 ( .A(n1511), .B(n8787), .Z(n8794) );
  XNOR U8151 ( .A(n8795), .B(n8785), .Z(n8787) );
  XOR U8152 ( .A(n8796), .B(n8797), .Z(n8785) );
  AND U8153 ( .A(n1515), .B(n8798), .Z(n8797) );
  XOR U8154 ( .A(p_input[1221]), .B(n8796), .Z(n8798) );
  XOR U8155 ( .A(n8799), .B(n8800), .Z(n8796) );
  AND U8156 ( .A(n1519), .B(n8801), .Z(n8800) );
  IV U8157 ( .A(n8793), .Z(n8795) );
  XOR U8158 ( .A(n8802), .B(n8803), .Z(n8793) );
  AND U8159 ( .A(n1523), .B(n8804), .Z(n8803) );
  XOR U8160 ( .A(n8805), .B(n8806), .Z(n8791) );
  AND U8161 ( .A(n1527), .B(n8804), .Z(n8806) );
  XNOR U8162 ( .A(n8805), .B(n8802), .Z(n8804) );
  XOR U8163 ( .A(n8807), .B(n8808), .Z(n8802) );
  AND U8164 ( .A(n1530), .B(n8801), .Z(n8808) );
  XNOR U8165 ( .A(n8809), .B(n8799), .Z(n8801) );
  XOR U8166 ( .A(n8810), .B(n8811), .Z(n8799) );
  AND U8167 ( .A(n1534), .B(n8812), .Z(n8811) );
  XOR U8168 ( .A(p_input[1237]), .B(n8810), .Z(n8812) );
  XOR U8169 ( .A(n8813), .B(n8814), .Z(n8810) );
  AND U8170 ( .A(n1538), .B(n8815), .Z(n8814) );
  IV U8171 ( .A(n8807), .Z(n8809) );
  XOR U8172 ( .A(n8816), .B(n8817), .Z(n8807) );
  AND U8173 ( .A(n1542), .B(n8818), .Z(n8817) );
  XOR U8174 ( .A(n8819), .B(n8820), .Z(n8805) );
  AND U8175 ( .A(n1546), .B(n8818), .Z(n8820) );
  XNOR U8176 ( .A(n8819), .B(n8816), .Z(n8818) );
  XOR U8177 ( .A(n8821), .B(n8822), .Z(n8816) );
  AND U8178 ( .A(n1549), .B(n8815), .Z(n8822) );
  XNOR U8179 ( .A(n8823), .B(n8813), .Z(n8815) );
  XOR U8180 ( .A(n8824), .B(n8825), .Z(n8813) );
  AND U8181 ( .A(n1553), .B(n8826), .Z(n8825) );
  XOR U8182 ( .A(p_input[1253]), .B(n8824), .Z(n8826) );
  XOR U8183 ( .A(n8827), .B(n8828), .Z(n8824) );
  AND U8184 ( .A(n1557), .B(n8829), .Z(n8828) );
  IV U8185 ( .A(n8821), .Z(n8823) );
  XOR U8186 ( .A(n8830), .B(n8831), .Z(n8821) );
  AND U8187 ( .A(n1561), .B(n8832), .Z(n8831) );
  XOR U8188 ( .A(n8833), .B(n8834), .Z(n8819) );
  AND U8189 ( .A(n1565), .B(n8832), .Z(n8834) );
  XNOR U8190 ( .A(n8833), .B(n8830), .Z(n8832) );
  XOR U8191 ( .A(n8835), .B(n8836), .Z(n8830) );
  AND U8192 ( .A(n1568), .B(n8829), .Z(n8836) );
  XNOR U8193 ( .A(n8837), .B(n8827), .Z(n8829) );
  XOR U8194 ( .A(n8838), .B(n8839), .Z(n8827) );
  AND U8195 ( .A(n1572), .B(n8840), .Z(n8839) );
  XOR U8196 ( .A(p_input[1269]), .B(n8838), .Z(n8840) );
  XOR U8197 ( .A(n8841), .B(n8842), .Z(n8838) );
  AND U8198 ( .A(n1576), .B(n8843), .Z(n8842) );
  IV U8199 ( .A(n8835), .Z(n8837) );
  XOR U8200 ( .A(n8844), .B(n8845), .Z(n8835) );
  AND U8201 ( .A(n1580), .B(n8846), .Z(n8845) );
  XOR U8202 ( .A(n8847), .B(n8848), .Z(n8833) );
  AND U8203 ( .A(n1584), .B(n8846), .Z(n8848) );
  XNOR U8204 ( .A(n8847), .B(n8844), .Z(n8846) );
  XOR U8205 ( .A(n8849), .B(n8850), .Z(n8844) );
  AND U8206 ( .A(n1587), .B(n8843), .Z(n8850) );
  XNOR U8207 ( .A(n8851), .B(n8841), .Z(n8843) );
  XOR U8208 ( .A(n8852), .B(n8853), .Z(n8841) );
  AND U8209 ( .A(n1591), .B(n8854), .Z(n8853) );
  XOR U8210 ( .A(p_input[1285]), .B(n8852), .Z(n8854) );
  XOR U8211 ( .A(n8855), .B(n8856), .Z(n8852) );
  AND U8212 ( .A(n1595), .B(n8857), .Z(n8856) );
  IV U8213 ( .A(n8849), .Z(n8851) );
  XOR U8214 ( .A(n8858), .B(n8859), .Z(n8849) );
  AND U8215 ( .A(n1599), .B(n8860), .Z(n8859) );
  XOR U8216 ( .A(n8861), .B(n8862), .Z(n8847) );
  AND U8217 ( .A(n1603), .B(n8860), .Z(n8862) );
  XNOR U8218 ( .A(n8861), .B(n8858), .Z(n8860) );
  XOR U8219 ( .A(n8863), .B(n8864), .Z(n8858) );
  AND U8220 ( .A(n1606), .B(n8857), .Z(n8864) );
  XNOR U8221 ( .A(n8865), .B(n8855), .Z(n8857) );
  XOR U8222 ( .A(n8866), .B(n8867), .Z(n8855) );
  AND U8223 ( .A(n1610), .B(n8868), .Z(n8867) );
  XOR U8224 ( .A(p_input[1301]), .B(n8866), .Z(n8868) );
  XOR U8225 ( .A(n8869), .B(n8870), .Z(n8866) );
  AND U8226 ( .A(n1614), .B(n8871), .Z(n8870) );
  IV U8227 ( .A(n8863), .Z(n8865) );
  XOR U8228 ( .A(n8872), .B(n8873), .Z(n8863) );
  AND U8229 ( .A(n1618), .B(n8874), .Z(n8873) );
  XOR U8230 ( .A(n8875), .B(n8876), .Z(n8861) );
  AND U8231 ( .A(n1622), .B(n8874), .Z(n8876) );
  XNOR U8232 ( .A(n8875), .B(n8872), .Z(n8874) );
  XOR U8233 ( .A(n8877), .B(n8878), .Z(n8872) );
  AND U8234 ( .A(n1625), .B(n8871), .Z(n8878) );
  XNOR U8235 ( .A(n8879), .B(n8869), .Z(n8871) );
  XOR U8236 ( .A(n8880), .B(n8881), .Z(n8869) );
  AND U8237 ( .A(n1629), .B(n8882), .Z(n8881) );
  XOR U8238 ( .A(p_input[1317]), .B(n8880), .Z(n8882) );
  XOR U8239 ( .A(n8883), .B(n8884), .Z(n8880) );
  AND U8240 ( .A(n1633), .B(n8885), .Z(n8884) );
  IV U8241 ( .A(n8877), .Z(n8879) );
  XOR U8242 ( .A(n8886), .B(n8887), .Z(n8877) );
  AND U8243 ( .A(n1637), .B(n8888), .Z(n8887) );
  XOR U8244 ( .A(n8889), .B(n8890), .Z(n8875) );
  AND U8245 ( .A(n1641), .B(n8888), .Z(n8890) );
  XNOR U8246 ( .A(n8889), .B(n8886), .Z(n8888) );
  XOR U8247 ( .A(n8891), .B(n8892), .Z(n8886) );
  AND U8248 ( .A(n1644), .B(n8885), .Z(n8892) );
  XNOR U8249 ( .A(n8893), .B(n8883), .Z(n8885) );
  XOR U8250 ( .A(n8894), .B(n8895), .Z(n8883) );
  AND U8251 ( .A(n1648), .B(n8896), .Z(n8895) );
  XOR U8252 ( .A(p_input[1333]), .B(n8894), .Z(n8896) );
  XOR U8253 ( .A(n8897), .B(n8898), .Z(n8894) );
  AND U8254 ( .A(n1652), .B(n8899), .Z(n8898) );
  IV U8255 ( .A(n8891), .Z(n8893) );
  XOR U8256 ( .A(n8900), .B(n8901), .Z(n8891) );
  AND U8257 ( .A(n1656), .B(n8902), .Z(n8901) );
  XOR U8258 ( .A(n8903), .B(n8904), .Z(n8889) );
  AND U8259 ( .A(n1660), .B(n8902), .Z(n8904) );
  XNOR U8260 ( .A(n8903), .B(n8900), .Z(n8902) );
  XOR U8261 ( .A(n8905), .B(n8906), .Z(n8900) );
  AND U8262 ( .A(n1663), .B(n8899), .Z(n8906) );
  XNOR U8263 ( .A(n8907), .B(n8897), .Z(n8899) );
  XOR U8264 ( .A(n8908), .B(n8909), .Z(n8897) );
  AND U8265 ( .A(n1667), .B(n8910), .Z(n8909) );
  XOR U8266 ( .A(p_input[1349]), .B(n8908), .Z(n8910) );
  XOR U8267 ( .A(n8911), .B(n8912), .Z(n8908) );
  AND U8268 ( .A(n1671), .B(n8913), .Z(n8912) );
  IV U8269 ( .A(n8905), .Z(n8907) );
  XOR U8270 ( .A(n8914), .B(n8915), .Z(n8905) );
  AND U8271 ( .A(n1675), .B(n8916), .Z(n8915) );
  XOR U8272 ( .A(n8917), .B(n8918), .Z(n8903) );
  AND U8273 ( .A(n1679), .B(n8916), .Z(n8918) );
  XNOR U8274 ( .A(n8917), .B(n8914), .Z(n8916) );
  XOR U8275 ( .A(n8919), .B(n8920), .Z(n8914) );
  AND U8276 ( .A(n1682), .B(n8913), .Z(n8920) );
  XNOR U8277 ( .A(n8921), .B(n8911), .Z(n8913) );
  XOR U8278 ( .A(n8922), .B(n8923), .Z(n8911) );
  AND U8279 ( .A(n1686), .B(n8924), .Z(n8923) );
  XOR U8280 ( .A(p_input[1365]), .B(n8922), .Z(n8924) );
  XOR U8281 ( .A(n8925), .B(n8926), .Z(n8922) );
  AND U8282 ( .A(n1690), .B(n8927), .Z(n8926) );
  IV U8283 ( .A(n8919), .Z(n8921) );
  XOR U8284 ( .A(n8928), .B(n8929), .Z(n8919) );
  AND U8285 ( .A(n1694), .B(n8930), .Z(n8929) );
  XOR U8286 ( .A(n8931), .B(n8932), .Z(n8917) );
  AND U8287 ( .A(n1698), .B(n8930), .Z(n8932) );
  XNOR U8288 ( .A(n8931), .B(n8928), .Z(n8930) );
  XOR U8289 ( .A(n8933), .B(n8934), .Z(n8928) );
  AND U8290 ( .A(n1701), .B(n8927), .Z(n8934) );
  XNOR U8291 ( .A(n8935), .B(n8925), .Z(n8927) );
  XOR U8292 ( .A(n8936), .B(n8937), .Z(n8925) );
  AND U8293 ( .A(n1705), .B(n8938), .Z(n8937) );
  XOR U8294 ( .A(p_input[1381]), .B(n8936), .Z(n8938) );
  XOR U8295 ( .A(n8939), .B(n8940), .Z(n8936) );
  AND U8296 ( .A(n1709), .B(n8941), .Z(n8940) );
  IV U8297 ( .A(n8933), .Z(n8935) );
  XOR U8298 ( .A(n8942), .B(n8943), .Z(n8933) );
  AND U8299 ( .A(n1713), .B(n8944), .Z(n8943) );
  XOR U8300 ( .A(n8945), .B(n8946), .Z(n8931) );
  AND U8301 ( .A(n1717), .B(n8944), .Z(n8946) );
  XNOR U8302 ( .A(n8945), .B(n8942), .Z(n8944) );
  XOR U8303 ( .A(n8947), .B(n8948), .Z(n8942) );
  AND U8304 ( .A(n1720), .B(n8941), .Z(n8948) );
  XNOR U8305 ( .A(n8949), .B(n8939), .Z(n8941) );
  XOR U8306 ( .A(n8950), .B(n8951), .Z(n8939) );
  AND U8307 ( .A(n1724), .B(n8952), .Z(n8951) );
  XOR U8308 ( .A(p_input[1397]), .B(n8950), .Z(n8952) );
  XOR U8309 ( .A(n8953), .B(n8954), .Z(n8950) );
  AND U8310 ( .A(n1728), .B(n8955), .Z(n8954) );
  IV U8311 ( .A(n8947), .Z(n8949) );
  XOR U8312 ( .A(n8956), .B(n8957), .Z(n8947) );
  AND U8313 ( .A(n1732), .B(n8958), .Z(n8957) );
  XOR U8314 ( .A(n8959), .B(n8960), .Z(n8945) );
  AND U8315 ( .A(n1736), .B(n8958), .Z(n8960) );
  XNOR U8316 ( .A(n8959), .B(n8956), .Z(n8958) );
  XOR U8317 ( .A(n8961), .B(n8962), .Z(n8956) );
  AND U8318 ( .A(n1739), .B(n8955), .Z(n8962) );
  XNOR U8319 ( .A(n8963), .B(n8953), .Z(n8955) );
  XOR U8320 ( .A(n8964), .B(n8965), .Z(n8953) );
  AND U8321 ( .A(n1743), .B(n8966), .Z(n8965) );
  XOR U8322 ( .A(p_input[1413]), .B(n8964), .Z(n8966) );
  XOR U8323 ( .A(n8967), .B(n8968), .Z(n8964) );
  AND U8324 ( .A(n1747), .B(n8969), .Z(n8968) );
  IV U8325 ( .A(n8961), .Z(n8963) );
  XOR U8326 ( .A(n8970), .B(n8971), .Z(n8961) );
  AND U8327 ( .A(n1751), .B(n8972), .Z(n8971) );
  XOR U8328 ( .A(n8973), .B(n8974), .Z(n8959) );
  AND U8329 ( .A(n1755), .B(n8972), .Z(n8974) );
  XNOR U8330 ( .A(n8973), .B(n8970), .Z(n8972) );
  XOR U8331 ( .A(n8975), .B(n8976), .Z(n8970) );
  AND U8332 ( .A(n1758), .B(n8969), .Z(n8976) );
  XNOR U8333 ( .A(n8977), .B(n8967), .Z(n8969) );
  XOR U8334 ( .A(n8978), .B(n8979), .Z(n8967) );
  AND U8335 ( .A(n1762), .B(n8980), .Z(n8979) );
  XOR U8336 ( .A(p_input[1429]), .B(n8978), .Z(n8980) );
  XOR U8337 ( .A(n8981), .B(n8982), .Z(n8978) );
  AND U8338 ( .A(n1766), .B(n8983), .Z(n8982) );
  IV U8339 ( .A(n8975), .Z(n8977) );
  XOR U8340 ( .A(n8984), .B(n8985), .Z(n8975) );
  AND U8341 ( .A(n1770), .B(n8986), .Z(n8985) );
  XOR U8342 ( .A(n8987), .B(n8988), .Z(n8973) );
  AND U8343 ( .A(n1774), .B(n8986), .Z(n8988) );
  XNOR U8344 ( .A(n8987), .B(n8984), .Z(n8986) );
  XOR U8345 ( .A(n8989), .B(n8990), .Z(n8984) );
  AND U8346 ( .A(n1777), .B(n8983), .Z(n8990) );
  XNOR U8347 ( .A(n8991), .B(n8981), .Z(n8983) );
  XOR U8348 ( .A(n8992), .B(n8993), .Z(n8981) );
  AND U8349 ( .A(n1781), .B(n8994), .Z(n8993) );
  XOR U8350 ( .A(p_input[1445]), .B(n8992), .Z(n8994) );
  XOR U8351 ( .A(n8995), .B(n8996), .Z(n8992) );
  AND U8352 ( .A(n1785), .B(n8997), .Z(n8996) );
  IV U8353 ( .A(n8989), .Z(n8991) );
  XOR U8354 ( .A(n8998), .B(n8999), .Z(n8989) );
  AND U8355 ( .A(n1789), .B(n9000), .Z(n8999) );
  XOR U8356 ( .A(n9001), .B(n9002), .Z(n8987) );
  AND U8357 ( .A(n1793), .B(n9000), .Z(n9002) );
  XNOR U8358 ( .A(n9001), .B(n8998), .Z(n9000) );
  XOR U8359 ( .A(n9003), .B(n9004), .Z(n8998) );
  AND U8360 ( .A(n1796), .B(n8997), .Z(n9004) );
  XNOR U8361 ( .A(n9005), .B(n8995), .Z(n8997) );
  XOR U8362 ( .A(n9006), .B(n9007), .Z(n8995) );
  AND U8363 ( .A(n1800), .B(n9008), .Z(n9007) );
  XOR U8364 ( .A(p_input[1461]), .B(n9006), .Z(n9008) );
  XOR U8365 ( .A(n9009), .B(n9010), .Z(n9006) );
  AND U8366 ( .A(n1804), .B(n9011), .Z(n9010) );
  IV U8367 ( .A(n9003), .Z(n9005) );
  XOR U8368 ( .A(n9012), .B(n9013), .Z(n9003) );
  AND U8369 ( .A(n1808), .B(n9014), .Z(n9013) );
  XOR U8370 ( .A(n9015), .B(n9016), .Z(n9001) );
  AND U8371 ( .A(n1812), .B(n9014), .Z(n9016) );
  XNOR U8372 ( .A(n9015), .B(n9012), .Z(n9014) );
  XOR U8373 ( .A(n9017), .B(n9018), .Z(n9012) );
  AND U8374 ( .A(n1815), .B(n9011), .Z(n9018) );
  XNOR U8375 ( .A(n9019), .B(n9009), .Z(n9011) );
  XOR U8376 ( .A(n9020), .B(n9021), .Z(n9009) );
  AND U8377 ( .A(n1819), .B(n9022), .Z(n9021) );
  XOR U8378 ( .A(p_input[1477]), .B(n9020), .Z(n9022) );
  XOR U8379 ( .A(n9023), .B(n9024), .Z(n9020) );
  AND U8380 ( .A(n1823), .B(n9025), .Z(n9024) );
  IV U8381 ( .A(n9017), .Z(n9019) );
  XOR U8382 ( .A(n9026), .B(n9027), .Z(n9017) );
  AND U8383 ( .A(n1827), .B(n9028), .Z(n9027) );
  XOR U8384 ( .A(n9029), .B(n9030), .Z(n9015) );
  AND U8385 ( .A(n1831), .B(n9028), .Z(n9030) );
  XNOR U8386 ( .A(n9029), .B(n9026), .Z(n9028) );
  XOR U8387 ( .A(n9031), .B(n9032), .Z(n9026) );
  AND U8388 ( .A(n1834), .B(n9025), .Z(n9032) );
  XNOR U8389 ( .A(n9033), .B(n9023), .Z(n9025) );
  XOR U8390 ( .A(n9034), .B(n9035), .Z(n9023) );
  AND U8391 ( .A(n1838), .B(n9036), .Z(n9035) );
  XOR U8392 ( .A(p_input[1493]), .B(n9034), .Z(n9036) );
  XOR U8393 ( .A(n9037), .B(n9038), .Z(n9034) );
  AND U8394 ( .A(n1842), .B(n9039), .Z(n9038) );
  IV U8395 ( .A(n9031), .Z(n9033) );
  XOR U8396 ( .A(n9040), .B(n9041), .Z(n9031) );
  AND U8397 ( .A(n1846), .B(n9042), .Z(n9041) );
  XOR U8398 ( .A(n9043), .B(n9044), .Z(n9029) );
  AND U8399 ( .A(n1850), .B(n9042), .Z(n9044) );
  XNOR U8400 ( .A(n9043), .B(n9040), .Z(n9042) );
  XOR U8401 ( .A(n9045), .B(n9046), .Z(n9040) );
  AND U8402 ( .A(n1853), .B(n9039), .Z(n9046) );
  XNOR U8403 ( .A(n9047), .B(n9037), .Z(n9039) );
  XOR U8404 ( .A(n9048), .B(n9049), .Z(n9037) );
  AND U8405 ( .A(n1857), .B(n9050), .Z(n9049) );
  XOR U8406 ( .A(p_input[1509]), .B(n9048), .Z(n9050) );
  XOR U8407 ( .A(n9051), .B(n9052), .Z(n9048) );
  AND U8408 ( .A(n1861), .B(n9053), .Z(n9052) );
  IV U8409 ( .A(n9045), .Z(n9047) );
  XOR U8410 ( .A(n9054), .B(n9055), .Z(n9045) );
  AND U8411 ( .A(n1865), .B(n9056), .Z(n9055) );
  XOR U8412 ( .A(n9057), .B(n9058), .Z(n9043) );
  AND U8413 ( .A(n1869), .B(n9056), .Z(n9058) );
  XNOR U8414 ( .A(n9057), .B(n9054), .Z(n9056) );
  XOR U8415 ( .A(n9059), .B(n9060), .Z(n9054) );
  AND U8416 ( .A(n1872), .B(n9053), .Z(n9060) );
  XNOR U8417 ( .A(n9061), .B(n9051), .Z(n9053) );
  XOR U8418 ( .A(n9062), .B(n9063), .Z(n9051) );
  AND U8419 ( .A(n1876), .B(n9064), .Z(n9063) );
  XOR U8420 ( .A(p_input[1525]), .B(n9062), .Z(n9064) );
  XOR U8421 ( .A(n9065), .B(n9066), .Z(n9062) );
  AND U8422 ( .A(n1880), .B(n9067), .Z(n9066) );
  IV U8423 ( .A(n9059), .Z(n9061) );
  XOR U8424 ( .A(n9068), .B(n9069), .Z(n9059) );
  AND U8425 ( .A(n1884), .B(n9070), .Z(n9069) );
  XOR U8426 ( .A(n9071), .B(n9072), .Z(n9057) );
  AND U8427 ( .A(n1888), .B(n9070), .Z(n9072) );
  XNOR U8428 ( .A(n9071), .B(n9068), .Z(n9070) );
  XOR U8429 ( .A(n9073), .B(n9074), .Z(n9068) );
  AND U8430 ( .A(n1891), .B(n9067), .Z(n9074) );
  XNOR U8431 ( .A(n9075), .B(n9065), .Z(n9067) );
  XOR U8432 ( .A(n9076), .B(n9077), .Z(n9065) );
  AND U8433 ( .A(n1895), .B(n9078), .Z(n9077) );
  XOR U8434 ( .A(p_input[1541]), .B(n9076), .Z(n9078) );
  XOR U8435 ( .A(n9079), .B(n9080), .Z(n9076) );
  AND U8436 ( .A(n1899), .B(n9081), .Z(n9080) );
  IV U8437 ( .A(n9073), .Z(n9075) );
  XOR U8438 ( .A(n9082), .B(n9083), .Z(n9073) );
  AND U8439 ( .A(n1903), .B(n9084), .Z(n9083) );
  XOR U8440 ( .A(n9085), .B(n9086), .Z(n9071) );
  AND U8441 ( .A(n1907), .B(n9084), .Z(n9086) );
  XNOR U8442 ( .A(n9085), .B(n9082), .Z(n9084) );
  XOR U8443 ( .A(n9087), .B(n9088), .Z(n9082) );
  AND U8444 ( .A(n1910), .B(n9081), .Z(n9088) );
  XNOR U8445 ( .A(n9089), .B(n9079), .Z(n9081) );
  XOR U8446 ( .A(n9090), .B(n9091), .Z(n9079) );
  AND U8447 ( .A(n1914), .B(n9092), .Z(n9091) );
  XOR U8448 ( .A(p_input[1557]), .B(n9090), .Z(n9092) );
  XOR U8449 ( .A(n9093), .B(n9094), .Z(n9090) );
  AND U8450 ( .A(n1918), .B(n9095), .Z(n9094) );
  IV U8451 ( .A(n9087), .Z(n9089) );
  XOR U8452 ( .A(n9096), .B(n9097), .Z(n9087) );
  AND U8453 ( .A(n1922), .B(n9098), .Z(n9097) );
  XOR U8454 ( .A(n9099), .B(n9100), .Z(n9085) );
  AND U8455 ( .A(n1926), .B(n9098), .Z(n9100) );
  XNOR U8456 ( .A(n9099), .B(n9096), .Z(n9098) );
  XOR U8457 ( .A(n9101), .B(n9102), .Z(n9096) );
  AND U8458 ( .A(n1929), .B(n9095), .Z(n9102) );
  XNOR U8459 ( .A(n9103), .B(n9093), .Z(n9095) );
  XOR U8460 ( .A(n9104), .B(n9105), .Z(n9093) );
  AND U8461 ( .A(n1933), .B(n9106), .Z(n9105) );
  XOR U8462 ( .A(p_input[1573]), .B(n9104), .Z(n9106) );
  XOR U8463 ( .A(n9107), .B(n9108), .Z(n9104) );
  AND U8464 ( .A(n1937), .B(n9109), .Z(n9108) );
  IV U8465 ( .A(n9101), .Z(n9103) );
  XOR U8466 ( .A(n9110), .B(n9111), .Z(n9101) );
  AND U8467 ( .A(n1941), .B(n9112), .Z(n9111) );
  XOR U8468 ( .A(n9113), .B(n9114), .Z(n9099) );
  AND U8469 ( .A(n1945), .B(n9112), .Z(n9114) );
  XNOR U8470 ( .A(n9113), .B(n9110), .Z(n9112) );
  XOR U8471 ( .A(n9115), .B(n9116), .Z(n9110) );
  AND U8472 ( .A(n1948), .B(n9109), .Z(n9116) );
  XNOR U8473 ( .A(n9117), .B(n9107), .Z(n9109) );
  XOR U8474 ( .A(n9118), .B(n9119), .Z(n9107) );
  AND U8475 ( .A(n1952), .B(n9120), .Z(n9119) );
  XOR U8476 ( .A(p_input[1589]), .B(n9118), .Z(n9120) );
  XOR U8477 ( .A(n9121), .B(n9122), .Z(n9118) );
  AND U8478 ( .A(n1956), .B(n9123), .Z(n9122) );
  IV U8479 ( .A(n9115), .Z(n9117) );
  XOR U8480 ( .A(n9124), .B(n9125), .Z(n9115) );
  AND U8481 ( .A(n1960), .B(n9126), .Z(n9125) );
  XOR U8482 ( .A(n9127), .B(n9128), .Z(n9113) );
  AND U8483 ( .A(n1964), .B(n9126), .Z(n9128) );
  XNOR U8484 ( .A(n9127), .B(n9124), .Z(n9126) );
  XOR U8485 ( .A(n9129), .B(n9130), .Z(n9124) );
  AND U8486 ( .A(n1967), .B(n9123), .Z(n9130) );
  XNOR U8487 ( .A(n9131), .B(n9121), .Z(n9123) );
  XOR U8488 ( .A(n9132), .B(n9133), .Z(n9121) );
  AND U8489 ( .A(n1971), .B(n9134), .Z(n9133) );
  XOR U8490 ( .A(p_input[1605]), .B(n9132), .Z(n9134) );
  XOR U8491 ( .A(n9135), .B(n9136), .Z(n9132) );
  AND U8492 ( .A(n1975), .B(n9137), .Z(n9136) );
  IV U8493 ( .A(n9129), .Z(n9131) );
  XOR U8494 ( .A(n9138), .B(n9139), .Z(n9129) );
  AND U8495 ( .A(n1979), .B(n9140), .Z(n9139) );
  XOR U8496 ( .A(n9141), .B(n9142), .Z(n9127) );
  AND U8497 ( .A(n1983), .B(n9140), .Z(n9142) );
  XNOR U8498 ( .A(n9141), .B(n9138), .Z(n9140) );
  XOR U8499 ( .A(n9143), .B(n9144), .Z(n9138) );
  AND U8500 ( .A(n1986), .B(n9137), .Z(n9144) );
  XNOR U8501 ( .A(n9145), .B(n9135), .Z(n9137) );
  XOR U8502 ( .A(n9146), .B(n9147), .Z(n9135) );
  AND U8503 ( .A(n1990), .B(n9148), .Z(n9147) );
  XOR U8504 ( .A(p_input[1621]), .B(n9146), .Z(n9148) );
  XOR U8505 ( .A(n9149), .B(n9150), .Z(n9146) );
  AND U8506 ( .A(n1994), .B(n9151), .Z(n9150) );
  IV U8507 ( .A(n9143), .Z(n9145) );
  XOR U8508 ( .A(n9152), .B(n9153), .Z(n9143) );
  AND U8509 ( .A(n1998), .B(n9154), .Z(n9153) );
  XOR U8510 ( .A(n9155), .B(n9156), .Z(n9141) );
  AND U8511 ( .A(n2002), .B(n9154), .Z(n9156) );
  XNOR U8512 ( .A(n9155), .B(n9152), .Z(n9154) );
  XOR U8513 ( .A(n9157), .B(n9158), .Z(n9152) );
  AND U8514 ( .A(n2005), .B(n9151), .Z(n9158) );
  XNOR U8515 ( .A(n9159), .B(n9149), .Z(n9151) );
  XOR U8516 ( .A(n9160), .B(n9161), .Z(n9149) );
  AND U8517 ( .A(n2009), .B(n9162), .Z(n9161) );
  XOR U8518 ( .A(p_input[1637]), .B(n9160), .Z(n9162) );
  XOR U8519 ( .A(n9163), .B(n9164), .Z(n9160) );
  AND U8520 ( .A(n2013), .B(n9165), .Z(n9164) );
  IV U8521 ( .A(n9157), .Z(n9159) );
  XOR U8522 ( .A(n9166), .B(n9167), .Z(n9157) );
  AND U8523 ( .A(n2017), .B(n9168), .Z(n9167) );
  XOR U8524 ( .A(n9169), .B(n9170), .Z(n9155) );
  AND U8525 ( .A(n2021), .B(n9168), .Z(n9170) );
  XNOR U8526 ( .A(n9169), .B(n9166), .Z(n9168) );
  XOR U8527 ( .A(n9171), .B(n9172), .Z(n9166) );
  AND U8528 ( .A(n2024), .B(n9165), .Z(n9172) );
  XNOR U8529 ( .A(n9173), .B(n9163), .Z(n9165) );
  XOR U8530 ( .A(n9174), .B(n9175), .Z(n9163) );
  AND U8531 ( .A(n2028), .B(n9176), .Z(n9175) );
  XOR U8532 ( .A(p_input[1653]), .B(n9174), .Z(n9176) );
  XOR U8533 ( .A(n9177), .B(n9178), .Z(n9174) );
  AND U8534 ( .A(n2032), .B(n9179), .Z(n9178) );
  IV U8535 ( .A(n9171), .Z(n9173) );
  XOR U8536 ( .A(n9180), .B(n9181), .Z(n9171) );
  AND U8537 ( .A(n2036), .B(n9182), .Z(n9181) );
  XOR U8538 ( .A(n9183), .B(n9184), .Z(n9169) );
  AND U8539 ( .A(n2040), .B(n9182), .Z(n9184) );
  XNOR U8540 ( .A(n9183), .B(n9180), .Z(n9182) );
  XOR U8541 ( .A(n9185), .B(n9186), .Z(n9180) );
  AND U8542 ( .A(n2043), .B(n9179), .Z(n9186) );
  XNOR U8543 ( .A(n9187), .B(n9177), .Z(n9179) );
  XOR U8544 ( .A(n9188), .B(n9189), .Z(n9177) );
  AND U8545 ( .A(n2047), .B(n9190), .Z(n9189) );
  XOR U8546 ( .A(p_input[1669]), .B(n9188), .Z(n9190) );
  XOR U8547 ( .A(n9191), .B(n9192), .Z(n9188) );
  AND U8548 ( .A(n2051), .B(n9193), .Z(n9192) );
  IV U8549 ( .A(n9185), .Z(n9187) );
  XOR U8550 ( .A(n9194), .B(n9195), .Z(n9185) );
  AND U8551 ( .A(n2055), .B(n9196), .Z(n9195) );
  XOR U8552 ( .A(n9197), .B(n9198), .Z(n9183) );
  AND U8553 ( .A(n2059), .B(n9196), .Z(n9198) );
  XNOR U8554 ( .A(n9197), .B(n9194), .Z(n9196) );
  XOR U8555 ( .A(n9199), .B(n9200), .Z(n9194) );
  AND U8556 ( .A(n2062), .B(n9193), .Z(n9200) );
  XNOR U8557 ( .A(n9201), .B(n9191), .Z(n9193) );
  XOR U8558 ( .A(n9202), .B(n9203), .Z(n9191) );
  AND U8559 ( .A(n2066), .B(n9204), .Z(n9203) );
  XOR U8560 ( .A(p_input[1685]), .B(n9202), .Z(n9204) );
  XOR U8561 ( .A(n9205), .B(n9206), .Z(n9202) );
  AND U8562 ( .A(n2070), .B(n9207), .Z(n9206) );
  IV U8563 ( .A(n9199), .Z(n9201) );
  XOR U8564 ( .A(n9208), .B(n9209), .Z(n9199) );
  AND U8565 ( .A(n2074), .B(n9210), .Z(n9209) );
  XOR U8566 ( .A(n9211), .B(n9212), .Z(n9197) );
  AND U8567 ( .A(n2078), .B(n9210), .Z(n9212) );
  XNOR U8568 ( .A(n9211), .B(n9208), .Z(n9210) );
  XOR U8569 ( .A(n9213), .B(n9214), .Z(n9208) );
  AND U8570 ( .A(n2081), .B(n9207), .Z(n9214) );
  XNOR U8571 ( .A(n9215), .B(n9205), .Z(n9207) );
  XOR U8572 ( .A(n9216), .B(n9217), .Z(n9205) );
  AND U8573 ( .A(n2085), .B(n9218), .Z(n9217) );
  XOR U8574 ( .A(p_input[1701]), .B(n9216), .Z(n9218) );
  XOR U8575 ( .A(n9219), .B(n9220), .Z(n9216) );
  AND U8576 ( .A(n2089), .B(n9221), .Z(n9220) );
  IV U8577 ( .A(n9213), .Z(n9215) );
  XOR U8578 ( .A(n9222), .B(n9223), .Z(n9213) );
  AND U8579 ( .A(n2093), .B(n9224), .Z(n9223) );
  XOR U8580 ( .A(n9225), .B(n9226), .Z(n9211) );
  AND U8581 ( .A(n2097), .B(n9224), .Z(n9226) );
  XNOR U8582 ( .A(n9225), .B(n9222), .Z(n9224) );
  XOR U8583 ( .A(n9227), .B(n9228), .Z(n9222) );
  AND U8584 ( .A(n2100), .B(n9221), .Z(n9228) );
  XNOR U8585 ( .A(n9229), .B(n9219), .Z(n9221) );
  XOR U8586 ( .A(n9230), .B(n9231), .Z(n9219) );
  AND U8587 ( .A(n2104), .B(n9232), .Z(n9231) );
  XOR U8588 ( .A(p_input[1717]), .B(n9230), .Z(n9232) );
  XOR U8589 ( .A(n9233), .B(n9234), .Z(n9230) );
  AND U8590 ( .A(n2108), .B(n9235), .Z(n9234) );
  IV U8591 ( .A(n9227), .Z(n9229) );
  XOR U8592 ( .A(n9236), .B(n9237), .Z(n9227) );
  AND U8593 ( .A(n2112), .B(n9238), .Z(n9237) );
  XOR U8594 ( .A(n9239), .B(n9240), .Z(n9225) );
  AND U8595 ( .A(n2116), .B(n9238), .Z(n9240) );
  XNOR U8596 ( .A(n9239), .B(n9236), .Z(n9238) );
  XOR U8597 ( .A(n9241), .B(n9242), .Z(n9236) );
  AND U8598 ( .A(n2119), .B(n9235), .Z(n9242) );
  XNOR U8599 ( .A(n9243), .B(n9233), .Z(n9235) );
  XOR U8600 ( .A(n9244), .B(n9245), .Z(n9233) );
  AND U8601 ( .A(n2123), .B(n9246), .Z(n9245) );
  XOR U8602 ( .A(p_input[1733]), .B(n9244), .Z(n9246) );
  XOR U8603 ( .A(n9247), .B(n9248), .Z(n9244) );
  AND U8604 ( .A(n2127), .B(n9249), .Z(n9248) );
  IV U8605 ( .A(n9241), .Z(n9243) );
  XOR U8606 ( .A(n9250), .B(n9251), .Z(n9241) );
  AND U8607 ( .A(n2131), .B(n9252), .Z(n9251) );
  XOR U8608 ( .A(n9253), .B(n9254), .Z(n9239) );
  AND U8609 ( .A(n2135), .B(n9252), .Z(n9254) );
  XNOR U8610 ( .A(n9253), .B(n9250), .Z(n9252) );
  XOR U8611 ( .A(n9255), .B(n9256), .Z(n9250) );
  AND U8612 ( .A(n2138), .B(n9249), .Z(n9256) );
  XNOR U8613 ( .A(n9257), .B(n9247), .Z(n9249) );
  XOR U8614 ( .A(n9258), .B(n9259), .Z(n9247) );
  AND U8615 ( .A(n2142), .B(n9260), .Z(n9259) );
  XOR U8616 ( .A(p_input[1749]), .B(n9258), .Z(n9260) );
  XOR U8617 ( .A(n9261), .B(n9262), .Z(n9258) );
  AND U8618 ( .A(n2146), .B(n9263), .Z(n9262) );
  IV U8619 ( .A(n9255), .Z(n9257) );
  XOR U8620 ( .A(n9264), .B(n9265), .Z(n9255) );
  AND U8621 ( .A(n2150), .B(n9266), .Z(n9265) );
  XOR U8622 ( .A(n9267), .B(n9268), .Z(n9253) );
  AND U8623 ( .A(n2154), .B(n9266), .Z(n9268) );
  XNOR U8624 ( .A(n9267), .B(n9264), .Z(n9266) );
  XOR U8625 ( .A(n9269), .B(n9270), .Z(n9264) );
  AND U8626 ( .A(n2157), .B(n9263), .Z(n9270) );
  XNOR U8627 ( .A(n9271), .B(n9261), .Z(n9263) );
  XOR U8628 ( .A(n9272), .B(n9273), .Z(n9261) );
  AND U8629 ( .A(n2161), .B(n9274), .Z(n9273) );
  XOR U8630 ( .A(p_input[1765]), .B(n9272), .Z(n9274) );
  XOR U8631 ( .A(n9275), .B(n9276), .Z(n9272) );
  AND U8632 ( .A(n2165), .B(n9277), .Z(n9276) );
  IV U8633 ( .A(n9269), .Z(n9271) );
  XOR U8634 ( .A(n9278), .B(n9279), .Z(n9269) );
  AND U8635 ( .A(n2169), .B(n9280), .Z(n9279) );
  XOR U8636 ( .A(n9281), .B(n9282), .Z(n9267) );
  AND U8637 ( .A(n2173), .B(n9280), .Z(n9282) );
  XNOR U8638 ( .A(n9281), .B(n9278), .Z(n9280) );
  XOR U8639 ( .A(n9283), .B(n9284), .Z(n9278) );
  AND U8640 ( .A(n2176), .B(n9277), .Z(n9284) );
  XNOR U8641 ( .A(n9285), .B(n9275), .Z(n9277) );
  XOR U8642 ( .A(n9286), .B(n9287), .Z(n9275) );
  AND U8643 ( .A(n2180), .B(n9288), .Z(n9287) );
  XOR U8644 ( .A(p_input[1781]), .B(n9286), .Z(n9288) );
  XOR U8645 ( .A(n9289), .B(n9290), .Z(n9286) );
  AND U8646 ( .A(n2184), .B(n9291), .Z(n9290) );
  IV U8647 ( .A(n9283), .Z(n9285) );
  XOR U8648 ( .A(n9292), .B(n9293), .Z(n9283) );
  AND U8649 ( .A(n2188), .B(n9294), .Z(n9293) );
  XOR U8650 ( .A(n9295), .B(n9296), .Z(n9281) );
  AND U8651 ( .A(n2192), .B(n9294), .Z(n9296) );
  XNOR U8652 ( .A(n9295), .B(n9292), .Z(n9294) );
  XOR U8653 ( .A(n9297), .B(n9298), .Z(n9292) );
  AND U8654 ( .A(n2195), .B(n9291), .Z(n9298) );
  XNOR U8655 ( .A(n9299), .B(n9289), .Z(n9291) );
  XOR U8656 ( .A(n9300), .B(n9301), .Z(n9289) );
  AND U8657 ( .A(n2199), .B(n9302), .Z(n9301) );
  XOR U8658 ( .A(p_input[1797]), .B(n9300), .Z(n9302) );
  XOR U8659 ( .A(n9303), .B(n9304), .Z(n9300) );
  AND U8660 ( .A(n2203), .B(n9305), .Z(n9304) );
  IV U8661 ( .A(n9297), .Z(n9299) );
  XOR U8662 ( .A(n9306), .B(n9307), .Z(n9297) );
  AND U8663 ( .A(n2207), .B(n9308), .Z(n9307) );
  XOR U8664 ( .A(n9309), .B(n9310), .Z(n9295) );
  AND U8665 ( .A(n2211), .B(n9308), .Z(n9310) );
  XNOR U8666 ( .A(n9309), .B(n9306), .Z(n9308) );
  XOR U8667 ( .A(n9311), .B(n9312), .Z(n9306) );
  AND U8668 ( .A(n2214), .B(n9305), .Z(n9312) );
  XNOR U8669 ( .A(n9313), .B(n9303), .Z(n9305) );
  XOR U8670 ( .A(n9314), .B(n9315), .Z(n9303) );
  AND U8671 ( .A(n2218), .B(n9316), .Z(n9315) );
  XOR U8672 ( .A(p_input[1813]), .B(n9314), .Z(n9316) );
  XOR U8673 ( .A(n9317), .B(n9318), .Z(n9314) );
  AND U8674 ( .A(n2222), .B(n9319), .Z(n9318) );
  IV U8675 ( .A(n9311), .Z(n9313) );
  XOR U8676 ( .A(n9320), .B(n9321), .Z(n9311) );
  AND U8677 ( .A(n2226), .B(n9322), .Z(n9321) );
  XOR U8678 ( .A(n9323), .B(n9324), .Z(n9309) );
  AND U8679 ( .A(n2230), .B(n9322), .Z(n9324) );
  XNOR U8680 ( .A(n9323), .B(n9320), .Z(n9322) );
  XOR U8681 ( .A(n9325), .B(n9326), .Z(n9320) );
  AND U8682 ( .A(n2233), .B(n9319), .Z(n9326) );
  XNOR U8683 ( .A(n9327), .B(n9317), .Z(n9319) );
  XOR U8684 ( .A(n9328), .B(n9329), .Z(n9317) );
  AND U8685 ( .A(n2237), .B(n9330), .Z(n9329) );
  XOR U8686 ( .A(p_input[1829]), .B(n9328), .Z(n9330) );
  XOR U8687 ( .A(n9331), .B(n9332), .Z(n9328) );
  AND U8688 ( .A(n2241), .B(n9333), .Z(n9332) );
  IV U8689 ( .A(n9325), .Z(n9327) );
  XOR U8690 ( .A(n9334), .B(n9335), .Z(n9325) );
  AND U8691 ( .A(n2245), .B(n9336), .Z(n9335) );
  XOR U8692 ( .A(n9337), .B(n9338), .Z(n9323) );
  AND U8693 ( .A(n2249), .B(n9336), .Z(n9338) );
  XNOR U8694 ( .A(n9337), .B(n9334), .Z(n9336) );
  XOR U8695 ( .A(n9339), .B(n9340), .Z(n9334) );
  AND U8696 ( .A(n2252), .B(n9333), .Z(n9340) );
  XNOR U8697 ( .A(n9341), .B(n9331), .Z(n9333) );
  XOR U8698 ( .A(n9342), .B(n9343), .Z(n9331) );
  AND U8699 ( .A(n2256), .B(n9344), .Z(n9343) );
  XOR U8700 ( .A(p_input[1845]), .B(n9342), .Z(n9344) );
  XOR U8701 ( .A(n9345), .B(n9346), .Z(n9342) );
  AND U8702 ( .A(n2260), .B(n9347), .Z(n9346) );
  IV U8703 ( .A(n9339), .Z(n9341) );
  XOR U8704 ( .A(n9348), .B(n9349), .Z(n9339) );
  AND U8705 ( .A(n2264), .B(n9350), .Z(n9349) );
  XOR U8706 ( .A(n9351), .B(n9352), .Z(n9337) );
  AND U8707 ( .A(n2268), .B(n9350), .Z(n9352) );
  XNOR U8708 ( .A(n9351), .B(n9348), .Z(n9350) );
  XOR U8709 ( .A(n9353), .B(n9354), .Z(n9348) );
  AND U8710 ( .A(n2271), .B(n9347), .Z(n9354) );
  XNOR U8711 ( .A(n9355), .B(n9345), .Z(n9347) );
  XOR U8712 ( .A(n9356), .B(n9357), .Z(n9345) );
  AND U8713 ( .A(n2275), .B(n9358), .Z(n9357) );
  XOR U8714 ( .A(p_input[1861]), .B(n9356), .Z(n9358) );
  XOR U8715 ( .A(n9359), .B(n9360), .Z(n9356) );
  AND U8716 ( .A(n2279), .B(n9361), .Z(n9360) );
  IV U8717 ( .A(n9353), .Z(n9355) );
  XOR U8718 ( .A(n9362), .B(n9363), .Z(n9353) );
  AND U8719 ( .A(n2283), .B(n9364), .Z(n9363) );
  XOR U8720 ( .A(n9365), .B(n9366), .Z(n9351) );
  AND U8721 ( .A(n2287), .B(n9364), .Z(n9366) );
  XNOR U8722 ( .A(n9365), .B(n9362), .Z(n9364) );
  XOR U8723 ( .A(n9367), .B(n9368), .Z(n9362) );
  AND U8724 ( .A(n2290), .B(n9361), .Z(n9368) );
  XNOR U8725 ( .A(n9369), .B(n9359), .Z(n9361) );
  XOR U8726 ( .A(n9370), .B(n9371), .Z(n9359) );
  AND U8727 ( .A(n2294), .B(n9372), .Z(n9371) );
  XOR U8728 ( .A(p_input[1877]), .B(n9370), .Z(n9372) );
  XOR U8729 ( .A(n9373), .B(n9374), .Z(n9370) );
  AND U8730 ( .A(n2298), .B(n9375), .Z(n9374) );
  IV U8731 ( .A(n9367), .Z(n9369) );
  XOR U8732 ( .A(n9376), .B(n9377), .Z(n9367) );
  AND U8733 ( .A(n2302), .B(n9378), .Z(n9377) );
  XOR U8734 ( .A(n9379), .B(n9380), .Z(n9365) );
  AND U8735 ( .A(n2306), .B(n9378), .Z(n9380) );
  XNOR U8736 ( .A(n9379), .B(n9376), .Z(n9378) );
  XOR U8737 ( .A(n9381), .B(n9382), .Z(n9376) );
  AND U8738 ( .A(n2309), .B(n9375), .Z(n9382) );
  XNOR U8739 ( .A(n9383), .B(n9373), .Z(n9375) );
  XOR U8740 ( .A(n9384), .B(n9385), .Z(n9373) );
  AND U8741 ( .A(n2313), .B(n9386), .Z(n9385) );
  XOR U8742 ( .A(p_input[1893]), .B(n9384), .Z(n9386) );
  XOR U8743 ( .A(n9387), .B(n9388), .Z(n9384) );
  AND U8744 ( .A(n2317), .B(n9389), .Z(n9388) );
  IV U8745 ( .A(n9381), .Z(n9383) );
  XOR U8746 ( .A(n9390), .B(n9391), .Z(n9381) );
  AND U8747 ( .A(n2321), .B(n9392), .Z(n9391) );
  XOR U8748 ( .A(n9393), .B(n9394), .Z(n9379) );
  AND U8749 ( .A(n2325), .B(n9392), .Z(n9394) );
  XNOR U8750 ( .A(n9393), .B(n9390), .Z(n9392) );
  XOR U8751 ( .A(n9395), .B(n9396), .Z(n9390) );
  AND U8752 ( .A(n2328), .B(n9389), .Z(n9396) );
  XNOR U8753 ( .A(n9397), .B(n9387), .Z(n9389) );
  XOR U8754 ( .A(n9398), .B(n9399), .Z(n9387) );
  AND U8755 ( .A(n2332), .B(n9400), .Z(n9399) );
  XOR U8756 ( .A(p_input[1909]), .B(n9398), .Z(n9400) );
  XOR U8757 ( .A(n9401), .B(n9402), .Z(n9398) );
  AND U8758 ( .A(n2336), .B(n9403), .Z(n9402) );
  IV U8759 ( .A(n9395), .Z(n9397) );
  XOR U8760 ( .A(n9404), .B(n9405), .Z(n9395) );
  AND U8761 ( .A(n2340), .B(n9406), .Z(n9405) );
  XOR U8762 ( .A(n9407), .B(n9408), .Z(n9393) );
  AND U8763 ( .A(n2344), .B(n9406), .Z(n9408) );
  XNOR U8764 ( .A(n9407), .B(n9404), .Z(n9406) );
  XOR U8765 ( .A(n9409), .B(n9410), .Z(n9404) );
  AND U8766 ( .A(n2347), .B(n9403), .Z(n9410) );
  XNOR U8767 ( .A(n9411), .B(n9401), .Z(n9403) );
  XOR U8768 ( .A(n9412), .B(n9413), .Z(n9401) );
  AND U8769 ( .A(n2351), .B(n9414), .Z(n9413) );
  XOR U8770 ( .A(p_input[1925]), .B(n9412), .Z(n9414) );
  XOR U8771 ( .A(n9415), .B(n9416), .Z(n9412) );
  AND U8772 ( .A(n2355), .B(n9417), .Z(n9416) );
  IV U8773 ( .A(n9409), .Z(n9411) );
  XOR U8774 ( .A(n9418), .B(n9419), .Z(n9409) );
  AND U8775 ( .A(n2359), .B(n9420), .Z(n9419) );
  XOR U8776 ( .A(n9421), .B(n9422), .Z(n9407) );
  AND U8777 ( .A(n2363), .B(n9420), .Z(n9422) );
  XNOR U8778 ( .A(n9421), .B(n9418), .Z(n9420) );
  XOR U8779 ( .A(n9423), .B(n9424), .Z(n9418) );
  AND U8780 ( .A(n2366), .B(n9417), .Z(n9424) );
  XNOR U8781 ( .A(n9425), .B(n9415), .Z(n9417) );
  XOR U8782 ( .A(n9426), .B(n9427), .Z(n9415) );
  AND U8783 ( .A(n2370), .B(n9428), .Z(n9427) );
  XOR U8784 ( .A(p_input[1941]), .B(n9426), .Z(n9428) );
  XOR U8785 ( .A(n9429), .B(n9430), .Z(n9426) );
  AND U8786 ( .A(n2374), .B(n9431), .Z(n9430) );
  IV U8787 ( .A(n9423), .Z(n9425) );
  XOR U8788 ( .A(n9432), .B(n9433), .Z(n9423) );
  AND U8789 ( .A(n2378), .B(n9434), .Z(n9433) );
  XOR U8790 ( .A(n9435), .B(n9436), .Z(n9421) );
  AND U8791 ( .A(n2382), .B(n9434), .Z(n9436) );
  XNOR U8792 ( .A(n9435), .B(n9432), .Z(n9434) );
  XOR U8793 ( .A(n9437), .B(n9438), .Z(n9432) );
  AND U8794 ( .A(n2385), .B(n9431), .Z(n9438) );
  XNOR U8795 ( .A(n9439), .B(n9429), .Z(n9431) );
  XOR U8796 ( .A(n9440), .B(n9441), .Z(n9429) );
  AND U8797 ( .A(n2389), .B(n9442), .Z(n9441) );
  XOR U8798 ( .A(p_input[1957]), .B(n9440), .Z(n9442) );
  XOR U8799 ( .A(n9443), .B(n9444), .Z(n9440) );
  AND U8800 ( .A(n2393), .B(n9445), .Z(n9444) );
  IV U8801 ( .A(n9437), .Z(n9439) );
  XOR U8802 ( .A(n9446), .B(n9447), .Z(n9437) );
  AND U8803 ( .A(n2397), .B(n9448), .Z(n9447) );
  XOR U8804 ( .A(n9449), .B(n9450), .Z(n9435) );
  AND U8805 ( .A(n2401), .B(n9448), .Z(n9450) );
  XNOR U8806 ( .A(n9449), .B(n9446), .Z(n9448) );
  XOR U8807 ( .A(n9451), .B(n9452), .Z(n9446) );
  AND U8808 ( .A(n2404), .B(n9445), .Z(n9452) );
  XNOR U8809 ( .A(n9453), .B(n9443), .Z(n9445) );
  XOR U8810 ( .A(n9454), .B(n9455), .Z(n9443) );
  AND U8811 ( .A(n2408), .B(n9456), .Z(n9455) );
  XOR U8812 ( .A(p_input[1973]), .B(n9454), .Z(n9456) );
  XOR U8813 ( .A(n9457), .B(n9458), .Z(n9454) );
  AND U8814 ( .A(n2412), .B(n9459), .Z(n9458) );
  IV U8815 ( .A(n9451), .Z(n9453) );
  XOR U8816 ( .A(n9460), .B(n9461), .Z(n9451) );
  AND U8817 ( .A(n2416), .B(n9462), .Z(n9461) );
  XOR U8818 ( .A(n9463), .B(n9464), .Z(n9449) );
  AND U8819 ( .A(n2420), .B(n9462), .Z(n9464) );
  XNOR U8820 ( .A(n9463), .B(n9460), .Z(n9462) );
  XOR U8821 ( .A(n9465), .B(n9466), .Z(n9460) );
  AND U8822 ( .A(n2423), .B(n9459), .Z(n9466) );
  XNOR U8823 ( .A(n9467), .B(n9457), .Z(n9459) );
  XOR U8824 ( .A(n9468), .B(n9469), .Z(n9457) );
  AND U8825 ( .A(n2427), .B(n9470), .Z(n9469) );
  XOR U8826 ( .A(p_input[1989]), .B(n9468), .Z(n9470) );
  XOR U8827 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n9471), 
        .Z(n9468) );
  AND U8828 ( .A(n2430), .B(n9472), .Z(n9471) );
  IV U8829 ( .A(n9465), .Z(n9467) );
  XOR U8830 ( .A(n9473), .B(n9474), .Z(n9465) );
  AND U8831 ( .A(n2434), .B(n9475), .Z(n9474) );
  XOR U8832 ( .A(n9476), .B(n9477), .Z(n9463) );
  AND U8833 ( .A(n2438), .B(n9475), .Z(n9477) );
  XNOR U8834 ( .A(n9476), .B(n9473), .Z(n9475) );
  XNOR U8835 ( .A(n9478), .B(n9479), .Z(n9473) );
  AND U8836 ( .A(n2441), .B(n9472), .Z(n9479) );
  XNOR U8837 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n9478), 
        .Z(n9472) );
  XNOR U8838 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n9480), 
        .Z(n9478) );
  AND U8839 ( .A(n2443), .B(n9481), .Z(n9480) );
  XNOR U8840 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n9482), .Z(n9476) );
  AND U8841 ( .A(n2446), .B(n9481), .Z(n9482) );
  XOR U8842 ( .A(n9483), .B(n9484), .Z(n9481) );
  XOR U8843 ( .A(n11), .B(n9485), .Z(o[20]) );
  AND U8844 ( .A(n62), .B(n9486), .Z(n11) );
  XOR U8845 ( .A(n12), .B(n9485), .Z(n9486) );
  XOR U8846 ( .A(n9487), .B(n37), .Z(n9485) );
  AND U8847 ( .A(n65), .B(n9488), .Z(n37) );
  XNOR U8848 ( .A(n9489), .B(n38), .Z(n9488) );
  XOR U8849 ( .A(n9490), .B(n9491), .Z(n38) );
  AND U8850 ( .A(n70), .B(n9492), .Z(n9491) );
  XOR U8851 ( .A(p_input[4]), .B(n9490), .Z(n9492) );
  XOR U8852 ( .A(n9493), .B(n9494), .Z(n9490) );
  AND U8853 ( .A(n74), .B(n9495), .Z(n9494) );
  IV U8854 ( .A(n9487), .Z(n9489) );
  XOR U8855 ( .A(n9496), .B(n9497), .Z(n9487) );
  AND U8856 ( .A(n78), .B(n9498), .Z(n9497) );
  XOR U8857 ( .A(n9499), .B(n9500), .Z(n12) );
  AND U8858 ( .A(n82), .B(n9498), .Z(n9500) );
  XNOR U8859 ( .A(n9501), .B(n9496), .Z(n9498) );
  XOR U8860 ( .A(n9502), .B(n9503), .Z(n9496) );
  AND U8861 ( .A(n86), .B(n9495), .Z(n9503) );
  XNOR U8862 ( .A(n9504), .B(n9493), .Z(n9495) );
  XOR U8863 ( .A(n9505), .B(n9506), .Z(n9493) );
  AND U8864 ( .A(n90), .B(n9507), .Z(n9506) );
  XOR U8865 ( .A(p_input[20]), .B(n9505), .Z(n9507) );
  XOR U8866 ( .A(n9508), .B(n9509), .Z(n9505) );
  AND U8867 ( .A(n94), .B(n9510), .Z(n9509) );
  IV U8868 ( .A(n9502), .Z(n9504) );
  XOR U8869 ( .A(n9511), .B(n9512), .Z(n9502) );
  AND U8870 ( .A(n98), .B(n9513), .Z(n9512) );
  IV U8871 ( .A(n9499), .Z(n9501) );
  XNOR U8872 ( .A(n9514), .B(n9515), .Z(n9499) );
  AND U8873 ( .A(n102), .B(n9513), .Z(n9515) );
  XNOR U8874 ( .A(n9514), .B(n9511), .Z(n9513) );
  XOR U8875 ( .A(n9516), .B(n9517), .Z(n9511) );
  AND U8876 ( .A(n105), .B(n9510), .Z(n9517) );
  XNOR U8877 ( .A(n9518), .B(n9508), .Z(n9510) );
  XOR U8878 ( .A(n9519), .B(n9520), .Z(n9508) );
  AND U8879 ( .A(n109), .B(n9521), .Z(n9520) );
  XOR U8880 ( .A(p_input[36]), .B(n9519), .Z(n9521) );
  XOR U8881 ( .A(n9522), .B(n9523), .Z(n9519) );
  AND U8882 ( .A(n113), .B(n9524), .Z(n9523) );
  IV U8883 ( .A(n9516), .Z(n9518) );
  XOR U8884 ( .A(n9525), .B(n9526), .Z(n9516) );
  AND U8885 ( .A(n117), .B(n9527), .Z(n9526) );
  XOR U8886 ( .A(n9528), .B(n9529), .Z(n9514) );
  AND U8887 ( .A(n121), .B(n9527), .Z(n9529) );
  XNOR U8888 ( .A(n9528), .B(n9525), .Z(n9527) );
  XOR U8889 ( .A(n9530), .B(n9531), .Z(n9525) );
  AND U8890 ( .A(n124), .B(n9524), .Z(n9531) );
  XNOR U8891 ( .A(n9532), .B(n9522), .Z(n9524) );
  XOR U8892 ( .A(n9533), .B(n9534), .Z(n9522) );
  AND U8893 ( .A(n128), .B(n9535), .Z(n9534) );
  XOR U8894 ( .A(p_input[52]), .B(n9533), .Z(n9535) );
  XOR U8895 ( .A(n9536), .B(n9537), .Z(n9533) );
  AND U8896 ( .A(n132), .B(n9538), .Z(n9537) );
  IV U8897 ( .A(n9530), .Z(n9532) );
  XOR U8898 ( .A(n9539), .B(n9540), .Z(n9530) );
  AND U8899 ( .A(n136), .B(n9541), .Z(n9540) );
  XOR U8900 ( .A(n9542), .B(n9543), .Z(n9528) );
  AND U8901 ( .A(n140), .B(n9541), .Z(n9543) );
  XNOR U8902 ( .A(n9542), .B(n9539), .Z(n9541) );
  XOR U8903 ( .A(n9544), .B(n9545), .Z(n9539) );
  AND U8904 ( .A(n143), .B(n9538), .Z(n9545) );
  XNOR U8905 ( .A(n9546), .B(n9536), .Z(n9538) );
  XOR U8906 ( .A(n9547), .B(n9548), .Z(n9536) );
  AND U8907 ( .A(n147), .B(n9549), .Z(n9548) );
  XOR U8908 ( .A(p_input[68]), .B(n9547), .Z(n9549) );
  XOR U8909 ( .A(n9550), .B(n9551), .Z(n9547) );
  AND U8910 ( .A(n151), .B(n9552), .Z(n9551) );
  IV U8911 ( .A(n9544), .Z(n9546) );
  XOR U8912 ( .A(n9553), .B(n9554), .Z(n9544) );
  AND U8913 ( .A(n155), .B(n9555), .Z(n9554) );
  XOR U8914 ( .A(n9556), .B(n9557), .Z(n9542) );
  AND U8915 ( .A(n159), .B(n9555), .Z(n9557) );
  XNOR U8916 ( .A(n9556), .B(n9553), .Z(n9555) );
  XOR U8917 ( .A(n9558), .B(n9559), .Z(n9553) );
  AND U8918 ( .A(n162), .B(n9552), .Z(n9559) );
  XNOR U8919 ( .A(n9560), .B(n9550), .Z(n9552) );
  XOR U8920 ( .A(n9561), .B(n9562), .Z(n9550) );
  AND U8921 ( .A(n166), .B(n9563), .Z(n9562) );
  XOR U8922 ( .A(p_input[84]), .B(n9561), .Z(n9563) );
  XOR U8923 ( .A(n9564), .B(n9565), .Z(n9561) );
  AND U8924 ( .A(n170), .B(n9566), .Z(n9565) );
  IV U8925 ( .A(n9558), .Z(n9560) );
  XOR U8926 ( .A(n9567), .B(n9568), .Z(n9558) );
  AND U8927 ( .A(n174), .B(n9569), .Z(n9568) );
  XOR U8928 ( .A(n9570), .B(n9571), .Z(n9556) );
  AND U8929 ( .A(n178), .B(n9569), .Z(n9571) );
  XNOR U8930 ( .A(n9570), .B(n9567), .Z(n9569) );
  XOR U8931 ( .A(n9572), .B(n9573), .Z(n9567) );
  AND U8932 ( .A(n181), .B(n9566), .Z(n9573) );
  XNOR U8933 ( .A(n9574), .B(n9564), .Z(n9566) );
  XOR U8934 ( .A(n9575), .B(n9576), .Z(n9564) );
  AND U8935 ( .A(n185), .B(n9577), .Z(n9576) );
  XOR U8936 ( .A(p_input[100]), .B(n9575), .Z(n9577) );
  XOR U8937 ( .A(n9578), .B(n9579), .Z(n9575) );
  AND U8938 ( .A(n189), .B(n9580), .Z(n9579) );
  IV U8939 ( .A(n9572), .Z(n9574) );
  XOR U8940 ( .A(n9581), .B(n9582), .Z(n9572) );
  AND U8941 ( .A(n193), .B(n9583), .Z(n9582) );
  XOR U8942 ( .A(n9584), .B(n9585), .Z(n9570) );
  AND U8943 ( .A(n197), .B(n9583), .Z(n9585) );
  XNOR U8944 ( .A(n9584), .B(n9581), .Z(n9583) );
  XOR U8945 ( .A(n9586), .B(n9587), .Z(n9581) );
  AND U8946 ( .A(n200), .B(n9580), .Z(n9587) );
  XNOR U8947 ( .A(n9588), .B(n9578), .Z(n9580) );
  XOR U8948 ( .A(n9589), .B(n9590), .Z(n9578) );
  AND U8949 ( .A(n204), .B(n9591), .Z(n9590) );
  XOR U8950 ( .A(p_input[116]), .B(n9589), .Z(n9591) );
  XOR U8951 ( .A(n9592), .B(n9593), .Z(n9589) );
  AND U8952 ( .A(n208), .B(n9594), .Z(n9593) );
  IV U8953 ( .A(n9586), .Z(n9588) );
  XOR U8954 ( .A(n9595), .B(n9596), .Z(n9586) );
  AND U8955 ( .A(n212), .B(n9597), .Z(n9596) );
  XOR U8956 ( .A(n9598), .B(n9599), .Z(n9584) );
  AND U8957 ( .A(n216), .B(n9597), .Z(n9599) );
  XNOR U8958 ( .A(n9598), .B(n9595), .Z(n9597) );
  XOR U8959 ( .A(n9600), .B(n9601), .Z(n9595) );
  AND U8960 ( .A(n219), .B(n9594), .Z(n9601) );
  XNOR U8961 ( .A(n9602), .B(n9592), .Z(n9594) );
  XOR U8962 ( .A(n9603), .B(n9604), .Z(n9592) );
  AND U8963 ( .A(n223), .B(n9605), .Z(n9604) );
  XOR U8964 ( .A(p_input[132]), .B(n9603), .Z(n9605) );
  XOR U8965 ( .A(n9606), .B(n9607), .Z(n9603) );
  AND U8966 ( .A(n227), .B(n9608), .Z(n9607) );
  IV U8967 ( .A(n9600), .Z(n9602) );
  XOR U8968 ( .A(n9609), .B(n9610), .Z(n9600) );
  AND U8969 ( .A(n231), .B(n9611), .Z(n9610) );
  XOR U8970 ( .A(n9612), .B(n9613), .Z(n9598) );
  AND U8971 ( .A(n235), .B(n9611), .Z(n9613) );
  XNOR U8972 ( .A(n9612), .B(n9609), .Z(n9611) );
  XOR U8973 ( .A(n9614), .B(n9615), .Z(n9609) );
  AND U8974 ( .A(n238), .B(n9608), .Z(n9615) );
  XNOR U8975 ( .A(n9616), .B(n9606), .Z(n9608) );
  XOR U8976 ( .A(n9617), .B(n9618), .Z(n9606) );
  AND U8977 ( .A(n242), .B(n9619), .Z(n9618) );
  XOR U8978 ( .A(p_input[148]), .B(n9617), .Z(n9619) );
  XOR U8979 ( .A(n9620), .B(n9621), .Z(n9617) );
  AND U8980 ( .A(n246), .B(n9622), .Z(n9621) );
  IV U8981 ( .A(n9614), .Z(n9616) );
  XOR U8982 ( .A(n9623), .B(n9624), .Z(n9614) );
  AND U8983 ( .A(n250), .B(n9625), .Z(n9624) );
  XOR U8984 ( .A(n9626), .B(n9627), .Z(n9612) );
  AND U8985 ( .A(n254), .B(n9625), .Z(n9627) );
  XNOR U8986 ( .A(n9626), .B(n9623), .Z(n9625) );
  XOR U8987 ( .A(n9628), .B(n9629), .Z(n9623) );
  AND U8988 ( .A(n257), .B(n9622), .Z(n9629) );
  XNOR U8989 ( .A(n9630), .B(n9620), .Z(n9622) );
  XOR U8990 ( .A(n9631), .B(n9632), .Z(n9620) );
  AND U8991 ( .A(n261), .B(n9633), .Z(n9632) );
  XOR U8992 ( .A(p_input[164]), .B(n9631), .Z(n9633) );
  XOR U8993 ( .A(n9634), .B(n9635), .Z(n9631) );
  AND U8994 ( .A(n265), .B(n9636), .Z(n9635) );
  IV U8995 ( .A(n9628), .Z(n9630) );
  XOR U8996 ( .A(n9637), .B(n9638), .Z(n9628) );
  AND U8997 ( .A(n269), .B(n9639), .Z(n9638) );
  XOR U8998 ( .A(n9640), .B(n9641), .Z(n9626) );
  AND U8999 ( .A(n273), .B(n9639), .Z(n9641) );
  XNOR U9000 ( .A(n9640), .B(n9637), .Z(n9639) );
  XOR U9001 ( .A(n9642), .B(n9643), .Z(n9637) );
  AND U9002 ( .A(n276), .B(n9636), .Z(n9643) );
  XNOR U9003 ( .A(n9644), .B(n9634), .Z(n9636) );
  XOR U9004 ( .A(n9645), .B(n9646), .Z(n9634) );
  AND U9005 ( .A(n280), .B(n9647), .Z(n9646) );
  XOR U9006 ( .A(p_input[180]), .B(n9645), .Z(n9647) );
  XOR U9007 ( .A(n9648), .B(n9649), .Z(n9645) );
  AND U9008 ( .A(n284), .B(n9650), .Z(n9649) );
  IV U9009 ( .A(n9642), .Z(n9644) );
  XOR U9010 ( .A(n9651), .B(n9652), .Z(n9642) );
  AND U9011 ( .A(n288), .B(n9653), .Z(n9652) );
  XOR U9012 ( .A(n9654), .B(n9655), .Z(n9640) );
  AND U9013 ( .A(n292), .B(n9653), .Z(n9655) );
  XNOR U9014 ( .A(n9654), .B(n9651), .Z(n9653) );
  XOR U9015 ( .A(n9656), .B(n9657), .Z(n9651) );
  AND U9016 ( .A(n295), .B(n9650), .Z(n9657) );
  XNOR U9017 ( .A(n9658), .B(n9648), .Z(n9650) );
  XOR U9018 ( .A(n9659), .B(n9660), .Z(n9648) );
  AND U9019 ( .A(n299), .B(n9661), .Z(n9660) );
  XOR U9020 ( .A(p_input[196]), .B(n9659), .Z(n9661) );
  XOR U9021 ( .A(n9662), .B(n9663), .Z(n9659) );
  AND U9022 ( .A(n303), .B(n9664), .Z(n9663) );
  IV U9023 ( .A(n9656), .Z(n9658) );
  XOR U9024 ( .A(n9665), .B(n9666), .Z(n9656) );
  AND U9025 ( .A(n307), .B(n9667), .Z(n9666) );
  XOR U9026 ( .A(n9668), .B(n9669), .Z(n9654) );
  AND U9027 ( .A(n311), .B(n9667), .Z(n9669) );
  XNOR U9028 ( .A(n9668), .B(n9665), .Z(n9667) );
  XOR U9029 ( .A(n9670), .B(n9671), .Z(n9665) );
  AND U9030 ( .A(n314), .B(n9664), .Z(n9671) );
  XNOR U9031 ( .A(n9672), .B(n9662), .Z(n9664) );
  XOR U9032 ( .A(n9673), .B(n9674), .Z(n9662) );
  AND U9033 ( .A(n318), .B(n9675), .Z(n9674) );
  XOR U9034 ( .A(p_input[212]), .B(n9673), .Z(n9675) );
  XOR U9035 ( .A(n9676), .B(n9677), .Z(n9673) );
  AND U9036 ( .A(n322), .B(n9678), .Z(n9677) );
  IV U9037 ( .A(n9670), .Z(n9672) );
  XOR U9038 ( .A(n9679), .B(n9680), .Z(n9670) );
  AND U9039 ( .A(n326), .B(n9681), .Z(n9680) );
  XOR U9040 ( .A(n9682), .B(n9683), .Z(n9668) );
  AND U9041 ( .A(n330), .B(n9681), .Z(n9683) );
  XNOR U9042 ( .A(n9682), .B(n9679), .Z(n9681) );
  XOR U9043 ( .A(n9684), .B(n9685), .Z(n9679) );
  AND U9044 ( .A(n333), .B(n9678), .Z(n9685) );
  XNOR U9045 ( .A(n9686), .B(n9676), .Z(n9678) );
  XOR U9046 ( .A(n9687), .B(n9688), .Z(n9676) );
  AND U9047 ( .A(n337), .B(n9689), .Z(n9688) );
  XOR U9048 ( .A(p_input[228]), .B(n9687), .Z(n9689) );
  XOR U9049 ( .A(n9690), .B(n9691), .Z(n9687) );
  AND U9050 ( .A(n341), .B(n9692), .Z(n9691) );
  IV U9051 ( .A(n9684), .Z(n9686) );
  XOR U9052 ( .A(n9693), .B(n9694), .Z(n9684) );
  AND U9053 ( .A(n345), .B(n9695), .Z(n9694) );
  XOR U9054 ( .A(n9696), .B(n9697), .Z(n9682) );
  AND U9055 ( .A(n349), .B(n9695), .Z(n9697) );
  XNOR U9056 ( .A(n9696), .B(n9693), .Z(n9695) );
  XOR U9057 ( .A(n9698), .B(n9699), .Z(n9693) );
  AND U9058 ( .A(n352), .B(n9692), .Z(n9699) );
  XNOR U9059 ( .A(n9700), .B(n9690), .Z(n9692) );
  XOR U9060 ( .A(n9701), .B(n9702), .Z(n9690) );
  AND U9061 ( .A(n356), .B(n9703), .Z(n9702) );
  XOR U9062 ( .A(p_input[244]), .B(n9701), .Z(n9703) );
  XOR U9063 ( .A(n9704), .B(n9705), .Z(n9701) );
  AND U9064 ( .A(n360), .B(n9706), .Z(n9705) );
  IV U9065 ( .A(n9698), .Z(n9700) );
  XOR U9066 ( .A(n9707), .B(n9708), .Z(n9698) );
  AND U9067 ( .A(n364), .B(n9709), .Z(n9708) );
  XOR U9068 ( .A(n9710), .B(n9711), .Z(n9696) );
  AND U9069 ( .A(n368), .B(n9709), .Z(n9711) );
  XNOR U9070 ( .A(n9710), .B(n9707), .Z(n9709) );
  XOR U9071 ( .A(n9712), .B(n9713), .Z(n9707) );
  AND U9072 ( .A(n371), .B(n9706), .Z(n9713) );
  XNOR U9073 ( .A(n9714), .B(n9704), .Z(n9706) );
  XOR U9074 ( .A(n9715), .B(n9716), .Z(n9704) );
  AND U9075 ( .A(n375), .B(n9717), .Z(n9716) );
  XOR U9076 ( .A(p_input[260]), .B(n9715), .Z(n9717) );
  XOR U9077 ( .A(n9718), .B(n9719), .Z(n9715) );
  AND U9078 ( .A(n379), .B(n9720), .Z(n9719) );
  IV U9079 ( .A(n9712), .Z(n9714) );
  XOR U9080 ( .A(n9721), .B(n9722), .Z(n9712) );
  AND U9081 ( .A(n383), .B(n9723), .Z(n9722) );
  XOR U9082 ( .A(n9724), .B(n9725), .Z(n9710) );
  AND U9083 ( .A(n387), .B(n9723), .Z(n9725) );
  XNOR U9084 ( .A(n9724), .B(n9721), .Z(n9723) );
  XOR U9085 ( .A(n9726), .B(n9727), .Z(n9721) );
  AND U9086 ( .A(n390), .B(n9720), .Z(n9727) );
  XNOR U9087 ( .A(n9728), .B(n9718), .Z(n9720) );
  XOR U9088 ( .A(n9729), .B(n9730), .Z(n9718) );
  AND U9089 ( .A(n394), .B(n9731), .Z(n9730) );
  XOR U9090 ( .A(p_input[276]), .B(n9729), .Z(n9731) );
  XOR U9091 ( .A(n9732), .B(n9733), .Z(n9729) );
  AND U9092 ( .A(n398), .B(n9734), .Z(n9733) );
  IV U9093 ( .A(n9726), .Z(n9728) );
  XOR U9094 ( .A(n9735), .B(n9736), .Z(n9726) );
  AND U9095 ( .A(n402), .B(n9737), .Z(n9736) );
  XOR U9096 ( .A(n9738), .B(n9739), .Z(n9724) );
  AND U9097 ( .A(n406), .B(n9737), .Z(n9739) );
  XNOR U9098 ( .A(n9738), .B(n9735), .Z(n9737) );
  XOR U9099 ( .A(n9740), .B(n9741), .Z(n9735) );
  AND U9100 ( .A(n409), .B(n9734), .Z(n9741) );
  XNOR U9101 ( .A(n9742), .B(n9732), .Z(n9734) );
  XOR U9102 ( .A(n9743), .B(n9744), .Z(n9732) );
  AND U9103 ( .A(n413), .B(n9745), .Z(n9744) );
  XOR U9104 ( .A(p_input[292]), .B(n9743), .Z(n9745) );
  XOR U9105 ( .A(n9746), .B(n9747), .Z(n9743) );
  AND U9106 ( .A(n417), .B(n9748), .Z(n9747) );
  IV U9107 ( .A(n9740), .Z(n9742) );
  XOR U9108 ( .A(n9749), .B(n9750), .Z(n9740) );
  AND U9109 ( .A(n421), .B(n9751), .Z(n9750) );
  XOR U9110 ( .A(n9752), .B(n9753), .Z(n9738) );
  AND U9111 ( .A(n425), .B(n9751), .Z(n9753) );
  XNOR U9112 ( .A(n9752), .B(n9749), .Z(n9751) );
  XOR U9113 ( .A(n9754), .B(n9755), .Z(n9749) );
  AND U9114 ( .A(n428), .B(n9748), .Z(n9755) );
  XNOR U9115 ( .A(n9756), .B(n9746), .Z(n9748) );
  XOR U9116 ( .A(n9757), .B(n9758), .Z(n9746) );
  AND U9117 ( .A(n432), .B(n9759), .Z(n9758) );
  XOR U9118 ( .A(p_input[308]), .B(n9757), .Z(n9759) );
  XOR U9119 ( .A(n9760), .B(n9761), .Z(n9757) );
  AND U9120 ( .A(n436), .B(n9762), .Z(n9761) );
  IV U9121 ( .A(n9754), .Z(n9756) );
  XOR U9122 ( .A(n9763), .B(n9764), .Z(n9754) );
  AND U9123 ( .A(n440), .B(n9765), .Z(n9764) );
  XOR U9124 ( .A(n9766), .B(n9767), .Z(n9752) );
  AND U9125 ( .A(n444), .B(n9765), .Z(n9767) );
  XNOR U9126 ( .A(n9766), .B(n9763), .Z(n9765) );
  XOR U9127 ( .A(n9768), .B(n9769), .Z(n9763) );
  AND U9128 ( .A(n447), .B(n9762), .Z(n9769) );
  XNOR U9129 ( .A(n9770), .B(n9760), .Z(n9762) );
  XOR U9130 ( .A(n9771), .B(n9772), .Z(n9760) );
  AND U9131 ( .A(n451), .B(n9773), .Z(n9772) );
  XOR U9132 ( .A(p_input[324]), .B(n9771), .Z(n9773) );
  XOR U9133 ( .A(n9774), .B(n9775), .Z(n9771) );
  AND U9134 ( .A(n455), .B(n9776), .Z(n9775) );
  IV U9135 ( .A(n9768), .Z(n9770) );
  XOR U9136 ( .A(n9777), .B(n9778), .Z(n9768) );
  AND U9137 ( .A(n459), .B(n9779), .Z(n9778) );
  XOR U9138 ( .A(n9780), .B(n9781), .Z(n9766) );
  AND U9139 ( .A(n463), .B(n9779), .Z(n9781) );
  XNOR U9140 ( .A(n9780), .B(n9777), .Z(n9779) );
  XOR U9141 ( .A(n9782), .B(n9783), .Z(n9777) );
  AND U9142 ( .A(n466), .B(n9776), .Z(n9783) );
  XNOR U9143 ( .A(n9784), .B(n9774), .Z(n9776) );
  XOR U9144 ( .A(n9785), .B(n9786), .Z(n9774) );
  AND U9145 ( .A(n470), .B(n9787), .Z(n9786) );
  XOR U9146 ( .A(p_input[340]), .B(n9785), .Z(n9787) );
  XOR U9147 ( .A(n9788), .B(n9789), .Z(n9785) );
  AND U9148 ( .A(n474), .B(n9790), .Z(n9789) );
  IV U9149 ( .A(n9782), .Z(n9784) );
  XOR U9150 ( .A(n9791), .B(n9792), .Z(n9782) );
  AND U9151 ( .A(n478), .B(n9793), .Z(n9792) );
  XOR U9152 ( .A(n9794), .B(n9795), .Z(n9780) );
  AND U9153 ( .A(n482), .B(n9793), .Z(n9795) );
  XNOR U9154 ( .A(n9794), .B(n9791), .Z(n9793) );
  XOR U9155 ( .A(n9796), .B(n9797), .Z(n9791) );
  AND U9156 ( .A(n485), .B(n9790), .Z(n9797) );
  XNOR U9157 ( .A(n9798), .B(n9788), .Z(n9790) );
  XOR U9158 ( .A(n9799), .B(n9800), .Z(n9788) );
  AND U9159 ( .A(n489), .B(n9801), .Z(n9800) );
  XOR U9160 ( .A(p_input[356]), .B(n9799), .Z(n9801) );
  XOR U9161 ( .A(n9802), .B(n9803), .Z(n9799) );
  AND U9162 ( .A(n493), .B(n9804), .Z(n9803) );
  IV U9163 ( .A(n9796), .Z(n9798) );
  XOR U9164 ( .A(n9805), .B(n9806), .Z(n9796) );
  AND U9165 ( .A(n497), .B(n9807), .Z(n9806) );
  XOR U9166 ( .A(n9808), .B(n9809), .Z(n9794) );
  AND U9167 ( .A(n501), .B(n9807), .Z(n9809) );
  XNOR U9168 ( .A(n9808), .B(n9805), .Z(n9807) );
  XOR U9169 ( .A(n9810), .B(n9811), .Z(n9805) );
  AND U9170 ( .A(n504), .B(n9804), .Z(n9811) );
  XNOR U9171 ( .A(n9812), .B(n9802), .Z(n9804) );
  XOR U9172 ( .A(n9813), .B(n9814), .Z(n9802) );
  AND U9173 ( .A(n508), .B(n9815), .Z(n9814) );
  XOR U9174 ( .A(p_input[372]), .B(n9813), .Z(n9815) );
  XOR U9175 ( .A(n9816), .B(n9817), .Z(n9813) );
  AND U9176 ( .A(n512), .B(n9818), .Z(n9817) );
  IV U9177 ( .A(n9810), .Z(n9812) );
  XOR U9178 ( .A(n9819), .B(n9820), .Z(n9810) );
  AND U9179 ( .A(n516), .B(n9821), .Z(n9820) );
  XOR U9180 ( .A(n9822), .B(n9823), .Z(n9808) );
  AND U9181 ( .A(n520), .B(n9821), .Z(n9823) );
  XNOR U9182 ( .A(n9822), .B(n9819), .Z(n9821) );
  XOR U9183 ( .A(n9824), .B(n9825), .Z(n9819) );
  AND U9184 ( .A(n523), .B(n9818), .Z(n9825) );
  XNOR U9185 ( .A(n9826), .B(n9816), .Z(n9818) );
  XOR U9186 ( .A(n9827), .B(n9828), .Z(n9816) );
  AND U9187 ( .A(n527), .B(n9829), .Z(n9828) );
  XOR U9188 ( .A(p_input[388]), .B(n9827), .Z(n9829) );
  XOR U9189 ( .A(n9830), .B(n9831), .Z(n9827) );
  AND U9190 ( .A(n531), .B(n9832), .Z(n9831) );
  IV U9191 ( .A(n9824), .Z(n9826) );
  XOR U9192 ( .A(n9833), .B(n9834), .Z(n9824) );
  AND U9193 ( .A(n535), .B(n9835), .Z(n9834) );
  XOR U9194 ( .A(n9836), .B(n9837), .Z(n9822) );
  AND U9195 ( .A(n539), .B(n9835), .Z(n9837) );
  XNOR U9196 ( .A(n9836), .B(n9833), .Z(n9835) );
  XOR U9197 ( .A(n9838), .B(n9839), .Z(n9833) );
  AND U9198 ( .A(n542), .B(n9832), .Z(n9839) );
  XNOR U9199 ( .A(n9840), .B(n9830), .Z(n9832) );
  XOR U9200 ( .A(n9841), .B(n9842), .Z(n9830) );
  AND U9201 ( .A(n546), .B(n9843), .Z(n9842) );
  XOR U9202 ( .A(p_input[404]), .B(n9841), .Z(n9843) );
  XOR U9203 ( .A(n9844), .B(n9845), .Z(n9841) );
  AND U9204 ( .A(n550), .B(n9846), .Z(n9845) );
  IV U9205 ( .A(n9838), .Z(n9840) );
  XOR U9206 ( .A(n9847), .B(n9848), .Z(n9838) );
  AND U9207 ( .A(n554), .B(n9849), .Z(n9848) );
  XOR U9208 ( .A(n9850), .B(n9851), .Z(n9836) );
  AND U9209 ( .A(n558), .B(n9849), .Z(n9851) );
  XNOR U9210 ( .A(n9850), .B(n9847), .Z(n9849) );
  XOR U9211 ( .A(n9852), .B(n9853), .Z(n9847) );
  AND U9212 ( .A(n561), .B(n9846), .Z(n9853) );
  XNOR U9213 ( .A(n9854), .B(n9844), .Z(n9846) );
  XOR U9214 ( .A(n9855), .B(n9856), .Z(n9844) );
  AND U9215 ( .A(n565), .B(n9857), .Z(n9856) );
  XOR U9216 ( .A(p_input[420]), .B(n9855), .Z(n9857) );
  XOR U9217 ( .A(n9858), .B(n9859), .Z(n9855) );
  AND U9218 ( .A(n569), .B(n9860), .Z(n9859) );
  IV U9219 ( .A(n9852), .Z(n9854) );
  XOR U9220 ( .A(n9861), .B(n9862), .Z(n9852) );
  AND U9221 ( .A(n573), .B(n9863), .Z(n9862) );
  XOR U9222 ( .A(n9864), .B(n9865), .Z(n9850) );
  AND U9223 ( .A(n577), .B(n9863), .Z(n9865) );
  XNOR U9224 ( .A(n9864), .B(n9861), .Z(n9863) );
  XOR U9225 ( .A(n9866), .B(n9867), .Z(n9861) );
  AND U9226 ( .A(n580), .B(n9860), .Z(n9867) );
  XNOR U9227 ( .A(n9868), .B(n9858), .Z(n9860) );
  XOR U9228 ( .A(n9869), .B(n9870), .Z(n9858) );
  AND U9229 ( .A(n584), .B(n9871), .Z(n9870) );
  XOR U9230 ( .A(p_input[436]), .B(n9869), .Z(n9871) );
  XOR U9231 ( .A(n9872), .B(n9873), .Z(n9869) );
  AND U9232 ( .A(n588), .B(n9874), .Z(n9873) );
  IV U9233 ( .A(n9866), .Z(n9868) );
  XOR U9234 ( .A(n9875), .B(n9876), .Z(n9866) );
  AND U9235 ( .A(n592), .B(n9877), .Z(n9876) );
  XOR U9236 ( .A(n9878), .B(n9879), .Z(n9864) );
  AND U9237 ( .A(n596), .B(n9877), .Z(n9879) );
  XNOR U9238 ( .A(n9878), .B(n9875), .Z(n9877) );
  XOR U9239 ( .A(n9880), .B(n9881), .Z(n9875) );
  AND U9240 ( .A(n599), .B(n9874), .Z(n9881) );
  XNOR U9241 ( .A(n9882), .B(n9872), .Z(n9874) );
  XOR U9242 ( .A(n9883), .B(n9884), .Z(n9872) );
  AND U9243 ( .A(n603), .B(n9885), .Z(n9884) );
  XOR U9244 ( .A(p_input[452]), .B(n9883), .Z(n9885) );
  XOR U9245 ( .A(n9886), .B(n9887), .Z(n9883) );
  AND U9246 ( .A(n607), .B(n9888), .Z(n9887) );
  IV U9247 ( .A(n9880), .Z(n9882) );
  XOR U9248 ( .A(n9889), .B(n9890), .Z(n9880) );
  AND U9249 ( .A(n611), .B(n9891), .Z(n9890) );
  XOR U9250 ( .A(n9892), .B(n9893), .Z(n9878) );
  AND U9251 ( .A(n615), .B(n9891), .Z(n9893) );
  XNOR U9252 ( .A(n9892), .B(n9889), .Z(n9891) );
  XOR U9253 ( .A(n9894), .B(n9895), .Z(n9889) );
  AND U9254 ( .A(n618), .B(n9888), .Z(n9895) );
  XNOR U9255 ( .A(n9896), .B(n9886), .Z(n9888) );
  XOR U9256 ( .A(n9897), .B(n9898), .Z(n9886) );
  AND U9257 ( .A(n622), .B(n9899), .Z(n9898) );
  XOR U9258 ( .A(p_input[468]), .B(n9897), .Z(n9899) );
  XOR U9259 ( .A(n9900), .B(n9901), .Z(n9897) );
  AND U9260 ( .A(n626), .B(n9902), .Z(n9901) );
  IV U9261 ( .A(n9894), .Z(n9896) );
  XOR U9262 ( .A(n9903), .B(n9904), .Z(n9894) );
  AND U9263 ( .A(n630), .B(n9905), .Z(n9904) );
  XOR U9264 ( .A(n9906), .B(n9907), .Z(n9892) );
  AND U9265 ( .A(n634), .B(n9905), .Z(n9907) );
  XNOR U9266 ( .A(n9906), .B(n9903), .Z(n9905) );
  XOR U9267 ( .A(n9908), .B(n9909), .Z(n9903) );
  AND U9268 ( .A(n637), .B(n9902), .Z(n9909) );
  XNOR U9269 ( .A(n9910), .B(n9900), .Z(n9902) );
  XOR U9270 ( .A(n9911), .B(n9912), .Z(n9900) );
  AND U9271 ( .A(n641), .B(n9913), .Z(n9912) );
  XOR U9272 ( .A(p_input[484]), .B(n9911), .Z(n9913) );
  XOR U9273 ( .A(n9914), .B(n9915), .Z(n9911) );
  AND U9274 ( .A(n645), .B(n9916), .Z(n9915) );
  IV U9275 ( .A(n9908), .Z(n9910) );
  XOR U9276 ( .A(n9917), .B(n9918), .Z(n9908) );
  AND U9277 ( .A(n649), .B(n9919), .Z(n9918) );
  XOR U9278 ( .A(n9920), .B(n9921), .Z(n9906) );
  AND U9279 ( .A(n653), .B(n9919), .Z(n9921) );
  XNOR U9280 ( .A(n9920), .B(n9917), .Z(n9919) );
  XOR U9281 ( .A(n9922), .B(n9923), .Z(n9917) );
  AND U9282 ( .A(n656), .B(n9916), .Z(n9923) );
  XNOR U9283 ( .A(n9924), .B(n9914), .Z(n9916) );
  XOR U9284 ( .A(n9925), .B(n9926), .Z(n9914) );
  AND U9285 ( .A(n660), .B(n9927), .Z(n9926) );
  XOR U9286 ( .A(p_input[500]), .B(n9925), .Z(n9927) );
  XOR U9287 ( .A(n9928), .B(n9929), .Z(n9925) );
  AND U9288 ( .A(n664), .B(n9930), .Z(n9929) );
  IV U9289 ( .A(n9922), .Z(n9924) );
  XOR U9290 ( .A(n9931), .B(n9932), .Z(n9922) );
  AND U9291 ( .A(n668), .B(n9933), .Z(n9932) );
  XOR U9292 ( .A(n9934), .B(n9935), .Z(n9920) );
  AND U9293 ( .A(n672), .B(n9933), .Z(n9935) );
  XNOR U9294 ( .A(n9934), .B(n9931), .Z(n9933) );
  XOR U9295 ( .A(n9936), .B(n9937), .Z(n9931) );
  AND U9296 ( .A(n675), .B(n9930), .Z(n9937) );
  XNOR U9297 ( .A(n9938), .B(n9928), .Z(n9930) );
  XOR U9298 ( .A(n9939), .B(n9940), .Z(n9928) );
  AND U9299 ( .A(n679), .B(n9941), .Z(n9940) );
  XOR U9300 ( .A(p_input[516]), .B(n9939), .Z(n9941) );
  XOR U9301 ( .A(n9942), .B(n9943), .Z(n9939) );
  AND U9302 ( .A(n683), .B(n9944), .Z(n9943) );
  IV U9303 ( .A(n9936), .Z(n9938) );
  XOR U9304 ( .A(n9945), .B(n9946), .Z(n9936) );
  AND U9305 ( .A(n687), .B(n9947), .Z(n9946) );
  XOR U9306 ( .A(n9948), .B(n9949), .Z(n9934) );
  AND U9307 ( .A(n691), .B(n9947), .Z(n9949) );
  XNOR U9308 ( .A(n9948), .B(n9945), .Z(n9947) );
  XOR U9309 ( .A(n9950), .B(n9951), .Z(n9945) );
  AND U9310 ( .A(n694), .B(n9944), .Z(n9951) );
  XNOR U9311 ( .A(n9952), .B(n9942), .Z(n9944) );
  XOR U9312 ( .A(n9953), .B(n9954), .Z(n9942) );
  AND U9313 ( .A(n698), .B(n9955), .Z(n9954) );
  XOR U9314 ( .A(p_input[532]), .B(n9953), .Z(n9955) );
  XOR U9315 ( .A(n9956), .B(n9957), .Z(n9953) );
  AND U9316 ( .A(n702), .B(n9958), .Z(n9957) );
  IV U9317 ( .A(n9950), .Z(n9952) );
  XOR U9318 ( .A(n9959), .B(n9960), .Z(n9950) );
  AND U9319 ( .A(n706), .B(n9961), .Z(n9960) );
  XOR U9320 ( .A(n9962), .B(n9963), .Z(n9948) );
  AND U9321 ( .A(n710), .B(n9961), .Z(n9963) );
  XNOR U9322 ( .A(n9962), .B(n9959), .Z(n9961) );
  XOR U9323 ( .A(n9964), .B(n9965), .Z(n9959) );
  AND U9324 ( .A(n713), .B(n9958), .Z(n9965) );
  XNOR U9325 ( .A(n9966), .B(n9956), .Z(n9958) );
  XOR U9326 ( .A(n9967), .B(n9968), .Z(n9956) );
  AND U9327 ( .A(n717), .B(n9969), .Z(n9968) );
  XOR U9328 ( .A(p_input[548]), .B(n9967), .Z(n9969) );
  XOR U9329 ( .A(n9970), .B(n9971), .Z(n9967) );
  AND U9330 ( .A(n721), .B(n9972), .Z(n9971) );
  IV U9331 ( .A(n9964), .Z(n9966) );
  XOR U9332 ( .A(n9973), .B(n9974), .Z(n9964) );
  AND U9333 ( .A(n725), .B(n9975), .Z(n9974) );
  XOR U9334 ( .A(n9976), .B(n9977), .Z(n9962) );
  AND U9335 ( .A(n729), .B(n9975), .Z(n9977) );
  XNOR U9336 ( .A(n9976), .B(n9973), .Z(n9975) );
  XOR U9337 ( .A(n9978), .B(n9979), .Z(n9973) );
  AND U9338 ( .A(n732), .B(n9972), .Z(n9979) );
  XNOR U9339 ( .A(n9980), .B(n9970), .Z(n9972) );
  XOR U9340 ( .A(n9981), .B(n9982), .Z(n9970) );
  AND U9341 ( .A(n736), .B(n9983), .Z(n9982) );
  XOR U9342 ( .A(p_input[564]), .B(n9981), .Z(n9983) );
  XOR U9343 ( .A(n9984), .B(n9985), .Z(n9981) );
  AND U9344 ( .A(n740), .B(n9986), .Z(n9985) );
  IV U9345 ( .A(n9978), .Z(n9980) );
  XOR U9346 ( .A(n9987), .B(n9988), .Z(n9978) );
  AND U9347 ( .A(n744), .B(n9989), .Z(n9988) );
  XOR U9348 ( .A(n9990), .B(n9991), .Z(n9976) );
  AND U9349 ( .A(n748), .B(n9989), .Z(n9991) );
  XNOR U9350 ( .A(n9990), .B(n9987), .Z(n9989) );
  XOR U9351 ( .A(n9992), .B(n9993), .Z(n9987) );
  AND U9352 ( .A(n751), .B(n9986), .Z(n9993) );
  XNOR U9353 ( .A(n9994), .B(n9984), .Z(n9986) );
  XOR U9354 ( .A(n9995), .B(n9996), .Z(n9984) );
  AND U9355 ( .A(n755), .B(n9997), .Z(n9996) );
  XOR U9356 ( .A(p_input[580]), .B(n9995), .Z(n9997) );
  XOR U9357 ( .A(n9998), .B(n9999), .Z(n9995) );
  AND U9358 ( .A(n759), .B(n10000), .Z(n9999) );
  IV U9359 ( .A(n9992), .Z(n9994) );
  XOR U9360 ( .A(n10001), .B(n10002), .Z(n9992) );
  AND U9361 ( .A(n763), .B(n10003), .Z(n10002) );
  XOR U9362 ( .A(n10004), .B(n10005), .Z(n9990) );
  AND U9363 ( .A(n767), .B(n10003), .Z(n10005) );
  XNOR U9364 ( .A(n10004), .B(n10001), .Z(n10003) );
  XOR U9365 ( .A(n10006), .B(n10007), .Z(n10001) );
  AND U9366 ( .A(n770), .B(n10000), .Z(n10007) );
  XNOR U9367 ( .A(n10008), .B(n9998), .Z(n10000) );
  XOR U9368 ( .A(n10009), .B(n10010), .Z(n9998) );
  AND U9369 ( .A(n774), .B(n10011), .Z(n10010) );
  XOR U9370 ( .A(p_input[596]), .B(n10009), .Z(n10011) );
  XOR U9371 ( .A(n10012), .B(n10013), .Z(n10009) );
  AND U9372 ( .A(n778), .B(n10014), .Z(n10013) );
  IV U9373 ( .A(n10006), .Z(n10008) );
  XOR U9374 ( .A(n10015), .B(n10016), .Z(n10006) );
  AND U9375 ( .A(n782), .B(n10017), .Z(n10016) );
  XOR U9376 ( .A(n10018), .B(n10019), .Z(n10004) );
  AND U9377 ( .A(n786), .B(n10017), .Z(n10019) );
  XNOR U9378 ( .A(n10018), .B(n10015), .Z(n10017) );
  XOR U9379 ( .A(n10020), .B(n10021), .Z(n10015) );
  AND U9380 ( .A(n789), .B(n10014), .Z(n10021) );
  XNOR U9381 ( .A(n10022), .B(n10012), .Z(n10014) );
  XOR U9382 ( .A(n10023), .B(n10024), .Z(n10012) );
  AND U9383 ( .A(n793), .B(n10025), .Z(n10024) );
  XOR U9384 ( .A(p_input[612]), .B(n10023), .Z(n10025) );
  XOR U9385 ( .A(n10026), .B(n10027), .Z(n10023) );
  AND U9386 ( .A(n797), .B(n10028), .Z(n10027) );
  IV U9387 ( .A(n10020), .Z(n10022) );
  XOR U9388 ( .A(n10029), .B(n10030), .Z(n10020) );
  AND U9389 ( .A(n801), .B(n10031), .Z(n10030) );
  XOR U9390 ( .A(n10032), .B(n10033), .Z(n10018) );
  AND U9391 ( .A(n805), .B(n10031), .Z(n10033) );
  XNOR U9392 ( .A(n10032), .B(n10029), .Z(n10031) );
  XOR U9393 ( .A(n10034), .B(n10035), .Z(n10029) );
  AND U9394 ( .A(n808), .B(n10028), .Z(n10035) );
  XNOR U9395 ( .A(n10036), .B(n10026), .Z(n10028) );
  XOR U9396 ( .A(n10037), .B(n10038), .Z(n10026) );
  AND U9397 ( .A(n812), .B(n10039), .Z(n10038) );
  XOR U9398 ( .A(p_input[628]), .B(n10037), .Z(n10039) );
  XOR U9399 ( .A(n10040), .B(n10041), .Z(n10037) );
  AND U9400 ( .A(n816), .B(n10042), .Z(n10041) );
  IV U9401 ( .A(n10034), .Z(n10036) );
  XOR U9402 ( .A(n10043), .B(n10044), .Z(n10034) );
  AND U9403 ( .A(n820), .B(n10045), .Z(n10044) );
  XOR U9404 ( .A(n10046), .B(n10047), .Z(n10032) );
  AND U9405 ( .A(n824), .B(n10045), .Z(n10047) );
  XNOR U9406 ( .A(n10046), .B(n10043), .Z(n10045) );
  XOR U9407 ( .A(n10048), .B(n10049), .Z(n10043) );
  AND U9408 ( .A(n827), .B(n10042), .Z(n10049) );
  XNOR U9409 ( .A(n10050), .B(n10040), .Z(n10042) );
  XOR U9410 ( .A(n10051), .B(n10052), .Z(n10040) );
  AND U9411 ( .A(n831), .B(n10053), .Z(n10052) );
  XOR U9412 ( .A(p_input[644]), .B(n10051), .Z(n10053) );
  XOR U9413 ( .A(n10054), .B(n10055), .Z(n10051) );
  AND U9414 ( .A(n835), .B(n10056), .Z(n10055) );
  IV U9415 ( .A(n10048), .Z(n10050) );
  XOR U9416 ( .A(n10057), .B(n10058), .Z(n10048) );
  AND U9417 ( .A(n839), .B(n10059), .Z(n10058) );
  XOR U9418 ( .A(n10060), .B(n10061), .Z(n10046) );
  AND U9419 ( .A(n843), .B(n10059), .Z(n10061) );
  XNOR U9420 ( .A(n10060), .B(n10057), .Z(n10059) );
  XOR U9421 ( .A(n10062), .B(n10063), .Z(n10057) );
  AND U9422 ( .A(n846), .B(n10056), .Z(n10063) );
  XNOR U9423 ( .A(n10064), .B(n10054), .Z(n10056) );
  XOR U9424 ( .A(n10065), .B(n10066), .Z(n10054) );
  AND U9425 ( .A(n850), .B(n10067), .Z(n10066) );
  XOR U9426 ( .A(p_input[660]), .B(n10065), .Z(n10067) );
  XOR U9427 ( .A(n10068), .B(n10069), .Z(n10065) );
  AND U9428 ( .A(n854), .B(n10070), .Z(n10069) );
  IV U9429 ( .A(n10062), .Z(n10064) );
  XOR U9430 ( .A(n10071), .B(n10072), .Z(n10062) );
  AND U9431 ( .A(n858), .B(n10073), .Z(n10072) );
  XOR U9432 ( .A(n10074), .B(n10075), .Z(n10060) );
  AND U9433 ( .A(n862), .B(n10073), .Z(n10075) );
  XNOR U9434 ( .A(n10074), .B(n10071), .Z(n10073) );
  XOR U9435 ( .A(n10076), .B(n10077), .Z(n10071) );
  AND U9436 ( .A(n865), .B(n10070), .Z(n10077) );
  XNOR U9437 ( .A(n10078), .B(n10068), .Z(n10070) );
  XOR U9438 ( .A(n10079), .B(n10080), .Z(n10068) );
  AND U9439 ( .A(n869), .B(n10081), .Z(n10080) );
  XOR U9440 ( .A(p_input[676]), .B(n10079), .Z(n10081) );
  XOR U9441 ( .A(n10082), .B(n10083), .Z(n10079) );
  AND U9442 ( .A(n873), .B(n10084), .Z(n10083) );
  IV U9443 ( .A(n10076), .Z(n10078) );
  XOR U9444 ( .A(n10085), .B(n10086), .Z(n10076) );
  AND U9445 ( .A(n877), .B(n10087), .Z(n10086) );
  XOR U9446 ( .A(n10088), .B(n10089), .Z(n10074) );
  AND U9447 ( .A(n881), .B(n10087), .Z(n10089) );
  XNOR U9448 ( .A(n10088), .B(n10085), .Z(n10087) );
  XOR U9449 ( .A(n10090), .B(n10091), .Z(n10085) );
  AND U9450 ( .A(n884), .B(n10084), .Z(n10091) );
  XNOR U9451 ( .A(n10092), .B(n10082), .Z(n10084) );
  XOR U9452 ( .A(n10093), .B(n10094), .Z(n10082) );
  AND U9453 ( .A(n888), .B(n10095), .Z(n10094) );
  XOR U9454 ( .A(p_input[692]), .B(n10093), .Z(n10095) );
  XOR U9455 ( .A(n10096), .B(n10097), .Z(n10093) );
  AND U9456 ( .A(n892), .B(n10098), .Z(n10097) );
  IV U9457 ( .A(n10090), .Z(n10092) );
  XOR U9458 ( .A(n10099), .B(n10100), .Z(n10090) );
  AND U9459 ( .A(n896), .B(n10101), .Z(n10100) );
  XOR U9460 ( .A(n10102), .B(n10103), .Z(n10088) );
  AND U9461 ( .A(n900), .B(n10101), .Z(n10103) );
  XNOR U9462 ( .A(n10102), .B(n10099), .Z(n10101) );
  XOR U9463 ( .A(n10104), .B(n10105), .Z(n10099) );
  AND U9464 ( .A(n903), .B(n10098), .Z(n10105) );
  XNOR U9465 ( .A(n10106), .B(n10096), .Z(n10098) );
  XOR U9466 ( .A(n10107), .B(n10108), .Z(n10096) );
  AND U9467 ( .A(n907), .B(n10109), .Z(n10108) );
  XOR U9468 ( .A(p_input[708]), .B(n10107), .Z(n10109) );
  XOR U9469 ( .A(n10110), .B(n10111), .Z(n10107) );
  AND U9470 ( .A(n911), .B(n10112), .Z(n10111) );
  IV U9471 ( .A(n10104), .Z(n10106) );
  XOR U9472 ( .A(n10113), .B(n10114), .Z(n10104) );
  AND U9473 ( .A(n915), .B(n10115), .Z(n10114) );
  XOR U9474 ( .A(n10116), .B(n10117), .Z(n10102) );
  AND U9475 ( .A(n919), .B(n10115), .Z(n10117) );
  XNOR U9476 ( .A(n10116), .B(n10113), .Z(n10115) );
  XOR U9477 ( .A(n10118), .B(n10119), .Z(n10113) );
  AND U9478 ( .A(n922), .B(n10112), .Z(n10119) );
  XNOR U9479 ( .A(n10120), .B(n10110), .Z(n10112) );
  XOR U9480 ( .A(n10121), .B(n10122), .Z(n10110) );
  AND U9481 ( .A(n926), .B(n10123), .Z(n10122) );
  XOR U9482 ( .A(p_input[724]), .B(n10121), .Z(n10123) );
  XOR U9483 ( .A(n10124), .B(n10125), .Z(n10121) );
  AND U9484 ( .A(n930), .B(n10126), .Z(n10125) );
  IV U9485 ( .A(n10118), .Z(n10120) );
  XOR U9486 ( .A(n10127), .B(n10128), .Z(n10118) );
  AND U9487 ( .A(n934), .B(n10129), .Z(n10128) );
  XOR U9488 ( .A(n10130), .B(n10131), .Z(n10116) );
  AND U9489 ( .A(n938), .B(n10129), .Z(n10131) );
  XNOR U9490 ( .A(n10130), .B(n10127), .Z(n10129) );
  XOR U9491 ( .A(n10132), .B(n10133), .Z(n10127) );
  AND U9492 ( .A(n941), .B(n10126), .Z(n10133) );
  XNOR U9493 ( .A(n10134), .B(n10124), .Z(n10126) );
  XOR U9494 ( .A(n10135), .B(n10136), .Z(n10124) );
  AND U9495 ( .A(n945), .B(n10137), .Z(n10136) );
  XOR U9496 ( .A(p_input[740]), .B(n10135), .Z(n10137) );
  XOR U9497 ( .A(n10138), .B(n10139), .Z(n10135) );
  AND U9498 ( .A(n949), .B(n10140), .Z(n10139) );
  IV U9499 ( .A(n10132), .Z(n10134) );
  XOR U9500 ( .A(n10141), .B(n10142), .Z(n10132) );
  AND U9501 ( .A(n953), .B(n10143), .Z(n10142) );
  XOR U9502 ( .A(n10144), .B(n10145), .Z(n10130) );
  AND U9503 ( .A(n957), .B(n10143), .Z(n10145) );
  XNOR U9504 ( .A(n10144), .B(n10141), .Z(n10143) );
  XOR U9505 ( .A(n10146), .B(n10147), .Z(n10141) );
  AND U9506 ( .A(n960), .B(n10140), .Z(n10147) );
  XNOR U9507 ( .A(n10148), .B(n10138), .Z(n10140) );
  XOR U9508 ( .A(n10149), .B(n10150), .Z(n10138) );
  AND U9509 ( .A(n964), .B(n10151), .Z(n10150) );
  XOR U9510 ( .A(p_input[756]), .B(n10149), .Z(n10151) );
  XOR U9511 ( .A(n10152), .B(n10153), .Z(n10149) );
  AND U9512 ( .A(n968), .B(n10154), .Z(n10153) );
  IV U9513 ( .A(n10146), .Z(n10148) );
  XOR U9514 ( .A(n10155), .B(n10156), .Z(n10146) );
  AND U9515 ( .A(n972), .B(n10157), .Z(n10156) );
  XOR U9516 ( .A(n10158), .B(n10159), .Z(n10144) );
  AND U9517 ( .A(n976), .B(n10157), .Z(n10159) );
  XNOR U9518 ( .A(n10158), .B(n10155), .Z(n10157) );
  XOR U9519 ( .A(n10160), .B(n10161), .Z(n10155) );
  AND U9520 ( .A(n979), .B(n10154), .Z(n10161) );
  XNOR U9521 ( .A(n10162), .B(n10152), .Z(n10154) );
  XOR U9522 ( .A(n10163), .B(n10164), .Z(n10152) );
  AND U9523 ( .A(n983), .B(n10165), .Z(n10164) );
  XOR U9524 ( .A(p_input[772]), .B(n10163), .Z(n10165) );
  XOR U9525 ( .A(n10166), .B(n10167), .Z(n10163) );
  AND U9526 ( .A(n987), .B(n10168), .Z(n10167) );
  IV U9527 ( .A(n10160), .Z(n10162) );
  XOR U9528 ( .A(n10169), .B(n10170), .Z(n10160) );
  AND U9529 ( .A(n991), .B(n10171), .Z(n10170) );
  XOR U9530 ( .A(n10172), .B(n10173), .Z(n10158) );
  AND U9531 ( .A(n995), .B(n10171), .Z(n10173) );
  XNOR U9532 ( .A(n10172), .B(n10169), .Z(n10171) );
  XOR U9533 ( .A(n10174), .B(n10175), .Z(n10169) );
  AND U9534 ( .A(n998), .B(n10168), .Z(n10175) );
  XNOR U9535 ( .A(n10176), .B(n10166), .Z(n10168) );
  XOR U9536 ( .A(n10177), .B(n10178), .Z(n10166) );
  AND U9537 ( .A(n1002), .B(n10179), .Z(n10178) );
  XOR U9538 ( .A(p_input[788]), .B(n10177), .Z(n10179) );
  XOR U9539 ( .A(n10180), .B(n10181), .Z(n10177) );
  AND U9540 ( .A(n1006), .B(n10182), .Z(n10181) );
  IV U9541 ( .A(n10174), .Z(n10176) );
  XOR U9542 ( .A(n10183), .B(n10184), .Z(n10174) );
  AND U9543 ( .A(n1010), .B(n10185), .Z(n10184) );
  XOR U9544 ( .A(n10186), .B(n10187), .Z(n10172) );
  AND U9545 ( .A(n1014), .B(n10185), .Z(n10187) );
  XNOR U9546 ( .A(n10186), .B(n10183), .Z(n10185) );
  XOR U9547 ( .A(n10188), .B(n10189), .Z(n10183) );
  AND U9548 ( .A(n1017), .B(n10182), .Z(n10189) );
  XNOR U9549 ( .A(n10190), .B(n10180), .Z(n10182) );
  XOR U9550 ( .A(n10191), .B(n10192), .Z(n10180) );
  AND U9551 ( .A(n1021), .B(n10193), .Z(n10192) );
  XOR U9552 ( .A(p_input[804]), .B(n10191), .Z(n10193) );
  XOR U9553 ( .A(n10194), .B(n10195), .Z(n10191) );
  AND U9554 ( .A(n1025), .B(n10196), .Z(n10195) );
  IV U9555 ( .A(n10188), .Z(n10190) );
  XOR U9556 ( .A(n10197), .B(n10198), .Z(n10188) );
  AND U9557 ( .A(n1029), .B(n10199), .Z(n10198) );
  XOR U9558 ( .A(n10200), .B(n10201), .Z(n10186) );
  AND U9559 ( .A(n1033), .B(n10199), .Z(n10201) );
  XNOR U9560 ( .A(n10200), .B(n10197), .Z(n10199) );
  XOR U9561 ( .A(n10202), .B(n10203), .Z(n10197) );
  AND U9562 ( .A(n1036), .B(n10196), .Z(n10203) );
  XNOR U9563 ( .A(n10204), .B(n10194), .Z(n10196) );
  XOR U9564 ( .A(n10205), .B(n10206), .Z(n10194) );
  AND U9565 ( .A(n1040), .B(n10207), .Z(n10206) );
  XOR U9566 ( .A(p_input[820]), .B(n10205), .Z(n10207) );
  XOR U9567 ( .A(n10208), .B(n10209), .Z(n10205) );
  AND U9568 ( .A(n1044), .B(n10210), .Z(n10209) );
  IV U9569 ( .A(n10202), .Z(n10204) );
  XOR U9570 ( .A(n10211), .B(n10212), .Z(n10202) );
  AND U9571 ( .A(n1048), .B(n10213), .Z(n10212) );
  XOR U9572 ( .A(n10214), .B(n10215), .Z(n10200) );
  AND U9573 ( .A(n1052), .B(n10213), .Z(n10215) );
  XNOR U9574 ( .A(n10214), .B(n10211), .Z(n10213) );
  XOR U9575 ( .A(n10216), .B(n10217), .Z(n10211) );
  AND U9576 ( .A(n1055), .B(n10210), .Z(n10217) );
  XNOR U9577 ( .A(n10218), .B(n10208), .Z(n10210) );
  XOR U9578 ( .A(n10219), .B(n10220), .Z(n10208) );
  AND U9579 ( .A(n1059), .B(n10221), .Z(n10220) );
  XOR U9580 ( .A(p_input[836]), .B(n10219), .Z(n10221) );
  XOR U9581 ( .A(n10222), .B(n10223), .Z(n10219) );
  AND U9582 ( .A(n1063), .B(n10224), .Z(n10223) );
  IV U9583 ( .A(n10216), .Z(n10218) );
  XOR U9584 ( .A(n10225), .B(n10226), .Z(n10216) );
  AND U9585 ( .A(n1067), .B(n10227), .Z(n10226) );
  XOR U9586 ( .A(n10228), .B(n10229), .Z(n10214) );
  AND U9587 ( .A(n1071), .B(n10227), .Z(n10229) );
  XNOR U9588 ( .A(n10228), .B(n10225), .Z(n10227) );
  XOR U9589 ( .A(n10230), .B(n10231), .Z(n10225) );
  AND U9590 ( .A(n1074), .B(n10224), .Z(n10231) );
  XNOR U9591 ( .A(n10232), .B(n10222), .Z(n10224) );
  XOR U9592 ( .A(n10233), .B(n10234), .Z(n10222) );
  AND U9593 ( .A(n1078), .B(n10235), .Z(n10234) );
  XOR U9594 ( .A(p_input[852]), .B(n10233), .Z(n10235) );
  XOR U9595 ( .A(n10236), .B(n10237), .Z(n10233) );
  AND U9596 ( .A(n1082), .B(n10238), .Z(n10237) );
  IV U9597 ( .A(n10230), .Z(n10232) );
  XOR U9598 ( .A(n10239), .B(n10240), .Z(n10230) );
  AND U9599 ( .A(n1086), .B(n10241), .Z(n10240) );
  XOR U9600 ( .A(n10242), .B(n10243), .Z(n10228) );
  AND U9601 ( .A(n1090), .B(n10241), .Z(n10243) );
  XNOR U9602 ( .A(n10242), .B(n10239), .Z(n10241) );
  XOR U9603 ( .A(n10244), .B(n10245), .Z(n10239) );
  AND U9604 ( .A(n1093), .B(n10238), .Z(n10245) );
  XNOR U9605 ( .A(n10246), .B(n10236), .Z(n10238) );
  XOR U9606 ( .A(n10247), .B(n10248), .Z(n10236) );
  AND U9607 ( .A(n1097), .B(n10249), .Z(n10248) );
  XOR U9608 ( .A(p_input[868]), .B(n10247), .Z(n10249) );
  XOR U9609 ( .A(n10250), .B(n10251), .Z(n10247) );
  AND U9610 ( .A(n1101), .B(n10252), .Z(n10251) );
  IV U9611 ( .A(n10244), .Z(n10246) );
  XOR U9612 ( .A(n10253), .B(n10254), .Z(n10244) );
  AND U9613 ( .A(n1105), .B(n10255), .Z(n10254) );
  XOR U9614 ( .A(n10256), .B(n10257), .Z(n10242) );
  AND U9615 ( .A(n1109), .B(n10255), .Z(n10257) );
  XNOR U9616 ( .A(n10256), .B(n10253), .Z(n10255) );
  XOR U9617 ( .A(n10258), .B(n10259), .Z(n10253) );
  AND U9618 ( .A(n1112), .B(n10252), .Z(n10259) );
  XNOR U9619 ( .A(n10260), .B(n10250), .Z(n10252) );
  XOR U9620 ( .A(n10261), .B(n10262), .Z(n10250) );
  AND U9621 ( .A(n1116), .B(n10263), .Z(n10262) );
  XOR U9622 ( .A(p_input[884]), .B(n10261), .Z(n10263) );
  XOR U9623 ( .A(n10264), .B(n10265), .Z(n10261) );
  AND U9624 ( .A(n1120), .B(n10266), .Z(n10265) );
  IV U9625 ( .A(n10258), .Z(n10260) );
  XOR U9626 ( .A(n10267), .B(n10268), .Z(n10258) );
  AND U9627 ( .A(n1124), .B(n10269), .Z(n10268) );
  XOR U9628 ( .A(n10270), .B(n10271), .Z(n10256) );
  AND U9629 ( .A(n1128), .B(n10269), .Z(n10271) );
  XNOR U9630 ( .A(n10270), .B(n10267), .Z(n10269) );
  XOR U9631 ( .A(n10272), .B(n10273), .Z(n10267) );
  AND U9632 ( .A(n1131), .B(n10266), .Z(n10273) );
  XNOR U9633 ( .A(n10274), .B(n10264), .Z(n10266) );
  XOR U9634 ( .A(n10275), .B(n10276), .Z(n10264) );
  AND U9635 ( .A(n1135), .B(n10277), .Z(n10276) );
  XOR U9636 ( .A(p_input[900]), .B(n10275), .Z(n10277) );
  XOR U9637 ( .A(n10278), .B(n10279), .Z(n10275) );
  AND U9638 ( .A(n1139), .B(n10280), .Z(n10279) );
  IV U9639 ( .A(n10272), .Z(n10274) );
  XOR U9640 ( .A(n10281), .B(n10282), .Z(n10272) );
  AND U9641 ( .A(n1143), .B(n10283), .Z(n10282) );
  XOR U9642 ( .A(n10284), .B(n10285), .Z(n10270) );
  AND U9643 ( .A(n1147), .B(n10283), .Z(n10285) );
  XNOR U9644 ( .A(n10284), .B(n10281), .Z(n10283) );
  XOR U9645 ( .A(n10286), .B(n10287), .Z(n10281) );
  AND U9646 ( .A(n1150), .B(n10280), .Z(n10287) );
  XNOR U9647 ( .A(n10288), .B(n10278), .Z(n10280) );
  XOR U9648 ( .A(n10289), .B(n10290), .Z(n10278) );
  AND U9649 ( .A(n1154), .B(n10291), .Z(n10290) );
  XOR U9650 ( .A(p_input[916]), .B(n10289), .Z(n10291) );
  XOR U9651 ( .A(n10292), .B(n10293), .Z(n10289) );
  AND U9652 ( .A(n1158), .B(n10294), .Z(n10293) );
  IV U9653 ( .A(n10286), .Z(n10288) );
  XOR U9654 ( .A(n10295), .B(n10296), .Z(n10286) );
  AND U9655 ( .A(n1162), .B(n10297), .Z(n10296) );
  XOR U9656 ( .A(n10298), .B(n10299), .Z(n10284) );
  AND U9657 ( .A(n1166), .B(n10297), .Z(n10299) );
  XNOR U9658 ( .A(n10298), .B(n10295), .Z(n10297) );
  XOR U9659 ( .A(n10300), .B(n10301), .Z(n10295) );
  AND U9660 ( .A(n1169), .B(n10294), .Z(n10301) );
  XNOR U9661 ( .A(n10302), .B(n10292), .Z(n10294) );
  XOR U9662 ( .A(n10303), .B(n10304), .Z(n10292) );
  AND U9663 ( .A(n1173), .B(n10305), .Z(n10304) );
  XOR U9664 ( .A(p_input[932]), .B(n10303), .Z(n10305) );
  XOR U9665 ( .A(n10306), .B(n10307), .Z(n10303) );
  AND U9666 ( .A(n1177), .B(n10308), .Z(n10307) );
  IV U9667 ( .A(n10300), .Z(n10302) );
  XOR U9668 ( .A(n10309), .B(n10310), .Z(n10300) );
  AND U9669 ( .A(n1181), .B(n10311), .Z(n10310) );
  XOR U9670 ( .A(n10312), .B(n10313), .Z(n10298) );
  AND U9671 ( .A(n1185), .B(n10311), .Z(n10313) );
  XNOR U9672 ( .A(n10312), .B(n10309), .Z(n10311) );
  XOR U9673 ( .A(n10314), .B(n10315), .Z(n10309) );
  AND U9674 ( .A(n1188), .B(n10308), .Z(n10315) );
  XNOR U9675 ( .A(n10316), .B(n10306), .Z(n10308) );
  XOR U9676 ( .A(n10317), .B(n10318), .Z(n10306) );
  AND U9677 ( .A(n1192), .B(n10319), .Z(n10318) );
  XOR U9678 ( .A(p_input[948]), .B(n10317), .Z(n10319) );
  XOR U9679 ( .A(n10320), .B(n10321), .Z(n10317) );
  AND U9680 ( .A(n1196), .B(n10322), .Z(n10321) );
  IV U9681 ( .A(n10314), .Z(n10316) );
  XOR U9682 ( .A(n10323), .B(n10324), .Z(n10314) );
  AND U9683 ( .A(n1200), .B(n10325), .Z(n10324) );
  XOR U9684 ( .A(n10326), .B(n10327), .Z(n10312) );
  AND U9685 ( .A(n1204), .B(n10325), .Z(n10327) );
  XNOR U9686 ( .A(n10326), .B(n10323), .Z(n10325) );
  XOR U9687 ( .A(n10328), .B(n10329), .Z(n10323) );
  AND U9688 ( .A(n1207), .B(n10322), .Z(n10329) );
  XNOR U9689 ( .A(n10330), .B(n10320), .Z(n10322) );
  XOR U9690 ( .A(n10331), .B(n10332), .Z(n10320) );
  AND U9691 ( .A(n1211), .B(n10333), .Z(n10332) );
  XOR U9692 ( .A(p_input[964]), .B(n10331), .Z(n10333) );
  XOR U9693 ( .A(n10334), .B(n10335), .Z(n10331) );
  AND U9694 ( .A(n1215), .B(n10336), .Z(n10335) );
  IV U9695 ( .A(n10328), .Z(n10330) );
  XOR U9696 ( .A(n10337), .B(n10338), .Z(n10328) );
  AND U9697 ( .A(n1219), .B(n10339), .Z(n10338) );
  XOR U9698 ( .A(n10340), .B(n10341), .Z(n10326) );
  AND U9699 ( .A(n1223), .B(n10339), .Z(n10341) );
  XNOR U9700 ( .A(n10340), .B(n10337), .Z(n10339) );
  XOR U9701 ( .A(n10342), .B(n10343), .Z(n10337) );
  AND U9702 ( .A(n1226), .B(n10336), .Z(n10343) );
  XNOR U9703 ( .A(n10344), .B(n10334), .Z(n10336) );
  XOR U9704 ( .A(n10345), .B(n10346), .Z(n10334) );
  AND U9705 ( .A(n1230), .B(n10347), .Z(n10346) );
  XOR U9706 ( .A(p_input[980]), .B(n10345), .Z(n10347) );
  XOR U9707 ( .A(n10348), .B(n10349), .Z(n10345) );
  AND U9708 ( .A(n1234), .B(n10350), .Z(n10349) );
  IV U9709 ( .A(n10342), .Z(n10344) );
  XOR U9710 ( .A(n10351), .B(n10352), .Z(n10342) );
  AND U9711 ( .A(n1238), .B(n10353), .Z(n10352) );
  XOR U9712 ( .A(n10354), .B(n10355), .Z(n10340) );
  AND U9713 ( .A(n1242), .B(n10353), .Z(n10355) );
  XNOR U9714 ( .A(n10354), .B(n10351), .Z(n10353) );
  XOR U9715 ( .A(n10356), .B(n10357), .Z(n10351) );
  AND U9716 ( .A(n1245), .B(n10350), .Z(n10357) );
  XNOR U9717 ( .A(n10358), .B(n10348), .Z(n10350) );
  XOR U9718 ( .A(n10359), .B(n10360), .Z(n10348) );
  AND U9719 ( .A(n1249), .B(n10361), .Z(n10360) );
  XOR U9720 ( .A(p_input[996]), .B(n10359), .Z(n10361) );
  XOR U9721 ( .A(n10362), .B(n10363), .Z(n10359) );
  AND U9722 ( .A(n1253), .B(n10364), .Z(n10363) );
  IV U9723 ( .A(n10356), .Z(n10358) );
  XOR U9724 ( .A(n10365), .B(n10366), .Z(n10356) );
  AND U9725 ( .A(n1257), .B(n10367), .Z(n10366) );
  XOR U9726 ( .A(n10368), .B(n10369), .Z(n10354) );
  AND U9727 ( .A(n1261), .B(n10367), .Z(n10369) );
  XNOR U9728 ( .A(n10368), .B(n10365), .Z(n10367) );
  XOR U9729 ( .A(n10370), .B(n10371), .Z(n10365) );
  AND U9730 ( .A(n1264), .B(n10364), .Z(n10371) );
  XNOR U9731 ( .A(n10372), .B(n10362), .Z(n10364) );
  XOR U9732 ( .A(n10373), .B(n10374), .Z(n10362) );
  AND U9733 ( .A(n1268), .B(n10375), .Z(n10374) );
  XOR U9734 ( .A(p_input[1012]), .B(n10373), .Z(n10375) );
  XOR U9735 ( .A(n10376), .B(n10377), .Z(n10373) );
  AND U9736 ( .A(n1272), .B(n10378), .Z(n10377) );
  IV U9737 ( .A(n10370), .Z(n10372) );
  XOR U9738 ( .A(n10379), .B(n10380), .Z(n10370) );
  AND U9739 ( .A(n1276), .B(n10381), .Z(n10380) );
  XOR U9740 ( .A(n10382), .B(n10383), .Z(n10368) );
  AND U9741 ( .A(n1280), .B(n10381), .Z(n10383) );
  XNOR U9742 ( .A(n10382), .B(n10379), .Z(n10381) );
  XOR U9743 ( .A(n10384), .B(n10385), .Z(n10379) );
  AND U9744 ( .A(n1283), .B(n10378), .Z(n10385) );
  XNOR U9745 ( .A(n10386), .B(n10376), .Z(n10378) );
  XOR U9746 ( .A(n10387), .B(n10388), .Z(n10376) );
  AND U9747 ( .A(n1287), .B(n10389), .Z(n10388) );
  XOR U9748 ( .A(p_input[1028]), .B(n10387), .Z(n10389) );
  XOR U9749 ( .A(n10390), .B(n10391), .Z(n10387) );
  AND U9750 ( .A(n1291), .B(n10392), .Z(n10391) );
  IV U9751 ( .A(n10384), .Z(n10386) );
  XOR U9752 ( .A(n10393), .B(n10394), .Z(n10384) );
  AND U9753 ( .A(n1295), .B(n10395), .Z(n10394) );
  XOR U9754 ( .A(n10396), .B(n10397), .Z(n10382) );
  AND U9755 ( .A(n1299), .B(n10395), .Z(n10397) );
  XNOR U9756 ( .A(n10396), .B(n10393), .Z(n10395) );
  XOR U9757 ( .A(n10398), .B(n10399), .Z(n10393) );
  AND U9758 ( .A(n1302), .B(n10392), .Z(n10399) );
  XNOR U9759 ( .A(n10400), .B(n10390), .Z(n10392) );
  XOR U9760 ( .A(n10401), .B(n10402), .Z(n10390) );
  AND U9761 ( .A(n1306), .B(n10403), .Z(n10402) );
  XOR U9762 ( .A(p_input[1044]), .B(n10401), .Z(n10403) );
  XOR U9763 ( .A(n10404), .B(n10405), .Z(n10401) );
  AND U9764 ( .A(n1310), .B(n10406), .Z(n10405) );
  IV U9765 ( .A(n10398), .Z(n10400) );
  XOR U9766 ( .A(n10407), .B(n10408), .Z(n10398) );
  AND U9767 ( .A(n1314), .B(n10409), .Z(n10408) );
  XOR U9768 ( .A(n10410), .B(n10411), .Z(n10396) );
  AND U9769 ( .A(n1318), .B(n10409), .Z(n10411) );
  XNOR U9770 ( .A(n10410), .B(n10407), .Z(n10409) );
  XOR U9771 ( .A(n10412), .B(n10413), .Z(n10407) );
  AND U9772 ( .A(n1321), .B(n10406), .Z(n10413) );
  XNOR U9773 ( .A(n10414), .B(n10404), .Z(n10406) );
  XOR U9774 ( .A(n10415), .B(n10416), .Z(n10404) );
  AND U9775 ( .A(n1325), .B(n10417), .Z(n10416) );
  XOR U9776 ( .A(p_input[1060]), .B(n10415), .Z(n10417) );
  XOR U9777 ( .A(n10418), .B(n10419), .Z(n10415) );
  AND U9778 ( .A(n1329), .B(n10420), .Z(n10419) );
  IV U9779 ( .A(n10412), .Z(n10414) );
  XOR U9780 ( .A(n10421), .B(n10422), .Z(n10412) );
  AND U9781 ( .A(n1333), .B(n10423), .Z(n10422) );
  XOR U9782 ( .A(n10424), .B(n10425), .Z(n10410) );
  AND U9783 ( .A(n1337), .B(n10423), .Z(n10425) );
  XNOR U9784 ( .A(n10424), .B(n10421), .Z(n10423) );
  XOR U9785 ( .A(n10426), .B(n10427), .Z(n10421) );
  AND U9786 ( .A(n1340), .B(n10420), .Z(n10427) );
  XNOR U9787 ( .A(n10428), .B(n10418), .Z(n10420) );
  XOR U9788 ( .A(n10429), .B(n10430), .Z(n10418) );
  AND U9789 ( .A(n1344), .B(n10431), .Z(n10430) );
  XOR U9790 ( .A(p_input[1076]), .B(n10429), .Z(n10431) );
  XOR U9791 ( .A(n10432), .B(n10433), .Z(n10429) );
  AND U9792 ( .A(n1348), .B(n10434), .Z(n10433) );
  IV U9793 ( .A(n10426), .Z(n10428) );
  XOR U9794 ( .A(n10435), .B(n10436), .Z(n10426) );
  AND U9795 ( .A(n1352), .B(n10437), .Z(n10436) );
  XOR U9796 ( .A(n10438), .B(n10439), .Z(n10424) );
  AND U9797 ( .A(n1356), .B(n10437), .Z(n10439) );
  XNOR U9798 ( .A(n10438), .B(n10435), .Z(n10437) );
  XOR U9799 ( .A(n10440), .B(n10441), .Z(n10435) );
  AND U9800 ( .A(n1359), .B(n10434), .Z(n10441) );
  XNOR U9801 ( .A(n10442), .B(n10432), .Z(n10434) );
  XOR U9802 ( .A(n10443), .B(n10444), .Z(n10432) );
  AND U9803 ( .A(n1363), .B(n10445), .Z(n10444) );
  XOR U9804 ( .A(p_input[1092]), .B(n10443), .Z(n10445) );
  XOR U9805 ( .A(n10446), .B(n10447), .Z(n10443) );
  AND U9806 ( .A(n1367), .B(n10448), .Z(n10447) );
  IV U9807 ( .A(n10440), .Z(n10442) );
  XOR U9808 ( .A(n10449), .B(n10450), .Z(n10440) );
  AND U9809 ( .A(n1371), .B(n10451), .Z(n10450) );
  XOR U9810 ( .A(n10452), .B(n10453), .Z(n10438) );
  AND U9811 ( .A(n1375), .B(n10451), .Z(n10453) );
  XNOR U9812 ( .A(n10452), .B(n10449), .Z(n10451) );
  XOR U9813 ( .A(n10454), .B(n10455), .Z(n10449) );
  AND U9814 ( .A(n1378), .B(n10448), .Z(n10455) );
  XNOR U9815 ( .A(n10456), .B(n10446), .Z(n10448) );
  XOR U9816 ( .A(n10457), .B(n10458), .Z(n10446) );
  AND U9817 ( .A(n1382), .B(n10459), .Z(n10458) );
  XOR U9818 ( .A(p_input[1108]), .B(n10457), .Z(n10459) );
  XOR U9819 ( .A(n10460), .B(n10461), .Z(n10457) );
  AND U9820 ( .A(n1386), .B(n10462), .Z(n10461) );
  IV U9821 ( .A(n10454), .Z(n10456) );
  XOR U9822 ( .A(n10463), .B(n10464), .Z(n10454) );
  AND U9823 ( .A(n1390), .B(n10465), .Z(n10464) );
  XOR U9824 ( .A(n10466), .B(n10467), .Z(n10452) );
  AND U9825 ( .A(n1394), .B(n10465), .Z(n10467) );
  XNOR U9826 ( .A(n10466), .B(n10463), .Z(n10465) );
  XOR U9827 ( .A(n10468), .B(n10469), .Z(n10463) );
  AND U9828 ( .A(n1397), .B(n10462), .Z(n10469) );
  XNOR U9829 ( .A(n10470), .B(n10460), .Z(n10462) );
  XOR U9830 ( .A(n10471), .B(n10472), .Z(n10460) );
  AND U9831 ( .A(n1401), .B(n10473), .Z(n10472) );
  XOR U9832 ( .A(p_input[1124]), .B(n10471), .Z(n10473) );
  XOR U9833 ( .A(n10474), .B(n10475), .Z(n10471) );
  AND U9834 ( .A(n1405), .B(n10476), .Z(n10475) );
  IV U9835 ( .A(n10468), .Z(n10470) );
  XOR U9836 ( .A(n10477), .B(n10478), .Z(n10468) );
  AND U9837 ( .A(n1409), .B(n10479), .Z(n10478) );
  XOR U9838 ( .A(n10480), .B(n10481), .Z(n10466) );
  AND U9839 ( .A(n1413), .B(n10479), .Z(n10481) );
  XNOR U9840 ( .A(n10480), .B(n10477), .Z(n10479) );
  XOR U9841 ( .A(n10482), .B(n10483), .Z(n10477) );
  AND U9842 ( .A(n1416), .B(n10476), .Z(n10483) );
  XNOR U9843 ( .A(n10484), .B(n10474), .Z(n10476) );
  XOR U9844 ( .A(n10485), .B(n10486), .Z(n10474) );
  AND U9845 ( .A(n1420), .B(n10487), .Z(n10486) );
  XOR U9846 ( .A(p_input[1140]), .B(n10485), .Z(n10487) );
  XOR U9847 ( .A(n10488), .B(n10489), .Z(n10485) );
  AND U9848 ( .A(n1424), .B(n10490), .Z(n10489) );
  IV U9849 ( .A(n10482), .Z(n10484) );
  XOR U9850 ( .A(n10491), .B(n10492), .Z(n10482) );
  AND U9851 ( .A(n1428), .B(n10493), .Z(n10492) );
  XOR U9852 ( .A(n10494), .B(n10495), .Z(n10480) );
  AND U9853 ( .A(n1432), .B(n10493), .Z(n10495) );
  XNOR U9854 ( .A(n10494), .B(n10491), .Z(n10493) );
  XOR U9855 ( .A(n10496), .B(n10497), .Z(n10491) );
  AND U9856 ( .A(n1435), .B(n10490), .Z(n10497) );
  XNOR U9857 ( .A(n10498), .B(n10488), .Z(n10490) );
  XOR U9858 ( .A(n10499), .B(n10500), .Z(n10488) );
  AND U9859 ( .A(n1439), .B(n10501), .Z(n10500) );
  XOR U9860 ( .A(p_input[1156]), .B(n10499), .Z(n10501) );
  XOR U9861 ( .A(n10502), .B(n10503), .Z(n10499) );
  AND U9862 ( .A(n1443), .B(n10504), .Z(n10503) );
  IV U9863 ( .A(n10496), .Z(n10498) );
  XOR U9864 ( .A(n10505), .B(n10506), .Z(n10496) );
  AND U9865 ( .A(n1447), .B(n10507), .Z(n10506) );
  XOR U9866 ( .A(n10508), .B(n10509), .Z(n10494) );
  AND U9867 ( .A(n1451), .B(n10507), .Z(n10509) );
  XNOR U9868 ( .A(n10508), .B(n10505), .Z(n10507) );
  XOR U9869 ( .A(n10510), .B(n10511), .Z(n10505) );
  AND U9870 ( .A(n1454), .B(n10504), .Z(n10511) );
  XNOR U9871 ( .A(n10512), .B(n10502), .Z(n10504) );
  XOR U9872 ( .A(n10513), .B(n10514), .Z(n10502) );
  AND U9873 ( .A(n1458), .B(n10515), .Z(n10514) );
  XOR U9874 ( .A(p_input[1172]), .B(n10513), .Z(n10515) );
  XOR U9875 ( .A(n10516), .B(n10517), .Z(n10513) );
  AND U9876 ( .A(n1462), .B(n10518), .Z(n10517) );
  IV U9877 ( .A(n10510), .Z(n10512) );
  XOR U9878 ( .A(n10519), .B(n10520), .Z(n10510) );
  AND U9879 ( .A(n1466), .B(n10521), .Z(n10520) );
  XOR U9880 ( .A(n10522), .B(n10523), .Z(n10508) );
  AND U9881 ( .A(n1470), .B(n10521), .Z(n10523) );
  XNOR U9882 ( .A(n10522), .B(n10519), .Z(n10521) );
  XOR U9883 ( .A(n10524), .B(n10525), .Z(n10519) );
  AND U9884 ( .A(n1473), .B(n10518), .Z(n10525) );
  XNOR U9885 ( .A(n10526), .B(n10516), .Z(n10518) );
  XOR U9886 ( .A(n10527), .B(n10528), .Z(n10516) );
  AND U9887 ( .A(n1477), .B(n10529), .Z(n10528) );
  XOR U9888 ( .A(p_input[1188]), .B(n10527), .Z(n10529) );
  XOR U9889 ( .A(n10530), .B(n10531), .Z(n10527) );
  AND U9890 ( .A(n1481), .B(n10532), .Z(n10531) );
  IV U9891 ( .A(n10524), .Z(n10526) );
  XOR U9892 ( .A(n10533), .B(n10534), .Z(n10524) );
  AND U9893 ( .A(n1485), .B(n10535), .Z(n10534) );
  XOR U9894 ( .A(n10536), .B(n10537), .Z(n10522) );
  AND U9895 ( .A(n1489), .B(n10535), .Z(n10537) );
  XNOR U9896 ( .A(n10536), .B(n10533), .Z(n10535) );
  XOR U9897 ( .A(n10538), .B(n10539), .Z(n10533) );
  AND U9898 ( .A(n1492), .B(n10532), .Z(n10539) );
  XNOR U9899 ( .A(n10540), .B(n10530), .Z(n10532) );
  XOR U9900 ( .A(n10541), .B(n10542), .Z(n10530) );
  AND U9901 ( .A(n1496), .B(n10543), .Z(n10542) );
  XOR U9902 ( .A(p_input[1204]), .B(n10541), .Z(n10543) );
  XOR U9903 ( .A(n10544), .B(n10545), .Z(n10541) );
  AND U9904 ( .A(n1500), .B(n10546), .Z(n10545) );
  IV U9905 ( .A(n10538), .Z(n10540) );
  XOR U9906 ( .A(n10547), .B(n10548), .Z(n10538) );
  AND U9907 ( .A(n1504), .B(n10549), .Z(n10548) );
  XOR U9908 ( .A(n10550), .B(n10551), .Z(n10536) );
  AND U9909 ( .A(n1508), .B(n10549), .Z(n10551) );
  XNOR U9910 ( .A(n10550), .B(n10547), .Z(n10549) );
  XOR U9911 ( .A(n10552), .B(n10553), .Z(n10547) );
  AND U9912 ( .A(n1511), .B(n10546), .Z(n10553) );
  XNOR U9913 ( .A(n10554), .B(n10544), .Z(n10546) );
  XOR U9914 ( .A(n10555), .B(n10556), .Z(n10544) );
  AND U9915 ( .A(n1515), .B(n10557), .Z(n10556) );
  XOR U9916 ( .A(p_input[1220]), .B(n10555), .Z(n10557) );
  XOR U9917 ( .A(n10558), .B(n10559), .Z(n10555) );
  AND U9918 ( .A(n1519), .B(n10560), .Z(n10559) );
  IV U9919 ( .A(n10552), .Z(n10554) );
  XOR U9920 ( .A(n10561), .B(n10562), .Z(n10552) );
  AND U9921 ( .A(n1523), .B(n10563), .Z(n10562) );
  XOR U9922 ( .A(n10564), .B(n10565), .Z(n10550) );
  AND U9923 ( .A(n1527), .B(n10563), .Z(n10565) );
  XNOR U9924 ( .A(n10564), .B(n10561), .Z(n10563) );
  XOR U9925 ( .A(n10566), .B(n10567), .Z(n10561) );
  AND U9926 ( .A(n1530), .B(n10560), .Z(n10567) );
  XNOR U9927 ( .A(n10568), .B(n10558), .Z(n10560) );
  XOR U9928 ( .A(n10569), .B(n10570), .Z(n10558) );
  AND U9929 ( .A(n1534), .B(n10571), .Z(n10570) );
  XOR U9930 ( .A(p_input[1236]), .B(n10569), .Z(n10571) );
  XOR U9931 ( .A(n10572), .B(n10573), .Z(n10569) );
  AND U9932 ( .A(n1538), .B(n10574), .Z(n10573) );
  IV U9933 ( .A(n10566), .Z(n10568) );
  XOR U9934 ( .A(n10575), .B(n10576), .Z(n10566) );
  AND U9935 ( .A(n1542), .B(n10577), .Z(n10576) );
  XOR U9936 ( .A(n10578), .B(n10579), .Z(n10564) );
  AND U9937 ( .A(n1546), .B(n10577), .Z(n10579) );
  XNOR U9938 ( .A(n10578), .B(n10575), .Z(n10577) );
  XOR U9939 ( .A(n10580), .B(n10581), .Z(n10575) );
  AND U9940 ( .A(n1549), .B(n10574), .Z(n10581) );
  XNOR U9941 ( .A(n10582), .B(n10572), .Z(n10574) );
  XOR U9942 ( .A(n10583), .B(n10584), .Z(n10572) );
  AND U9943 ( .A(n1553), .B(n10585), .Z(n10584) );
  XOR U9944 ( .A(p_input[1252]), .B(n10583), .Z(n10585) );
  XOR U9945 ( .A(n10586), .B(n10587), .Z(n10583) );
  AND U9946 ( .A(n1557), .B(n10588), .Z(n10587) );
  IV U9947 ( .A(n10580), .Z(n10582) );
  XOR U9948 ( .A(n10589), .B(n10590), .Z(n10580) );
  AND U9949 ( .A(n1561), .B(n10591), .Z(n10590) );
  XOR U9950 ( .A(n10592), .B(n10593), .Z(n10578) );
  AND U9951 ( .A(n1565), .B(n10591), .Z(n10593) );
  XNOR U9952 ( .A(n10592), .B(n10589), .Z(n10591) );
  XOR U9953 ( .A(n10594), .B(n10595), .Z(n10589) );
  AND U9954 ( .A(n1568), .B(n10588), .Z(n10595) );
  XNOR U9955 ( .A(n10596), .B(n10586), .Z(n10588) );
  XOR U9956 ( .A(n10597), .B(n10598), .Z(n10586) );
  AND U9957 ( .A(n1572), .B(n10599), .Z(n10598) );
  XOR U9958 ( .A(p_input[1268]), .B(n10597), .Z(n10599) );
  XOR U9959 ( .A(n10600), .B(n10601), .Z(n10597) );
  AND U9960 ( .A(n1576), .B(n10602), .Z(n10601) );
  IV U9961 ( .A(n10594), .Z(n10596) );
  XOR U9962 ( .A(n10603), .B(n10604), .Z(n10594) );
  AND U9963 ( .A(n1580), .B(n10605), .Z(n10604) );
  XOR U9964 ( .A(n10606), .B(n10607), .Z(n10592) );
  AND U9965 ( .A(n1584), .B(n10605), .Z(n10607) );
  XNOR U9966 ( .A(n10606), .B(n10603), .Z(n10605) );
  XOR U9967 ( .A(n10608), .B(n10609), .Z(n10603) );
  AND U9968 ( .A(n1587), .B(n10602), .Z(n10609) );
  XNOR U9969 ( .A(n10610), .B(n10600), .Z(n10602) );
  XOR U9970 ( .A(n10611), .B(n10612), .Z(n10600) );
  AND U9971 ( .A(n1591), .B(n10613), .Z(n10612) );
  XOR U9972 ( .A(p_input[1284]), .B(n10611), .Z(n10613) );
  XOR U9973 ( .A(n10614), .B(n10615), .Z(n10611) );
  AND U9974 ( .A(n1595), .B(n10616), .Z(n10615) );
  IV U9975 ( .A(n10608), .Z(n10610) );
  XOR U9976 ( .A(n10617), .B(n10618), .Z(n10608) );
  AND U9977 ( .A(n1599), .B(n10619), .Z(n10618) );
  XOR U9978 ( .A(n10620), .B(n10621), .Z(n10606) );
  AND U9979 ( .A(n1603), .B(n10619), .Z(n10621) );
  XNOR U9980 ( .A(n10620), .B(n10617), .Z(n10619) );
  XOR U9981 ( .A(n10622), .B(n10623), .Z(n10617) );
  AND U9982 ( .A(n1606), .B(n10616), .Z(n10623) );
  XNOR U9983 ( .A(n10624), .B(n10614), .Z(n10616) );
  XOR U9984 ( .A(n10625), .B(n10626), .Z(n10614) );
  AND U9985 ( .A(n1610), .B(n10627), .Z(n10626) );
  XOR U9986 ( .A(p_input[1300]), .B(n10625), .Z(n10627) );
  XOR U9987 ( .A(n10628), .B(n10629), .Z(n10625) );
  AND U9988 ( .A(n1614), .B(n10630), .Z(n10629) );
  IV U9989 ( .A(n10622), .Z(n10624) );
  XOR U9990 ( .A(n10631), .B(n10632), .Z(n10622) );
  AND U9991 ( .A(n1618), .B(n10633), .Z(n10632) );
  XOR U9992 ( .A(n10634), .B(n10635), .Z(n10620) );
  AND U9993 ( .A(n1622), .B(n10633), .Z(n10635) );
  XNOR U9994 ( .A(n10634), .B(n10631), .Z(n10633) );
  XOR U9995 ( .A(n10636), .B(n10637), .Z(n10631) );
  AND U9996 ( .A(n1625), .B(n10630), .Z(n10637) );
  XNOR U9997 ( .A(n10638), .B(n10628), .Z(n10630) );
  XOR U9998 ( .A(n10639), .B(n10640), .Z(n10628) );
  AND U9999 ( .A(n1629), .B(n10641), .Z(n10640) );
  XOR U10000 ( .A(p_input[1316]), .B(n10639), .Z(n10641) );
  XOR U10001 ( .A(n10642), .B(n10643), .Z(n10639) );
  AND U10002 ( .A(n1633), .B(n10644), .Z(n10643) );
  IV U10003 ( .A(n10636), .Z(n10638) );
  XOR U10004 ( .A(n10645), .B(n10646), .Z(n10636) );
  AND U10005 ( .A(n1637), .B(n10647), .Z(n10646) );
  XOR U10006 ( .A(n10648), .B(n10649), .Z(n10634) );
  AND U10007 ( .A(n1641), .B(n10647), .Z(n10649) );
  XNOR U10008 ( .A(n10648), .B(n10645), .Z(n10647) );
  XOR U10009 ( .A(n10650), .B(n10651), .Z(n10645) );
  AND U10010 ( .A(n1644), .B(n10644), .Z(n10651) );
  XNOR U10011 ( .A(n10652), .B(n10642), .Z(n10644) );
  XOR U10012 ( .A(n10653), .B(n10654), .Z(n10642) );
  AND U10013 ( .A(n1648), .B(n10655), .Z(n10654) );
  XOR U10014 ( .A(p_input[1332]), .B(n10653), .Z(n10655) );
  XOR U10015 ( .A(n10656), .B(n10657), .Z(n10653) );
  AND U10016 ( .A(n1652), .B(n10658), .Z(n10657) );
  IV U10017 ( .A(n10650), .Z(n10652) );
  XOR U10018 ( .A(n10659), .B(n10660), .Z(n10650) );
  AND U10019 ( .A(n1656), .B(n10661), .Z(n10660) );
  XOR U10020 ( .A(n10662), .B(n10663), .Z(n10648) );
  AND U10021 ( .A(n1660), .B(n10661), .Z(n10663) );
  XNOR U10022 ( .A(n10662), .B(n10659), .Z(n10661) );
  XOR U10023 ( .A(n10664), .B(n10665), .Z(n10659) );
  AND U10024 ( .A(n1663), .B(n10658), .Z(n10665) );
  XNOR U10025 ( .A(n10666), .B(n10656), .Z(n10658) );
  XOR U10026 ( .A(n10667), .B(n10668), .Z(n10656) );
  AND U10027 ( .A(n1667), .B(n10669), .Z(n10668) );
  XOR U10028 ( .A(p_input[1348]), .B(n10667), .Z(n10669) );
  XOR U10029 ( .A(n10670), .B(n10671), .Z(n10667) );
  AND U10030 ( .A(n1671), .B(n10672), .Z(n10671) );
  IV U10031 ( .A(n10664), .Z(n10666) );
  XOR U10032 ( .A(n10673), .B(n10674), .Z(n10664) );
  AND U10033 ( .A(n1675), .B(n10675), .Z(n10674) );
  XOR U10034 ( .A(n10676), .B(n10677), .Z(n10662) );
  AND U10035 ( .A(n1679), .B(n10675), .Z(n10677) );
  XNOR U10036 ( .A(n10676), .B(n10673), .Z(n10675) );
  XOR U10037 ( .A(n10678), .B(n10679), .Z(n10673) );
  AND U10038 ( .A(n1682), .B(n10672), .Z(n10679) );
  XNOR U10039 ( .A(n10680), .B(n10670), .Z(n10672) );
  XOR U10040 ( .A(n10681), .B(n10682), .Z(n10670) );
  AND U10041 ( .A(n1686), .B(n10683), .Z(n10682) );
  XOR U10042 ( .A(p_input[1364]), .B(n10681), .Z(n10683) );
  XOR U10043 ( .A(n10684), .B(n10685), .Z(n10681) );
  AND U10044 ( .A(n1690), .B(n10686), .Z(n10685) );
  IV U10045 ( .A(n10678), .Z(n10680) );
  XOR U10046 ( .A(n10687), .B(n10688), .Z(n10678) );
  AND U10047 ( .A(n1694), .B(n10689), .Z(n10688) );
  XOR U10048 ( .A(n10690), .B(n10691), .Z(n10676) );
  AND U10049 ( .A(n1698), .B(n10689), .Z(n10691) );
  XNOR U10050 ( .A(n10690), .B(n10687), .Z(n10689) );
  XOR U10051 ( .A(n10692), .B(n10693), .Z(n10687) );
  AND U10052 ( .A(n1701), .B(n10686), .Z(n10693) );
  XNOR U10053 ( .A(n10694), .B(n10684), .Z(n10686) );
  XOR U10054 ( .A(n10695), .B(n10696), .Z(n10684) );
  AND U10055 ( .A(n1705), .B(n10697), .Z(n10696) );
  XOR U10056 ( .A(p_input[1380]), .B(n10695), .Z(n10697) );
  XOR U10057 ( .A(n10698), .B(n10699), .Z(n10695) );
  AND U10058 ( .A(n1709), .B(n10700), .Z(n10699) );
  IV U10059 ( .A(n10692), .Z(n10694) );
  XOR U10060 ( .A(n10701), .B(n10702), .Z(n10692) );
  AND U10061 ( .A(n1713), .B(n10703), .Z(n10702) );
  XOR U10062 ( .A(n10704), .B(n10705), .Z(n10690) );
  AND U10063 ( .A(n1717), .B(n10703), .Z(n10705) );
  XNOR U10064 ( .A(n10704), .B(n10701), .Z(n10703) );
  XOR U10065 ( .A(n10706), .B(n10707), .Z(n10701) );
  AND U10066 ( .A(n1720), .B(n10700), .Z(n10707) );
  XNOR U10067 ( .A(n10708), .B(n10698), .Z(n10700) );
  XOR U10068 ( .A(n10709), .B(n10710), .Z(n10698) );
  AND U10069 ( .A(n1724), .B(n10711), .Z(n10710) );
  XOR U10070 ( .A(p_input[1396]), .B(n10709), .Z(n10711) );
  XOR U10071 ( .A(n10712), .B(n10713), .Z(n10709) );
  AND U10072 ( .A(n1728), .B(n10714), .Z(n10713) );
  IV U10073 ( .A(n10706), .Z(n10708) );
  XOR U10074 ( .A(n10715), .B(n10716), .Z(n10706) );
  AND U10075 ( .A(n1732), .B(n10717), .Z(n10716) );
  XOR U10076 ( .A(n10718), .B(n10719), .Z(n10704) );
  AND U10077 ( .A(n1736), .B(n10717), .Z(n10719) );
  XNOR U10078 ( .A(n10718), .B(n10715), .Z(n10717) );
  XOR U10079 ( .A(n10720), .B(n10721), .Z(n10715) );
  AND U10080 ( .A(n1739), .B(n10714), .Z(n10721) );
  XNOR U10081 ( .A(n10722), .B(n10712), .Z(n10714) );
  XOR U10082 ( .A(n10723), .B(n10724), .Z(n10712) );
  AND U10083 ( .A(n1743), .B(n10725), .Z(n10724) );
  XOR U10084 ( .A(p_input[1412]), .B(n10723), .Z(n10725) );
  XOR U10085 ( .A(n10726), .B(n10727), .Z(n10723) );
  AND U10086 ( .A(n1747), .B(n10728), .Z(n10727) );
  IV U10087 ( .A(n10720), .Z(n10722) );
  XOR U10088 ( .A(n10729), .B(n10730), .Z(n10720) );
  AND U10089 ( .A(n1751), .B(n10731), .Z(n10730) );
  XOR U10090 ( .A(n10732), .B(n10733), .Z(n10718) );
  AND U10091 ( .A(n1755), .B(n10731), .Z(n10733) );
  XNOR U10092 ( .A(n10732), .B(n10729), .Z(n10731) );
  XOR U10093 ( .A(n10734), .B(n10735), .Z(n10729) );
  AND U10094 ( .A(n1758), .B(n10728), .Z(n10735) );
  XNOR U10095 ( .A(n10736), .B(n10726), .Z(n10728) );
  XOR U10096 ( .A(n10737), .B(n10738), .Z(n10726) );
  AND U10097 ( .A(n1762), .B(n10739), .Z(n10738) );
  XOR U10098 ( .A(p_input[1428]), .B(n10737), .Z(n10739) );
  XOR U10099 ( .A(n10740), .B(n10741), .Z(n10737) );
  AND U10100 ( .A(n1766), .B(n10742), .Z(n10741) );
  IV U10101 ( .A(n10734), .Z(n10736) );
  XOR U10102 ( .A(n10743), .B(n10744), .Z(n10734) );
  AND U10103 ( .A(n1770), .B(n10745), .Z(n10744) );
  XOR U10104 ( .A(n10746), .B(n10747), .Z(n10732) );
  AND U10105 ( .A(n1774), .B(n10745), .Z(n10747) );
  XNOR U10106 ( .A(n10746), .B(n10743), .Z(n10745) );
  XOR U10107 ( .A(n10748), .B(n10749), .Z(n10743) );
  AND U10108 ( .A(n1777), .B(n10742), .Z(n10749) );
  XNOR U10109 ( .A(n10750), .B(n10740), .Z(n10742) );
  XOR U10110 ( .A(n10751), .B(n10752), .Z(n10740) );
  AND U10111 ( .A(n1781), .B(n10753), .Z(n10752) );
  XOR U10112 ( .A(p_input[1444]), .B(n10751), .Z(n10753) );
  XOR U10113 ( .A(n10754), .B(n10755), .Z(n10751) );
  AND U10114 ( .A(n1785), .B(n10756), .Z(n10755) );
  IV U10115 ( .A(n10748), .Z(n10750) );
  XOR U10116 ( .A(n10757), .B(n10758), .Z(n10748) );
  AND U10117 ( .A(n1789), .B(n10759), .Z(n10758) );
  XOR U10118 ( .A(n10760), .B(n10761), .Z(n10746) );
  AND U10119 ( .A(n1793), .B(n10759), .Z(n10761) );
  XNOR U10120 ( .A(n10760), .B(n10757), .Z(n10759) );
  XOR U10121 ( .A(n10762), .B(n10763), .Z(n10757) );
  AND U10122 ( .A(n1796), .B(n10756), .Z(n10763) );
  XNOR U10123 ( .A(n10764), .B(n10754), .Z(n10756) );
  XOR U10124 ( .A(n10765), .B(n10766), .Z(n10754) );
  AND U10125 ( .A(n1800), .B(n10767), .Z(n10766) );
  XOR U10126 ( .A(p_input[1460]), .B(n10765), .Z(n10767) );
  XOR U10127 ( .A(n10768), .B(n10769), .Z(n10765) );
  AND U10128 ( .A(n1804), .B(n10770), .Z(n10769) );
  IV U10129 ( .A(n10762), .Z(n10764) );
  XOR U10130 ( .A(n10771), .B(n10772), .Z(n10762) );
  AND U10131 ( .A(n1808), .B(n10773), .Z(n10772) );
  XOR U10132 ( .A(n10774), .B(n10775), .Z(n10760) );
  AND U10133 ( .A(n1812), .B(n10773), .Z(n10775) );
  XNOR U10134 ( .A(n10774), .B(n10771), .Z(n10773) );
  XOR U10135 ( .A(n10776), .B(n10777), .Z(n10771) );
  AND U10136 ( .A(n1815), .B(n10770), .Z(n10777) );
  XNOR U10137 ( .A(n10778), .B(n10768), .Z(n10770) );
  XOR U10138 ( .A(n10779), .B(n10780), .Z(n10768) );
  AND U10139 ( .A(n1819), .B(n10781), .Z(n10780) );
  XOR U10140 ( .A(p_input[1476]), .B(n10779), .Z(n10781) );
  XOR U10141 ( .A(n10782), .B(n10783), .Z(n10779) );
  AND U10142 ( .A(n1823), .B(n10784), .Z(n10783) );
  IV U10143 ( .A(n10776), .Z(n10778) );
  XOR U10144 ( .A(n10785), .B(n10786), .Z(n10776) );
  AND U10145 ( .A(n1827), .B(n10787), .Z(n10786) );
  XOR U10146 ( .A(n10788), .B(n10789), .Z(n10774) );
  AND U10147 ( .A(n1831), .B(n10787), .Z(n10789) );
  XNOR U10148 ( .A(n10788), .B(n10785), .Z(n10787) );
  XOR U10149 ( .A(n10790), .B(n10791), .Z(n10785) );
  AND U10150 ( .A(n1834), .B(n10784), .Z(n10791) );
  XNOR U10151 ( .A(n10792), .B(n10782), .Z(n10784) );
  XOR U10152 ( .A(n10793), .B(n10794), .Z(n10782) );
  AND U10153 ( .A(n1838), .B(n10795), .Z(n10794) );
  XOR U10154 ( .A(p_input[1492]), .B(n10793), .Z(n10795) );
  XOR U10155 ( .A(n10796), .B(n10797), .Z(n10793) );
  AND U10156 ( .A(n1842), .B(n10798), .Z(n10797) );
  IV U10157 ( .A(n10790), .Z(n10792) );
  XOR U10158 ( .A(n10799), .B(n10800), .Z(n10790) );
  AND U10159 ( .A(n1846), .B(n10801), .Z(n10800) );
  XOR U10160 ( .A(n10802), .B(n10803), .Z(n10788) );
  AND U10161 ( .A(n1850), .B(n10801), .Z(n10803) );
  XNOR U10162 ( .A(n10802), .B(n10799), .Z(n10801) );
  XOR U10163 ( .A(n10804), .B(n10805), .Z(n10799) );
  AND U10164 ( .A(n1853), .B(n10798), .Z(n10805) );
  XNOR U10165 ( .A(n10806), .B(n10796), .Z(n10798) );
  XOR U10166 ( .A(n10807), .B(n10808), .Z(n10796) );
  AND U10167 ( .A(n1857), .B(n10809), .Z(n10808) );
  XOR U10168 ( .A(p_input[1508]), .B(n10807), .Z(n10809) );
  XOR U10169 ( .A(n10810), .B(n10811), .Z(n10807) );
  AND U10170 ( .A(n1861), .B(n10812), .Z(n10811) );
  IV U10171 ( .A(n10804), .Z(n10806) );
  XOR U10172 ( .A(n10813), .B(n10814), .Z(n10804) );
  AND U10173 ( .A(n1865), .B(n10815), .Z(n10814) );
  XOR U10174 ( .A(n10816), .B(n10817), .Z(n10802) );
  AND U10175 ( .A(n1869), .B(n10815), .Z(n10817) );
  XNOR U10176 ( .A(n10816), .B(n10813), .Z(n10815) );
  XOR U10177 ( .A(n10818), .B(n10819), .Z(n10813) );
  AND U10178 ( .A(n1872), .B(n10812), .Z(n10819) );
  XNOR U10179 ( .A(n10820), .B(n10810), .Z(n10812) );
  XOR U10180 ( .A(n10821), .B(n10822), .Z(n10810) );
  AND U10181 ( .A(n1876), .B(n10823), .Z(n10822) );
  XOR U10182 ( .A(p_input[1524]), .B(n10821), .Z(n10823) );
  XOR U10183 ( .A(n10824), .B(n10825), .Z(n10821) );
  AND U10184 ( .A(n1880), .B(n10826), .Z(n10825) );
  IV U10185 ( .A(n10818), .Z(n10820) );
  XOR U10186 ( .A(n10827), .B(n10828), .Z(n10818) );
  AND U10187 ( .A(n1884), .B(n10829), .Z(n10828) );
  XOR U10188 ( .A(n10830), .B(n10831), .Z(n10816) );
  AND U10189 ( .A(n1888), .B(n10829), .Z(n10831) );
  XNOR U10190 ( .A(n10830), .B(n10827), .Z(n10829) );
  XOR U10191 ( .A(n10832), .B(n10833), .Z(n10827) );
  AND U10192 ( .A(n1891), .B(n10826), .Z(n10833) );
  XNOR U10193 ( .A(n10834), .B(n10824), .Z(n10826) );
  XOR U10194 ( .A(n10835), .B(n10836), .Z(n10824) );
  AND U10195 ( .A(n1895), .B(n10837), .Z(n10836) );
  XOR U10196 ( .A(p_input[1540]), .B(n10835), .Z(n10837) );
  XOR U10197 ( .A(n10838), .B(n10839), .Z(n10835) );
  AND U10198 ( .A(n1899), .B(n10840), .Z(n10839) );
  IV U10199 ( .A(n10832), .Z(n10834) );
  XOR U10200 ( .A(n10841), .B(n10842), .Z(n10832) );
  AND U10201 ( .A(n1903), .B(n10843), .Z(n10842) );
  XOR U10202 ( .A(n10844), .B(n10845), .Z(n10830) );
  AND U10203 ( .A(n1907), .B(n10843), .Z(n10845) );
  XNOR U10204 ( .A(n10844), .B(n10841), .Z(n10843) );
  XOR U10205 ( .A(n10846), .B(n10847), .Z(n10841) );
  AND U10206 ( .A(n1910), .B(n10840), .Z(n10847) );
  XNOR U10207 ( .A(n10848), .B(n10838), .Z(n10840) );
  XOR U10208 ( .A(n10849), .B(n10850), .Z(n10838) );
  AND U10209 ( .A(n1914), .B(n10851), .Z(n10850) );
  XOR U10210 ( .A(p_input[1556]), .B(n10849), .Z(n10851) );
  XOR U10211 ( .A(n10852), .B(n10853), .Z(n10849) );
  AND U10212 ( .A(n1918), .B(n10854), .Z(n10853) );
  IV U10213 ( .A(n10846), .Z(n10848) );
  XOR U10214 ( .A(n10855), .B(n10856), .Z(n10846) );
  AND U10215 ( .A(n1922), .B(n10857), .Z(n10856) );
  XOR U10216 ( .A(n10858), .B(n10859), .Z(n10844) );
  AND U10217 ( .A(n1926), .B(n10857), .Z(n10859) );
  XNOR U10218 ( .A(n10858), .B(n10855), .Z(n10857) );
  XOR U10219 ( .A(n10860), .B(n10861), .Z(n10855) );
  AND U10220 ( .A(n1929), .B(n10854), .Z(n10861) );
  XNOR U10221 ( .A(n10862), .B(n10852), .Z(n10854) );
  XOR U10222 ( .A(n10863), .B(n10864), .Z(n10852) );
  AND U10223 ( .A(n1933), .B(n10865), .Z(n10864) );
  XOR U10224 ( .A(p_input[1572]), .B(n10863), .Z(n10865) );
  XOR U10225 ( .A(n10866), .B(n10867), .Z(n10863) );
  AND U10226 ( .A(n1937), .B(n10868), .Z(n10867) );
  IV U10227 ( .A(n10860), .Z(n10862) );
  XOR U10228 ( .A(n10869), .B(n10870), .Z(n10860) );
  AND U10229 ( .A(n1941), .B(n10871), .Z(n10870) );
  XOR U10230 ( .A(n10872), .B(n10873), .Z(n10858) );
  AND U10231 ( .A(n1945), .B(n10871), .Z(n10873) );
  XNOR U10232 ( .A(n10872), .B(n10869), .Z(n10871) );
  XOR U10233 ( .A(n10874), .B(n10875), .Z(n10869) );
  AND U10234 ( .A(n1948), .B(n10868), .Z(n10875) );
  XNOR U10235 ( .A(n10876), .B(n10866), .Z(n10868) );
  XOR U10236 ( .A(n10877), .B(n10878), .Z(n10866) );
  AND U10237 ( .A(n1952), .B(n10879), .Z(n10878) );
  XOR U10238 ( .A(p_input[1588]), .B(n10877), .Z(n10879) );
  XOR U10239 ( .A(n10880), .B(n10881), .Z(n10877) );
  AND U10240 ( .A(n1956), .B(n10882), .Z(n10881) );
  IV U10241 ( .A(n10874), .Z(n10876) );
  XOR U10242 ( .A(n10883), .B(n10884), .Z(n10874) );
  AND U10243 ( .A(n1960), .B(n10885), .Z(n10884) );
  XOR U10244 ( .A(n10886), .B(n10887), .Z(n10872) );
  AND U10245 ( .A(n1964), .B(n10885), .Z(n10887) );
  XNOR U10246 ( .A(n10886), .B(n10883), .Z(n10885) );
  XOR U10247 ( .A(n10888), .B(n10889), .Z(n10883) );
  AND U10248 ( .A(n1967), .B(n10882), .Z(n10889) );
  XNOR U10249 ( .A(n10890), .B(n10880), .Z(n10882) );
  XOR U10250 ( .A(n10891), .B(n10892), .Z(n10880) );
  AND U10251 ( .A(n1971), .B(n10893), .Z(n10892) );
  XOR U10252 ( .A(p_input[1604]), .B(n10891), .Z(n10893) );
  XOR U10253 ( .A(n10894), .B(n10895), .Z(n10891) );
  AND U10254 ( .A(n1975), .B(n10896), .Z(n10895) );
  IV U10255 ( .A(n10888), .Z(n10890) );
  XOR U10256 ( .A(n10897), .B(n10898), .Z(n10888) );
  AND U10257 ( .A(n1979), .B(n10899), .Z(n10898) );
  XOR U10258 ( .A(n10900), .B(n10901), .Z(n10886) );
  AND U10259 ( .A(n1983), .B(n10899), .Z(n10901) );
  XNOR U10260 ( .A(n10900), .B(n10897), .Z(n10899) );
  XOR U10261 ( .A(n10902), .B(n10903), .Z(n10897) );
  AND U10262 ( .A(n1986), .B(n10896), .Z(n10903) );
  XNOR U10263 ( .A(n10904), .B(n10894), .Z(n10896) );
  XOR U10264 ( .A(n10905), .B(n10906), .Z(n10894) );
  AND U10265 ( .A(n1990), .B(n10907), .Z(n10906) );
  XOR U10266 ( .A(p_input[1620]), .B(n10905), .Z(n10907) );
  XOR U10267 ( .A(n10908), .B(n10909), .Z(n10905) );
  AND U10268 ( .A(n1994), .B(n10910), .Z(n10909) );
  IV U10269 ( .A(n10902), .Z(n10904) );
  XOR U10270 ( .A(n10911), .B(n10912), .Z(n10902) );
  AND U10271 ( .A(n1998), .B(n10913), .Z(n10912) );
  XOR U10272 ( .A(n10914), .B(n10915), .Z(n10900) );
  AND U10273 ( .A(n2002), .B(n10913), .Z(n10915) );
  XNOR U10274 ( .A(n10914), .B(n10911), .Z(n10913) );
  XOR U10275 ( .A(n10916), .B(n10917), .Z(n10911) );
  AND U10276 ( .A(n2005), .B(n10910), .Z(n10917) );
  XNOR U10277 ( .A(n10918), .B(n10908), .Z(n10910) );
  XOR U10278 ( .A(n10919), .B(n10920), .Z(n10908) );
  AND U10279 ( .A(n2009), .B(n10921), .Z(n10920) );
  XOR U10280 ( .A(p_input[1636]), .B(n10919), .Z(n10921) );
  XOR U10281 ( .A(n10922), .B(n10923), .Z(n10919) );
  AND U10282 ( .A(n2013), .B(n10924), .Z(n10923) );
  IV U10283 ( .A(n10916), .Z(n10918) );
  XOR U10284 ( .A(n10925), .B(n10926), .Z(n10916) );
  AND U10285 ( .A(n2017), .B(n10927), .Z(n10926) );
  XOR U10286 ( .A(n10928), .B(n10929), .Z(n10914) );
  AND U10287 ( .A(n2021), .B(n10927), .Z(n10929) );
  XNOR U10288 ( .A(n10928), .B(n10925), .Z(n10927) );
  XOR U10289 ( .A(n10930), .B(n10931), .Z(n10925) );
  AND U10290 ( .A(n2024), .B(n10924), .Z(n10931) );
  XNOR U10291 ( .A(n10932), .B(n10922), .Z(n10924) );
  XOR U10292 ( .A(n10933), .B(n10934), .Z(n10922) );
  AND U10293 ( .A(n2028), .B(n10935), .Z(n10934) );
  XOR U10294 ( .A(p_input[1652]), .B(n10933), .Z(n10935) );
  XOR U10295 ( .A(n10936), .B(n10937), .Z(n10933) );
  AND U10296 ( .A(n2032), .B(n10938), .Z(n10937) );
  IV U10297 ( .A(n10930), .Z(n10932) );
  XOR U10298 ( .A(n10939), .B(n10940), .Z(n10930) );
  AND U10299 ( .A(n2036), .B(n10941), .Z(n10940) );
  XOR U10300 ( .A(n10942), .B(n10943), .Z(n10928) );
  AND U10301 ( .A(n2040), .B(n10941), .Z(n10943) );
  XNOR U10302 ( .A(n10942), .B(n10939), .Z(n10941) );
  XOR U10303 ( .A(n10944), .B(n10945), .Z(n10939) );
  AND U10304 ( .A(n2043), .B(n10938), .Z(n10945) );
  XNOR U10305 ( .A(n10946), .B(n10936), .Z(n10938) );
  XOR U10306 ( .A(n10947), .B(n10948), .Z(n10936) );
  AND U10307 ( .A(n2047), .B(n10949), .Z(n10948) );
  XOR U10308 ( .A(p_input[1668]), .B(n10947), .Z(n10949) );
  XOR U10309 ( .A(n10950), .B(n10951), .Z(n10947) );
  AND U10310 ( .A(n2051), .B(n10952), .Z(n10951) );
  IV U10311 ( .A(n10944), .Z(n10946) );
  XOR U10312 ( .A(n10953), .B(n10954), .Z(n10944) );
  AND U10313 ( .A(n2055), .B(n10955), .Z(n10954) );
  XOR U10314 ( .A(n10956), .B(n10957), .Z(n10942) );
  AND U10315 ( .A(n2059), .B(n10955), .Z(n10957) );
  XNOR U10316 ( .A(n10956), .B(n10953), .Z(n10955) );
  XOR U10317 ( .A(n10958), .B(n10959), .Z(n10953) );
  AND U10318 ( .A(n2062), .B(n10952), .Z(n10959) );
  XNOR U10319 ( .A(n10960), .B(n10950), .Z(n10952) );
  XOR U10320 ( .A(n10961), .B(n10962), .Z(n10950) );
  AND U10321 ( .A(n2066), .B(n10963), .Z(n10962) );
  XOR U10322 ( .A(p_input[1684]), .B(n10961), .Z(n10963) );
  XOR U10323 ( .A(n10964), .B(n10965), .Z(n10961) );
  AND U10324 ( .A(n2070), .B(n10966), .Z(n10965) );
  IV U10325 ( .A(n10958), .Z(n10960) );
  XOR U10326 ( .A(n10967), .B(n10968), .Z(n10958) );
  AND U10327 ( .A(n2074), .B(n10969), .Z(n10968) );
  XOR U10328 ( .A(n10970), .B(n10971), .Z(n10956) );
  AND U10329 ( .A(n2078), .B(n10969), .Z(n10971) );
  XNOR U10330 ( .A(n10970), .B(n10967), .Z(n10969) );
  XOR U10331 ( .A(n10972), .B(n10973), .Z(n10967) );
  AND U10332 ( .A(n2081), .B(n10966), .Z(n10973) );
  XNOR U10333 ( .A(n10974), .B(n10964), .Z(n10966) );
  XOR U10334 ( .A(n10975), .B(n10976), .Z(n10964) );
  AND U10335 ( .A(n2085), .B(n10977), .Z(n10976) );
  XOR U10336 ( .A(p_input[1700]), .B(n10975), .Z(n10977) );
  XOR U10337 ( .A(n10978), .B(n10979), .Z(n10975) );
  AND U10338 ( .A(n2089), .B(n10980), .Z(n10979) );
  IV U10339 ( .A(n10972), .Z(n10974) );
  XOR U10340 ( .A(n10981), .B(n10982), .Z(n10972) );
  AND U10341 ( .A(n2093), .B(n10983), .Z(n10982) );
  XOR U10342 ( .A(n10984), .B(n10985), .Z(n10970) );
  AND U10343 ( .A(n2097), .B(n10983), .Z(n10985) );
  XNOR U10344 ( .A(n10984), .B(n10981), .Z(n10983) );
  XOR U10345 ( .A(n10986), .B(n10987), .Z(n10981) );
  AND U10346 ( .A(n2100), .B(n10980), .Z(n10987) );
  XNOR U10347 ( .A(n10988), .B(n10978), .Z(n10980) );
  XOR U10348 ( .A(n10989), .B(n10990), .Z(n10978) );
  AND U10349 ( .A(n2104), .B(n10991), .Z(n10990) );
  XOR U10350 ( .A(p_input[1716]), .B(n10989), .Z(n10991) );
  XOR U10351 ( .A(n10992), .B(n10993), .Z(n10989) );
  AND U10352 ( .A(n2108), .B(n10994), .Z(n10993) );
  IV U10353 ( .A(n10986), .Z(n10988) );
  XOR U10354 ( .A(n10995), .B(n10996), .Z(n10986) );
  AND U10355 ( .A(n2112), .B(n10997), .Z(n10996) );
  XOR U10356 ( .A(n10998), .B(n10999), .Z(n10984) );
  AND U10357 ( .A(n2116), .B(n10997), .Z(n10999) );
  XNOR U10358 ( .A(n10998), .B(n10995), .Z(n10997) );
  XOR U10359 ( .A(n11000), .B(n11001), .Z(n10995) );
  AND U10360 ( .A(n2119), .B(n10994), .Z(n11001) );
  XNOR U10361 ( .A(n11002), .B(n10992), .Z(n10994) );
  XOR U10362 ( .A(n11003), .B(n11004), .Z(n10992) );
  AND U10363 ( .A(n2123), .B(n11005), .Z(n11004) );
  XOR U10364 ( .A(p_input[1732]), .B(n11003), .Z(n11005) );
  XOR U10365 ( .A(n11006), .B(n11007), .Z(n11003) );
  AND U10366 ( .A(n2127), .B(n11008), .Z(n11007) );
  IV U10367 ( .A(n11000), .Z(n11002) );
  XOR U10368 ( .A(n11009), .B(n11010), .Z(n11000) );
  AND U10369 ( .A(n2131), .B(n11011), .Z(n11010) );
  XOR U10370 ( .A(n11012), .B(n11013), .Z(n10998) );
  AND U10371 ( .A(n2135), .B(n11011), .Z(n11013) );
  XNOR U10372 ( .A(n11012), .B(n11009), .Z(n11011) );
  XOR U10373 ( .A(n11014), .B(n11015), .Z(n11009) );
  AND U10374 ( .A(n2138), .B(n11008), .Z(n11015) );
  XNOR U10375 ( .A(n11016), .B(n11006), .Z(n11008) );
  XOR U10376 ( .A(n11017), .B(n11018), .Z(n11006) );
  AND U10377 ( .A(n2142), .B(n11019), .Z(n11018) );
  XOR U10378 ( .A(p_input[1748]), .B(n11017), .Z(n11019) );
  XOR U10379 ( .A(n11020), .B(n11021), .Z(n11017) );
  AND U10380 ( .A(n2146), .B(n11022), .Z(n11021) );
  IV U10381 ( .A(n11014), .Z(n11016) );
  XOR U10382 ( .A(n11023), .B(n11024), .Z(n11014) );
  AND U10383 ( .A(n2150), .B(n11025), .Z(n11024) );
  XOR U10384 ( .A(n11026), .B(n11027), .Z(n11012) );
  AND U10385 ( .A(n2154), .B(n11025), .Z(n11027) );
  XNOR U10386 ( .A(n11026), .B(n11023), .Z(n11025) );
  XOR U10387 ( .A(n11028), .B(n11029), .Z(n11023) );
  AND U10388 ( .A(n2157), .B(n11022), .Z(n11029) );
  XNOR U10389 ( .A(n11030), .B(n11020), .Z(n11022) );
  XOR U10390 ( .A(n11031), .B(n11032), .Z(n11020) );
  AND U10391 ( .A(n2161), .B(n11033), .Z(n11032) );
  XOR U10392 ( .A(p_input[1764]), .B(n11031), .Z(n11033) );
  XOR U10393 ( .A(n11034), .B(n11035), .Z(n11031) );
  AND U10394 ( .A(n2165), .B(n11036), .Z(n11035) );
  IV U10395 ( .A(n11028), .Z(n11030) );
  XOR U10396 ( .A(n11037), .B(n11038), .Z(n11028) );
  AND U10397 ( .A(n2169), .B(n11039), .Z(n11038) );
  XOR U10398 ( .A(n11040), .B(n11041), .Z(n11026) );
  AND U10399 ( .A(n2173), .B(n11039), .Z(n11041) );
  XNOR U10400 ( .A(n11040), .B(n11037), .Z(n11039) );
  XOR U10401 ( .A(n11042), .B(n11043), .Z(n11037) );
  AND U10402 ( .A(n2176), .B(n11036), .Z(n11043) );
  XNOR U10403 ( .A(n11044), .B(n11034), .Z(n11036) );
  XOR U10404 ( .A(n11045), .B(n11046), .Z(n11034) );
  AND U10405 ( .A(n2180), .B(n11047), .Z(n11046) );
  XOR U10406 ( .A(p_input[1780]), .B(n11045), .Z(n11047) );
  XOR U10407 ( .A(n11048), .B(n11049), .Z(n11045) );
  AND U10408 ( .A(n2184), .B(n11050), .Z(n11049) );
  IV U10409 ( .A(n11042), .Z(n11044) );
  XOR U10410 ( .A(n11051), .B(n11052), .Z(n11042) );
  AND U10411 ( .A(n2188), .B(n11053), .Z(n11052) );
  XOR U10412 ( .A(n11054), .B(n11055), .Z(n11040) );
  AND U10413 ( .A(n2192), .B(n11053), .Z(n11055) );
  XNOR U10414 ( .A(n11054), .B(n11051), .Z(n11053) );
  XOR U10415 ( .A(n11056), .B(n11057), .Z(n11051) );
  AND U10416 ( .A(n2195), .B(n11050), .Z(n11057) );
  XNOR U10417 ( .A(n11058), .B(n11048), .Z(n11050) );
  XOR U10418 ( .A(n11059), .B(n11060), .Z(n11048) );
  AND U10419 ( .A(n2199), .B(n11061), .Z(n11060) );
  XOR U10420 ( .A(p_input[1796]), .B(n11059), .Z(n11061) );
  XOR U10421 ( .A(n11062), .B(n11063), .Z(n11059) );
  AND U10422 ( .A(n2203), .B(n11064), .Z(n11063) );
  IV U10423 ( .A(n11056), .Z(n11058) );
  XOR U10424 ( .A(n11065), .B(n11066), .Z(n11056) );
  AND U10425 ( .A(n2207), .B(n11067), .Z(n11066) );
  XOR U10426 ( .A(n11068), .B(n11069), .Z(n11054) );
  AND U10427 ( .A(n2211), .B(n11067), .Z(n11069) );
  XNOR U10428 ( .A(n11068), .B(n11065), .Z(n11067) );
  XOR U10429 ( .A(n11070), .B(n11071), .Z(n11065) );
  AND U10430 ( .A(n2214), .B(n11064), .Z(n11071) );
  XNOR U10431 ( .A(n11072), .B(n11062), .Z(n11064) );
  XOR U10432 ( .A(n11073), .B(n11074), .Z(n11062) );
  AND U10433 ( .A(n2218), .B(n11075), .Z(n11074) );
  XOR U10434 ( .A(p_input[1812]), .B(n11073), .Z(n11075) );
  XOR U10435 ( .A(n11076), .B(n11077), .Z(n11073) );
  AND U10436 ( .A(n2222), .B(n11078), .Z(n11077) );
  IV U10437 ( .A(n11070), .Z(n11072) );
  XOR U10438 ( .A(n11079), .B(n11080), .Z(n11070) );
  AND U10439 ( .A(n2226), .B(n11081), .Z(n11080) );
  XOR U10440 ( .A(n11082), .B(n11083), .Z(n11068) );
  AND U10441 ( .A(n2230), .B(n11081), .Z(n11083) );
  XNOR U10442 ( .A(n11082), .B(n11079), .Z(n11081) );
  XOR U10443 ( .A(n11084), .B(n11085), .Z(n11079) );
  AND U10444 ( .A(n2233), .B(n11078), .Z(n11085) );
  XNOR U10445 ( .A(n11086), .B(n11076), .Z(n11078) );
  XOR U10446 ( .A(n11087), .B(n11088), .Z(n11076) );
  AND U10447 ( .A(n2237), .B(n11089), .Z(n11088) );
  XOR U10448 ( .A(p_input[1828]), .B(n11087), .Z(n11089) );
  XOR U10449 ( .A(n11090), .B(n11091), .Z(n11087) );
  AND U10450 ( .A(n2241), .B(n11092), .Z(n11091) );
  IV U10451 ( .A(n11084), .Z(n11086) );
  XOR U10452 ( .A(n11093), .B(n11094), .Z(n11084) );
  AND U10453 ( .A(n2245), .B(n11095), .Z(n11094) );
  XOR U10454 ( .A(n11096), .B(n11097), .Z(n11082) );
  AND U10455 ( .A(n2249), .B(n11095), .Z(n11097) );
  XNOR U10456 ( .A(n11096), .B(n11093), .Z(n11095) );
  XOR U10457 ( .A(n11098), .B(n11099), .Z(n11093) );
  AND U10458 ( .A(n2252), .B(n11092), .Z(n11099) );
  XNOR U10459 ( .A(n11100), .B(n11090), .Z(n11092) );
  XOR U10460 ( .A(n11101), .B(n11102), .Z(n11090) );
  AND U10461 ( .A(n2256), .B(n11103), .Z(n11102) );
  XOR U10462 ( .A(p_input[1844]), .B(n11101), .Z(n11103) );
  XOR U10463 ( .A(n11104), .B(n11105), .Z(n11101) );
  AND U10464 ( .A(n2260), .B(n11106), .Z(n11105) );
  IV U10465 ( .A(n11098), .Z(n11100) );
  XOR U10466 ( .A(n11107), .B(n11108), .Z(n11098) );
  AND U10467 ( .A(n2264), .B(n11109), .Z(n11108) );
  XOR U10468 ( .A(n11110), .B(n11111), .Z(n11096) );
  AND U10469 ( .A(n2268), .B(n11109), .Z(n11111) );
  XNOR U10470 ( .A(n11110), .B(n11107), .Z(n11109) );
  XOR U10471 ( .A(n11112), .B(n11113), .Z(n11107) );
  AND U10472 ( .A(n2271), .B(n11106), .Z(n11113) );
  XNOR U10473 ( .A(n11114), .B(n11104), .Z(n11106) );
  XOR U10474 ( .A(n11115), .B(n11116), .Z(n11104) );
  AND U10475 ( .A(n2275), .B(n11117), .Z(n11116) );
  XOR U10476 ( .A(p_input[1860]), .B(n11115), .Z(n11117) );
  XOR U10477 ( .A(n11118), .B(n11119), .Z(n11115) );
  AND U10478 ( .A(n2279), .B(n11120), .Z(n11119) );
  IV U10479 ( .A(n11112), .Z(n11114) );
  XOR U10480 ( .A(n11121), .B(n11122), .Z(n11112) );
  AND U10481 ( .A(n2283), .B(n11123), .Z(n11122) );
  XOR U10482 ( .A(n11124), .B(n11125), .Z(n11110) );
  AND U10483 ( .A(n2287), .B(n11123), .Z(n11125) );
  XNOR U10484 ( .A(n11124), .B(n11121), .Z(n11123) );
  XOR U10485 ( .A(n11126), .B(n11127), .Z(n11121) );
  AND U10486 ( .A(n2290), .B(n11120), .Z(n11127) );
  XNOR U10487 ( .A(n11128), .B(n11118), .Z(n11120) );
  XOR U10488 ( .A(n11129), .B(n11130), .Z(n11118) );
  AND U10489 ( .A(n2294), .B(n11131), .Z(n11130) );
  XOR U10490 ( .A(p_input[1876]), .B(n11129), .Z(n11131) );
  XOR U10491 ( .A(n11132), .B(n11133), .Z(n11129) );
  AND U10492 ( .A(n2298), .B(n11134), .Z(n11133) );
  IV U10493 ( .A(n11126), .Z(n11128) );
  XOR U10494 ( .A(n11135), .B(n11136), .Z(n11126) );
  AND U10495 ( .A(n2302), .B(n11137), .Z(n11136) );
  XOR U10496 ( .A(n11138), .B(n11139), .Z(n11124) );
  AND U10497 ( .A(n2306), .B(n11137), .Z(n11139) );
  XNOR U10498 ( .A(n11138), .B(n11135), .Z(n11137) );
  XOR U10499 ( .A(n11140), .B(n11141), .Z(n11135) );
  AND U10500 ( .A(n2309), .B(n11134), .Z(n11141) );
  XNOR U10501 ( .A(n11142), .B(n11132), .Z(n11134) );
  XOR U10502 ( .A(n11143), .B(n11144), .Z(n11132) );
  AND U10503 ( .A(n2313), .B(n11145), .Z(n11144) );
  XOR U10504 ( .A(p_input[1892]), .B(n11143), .Z(n11145) );
  XOR U10505 ( .A(n11146), .B(n11147), .Z(n11143) );
  AND U10506 ( .A(n2317), .B(n11148), .Z(n11147) );
  IV U10507 ( .A(n11140), .Z(n11142) );
  XOR U10508 ( .A(n11149), .B(n11150), .Z(n11140) );
  AND U10509 ( .A(n2321), .B(n11151), .Z(n11150) );
  XOR U10510 ( .A(n11152), .B(n11153), .Z(n11138) );
  AND U10511 ( .A(n2325), .B(n11151), .Z(n11153) );
  XNOR U10512 ( .A(n11152), .B(n11149), .Z(n11151) );
  XOR U10513 ( .A(n11154), .B(n11155), .Z(n11149) );
  AND U10514 ( .A(n2328), .B(n11148), .Z(n11155) );
  XNOR U10515 ( .A(n11156), .B(n11146), .Z(n11148) );
  XOR U10516 ( .A(n11157), .B(n11158), .Z(n11146) );
  AND U10517 ( .A(n2332), .B(n11159), .Z(n11158) );
  XOR U10518 ( .A(p_input[1908]), .B(n11157), .Z(n11159) );
  XOR U10519 ( .A(n11160), .B(n11161), .Z(n11157) );
  AND U10520 ( .A(n2336), .B(n11162), .Z(n11161) );
  IV U10521 ( .A(n11154), .Z(n11156) );
  XOR U10522 ( .A(n11163), .B(n11164), .Z(n11154) );
  AND U10523 ( .A(n2340), .B(n11165), .Z(n11164) );
  XOR U10524 ( .A(n11166), .B(n11167), .Z(n11152) );
  AND U10525 ( .A(n2344), .B(n11165), .Z(n11167) );
  XNOR U10526 ( .A(n11166), .B(n11163), .Z(n11165) );
  XOR U10527 ( .A(n11168), .B(n11169), .Z(n11163) );
  AND U10528 ( .A(n2347), .B(n11162), .Z(n11169) );
  XNOR U10529 ( .A(n11170), .B(n11160), .Z(n11162) );
  XOR U10530 ( .A(n11171), .B(n11172), .Z(n11160) );
  AND U10531 ( .A(n2351), .B(n11173), .Z(n11172) );
  XOR U10532 ( .A(p_input[1924]), .B(n11171), .Z(n11173) );
  XOR U10533 ( .A(n11174), .B(n11175), .Z(n11171) );
  AND U10534 ( .A(n2355), .B(n11176), .Z(n11175) );
  IV U10535 ( .A(n11168), .Z(n11170) );
  XOR U10536 ( .A(n11177), .B(n11178), .Z(n11168) );
  AND U10537 ( .A(n2359), .B(n11179), .Z(n11178) );
  XOR U10538 ( .A(n11180), .B(n11181), .Z(n11166) );
  AND U10539 ( .A(n2363), .B(n11179), .Z(n11181) );
  XNOR U10540 ( .A(n11180), .B(n11177), .Z(n11179) );
  XOR U10541 ( .A(n11182), .B(n11183), .Z(n11177) );
  AND U10542 ( .A(n2366), .B(n11176), .Z(n11183) );
  XNOR U10543 ( .A(n11184), .B(n11174), .Z(n11176) );
  XOR U10544 ( .A(n11185), .B(n11186), .Z(n11174) );
  AND U10545 ( .A(n2370), .B(n11187), .Z(n11186) );
  XOR U10546 ( .A(p_input[1940]), .B(n11185), .Z(n11187) );
  XOR U10547 ( .A(n11188), .B(n11189), .Z(n11185) );
  AND U10548 ( .A(n2374), .B(n11190), .Z(n11189) );
  IV U10549 ( .A(n11182), .Z(n11184) );
  XOR U10550 ( .A(n11191), .B(n11192), .Z(n11182) );
  AND U10551 ( .A(n2378), .B(n11193), .Z(n11192) );
  XOR U10552 ( .A(n11194), .B(n11195), .Z(n11180) );
  AND U10553 ( .A(n2382), .B(n11193), .Z(n11195) );
  XNOR U10554 ( .A(n11194), .B(n11191), .Z(n11193) );
  XOR U10555 ( .A(n11196), .B(n11197), .Z(n11191) );
  AND U10556 ( .A(n2385), .B(n11190), .Z(n11197) );
  XNOR U10557 ( .A(n11198), .B(n11188), .Z(n11190) );
  XOR U10558 ( .A(n11199), .B(n11200), .Z(n11188) );
  AND U10559 ( .A(n2389), .B(n11201), .Z(n11200) );
  XOR U10560 ( .A(p_input[1956]), .B(n11199), .Z(n11201) );
  XOR U10561 ( .A(n11202), .B(n11203), .Z(n11199) );
  AND U10562 ( .A(n2393), .B(n11204), .Z(n11203) );
  IV U10563 ( .A(n11196), .Z(n11198) );
  XOR U10564 ( .A(n11205), .B(n11206), .Z(n11196) );
  AND U10565 ( .A(n2397), .B(n11207), .Z(n11206) );
  XOR U10566 ( .A(n11208), .B(n11209), .Z(n11194) );
  AND U10567 ( .A(n2401), .B(n11207), .Z(n11209) );
  XNOR U10568 ( .A(n11208), .B(n11205), .Z(n11207) );
  XOR U10569 ( .A(n11210), .B(n11211), .Z(n11205) );
  AND U10570 ( .A(n2404), .B(n11204), .Z(n11211) );
  XNOR U10571 ( .A(n11212), .B(n11202), .Z(n11204) );
  XOR U10572 ( .A(n11213), .B(n11214), .Z(n11202) );
  AND U10573 ( .A(n2408), .B(n11215), .Z(n11214) );
  XOR U10574 ( .A(p_input[1972]), .B(n11213), .Z(n11215) );
  XOR U10575 ( .A(n11216), .B(n11217), .Z(n11213) );
  AND U10576 ( .A(n2412), .B(n11218), .Z(n11217) );
  IV U10577 ( .A(n11210), .Z(n11212) );
  XOR U10578 ( .A(n11219), .B(n11220), .Z(n11210) );
  AND U10579 ( .A(n2416), .B(n11221), .Z(n11220) );
  XOR U10580 ( .A(n11222), .B(n11223), .Z(n11208) );
  AND U10581 ( .A(n2420), .B(n11221), .Z(n11223) );
  XNOR U10582 ( .A(n11222), .B(n11219), .Z(n11221) );
  XOR U10583 ( .A(n11224), .B(n11225), .Z(n11219) );
  AND U10584 ( .A(n2423), .B(n11218), .Z(n11225) );
  XNOR U10585 ( .A(n11226), .B(n11216), .Z(n11218) );
  XOR U10586 ( .A(n11227), .B(n11228), .Z(n11216) );
  AND U10587 ( .A(n2427), .B(n11229), .Z(n11228) );
  XOR U10588 ( .A(p_input[1988]), .B(n11227), .Z(n11229) );
  XOR U10589 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n11230), 
        .Z(n11227) );
  AND U10590 ( .A(n2430), .B(n11231), .Z(n11230) );
  IV U10591 ( .A(n11224), .Z(n11226) );
  XOR U10592 ( .A(n11232), .B(n11233), .Z(n11224) );
  AND U10593 ( .A(n2434), .B(n11234), .Z(n11233) );
  XOR U10594 ( .A(n11235), .B(n11236), .Z(n11222) );
  AND U10595 ( .A(n2438), .B(n11234), .Z(n11236) );
  XNOR U10596 ( .A(n11235), .B(n11232), .Z(n11234) );
  XNOR U10597 ( .A(n11237), .B(n11238), .Z(n11232) );
  AND U10598 ( .A(n2441), .B(n11231), .Z(n11238) );
  XNOR U10599 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n11237), 
        .Z(n11231) );
  XNOR U10600 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n11239), 
        .Z(n11237) );
  AND U10601 ( .A(n2443), .B(n11240), .Z(n11239) );
  XNOR U10602 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n11241), .Z(n11235) );
  AND U10603 ( .A(n2446), .B(n11240), .Z(n11241) );
  XOR U10604 ( .A(n11242), .B(n11243), .Z(n11240) );
  IV U10605 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n11243) );
  IV U10606 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n11242) );
  XOR U10607 ( .A(n11244), .B(n11245), .Z(o[1]) );
  XOR U10608 ( .A(n29), .B(n11246), .Z(o[19]) );
  AND U10609 ( .A(n62), .B(n11247), .Z(n29) );
  XOR U10610 ( .A(n30), .B(n11246), .Z(n11247) );
  XOR U10611 ( .A(n11248), .B(n39), .Z(n11246) );
  AND U10612 ( .A(n65), .B(n11249), .Z(n39) );
  XNOR U10613 ( .A(n11250), .B(n40), .Z(n11249) );
  XOR U10614 ( .A(n11251), .B(n11252), .Z(n40) );
  AND U10615 ( .A(n70), .B(n11253), .Z(n11252) );
  XOR U10616 ( .A(p_input[3]), .B(n11251), .Z(n11253) );
  XOR U10617 ( .A(n11254), .B(n11255), .Z(n11251) );
  AND U10618 ( .A(n74), .B(n11256), .Z(n11255) );
  IV U10619 ( .A(n11248), .Z(n11250) );
  XOR U10620 ( .A(n11257), .B(n11258), .Z(n11248) );
  AND U10621 ( .A(n78), .B(n11259), .Z(n11258) );
  XOR U10622 ( .A(n11260), .B(n11261), .Z(n30) );
  AND U10623 ( .A(n82), .B(n11259), .Z(n11261) );
  XNOR U10624 ( .A(n11262), .B(n11257), .Z(n11259) );
  XOR U10625 ( .A(n11263), .B(n11264), .Z(n11257) );
  AND U10626 ( .A(n86), .B(n11256), .Z(n11264) );
  XNOR U10627 ( .A(n11265), .B(n11254), .Z(n11256) );
  XOR U10628 ( .A(n11266), .B(n11267), .Z(n11254) );
  AND U10629 ( .A(n90), .B(n11268), .Z(n11267) );
  XOR U10630 ( .A(p_input[19]), .B(n11266), .Z(n11268) );
  XOR U10631 ( .A(n11269), .B(n11270), .Z(n11266) );
  AND U10632 ( .A(n94), .B(n11271), .Z(n11270) );
  IV U10633 ( .A(n11263), .Z(n11265) );
  XOR U10634 ( .A(n11272), .B(n11273), .Z(n11263) );
  AND U10635 ( .A(n98), .B(n11274), .Z(n11273) );
  IV U10636 ( .A(n11260), .Z(n11262) );
  XNOR U10637 ( .A(n11275), .B(n11276), .Z(n11260) );
  AND U10638 ( .A(n102), .B(n11274), .Z(n11276) );
  XNOR U10639 ( .A(n11275), .B(n11272), .Z(n11274) );
  XOR U10640 ( .A(n11277), .B(n11278), .Z(n11272) );
  AND U10641 ( .A(n105), .B(n11271), .Z(n11278) );
  XNOR U10642 ( .A(n11279), .B(n11269), .Z(n11271) );
  XOR U10643 ( .A(n11280), .B(n11281), .Z(n11269) );
  AND U10644 ( .A(n109), .B(n11282), .Z(n11281) );
  XOR U10645 ( .A(p_input[35]), .B(n11280), .Z(n11282) );
  XOR U10646 ( .A(n11283), .B(n11284), .Z(n11280) );
  AND U10647 ( .A(n113), .B(n11285), .Z(n11284) );
  IV U10648 ( .A(n11277), .Z(n11279) );
  XOR U10649 ( .A(n11286), .B(n11287), .Z(n11277) );
  AND U10650 ( .A(n117), .B(n11288), .Z(n11287) );
  XOR U10651 ( .A(n11289), .B(n11290), .Z(n11275) );
  AND U10652 ( .A(n121), .B(n11288), .Z(n11290) );
  XNOR U10653 ( .A(n11289), .B(n11286), .Z(n11288) );
  XOR U10654 ( .A(n11291), .B(n11292), .Z(n11286) );
  AND U10655 ( .A(n124), .B(n11285), .Z(n11292) );
  XNOR U10656 ( .A(n11293), .B(n11283), .Z(n11285) );
  XOR U10657 ( .A(n11294), .B(n11295), .Z(n11283) );
  AND U10658 ( .A(n128), .B(n11296), .Z(n11295) );
  XOR U10659 ( .A(p_input[51]), .B(n11294), .Z(n11296) );
  XOR U10660 ( .A(n11297), .B(n11298), .Z(n11294) );
  AND U10661 ( .A(n132), .B(n11299), .Z(n11298) );
  IV U10662 ( .A(n11291), .Z(n11293) );
  XOR U10663 ( .A(n11300), .B(n11301), .Z(n11291) );
  AND U10664 ( .A(n136), .B(n11302), .Z(n11301) );
  XOR U10665 ( .A(n11303), .B(n11304), .Z(n11289) );
  AND U10666 ( .A(n140), .B(n11302), .Z(n11304) );
  XNOR U10667 ( .A(n11303), .B(n11300), .Z(n11302) );
  XOR U10668 ( .A(n11305), .B(n11306), .Z(n11300) );
  AND U10669 ( .A(n143), .B(n11299), .Z(n11306) );
  XNOR U10670 ( .A(n11307), .B(n11297), .Z(n11299) );
  XOR U10671 ( .A(n11308), .B(n11309), .Z(n11297) );
  AND U10672 ( .A(n147), .B(n11310), .Z(n11309) );
  XOR U10673 ( .A(p_input[67]), .B(n11308), .Z(n11310) );
  XOR U10674 ( .A(n11311), .B(n11312), .Z(n11308) );
  AND U10675 ( .A(n151), .B(n11313), .Z(n11312) );
  IV U10676 ( .A(n11305), .Z(n11307) );
  XOR U10677 ( .A(n11314), .B(n11315), .Z(n11305) );
  AND U10678 ( .A(n155), .B(n11316), .Z(n11315) );
  XOR U10679 ( .A(n11317), .B(n11318), .Z(n11303) );
  AND U10680 ( .A(n159), .B(n11316), .Z(n11318) );
  XNOR U10681 ( .A(n11317), .B(n11314), .Z(n11316) );
  XOR U10682 ( .A(n11319), .B(n11320), .Z(n11314) );
  AND U10683 ( .A(n162), .B(n11313), .Z(n11320) );
  XNOR U10684 ( .A(n11321), .B(n11311), .Z(n11313) );
  XOR U10685 ( .A(n11322), .B(n11323), .Z(n11311) );
  AND U10686 ( .A(n166), .B(n11324), .Z(n11323) );
  XOR U10687 ( .A(p_input[83]), .B(n11322), .Z(n11324) );
  XOR U10688 ( .A(n11325), .B(n11326), .Z(n11322) );
  AND U10689 ( .A(n170), .B(n11327), .Z(n11326) );
  IV U10690 ( .A(n11319), .Z(n11321) );
  XOR U10691 ( .A(n11328), .B(n11329), .Z(n11319) );
  AND U10692 ( .A(n174), .B(n11330), .Z(n11329) );
  XOR U10693 ( .A(n11331), .B(n11332), .Z(n11317) );
  AND U10694 ( .A(n178), .B(n11330), .Z(n11332) );
  XNOR U10695 ( .A(n11331), .B(n11328), .Z(n11330) );
  XOR U10696 ( .A(n11333), .B(n11334), .Z(n11328) );
  AND U10697 ( .A(n181), .B(n11327), .Z(n11334) );
  XNOR U10698 ( .A(n11335), .B(n11325), .Z(n11327) );
  XOR U10699 ( .A(n11336), .B(n11337), .Z(n11325) );
  AND U10700 ( .A(n185), .B(n11338), .Z(n11337) );
  XOR U10701 ( .A(p_input[99]), .B(n11336), .Z(n11338) );
  XOR U10702 ( .A(n11339), .B(n11340), .Z(n11336) );
  AND U10703 ( .A(n189), .B(n11341), .Z(n11340) );
  IV U10704 ( .A(n11333), .Z(n11335) );
  XOR U10705 ( .A(n11342), .B(n11343), .Z(n11333) );
  AND U10706 ( .A(n193), .B(n11344), .Z(n11343) );
  XOR U10707 ( .A(n11345), .B(n11346), .Z(n11331) );
  AND U10708 ( .A(n197), .B(n11344), .Z(n11346) );
  XNOR U10709 ( .A(n11345), .B(n11342), .Z(n11344) );
  XOR U10710 ( .A(n11347), .B(n11348), .Z(n11342) );
  AND U10711 ( .A(n200), .B(n11341), .Z(n11348) );
  XNOR U10712 ( .A(n11349), .B(n11339), .Z(n11341) );
  XOR U10713 ( .A(n11350), .B(n11351), .Z(n11339) );
  AND U10714 ( .A(n204), .B(n11352), .Z(n11351) );
  XOR U10715 ( .A(p_input[115]), .B(n11350), .Z(n11352) );
  XOR U10716 ( .A(n11353), .B(n11354), .Z(n11350) );
  AND U10717 ( .A(n208), .B(n11355), .Z(n11354) );
  IV U10718 ( .A(n11347), .Z(n11349) );
  XOR U10719 ( .A(n11356), .B(n11357), .Z(n11347) );
  AND U10720 ( .A(n212), .B(n11358), .Z(n11357) );
  XOR U10721 ( .A(n11359), .B(n11360), .Z(n11345) );
  AND U10722 ( .A(n216), .B(n11358), .Z(n11360) );
  XNOR U10723 ( .A(n11359), .B(n11356), .Z(n11358) );
  XOR U10724 ( .A(n11361), .B(n11362), .Z(n11356) );
  AND U10725 ( .A(n219), .B(n11355), .Z(n11362) );
  XNOR U10726 ( .A(n11363), .B(n11353), .Z(n11355) );
  XOR U10727 ( .A(n11364), .B(n11365), .Z(n11353) );
  AND U10728 ( .A(n223), .B(n11366), .Z(n11365) );
  XOR U10729 ( .A(p_input[131]), .B(n11364), .Z(n11366) );
  XOR U10730 ( .A(n11367), .B(n11368), .Z(n11364) );
  AND U10731 ( .A(n227), .B(n11369), .Z(n11368) );
  IV U10732 ( .A(n11361), .Z(n11363) );
  XOR U10733 ( .A(n11370), .B(n11371), .Z(n11361) );
  AND U10734 ( .A(n231), .B(n11372), .Z(n11371) );
  XOR U10735 ( .A(n11373), .B(n11374), .Z(n11359) );
  AND U10736 ( .A(n235), .B(n11372), .Z(n11374) );
  XNOR U10737 ( .A(n11373), .B(n11370), .Z(n11372) );
  XOR U10738 ( .A(n11375), .B(n11376), .Z(n11370) );
  AND U10739 ( .A(n238), .B(n11369), .Z(n11376) );
  XNOR U10740 ( .A(n11377), .B(n11367), .Z(n11369) );
  XOR U10741 ( .A(n11378), .B(n11379), .Z(n11367) );
  AND U10742 ( .A(n242), .B(n11380), .Z(n11379) );
  XOR U10743 ( .A(p_input[147]), .B(n11378), .Z(n11380) );
  XOR U10744 ( .A(n11381), .B(n11382), .Z(n11378) );
  AND U10745 ( .A(n246), .B(n11383), .Z(n11382) );
  IV U10746 ( .A(n11375), .Z(n11377) );
  XOR U10747 ( .A(n11384), .B(n11385), .Z(n11375) );
  AND U10748 ( .A(n250), .B(n11386), .Z(n11385) );
  XOR U10749 ( .A(n11387), .B(n11388), .Z(n11373) );
  AND U10750 ( .A(n254), .B(n11386), .Z(n11388) );
  XNOR U10751 ( .A(n11387), .B(n11384), .Z(n11386) );
  XOR U10752 ( .A(n11389), .B(n11390), .Z(n11384) );
  AND U10753 ( .A(n257), .B(n11383), .Z(n11390) );
  XNOR U10754 ( .A(n11391), .B(n11381), .Z(n11383) );
  XOR U10755 ( .A(n11392), .B(n11393), .Z(n11381) );
  AND U10756 ( .A(n261), .B(n11394), .Z(n11393) );
  XOR U10757 ( .A(p_input[163]), .B(n11392), .Z(n11394) );
  XOR U10758 ( .A(n11395), .B(n11396), .Z(n11392) );
  AND U10759 ( .A(n265), .B(n11397), .Z(n11396) );
  IV U10760 ( .A(n11389), .Z(n11391) );
  XOR U10761 ( .A(n11398), .B(n11399), .Z(n11389) );
  AND U10762 ( .A(n269), .B(n11400), .Z(n11399) );
  XOR U10763 ( .A(n11401), .B(n11402), .Z(n11387) );
  AND U10764 ( .A(n273), .B(n11400), .Z(n11402) );
  XNOR U10765 ( .A(n11401), .B(n11398), .Z(n11400) );
  XOR U10766 ( .A(n11403), .B(n11404), .Z(n11398) );
  AND U10767 ( .A(n276), .B(n11397), .Z(n11404) );
  XNOR U10768 ( .A(n11405), .B(n11395), .Z(n11397) );
  XOR U10769 ( .A(n11406), .B(n11407), .Z(n11395) );
  AND U10770 ( .A(n280), .B(n11408), .Z(n11407) );
  XOR U10771 ( .A(p_input[179]), .B(n11406), .Z(n11408) );
  XOR U10772 ( .A(n11409), .B(n11410), .Z(n11406) );
  AND U10773 ( .A(n284), .B(n11411), .Z(n11410) );
  IV U10774 ( .A(n11403), .Z(n11405) );
  XOR U10775 ( .A(n11412), .B(n11413), .Z(n11403) );
  AND U10776 ( .A(n288), .B(n11414), .Z(n11413) );
  XOR U10777 ( .A(n11415), .B(n11416), .Z(n11401) );
  AND U10778 ( .A(n292), .B(n11414), .Z(n11416) );
  XNOR U10779 ( .A(n11415), .B(n11412), .Z(n11414) );
  XOR U10780 ( .A(n11417), .B(n11418), .Z(n11412) );
  AND U10781 ( .A(n295), .B(n11411), .Z(n11418) );
  XNOR U10782 ( .A(n11419), .B(n11409), .Z(n11411) );
  XOR U10783 ( .A(n11420), .B(n11421), .Z(n11409) );
  AND U10784 ( .A(n299), .B(n11422), .Z(n11421) );
  XOR U10785 ( .A(p_input[195]), .B(n11420), .Z(n11422) );
  XOR U10786 ( .A(n11423), .B(n11424), .Z(n11420) );
  AND U10787 ( .A(n303), .B(n11425), .Z(n11424) );
  IV U10788 ( .A(n11417), .Z(n11419) );
  XOR U10789 ( .A(n11426), .B(n11427), .Z(n11417) );
  AND U10790 ( .A(n307), .B(n11428), .Z(n11427) );
  XOR U10791 ( .A(n11429), .B(n11430), .Z(n11415) );
  AND U10792 ( .A(n311), .B(n11428), .Z(n11430) );
  XNOR U10793 ( .A(n11429), .B(n11426), .Z(n11428) );
  XOR U10794 ( .A(n11431), .B(n11432), .Z(n11426) );
  AND U10795 ( .A(n314), .B(n11425), .Z(n11432) );
  XNOR U10796 ( .A(n11433), .B(n11423), .Z(n11425) );
  XOR U10797 ( .A(n11434), .B(n11435), .Z(n11423) );
  AND U10798 ( .A(n318), .B(n11436), .Z(n11435) );
  XOR U10799 ( .A(p_input[211]), .B(n11434), .Z(n11436) );
  XOR U10800 ( .A(n11437), .B(n11438), .Z(n11434) );
  AND U10801 ( .A(n322), .B(n11439), .Z(n11438) );
  IV U10802 ( .A(n11431), .Z(n11433) );
  XOR U10803 ( .A(n11440), .B(n11441), .Z(n11431) );
  AND U10804 ( .A(n326), .B(n11442), .Z(n11441) );
  XOR U10805 ( .A(n11443), .B(n11444), .Z(n11429) );
  AND U10806 ( .A(n330), .B(n11442), .Z(n11444) );
  XNOR U10807 ( .A(n11443), .B(n11440), .Z(n11442) );
  XOR U10808 ( .A(n11445), .B(n11446), .Z(n11440) );
  AND U10809 ( .A(n333), .B(n11439), .Z(n11446) );
  XNOR U10810 ( .A(n11447), .B(n11437), .Z(n11439) );
  XOR U10811 ( .A(n11448), .B(n11449), .Z(n11437) );
  AND U10812 ( .A(n337), .B(n11450), .Z(n11449) );
  XOR U10813 ( .A(p_input[227]), .B(n11448), .Z(n11450) );
  XOR U10814 ( .A(n11451), .B(n11452), .Z(n11448) );
  AND U10815 ( .A(n341), .B(n11453), .Z(n11452) );
  IV U10816 ( .A(n11445), .Z(n11447) );
  XOR U10817 ( .A(n11454), .B(n11455), .Z(n11445) );
  AND U10818 ( .A(n345), .B(n11456), .Z(n11455) );
  XOR U10819 ( .A(n11457), .B(n11458), .Z(n11443) );
  AND U10820 ( .A(n349), .B(n11456), .Z(n11458) );
  XNOR U10821 ( .A(n11457), .B(n11454), .Z(n11456) );
  XOR U10822 ( .A(n11459), .B(n11460), .Z(n11454) );
  AND U10823 ( .A(n352), .B(n11453), .Z(n11460) );
  XNOR U10824 ( .A(n11461), .B(n11451), .Z(n11453) );
  XOR U10825 ( .A(n11462), .B(n11463), .Z(n11451) );
  AND U10826 ( .A(n356), .B(n11464), .Z(n11463) );
  XOR U10827 ( .A(p_input[243]), .B(n11462), .Z(n11464) );
  XOR U10828 ( .A(n11465), .B(n11466), .Z(n11462) );
  AND U10829 ( .A(n360), .B(n11467), .Z(n11466) );
  IV U10830 ( .A(n11459), .Z(n11461) );
  XOR U10831 ( .A(n11468), .B(n11469), .Z(n11459) );
  AND U10832 ( .A(n364), .B(n11470), .Z(n11469) );
  XOR U10833 ( .A(n11471), .B(n11472), .Z(n11457) );
  AND U10834 ( .A(n368), .B(n11470), .Z(n11472) );
  XNOR U10835 ( .A(n11471), .B(n11468), .Z(n11470) );
  XOR U10836 ( .A(n11473), .B(n11474), .Z(n11468) );
  AND U10837 ( .A(n371), .B(n11467), .Z(n11474) );
  XNOR U10838 ( .A(n11475), .B(n11465), .Z(n11467) );
  XOR U10839 ( .A(n11476), .B(n11477), .Z(n11465) );
  AND U10840 ( .A(n375), .B(n11478), .Z(n11477) );
  XOR U10841 ( .A(p_input[259]), .B(n11476), .Z(n11478) );
  XOR U10842 ( .A(n11479), .B(n11480), .Z(n11476) );
  AND U10843 ( .A(n379), .B(n11481), .Z(n11480) );
  IV U10844 ( .A(n11473), .Z(n11475) );
  XOR U10845 ( .A(n11482), .B(n11483), .Z(n11473) );
  AND U10846 ( .A(n383), .B(n11484), .Z(n11483) );
  XOR U10847 ( .A(n11485), .B(n11486), .Z(n11471) );
  AND U10848 ( .A(n387), .B(n11484), .Z(n11486) );
  XNOR U10849 ( .A(n11485), .B(n11482), .Z(n11484) );
  XOR U10850 ( .A(n11487), .B(n11488), .Z(n11482) );
  AND U10851 ( .A(n390), .B(n11481), .Z(n11488) );
  XNOR U10852 ( .A(n11489), .B(n11479), .Z(n11481) );
  XOR U10853 ( .A(n11490), .B(n11491), .Z(n11479) );
  AND U10854 ( .A(n394), .B(n11492), .Z(n11491) );
  XOR U10855 ( .A(p_input[275]), .B(n11490), .Z(n11492) );
  XOR U10856 ( .A(n11493), .B(n11494), .Z(n11490) );
  AND U10857 ( .A(n398), .B(n11495), .Z(n11494) );
  IV U10858 ( .A(n11487), .Z(n11489) );
  XOR U10859 ( .A(n11496), .B(n11497), .Z(n11487) );
  AND U10860 ( .A(n402), .B(n11498), .Z(n11497) );
  XOR U10861 ( .A(n11499), .B(n11500), .Z(n11485) );
  AND U10862 ( .A(n406), .B(n11498), .Z(n11500) );
  XNOR U10863 ( .A(n11499), .B(n11496), .Z(n11498) );
  XOR U10864 ( .A(n11501), .B(n11502), .Z(n11496) );
  AND U10865 ( .A(n409), .B(n11495), .Z(n11502) );
  XNOR U10866 ( .A(n11503), .B(n11493), .Z(n11495) );
  XOR U10867 ( .A(n11504), .B(n11505), .Z(n11493) );
  AND U10868 ( .A(n413), .B(n11506), .Z(n11505) );
  XOR U10869 ( .A(p_input[291]), .B(n11504), .Z(n11506) );
  XOR U10870 ( .A(n11507), .B(n11508), .Z(n11504) );
  AND U10871 ( .A(n417), .B(n11509), .Z(n11508) );
  IV U10872 ( .A(n11501), .Z(n11503) );
  XOR U10873 ( .A(n11510), .B(n11511), .Z(n11501) );
  AND U10874 ( .A(n421), .B(n11512), .Z(n11511) );
  XOR U10875 ( .A(n11513), .B(n11514), .Z(n11499) );
  AND U10876 ( .A(n425), .B(n11512), .Z(n11514) );
  XNOR U10877 ( .A(n11513), .B(n11510), .Z(n11512) );
  XOR U10878 ( .A(n11515), .B(n11516), .Z(n11510) );
  AND U10879 ( .A(n428), .B(n11509), .Z(n11516) );
  XNOR U10880 ( .A(n11517), .B(n11507), .Z(n11509) );
  XOR U10881 ( .A(n11518), .B(n11519), .Z(n11507) );
  AND U10882 ( .A(n432), .B(n11520), .Z(n11519) );
  XOR U10883 ( .A(p_input[307]), .B(n11518), .Z(n11520) );
  XOR U10884 ( .A(n11521), .B(n11522), .Z(n11518) );
  AND U10885 ( .A(n436), .B(n11523), .Z(n11522) );
  IV U10886 ( .A(n11515), .Z(n11517) );
  XOR U10887 ( .A(n11524), .B(n11525), .Z(n11515) );
  AND U10888 ( .A(n440), .B(n11526), .Z(n11525) );
  XOR U10889 ( .A(n11527), .B(n11528), .Z(n11513) );
  AND U10890 ( .A(n444), .B(n11526), .Z(n11528) );
  XNOR U10891 ( .A(n11527), .B(n11524), .Z(n11526) );
  XOR U10892 ( .A(n11529), .B(n11530), .Z(n11524) );
  AND U10893 ( .A(n447), .B(n11523), .Z(n11530) );
  XNOR U10894 ( .A(n11531), .B(n11521), .Z(n11523) );
  XOR U10895 ( .A(n11532), .B(n11533), .Z(n11521) );
  AND U10896 ( .A(n451), .B(n11534), .Z(n11533) );
  XOR U10897 ( .A(p_input[323]), .B(n11532), .Z(n11534) );
  XOR U10898 ( .A(n11535), .B(n11536), .Z(n11532) );
  AND U10899 ( .A(n455), .B(n11537), .Z(n11536) );
  IV U10900 ( .A(n11529), .Z(n11531) );
  XOR U10901 ( .A(n11538), .B(n11539), .Z(n11529) );
  AND U10902 ( .A(n459), .B(n11540), .Z(n11539) );
  XOR U10903 ( .A(n11541), .B(n11542), .Z(n11527) );
  AND U10904 ( .A(n463), .B(n11540), .Z(n11542) );
  XNOR U10905 ( .A(n11541), .B(n11538), .Z(n11540) );
  XOR U10906 ( .A(n11543), .B(n11544), .Z(n11538) );
  AND U10907 ( .A(n466), .B(n11537), .Z(n11544) );
  XNOR U10908 ( .A(n11545), .B(n11535), .Z(n11537) );
  XOR U10909 ( .A(n11546), .B(n11547), .Z(n11535) );
  AND U10910 ( .A(n470), .B(n11548), .Z(n11547) );
  XOR U10911 ( .A(p_input[339]), .B(n11546), .Z(n11548) );
  XOR U10912 ( .A(n11549), .B(n11550), .Z(n11546) );
  AND U10913 ( .A(n474), .B(n11551), .Z(n11550) );
  IV U10914 ( .A(n11543), .Z(n11545) );
  XOR U10915 ( .A(n11552), .B(n11553), .Z(n11543) );
  AND U10916 ( .A(n478), .B(n11554), .Z(n11553) );
  XOR U10917 ( .A(n11555), .B(n11556), .Z(n11541) );
  AND U10918 ( .A(n482), .B(n11554), .Z(n11556) );
  XNOR U10919 ( .A(n11555), .B(n11552), .Z(n11554) );
  XOR U10920 ( .A(n11557), .B(n11558), .Z(n11552) );
  AND U10921 ( .A(n485), .B(n11551), .Z(n11558) );
  XNOR U10922 ( .A(n11559), .B(n11549), .Z(n11551) );
  XOR U10923 ( .A(n11560), .B(n11561), .Z(n11549) );
  AND U10924 ( .A(n489), .B(n11562), .Z(n11561) );
  XOR U10925 ( .A(p_input[355]), .B(n11560), .Z(n11562) );
  XOR U10926 ( .A(n11563), .B(n11564), .Z(n11560) );
  AND U10927 ( .A(n493), .B(n11565), .Z(n11564) );
  IV U10928 ( .A(n11557), .Z(n11559) );
  XOR U10929 ( .A(n11566), .B(n11567), .Z(n11557) );
  AND U10930 ( .A(n497), .B(n11568), .Z(n11567) );
  XOR U10931 ( .A(n11569), .B(n11570), .Z(n11555) );
  AND U10932 ( .A(n501), .B(n11568), .Z(n11570) );
  XNOR U10933 ( .A(n11569), .B(n11566), .Z(n11568) );
  XOR U10934 ( .A(n11571), .B(n11572), .Z(n11566) );
  AND U10935 ( .A(n504), .B(n11565), .Z(n11572) );
  XNOR U10936 ( .A(n11573), .B(n11563), .Z(n11565) );
  XOR U10937 ( .A(n11574), .B(n11575), .Z(n11563) );
  AND U10938 ( .A(n508), .B(n11576), .Z(n11575) );
  XOR U10939 ( .A(p_input[371]), .B(n11574), .Z(n11576) );
  XOR U10940 ( .A(n11577), .B(n11578), .Z(n11574) );
  AND U10941 ( .A(n512), .B(n11579), .Z(n11578) );
  IV U10942 ( .A(n11571), .Z(n11573) );
  XOR U10943 ( .A(n11580), .B(n11581), .Z(n11571) );
  AND U10944 ( .A(n516), .B(n11582), .Z(n11581) );
  XOR U10945 ( .A(n11583), .B(n11584), .Z(n11569) );
  AND U10946 ( .A(n520), .B(n11582), .Z(n11584) );
  XNOR U10947 ( .A(n11583), .B(n11580), .Z(n11582) );
  XOR U10948 ( .A(n11585), .B(n11586), .Z(n11580) );
  AND U10949 ( .A(n523), .B(n11579), .Z(n11586) );
  XNOR U10950 ( .A(n11587), .B(n11577), .Z(n11579) );
  XOR U10951 ( .A(n11588), .B(n11589), .Z(n11577) );
  AND U10952 ( .A(n527), .B(n11590), .Z(n11589) );
  XOR U10953 ( .A(p_input[387]), .B(n11588), .Z(n11590) );
  XOR U10954 ( .A(n11591), .B(n11592), .Z(n11588) );
  AND U10955 ( .A(n531), .B(n11593), .Z(n11592) );
  IV U10956 ( .A(n11585), .Z(n11587) );
  XOR U10957 ( .A(n11594), .B(n11595), .Z(n11585) );
  AND U10958 ( .A(n535), .B(n11596), .Z(n11595) );
  XOR U10959 ( .A(n11597), .B(n11598), .Z(n11583) );
  AND U10960 ( .A(n539), .B(n11596), .Z(n11598) );
  XNOR U10961 ( .A(n11597), .B(n11594), .Z(n11596) );
  XOR U10962 ( .A(n11599), .B(n11600), .Z(n11594) );
  AND U10963 ( .A(n542), .B(n11593), .Z(n11600) );
  XNOR U10964 ( .A(n11601), .B(n11591), .Z(n11593) );
  XOR U10965 ( .A(n11602), .B(n11603), .Z(n11591) );
  AND U10966 ( .A(n546), .B(n11604), .Z(n11603) );
  XOR U10967 ( .A(p_input[403]), .B(n11602), .Z(n11604) );
  XOR U10968 ( .A(n11605), .B(n11606), .Z(n11602) );
  AND U10969 ( .A(n550), .B(n11607), .Z(n11606) );
  IV U10970 ( .A(n11599), .Z(n11601) );
  XOR U10971 ( .A(n11608), .B(n11609), .Z(n11599) );
  AND U10972 ( .A(n554), .B(n11610), .Z(n11609) );
  XOR U10973 ( .A(n11611), .B(n11612), .Z(n11597) );
  AND U10974 ( .A(n558), .B(n11610), .Z(n11612) );
  XNOR U10975 ( .A(n11611), .B(n11608), .Z(n11610) );
  XOR U10976 ( .A(n11613), .B(n11614), .Z(n11608) );
  AND U10977 ( .A(n561), .B(n11607), .Z(n11614) );
  XNOR U10978 ( .A(n11615), .B(n11605), .Z(n11607) );
  XOR U10979 ( .A(n11616), .B(n11617), .Z(n11605) );
  AND U10980 ( .A(n565), .B(n11618), .Z(n11617) );
  XOR U10981 ( .A(p_input[419]), .B(n11616), .Z(n11618) );
  XOR U10982 ( .A(n11619), .B(n11620), .Z(n11616) );
  AND U10983 ( .A(n569), .B(n11621), .Z(n11620) );
  IV U10984 ( .A(n11613), .Z(n11615) );
  XOR U10985 ( .A(n11622), .B(n11623), .Z(n11613) );
  AND U10986 ( .A(n573), .B(n11624), .Z(n11623) );
  XOR U10987 ( .A(n11625), .B(n11626), .Z(n11611) );
  AND U10988 ( .A(n577), .B(n11624), .Z(n11626) );
  XNOR U10989 ( .A(n11625), .B(n11622), .Z(n11624) );
  XOR U10990 ( .A(n11627), .B(n11628), .Z(n11622) );
  AND U10991 ( .A(n580), .B(n11621), .Z(n11628) );
  XNOR U10992 ( .A(n11629), .B(n11619), .Z(n11621) );
  XOR U10993 ( .A(n11630), .B(n11631), .Z(n11619) );
  AND U10994 ( .A(n584), .B(n11632), .Z(n11631) );
  XOR U10995 ( .A(p_input[435]), .B(n11630), .Z(n11632) );
  XOR U10996 ( .A(n11633), .B(n11634), .Z(n11630) );
  AND U10997 ( .A(n588), .B(n11635), .Z(n11634) );
  IV U10998 ( .A(n11627), .Z(n11629) );
  XOR U10999 ( .A(n11636), .B(n11637), .Z(n11627) );
  AND U11000 ( .A(n592), .B(n11638), .Z(n11637) );
  XOR U11001 ( .A(n11639), .B(n11640), .Z(n11625) );
  AND U11002 ( .A(n596), .B(n11638), .Z(n11640) );
  XNOR U11003 ( .A(n11639), .B(n11636), .Z(n11638) );
  XOR U11004 ( .A(n11641), .B(n11642), .Z(n11636) );
  AND U11005 ( .A(n599), .B(n11635), .Z(n11642) );
  XNOR U11006 ( .A(n11643), .B(n11633), .Z(n11635) );
  XOR U11007 ( .A(n11644), .B(n11645), .Z(n11633) );
  AND U11008 ( .A(n603), .B(n11646), .Z(n11645) );
  XOR U11009 ( .A(p_input[451]), .B(n11644), .Z(n11646) );
  XOR U11010 ( .A(n11647), .B(n11648), .Z(n11644) );
  AND U11011 ( .A(n607), .B(n11649), .Z(n11648) );
  IV U11012 ( .A(n11641), .Z(n11643) );
  XOR U11013 ( .A(n11650), .B(n11651), .Z(n11641) );
  AND U11014 ( .A(n611), .B(n11652), .Z(n11651) );
  XOR U11015 ( .A(n11653), .B(n11654), .Z(n11639) );
  AND U11016 ( .A(n615), .B(n11652), .Z(n11654) );
  XNOR U11017 ( .A(n11653), .B(n11650), .Z(n11652) );
  XOR U11018 ( .A(n11655), .B(n11656), .Z(n11650) );
  AND U11019 ( .A(n618), .B(n11649), .Z(n11656) );
  XNOR U11020 ( .A(n11657), .B(n11647), .Z(n11649) );
  XOR U11021 ( .A(n11658), .B(n11659), .Z(n11647) );
  AND U11022 ( .A(n622), .B(n11660), .Z(n11659) );
  XOR U11023 ( .A(p_input[467]), .B(n11658), .Z(n11660) );
  XOR U11024 ( .A(n11661), .B(n11662), .Z(n11658) );
  AND U11025 ( .A(n626), .B(n11663), .Z(n11662) );
  IV U11026 ( .A(n11655), .Z(n11657) );
  XOR U11027 ( .A(n11664), .B(n11665), .Z(n11655) );
  AND U11028 ( .A(n630), .B(n11666), .Z(n11665) );
  XOR U11029 ( .A(n11667), .B(n11668), .Z(n11653) );
  AND U11030 ( .A(n634), .B(n11666), .Z(n11668) );
  XNOR U11031 ( .A(n11667), .B(n11664), .Z(n11666) );
  XOR U11032 ( .A(n11669), .B(n11670), .Z(n11664) );
  AND U11033 ( .A(n637), .B(n11663), .Z(n11670) );
  XNOR U11034 ( .A(n11671), .B(n11661), .Z(n11663) );
  XOR U11035 ( .A(n11672), .B(n11673), .Z(n11661) );
  AND U11036 ( .A(n641), .B(n11674), .Z(n11673) );
  XOR U11037 ( .A(p_input[483]), .B(n11672), .Z(n11674) );
  XOR U11038 ( .A(n11675), .B(n11676), .Z(n11672) );
  AND U11039 ( .A(n645), .B(n11677), .Z(n11676) );
  IV U11040 ( .A(n11669), .Z(n11671) );
  XOR U11041 ( .A(n11678), .B(n11679), .Z(n11669) );
  AND U11042 ( .A(n649), .B(n11680), .Z(n11679) );
  XOR U11043 ( .A(n11681), .B(n11682), .Z(n11667) );
  AND U11044 ( .A(n653), .B(n11680), .Z(n11682) );
  XNOR U11045 ( .A(n11681), .B(n11678), .Z(n11680) );
  XOR U11046 ( .A(n11683), .B(n11684), .Z(n11678) );
  AND U11047 ( .A(n656), .B(n11677), .Z(n11684) );
  XNOR U11048 ( .A(n11685), .B(n11675), .Z(n11677) );
  XOR U11049 ( .A(n11686), .B(n11687), .Z(n11675) );
  AND U11050 ( .A(n660), .B(n11688), .Z(n11687) );
  XOR U11051 ( .A(p_input[499]), .B(n11686), .Z(n11688) );
  XOR U11052 ( .A(n11689), .B(n11690), .Z(n11686) );
  AND U11053 ( .A(n664), .B(n11691), .Z(n11690) );
  IV U11054 ( .A(n11683), .Z(n11685) );
  XOR U11055 ( .A(n11692), .B(n11693), .Z(n11683) );
  AND U11056 ( .A(n668), .B(n11694), .Z(n11693) );
  XOR U11057 ( .A(n11695), .B(n11696), .Z(n11681) );
  AND U11058 ( .A(n672), .B(n11694), .Z(n11696) );
  XNOR U11059 ( .A(n11695), .B(n11692), .Z(n11694) );
  XOR U11060 ( .A(n11697), .B(n11698), .Z(n11692) );
  AND U11061 ( .A(n675), .B(n11691), .Z(n11698) );
  XNOR U11062 ( .A(n11699), .B(n11689), .Z(n11691) );
  XOR U11063 ( .A(n11700), .B(n11701), .Z(n11689) );
  AND U11064 ( .A(n679), .B(n11702), .Z(n11701) );
  XOR U11065 ( .A(p_input[515]), .B(n11700), .Z(n11702) );
  XOR U11066 ( .A(n11703), .B(n11704), .Z(n11700) );
  AND U11067 ( .A(n683), .B(n11705), .Z(n11704) );
  IV U11068 ( .A(n11697), .Z(n11699) );
  XOR U11069 ( .A(n11706), .B(n11707), .Z(n11697) );
  AND U11070 ( .A(n687), .B(n11708), .Z(n11707) );
  XOR U11071 ( .A(n11709), .B(n11710), .Z(n11695) );
  AND U11072 ( .A(n691), .B(n11708), .Z(n11710) );
  XNOR U11073 ( .A(n11709), .B(n11706), .Z(n11708) );
  XOR U11074 ( .A(n11711), .B(n11712), .Z(n11706) );
  AND U11075 ( .A(n694), .B(n11705), .Z(n11712) );
  XNOR U11076 ( .A(n11713), .B(n11703), .Z(n11705) );
  XOR U11077 ( .A(n11714), .B(n11715), .Z(n11703) );
  AND U11078 ( .A(n698), .B(n11716), .Z(n11715) );
  XOR U11079 ( .A(p_input[531]), .B(n11714), .Z(n11716) );
  XOR U11080 ( .A(n11717), .B(n11718), .Z(n11714) );
  AND U11081 ( .A(n702), .B(n11719), .Z(n11718) );
  IV U11082 ( .A(n11711), .Z(n11713) );
  XOR U11083 ( .A(n11720), .B(n11721), .Z(n11711) );
  AND U11084 ( .A(n706), .B(n11722), .Z(n11721) );
  XOR U11085 ( .A(n11723), .B(n11724), .Z(n11709) );
  AND U11086 ( .A(n710), .B(n11722), .Z(n11724) );
  XNOR U11087 ( .A(n11723), .B(n11720), .Z(n11722) );
  XOR U11088 ( .A(n11725), .B(n11726), .Z(n11720) );
  AND U11089 ( .A(n713), .B(n11719), .Z(n11726) );
  XNOR U11090 ( .A(n11727), .B(n11717), .Z(n11719) );
  XOR U11091 ( .A(n11728), .B(n11729), .Z(n11717) );
  AND U11092 ( .A(n717), .B(n11730), .Z(n11729) );
  XOR U11093 ( .A(p_input[547]), .B(n11728), .Z(n11730) );
  XOR U11094 ( .A(n11731), .B(n11732), .Z(n11728) );
  AND U11095 ( .A(n721), .B(n11733), .Z(n11732) );
  IV U11096 ( .A(n11725), .Z(n11727) );
  XOR U11097 ( .A(n11734), .B(n11735), .Z(n11725) );
  AND U11098 ( .A(n725), .B(n11736), .Z(n11735) );
  XOR U11099 ( .A(n11737), .B(n11738), .Z(n11723) );
  AND U11100 ( .A(n729), .B(n11736), .Z(n11738) );
  XNOR U11101 ( .A(n11737), .B(n11734), .Z(n11736) );
  XOR U11102 ( .A(n11739), .B(n11740), .Z(n11734) );
  AND U11103 ( .A(n732), .B(n11733), .Z(n11740) );
  XNOR U11104 ( .A(n11741), .B(n11731), .Z(n11733) );
  XOR U11105 ( .A(n11742), .B(n11743), .Z(n11731) );
  AND U11106 ( .A(n736), .B(n11744), .Z(n11743) );
  XOR U11107 ( .A(p_input[563]), .B(n11742), .Z(n11744) );
  XOR U11108 ( .A(n11745), .B(n11746), .Z(n11742) );
  AND U11109 ( .A(n740), .B(n11747), .Z(n11746) );
  IV U11110 ( .A(n11739), .Z(n11741) );
  XOR U11111 ( .A(n11748), .B(n11749), .Z(n11739) );
  AND U11112 ( .A(n744), .B(n11750), .Z(n11749) );
  XOR U11113 ( .A(n11751), .B(n11752), .Z(n11737) );
  AND U11114 ( .A(n748), .B(n11750), .Z(n11752) );
  XNOR U11115 ( .A(n11751), .B(n11748), .Z(n11750) );
  XOR U11116 ( .A(n11753), .B(n11754), .Z(n11748) );
  AND U11117 ( .A(n751), .B(n11747), .Z(n11754) );
  XNOR U11118 ( .A(n11755), .B(n11745), .Z(n11747) );
  XOR U11119 ( .A(n11756), .B(n11757), .Z(n11745) );
  AND U11120 ( .A(n755), .B(n11758), .Z(n11757) );
  XOR U11121 ( .A(p_input[579]), .B(n11756), .Z(n11758) );
  XOR U11122 ( .A(n11759), .B(n11760), .Z(n11756) );
  AND U11123 ( .A(n759), .B(n11761), .Z(n11760) );
  IV U11124 ( .A(n11753), .Z(n11755) );
  XOR U11125 ( .A(n11762), .B(n11763), .Z(n11753) );
  AND U11126 ( .A(n763), .B(n11764), .Z(n11763) );
  XOR U11127 ( .A(n11765), .B(n11766), .Z(n11751) );
  AND U11128 ( .A(n767), .B(n11764), .Z(n11766) );
  XNOR U11129 ( .A(n11765), .B(n11762), .Z(n11764) );
  XOR U11130 ( .A(n11767), .B(n11768), .Z(n11762) );
  AND U11131 ( .A(n770), .B(n11761), .Z(n11768) );
  XNOR U11132 ( .A(n11769), .B(n11759), .Z(n11761) );
  XOR U11133 ( .A(n11770), .B(n11771), .Z(n11759) );
  AND U11134 ( .A(n774), .B(n11772), .Z(n11771) );
  XOR U11135 ( .A(p_input[595]), .B(n11770), .Z(n11772) );
  XOR U11136 ( .A(n11773), .B(n11774), .Z(n11770) );
  AND U11137 ( .A(n778), .B(n11775), .Z(n11774) );
  IV U11138 ( .A(n11767), .Z(n11769) );
  XOR U11139 ( .A(n11776), .B(n11777), .Z(n11767) );
  AND U11140 ( .A(n782), .B(n11778), .Z(n11777) );
  XOR U11141 ( .A(n11779), .B(n11780), .Z(n11765) );
  AND U11142 ( .A(n786), .B(n11778), .Z(n11780) );
  XNOR U11143 ( .A(n11779), .B(n11776), .Z(n11778) );
  XOR U11144 ( .A(n11781), .B(n11782), .Z(n11776) );
  AND U11145 ( .A(n789), .B(n11775), .Z(n11782) );
  XNOR U11146 ( .A(n11783), .B(n11773), .Z(n11775) );
  XOR U11147 ( .A(n11784), .B(n11785), .Z(n11773) );
  AND U11148 ( .A(n793), .B(n11786), .Z(n11785) );
  XOR U11149 ( .A(p_input[611]), .B(n11784), .Z(n11786) );
  XOR U11150 ( .A(n11787), .B(n11788), .Z(n11784) );
  AND U11151 ( .A(n797), .B(n11789), .Z(n11788) );
  IV U11152 ( .A(n11781), .Z(n11783) );
  XOR U11153 ( .A(n11790), .B(n11791), .Z(n11781) );
  AND U11154 ( .A(n801), .B(n11792), .Z(n11791) );
  XOR U11155 ( .A(n11793), .B(n11794), .Z(n11779) );
  AND U11156 ( .A(n805), .B(n11792), .Z(n11794) );
  XNOR U11157 ( .A(n11793), .B(n11790), .Z(n11792) );
  XOR U11158 ( .A(n11795), .B(n11796), .Z(n11790) );
  AND U11159 ( .A(n808), .B(n11789), .Z(n11796) );
  XNOR U11160 ( .A(n11797), .B(n11787), .Z(n11789) );
  XOR U11161 ( .A(n11798), .B(n11799), .Z(n11787) );
  AND U11162 ( .A(n812), .B(n11800), .Z(n11799) );
  XOR U11163 ( .A(p_input[627]), .B(n11798), .Z(n11800) );
  XOR U11164 ( .A(n11801), .B(n11802), .Z(n11798) );
  AND U11165 ( .A(n816), .B(n11803), .Z(n11802) );
  IV U11166 ( .A(n11795), .Z(n11797) );
  XOR U11167 ( .A(n11804), .B(n11805), .Z(n11795) );
  AND U11168 ( .A(n820), .B(n11806), .Z(n11805) );
  XOR U11169 ( .A(n11807), .B(n11808), .Z(n11793) );
  AND U11170 ( .A(n824), .B(n11806), .Z(n11808) );
  XNOR U11171 ( .A(n11807), .B(n11804), .Z(n11806) );
  XOR U11172 ( .A(n11809), .B(n11810), .Z(n11804) );
  AND U11173 ( .A(n827), .B(n11803), .Z(n11810) );
  XNOR U11174 ( .A(n11811), .B(n11801), .Z(n11803) );
  XOR U11175 ( .A(n11812), .B(n11813), .Z(n11801) );
  AND U11176 ( .A(n831), .B(n11814), .Z(n11813) );
  XOR U11177 ( .A(p_input[643]), .B(n11812), .Z(n11814) );
  XOR U11178 ( .A(n11815), .B(n11816), .Z(n11812) );
  AND U11179 ( .A(n835), .B(n11817), .Z(n11816) );
  IV U11180 ( .A(n11809), .Z(n11811) );
  XOR U11181 ( .A(n11818), .B(n11819), .Z(n11809) );
  AND U11182 ( .A(n839), .B(n11820), .Z(n11819) );
  XOR U11183 ( .A(n11821), .B(n11822), .Z(n11807) );
  AND U11184 ( .A(n843), .B(n11820), .Z(n11822) );
  XNOR U11185 ( .A(n11821), .B(n11818), .Z(n11820) );
  XOR U11186 ( .A(n11823), .B(n11824), .Z(n11818) );
  AND U11187 ( .A(n846), .B(n11817), .Z(n11824) );
  XNOR U11188 ( .A(n11825), .B(n11815), .Z(n11817) );
  XOR U11189 ( .A(n11826), .B(n11827), .Z(n11815) );
  AND U11190 ( .A(n850), .B(n11828), .Z(n11827) );
  XOR U11191 ( .A(p_input[659]), .B(n11826), .Z(n11828) );
  XOR U11192 ( .A(n11829), .B(n11830), .Z(n11826) );
  AND U11193 ( .A(n854), .B(n11831), .Z(n11830) );
  IV U11194 ( .A(n11823), .Z(n11825) );
  XOR U11195 ( .A(n11832), .B(n11833), .Z(n11823) );
  AND U11196 ( .A(n858), .B(n11834), .Z(n11833) );
  XOR U11197 ( .A(n11835), .B(n11836), .Z(n11821) );
  AND U11198 ( .A(n862), .B(n11834), .Z(n11836) );
  XNOR U11199 ( .A(n11835), .B(n11832), .Z(n11834) );
  XOR U11200 ( .A(n11837), .B(n11838), .Z(n11832) );
  AND U11201 ( .A(n865), .B(n11831), .Z(n11838) );
  XNOR U11202 ( .A(n11839), .B(n11829), .Z(n11831) );
  XOR U11203 ( .A(n11840), .B(n11841), .Z(n11829) );
  AND U11204 ( .A(n869), .B(n11842), .Z(n11841) );
  XOR U11205 ( .A(p_input[675]), .B(n11840), .Z(n11842) );
  XOR U11206 ( .A(n11843), .B(n11844), .Z(n11840) );
  AND U11207 ( .A(n873), .B(n11845), .Z(n11844) );
  IV U11208 ( .A(n11837), .Z(n11839) );
  XOR U11209 ( .A(n11846), .B(n11847), .Z(n11837) );
  AND U11210 ( .A(n877), .B(n11848), .Z(n11847) );
  XOR U11211 ( .A(n11849), .B(n11850), .Z(n11835) );
  AND U11212 ( .A(n881), .B(n11848), .Z(n11850) );
  XNOR U11213 ( .A(n11849), .B(n11846), .Z(n11848) );
  XOR U11214 ( .A(n11851), .B(n11852), .Z(n11846) );
  AND U11215 ( .A(n884), .B(n11845), .Z(n11852) );
  XNOR U11216 ( .A(n11853), .B(n11843), .Z(n11845) );
  XOR U11217 ( .A(n11854), .B(n11855), .Z(n11843) );
  AND U11218 ( .A(n888), .B(n11856), .Z(n11855) );
  XOR U11219 ( .A(p_input[691]), .B(n11854), .Z(n11856) );
  XOR U11220 ( .A(n11857), .B(n11858), .Z(n11854) );
  AND U11221 ( .A(n892), .B(n11859), .Z(n11858) );
  IV U11222 ( .A(n11851), .Z(n11853) );
  XOR U11223 ( .A(n11860), .B(n11861), .Z(n11851) );
  AND U11224 ( .A(n896), .B(n11862), .Z(n11861) );
  XOR U11225 ( .A(n11863), .B(n11864), .Z(n11849) );
  AND U11226 ( .A(n900), .B(n11862), .Z(n11864) );
  XNOR U11227 ( .A(n11863), .B(n11860), .Z(n11862) );
  XOR U11228 ( .A(n11865), .B(n11866), .Z(n11860) );
  AND U11229 ( .A(n903), .B(n11859), .Z(n11866) );
  XNOR U11230 ( .A(n11867), .B(n11857), .Z(n11859) );
  XOR U11231 ( .A(n11868), .B(n11869), .Z(n11857) );
  AND U11232 ( .A(n907), .B(n11870), .Z(n11869) );
  XOR U11233 ( .A(p_input[707]), .B(n11868), .Z(n11870) );
  XOR U11234 ( .A(n11871), .B(n11872), .Z(n11868) );
  AND U11235 ( .A(n911), .B(n11873), .Z(n11872) );
  IV U11236 ( .A(n11865), .Z(n11867) );
  XOR U11237 ( .A(n11874), .B(n11875), .Z(n11865) );
  AND U11238 ( .A(n915), .B(n11876), .Z(n11875) );
  XOR U11239 ( .A(n11877), .B(n11878), .Z(n11863) );
  AND U11240 ( .A(n919), .B(n11876), .Z(n11878) );
  XNOR U11241 ( .A(n11877), .B(n11874), .Z(n11876) );
  XOR U11242 ( .A(n11879), .B(n11880), .Z(n11874) );
  AND U11243 ( .A(n922), .B(n11873), .Z(n11880) );
  XNOR U11244 ( .A(n11881), .B(n11871), .Z(n11873) );
  XOR U11245 ( .A(n11882), .B(n11883), .Z(n11871) );
  AND U11246 ( .A(n926), .B(n11884), .Z(n11883) );
  XOR U11247 ( .A(p_input[723]), .B(n11882), .Z(n11884) );
  XOR U11248 ( .A(n11885), .B(n11886), .Z(n11882) );
  AND U11249 ( .A(n930), .B(n11887), .Z(n11886) );
  IV U11250 ( .A(n11879), .Z(n11881) );
  XOR U11251 ( .A(n11888), .B(n11889), .Z(n11879) );
  AND U11252 ( .A(n934), .B(n11890), .Z(n11889) );
  XOR U11253 ( .A(n11891), .B(n11892), .Z(n11877) );
  AND U11254 ( .A(n938), .B(n11890), .Z(n11892) );
  XNOR U11255 ( .A(n11891), .B(n11888), .Z(n11890) );
  XOR U11256 ( .A(n11893), .B(n11894), .Z(n11888) );
  AND U11257 ( .A(n941), .B(n11887), .Z(n11894) );
  XNOR U11258 ( .A(n11895), .B(n11885), .Z(n11887) );
  XOR U11259 ( .A(n11896), .B(n11897), .Z(n11885) );
  AND U11260 ( .A(n945), .B(n11898), .Z(n11897) );
  XOR U11261 ( .A(p_input[739]), .B(n11896), .Z(n11898) );
  XOR U11262 ( .A(n11899), .B(n11900), .Z(n11896) );
  AND U11263 ( .A(n949), .B(n11901), .Z(n11900) );
  IV U11264 ( .A(n11893), .Z(n11895) );
  XOR U11265 ( .A(n11902), .B(n11903), .Z(n11893) );
  AND U11266 ( .A(n953), .B(n11904), .Z(n11903) );
  XOR U11267 ( .A(n11905), .B(n11906), .Z(n11891) );
  AND U11268 ( .A(n957), .B(n11904), .Z(n11906) );
  XNOR U11269 ( .A(n11905), .B(n11902), .Z(n11904) );
  XOR U11270 ( .A(n11907), .B(n11908), .Z(n11902) );
  AND U11271 ( .A(n960), .B(n11901), .Z(n11908) );
  XNOR U11272 ( .A(n11909), .B(n11899), .Z(n11901) );
  XOR U11273 ( .A(n11910), .B(n11911), .Z(n11899) );
  AND U11274 ( .A(n964), .B(n11912), .Z(n11911) );
  XOR U11275 ( .A(p_input[755]), .B(n11910), .Z(n11912) );
  XOR U11276 ( .A(n11913), .B(n11914), .Z(n11910) );
  AND U11277 ( .A(n968), .B(n11915), .Z(n11914) );
  IV U11278 ( .A(n11907), .Z(n11909) );
  XOR U11279 ( .A(n11916), .B(n11917), .Z(n11907) );
  AND U11280 ( .A(n972), .B(n11918), .Z(n11917) );
  XOR U11281 ( .A(n11919), .B(n11920), .Z(n11905) );
  AND U11282 ( .A(n976), .B(n11918), .Z(n11920) );
  XNOR U11283 ( .A(n11919), .B(n11916), .Z(n11918) );
  XOR U11284 ( .A(n11921), .B(n11922), .Z(n11916) );
  AND U11285 ( .A(n979), .B(n11915), .Z(n11922) );
  XNOR U11286 ( .A(n11923), .B(n11913), .Z(n11915) );
  XOR U11287 ( .A(n11924), .B(n11925), .Z(n11913) );
  AND U11288 ( .A(n983), .B(n11926), .Z(n11925) );
  XOR U11289 ( .A(p_input[771]), .B(n11924), .Z(n11926) );
  XOR U11290 ( .A(n11927), .B(n11928), .Z(n11924) );
  AND U11291 ( .A(n987), .B(n11929), .Z(n11928) );
  IV U11292 ( .A(n11921), .Z(n11923) );
  XOR U11293 ( .A(n11930), .B(n11931), .Z(n11921) );
  AND U11294 ( .A(n991), .B(n11932), .Z(n11931) );
  XOR U11295 ( .A(n11933), .B(n11934), .Z(n11919) );
  AND U11296 ( .A(n995), .B(n11932), .Z(n11934) );
  XNOR U11297 ( .A(n11933), .B(n11930), .Z(n11932) );
  XOR U11298 ( .A(n11935), .B(n11936), .Z(n11930) );
  AND U11299 ( .A(n998), .B(n11929), .Z(n11936) );
  XNOR U11300 ( .A(n11937), .B(n11927), .Z(n11929) );
  XOR U11301 ( .A(n11938), .B(n11939), .Z(n11927) );
  AND U11302 ( .A(n1002), .B(n11940), .Z(n11939) );
  XOR U11303 ( .A(p_input[787]), .B(n11938), .Z(n11940) );
  XOR U11304 ( .A(n11941), .B(n11942), .Z(n11938) );
  AND U11305 ( .A(n1006), .B(n11943), .Z(n11942) );
  IV U11306 ( .A(n11935), .Z(n11937) );
  XOR U11307 ( .A(n11944), .B(n11945), .Z(n11935) );
  AND U11308 ( .A(n1010), .B(n11946), .Z(n11945) );
  XOR U11309 ( .A(n11947), .B(n11948), .Z(n11933) );
  AND U11310 ( .A(n1014), .B(n11946), .Z(n11948) );
  XNOR U11311 ( .A(n11947), .B(n11944), .Z(n11946) );
  XOR U11312 ( .A(n11949), .B(n11950), .Z(n11944) );
  AND U11313 ( .A(n1017), .B(n11943), .Z(n11950) );
  XNOR U11314 ( .A(n11951), .B(n11941), .Z(n11943) );
  XOR U11315 ( .A(n11952), .B(n11953), .Z(n11941) );
  AND U11316 ( .A(n1021), .B(n11954), .Z(n11953) );
  XOR U11317 ( .A(p_input[803]), .B(n11952), .Z(n11954) );
  XOR U11318 ( .A(n11955), .B(n11956), .Z(n11952) );
  AND U11319 ( .A(n1025), .B(n11957), .Z(n11956) );
  IV U11320 ( .A(n11949), .Z(n11951) );
  XOR U11321 ( .A(n11958), .B(n11959), .Z(n11949) );
  AND U11322 ( .A(n1029), .B(n11960), .Z(n11959) );
  XOR U11323 ( .A(n11961), .B(n11962), .Z(n11947) );
  AND U11324 ( .A(n1033), .B(n11960), .Z(n11962) );
  XNOR U11325 ( .A(n11961), .B(n11958), .Z(n11960) );
  XOR U11326 ( .A(n11963), .B(n11964), .Z(n11958) );
  AND U11327 ( .A(n1036), .B(n11957), .Z(n11964) );
  XNOR U11328 ( .A(n11965), .B(n11955), .Z(n11957) );
  XOR U11329 ( .A(n11966), .B(n11967), .Z(n11955) );
  AND U11330 ( .A(n1040), .B(n11968), .Z(n11967) );
  XOR U11331 ( .A(p_input[819]), .B(n11966), .Z(n11968) );
  XOR U11332 ( .A(n11969), .B(n11970), .Z(n11966) );
  AND U11333 ( .A(n1044), .B(n11971), .Z(n11970) );
  IV U11334 ( .A(n11963), .Z(n11965) );
  XOR U11335 ( .A(n11972), .B(n11973), .Z(n11963) );
  AND U11336 ( .A(n1048), .B(n11974), .Z(n11973) );
  XOR U11337 ( .A(n11975), .B(n11976), .Z(n11961) );
  AND U11338 ( .A(n1052), .B(n11974), .Z(n11976) );
  XNOR U11339 ( .A(n11975), .B(n11972), .Z(n11974) );
  XOR U11340 ( .A(n11977), .B(n11978), .Z(n11972) );
  AND U11341 ( .A(n1055), .B(n11971), .Z(n11978) );
  XNOR U11342 ( .A(n11979), .B(n11969), .Z(n11971) );
  XOR U11343 ( .A(n11980), .B(n11981), .Z(n11969) );
  AND U11344 ( .A(n1059), .B(n11982), .Z(n11981) );
  XOR U11345 ( .A(p_input[835]), .B(n11980), .Z(n11982) );
  XOR U11346 ( .A(n11983), .B(n11984), .Z(n11980) );
  AND U11347 ( .A(n1063), .B(n11985), .Z(n11984) );
  IV U11348 ( .A(n11977), .Z(n11979) );
  XOR U11349 ( .A(n11986), .B(n11987), .Z(n11977) );
  AND U11350 ( .A(n1067), .B(n11988), .Z(n11987) );
  XOR U11351 ( .A(n11989), .B(n11990), .Z(n11975) );
  AND U11352 ( .A(n1071), .B(n11988), .Z(n11990) );
  XNOR U11353 ( .A(n11989), .B(n11986), .Z(n11988) );
  XOR U11354 ( .A(n11991), .B(n11992), .Z(n11986) );
  AND U11355 ( .A(n1074), .B(n11985), .Z(n11992) );
  XNOR U11356 ( .A(n11993), .B(n11983), .Z(n11985) );
  XOR U11357 ( .A(n11994), .B(n11995), .Z(n11983) );
  AND U11358 ( .A(n1078), .B(n11996), .Z(n11995) );
  XOR U11359 ( .A(p_input[851]), .B(n11994), .Z(n11996) );
  XOR U11360 ( .A(n11997), .B(n11998), .Z(n11994) );
  AND U11361 ( .A(n1082), .B(n11999), .Z(n11998) );
  IV U11362 ( .A(n11991), .Z(n11993) );
  XOR U11363 ( .A(n12000), .B(n12001), .Z(n11991) );
  AND U11364 ( .A(n1086), .B(n12002), .Z(n12001) );
  XOR U11365 ( .A(n12003), .B(n12004), .Z(n11989) );
  AND U11366 ( .A(n1090), .B(n12002), .Z(n12004) );
  XNOR U11367 ( .A(n12003), .B(n12000), .Z(n12002) );
  XOR U11368 ( .A(n12005), .B(n12006), .Z(n12000) );
  AND U11369 ( .A(n1093), .B(n11999), .Z(n12006) );
  XNOR U11370 ( .A(n12007), .B(n11997), .Z(n11999) );
  XOR U11371 ( .A(n12008), .B(n12009), .Z(n11997) );
  AND U11372 ( .A(n1097), .B(n12010), .Z(n12009) );
  XOR U11373 ( .A(p_input[867]), .B(n12008), .Z(n12010) );
  XOR U11374 ( .A(n12011), .B(n12012), .Z(n12008) );
  AND U11375 ( .A(n1101), .B(n12013), .Z(n12012) );
  IV U11376 ( .A(n12005), .Z(n12007) );
  XOR U11377 ( .A(n12014), .B(n12015), .Z(n12005) );
  AND U11378 ( .A(n1105), .B(n12016), .Z(n12015) );
  XOR U11379 ( .A(n12017), .B(n12018), .Z(n12003) );
  AND U11380 ( .A(n1109), .B(n12016), .Z(n12018) );
  XNOR U11381 ( .A(n12017), .B(n12014), .Z(n12016) );
  XOR U11382 ( .A(n12019), .B(n12020), .Z(n12014) );
  AND U11383 ( .A(n1112), .B(n12013), .Z(n12020) );
  XNOR U11384 ( .A(n12021), .B(n12011), .Z(n12013) );
  XOR U11385 ( .A(n12022), .B(n12023), .Z(n12011) );
  AND U11386 ( .A(n1116), .B(n12024), .Z(n12023) );
  XOR U11387 ( .A(p_input[883]), .B(n12022), .Z(n12024) );
  XOR U11388 ( .A(n12025), .B(n12026), .Z(n12022) );
  AND U11389 ( .A(n1120), .B(n12027), .Z(n12026) );
  IV U11390 ( .A(n12019), .Z(n12021) );
  XOR U11391 ( .A(n12028), .B(n12029), .Z(n12019) );
  AND U11392 ( .A(n1124), .B(n12030), .Z(n12029) );
  XOR U11393 ( .A(n12031), .B(n12032), .Z(n12017) );
  AND U11394 ( .A(n1128), .B(n12030), .Z(n12032) );
  XNOR U11395 ( .A(n12031), .B(n12028), .Z(n12030) );
  XOR U11396 ( .A(n12033), .B(n12034), .Z(n12028) );
  AND U11397 ( .A(n1131), .B(n12027), .Z(n12034) );
  XNOR U11398 ( .A(n12035), .B(n12025), .Z(n12027) );
  XOR U11399 ( .A(n12036), .B(n12037), .Z(n12025) );
  AND U11400 ( .A(n1135), .B(n12038), .Z(n12037) );
  XOR U11401 ( .A(p_input[899]), .B(n12036), .Z(n12038) );
  XOR U11402 ( .A(n12039), .B(n12040), .Z(n12036) );
  AND U11403 ( .A(n1139), .B(n12041), .Z(n12040) );
  IV U11404 ( .A(n12033), .Z(n12035) );
  XOR U11405 ( .A(n12042), .B(n12043), .Z(n12033) );
  AND U11406 ( .A(n1143), .B(n12044), .Z(n12043) );
  XOR U11407 ( .A(n12045), .B(n12046), .Z(n12031) );
  AND U11408 ( .A(n1147), .B(n12044), .Z(n12046) );
  XNOR U11409 ( .A(n12045), .B(n12042), .Z(n12044) );
  XOR U11410 ( .A(n12047), .B(n12048), .Z(n12042) );
  AND U11411 ( .A(n1150), .B(n12041), .Z(n12048) );
  XNOR U11412 ( .A(n12049), .B(n12039), .Z(n12041) );
  XOR U11413 ( .A(n12050), .B(n12051), .Z(n12039) );
  AND U11414 ( .A(n1154), .B(n12052), .Z(n12051) );
  XOR U11415 ( .A(p_input[915]), .B(n12050), .Z(n12052) );
  XOR U11416 ( .A(n12053), .B(n12054), .Z(n12050) );
  AND U11417 ( .A(n1158), .B(n12055), .Z(n12054) );
  IV U11418 ( .A(n12047), .Z(n12049) );
  XOR U11419 ( .A(n12056), .B(n12057), .Z(n12047) );
  AND U11420 ( .A(n1162), .B(n12058), .Z(n12057) );
  XOR U11421 ( .A(n12059), .B(n12060), .Z(n12045) );
  AND U11422 ( .A(n1166), .B(n12058), .Z(n12060) );
  XNOR U11423 ( .A(n12059), .B(n12056), .Z(n12058) );
  XOR U11424 ( .A(n12061), .B(n12062), .Z(n12056) );
  AND U11425 ( .A(n1169), .B(n12055), .Z(n12062) );
  XNOR U11426 ( .A(n12063), .B(n12053), .Z(n12055) );
  XOR U11427 ( .A(n12064), .B(n12065), .Z(n12053) );
  AND U11428 ( .A(n1173), .B(n12066), .Z(n12065) );
  XOR U11429 ( .A(p_input[931]), .B(n12064), .Z(n12066) );
  XOR U11430 ( .A(n12067), .B(n12068), .Z(n12064) );
  AND U11431 ( .A(n1177), .B(n12069), .Z(n12068) );
  IV U11432 ( .A(n12061), .Z(n12063) );
  XOR U11433 ( .A(n12070), .B(n12071), .Z(n12061) );
  AND U11434 ( .A(n1181), .B(n12072), .Z(n12071) );
  XOR U11435 ( .A(n12073), .B(n12074), .Z(n12059) );
  AND U11436 ( .A(n1185), .B(n12072), .Z(n12074) );
  XNOR U11437 ( .A(n12073), .B(n12070), .Z(n12072) );
  XOR U11438 ( .A(n12075), .B(n12076), .Z(n12070) );
  AND U11439 ( .A(n1188), .B(n12069), .Z(n12076) );
  XNOR U11440 ( .A(n12077), .B(n12067), .Z(n12069) );
  XOR U11441 ( .A(n12078), .B(n12079), .Z(n12067) );
  AND U11442 ( .A(n1192), .B(n12080), .Z(n12079) );
  XOR U11443 ( .A(p_input[947]), .B(n12078), .Z(n12080) );
  XOR U11444 ( .A(n12081), .B(n12082), .Z(n12078) );
  AND U11445 ( .A(n1196), .B(n12083), .Z(n12082) );
  IV U11446 ( .A(n12075), .Z(n12077) );
  XOR U11447 ( .A(n12084), .B(n12085), .Z(n12075) );
  AND U11448 ( .A(n1200), .B(n12086), .Z(n12085) );
  XOR U11449 ( .A(n12087), .B(n12088), .Z(n12073) );
  AND U11450 ( .A(n1204), .B(n12086), .Z(n12088) );
  XNOR U11451 ( .A(n12087), .B(n12084), .Z(n12086) );
  XOR U11452 ( .A(n12089), .B(n12090), .Z(n12084) );
  AND U11453 ( .A(n1207), .B(n12083), .Z(n12090) );
  XNOR U11454 ( .A(n12091), .B(n12081), .Z(n12083) );
  XOR U11455 ( .A(n12092), .B(n12093), .Z(n12081) );
  AND U11456 ( .A(n1211), .B(n12094), .Z(n12093) );
  XOR U11457 ( .A(p_input[963]), .B(n12092), .Z(n12094) );
  XOR U11458 ( .A(n12095), .B(n12096), .Z(n12092) );
  AND U11459 ( .A(n1215), .B(n12097), .Z(n12096) );
  IV U11460 ( .A(n12089), .Z(n12091) );
  XOR U11461 ( .A(n12098), .B(n12099), .Z(n12089) );
  AND U11462 ( .A(n1219), .B(n12100), .Z(n12099) );
  XOR U11463 ( .A(n12101), .B(n12102), .Z(n12087) );
  AND U11464 ( .A(n1223), .B(n12100), .Z(n12102) );
  XNOR U11465 ( .A(n12101), .B(n12098), .Z(n12100) );
  XOR U11466 ( .A(n12103), .B(n12104), .Z(n12098) );
  AND U11467 ( .A(n1226), .B(n12097), .Z(n12104) );
  XNOR U11468 ( .A(n12105), .B(n12095), .Z(n12097) );
  XOR U11469 ( .A(n12106), .B(n12107), .Z(n12095) );
  AND U11470 ( .A(n1230), .B(n12108), .Z(n12107) );
  XOR U11471 ( .A(p_input[979]), .B(n12106), .Z(n12108) );
  XOR U11472 ( .A(n12109), .B(n12110), .Z(n12106) );
  AND U11473 ( .A(n1234), .B(n12111), .Z(n12110) );
  IV U11474 ( .A(n12103), .Z(n12105) );
  XOR U11475 ( .A(n12112), .B(n12113), .Z(n12103) );
  AND U11476 ( .A(n1238), .B(n12114), .Z(n12113) );
  XOR U11477 ( .A(n12115), .B(n12116), .Z(n12101) );
  AND U11478 ( .A(n1242), .B(n12114), .Z(n12116) );
  XNOR U11479 ( .A(n12115), .B(n12112), .Z(n12114) );
  XOR U11480 ( .A(n12117), .B(n12118), .Z(n12112) );
  AND U11481 ( .A(n1245), .B(n12111), .Z(n12118) );
  XNOR U11482 ( .A(n12119), .B(n12109), .Z(n12111) );
  XOR U11483 ( .A(n12120), .B(n12121), .Z(n12109) );
  AND U11484 ( .A(n1249), .B(n12122), .Z(n12121) );
  XOR U11485 ( .A(p_input[995]), .B(n12120), .Z(n12122) );
  XOR U11486 ( .A(n12123), .B(n12124), .Z(n12120) );
  AND U11487 ( .A(n1253), .B(n12125), .Z(n12124) );
  IV U11488 ( .A(n12117), .Z(n12119) );
  XOR U11489 ( .A(n12126), .B(n12127), .Z(n12117) );
  AND U11490 ( .A(n1257), .B(n12128), .Z(n12127) );
  XOR U11491 ( .A(n12129), .B(n12130), .Z(n12115) );
  AND U11492 ( .A(n1261), .B(n12128), .Z(n12130) );
  XNOR U11493 ( .A(n12129), .B(n12126), .Z(n12128) );
  XOR U11494 ( .A(n12131), .B(n12132), .Z(n12126) );
  AND U11495 ( .A(n1264), .B(n12125), .Z(n12132) );
  XNOR U11496 ( .A(n12133), .B(n12123), .Z(n12125) );
  XOR U11497 ( .A(n12134), .B(n12135), .Z(n12123) );
  AND U11498 ( .A(n1268), .B(n12136), .Z(n12135) );
  XOR U11499 ( .A(p_input[1011]), .B(n12134), .Z(n12136) );
  XOR U11500 ( .A(n12137), .B(n12138), .Z(n12134) );
  AND U11501 ( .A(n1272), .B(n12139), .Z(n12138) );
  IV U11502 ( .A(n12131), .Z(n12133) );
  XOR U11503 ( .A(n12140), .B(n12141), .Z(n12131) );
  AND U11504 ( .A(n1276), .B(n12142), .Z(n12141) );
  XOR U11505 ( .A(n12143), .B(n12144), .Z(n12129) );
  AND U11506 ( .A(n1280), .B(n12142), .Z(n12144) );
  XNOR U11507 ( .A(n12143), .B(n12140), .Z(n12142) );
  XOR U11508 ( .A(n12145), .B(n12146), .Z(n12140) );
  AND U11509 ( .A(n1283), .B(n12139), .Z(n12146) );
  XNOR U11510 ( .A(n12147), .B(n12137), .Z(n12139) );
  XOR U11511 ( .A(n12148), .B(n12149), .Z(n12137) );
  AND U11512 ( .A(n1287), .B(n12150), .Z(n12149) );
  XOR U11513 ( .A(p_input[1027]), .B(n12148), .Z(n12150) );
  XOR U11514 ( .A(n12151), .B(n12152), .Z(n12148) );
  AND U11515 ( .A(n1291), .B(n12153), .Z(n12152) );
  IV U11516 ( .A(n12145), .Z(n12147) );
  XOR U11517 ( .A(n12154), .B(n12155), .Z(n12145) );
  AND U11518 ( .A(n1295), .B(n12156), .Z(n12155) );
  XOR U11519 ( .A(n12157), .B(n12158), .Z(n12143) );
  AND U11520 ( .A(n1299), .B(n12156), .Z(n12158) );
  XNOR U11521 ( .A(n12157), .B(n12154), .Z(n12156) );
  XOR U11522 ( .A(n12159), .B(n12160), .Z(n12154) );
  AND U11523 ( .A(n1302), .B(n12153), .Z(n12160) );
  XNOR U11524 ( .A(n12161), .B(n12151), .Z(n12153) );
  XOR U11525 ( .A(n12162), .B(n12163), .Z(n12151) );
  AND U11526 ( .A(n1306), .B(n12164), .Z(n12163) );
  XOR U11527 ( .A(p_input[1043]), .B(n12162), .Z(n12164) );
  XOR U11528 ( .A(n12165), .B(n12166), .Z(n12162) );
  AND U11529 ( .A(n1310), .B(n12167), .Z(n12166) );
  IV U11530 ( .A(n12159), .Z(n12161) );
  XOR U11531 ( .A(n12168), .B(n12169), .Z(n12159) );
  AND U11532 ( .A(n1314), .B(n12170), .Z(n12169) );
  XOR U11533 ( .A(n12171), .B(n12172), .Z(n12157) );
  AND U11534 ( .A(n1318), .B(n12170), .Z(n12172) );
  XNOR U11535 ( .A(n12171), .B(n12168), .Z(n12170) );
  XOR U11536 ( .A(n12173), .B(n12174), .Z(n12168) );
  AND U11537 ( .A(n1321), .B(n12167), .Z(n12174) );
  XNOR U11538 ( .A(n12175), .B(n12165), .Z(n12167) );
  XOR U11539 ( .A(n12176), .B(n12177), .Z(n12165) );
  AND U11540 ( .A(n1325), .B(n12178), .Z(n12177) );
  XOR U11541 ( .A(p_input[1059]), .B(n12176), .Z(n12178) );
  XOR U11542 ( .A(n12179), .B(n12180), .Z(n12176) );
  AND U11543 ( .A(n1329), .B(n12181), .Z(n12180) );
  IV U11544 ( .A(n12173), .Z(n12175) );
  XOR U11545 ( .A(n12182), .B(n12183), .Z(n12173) );
  AND U11546 ( .A(n1333), .B(n12184), .Z(n12183) );
  XOR U11547 ( .A(n12185), .B(n12186), .Z(n12171) );
  AND U11548 ( .A(n1337), .B(n12184), .Z(n12186) );
  XNOR U11549 ( .A(n12185), .B(n12182), .Z(n12184) );
  XOR U11550 ( .A(n12187), .B(n12188), .Z(n12182) );
  AND U11551 ( .A(n1340), .B(n12181), .Z(n12188) );
  XNOR U11552 ( .A(n12189), .B(n12179), .Z(n12181) );
  XOR U11553 ( .A(n12190), .B(n12191), .Z(n12179) );
  AND U11554 ( .A(n1344), .B(n12192), .Z(n12191) );
  XOR U11555 ( .A(p_input[1075]), .B(n12190), .Z(n12192) );
  XOR U11556 ( .A(n12193), .B(n12194), .Z(n12190) );
  AND U11557 ( .A(n1348), .B(n12195), .Z(n12194) );
  IV U11558 ( .A(n12187), .Z(n12189) );
  XOR U11559 ( .A(n12196), .B(n12197), .Z(n12187) );
  AND U11560 ( .A(n1352), .B(n12198), .Z(n12197) );
  XOR U11561 ( .A(n12199), .B(n12200), .Z(n12185) );
  AND U11562 ( .A(n1356), .B(n12198), .Z(n12200) );
  XNOR U11563 ( .A(n12199), .B(n12196), .Z(n12198) );
  XOR U11564 ( .A(n12201), .B(n12202), .Z(n12196) );
  AND U11565 ( .A(n1359), .B(n12195), .Z(n12202) );
  XNOR U11566 ( .A(n12203), .B(n12193), .Z(n12195) );
  XOR U11567 ( .A(n12204), .B(n12205), .Z(n12193) );
  AND U11568 ( .A(n1363), .B(n12206), .Z(n12205) );
  XOR U11569 ( .A(p_input[1091]), .B(n12204), .Z(n12206) );
  XOR U11570 ( .A(n12207), .B(n12208), .Z(n12204) );
  AND U11571 ( .A(n1367), .B(n12209), .Z(n12208) );
  IV U11572 ( .A(n12201), .Z(n12203) );
  XOR U11573 ( .A(n12210), .B(n12211), .Z(n12201) );
  AND U11574 ( .A(n1371), .B(n12212), .Z(n12211) );
  XOR U11575 ( .A(n12213), .B(n12214), .Z(n12199) );
  AND U11576 ( .A(n1375), .B(n12212), .Z(n12214) );
  XNOR U11577 ( .A(n12213), .B(n12210), .Z(n12212) );
  XOR U11578 ( .A(n12215), .B(n12216), .Z(n12210) );
  AND U11579 ( .A(n1378), .B(n12209), .Z(n12216) );
  XNOR U11580 ( .A(n12217), .B(n12207), .Z(n12209) );
  XOR U11581 ( .A(n12218), .B(n12219), .Z(n12207) );
  AND U11582 ( .A(n1382), .B(n12220), .Z(n12219) );
  XOR U11583 ( .A(p_input[1107]), .B(n12218), .Z(n12220) );
  XOR U11584 ( .A(n12221), .B(n12222), .Z(n12218) );
  AND U11585 ( .A(n1386), .B(n12223), .Z(n12222) );
  IV U11586 ( .A(n12215), .Z(n12217) );
  XOR U11587 ( .A(n12224), .B(n12225), .Z(n12215) );
  AND U11588 ( .A(n1390), .B(n12226), .Z(n12225) );
  XOR U11589 ( .A(n12227), .B(n12228), .Z(n12213) );
  AND U11590 ( .A(n1394), .B(n12226), .Z(n12228) );
  XNOR U11591 ( .A(n12227), .B(n12224), .Z(n12226) );
  XOR U11592 ( .A(n12229), .B(n12230), .Z(n12224) );
  AND U11593 ( .A(n1397), .B(n12223), .Z(n12230) );
  XNOR U11594 ( .A(n12231), .B(n12221), .Z(n12223) );
  XOR U11595 ( .A(n12232), .B(n12233), .Z(n12221) );
  AND U11596 ( .A(n1401), .B(n12234), .Z(n12233) );
  XOR U11597 ( .A(p_input[1123]), .B(n12232), .Z(n12234) );
  XOR U11598 ( .A(n12235), .B(n12236), .Z(n12232) );
  AND U11599 ( .A(n1405), .B(n12237), .Z(n12236) );
  IV U11600 ( .A(n12229), .Z(n12231) );
  XOR U11601 ( .A(n12238), .B(n12239), .Z(n12229) );
  AND U11602 ( .A(n1409), .B(n12240), .Z(n12239) );
  XOR U11603 ( .A(n12241), .B(n12242), .Z(n12227) );
  AND U11604 ( .A(n1413), .B(n12240), .Z(n12242) );
  XNOR U11605 ( .A(n12241), .B(n12238), .Z(n12240) );
  XOR U11606 ( .A(n12243), .B(n12244), .Z(n12238) );
  AND U11607 ( .A(n1416), .B(n12237), .Z(n12244) );
  XNOR U11608 ( .A(n12245), .B(n12235), .Z(n12237) );
  XOR U11609 ( .A(n12246), .B(n12247), .Z(n12235) );
  AND U11610 ( .A(n1420), .B(n12248), .Z(n12247) );
  XOR U11611 ( .A(p_input[1139]), .B(n12246), .Z(n12248) );
  XOR U11612 ( .A(n12249), .B(n12250), .Z(n12246) );
  AND U11613 ( .A(n1424), .B(n12251), .Z(n12250) );
  IV U11614 ( .A(n12243), .Z(n12245) );
  XOR U11615 ( .A(n12252), .B(n12253), .Z(n12243) );
  AND U11616 ( .A(n1428), .B(n12254), .Z(n12253) );
  XOR U11617 ( .A(n12255), .B(n12256), .Z(n12241) );
  AND U11618 ( .A(n1432), .B(n12254), .Z(n12256) );
  XNOR U11619 ( .A(n12255), .B(n12252), .Z(n12254) );
  XOR U11620 ( .A(n12257), .B(n12258), .Z(n12252) );
  AND U11621 ( .A(n1435), .B(n12251), .Z(n12258) );
  XNOR U11622 ( .A(n12259), .B(n12249), .Z(n12251) );
  XOR U11623 ( .A(n12260), .B(n12261), .Z(n12249) );
  AND U11624 ( .A(n1439), .B(n12262), .Z(n12261) );
  XOR U11625 ( .A(p_input[1155]), .B(n12260), .Z(n12262) );
  XOR U11626 ( .A(n12263), .B(n12264), .Z(n12260) );
  AND U11627 ( .A(n1443), .B(n12265), .Z(n12264) );
  IV U11628 ( .A(n12257), .Z(n12259) );
  XOR U11629 ( .A(n12266), .B(n12267), .Z(n12257) );
  AND U11630 ( .A(n1447), .B(n12268), .Z(n12267) );
  XOR U11631 ( .A(n12269), .B(n12270), .Z(n12255) );
  AND U11632 ( .A(n1451), .B(n12268), .Z(n12270) );
  XNOR U11633 ( .A(n12269), .B(n12266), .Z(n12268) );
  XOR U11634 ( .A(n12271), .B(n12272), .Z(n12266) );
  AND U11635 ( .A(n1454), .B(n12265), .Z(n12272) );
  XNOR U11636 ( .A(n12273), .B(n12263), .Z(n12265) );
  XOR U11637 ( .A(n12274), .B(n12275), .Z(n12263) );
  AND U11638 ( .A(n1458), .B(n12276), .Z(n12275) );
  XOR U11639 ( .A(p_input[1171]), .B(n12274), .Z(n12276) );
  XOR U11640 ( .A(n12277), .B(n12278), .Z(n12274) );
  AND U11641 ( .A(n1462), .B(n12279), .Z(n12278) );
  IV U11642 ( .A(n12271), .Z(n12273) );
  XOR U11643 ( .A(n12280), .B(n12281), .Z(n12271) );
  AND U11644 ( .A(n1466), .B(n12282), .Z(n12281) );
  XOR U11645 ( .A(n12283), .B(n12284), .Z(n12269) );
  AND U11646 ( .A(n1470), .B(n12282), .Z(n12284) );
  XNOR U11647 ( .A(n12283), .B(n12280), .Z(n12282) );
  XOR U11648 ( .A(n12285), .B(n12286), .Z(n12280) );
  AND U11649 ( .A(n1473), .B(n12279), .Z(n12286) );
  XNOR U11650 ( .A(n12287), .B(n12277), .Z(n12279) );
  XOR U11651 ( .A(n12288), .B(n12289), .Z(n12277) );
  AND U11652 ( .A(n1477), .B(n12290), .Z(n12289) );
  XOR U11653 ( .A(p_input[1187]), .B(n12288), .Z(n12290) );
  XOR U11654 ( .A(n12291), .B(n12292), .Z(n12288) );
  AND U11655 ( .A(n1481), .B(n12293), .Z(n12292) );
  IV U11656 ( .A(n12285), .Z(n12287) );
  XOR U11657 ( .A(n12294), .B(n12295), .Z(n12285) );
  AND U11658 ( .A(n1485), .B(n12296), .Z(n12295) );
  XOR U11659 ( .A(n12297), .B(n12298), .Z(n12283) );
  AND U11660 ( .A(n1489), .B(n12296), .Z(n12298) );
  XNOR U11661 ( .A(n12297), .B(n12294), .Z(n12296) );
  XOR U11662 ( .A(n12299), .B(n12300), .Z(n12294) );
  AND U11663 ( .A(n1492), .B(n12293), .Z(n12300) );
  XNOR U11664 ( .A(n12301), .B(n12291), .Z(n12293) );
  XOR U11665 ( .A(n12302), .B(n12303), .Z(n12291) );
  AND U11666 ( .A(n1496), .B(n12304), .Z(n12303) );
  XOR U11667 ( .A(p_input[1203]), .B(n12302), .Z(n12304) );
  XOR U11668 ( .A(n12305), .B(n12306), .Z(n12302) );
  AND U11669 ( .A(n1500), .B(n12307), .Z(n12306) );
  IV U11670 ( .A(n12299), .Z(n12301) );
  XOR U11671 ( .A(n12308), .B(n12309), .Z(n12299) );
  AND U11672 ( .A(n1504), .B(n12310), .Z(n12309) );
  XOR U11673 ( .A(n12311), .B(n12312), .Z(n12297) );
  AND U11674 ( .A(n1508), .B(n12310), .Z(n12312) );
  XNOR U11675 ( .A(n12311), .B(n12308), .Z(n12310) );
  XOR U11676 ( .A(n12313), .B(n12314), .Z(n12308) );
  AND U11677 ( .A(n1511), .B(n12307), .Z(n12314) );
  XNOR U11678 ( .A(n12315), .B(n12305), .Z(n12307) );
  XOR U11679 ( .A(n12316), .B(n12317), .Z(n12305) );
  AND U11680 ( .A(n1515), .B(n12318), .Z(n12317) );
  XOR U11681 ( .A(p_input[1219]), .B(n12316), .Z(n12318) );
  XOR U11682 ( .A(n12319), .B(n12320), .Z(n12316) );
  AND U11683 ( .A(n1519), .B(n12321), .Z(n12320) );
  IV U11684 ( .A(n12313), .Z(n12315) );
  XOR U11685 ( .A(n12322), .B(n12323), .Z(n12313) );
  AND U11686 ( .A(n1523), .B(n12324), .Z(n12323) );
  XOR U11687 ( .A(n12325), .B(n12326), .Z(n12311) );
  AND U11688 ( .A(n1527), .B(n12324), .Z(n12326) );
  XNOR U11689 ( .A(n12325), .B(n12322), .Z(n12324) );
  XOR U11690 ( .A(n12327), .B(n12328), .Z(n12322) );
  AND U11691 ( .A(n1530), .B(n12321), .Z(n12328) );
  XNOR U11692 ( .A(n12329), .B(n12319), .Z(n12321) );
  XOR U11693 ( .A(n12330), .B(n12331), .Z(n12319) );
  AND U11694 ( .A(n1534), .B(n12332), .Z(n12331) );
  XOR U11695 ( .A(p_input[1235]), .B(n12330), .Z(n12332) );
  XOR U11696 ( .A(n12333), .B(n12334), .Z(n12330) );
  AND U11697 ( .A(n1538), .B(n12335), .Z(n12334) );
  IV U11698 ( .A(n12327), .Z(n12329) );
  XOR U11699 ( .A(n12336), .B(n12337), .Z(n12327) );
  AND U11700 ( .A(n1542), .B(n12338), .Z(n12337) );
  XOR U11701 ( .A(n12339), .B(n12340), .Z(n12325) );
  AND U11702 ( .A(n1546), .B(n12338), .Z(n12340) );
  XNOR U11703 ( .A(n12339), .B(n12336), .Z(n12338) );
  XOR U11704 ( .A(n12341), .B(n12342), .Z(n12336) );
  AND U11705 ( .A(n1549), .B(n12335), .Z(n12342) );
  XNOR U11706 ( .A(n12343), .B(n12333), .Z(n12335) );
  XOR U11707 ( .A(n12344), .B(n12345), .Z(n12333) );
  AND U11708 ( .A(n1553), .B(n12346), .Z(n12345) );
  XOR U11709 ( .A(p_input[1251]), .B(n12344), .Z(n12346) );
  XOR U11710 ( .A(n12347), .B(n12348), .Z(n12344) );
  AND U11711 ( .A(n1557), .B(n12349), .Z(n12348) );
  IV U11712 ( .A(n12341), .Z(n12343) );
  XOR U11713 ( .A(n12350), .B(n12351), .Z(n12341) );
  AND U11714 ( .A(n1561), .B(n12352), .Z(n12351) );
  XOR U11715 ( .A(n12353), .B(n12354), .Z(n12339) );
  AND U11716 ( .A(n1565), .B(n12352), .Z(n12354) );
  XNOR U11717 ( .A(n12353), .B(n12350), .Z(n12352) );
  XOR U11718 ( .A(n12355), .B(n12356), .Z(n12350) );
  AND U11719 ( .A(n1568), .B(n12349), .Z(n12356) );
  XNOR U11720 ( .A(n12357), .B(n12347), .Z(n12349) );
  XOR U11721 ( .A(n12358), .B(n12359), .Z(n12347) );
  AND U11722 ( .A(n1572), .B(n12360), .Z(n12359) );
  XOR U11723 ( .A(p_input[1267]), .B(n12358), .Z(n12360) );
  XOR U11724 ( .A(n12361), .B(n12362), .Z(n12358) );
  AND U11725 ( .A(n1576), .B(n12363), .Z(n12362) );
  IV U11726 ( .A(n12355), .Z(n12357) );
  XOR U11727 ( .A(n12364), .B(n12365), .Z(n12355) );
  AND U11728 ( .A(n1580), .B(n12366), .Z(n12365) );
  XOR U11729 ( .A(n12367), .B(n12368), .Z(n12353) );
  AND U11730 ( .A(n1584), .B(n12366), .Z(n12368) );
  XNOR U11731 ( .A(n12367), .B(n12364), .Z(n12366) );
  XOR U11732 ( .A(n12369), .B(n12370), .Z(n12364) );
  AND U11733 ( .A(n1587), .B(n12363), .Z(n12370) );
  XNOR U11734 ( .A(n12371), .B(n12361), .Z(n12363) );
  XOR U11735 ( .A(n12372), .B(n12373), .Z(n12361) );
  AND U11736 ( .A(n1591), .B(n12374), .Z(n12373) );
  XOR U11737 ( .A(p_input[1283]), .B(n12372), .Z(n12374) );
  XOR U11738 ( .A(n12375), .B(n12376), .Z(n12372) );
  AND U11739 ( .A(n1595), .B(n12377), .Z(n12376) );
  IV U11740 ( .A(n12369), .Z(n12371) );
  XOR U11741 ( .A(n12378), .B(n12379), .Z(n12369) );
  AND U11742 ( .A(n1599), .B(n12380), .Z(n12379) );
  XOR U11743 ( .A(n12381), .B(n12382), .Z(n12367) );
  AND U11744 ( .A(n1603), .B(n12380), .Z(n12382) );
  XNOR U11745 ( .A(n12381), .B(n12378), .Z(n12380) );
  XOR U11746 ( .A(n12383), .B(n12384), .Z(n12378) );
  AND U11747 ( .A(n1606), .B(n12377), .Z(n12384) );
  XNOR U11748 ( .A(n12385), .B(n12375), .Z(n12377) );
  XOR U11749 ( .A(n12386), .B(n12387), .Z(n12375) );
  AND U11750 ( .A(n1610), .B(n12388), .Z(n12387) );
  XOR U11751 ( .A(p_input[1299]), .B(n12386), .Z(n12388) );
  XOR U11752 ( .A(n12389), .B(n12390), .Z(n12386) );
  AND U11753 ( .A(n1614), .B(n12391), .Z(n12390) );
  IV U11754 ( .A(n12383), .Z(n12385) );
  XOR U11755 ( .A(n12392), .B(n12393), .Z(n12383) );
  AND U11756 ( .A(n1618), .B(n12394), .Z(n12393) );
  XOR U11757 ( .A(n12395), .B(n12396), .Z(n12381) );
  AND U11758 ( .A(n1622), .B(n12394), .Z(n12396) );
  XNOR U11759 ( .A(n12395), .B(n12392), .Z(n12394) );
  XOR U11760 ( .A(n12397), .B(n12398), .Z(n12392) );
  AND U11761 ( .A(n1625), .B(n12391), .Z(n12398) );
  XNOR U11762 ( .A(n12399), .B(n12389), .Z(n12391) );
  XOR U11763 ( .A(n12400), .B(n12401), .Z(n12389) );
  AND U11764 ( .A(n1629), .B(n12402), .Z(n12401) );
  XOR U11765 ( .A(p_input[1315]), .B(n12400), .Z(n12402) );
  XOR U11766 ( .A(n12403), .B(n12404), .Z(n12400) );
  AND U11767 ( .A(n1633), .B(n12405), .Z(n12404) );
  IV U11768 ( .A(n12397), .Z(n12399) );
  XOR U11769 ( .A(n12406), .B(n12407), .Z(n12397) );
  AND U11770 ( .A(n1637), .B(n12408), .Z(n12407) );
  XOR U11771 ( .A(n12409), .B(n12410), .Z(n12395) );
  AND U11772 ( .A(n1641), .B(n12408), .Z(n12410) );
  XNOR U11773 ( .A(n12409), .B(n12406), .Z(n12408) );
  XOR U11774 ( .A(n12411), .B(n12412), .Z(n12406) );
  AND U11775 ( .A(n1644), .B(n12405), .Z(n12412) );
  XNOR U11776 ( .A(n12413), .B(n12403), .Z(n12405) );
  XOR U11777 ( .A(n12414), .B(n12415), .Z(n12403) );
  AND U11778 ( .A(n1648), .B(n12416), .Z(n12415) );
  XOR U11779 ( .A(p_input[1331]), .B(n12414), .Z(n12416) );
  XOR U11780 ( .A(n12417), .B(n12418), .Z(n12414) );
  AND U11781 ( .A(n1652), .B(n12419), .Z(n12418) );
  IV U11782 ( .A(n12411), .Z(n12413) );
  XOR U11783 ( .A(n12420), .B(n12421), .Z(n12411) );
  AND U11784 ( .A(n1656), .B(n12422), .Z(n12421) );
  XOR U11785 ( .A(n12423), .B(n12424), .Z(n12409) );
  AND U11786 ( .A(n1660), .B(n12422), .Z(n12424) );
  XNOR U11787 ( .A(n12423), .B(n12420), .Z(n12422) );
  XOR U11788 ( .A(n12425), .B(n12426), .Z(n12420) );
  AND U11789 ( .A(n1663), .B(n12419), .Z(n12426) );
  XNOR U11790 ( .A(n12427), .B(n12417), .Z(n12419) );
  XOR U11791 ( .A(n12428), .B(n12429), .Z(n12417) );
  AND U11792 ( .A(n1667), .B(n12430), .Z(n12429) );
  XOR U11793 ( .A(p_input[1347]), .B(n12428), .Z(n12430) );
  XOR U11794 ( .A(n12431), .B(n12432), .Z(n12428) );
  AND U11795 ( .A(n1671), .B(n12433), .Z(n12432) );
  IV U11796 ( .A(n12425), .Z(n12427) );
  XOR U11797 ( .A(n12434), .B(n12435), .Z(n12425) );
  AND U11798 ( .A(n1675), .B(n12436), .Z(n12435) );
  XOR U11799 ( .A(n12437), .B(n12438), .Z(n12423) );
  AND U11800 ( .A(n1679), .B(n12436), .Z(n12438) );
  XNOR U11801 ( .A(n12437), .B(n12434), .Z(n12436) );
  XOR U11802 ( .A(n12439), .B(n12440), .Z(n12434) );
  AND U11803 ( .A(n1682), .B(n12433), .Z(n12440) );
  XNOR U11804 ( .A(n12441), .B(n12431), .Z(n12433) );
  XOR U11805 ( .A(n12442), .B(n12443), .Z(n12431) );
  AND U11806 ( .A(n1686), .B(n12444), .Z(n12443) );
  XOR U11807 ( .A(p_input[1363]), .B(n12442), .Z(n12444) );
  XOR U11808 ( .A(n12445), .B(n12446), .Z(n12442) );
  AND U11809 ( .A(n1690), .B(n12447), .Z(n12446) );
  IV U11810 ( .A(n12439), .Z(n12441) );
  XOR U11811 ( .A(n12448), .B(n12449), .Z(n12439) );
  AND U11812 ( .A(n1694), .B(n12450), .Z(n12449) );
  XOR U11813 ( .A(n12451), .B(n12452), .Z(n12437) );
  AND U11814 ( .A(n1698), .B(n12450), .Z(n12452) );
  XNOR U11815 ( .A(n12451), .B(n12448), .Z(n12450) );
  XOR U11816 ( .A(n12453), .B(n12454), .Z(n12448) );
  AND U11817 ( .A(n1701), .B(n12447), .Z(n12454) );
  XNOR U11818 ( .A(n12455), .B(n12445), .Z(n12447) );
  XOR U11819 ( .A(n12456), .B(n12457), .Z(n12445) );
  AND U11820 ( .A(n1705), .B(n12458), .Z(n12457) );
  XOR U11821 ( .A(p_input[1379]), .B(n12456), .Z(n12458) );
  XOR U11822 ( .A(n12459), .B(n12460), .Z(n12456) );
  AND U11823 ( .A(n1709), .B(n12461), .Z(n12460) );
  IV U11824 ( .A(n12453), .Z(n12455) );
  XOR U11825 ( .A(n12462), .B(n12463), .Z(n12453) );
  AND U11826 ( .A(n1713), .B(n12464), .Z(n12463) );
  XOR U11827 ( .A(n12465), .B(n12466), .Z(n12451) );
  AND U11828 ( .A(n1717), .B(n12464), .Z(n12466) );
  XNOR U11829 ( .A(n12465), .B(n12462), .Z(n12464) );
  XOR U11830 ( .A(n12467), .B(n12468), .Z(n12462) );
  AND U11831 ( .A(n1720), .B(n12461), .Z(n12468) );
  XNOR U11832 ( .A(n12469), .B(n12459), .Z(n12461) );
  XOR U11833 ( .A(n12470), .B(n12471), .Z(n12459) );
  AND U11834 ( .A(n1724), .B(n12472), .Z(n12471) );
  XOR U11835 ( .A(p_input[1395]), .B(n12470), .Z(n12472) );
  XOR U11836 ( .A(n12473), .B(n12474), .Z(n12470) );
  AND U11837 ( .A(n1728), .B(n12475), .Z(n12474) );
  IV U11838 ( .A(n12467), .Z(n12469) );
  XOR U11839 ( .A(n12476), .B(n12477), .Z(n12467) );
  AND U11840 ( .A(n1732), .B(n12478), .Z(n12477) );
  XOR U11841 ( .A(n12479), .B(n12480), .Z(n12465) );
  AND U11842 ( .A(n1736), .B(n12478), .Z(n12480) );
  XNOR U11843 ( .A(n12479), .B(n12476), .Z(n12478) );
  XOR U11844 ( .A(n12481), .B(n12482), .Z(n12476) );
  AND U11845 ( .A(n1739), .B(n12475), .Z(n12482) );
  XNOR U11846 ( .A(n12483), .B(n12473), .Z(n12475) );
  XOR U11847 ( .A(n12484), .B(n12485), .Z(n12473) );
  AND U11848 ( .A(n1743), .B(n12486), .Z(n12485) );
  XOR U11849 ( .A(p_input[1411]), .B(n12484), .Z(n12486) );
  XOR U11850 ( .A(n12487), .B(n12488), .Z(n12484) );
  AND U11851 ( .A(n1747), .B(n12489), .Z(n12488) );
  IV U11852 ( .A(n12481), .Z(n12483) );
  XOR U11853 ( .A(n12490), .B(n12491), .Z(n12481) );
  AND U11854 ( .A(n1751), .B(n12492), .Z(n12491) );
  XOR U11855 ( .A(n12493), .B(n12494), .Z(n12479) );
  AND U11856 ( .A(n1755), .B(n12492), .Z(n12494) );
  XNOR U11857 ( .A(n12493), .B(n12490), .Z(n12492) );
  XOR U11858 ( .A(n12495), .B(n12496), .Z(n12490) );
  AND U11859 ( .A(n1758), .B(n12489), .Z(n12496) );
  XNOR U11860 ( .A(n12497), .B(n12487), .Z(n12489) );
  XOR U11861 ( .A(n12498), .B(n12499), .Z(n12487) );
  AND U11862 ( .A(n1762), .B(n12500), .Z(n12499) );
  XOR U11863 ( .A(p_input[1427]), .B(n12498), .Z(n12500) );
  XOR U11864 ( .A(n12501), .B(n12502), .Z(n12498) );
  AND U11865 ( .A(n1766), .B(n12503), .Z(n12502) );
  IV U11866 ( .A(n12495), .Z(n12497) );
  XOR U11867 ( .A(n12504), .B(n12505), .Z(n12495) );
  AND U11868 ( .A(n1770), .B(n12506), .Z(n12505) );
  XOR U11869 ( .A(n12507), .B(n12508), .Z(n12493) );
  AND U11870 ( .A(n1774), .B(n12506), .Z(n12508) );
  XNOR U11871 ( .A(n12507), .B(n12504), .Z(n12506) );
  XOR U11872 ( .A(n12509), .B(n12510), .Z(n12504) );
  AND U11873 ( .A(n1777), .B(n12503), .Z(n12510) );
  XNOR U11874 ( .A(n12511), .B(n12501), .Z(n12503) );
  XOR U11875 ( .A(n12512), .B(n12513), .Z(n12501) );
  AND U11876 ( .A(n1781), .B(n12514), .Z(n12513) );
  XOR U11877 ( .A(p_input[1443]), .B(n12512), .Z(n12514) );
  XOR U11878 ( .A(n12515), .B(n12516), .Z(n12512) );
  AND U11879 ( .A(n1785), .B(n12517), .Z(n12516) );
  IV U11880 ( .A(n12509), .Z(n12511) );
  XOR U11881 ( .A(n12518), .B(n12519), .Z(n12509) );
  AND U11882 ( .A(n1789), .B(n12520), .Z(n12519) );
  XOR U11883 ( .A(n12521), .B(n12522), .Z(n12507) );
  AND U11884 ( .A(n1793), .B(n12520), .Z(n12522) );
  XNOR U11885 ( .A(n12521), .B(n12518), .Z(n12520) );
  XOR U11886 ( .A(n12523), .B(n12524), .Z(n12518) );
  AND U11887 ( .A(n1796), .B(n12517), .Z(n12524) );
  XNOR U11888 ( .A(n12525), .B(n12515), .Z(n12517) );
  XOR U11889 ( .A(n12526), .B(n12527), .Z(n12515) );
  AND U11890 ( .A(n1800), .B(n12528), .Z(n12527) );
  XOR U11891 ( .A(p_input[1459]), .B(n12526), .Z(n12528) );
  XOR U11892 ( .A(n12529), .B(n12530), .Z(n12526) );
  AND U11893 ( .A(n1804), .B(n12531), .Z(n12530) );
  IV U11894 ( .A(n12523), .Z(n12525) );
  XOR U11895 ( .A(n12532), .B(n12533), .Z(n12523) );
  AND U11896 ( .A(n1808), .B(n12534), .Z(n12533) );
  XOR U11897 ( .A(n12535), .B(n12536), .Z(n12521) );
  AND U11898 ( .A(n1812), .B(n12534), .Z(n12536) );
  XNOR U11899 ( .A(n12535), .B(n12532), .Z(n12534) );
  XOR U11900 ( .A(n12537), .B(n12538), .Z(n12532) );
  AND U11901 ( .A(n1815), .B(n12531), .Z(n12538) );
  XNOR U11902 ( .A(n12539), .B(n12529), .Z(n12531) );
  XOR U11903 ( .A(n12540), .B(n12541), .Z(n12529) );
  AND U11904 ( .A(n1819), .B(n12542), .Z(n12541) );
  XOR U11905 ( .A(p_input[1475]), .B(n12540), .Z(n12542) );
  XOR U11906 ( .A(n12543), .B(n12544), .Z(n12540) );
  AND U11907 ( .A(n1823), .B(n12545), .Z(n12544) );
  IV U11908 ( .A(n12537), .Z(n12539) );
  XOR U11909 ( .A(n12546), .B(n12547), .Z(n12537) );
  AND U11910 ( .A(n1827), .B(n12548), .Z(n12547) );
  XOR U11911 ( .A(n12549), .B(n12550), .Z(n12535) );
  AND U11912 ( .A(n1831), .B(n12548), .Z(n12550) );
  XNOR U11913 ( .A(n12549), .B(n12546), .Z(n12548) );
  XOR U11914 ( .A(n12551), .B(n12552), .Z(n12546) );
  AND U11915 ( .A(n1834), .B(n12545), .Z(n12552) );
  XNOR U11916 ( .A(n12553), .B(n12543), .Z(n12545) );
  XOR U11917 ( .A(n12554), .B(n12555), .Z(n12543) );
  AND U11918 ( .A(n1838), .B(n12556), .Z(n12555) );
  XOR U11919 ( .A(p_input[1491]), .B(n12554), .Z(n12556) );
  XOR U11920 ( .A(n12557), .B(n12558), .Z(n12554) );
  AND U11921 ( .A(n1842), .B(n12559), .Z(n12558) );
  IV U11922 ( .A(n12551), .Z(n12553) );
  XOR U11923 ( .A(n12560), .B(n12561), .Z(n12551) );
  AND U11924 ( .A(n1846), .B(n12562), .Z(n12561) );
  XOR U11925 ( .A(n12563), .B(n12564), .Z(n12549) );
  AND U11926 ( .A(n1850), .B(n12562), .Z(n12564) );
  XNOR U11927 ( .A(n12563), .B(n12560), .Z(n12562) );
  XOR U11928 ( .A(n12565), .B(n12566), .Z(n12560) );
  AND U11929 ( .A(n1853), .B(n12559), .Z(n12566) );
  XNOR U11930 ( .A(n12567), .B(n12557), .Z(n12559) );
  XOR U11931 ( .A(n12568), .B(n12569), .Z(n12557) );
  AND U11932 ( .A(n1857), .B(n12570), .Z(n12569) );
  XOR U11933 ( .A(p_input[1507]), .B(n12568), .Z(n12570) );
  XOR U11934 ( .A(n12571), .B(n12572), .Z(n12568) );
  AND U11935 ( .A(n1861), .B(n12573), .Z(n12572) );
  IV U11936 ( .A(n12565), .Z(n12567) );
  XOR U11937 ( .A(n12574), .B(n12575), .Z(n12565) );
  AND U11938 ( .A(n1865), .B(n12576), .Z(n12575) );
  XOR U11939 ( .A(n12577), .B(n12578), .Z(n12563) );
  AND U11940 ( .A(n1869), .B(n12576), .Z(n12578) );
  XNOR U11941 ( .A(n12577), .B(n12574), .Z(n12576) );
  XOR U11942 ( .A(n12579), .B(n12580), .Z(n12574) );
  AND U11943 ( .A(n1872), .B(n12573), .Z(n12580) );
  XNOR U11944 ( .A(n12581), .B(n12571), .Z(n12573) );
  XOR U11945 ( .A(n12582), .B(n12583), .Z(n12571) );
  AND U11946 ( .A(n1876), .B(n12584), .Z(n12583) );
  XOR U11947 ( .A(p_input[1523]), .B(n12582), .Z(n12584) );
  XOR U11948 ( .A(n12585), .B(n12586), .Z(n12582) );
  AND U11949 ( .A(n1880), .B(n12587), .Z(n12586) );
  IV U11950 ( .A(n12579), .Z(n12581) );
  XOR U11951 ( .A(n12588), .B(n12589), .Z(n12579) );
  AND U11952 ( .A(n1884), .B(n12590), .Z(n12589) );
  XOR U11953 ( .A(n12591), .B(n12592), .Z(n12577) );
  AND U11954 ( .A(n1888), .B(n12590), .Z(n12592) );
  XNOR U11955 ( .A(n12591), .B(n12588), .Z(n12590) );
  XOR U11956 ( .A(n12593), .B(n12594), .Z(n12588) );
  AND U11957 ( .A(n1891), .B(n12587), .Z(n12594) );
  XNOR U11958 ( .A(n12595), .B(n12585), .Z(n12587) );
  XOR U11959 ( .A(n12596), .B(n12597), .Z(n12585) );
  AND U11960 ( .A(n1895), .B(n12598), .Z(n12597) );
  XOR U11961 ( .A(p_input[1539]), .B(n12596), .Z(n12598) );
  XOR U11962 ( .A(n12599), .B(n12600), .Z(n12596) );
  AND U11963 ( .A(n1899), .B(n12601), .Z(n12600) );
  IV U11964 ( .A(n12593), .Z(n12595) );
  XOR U11965 ( .A(n12602), .B(n12603), .Z(n12593) );
  AND U11966 ( .A(n1903), .B(n12604), .Z(n12603) );
  XOR U11967 ( .A(n12605), .B(n12606), .Z(n12591) );
  AND U11968 ( .A(n1907), .B(n12604), .Z(n12606) );
  XNOR U11969 ( .A(n12605), .B(n12602), .Z(n12604) );
  XOR U11970 ( .A(n12607), .B(n12608), .Z(n12602) );
  AND U11971 ( .A(n1910), .B(n12601), .Z(n12608) );
  XNOR U11972 ( .A(n12609), .B(n12599), .Z(n12601) );
  XOR U11973 ( .A(n12610), .B(n12611), .Z(n12599) );
  AND U11974 ( .A(n1914), .B(n12612), .Z(n12611) );
  XOR U11975 ( .A(p_input[1555]), .B(n12610), .Z(n12612) );
  XOR U11976 ( .A(n12613), .B(n12614), .Z(n12610) );
  AND U11977 ( .A(n1918), .B(n12615), .Z(n12614) );
  IV U11978 ( .A(n12607), .Z(n12609) );
  XOR U11979 ( .A(n12616), .B(n12617), .Z(n12607) );
  AND U11980 ( .A(n1922), .B(n12618), .Z(n12617) );
  XOR U11981 ( .A(n12619), .B(n12620), .Z(n12605) );
  AND U11982 ( .A(n1926), .B(n12618), .Z(n12620) );
  XNOR U11983 ( .A(n12619), .B(n12616), .Z(n12618) );
  XOR U11984 ( .A(n12621), .B(n12622), .Z(n12616) );
  AND U11985 ( .A(n1929), .B(n12615), .Z(n12622) );
  XNOR U11986 ( .A(n12623), .B(n12613), .Z(n12615) );
  XOR U11987 ( .A(n12624), .B(n12625), .Z(n12613) );
  AND U11988 ( .A(n1933), .B(n12626), .Z(n12625) );
  XOR U11989 ( .A(p_input[1571]), .B(n12624), .Z(n12626) );
  XOR U11990 ( .A(n12627), .B(n12628), .Z(n12624) );
  AND U11991 ( .A(n1937), .B(n12629), .Z(n12628) );
  IV U11992 ( .A(n12621), .Z(n12623) );
  XOR U11993 ( .A(n12630), .B(n12631), .Z(n12621) );
  AND U11994 ( .A(n1941), .B(n12632), .Z(n12631) );
  XOR U11995 ( .A(n12633), .B(n12634), .Z(n12619) );
  AND U11996 ( .A(n1945), .B(n12632), .Z(n12634) );
  XNOR U11997 ( .A(n12633), .B(n12630), .Z(n12632) );
  XOR U11998 ( .A(n12635), .B(n12636), .Z(n12630) );
  AND U11999 ( .A(n1948), .B(n12629), .Z(n12636) );
  XNOR U12000 ( .A(n12637), .B(n12627), .Z(n12629) );
  XOR U12001 ( .A(n12638), .B(n12639), .Z(n12627) );
  AND U12002 ( .A(n1952), .B(n12640), .Z(n12639) );
  XOR U12003 ( .A(p_input[1587]), .B(n12638), .Z(n12640) );
  XOR U12004 ( .A(n12641), .B(n12642), .Z(n12638) );
  AND U12005 ( .A(n1956), .B(n12643), .Z(n12642) );
  IV U12006 ( .A(n12635), .Z(n12637) );
  XOR U12007 ( .A(n12644), .B(n12645), .Z(n12635) );
  AND U12008 ( .A(n1960), .B(n12646), .Z(n12645) );
  XOR U12009 ( .A(n12647), .B(n12648), .Z(n12633) );
  AND U12010 ( .A(n1964), .B(n12646), .Z(n12648) );
  XNOR U12011 ( .A(n12647), .B(n12644), .Z(n12646) );
  XOR U12012 ( .A(n12649), .B(n12650), .Z(n12644) );
  AND U12013 ( .A(n1967), .B(n12643), .Z(n12650) );
  XNOR U12014 ( .A(n12651), .B(n12641), .Z(n12643) );
  XOR U12015 ( .A(n12652), .B(n12653), .Z(n12641) );
  AND U12016 ( .A(n1971), .B(n12654), .Z(n12653) );
  XOR U12017 ( .A(p_input[1603]), .B(n12652), .Z(n12654) );
  XOR U12018 ( .A(n12655), .B(n12656), .Z(n12652) );
  AND U12019 ( .A(n1975), .B(n12657), .Z(n12656) );
  IV U12020 ( .A(n12649), .Z(n12651) );
  XOR U12021 ( .A(n12658), .B(n12659), .Z(n12649) );
  AND U12022 ( .A(n1979), .B(n12660), .Z(n12659) );
  XOR U12023 ( .A(n12661), .B(n12662), .Z(n12647) );
  AND U12024 ( .A(n1983), .B(n12660), .Z(n12662) );
  XNOR U12025 ( .A(n12661), .B(n12658), .Z(n12660) );
  XOR U12026 ( .A(n12663), .B(n12664), .Z(n12658) );
  AND U12027 ( .A(n1986), .B(n12657), .Z(n12664) );
  XNOR U12028 ( .A(n12665), .B(n12655), .Z(n12657) );
  XOR U12029 ( .A(n12666), .B(n12667), .Z(n12655) );
  AND U12030 ( .A(n1990), .B(n12668), .Z(n12667) );
  XOR U12031 ( .A(p_input[1619]), .B(n12666), .Z(n12668) );
  XOR U12032 ( .A(n12669), .B(n12670), .Z(n12666) );
  AND U12033 ( .A(n1994), .B(n12671), .Z(n12670) );
  IV U12034 ( .A(n12663), .Z(n12665) );
  XOR U12035 ( .A(n12672), .B(n12673), .Z(n12663) );
  AND U12036 ( .A(n1998), .B(n12674), .Z(n12673) );
  XOR U12037 ( .A(n12675), .B(n12676), .Z(n12661) );
  AND U12038 ( .A(n2002), .B(n12674), .Z(n12676) );
  XNOR U12039 ( .A(n12675), .B(n12672), .Z(n12674) );
  XOR U12040 ( .A(n12677), .B(n12678), .Z(n12672) );
  AND U12041 ( .A(n2005), .B(n12671), .Z(n12678) );
  XNOR U12042 ( .A(n12679), .B(n12669), .Z(n12671) );
  XOR U12043 ( .A(n12680), .B(n12681), .Z(n12669) );
  AND U12044 ( .A(n2009), .B(n12682), .Z(n12681) );
  XOR U12045 ( .A(p_input[1635]), .B(n12680), .Z(n12682) );
  XOR U12046 ( .A(n12683), .B(n12684), .Z(n12680) );
  AND U12047 ( .A(n2013), .B(n12685), .Z(n12684) );
  IV U12048 ( .A(n12677), .Z(n12679) );
  XOR U12049 ( .A(n12686), .B(n12687), .Z(n12677) );
  AND U12050 ( .A(n2017), .B(n12688), .Z(n12687) );
  XOR U12051 ( .A(n12689), .B(n12690), .Z(n12675) );
  AND U12052 ( .A(n2021), .B(n12688), .Z(n12690) );
  XNOR U12053 ( .A(n12689), .B(n12686), .Z(n12688) );
  XOR U12054 ( .A(n12691), .B(n12692), .Z(n12686) );
  AND U12055 ( .A(n2024), .B(n12685), .Z(n12692) );
  XNOR U12056 ( .A(n12693), .B(n12683), .Z(n12685) );
  XOR U12057 ( .A(n12694), .B(n12695), .Z(n12683) );
  AND U12058 ( .A(n2028), .B(n12696), .Z(n12695) );
  XOR U12059 ( .A(p_input[1651]), .B(n12694), .Z(n12696) );
  XOR U12060 ( .A(n12697), .B(n12698), .Z(n12694) );
  AND U12061 ( .A(n2032), .B(n12699), .Z(n12698) );
  IV U12062 ( .A(n12691), .Z(n12693) );
  XOR U12063 ( .A(n12700), .B(n12701), .Z(n12691) );
  AND U12064 ( .A(n2036), .B(n12702), .Z(n12701) );
  XOR U12065 ( .A(n12703), .B(n12704), .Z(n12689) );
  AND U12066 ( .A(n2040), .B(n12702), .Z(n12704) );
  XNOR U12067 ( .A(n12703), .B(n12700), .Z(n12702) );
  XOR U12068 ( .A(n12705), .B(n12706), .Z(n12700) );
  AND U12069 ( .A(n2043), .B(n12699), .Z(n12706) );
  XNOR U12070 ( .A(n12707), .B(n12697), .Z(n12699) );
  XOR U12071 ( .A(n12708), .B(n12709), .Z(n12697) );
  AND U12072 ( .A(n2047), .B(n12710), .Z(n12709) );
  XOR U12073 ( .A(p_input[1667]), .B(n12708), .Z(n12710) );
  XOR U12074 ( .A(n12711), .B(n12712), .Z(n12708) );
  AND U12075 ( .A(n2051), .B(n12713), .Z(n12712) );
  IV U12076 ( .A(n12705), .Z(n12707) );
  XOR U12077 ( .A(n12714), .B(n12715), .Z(n12705) );
  AND U12078 ( .A(n2055), .B(n12716), .Z(n12715) );
  XOR U12079 ( .A(n12717), .B(n12718), .Z(n12703) );
  AND U12080 ( .A(n2059), .B(n12716), .Z(n12718) );
  XNOR U12081 ( .A(n12717), .B(n12714), .Z(n12716) );
  XOR U12082 ( .A(n12719), .B(n12720), .Z(n12714) );
  AND U12083 ( .A(n2062), .B(n12713), .Z(n12720) );
  XNOR U12084 ( .A(n12721), .B(n12711), .Z(n12713) );
  XOR U12085 ( .A(n12722), .B(n12723), .Z(n12711) );
  AND U12086 ( .A(n2066), .B(n12724), .Z(n12723) );
  XOR U12087 ( .A(p_input[1683]), .B(n12722), .Z(n12724) );
  XOR U12088 ( .A(n12725), .B(n12726), .Z(n12722) );
  AND U12089 ( .A(n2070), .B(n12727), .Z(n12726) );
  IV U12090 ( .A(n12719), .Z(n12721) );
  XOR U12091 ( .A(n12728), .B(n12729), .Z(n12719) );
  AND U12092 ( .A(n2074), .B(n12730), .Z(n12729) );
  XOR U12093 ( .A(n12731), .B(n12732), .Z(n12717) );
  AND U12094 ( .A(n2078), .B(n12730), .Z(n12732) );
  XNOR U12095 ( .A(n12731), .B(n12728), .Z(n12730) );
  XOR U12096 ( .A(n12733), .B(n12734), .Z(n12728) );
  AND U12097 ( .A(n2081), .B(n12727), .Z(n12734) );
  XNOR U12098 ( .A(n12735), .B(n12725), .Z(n12727) );
  XOR U12099 ( .A(n12736), .B(n12737), .Z(n12725) );
  AND U12100 ( .A(n2085), .B(n12738), .Z(n12737) );
  XOR U12101 ( .A(p_input[1699]), .B(n12736), .Z(n12738) );
  XOR U12102 ( .A(n12739), .B(n12740), .Z(n12736) );
  AND U12103 ( .A(n2089), .B(n12741), .Z(n12740) );
  IV U12104 ( .A(n12733), .Z(n12735) );
  XOR U12105 ( .A(n12742), .B(n12743), .Z(n12733) );
  AND U12106 ( .A(n2093), .B(n12744), .Z(n12743) );
  XOR U12107 ( .A(n12745), .B(n12746), .Z(n12731) );
  AND U12108 ( .A(n2097), .B(n12744), .Z(n12746) );
  XNOR U12109 ( .A(n12745), .B(n12742), .Z(n12744) );
  XOR U12110 ( .A(n12747), .B(n12748), .Z(n12742) );
  AND U12111 ( .A(n2100), .B(n12741), .Z(n12748) );
  XNOR U12112 ( .A(n12749), .B(n12739), .Z(n12741) );
  XOR U12113 ( .A(n12750), .B(n12751), .Z(n12739) );
  AND U12114 ( .A(n2104), .B(n12752), .Z(n12751) );
  XOR U12115 ( .A(p_input[1715]), .B(n12750), .Z(n12752) );
  XOR U12116 ( .A(n12753), .B(n12754), .Z(n12750) );
  AND U12117 ( .A(n2108), .B(n12755), .Z(n12754) );
  IV U12118 ( .A(n12747), .Z(n12749) );
  XOR U12119 ( .A(n12756), .B(n12757), .Z(n12747) );
  AND U12120 ( .A(n2112), .B(n12758), .Z(n12757) );
  XOR U12121 ( .A(n12759), .B(n12760), .Z(n12745) );
  AND U12122 ( .A(n2116), .B(n12758), .Z(n12760) );
  XNOR U12123 ( .A(n12759), .B(n12756), .Z(n12758) );
  XOR U12124 ( .A(n12761), .B(n12762), .Z(n12756) );
  AND U12125 ( .A(n2119), .B(n12755), .Z(n12762) );
  XNOR U12126 ( .A(n12763), .B(n12753), .Z(n12755) );
  XOR U12127 ( .A(n12764), .B(n12765), .Z(n12753) );
  AND U12128 ( .A(n2123), .B(n12766), .Z(n12765) );
  XOR U12129 ( .A(p_input[1731]), .B(n12764), .Z(n12766) );
  XOR U12130 ( .A(n12767), .B(n12768), .Z(n12764) );
  AND U12131 ( .A(n2127), .B(n12769), .Z(n12768) );
  IV U12132 ( .A(n12761), .Z(n12763) );
  XOR U12133 ( .A(n12770), .B(n12771), .Z(n12761) );
  AND U12134 ( .A(n2131), .B(n12772), .Z(n12771) );
  XOR U12135 ( .A(n12773), .B(n12774), .Z(n12759) );
  AND U12136 ( .A(n2135), .B(n12772), .Z(n12774) );
  XNOR U12137 ( .A(n12773), .B(n12770), .Z(n12772) );
  XOR U12138 ( .A(n12775), .B(n12776), .Z(n12770) );
  AND U12139 ( .A(n2138), .B(n12769), .Z(n12776) );
  XNOR U12140 ( .A(n12777), .B(n12767), .Z(n12769) );
  XOR U12141 ( .A(n12778), .B(n12779), .Z(n12767) );
  AND U12142 ( .A(n2142), .B(n12780), .Z(n12779) );
  XOR U12143 ( .A(p_input[1747]), .B(n12778), .Z(n12780) );
  XOR U12144 ( .A(n12781), .B(n12782), .Z(n12778) );
  AND U12145 ( .A(n2146), .B(n12783), .Z(n12782) );
  IV U12146 ( .A(n12775), .Z(n12777) );
  XOR U12147 ( .A(n12784), .B(n12785), .Z(n12775) );
  AND U12148 ( .A(n2150), .B(n12786), .Z(n12785) );
  XOR U12149 ( .A(n12787), .B(n12788), .Z(n12773) );
  AND U12150 ( .A(n2154), .B(n12786), .Z(n12788) );
  XNOR U12151 ( .A(n12787), .B(n12784), .Z(n12786) );
  XOR U12152 ( .A(n12789), .B(n12790), .Z(n12784) );
  AND U12153 ( .A(n2157), .B(n12783), .Z(n12790) );
  XNOR U12154 ( .A(n12791), .B(n12781), .Z(n12783) );
  XOR U12155 ( .A(n12792), .B(n12793), .Z(n12781) );
  AND U12156 ( .A(n2161), .B(n12794), .Z(n12793) );
  XOR U12157 ( .A(p_input[1763]), .B(n12792), .Z(n12794) );
  XOR U12158 ( .A(n12795), .B(n12796), .Z(n12792) );
  AND U12159 ( .A(n2165), .B(n12797), .Z(n12796) );
  IV U12160 ( .A(n12789), .Z(n12791) );
  XOR U12161 ( .A(n12798), .B(n12799), .Z(n12789) );
  AND U12162 ( .A(n2169), .B(n12800), .Z(n12799) );
  XOR U12163 ( .A(n12801), .B(n12802), .Z(n12787) );
  AND U12164 ( .A(n2173), .B(n12800), .Z(n12802) );
  XNOR U12165 ( .A(n12801), .B(n12798), .Z(n12800) );
  XOR U12166 ( .A(n12803), .B(n12804), .Z(n12798) );
  AND U12167 ( .A(n2176), .B(n12797), .Z(n12804) );
  XNOR U12168 ( .A(n12805), .B(n12795), .Z(n12797) );
  XOR U12169 ( .A(n12806), .B(n12807), .Z(n12795) );
  AND U12170 ( .A(n2180), .B(n12808), .Z(n12807) );
  XOR U12171 ( .A(p_input[1779]), .B(n12806), .Z(n12808) );
  XOR U12172 ( .A(n12809), .B(n12810), .Z(n12806) );
  AND U12173 ( .A(n2184), .B(n12811), .Z(n12810) );
  IV U12174 ( .A(n12803), .Z(n12805) );
  XOR U12175 ( .A(n12812), .B(n12813), .Z(n12803) );
  AND U12176 ( .A(n2188), .B(n12814), .Z(n12813) );
  XOR U12177 ( .A(n12815), .B(n12816), .Z(n12801) );
  AND U12178 ( .A(n2192), .B(n12814), .Z(n12816) );
  XNOR U12179 ( .A(n12815), .B(n12812), .Z(n12814) );
  XOR U12180 ( .A(n12817), .B(n12818), .Z(n12812) );
  AND U12181 ( .A(n2195), .B(n12811), .Z(n12818) );
  XNOR U12182 ( .A(n12819), .B(n12809), .Z(n12811) );
  XOR U12183 ( .A(n12820), .B(n12821), .Z(n12809) );
  AND U12184 ( .A(n2199), .B(n12822), .Z(n12821) );
  XOR U12185 ( .A(p_input[1795]), .B(n12820), .Z(n12822) );
  XOR U12186 ( .A(n12823), .B(n12824), .Z(n12820) );
  AND U12187 ( .A(n2203), .B(n12825), .Z(n12824) );
  IV U12188 ( .A(n12817), .Z(n12819) );
  XOR U12189 ( .A(n12826), .B(n12827), .Z(n12817) );
  AND U12190 ( .A(n2207), .B(n12828), .Z(n12827) );
  XOR U12191 ( .A(n12829), .B(n12830), .Z(n12815) );
  AND U12192 ( .A(n2211), .B(n12828), .Z(n12830) );
  XNOR U12193 ( .A(n12829), .B(n12826), .Z(n12828) );
  XOR U12194 ( .A(n12831), .B(n12832), .Z(n12826) );
  AND U12195 ( .A(n2214), .B(n12825), .Z(n12832) );
  XNOR U12196 ( .A(n12833), .B(n12823), .Z(n12825) );
  XOR U12197 ( .A(n12834), .B(n12835), .Z(n12823) );
  AND U12198 ( .A(n2218), .B(n12836), .Z(n12835) );
  XOR U12199 ( .A(p_input[1811]), .B(n12834), .Z(n12836) );
  XOR U12200 ( .A(n12837), .B(n12838), .Z(n12834) );
  AND U12201 ( .A(n2222), .B(n12839), .Z(n12838) );
  IV U12202 ( .A(n12831), .Z(n12833) );
  XOR U12203 ( .A(n12840), .B(n12841), .Z(n12831) );
  AND U12204 ( .A(n2226), .B(n12842), .Z(n12841) );
  XOR U12205 ( .A(n12843), .B(n12844), .Z(n12829) );
  AND U12206 ( .A(n2230), .B(n12842), .Z(n12844) );
  XNOR U12207 ( .A(n12843), .B(n12840), .Z(n12842) );
  XOR U12208 ( .A(n12845), .B(n12846), .Z(n12840) );
  AND U12209 ( .A(n2233), .B(n12839), .Z(n12846) );
  XNOR U12210 ( .A(n12847), .B(n12837), .Z(n12839) );
  XOR U12211 ( .A(n12848), .B(n12849), .Z(n12837) );
  AND U12212 ( .A(n2237), .B(n12850), .Z(n12849) );
  XOR U12213 ( .A(p_input[1827]), .B(n12848), .Z(n12850) );
  XOR U12214 ( .A(n12851), .B(n12852), .Z(n12848) );
  AND U12215 ( .A(n2241), .B(n12853), .Z(n12852) );
  IV U12216 ( .A(n12845), .Z(n12847) );
  XOR U12217 ( .A(n12854), .B(n12855), .Z(n12845) );
  AND U12218 ( .A(n2245), .B(n12856), .Z(n12855) );
  XOR U12219 ( .A(n12857), .B(n12858), .Z(n12843) );
  AND U12220 ( .A(n2249), .B(n12856), .Z(n12858) );
  XNOR U12221 ( .A(n12857), .B(n12854), .Z(n12856) );
  XOR U12222 ( .A(n12859), .B(n12860), .Z(n12854) );
  AND U12223 ( .A(n2252), .B(n12853), .Z(n12860) );
  XNOR U12224 ( .A(n12861), .B(n12851), .Z(n12853) );
  XOR U12225 ( .A(n12862), .B(n12863), .Z(n12851) );
  AND U12226 ( .A(n2256), .B(n12864), .Z(n12863) );
  XOR U12227 ( .A(p_input[1843]), .B(n12862), .Z(n12864) );
  XOR U12228 ( .A(n12865), .B(n12866), .Z(n12862) );
  AND U12229 ( .A(n2260), .B(n12867), .Z(n12866) );
  IV U12230 ( .A(n12859), .Z(n12861) );
  XOR U12231 ( .A(n12868), .B(n12869), .Z(n12859) );
  AND U12232 ( .A(n2264), .B(n12870), .Z(n12869) );
  XOR U12233 ( .A(n12871), .B(n12872), .Z(n12857) );
  AND U12234 ( .A(n2268), .B(n12870), .Z(n12872) );
  XNOR U12235 ( .A(n12871), .B(n12868), .Z(n12870) );
  XOR U12236 ( .A(n12873), .B(n12874), .Z(n12868) );
  AND U12237 ( .A(n2271), .B(n12867), .Z(n12874) );
  XNOR U12238 ( .A(n12875), .B(n12865), .Z(n12867) );
  XOR U12239 ( .A(n12876), .B(n12877), .Z(n12865) );
  AND U12240 ( .A(n2275), .B(n12878), .Z(n12877) );
  XOR U12241 ( .A(p_input[1859]), .B(n12876), .Z(n12878) );
  XOR U12242 ( .A(n12879), .B(n12880), .Z(n12876) );
  AND U12243 ( .A(n2279), .B(n12881), .Z(n12880) );
  IV U12244 ( .A(n12873), .Z(n12875) );
  XOR U12245 ( .A(n12882), .B(n12883), .Z(n12873) );
  AND U12246 ( .A(n2283), .B(n12884), .Z(n12883) );
  XOR U12247 ( .A(n12885), .B(n12886), .Z(n12871) );
  AND U12248 ( .A(n2287), .B(n12884), .Z(n12886) );
  XNOR U12249 ( .A(n12885), .B(n12882), .Z(n12884) );
  XOR U12250 ( .A(n12887), .B(n12888), .Z(n12882) );
  AND U12251 ( .A(n2290), .B(n12881), .Z(n12888) );
  XNOR U12252 ( .A(n12889), .B(n12879), .Z(n12881) );
  XOR U12253 ( .A(n12890), .B(n12891), .Z(n12879) );
  AND U12254 ( .A(n2294), .B(n12892), .Z(n12891) );
  XOR U12255 ( .A(p_input[1875]), .B(n12890), .Z(n12892) );
  XOR U12256 ( .A(n12893), .B(n12894), .Z(n12890) );
  AND U12257 ( .A(n2298), .B(n12895), .Z(n12894) );
  IV U12258 ( .A(n12887), .Z(n12889) );
  XOR U12259 ( .A(n12896), .B(n12897), .Z(n12887) );
  AND U12260 ( .A(n2302), .B(n12898), .Z(n12897) );
  XOR U12261 ( .A(n12899), .B(n12900), .Z(n12885) );
  AND U12262 ( .A(n2306), .B(n12898), .Z(n12900) );
  XNOR U12263 ( .A(n12899), .B(n12896), .Z(n12898) );
  XOR U12264 ( .A(n12901), .B(n12902), .Z(n12896) );
  AND U12265 ( .A(n2309), .B(n12895), .Z(n12902) );
  XNOR U12266 ( .A(n12903), .B(n12893), .Z(n12895) );
  XOR U12267 ( .A(n12904), .B(n12905), .Z(n12893) );
  AND U12268 ( .A(n2313), .B(n12906), .Z(n12905) );
  XOR U12269 ( .A(p_input[1891]), .B(n12904), .Z(n12906) );
  XOR U12270 ( .A(n12907), .B(n12908), .Z(n12904) );
  AND U12271 ( .A(n2317), .B(n12909), .Z(n12908) );
  IV U12272 ( .A(n12901), .Z(n12903) );
  XOR U12273 ( .A(n12910), .B(n12911), .Z(n12901) );
  AND U12274 ( .A(n2321), .B(n12912), .Z(n12911) );
  XOR U12275 ( .A(n12913), .B(n12914), .Z(n12899) );
  AND U12276 ( .A(n2325), .B(n12912), .Z(n12914) );
  XNOR U12277 ( .A(n12913), .B(n12910), .Z(n12912) );
  XOR U12278 ( .A(n12915), .B(n12916), .Z(n12910) );
  AND U12279 ( .A(n2328), .B(n12909), .Z(n12916) );
  XNOR U12280 ( .A(n12917), .B(n12907), .Z(n12909) );
  XOR U12281 ( .A(n12918), .B(n12919), .Z(n12907) );
  AND U12282 ( .A(n2332), .B(n12920), .Z(n12919) );
  XOR U12283 ( .A(p_input[1907]), .B(n12918), .Z(n12920) );
  XOR U12284 ( .A(n12921), .B(n12922), .Z(n12918) );
  AND U12285 ( .A(n2336), .B(n12923), .Z(n12922) );
  IV U12286 ( .A(n12915), .Z(n12917) );
  XOR U12287 ( .A(n12924), .B(n12925), .Z(n12915) );
  AND U12288 ( .A(n2340), .B(n12926), .Z(n12925) );
  XOR U12289 ( .A(n12927), .B(n12928), .Z(n12913) );
  AND U12290 ( .A(n2344), .B(n12926), .Z(n12928) );
  XNOR U12291 ( .A(n12927), .B(n12924), .Z(n12926) );
  XOR U12292 ( .A(n12929), .B(n12930), .Z(n12924) );
  AND U12293 ( .A(n2347), .B(n12923), .Z(n12930) );
  XNOR U12294 ( .A(n12931), .B(n12921), .Z(n12923) );
  XOR U12295 ( .A(n12932), .B(n12933), .Z(n12921) );
  AND U12296 ( .A(n2351), .B(n12934), .Z(n12933) );
  XOR U12297 ( .A(p_input[1923]), .B(n12932), .Z(n12934) );
  XOR U12298 ( .A(n12935), .B(n12936), .Z(n12932) );
  AND U12299 ( .A(n2355), .B(n12937), .Z(n12936) );
  IV U12300 ( .A(n12929), .Z(n12931) );
  XOR U12301 ( .A(n12938), .B(n12939), .Z(n12929) );
  AND U12302 ( .A(n2359), .B(n12940), .Z(n12939) );
  XOR U12303 ( .A(n12941), .B(n12942), .Z(n12927) );
  AND U12304 ( .A(n2363), .B(n12940), .Z(n12942) );
  XNOR U12305 ( .A(n12941), .B(n12938), .Z(n12940) );
  XOR U12306 ( .A(n12943), .B(n12944), .Z(n12938) );
  AND U12307 ( .A(n2366), .B(n12937), .Z(n12944) );
  XNOR U12308 ( .A(n12945), .B(n12935), .Z(n12937) );
  XOR U12309 ( .A(n12946), .B(n12947), .Z(n12935) );
  AND U12310 ( .A(n2370), .B(n12948), .Z(n12947) );
  XOR U12311 ( .A(p_input[1939]), .B(n12946), .Z(n12948) );
  XOR U12312 ( .A(n12949), .B(n12950), .Z(n12946) );
  AND U12313 ( .A(n2374), .B(n12951), .Z(n12950) );
  IV U12314 ( .A(n12943), .Z(n12945) );
  XOR U12315 ( .A(n12952), .B(n12953), .Z(n12943) );
  AND U12316 ( .A(n2378), .B(n12954), .Z(n12953) );
  XOR U12317 ( .A(n12955), .B(n12956), .Z(n12941) );
  AND U12318 ( .A(n2382), .B(n12954), .Z(n12956) );
  XNOR U12319 ( .A(n12955), .B(n12952), .Z(n12954) );
  XOR U12320 ( .A(n12957), .B(n12958), .Z(n12952) );
  AND U12321 ( .A(n2385), .B(n12951), .Z(n12958) );
  XNOR U12322 ( .A(n12959), .B(n12949), .Z(n12951) );
  XOR U12323 ( .A(n12960), .B(n12961), .Z(n12949) );
  AND U12324 ( .A(n2389), .B(n12962), .Z(n12961) );
  XOR U12325 ( .A(p_input[1955]), .B(n12960), .Z(n12962) );
  XOR U12326 ( .A(n12963), .B(n12964), .Z(n12960) );
  AND U12327 ( .A(n2393), .B(n12965), .Z(n12964) );
  IV U12328 ( .A(n12957), .Z(n12959) );
  XOR U12329 ( .A(n12966), .B(n12967), .Z(n12957) );
  AND U12330 ( .A(n2397), .B(n12968), .Z(n12967) );
  XOR U12331 ( .A(n12969), .B(n12970), .Z(n12955) );
  AND U12332 ( .A(n2401), .B(n12968), .Z(n12970) );
  XNOR U12333 ( .A(n12969), .B(n12966), .Z(n12968) );
  XOR U12334 ( .A(n12971), .B(n12972), .Z(n12966) );
  AND U12335 ( .A(n2404), .B(n12965), .Z(n12972) );
  XNOR U12336 ( .A(n12973), .B(n12963), .Z(n12965) );
  XOR U12337 ( .A(n12974), .B(n12975), .Z(n12963) );
  AND U12338 ( .A(n2408), .B(n12976), .Z(n12975) );
  XOR U12339 ( .A(p_input[1971]), .B(n12974), .Z(n12976) );
  XOR U12340 ( .A(n12977), .B(n12978), .Z(n12974) );
  AND U12341 ( .A(n2412), .B(n12979), .Z(n12978) );
  IV U12342 ( .A(n12971), .Z(n12973) );
  XOR U12343 ( .A(n12980), .B(n12981), .Z(n12971) );
  AND U12344 ( .A(n2416), .B(n12982), .Z(n12981) );
  XOR U12345 ( .A(n12983), .B(n12984), .Z(n12969) );
  AND U12346 ( .A(n2420), .B(n12982), .Z(n12984) );
  XNOR U12347 ( .A(n12983), .B(n12980), .Z(n12982) );
  XOR U12348 ( .A(n12985), .B(n12986), .Z(n12980) );
  AND U12349 ( .A(n2423), .B(n12979), .Z(n12986) );
  XNOR U12350 ( .A(n12987), .B(n12977), .Z(n12979) );
  XOR U12351 ( .A(n12988), .B(n12989), .Z(n12977) );
  AND U12352 ( .A(n2427), .B(n12990), .Z(n12989) );
  XOR U12353 ( .A(p_input[1987]), .B(n12988), .Z(n12990) );
  XOR U12354 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n12991), 
        .Z(n12988) );
  AND U12355 ( .A(n2430), .B(n12992), .Z(n12991) );
  IV U12356 ( .A(n12985), .Z(n12987) );
  XOR U12357 ( .A(n12993), .B(n12994), .Z(n12985) );
  AND U12358 ( .A(n2434), .B(n12995), .Z(n12994) );
  XOR U12359 ( .A(n12996), .B(n12997), .Z(n12983) );
  AND U12360 ( .A(n2438), .B(n12995), .Z(n12997) );
  XNOR U12361 ( .A(n12996), .B(n12993), .Z(n12995) );
  XNOR U12362 ( .A(n12998), .B(n12999), .Z(n12993) );
  AND U12363 ( .A(n2441), .B(n12992), .Z(n12999) );
  XNOR U12364 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n12998), 
        .Z(n12992) );
  XNOR U12365 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n13000), 
        .Z(n12998) );
  AND U12366 ( .A(n2443), .B(n13001), .Z(n13000) );
  XNOR U12367 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n13002), .Z(n12996) );
  AND U12368 ( .A(n2446), .B(n13001), .Z(n13002) );
  XOR U12369 ( .A(n13003), .B(n13004), .Z(n13001) );
  XOR U12370 ( .A(n51), .B(n13005), .Z(o[18]) );
  AND U12371 ( .A(n62), .B(n13006), .Z(n51) );
  XOR U12372 ( .A(n52), .B(n13005), .Z(n13006) );
  XOR U12373 ( .A(n13007), .B(n41), .Z(n13005) );
  AND U12374 ( .A(n65), .B(n13008), .Z(n41) );
  XOR U12375 ( .A(n42), .B(n13007), .Z(n13008) );
  XOR U12376 ( .A(n13009), .B(n13010), .Z(n42) );
  AND U12377 ( .A(n70), .B(n13011), .Z(n13010) );
  XOR U12378 ( .A(p_input[2]), .B(n13009), .Z(n13011) );
  XNOR U12379 ( .A(n13012), .B(n13013), .Z(n13009) );
  AND U12380 ( .A(n74), .B(n13014), .Z(n13013) );
  XOR U12381 ( .A(n13015), .B(n13016), .Z(n13007) );
  AND U12382 ( .A(n78), .B(n13017), .Z(n13016) );
  XOR U12383 ( .A(n13018), .B(n13019), .Z(n52) );
  AND U12384 ( .A(n82), .B(n13017), .Z(n13019) );
  XNOR U12385 ( .A(n13020), .B(n13018), .Z(n13017) );
  IV U12386 ( .A(n13015), .Z(n13020) );
  XOR U12387 ( .A(n13021), .B(n13022), .Z(n13015) );
  AND U12388 ( .A(n86), .B(n13014), .Z(n13022) );
  XNOR U12389 ( .A(n13012), .B(n13021), .Z(n13014) );
  XNOR U12390 ( .A(n13023), .B(n13024), .Z(n13012) );
  AND U12391 ( .A(n90), .B(n13025), .Z(n13024) );
  XOR U12392 ( .A(p_input[18]), .B(n13023), .Z(n13025) );
  XNOR U12393 ( .A(n13026), .B(n13027), .Z(n13023) );
  AND U12394 ( .A(n94), .B(n13028), .Z(n13027) );
  XOR U12395 ( .A(n13029), .B(n13030), .Z(n13021) );
  AND U12396 ( .A(n98), .B(n13031), .Z(n13030) );
  XOR U12397 ( .A(n13032), .B(n13033), .Z(n13018) );
  AND U12398 ( .A(n102), .B(n13031), .Z(n13033) );
  XNOR U12399 ( .A(n13034), .B(n13032), .Z(n13031) );
  IV U12400 ( .A(n13029), .Z(n13034) );
  XOR U12401 ( .A(n13035), .B(n13036), .Z(n13029) );
  AND U12402 ( .A(n105), .B(n13028), .Z(n13036) );
  XNOR U12403 ( .A(n13026), .B(n13035), .Z(n13028) );
  XNOR U12404 ( .A(n13037), .B(n13038), .Z(n13026) );
  AND U12405 ( .A(n109), .B(n13039), .Z(n13038) );
  XOR U12406 ( .A(p_input[34]), .B(n13037), .Z(n13039) );
  XNOR U12407 ( .A(n13040), .B(n13041), .Z(n13037) );
  AND U12408 ( .A(n113), .B(n13042), .Z(n13041) );
  XOR U12409 ( .A(n13043), .B(n13044), .Z(n13035) );
  AND U12410 ( .A(n117), .B(n13045), .Z(n13044) );
  XOR U12411 ( .A(n13046), .B(n13047), .Z(n13032) );
  AND U12412 ( .A(n121), .B(n13045), .Z(n13047) );
  XNOR U12413 ( .A(n13048), .B(n13046), .Z(n13045) );
  IV U12414 ( .A(n13043), .Z(n13048) );
  XOR U12415 ( .A(n13049), .B(n13050), .Z(n13043) );
  AND U12416 ( .A(n124), .B(n13042), .Z(n13050) );
  XNOR U12417 ( .A(n13040), .B(n13049), .Z(n13042) );
  XNOR U12418 ( .A(n13051), .B(n13052), .Z(n13040) );
  AND U12419 ( .A(n128), .B(n13053), .Z(n13052) );
  XOR U12420 ( .A(p_input[50]), .B(n13051), .Z(n13053) );
  XNOR U12421 ( .A(n13054), .B(n13055), .Z(n13051) );
  AND U12422 ( .A(n132), .B(n13056), .Z(n13055) );
  XOR U12423 ( .A(n13057), .B(n13058), .Z(n13049) );
  AND U12424 ( .A(n136), .B(n13059), .Z(n13058) );
  XOR U12425 ( .A(n13060), .B(n13061), .Z(n13046) );
  AND U12426 ( .A(n140), .B(n13059), .Z(n13061) );
  XNOR U12427 ( .A(n13062), .B(n13060), .Z(n13059) );
  IV U12428 ( .A(n13057), .Z(n13062) );
  XOR U12429 ( .A(n13063), .B(n13064), .Z(n13057) );
  AND U12430 ( .A(n143), .B(n13056), .Z(n13064) );
  XNOR U12431 ( .A(n13054), .B(n13063), .Z(n13056) );
  XNOR U12432 ( .A(n13065), .B(n13066), .Z(n13054) );
  AND U12433 ( .A(n147), .B(n13067), .Z(n13066) );
  XOR U12434 ( .A(p_input[66]), .B(n13065), .Z(n13067) );
  XNOR U12435 ( .A(n13068), .B(n13069), .Z(n13065) );
  AND U12436 ( .A(n151), .B(n13070), .Z(n13069) );
  XOR U12437 ( .A(n13071), .B(n13072), .Z(n13063) );
  AND U12438 ( .A(n155), .B(n13073), .Z(n13072) );
  XOR U12439 ( .A(n13074), .B(n13075), .Z(n13060) );
  AND U12440 ( .A(n159), .B(n13073), .Z(n13075) );
  XNOR U12441 ( .A(n13076), .B(n13074), .Z(n13073) );
  IV U12442 ( .A(n13071), .Z(n13076) );
  XOR U12443 ( .A(n13077), .B(n13078), .Z(n13071) );
  AND U12444 ( .A(n162), .B(n13070), .Z(n13078) );
  XNOR U12445 ( .A(n13068), .B(n13077), .Z(n13070) );
  XNOR U12446 ( .A(n13079), .B(n13080), .Z(n13068) );
  AND U12447 ( .A(n166), .B(n13081), .Z(n13080) );
  XOR U12448 ( .A(p_input[82]), .B(n13079), .Z(n13081) );
  XNOR U12449 ( .A(n13082), .B(n13083), .Z(n13079) );
  AND U12450 ( .A(n170), .B(n13084), .Z(n13083) );
  XOR U12451 ( .A(n13085), .B(n13086), .Z(n13077) );
  AND U12452 ( .A(n174), .B(n13087), .Z(n13086) );
  XOR U12453 ( .A(n13088), .B(n13089), .Z(n13074) );
  AND U12454 ( .A(n178), .B(n13087), .Z(n13089) );
  XNOR U12455 ( .A(n13090), .B(n13088), .Z(n13087) );
  IV U12456 ( .A(n13085), .Z(n13090) );
  XOR U12457 ( .A(n13091), .B(n13092), .Z(n13085) );
  AND U12458 ( .A(n181), .B(n13084), .Z(n13092) );
  XNOR U12459 ( .A(n13082), .B(n13091), .Z(n13084) );
  XNOR U12460 ( .A(n13093), .B(n13094), .Z(n13082) );
  AND U12461 ( .A(n185), .B(n13095), .Z(n13094) );
  XOR U12462 ( .A(p_input[98]), .B(n13093), .Z(n13095) );
  XNOR U12463 ( .A(n13096), .B(n13097), .Z(n13093) );
  AND U12464 ( .A(n189), .B(n13098), .Z(n13097) );
  XOR U12465 ( .A(n13099), .B(n13100), .Z(n13091) );
  AND U12466 ( .A(n193), .B(n13101), .Z(n13100) );
  XOR U12467 ( .A(n13102), .B(n13103), .Z(n13088) );
  AND U12468 ( .A(n197), .B(n13101), .Z(n13103) );
  XNOR U12469 ( .A(n13104), .B(n13102), .Z(n13101) );
  IV U12470 ( .A(n13099), .Z(n13104) );
  XOR U12471 ( .A(n13105), .B(n13106), .Z(n13099) );
  AND U12472 ( .A(n200), .B(n13098), .Z(n13106) );
  XNOR U12473 ( .A(n13096), .B(n13105), .Z(n13098) );
  XNOR U12474 ( .A(n13107), .B(n13108), .Z(n13096) );
  AND U12475 ( .A(n204), .B(n13109), .Z(n13108) );
  XOR U12476 ( .A(p_input[114]), .B(n13107), .Z(n13109) );
  XNOR U12477 ( .A(n13110), .B(n13111), .Z(n13107) );
  AND U12478 ( .A(n208), .B(n13112), .Z(n13111) );
  XOR U12479 ( .A(n13113), .B(n13114), .Z(n13105) );
  AND U12480 ( .A(n212), .B(n13115), .Z(n13114) );
  XOR U12481 ( .A(n13116), .B(n13117), .Z(n13102) );
  AND U12482 ( .A(n216), .B(n13115), .Z(n13117) );
  XNOR U12483 ( .A(n13118), .B(n13116), .Z(n13115) );
  IV U12484 ( .A(n13113), .Z(n13118) );
  XOR U12485 ( .A(n13119), .B(n13120), .Z(n13113) );
  AND U12486 ( .A(n219), .B(n13112), .Z(n13120) );
  XNOR U12487 ( .A(n13110), .B(n13119), .Z(n13112) );
  XNOR U12488 ( .A(n13121), .B(n13122), .Z(n13110) );
  AND U12489 ( .A(n223), .B(n13123), .Z(n13122) );
  XOR U12490 ( .A(p_input[130]), .B(n13121), .Z(n13123) );
  XNOR U12491 ( .A(n13124), .B(n13125), .Z(n13121) );
  AND U12492 ( .A(n227), .B(n13126), .Z(n13125) );
  XOR U12493 ( .A(n13127), .B(n13128), .Z(n13119) );
  AND U12494 ( .A(n231), .B(n13129), .Z(n13128) );
  XOR U12495 ( .A(n13130), .B(n13131), .Z(n13116) );
  AND U12496 ( .A(n235), .B(n13129), .Z(n13131) );
  XNOR U12497 ( .A(n13132), .B(n13130), .Z(n13129) );
  IV U12498 ( .A(n13127), .Z(n13132) );
  XOR U12499 ( .A(n13133), .B(n13134), .Z(n13127) );
  AND U12500 ( .A(n238), .B(n13126), .Z(n13134) );
  XNOR U12501 ( .A(n13124), .B(n13133), .Z(n13126) );
  XNOR U12502 ( .A(n13135), .B(n13136), .Z(n13124) );
  AND U12503 ( .A(n242), .B(n13137), .Z(n13136) );
  XOR U12504 ( .A(p_input[146]), .B(n13135), .Z(n13137) );
  XNOR U12505 ( .A(n13138), .B(n13139), .Z(n13135) );
  AND U12506 ( .A(n246), .B(n13140), .Z(n13139) );
  XOR U12507 ( .A(n13141), .B(n13142), .Z(n13133) );
  AND U12508 ( .A(n250), .B(n13143), .Z(n13142) );
  XOR U12509 ( .A(n13144), .B(n13145), .Z(n13130) );
  AND U12510 ( .A(n254), .B(n13143), .Z(n13145) );
  XNOR U12511 ( .A(n13146), .B(n13144), .Z(n13143) );
  IV U12512 ( .A(n13141), .Z(n13146) );
  XOR U12513 ( .A(n13147), .B(n13148), .Z(n13141) );
  AND U12514 ( .A(n257), .B(n13140), .Z(n13148) );
  XNOR U12515 ( .A(n13138), .B(n13147), .Z(n13140) );
  XNOR U12516 ( .A(n13149), .B(n13150), .Z(n13138) );
  AND U12517 ( .A(n261), .B(n13151), .Z(n13150) );
  XOR U12518 ( .A(p_input[162]), .B(n13149), .Z(n13151) );
  XNOR U12519 ( .A(n13152), .B(n13153), .Z(n13149) );
  AND U12520 ( .A(n265), .B(n13154), .Z(n13153) );
  XOR U12521 ( .A(n13155), .B(n13156), .Z(n13147) );
  AND U12522 ( .A(n269), .B(n13157), .Z(n13156) );
  XOR U12523 ( .A(n13158), .B(n13159), .Z(n13144) );
  AND U12524 ( .A(n273), .B(n13157), .Z(n13159) );
  XNOR U12525 ( .A(n13160), .B(n13158), .Z(n13157) );
  IV U12526 ( .A(n13155), .Z(n13160) );
  XOR U12527 ( .A(n13161), .B(n13162), .Z(n13155) );
  AND U12528 ( .A(n276), .B(n13154), .Z(n13162) );
  XNOR U12529 ( .A(n13152), .B(n13161), .Z(n13154) );
  XNOR U12530 ( .A(n13163), .B(n13164), .Z(n13152) );
  AND U12531 ( .A(n280), .B(n13165), .Z(n13164) );
  XOR U12532 ( .A(p_input[178]), .B(n13163), .Z(n13165) );
  XNOR U12533 ( .A(n13166), .B(n13167), .Z(n13163) );
  AND U12534 ( .A(n284), .B(n13168), .Z(n13167) );
  XOR U12535 ( .A(n13169), .B(n13170), .Z(n13161) );
  AND U12536 ( .A(n288), .B(n13171), .Z(n13170) );
  XOR U12537 ( .A(n13172), .B(n13173), .Z(n13158) );
  AND U12538 ( .A(n292), .B(n13171), .Z(n13173) );
  XNOR U12539 ( .A(n13174), .B(n13172), .Z(n13171) );
  IV U12540 ( .A(n13169), .Z(n13174) );
  XOR U12541 ( .A(n13175), .B(n13176), .Z(n13169) );
  AND U12542 ( .A(n295), .B(n13168), .Z(n13176) );
  XNOR U12543 ( .A(n13166), .B(n13175), .Z(n13168) );
  XNOR U12544 ( .A(n13177), .B(n13178), .Z(n13166) );
  AND U12545 ( .A(n299), .B(n13179), .Z(n13178) );
  XOR U12546 ( .A(p_input[194]), .B(n13177), .Z(n13179) );
  XNOR U12547 ( .A(n13180), .B(n13181), .Z(n13177) );
  AND U12548 ( .A(n303), .B(n13182), .Z(n13181) );
  XOR U12549 ( .A(n13183), .B(n13184), .Z(n13175) );
  AND U12550 ( .A(n307), .B(n13185), .Z(n13184) );
  XOR U12551 ( .A(n13186), .B(n13187), .Z(n13172) );
  AND U12552 ( .A(n311), .B(n13185), .Z(n13187) );
  XNOR U12553 ( .A(n13188), .B(n13186), .Z(n13185) );
  IV U12554 ( .A(n13183), .Z(n13188) );
  XOR U12555 ( .A(n13189), .B(n13190), .Z(n13183) );
  AND U12556 ( .A(n314), .B(n13182), .Z(n13190) );
  XNOR U12557 ( .A(n13180), .B(n13189), .Z(n13182) );
  XNOR U12558 ( .A(n13191), .B(n13192), .Z(n13180) );
  AND U12559 ( .A(n318), .B(n13193), .Z(n13192) );
  XOR U12560 ( .A(p_input[210]), .B(n13191), .Z(n13193) );
  XNOR U12561 ( .A(n13194), .B(n13195), .Z(n13191) );
  AND U12562 ( .A(n322), .B(n13196), .Z(n13195) );
  XOR U12563 ( .A(n13197), .B(n13198), .Z(n13189) );
  AND U12564 ( .A(n326), .B(n13199), .Z(n13198) );
  XOR U12565 ( .A(n13200), .B(n13201), .Z(n13186) );
  AND U12566 ( .A(n330), .B(n13199), .Z(n13201) );
  XNOR U12567 ( .A(n13202), .B(n13200), .Z(n13199) );
  IV U12568 ( .A(n13197), .Z(n13202) );
  XOR U12569 ( .A(n13203), .B(n13204), .Z(n13197) );
  AND U12570 ( .A(n333), .B(n13196), .Z(n13204) );
  XNOR U12571 ( .A(n13194), .B(n13203), .Z(n13196) );
  XNOR U12572 ( .A(n13205), .B(n13206), .Z(n13194) );
  AND U12573 ( .A(n337), .B(n13207), .Z(n13206) );
  XOR U12574 ( .A(p_input[226]), .B(n13205), .Z(n13207) );
  XNOR U12575 ( .A(n13208), .B(n13209), .Z(n13205) );
  AND U12576 ( .A(n341), .B(n13210), .Z(n13209) );
  XOR U12577 ( .A(n13211), .B(n13212), .Z(n13203) );
  AND U12578 ( .A(n345), .B(n13213), .Z(n13212) );
  XOR U12579 ( .A(n13214), .B(n13215), .Z(n13200) );
  AND U12580 ( .A(n349), .B(n13213), .Z(n13215) );
  XNOR U12581 ( .A(n13216), .B(n13214), .Z(n13213) );
  IV U12582 ( .A(n13211), .Z(n13216) );
  XOR U12583 ( .A(n13217), .B(n13218), .Z(n13211) );
  AND U12584 ( .A(n352), .B(n13210), .Z(n13218) );
  XNOR U12585 ( .A(n13208), .B(n13217), .Z(n13210) );
  XNOR U12586 ( .A(n13219), .B(n13220), .Z(n13208) );
  AND U12587 ( .A(n356), .B(n13221), .Z(n13220) );
  XOR U12588 ( .A(p_input[242]), .B(n13219), .Z(n13221) );
  XNOR U12589 ( .A(n13222), .B(n13223), .Z(n13219) );
  AND U12590 ( .A(n360), .B(n13224), .Z(n13223) );
  XOR U12591 ( .A(n13225), .B(n13226), .Z(n13217) );
  AND U12592 ( .A(n364), .B(n13227), .Z(n13226) );
  XOR U12593 ( .A(n13228), .B(n13229), .Z(n13214) );
  AND U12594 ( .A(n368), .B(n13227), .Z(n13229) );
  XNOR U12595 ( .A(n13230), .B(n13228), .Z(n13227) );
  IV U12596 ( .A(n13225), .Z(n13230) );
  XOR U12597 ( .A(n13231), .B(n13232), .Z(n13225) );
  AND U12598 ( .A(n371), .B(n13224), .Z(n13232) );
  XNOR U12599 ( .A(n13222), .B(n13231), .Z(n13224) );
  XNOR U12600 ( .A(n13233), .B(n13234), .Z(n13222) );
  AND U12601 ( .A(n375), .B(n13235), .Z(n13234) );
  XOR U12602 ( .A(p_input[258]), .B(n13233), .Z(n13235) );
  XNOR U12603 ( .A(n13236), .B(n13237), .Z(n13233) );
  AND U12604 ( .A(n379), .B(n13238), .Z(n13237) );
  XOR U12605 ( .A(n13239), .B(n13240), .Z(n13231) );
  AND U12606 ( .A(n383), .B(n13241), .Z(n13240) );
  XOR U12607 ( .A(n13242), .B(n13243), .Z(n13228) );
  AND U12608 ( .A(n387), .B(n13241), .Z(n13243) );
  XNOR U12609 ( .A(n13244), .B(n13242), .Z(n13241) );
  IV U12610 ( .A(n13239), .Z(n13244) );
  XOR U12611 ( .A(n13245), .B(n13246), .Z(n13239) );
  AND U12612 ( .A(n390), .B(n13238), .Z(n13246) );
  XNOR U12613 ( .A(n13236), .B(n13245), .Z(n13238) );
  XNOR U12614 ( .A(n13247), .B(n13248), .Z(n13236) );
  AND U12615 ( .A(n394), .B(n13249), .Z(n13248) );
  XOR U12616 ( .A(p_input[274]), .B(n13247), .Z(n13249) );
  XNOR U12617 ( .A(n13250), .B(n13251), .Z(n13247) );
  AND U12618 ( .A(n398), .B(n13252), .Z(n13251) );
  XOR U12619 ( .A(n13253), .B(n13254), .Z(n13245) );
  AND U12620 ( .A(n402), .B(n13255), .Z(n13254) );
  XOR U12621 ( .A(n13256), .B(n13257), .Z(n13242) );
  AND U12622 ( .A(n406), .B(n13255), .Z(n13257) );
  XNOR U12623 ( .A(n13258), .B(n13256), .Z(n13255) );
  IV U12624 ( .A(n13253), .Z(n13258) );
  XOR U12625 ( .A(n13259), .B(n13260), .Z(n13253) );
  AND U12626 ( .A(n409), .B(n13252), .Z(n13260) );
  XNOR U12627 ( .A(n13250), .B(n13259), .Z(n13252) );
  XNOR U12628 ( .A(n13261), .B(n13262), .Z(n13250) );
  AND U12629 ( .A(n413), .B(n13263), .Z(n13262) );
  XOR U12630 ( .A(p_input[290]), .B(n13261), .Z(n13263) );
  XNOR U12631 ( .A(n13264), .B(n13265), .Z(n13261) );
  AND U12632 ( .A(n417), .B(n13266), .Z(n13265) );
  XOR U12633 ( .A(n13267), .B(n13268), .Z(n13259) );
  AND U12634 ( .A(n421), .B(n13269), .Z(n13268) );
  XOR U12635 ( .A(n13270), .B(n13271), .Z(n13256) );
  AND U12636 ( .A(n425), .B(n13269), .Z(n13271) );
  XNOR U12637 ( .A(n13272), .B(n13270), .Z(n13269) );
  IV U12638 ( .A(n13267), .Z(n13272) );
  XOR U12639 ( .A(n13273), .B(n13274), .Z(n13267) );
  AND U12640 ( .A(n428), .B(n13266), .Z(n13274) );
  XNOR U12641 ( .A(n13264), .B(n13273), .Z(n13266) );
  XNOR U12642 ( .A(n13275), .B(n13276), .Z(n13264) );
  AND U12643 ( .A(n432), .B(n13277), .Z(n13276) );
  XOR U12644 ( .A(p_input[306]), .B(n13275), .Z(n13277) );
  XNOR U12645 ( .A(n13278), .B(n13279), .Z(n13275) );
  AND U12646 ( .A(n436), .B(n13280), .Z(n13279) );
  XOR U12647 ( .A(n13281), .B(n13282), .Z(n13273) );
  AND U12648 ( .A(n440), .B(n13283), .Z(n13282) );
  XOR U12649 ( .A(n13284), .B(n13285), .Z(n13270) );
  AND U12650 ( .A(n444), .B(n13283), .Z(n13285) );
  XNOR U12651 ( .A(n13286), .B(n13284), .Z(n13283) );
  IV U12652 ( .A(n13281), .Z(n13286) );
  XOR U12653 ( .A(n13287), .B(n13288), .Z(n13281) );
  AND U12654 ( .A(n447), .B(n13280), .Z(n13288) );
  XNOR U12655 ( .A(n13278), .B(n13287), .Z(n13280) );
  XNOR U12656 ( .A(n13289), .B(n13290), .Z(n13278) );
  AND U12657 ( .A(n451), .B(n13291), .Z(n13290) );
  XOR U12658 ( .A(p_input[322]), .B(n13289), .Z(n13291) );
  XNOR U12659 ( .A(n13292), .B(n13293), .Z(n13289) );
  AND U12660 ( .A(n455), .B(n13294), .Z(n13293) );
  XOR U12661 ( .A(n13295), .B(n13296), .Z(n13287) );
  AND U12662 ( .A(n459), .B(n13297), .Z(n13296) );
  XOR U12663 ( .A(n13298), .B(n13299), .Z(n13284) );
  AND U12664 ( .A(n463), .B(n13297), .Z(n13299) );
  XNOR U12665 ( .A(n13300), .B(n13298), .Z(n13297) );
  IV U12666 ( .A(n13295), .Z(n13300) );
  XOR U12667 ( .A(n13301), .B(n13302), .Z(n13295) );
  AND U12668 ( .A(n466), .B(n13294), .Z(n13302) );
  XNOR U12669 ( .A(n13292), .B(n13301), .Z(n13294) );
  XNOR U12670 ( .A(n13303), .B(n13304), .Z(n13292) );
  AND U12671 ( .A(n470), .B(n13305), .Z(n13304) );
  XOR U12672 ( .A(p_input[338]), .B(n13303), .Z(n13305) );
  XNOR U12673 ( .A(n13306), .B(n13307), .Z(n13303) );
  AND U12674 ( .A(n474), .B(n13308), .Z(n13307) );
  XOR U12675 ( .A(n13309), .B(n13310), .Z(n13301) );
  AND U12676 ( .A(n478), .B(n13311), .Z(n13310) );
  XOR U12677 ( .A(n13312), .B(n13313), .Z(n13298) );
  AND U12678 ( .A(n482), .B(n13311), .Z(n13313) );
  XNOR U12679 ( .A(n13314), .B(n13312), .Z(n13311) );
  IV U12680 ( .A(n13309), .Z(n13314) );
  XOR U12681 ( .A(n13315), .B(n13316), .Z(n13309) );
  AND U12682 ( .A(n485), .B(n13308), .Z(n13316) );
  XNOR U12683 ( .A(n13306), .B(n13315), .Z(n13308) );
  XNOR U12684 ( .A(n13317), .B(n13318), .Z(n13306) );
  AND U12685 ( .A(n489), .B(n13319), .Z(n13318) );
  XOR U12686 ( .A(p_input[354]), .B(n13317), .Z(n13319) );
  XNOR U12687 ( .A(n13320), .B(n13321), .Z(n13317) );
  AND U12688 ( .A(n493), .B(n13322), .Z(n13321) );
  XOR U12689 ( .A(n13323), .B(n13324), .Z(n13315) );
  AND U12690 ( .A(n497), .B(n13325), .Z(n13324) );
  XOR U12691 ( .A(n13326), .B(n13327), .Z(n13312) );
  AND U12692 ( .A(n501), .B(n13325), .Z(n13327) );
  XNOR U12693 ( .A(n13328), .B(n13326), .Z(n13325) );
  IV U12694 ( .A(n13323), .Z(n13328) );
  XOR U12695 ( .A(n13329), .B(n13330), .Z(n13323) );
  AND U12696 ( .A(n504), .B(n13322), .Z(n13330) );
  XNOR U12697 ( .A(n13320), .B(n13329), .Z(n13322) );
  XNOR U12698 ( .A(n13331), .B(n13332), .Z(n13320) );
  AND U12699 ( .A(n508), .B(n13333), .Z(n13332) );
  XOR U12700 ( .A(p_input[370]), .B(n13331), .Z(n13333) );
  XNOR U12701 ( .A(n13334), .B(n13335), .Z(n13331) );
  AND U12702 ( .A(n512), .B(n13336), .Z(n13335) );
  XOR U12703 ( .A(n13337), .B(n13338), .Z(n13329) );
  AND U12704 ( .A(n516), .B(n13339), .Z(n13338) );
  XOR U12705 ( .A(n13340), .B(n13341), .Z(n13326) );
  AND U12706 ( .A(n520), .B(n13339), .Z(n13341) );
  XNOR U12707 ( .A(n13342), .B(n13340), .Z(n13339) );
  IV U12708 ( .A(n13337), .Z(n13342) );
  XOR U12709 ( .A(n13343), .B(n13344), .Z(n13337) );
  AND U12710 ( .A(n523), .B(n13336), .Z(n13344) );
  XNOR U12711 ( .A(n13334), .B(n13343), .Z(n13336) );
  XNOR U12712 ( .A(n13345), .B(n13346), .Z(n13334) );
  AND U12713 ( .A(n527), .B(n13347), .Z(n13346) );
  XOR U12714 ( .A(p_input[386]), .B(n13345), .Z(n13347) );
  XNOR U12715 ( .A(n13348), .B(n13349), .Z(n13345) );
  AND U12716 ( .A(n531), .B(n13350), .Z(n13349) );
  XOR U12717 ( .A(n13351), .B(n13352), .Z(n13343) );
  AND U12718 ( .A(n535), .B(n13353), .Z(n13352) );
  XOR U12719 ( .A(n13354), .B(n13355), .Z(n13340) );
  AND U12720 ( .A(n539), .B(n13353), .Z(n13355) );
  XNOR U12721 ( .A(n13356), .B(n13354), .Z(n13353) );
  IV U12722 ( .A(n13351), .Z(n13356) );
  XOR U12723 ( .A(n13357), .B(n13358), .Z(n13351) );
  AND U12724 ( .A(n542), .B(n13350), .Z(n13358) );
  XNOR U12725 ( .A(n13348), .B(n13357), .Z(n13350) );
  XNOR U12726 ( .A(n13359), .B(n13360), .Z(n13348) );
  AND U12727 ( .A(n546), .B(n13361), .Z(n13360) );
  XOR U12728 ( .A(p_input[402]), .B(n13359), .Z(n13361) );
  XNOR U12729 ( .A(n13362), .B(n13363), .Z(n13359) );
  AND U12730 ( .A(n550), .B(n13364), .Z(n13363) );
  XOR U12731 ( .A(n13365), .B(n13366), .Z(n13357) );
  AND U12732 ( .A(n554), .B(n13367), .Z(n13366) );
  XOR U12733 ( .A(n13368), .B(n13369), .Z(n13354) );
  AND U12734 ( .A(n558), .B(n13367), .Z(n13369) );
  XNOR U12735 ( .A(n13370), .B(n13368), .Z(n13367) );
  IV U12736 ( .A(n13365), .Z(n13370) );
  XOR U12737 ( .A(n13371), .B(n13372), .Z(n13365) );
  AND U12738 ( .A(n561), .B(n13364), .Z(n13372) );
  XNOR U12739 ( .A(n13362), .B(n13371), .Z(n13364) );
  XNOR U12740 ( .A(n13373), .B(n13374), .Z(n13362) );
  AND U12741 ( .A(n565), .B(n13375), .Z(n13374) );
  XOR U12742 ( .A(p_input[418]), .B(n13373), .Z(n13375) );
  XNOR U12743 ( .A(n13376), .B(n13377), .Z(n13373) );
  AND U12744 ( .A(n569), .B(n13378), .Z(n13377) );
  XOR U12745 ( .A(n13379), .B(n13380), .Z(n13371) );
  AND U12746 ( .A(n573), .B(n13381), .Z(n13380) );
  XOR U12747 ( .A(n13382), .B(n13383), .Z(n13368) );
  AND U12748 ( .A(n577), .B(n13381), .Z(n13383) );
  XNOR U12749 ( .A(n13384), .B(n13382), .Z(n13381) );
  IV U12750 ( .A(n13379), .Z(n13384) );
  XOR U12751 ( .A(n13385), .B(n13386), .Z(n13379) );
  AND U12752 ( .A(n580), .B(n13378), .Z(n13386) );
  XNOR U12753 ( .A(n13376), .B(n13385), .Z(n13378) );
  XNOR U12754 ( .A(n13387), .B(n13388), .Z(n13376) );
  AND U12755 ( .A(n584), .B(n13389), .Z(n13388) );
  XOR U12756 ( .A(p_input[434]), .B(n13387), .Z(n13389) );
  XNOR U12757 ( .A(n13390), .B(n13391), .Z(n13387) );
  AND U12758 ( .A(n588), .B(n13392), .Z(n13391) );
  XOR U12759 ( .A(n13393), .B(n13394), .Z(n13385) );
  AND U12760 ( .A(n592), .B(n13395), .Z(n13394) );
  XOR U12761 ( .A(n13396), .B(n13397), .Z(n13382) );
  AND U12762 ( .A(n596), .B(n13395), .Z(n13397) );
  XNOR U12763 ( .A(n13398), .B(n13396), .Z(n13395) );
  IV U12764 ( .A(n13393), .Z(n13398) );
  XOR U12765 ( .A(n13399), .B(n13400), .Z(n13393) );
  AND U12766 ( .A(n599), .B(n13392), .Z(n13400) );
  XNOR U12767 ( .A(n13390), .B(n13399), .Z(n13392) );
  XNOR U12768 ( .A(n13401), .B(n13402), .Z(n13390) );
  AND U12769 ( .A(n603), .B(n13403), .Z(n13402) );
  XOR U12770 ( .A(p_input[450]), .B(n13401), .Z(n13403) );
  XNOR U12771 ( .A(n13404), .B(n13405), .Z(n13401) );
  AND U12772 ( .A(n607), .B(n13406), .Z(n13405) );
  XOR U12773 ( .A(n13407), .B(n13408), .Z(n13399) );
  AND U12774 ( .A(n611), .B(n13409), .Z(n13408) );
  XOR U12775 ( .A(n13410), .B(n13411), .Z(n13396) );
  AND U12776 ( .A(n615), .B(n13409), .Z(n13411) );
  XNOR U12777 ( .A(n13412), .B(n13410), .Z(n13409) );
  IV U12778 ( .A(n13407), .Z(n13412) );
  XOR U12779 ( .A(n13413), .B(n13414), .Z(n13407) );
  AND U12780 ( .A(n618), .B(n13406), .Z(n13414) );
  XNOR U12781 ( .A(n13404), .B(n13413), .Z(n13406) );
  XNOR U12782 ( .A(n13415), .B(n13416), .Z(n13404) );
  AND U12783 ( .A(n622), .B(n13417), .Z(n13416) );
  XOR U12784 ( .A(p_input[466]), .B(n13415), .Z(n13417) );
  XNOR U12785 ( .A(n13418), .B(n13419), .Z(n13415) );
  AND U12786 ( .A(n626), .B(n13420), .Z(n13419) );
  XOR U12787 ( .A(n13421), .B(n13422), .Z(n13413) );
  AND U12788 ( .A(n630), .B(n13423), .Z(n13422) );
  XOR U12789 ( .A(n13424), .B(n13425), .Z(n13410) );
  AND U12790 ( .A(n634), .B(n13423), .Z(n13425) );
  XNOR U12791 ( .A(n13426), .B(n13424), .Z(n13423) );
  IV U12792 ( .A(n13421), .Z(n13426) );
  XOR U12793 ( .A(n13427), .B(n13428), .Z(n13421) );
  AND U12794 ( .A(n637), .B(n13420), .Z(n13428) );
  XNOR U12795 ( .A(n13418), .B(n13427), .Z(n13420) );
  XNOR U12796 ( .A(n13429), .B(n13430), .Z(n13418) );
  AND U12797 ( .A(n641), .B(n13431), .Z(n13430) );
  XOR U12798 ( .A(p_input[482]), .B(n13429), .Z(n13431) );
  XNOR U12799 ( .A(n13432), .B(n13433), .Z(n13429) );
  AND U12800 ( .A(n645), .B(n13434), .Z(n13433) );
  XOR U12801 ( .A(n13435), .B(n13436), .Z(n13427) );
  AND U12802 ( .A(n649), .B(n13437), .Z(n13436) );
  XOR U12803 ( .A(n13438), .B(n13439), .Z(n13424) );
  AND U12804 ( .A(n653), .B(n13437), .Z(n13439) );
  XNOR U12805 ( .A(n13440), .B(n13438), .Z(n13437) );
  IV U12806 ( .A(n13435), .Z(n13440) );
  XOR U12807 ( .A(n13441), .B(n13442), .Z(n13435) );
  AND U12808 ( .A(n656), .B(n13434), .Z(n13442) );
  XNOR U12809 ( .A(n13432), .B(n13441), .Z(n13434) );
  XNOR U12810 ( .A(n13443), .B(n13444), .Z(n13432) );
  AND U12811 ( .A(n660), .B(n13445), .Z(n13444) );
  XOR U12812 ( .A(p_input[498]), .B(n13443), .Z(n13445) );
  XNOR U12813 ( .A(n13446), .B(n13447), .Z(n13443) );
  AND U12814 ( .A(n664), .B(n13448), .Z(n13447) );
  XOR U12815 ( .A(n13449), .B(n13450), .Z(n13441) );
  AND U12816 ( .A(n668), .B(n13451), .Z(n13450) );
  XOR U12817 ( .A(n13452), .B(n13453), .Z(n13438) );
  AND U12818 ( .A(n672), .B(n13451), .Z(n13453) );
  XNOR U12819 ( .A(n13454), .B(n13452), .Z(n13451) );
  IV U12820 ( .A(n13449), .Z(n13454) );
  XOR U12821 ( .A(n13455), .B(n13456), .Z(n13449) );
  AND U12822 ( .A(n675), .B(n13448), .Z(n13456) );
  XNOR U12823 ( .A(n13446), .B(n13455), .Z(n13448) );
  XNOR U12824 ( .A(n13457), .B(n13458), .Z(n13446) );
  AND U12825 ( .A(n679), .B(n13459), .Z(n13458) );
  XOR U12826 ( .A(p_input[514]), .B(n13457), .Z(n13459) );
  XNOR U12827 ( .A(n13460), .B(n13461), .Z(n13457) );
  AND U12828 ( .A(n683), .B(n13462), .Z(n13461) );
  XOR U12829 ( .A(n13463), .B(n13464), .Z(n13455) );
  AND U12830 ( .A(n687), .B(n13465), .Z(n13464) );
  XOR U12831 ( .A(n13466), .B(n13467), .Z(n13452) );
  AND U12832 ( .A(n691), .B(n13465), .Z(n13467) );
  XNOR U12833 ( .A(n13468), .B(n13466), .Z(n13465) );
  IV U12834 ( .A(n13463), .Z(n13468) );
  XOR U12835 ( .A(n13469), .B(n13470), .Z(n13463) );
  AND U12836 ( .A(n694), .B(n13462), .Z(n13470) );
  XNOR U12837 ( .A(n13460), .B(n13469), .Z(n13462) );
  XNOR U12838 ( .A(n13471), .B(n13472), .Z(n13460) );
  AND U12839 ( .A(n698), .B(n13473), .Z(n13472) );
  XOR U12840 ( .A(p_input[530]), .B(n13471), .Z(n13473) );
  XNOR U12841 ( .A(n13474), .B(n13475), .Z(n13471) );
  AND U12842 ( .A(n702), .B(n13476), .Z(n13475) );
  XOR U12843 ( .A(n13477), .B(n13478), .Z(n13469) );
  AND U12844 ( .A(n706), .B(n13479), .Z(n13478) );
  XOR U12845 ( .A(n13480), .B(n13481), .Z(n13466) );
  AND U12846 ( .A(n710), .B(n13479), .Z(n13481) );
  XNOR U12847 ( .A(n13482), .B(n13480), .Z(n13479) );
  IV U12848 ( .A(n13477), .Z(n13482) );
  XOR U12849 ( .A(n13483), .B(n13484), .Z(n13477) );
  AND U12850 ( .A(n713), .B(n13476), .Z(n13484) );
  XNOR U12851 ( .A(n13474), .B(n13483), .Z(n13476) );
  XNOR U12852 ( .A(n13485), .B(n13486), .Z(n13474) );
  AND U12853 ( .A(n717), .B(n13487), .Z(n13486) );
  XOR U12854 ( .A(p_input[546]), .B(n13485), .Z(n13487) );
  XNOR U12855 ( .A(n13488), .B(n13489), .Z(n13485) );
  AND U12856 ( .A(n721), .B(n13490), .Z(n13489) );
  XOR U12857 ( .A(n13491), .B(n13492), .Z(n13483) );
  AND U12858 ( .A(n725), .B(n13493), .Z(n13492) );
  XOR U12859 ( .A(n13494), .B(n13495), .Z(n13480) );
  AND U12860 ( .A(n729), .B(n13493), .Z(n13495) );
  XNOR U12861 ( .A(n13496), .B(n13494), .Z(n13493) );
  IV U12862 ( .A(n13491), .Z(n13496) );
  XOR U12863 ( .A(n13497), .B(n13498), .Z(n13491) );
  AND U12864 ( .A(n732), .B(n13490), .Z(n13498) );
  XNOR U12865 ( .A(n13488), .B(n13497), .Z(n13490) );
  XNOR U12866 ( .A(n13499), .B(n13500), .Z(n13488) );
  AND U12867 ( .A(n736), .B(n13501), .Z(n13500) );
  XOR U12868 ( .A(p_input[562]), .B(n13499), .Z(n13501) );
  XNOR U12869 ( .A(n13502), .B(n13503), .Z(n13499) );
  AND U12870 ( .A(n740), .B(n13504), .Z(n13503) );
  XOR U12871 ( .A(n13505), .B(n13506), .Z(n13497) );
  AND U12872 ( .A(n744), .B(n13507), .Z(n13506) );
  XOR U12873 ( .A(n13508), .B(n13509), .Z(n13494) );
  AND U12874 ( .A(n748), .B(n13507), .Z(n13509) );
  XNOR U12875 ( .A(n13510), .B(n13508), .Z(n13507) );
  IV U12876 ( .A(n13505), .Z(n13510) );
  XOR U12877 ( .A(n13511), .B(n13512), .Z(n13505) );
  AND U12878 ( .A(n751), .B(n13504), .Z(n13512) );
  XNOR U12879 ( .A(n13502), .B(n13511), .Z(n13504) );
  XNOR U12880 ( .A(n13513), .B(n13514), .Z(n13502) );
  AND U12881 ( .A(n755), .B(n13515), .Z(n13514) );
  XOR U12882 ( .A(p_input[578]), .B(n13513), .Z(n13515) );
  XNOR U12883 ( .A(n13516), .B(n13517), .Z(n13513) );
  AND U12884 ( .A(n759), .B(n13518), .Z(n13517) );
  XOR U12885 ( .A(n13519), .B(n13520), .Z(n13511) );
  AND U12886 ( .A(n763), .B(n13521), .Z(n13520) );
  XOR U12887 ( .A(n13522), .B(n13523), .Z(n13508) );
  AND U12888 ( .A(n767), .B(n13521), .Z(n13523) );
  XNOR U12889 ( .A(n13524), .B(n13522), .Z(n13521) );
  IV U12890 ( .A(n13519), .Z(n13524) );
  XOR U12891 ( .A(n13525), .B(n13526), .Z(n13519) );
  AND U12892 ( .A(n770), .B(n13518), .Z(n13526) );
  XNOR U12893 ( .A(n13516), .B(n13525), .Z(n13518) );
  XNOR U12894 ( .A(n13527), .B(n13528), .Z(n13516) );
  AND U12895 ( .A(n774), .B(n13529), .Z(n13528) );
  XOR U12896 ( .A(p_input[594]), .B(n13527), .Z(n13529) );
  XNOR U12897 ( .A(n13530), .B(n13531), .Z(n13527) );
  AND U12898 ( .A(n778), .B(n13532), .Z(n13531) );
  XOR U12899 ( .A(n13533), .B(n13534), .Z(n13525) );
  AND U12900 ( .A(n782), .B(n13535), .Z(n13534) );
  XOR U12901 ( .A(n13536), .B(n13537), .Z(n13522) );
  AND U12902 ( .A(n786), .B(n13535), .Z(n13537) );
  XNOR U12903 ( .A(n13538), .B(n13536), .Z(n13535) );
  IV U12904 ( .A(n13533), .Z(n13538) );
  XOR U12905 ( .A(n13539), .B(n13540), .Z(n13533) );
  AND U12906 ( .A(n789), .B(n13532), .Z(n13540) );
  XNOR U12907 ( .A(n13530), .B(n13539), .Z(n13532) );
  XNOR U12908 ( .A(n13541), .B(n13542), .Z(n13530) );
  AND U12909 ( .A(n793), .B(n13543), .Z(n13542) );
  XOR U12910 ( .A(p_input[610]), .B(n13541), .Z(n13543) );
  XNOR U12911 ( .A(n13544), .B(n13545), .Z(n13541) );
  AND U12912 ( .A(n797), .B(n13546), .Z(n13545) );
  XOR U12913 ( .A(n13547), .B(n13548), .Z(n13539) );
  AND U12914 ( .A(n801), .B(n13549), .Z(n13548) );
  XOR U12915 ( .A(n13550), .B(n13551), .Z(n13536) );
  AND U12916 ( .A(n805), .B(n13549), .Z(n13551) );
  XNOR U12917 ( .A(n13552), .B(n13550), .Z(n13549) );
  IV U12918 ( .A(n13547), .Z(n13552) );
  XOR U12919 ( .A(n13553), .B(n13554), .Z(n13547) );
  AND U12920 ( .A(n808), .B(n13546), .Z(n13554) );
  XNOR U12921 ( .A(n13544), .B(n13553), .Z(n13546) );
  XNOR U12922 ( .A(n13555), .B(n13556), .Z(n13544) );
  AND U12923 ( .A(n812), .B(n13557), .Z(n13556) );
  XOR U12924 ( .A(p_input[626]), .B(n13555), .Z(n13557) );
  XNOR U12925 ( .A(n13558), .B(n13559), .Z(n13555) );
  AND U12926 ( .A(n816), .B(n13560), .Z(n13559) );
  XOR U12927 ( .A(n13561), .B(n13562), .Z(n13553) );
  AND U12928 ( .A(n820), .B(n13563), .Z(n13562) );
  XOR U12929 ( .A(n13564), .B(n13565), .Z(n13550) );
  AND U12930 ( .A(n824), .B(n13563), .Z(n13565) );
  XNOR U12931 ( .A(n13566), .B(n13564), .Z(n13563) );
  IV U12932 ( .A(n13561), .Z(n13566) );
  XOR U12933 ( .A(n13567), .B(n13568), .Z(n13561) );
  AND U12934 ( .A(n827), .B(n13560), .Z(n13568) );
  XNOR U12935 ( .A(n13558), .B(n13567), .Z(n13560) );
  XNOR U12936 ( .A(n13569), .B(n13570), .Z(n13558) );
  AND U12937 ( .A(n831), .B(n13571), .Z(n13570) );
  XOR U12938 ( .A(p_input[642]), .B(n13569), .Z(n13571) );
  XNOR U12939 ( .A(n13572), .B(n13573), .Z(n13569) );
  AND U12940 ( .A(n835), .B(n13574), .Z(n13573) );
  XOR U12941 ( .A(n13575), .B(n13576), .Z(n13567) );
  AND U12942 ( .A(n839), .B(n13577), .Z(n13576) );
  XOR U12943 ( .A(n13578), .B(n13579), .Z(n13564) );
  AND U12944 ( .A(n843), .B(n13577), .Z(n13579) );
  XNOR U12945 ( .A(n13580), .B(n13578), .Z(n13577) );
  IV U12946 ( .A(n13575), .Z(n13580) );
  XOR U12947 ( .A(n13581), .B(n13582), .Z(n13575) );
  AND U12948 ( .A(n846), .B(n13574), .Z(n13582) );
  XNOR U12949 ( .A(n13572), .B(n13581), .Z(n13574) );
  XNOR U12950 ( .A(n13583), .B(n13584), .Z(n13572) );
  AND U12951 ( .A(n850), .B(n13585), .Z(n13584) );
  XOR U12952 ( .A(p_input[658]), .B(n13583), .Z(n13585) );
  XNOR U12953 ( .A(n13586), .B(n13587), .Z(n13583) );
  AND U12954 ( .A(n854), .B(n13588), .Z(n13587) );
  XOR U12955 ( .A(n13589), .B(n13590), .Z(n13581) );
  AND U12956 ( .A(n858), .B(n13591), .Z(n13590) );
  XOR U12957 ( .A(n13592), .B(n13593), .Z(n13578) );
  AND U12958 ( .A(n862), .B(n13591), .Z(n13593) );
  XNOR U12959 ( .A(n13594), .B(n13592), .Z(n13591) );
  IV U12960 ( .A(n13589), .Z(n13594) );
  XOR U12961 ( .A(n13595), .B(n13596), .Z(n13589) );
  AND U12962 ( .A(n865), .B(n13588), .Z(n13596) );
  XNOR U12963 ( .A(n13586), .B(n13595), .Z(n13588) );
  XNOR U12964 ( .A(n13597), .B(n13598), .Z(n13586) );
  AND U12965 ( .A(n869), .B(n13599), .Z(n13598) );
  XOR U12966 ( .A(p_input[674]), .B(n13597), .Z(n13599) );
  XNOR U12967 ( .A(n13600), .B(n13601), .Z(n13597) );
  AND U12968 ( .A(n873), .B(n13602), .Z(n13601) );
  XOR U12969 ( .A(n13603), .B(n13604), .Z(n13595) );
  AND U12970 ( .A(n877), .B(n13605), .Z(n13604) );
  XOR U12971 ( .A(n13606), .B(n13607), .Z(n13592) );
  AND U12972 ( .A(n881), .B(n13605), .Z(n13607) );
  XNOR U12973 ( .A(n13608), .B(n13606), .Z(n13605) );
  IV U12974 ( .A(n13603), .Z(n13608) );
  XOR U12975 ( .A(n13609), .B(n13610), .Z(n13603) );
  AND U12976 ( .A(n884), .B(n13602), .Z(n13610) );
  XNOR U12977 ( .A(n13600), .B(n13609), .Z(n13602) );
  XNOR U12978 ( .A(n13611), .B(n13612), .Z(n13600) );
  AND U12979 ( .A(n888), .B(n13613), .Z(n13612) );
  XOR U12980 ( .A(p_input[690]), .B(n13611), .Z(n13613) );
  XNOR U12981 ( .A(n13614), .B(n13615), .Z(n13611) );
  AND U12982 ( .A(n892), .B(n13616), .Z(n13615) );
  XOR U12983 ( .A(n13617), .B(n13618), .Z(n13609) );
  AND U12984 ( .A(n896), .B(n13619), .Z(n13618) );
  XOR U12985 ( .A(n13620), .B(n13621), .Z(n13606) );
  AND U12986 ( .A(n900), .B(n13619), .Z(n13621) );
  XNOR U12987 ( .A(n13622), .B(n13620), .Z(n13619) );
  IV U12988 ( .A(n13617), .Z(n13622) );
  XOR U12989 ( .A(n13623), .B(n13624), .Z(n13617) );
  AND U12990 ( .A(n903), .B(n13616), .Z(n13624) );
  XNOR U12991 ( .A(n13614), .B(n13623), .Z(n13616) );
  XNOR U12992 ( .A(n13625), .B(n13626), .Z(n13614) );
  AND U12993 ( .A(n907), .B(n13627), .Z(n13626) );
  XOR U12994 ( .A(p_input[706]), .B(n13625), .Z(n13627) );
  XNOR U12995 ( .A(n13628), .B(n13629), .Z(n13625) );
  AND U12996 ( .A(n911), .B(n13630), .Z(n13629) );
  XOR U12997 ( .A(n13631), .B(n13632), .Z(n13623) );
  AND U12998 ( .A(n915), .B(n13633), .Z(n13632) );
  XOR U12999 ( .A(n13634), .B(n13635), .Z(n13620) );
  AND U13000 ( .A(n919), .B(n13633), .Z(n13635) );
  XNOR U13001 ( .A(n13636), .B(n13634), .Z(n13633) );
  IV U13002 ( .A(n13631), .Z(n13636) );
  XOR U13003 ( .A(n13637), .B(n13638), .Z(n13631) );
  AND U13004 ( .A(n922), .B(n13630), .Z(n13638) );
  XNOR U13005 ( .A(n13628), .B(n13637), .Z(n13630) );
  XNOR U13006 ( .A(n13639), .B(n13640), .Z(n13628) );
  AND U13007 ( .A(n926), .B(n13641), .Z(n13640) );
  XOR U13008 ( .A(p_input[722]), .B(n13639), .Z(n13641) );
  XNOR U13009 ( .A(n13642), .B(n13643), .Z(n13639) );
  AND U13010 ( .A(n930), .B(n13644), .Z(n13643) );
  XOR U13011 ( .A(n13645), .B(n13646), .Z(n13637) );
  AND U13012 ( .A(n934), .B(n13647), .Z(n13646) );
  XOR U13013 ( .A(n13648), .B(n13649), .Z(n13634) );
  AND U13014 ( .A(n938), .B(n13647), .Z(n13649) );
  XNOR U13015 ( .A(n13650), .B(n13648), .Z(n13647) );
  IV U13016 ( .A(n13645), .Z(n13650) );
  XOR U13017 ( .A(n13651), .B(n13652), .Z(n13645) );
  AND U13018 ( .A(n941), .B(n13644), .Z(n13652) );
  XNOR U13019 ( .A(n13642), .B(n13651), .Z(n13644) );
  XNOR U13020 ( .A(n13653), .B(n13654), .Z(n13642) );
  AND U13021 ( .A(n945), .B(n13655), .Z(n13654) );
  XOR U13022 ( .A(p_input[738]), .B(n13653), .Z(n13655) );
  XNOR U13023 ( .A(n13656), .B(n13657), .Z(n13653) );
  AND U13024 ( .A(n949), .B(n13658), .Z(n13657) );
  XOR U13025 ( .A(n13659), .B(n13660), .Z(n13651) );
  AND U13026 ( .A(n953), .B(n13661), .Z(n13660) );
  XOR U13027 ( .A(n13662), .B(n13663), .Z(n13648) );
  AND U13028 ( .A(n957), .B(n13661), .Z(n13663) );
  XNOR U13029 ( .A(n13664), .B(n13662), .Z(n13661) );
  IV U13030 ( .A(n13659), .Z(n13664) );
  XOR U13031 ( .A(n13665), .B(n13666), .Z(n13659) );
  AND U13032 ( .A(n960), .B(n13658), .Z(n13666) );
  XNOR U13033 ( .A(n13656), .B(n13665), .Z(n13658) );
  XNOR U13034 ( .A(n13667), .B(n13668), .Z(n13656) );
  AND U13035 ( .A(n964), .B(n13669), .Z(n13668) );
  XOR U13036 ( .A(p_input[754]), .B(n13667), .Z(n13669) );
  XNOR U13037 ( .A(n13670), .B(n13671), .Z(n13667) );
  AND U13038 ( .A(n968), .B(n13672), .Z(n13671) );
  XOR U13039 ( .A(n13673), .B(n13674), .Z(n13665) );
  AND U13040 ( .A(n972), .B(n13675), .Z(n13674) );
  XOR U13041 ( .A(n13676), .B(n13677), .Z(n13662) );
  AND U13042 ( .A(n976), .B(n13675), .Z(n13677) );
  XNOR U13043 ( .A(n13678), .B(n13676), .Z(n13675) );
  IV U13044 ( .A(n13673), .Z(n13678) );
  XOR U13045 ( .A(n13679), .B(n13680), .Z(n13673) );
  AND U13046 ( .A(n979), .B(n13672), .Z(n13680) );
  XNOR U13047 ( .A(n13670), .B(n13679), .Z(n13672) );
  XNOR U13048 ( .A(n13681), .B(n13682), .Z(n13670) );
  AND U13049 ( .A(n983), .B(n13683), .Z(n13682) );
  XOR U13050 ( .A(p_input[770]), .B(n13681), .Z(n13683) );
  XNOR U13051 ( .A(n13684), .B(n13685), .Z(n13681) );
  AND U13052 ( .A(n987), .B(n13686), .Z(n13685) );
  XOR U13053 ( .A(n13687), .B(n13688), .Z(n13679) );
  AND U13054 ( .A(n991), .B(n13689), .Z(n13688) );
  XOR U13055 ( .A(n13690), .B(n13691), .Z(n13676) );
  AND U13056 ( .A(n995), .B(n13689), .Z(n13691) );
  XNOR U13057 ( .A(n13692), .B(n13690), .Z(n13689) );
  IV U13058 ( .A(n13687), .Z(n13692) );
  XOR U13059 ( .A(n13693), .B(n13694), .Z(n13687) );
  AND U13060 ( .A(n998), .B(n13686), .Z(n13694) );
  XNOR U13061 ( .A(n13684), .B(n13693), .Z(n13686) );
  XNOR U13062 ( .A(n13695), .B(n13696), .Z(n13684) );
  AND U13063 ( .A(n1002), .B(n13697), .Z(n13696) );
  XOR U13064 ( .A(p_input[786]), .B(n13695), .Z(n13697) );
  XNOR U13065 ( .A(n13698), .B(n13699), .Z(n13695) );
  AND U13066 ( .A(n1006), .B(n13700), .Z(n13699) );
  XOR U13067 ( .A(n13701), .B(n13702), .Z(n13693) );
  AND U13068 ( .A(n1010), .B(n13703), .Z(n13702) );
  XOR U13069 ( .A(n13704), .B(n13705), .Z(n13690) );
  AND U13070 ( .A(n1014), .B(n13703), .Z(n13705) );
  XNOR U13071 ( .A(n13706), .B(n13704), .Z(n13703) );
  IV U13072 ( .A(n13701), .Z(n13706) );
  XOR U13073 ( .A(n13707), .B(n13708), .Z(n13701) );
  AND U13074 ( .A(n1017), .B(n13700), .Z(n13708) );
  XNOR U13075 ( .A(n13698), .B(n13707), .Z(n13700) );
  XNOR U13076 ( .A(n13709), .B(n13710), .Z(n13698) );
  AND U13077 ( .A(n1021), .B(n13711), .Z(n13710) );
  XOR U13078 ( .A(p_input[802]), .B(n13709), .Z(n13711) );
  XNOR U13079 ( .A(n13712), .B(n13713), .Z(n13709) );
  AND U13080 ( .A(n1025), .B(n13714), .Z(n13713) );
  XOR U13081 ( .A(n13715), .B(n13716), .Z(n13707) );
  AND U13082 ( .A(n1029), .B(n13717), .Z(n13716) );
  XOR U13083 ( .A(n13718), .B(n13719), .Z(n13704) );
  AND U13084 ( .A(n1033), .B(n13717), .Z(n13719) );
  XNOR U13085 ( .A(n13720), .B(n13718), .Z(n13717) );
  IV U13086 ( .A(n13715), .Z(n13720) );
  XOR U13087 ( .A(n13721), .B(n13722), .Z(n13715) );
  AND U13088 ( .A(n1036), .B(n13714), .Z(n13722) );
  XNOR U13089 ( .A(n13712), .B(n13721), .Z(n13714) );
  XNOR U13090 ( .A(n13723), .B(n13724), .Z(n13712) );
  AND U13091 ( .A(n1040), .B(n13725), .Z(n13724) );
  XOR U13092 ( .A(p_input[818]), .B(n13723), .Z(n13725) );
  XNOR U13093 ( .A(n13726), .B(n13727), .Z(n13723) );
  AND U13094 ( .A(n1044), .B(n13728), .Z(n13727) );
  XOR U13095 ( .A(n13729), .B(n13730), .Z(n13721) );
  AND U13096 ( .A(n1048), .B(n13731), .Z(n13730) );
  XOR U13097 ( .A(n13732), .B(n13733), .Z(n13718) );
  AND U13098 ( .A(n1052), .B(n13731), .Z(n13733) );
  XNOR U13099 ( .A(n13734), .B(n13732), .Z(n13731) );
  IV U13100 ( .A(n13729), .Z(n13734) );
  XOR U13101 ( .A(n13735), .B(n13736), .Z(n13729) );
  AND U13102 ( .A(n1055), .B(n13728), .Z(n13736) );
  XNOR U13103 ( .A(n13726), .B(n13735), .Z(n13728) );
  XNOR U13104 ( .A(n13737), .B(n13738), .Z(n13726) );
  AND U13105 ( .A(n1059), .B(n13739), .Z(n13738) );
  XOR U13106 ( .A(p_input[834]), .B(n13737), .Z(n13739) );
  XNOR U13107 ( .A(n13740), .B(n13741), .Z(n13737) );
  AND U13108 ( .A(n1063), .B(n13742), .Z(n13741) );
  XOR U13109 ( .A(n13743), .B(n13744), .Z(n13735) );
  AND U13110 ( .A(n1067), .B(n13745), .Z(n13744) );
  XOR U13111 ( .A(n13746), .B(n13747), .Z(n13732) );
  AND U13112 ( .A(n1071), .B(n13745), .Z(n13747) );
  XNOR U13113 ( .A(n13748), .B(n13746), .Z(n13745) );
  IV U13114 ( .A(n13743), .Z(n13748) );
  XOR U13115 ( .A(n13749), .B(n13750), .Z(n13743) );
  AND U13116 ( .A(n1074), .B(n13742), .Z(n13750) );
  XNOR U13117 ( .A(n13740), .B(n13749), .Z(n13742) );
  XNOR U13118 ( .A(n13751), .B(n13752), .Z(n13740) );
  AND U13119 ( .A(n1078), .B(n13753), .Z(n13752) );
  XOR U13120 ( .A(p_input[850]), .B(n13751), .Z(n13753) );
  XNOR U13121 ( .A(n13754), .B(n13755), .Z(n13751) );
  AND U13122 ( .A(n1082), .B(n13756), .Z(n13755) );
  XOR U13123 ( .A(n13757), .B(n13758), .Z(n13749) );
  AND U13124 ( .A(n1086), .B(n13759), .Z(n13758) );
  XOR U13125 ( .A(n13760), .B(n13761), .Z(n13746) );
  AND U13126 ( .A(n1090), .B(n13759), .Z(n13761) );
  XNOR U13127 ( .A(n13762), .B(n13760), .Z(n13759) );
  IV U13128 ( .A(n13757), .Z(n13762) );
  XOR U13129 ( .A(n13763), .B(n13764), .Z(n13757) );
  AND U13130 ( .A(n1093), .B(n13756), .Z(n13764) );
  XNOR U13131 ( .A(n13754), .B(n13763), .Z(n13756) );
  XNOR U13132 ( .A(n13765), .B(n13766), .Z(n13754) );
  AND U13133 ( .A(n1097), .B(n13767), .Z(n13766) );
  XOR U13134 ( .A(p_input[866]), .B(n13765), .Z(n13767) );
  XNOR U13135 ( .A(n13768), .B(n13769), .Z(n13765) );
  AND U13136 ( .A(n1101), .B(n13770), .Z(n13769) );
  XOR U13137 ( .A(n13771), .B(n13772), .Z(n13763) );
  AND U13138 ( .A(n1105), .B(n13773), .Z(n13772) );
  XOR U13139 ( .A(n13774), .B(n13775), .Z(n13760) );
  AND U13140 ( .A(n1109), .B(n13773), .Z(n13775) );
  XNOR U13141 ( .A(n13776), .B(n13774), .Z(n13773) );
  IV U13142 ( .A(n13771), .Z(n13776) );
  XOR U13143 ( .A(n13777), .B(n13778), .Z(n13771) );
  AND U13144 ( .A(n1112), .B(n13770), .Z(n13778) );
  XNOR U13145 ( .A(n13768), .B(n13777), .Z(n13770) );
  XNOR U13146 ( .A(n13779), .B(n13780), .Z(n13768) );
  AND U13147 ( .A(n1116), .B(n13781), .Z(n13780) );
  XOR U13148 ( .A(p_input[882]), .B(n13779), .Z(n13781) );
  XNOR U13149 ( .A(n13782), .B(n13783), .Z(n13779) );
  AND U13150 ( .A(n1120), .B(n13784), .Z(n13783) );
  XOR U13151 ( .A(n13785), .B(n13786), .Z(n13777) );
  AND U13152 ( .A(n1124), .B(n13787), .Z(n13786) );
  XOR U13153 ( .A(n13788), .B(n13789), .Z(n13774) );
  AND U13154 ( .A(n1128), .B(n13787), .Z(n13789) );
  XNOR U13155 ( .A(n13790), .B(n13788), .Z(n13787) );
  IV U13156 ( .A(n13785), .Z(n13790) );
  XOR U13157 ( .A(n13791), .B(n13792), .Z(n13785) );
  AND U13158 ( .A(n1131), .B(n13784), .Z(n13792) );
  XNOR U13159 ( .A(n13782), .B(n13791), .Z(n13784) );
  XNOR U13160 ( .A(n13793), .B(n13794), .Z(n13782) );
  AND U13161 ( .A(n1135), .B(n13795), .Z(n13794) );
  XOR U13162 ( .A(p_input[898]), .B(n13793), .Z(n13795) );
  XNOR U13163 ( .A(n13796), .B(n13797), .Z(n13793) );
  AND U13164 ( .A(n1139), .B(n13798), .Z(n13797) );
  XOR U13165 ( .A(n13799), .B(n13800), .Z(n13791) );
  AND U13166 ( .A(n1143), .B(n13801), .Z(n13800) );
  XOR U13167 ( .A(n13802), .B(n13803), .Z(n13788) );
  AND U13168 ( .A(n1147), .B(n13801), .Z(n13803) );
  XNOR U13169 ( .A(n13804), .B(n13802), .Z(n13801) );
  IV U13170 ( .A(n13799), .Z(n13804) );
  XOR U13171 ( .A(n13805), .B(n13806), .Z(n13799) );
  AND U13172 ( .A(n1150), .B(n13798), .Z(n13806) );
  XNOR U13173 ( .A(n13796), .B(n13805), .Z(n13798) );
  XNOR U13174 ( .A(n13807), .B(n13808), .Z(n13796) );
  AND U13175 ( .A(n1154), .B(n13809), .Z(n13808) );
  XOR U13176 ( .A(p_input[914]), .B(n13807), .Z(n13809) );
  XNOR U13177 ( .A(n13810), .B(n13811), .Z(n13807) );
  AND U13178 ( .A(n1158), .B(n13812), .Z(n13811) );
  XOR U13179 ( .A(n13813), .B(n13814), .Z(n13805) );
  AND U13180 ( .A(n1162), .B(n13815), .Z(n13814) );
  XOR U13181 ( .A(n13816), .B(n13817), .Z(n13802) );
  AND U13182 ( .A(n1166), .B(n13815), .Z(n13817) );
  XNOR U13183 ( .A(n13818), .B(n13816), .Z(n13815) );
  IV U13184 ( .A(n13813), .Z(n13818) );
  XOR U13185 ( .A(n13819), .B(n13820), .Z(n13813) );
  AND U13186 ( .A(n1169), .B(n13812), .Z(n13820) );
  XNOR U13187 ( .A(n13810), .B(n13819), .Z(n13812) );
  XNOR U13188 ( .A(n13821), .B(n13822), .Z(n13810) );
  AND U13189 ( .A(n1173), .B(n13823), .Z(n13822) );
  XOR U13190 ( .A(p_input[930]), .B(n13821), .Z(n13823) );
  XNOR U13191 ( .A(n13824), .B(n13825), .Z(n13821) );
  AND U13192 ( .A(n1177), .B(n13826), .Z(n13825) );
  XOR U13193 ( .A(n13827), .B(n13828), .Z(n13819) );
  AND U13194 ( .A(n1181), .B(n13829), .Z(n13828) );
  XOR U13195 ( .A(n13830), .B(n13831), .Z(n13816) );
  AND U13196 ( .A(n1185), .B(n13829), .Z(n13831) );
  XNOR U13197 ( .A(n13832), .B(n13830), .Z(n13829) );
  IV U13198 ( .A(n13827), .Z(n13832) );
  XOR U13199 ( .A(n13833), .B(n13834), .Z(n13827) );
  AND U13200 ( .A(n1188), .B(n13826), .Z(n13834) );
  XNOR U13201 ( .A(n13824), .B(n13833), .Z(n13826) );
  XNOR U13202 ( .A(n13835), .B(n13836), .Z(n13824) );
  AND U13203 ( .A(n1192), .B(n13837), .Z(n13836) );
  XOR U13204 ( .A(p_input[946]), .B(n13835), .Z(n13837) );
  XNOR U13205 ( .A(n13838), .B(n13839), .Z(n13835) );
  AND U13206 ( .A(n1196), .B(n13840), .Z(n13839) );
  XOR U13207 ( .A(n13841), .B(n13842), .Z(n13833) );
  AND U13208 ( .A(n1200), .B(n13843), .Z(n13842) );
  XOR U13209 ( .A(n13844), .B(n13845), .Z(n13830) );
  AND U13210 ( .A(n1204), .B(n13843), .Z(n13845) );
  XNOR U13211 ( .A(n13846), .B(n13844), .Z(n13843) );
  IV U13212 ( .A(n13841), .Z(n13846) );
  XOR U13213 ( .A(n13847), .B(n13848), .Z(n13841) );
  AND U13214 ( .A(n1207), .B(n13840), .Z(n13848) );
  XNOR U13215 ( .A(n13838), .B(n13847), .Z(n13840) );
  XNOR U13216 ( .A(n13849), .B(n13850), .Z(n13838) );
  AND U13217 ( .A(n1211), .B(n13851), .Z(n13850) );
  XOR U13218 ( .A(p_input[962]), .B(n13849), .Z(n13851) );
  XNOR U13219 ( .A(n13852), .B(n13853), .Z(n13849) );
  AND U13220 ( .A(n1215), .B(n13854), .Z(n13853) );
  XOR U13221 ( .A(n13855), .B(n13856), .Z(n13847) );
  AND U13222 ( .A(n1219), .B(n13857), .Z(n13856) );
  XOR U13223 ( .A(n13858), .B(n13859), .Z(n13844) );
  AND U13224 ( .A(n1223), .B(n13857), .Z(n13859) );
  XNOR U13225 ( .A(n13860), .B(n13858), .Z(n13857) );
  IV U13226 ( .A(n13855), .Z(n13860) );
  XOR U13227 ( .A(n13861), .B(n13862), .Z(n13855) );
  AND U13228 ( .A(n1226), .B(n13854), .Z(n13862) );
  XNOR U13229 ( .A(n13852), .B(n13861), .Z(n13854) );
  XNOR U13230 ( .A(n13863), .B(n13864), .Z(n13852) );
  AND U13231 ( .A(n1230), .B(n13865), .Z(n13864) );
  XOR U13232 ( .A(p_input[978]), .B(n13863), .Z(n13865) );
  XNOR U13233 ( .A(n13866), .B(n13867), .Z(n13863) );
  AND U13234 ( .A(n1234), .B(n13868), .Z(n13867) );
  XOR U13235 ( .A(n13869), .B(n13870), .Z(n13861) );
  AND U13236 ( .A(n1238), .B(n13871), .Z(n13870) );
  XOR U13237 ( .A(n13872), .B(n13873), .Z(n13858) );
  AND U13238 ( .A(n1242), .B(n13871), .Z(n13873) );
  XNOR U13239 ( .A(n13874), .B(n13872), .Z(n13871) );
  IV U13240 ( .A(n13869), .Z(n13874) );
  XOR U13241 ( .A(n13875), .B(n13876), .Z(n13869) );
  AND U13242 ( .A(n1245), .B(n13868), .Z(n13876) );
  XNOR U13243 ( .A(n13866), .B(n13875), .Z(n13868) );
  XNOR U13244 ( .A(n13877), .B(n13878), .Z(n13866) );
  AND U13245 ( .A(n1249), .B(n13879), .Z(n13878) );
  XOR U13246 ( .A(p_input[994]), .B(n13877), .Z(n13879) );
  XNOR U13247 ( .A(n13880), .B(n13881), .Z(n13877) );
  AND U13248 ( .A(n1253), .B(n13882), .Z(n13881) );
  XOR U13249 ( .A(n13883), .B(n13884), .Z(n13875) );
  AND U13250 ( .A(n1257), .B(n13885), .Z(n13884) );
  XOR U13251 ( .A(n13886), .B(n13887), .Z(n13872) );
  AND U13252 ( .A(n1261), .B(n13885), .Z(n13887) );
  XNOR U13253 ( .A(n13888), .B(n13886), .Z(n13885) );
  IV U13254 ( .A(n13883), .Z(n13888) );
  XOR U13255 ( .A(n13889), .B(n13890), .Z(n13883) );
  AND U13256 ( .A(n1264), .B(n13882), .Z(n13890) );
  XNOR U13257 ( .A(n13880), .B(n13889), .Z(n13882) );
  XNOR U13258 ( .A(n13891), .B(n13892), .Z(n13880) );
  AND U13259 ( .A(n1268), .B(n13893), .Z(n13892) );
  XOR U13260 ( .A(p_input[1010]), .B(n13891), .Z(n13893) );
  XNOR U13261 ( .A(n13894), .B(n13895), .Z(n13891) );
  AND U13262 ( .A(n1272), .B(n13896), .Z(n13895) );
  XOR U13263 ( .A(n13897), .B(n13898), .Z(n13889) );
  AND U13264 ( .A(n1276), .B(n13899), .Z(n13898) );
  XOR U13265 ( .A(n13900), .B(n13901), .Z(n13886) );
  AND U13266 ( .A(n1280), .B(n13899), .Z(n13901) );
  XNOR U13267 ( .A(n13902), .B(n13900), .Z(n13899) );
  IV U13268 ( .A(n13897), .Z(n13902) );
  XOR U13269 ( .A(n13903), .B(n13904), .Z(n13897) );
  AND U13270 ( .A(n1283), .B(n13896), .Z(n13904) );
  XNOR U13271 ( .A(n13894), .B(n13903), .Z(n13896) );
  XNOR U13272 ( .A(n13905), .B(n13906), .Z(n13894) );
  AND U13273 ( .A(n1287), .B(n13907), .Z(n13906) );
  XOR U13274 ( .A(p_input[1026]), .B(n13905), .Z(n13907) );
  XNOR U13275 ( .A(n13908), .B(n13909), .Z(n13905) );
  AND U13276 ( .A(n1291), .B(n13910), .Z(n13909) );
  XOR U13277 ( .A(n13911), .B(n13912), .Z(n13903) );
  AND U13278 ( .A(n1295), .B(n13913), .Z(n13912) );
  XOR U13279 ( .A(n13914), .B(n13915), .Z(n13900) );
  AND U13280 ( .A(n1299), .B(n13913), .Z(n13915) );
  XNOR U13281 ( .A(n13916), .B(n13914), .Z(n13913) );
  IV U13282 ( .A(n13911), .Z(n13916) );
  XOR U13283 ( .A(n13917), .B(n13918), .Z(n13911) );
  AND U13284 ( .A(n1302), .B(n13910), .Z(n13918) );
  XNOR U13285 ( .A(n13908), .B(n13917), .Z(n13910) );
  XNOR U13286 ( .A(n13919), .B(n13920), .Z(n13908) );
  AND U13287 ( .A(n1306), .B(n13921), .Z(n13920) );
  XOR U13288 ( .A(p_input[1042]), .B(n13919), .Z(n13921) );
  XNOR U13289 ( .A(n13922), .B(n13923), .Z(n13919) );
  AND U13290 ( .A(n1310), .B(n13924), .Z(n13923) );
  XOR U13291 ( .A(n13925), .B(n13926), .Z(n13917) );
  AND U13292 ( .A(n1314), .B(n13927), .Z(n13926) );
  XOR U13293 ( .A(n13928), .B(n13929), .Z(n13914) );
  AND U13294 ( .A(n1318), .B(n13927), .Z(n13929) );
  XNOR U13295 ( .A(n13930), .B(n13928), .Z(n13927) );
  IV U13296 ( .A(n13925), .Z(n13930) );
  XOR U13297 ( .A(n13931), .B(n13932), .Z(n13925) );
  AND U13298 ( .A(n1321), .B(n13924), .Z(n13932) );
  XNOR U13299 ( .A(n13922), .B(n13931), .Z(n13924) );
  XNOR U13300 ( .A(n13933), .B(n13934), .Z(n13922) );
  AND U13301 ( .A(n1325), .B(n13935), .Z(n13934) );
  XOR U13302 ( .A(p_input[1058]), .B(n13933), .Z(n13935) );
  XNOR U13303 ( .A(n13936), .B(n13937), .Z(n13933) );
  AND U13304 ( .A(n1329), .B(n13938), .Z(n13937) );
  XOR U13305 ( .A(n13939), .B(n13940), .Z(n13931) );
  AND U13306 ( .A(n1333), .B(n13941), .Z(n13940) );
  XOR U13307 ( .A(n13942), .B(n13943), .Z(n13928) );
  AND U13308 ( .A(n1337), .B(n13941), .Z(n13943) );
  XNOR U13309 ( .A(n13944), .B(n13942), .Z(n13941) );
  IV U13310 ( .A(n13939), .Z(n13944) );
  XOR U13311 ( .A(n13945), .B(n13946), .Z(n13939) );
  AND U13312 ( .A(n1340), .B(n13938), .Z(n13946) );
  XNOR U13313 ( .A(n13936), .B(n13945), .Z(n13938) );
  XNOR U13314 ( .A(n13947), .B(n13948), .Z(n13936) );
  AND U13315 ( .A(n1344), .B(n13949), .Z(n13948) );
  XOR U13316 ( .A(p_input[1074]), .B(n13947), .Z(n13949) );
  XNOR U13317 ( .A(n13950), .B(n13951), .Z(n13947) );
  AND U13318 ( .A(n1348), .B(n13952), .Z(n13951) );
  XOR U13319 ( .A(n13953), .B(n13954), .Z(n13945) );
  AND U13320 ( .A(n1352), .B(n13955), .Z(n13954) );
  XOR U13321 ( .A(n13956), .B(n13957), .Z(n13942) );
  AND U13322 ( .A(n1356), .B(n13955), .Z(n13957) );
  XNOR U13323 ( .A(n13958), .B(n13956), .Z(n13955) );
  IV U13324 ( .A(n13953), .Z(n13958) );
  XOR U13325 ( .A(n13959), .B(n13960), .Z(n13953) );
  AND U13326 ( .A(n1359), .B(n13952), .Z(n13960) );
  XNOR U13327 ( .A(n13950), .B(n13959), .Z(n13952) );
  XNOR U13328 ( .A(n13961), .B(n13962), .Z(n13950) );
  AND U13329 ( .A(n1363), .B(n13963), .Z(n13962) );
  XOR U13330 ( .A(p_input[1090]), .B(n13961), .Z(n13963) );
  XNOR U13331 ( .A(n13964), .B(n13965), .Z(n13961) );
  AND U13332 ( .A(n1367), .B(n13966), .Z(n13965) );
  XOR U13333 ( .A(n13967), .B(n13968), .Z(n13959) );
  AND U13334 ( .A(n1371), .B(n13969), .Z(n13968) );
  XOR U13335 ( .A(n13970), .B(n13971), .Z(n13956) );
  AND U13336 ( .A(n1375), .B(n13969), .Z(n13971) );
  XNOR U13337 ( .A(n13972), .B(n13970), .Z(n13969) );
  IV U13338 ( .A(n13967), .Z(n13972) );
  XOR U13339 ( .A(n13973), .B(n13974), .Z(n13967) );
  AND U13340 ( .A(n1378), .B(n13966), .Z(n13974) );
  XNOR U13341 ( .A(n13964), .B(n13973), .Z(n13966) );
  XNOR U13342 ( .A(n13975), .B(n13976), .Z(n13964) );
  AND U13343 ( .A(n1382), .B(n13977), .Z(n13976) );
  XOR U13344 ( .A(p_input[1106]), .B(n13975), .Z(n13977) );
  XNOR U13345 ( .A(n13978), .B(n13979), .Z(n13975) );
  AND U13346 ( .A(n1386), .B(n13980), .Z(n13979) );
  XOR U13347 ( .A(n13981), .B(n13982), .Z(n13973) );
  AND U13348 ( .A(n1390), .B(n13983), .Z(n13982) );
  XOR U13349 ( .A(n13984), .B(n13985), .Z(n13970) );
  AND U13350 ( .A(n1394), .B(n13983), .Z(n13985) );
  XNOR U13351 ( .A(n13986), .B(n13984), .Z(n13983) );
  IV U13352 ( .A(n13981), .Z(n13986) );
  XOR U13353 ( .A(n13987), .B(n13988), .Z(n13981) );
  AND U13354 ( .A(n1397), .B(n13980), .Z(n13988) );
  XNOR U13355 ( .A(n13978), .B(n13987), .Z(n13980) );
  XNOR U13356 ( .A(n13989), .B(n13990), .Z(n13978) );
  AND U13357 ( .A(n1401), .B(n13991), .Z(n13990) );
  XOR U13358 ( .A(p_input[1122]), .B(n13989), .Z(n13991) );
  XNOR U13359 ( .A(n13992), .B(n13993), .Z(n13989) );
  AND U13360 ( .A(n1405), .B(n13994), .Z(n13993) );
  XOR U13361 ( .A(n13995), .B(n13996), .Z(n13987) );
  AND U13362 ( .A(n1409), .B(n13997), .Z(n13996) );
  XOR U13363 ( .A(n13998), .B(n13999), .Z(n13984) );
  AND U13364 ( .A(n1413), .B(n13997), .Z(n13999) );
  XNOR U13365 ( .A(n14000), .B(n13998), .Z(n13997) );
  IV U13366 ( .A(n13995), .Z(n14000) );
  XOR U13367 ( .A(n14001), .B(n14002), .Z(n13995) );
  AND U13368 ( .A(n1416), .B(n13994), .Z(n14002) );
  XNOR U13369 ( .A(n13992), .B(n14001), .Z(n13994) );
  XNOR U13370 ( .A(n14003), .B(n14004), .Z(n13992) );
  AND U13371 ( .A(n1420), .B(n14005), .Z(n14004) );
  XOR U13372 ( .A(p_input[1138]), .B(n14003), .Z(n14005) );
  XNOR U13373 ( .A(n14006), .B(n14007), .Z(n14003) );
  AND U13374 ( .A(n1424), .B(n14008), .Z(n14007) );
  XOR U13375 ( .A(n14009), .B(n14010), .Z(n14001) );
  AND U13376 ( .A(n1428), .B(n14011), .Z(n14010) );
  XOR U13377 ( .A(n14012), .B(n14013), .Z(n13998) );
  AND U13378 ( .A(n1432), .B(n14011), .Z(n14013) );
  XNOR U13379 ( .A(n14014), .B(n14012), .Z(n14011) );
  IV U13380 ( .A(n14009), .Z(n14014) );
  XOR U13381 ( .A(n14015), .B(n14016), .Z(n14009) );
  AND U13382 ( .A(n1435), .B(n14008), .Z(n14016) );
  XNOR U13383 ( .A(n14006), .B(n14015), .Z(n14008) );
  XNOR U13384 ( .A(n14017), .B(n14018), .Z(n14006) );
  AND U13385 ( .A(n1439), .B(n14019), .Z(n14018) );
  XOR U13386 ( .A(p_input[1154]), .B(n14017), .Z(n14019) );
  XNOR U13387 ( .A(n14020), .B(n14021), .Z(n14017) );
  AND U13388 ( .A(n1443), .B(n14022), .Z(n14021) );
  XOR U13389 ( .A(n14023), .B(n14024), .Z(n14015) );
  AND U13390 ( .A(n1447), .B(n14025), .Z(n14024) );
  XOR U13391 ( .A(n14026), .B(n14027), .Z(n14012) );
  AND U13392 ( .A(n1451), .B(n14025), .Z(n14027) );
  XNOR U13393 ( .A(n14028), .B(n14026), .Z(n14025) );
  IV U13394 ( .A(n14023), .Z(n14028) );
  XOR U13395 ( .A(n14029), .B(n14030), .Z(n14023) );
  AND U13396 ( .A(n1454), .B(n14022), .Z(n14030) );
  XNOR U13397 ( .A(n14020), .B(n14029), .Z(n14022) );
  XNOR U13398 ( .A(n14031), .B(n14032), .Z(n14020) );
  AND U13399 ( .A(n1458), .B(n14033), .Z(n14032) );
  XOR U13400 ( .A(p_input[1170]), .B(n14031), .Z(n14033) );
  XNOR U13401 ( .A(n14034), .B(n14035), .Z(n14031) );
  AND U13402 ( .A(n1462), .B(n14036), .Z(n14035) );
  XOR U13403 ( .A(n14037), .B(n14038), .Z(n14029) );
  AND U13404 ( .A(n1466), .B(n14039), .Z(n14038) );
  XOR U13405 ( .A(n14040), .B(n14041), .Z(n14026) );
  AND U13406 ( .A(n1470), .B(n14039), .Z(n14041) );
  XNOR U13407 ( .A(n14042), .B(n14040), .Z(n14039) );
  IV U13408 ( .A(n14037), .Z(n14042) );
  XOR U13409 ( .A(n14043), .B(n14044), .Z(n14037) );
  AND U13410 ( .A(n1473), .B(n14036), .Z(n14044) );
  XNOR U13411 ( .A(n14034), .B(n14043), .Z(n14036) );
  XNOR U13412 ( .A(n14045), .B(n14046), .Z(n14034) );
  AND U13413 ( .A(n1477), .B(n14047), .Z(n14046) );
  XOR U13414 ( .A(p_input[1186]), .B(n14045), .Z(n14047) );
  XNOR U13415 ( .A(n14048), .B(n14049), .Z(n14045) );
  AND U13416 ( .A(n1481), .B(n14050), .Z(n14049) );
  XOR U13417 ( .A(n14051), .B(n14052), .Z(n14043) );
  AND U13418 ( .A(n1485), .B(n14053), .Z(n14052) );
  XOR U13419 ( .A(n14054), .B(n14055), .Z(n14040) );
  AND U13420 ( .A(n1489), .B(n14053), .Z(n14055) );
  XNOR U13421 ( .A(n14056), .B(n14054), .Z(n14053) );
  IV U13422 ( .A(n14051), .Z(n14056) );
  XOR U13423 ( .A(n14057), .B(n14058), .Z(n14051) );
  AND U13424 ( .A(n1492), .B(n14050), .Z(n14058) );
  XNOR U13425 ( .A(n14048), .B(n14057), .Z(n14050) );
  XNOR U13426 ( .A(n14059), .B(n14060), .Z(n14048) );
  AND U13427 ( .A(n1496), .B(n14061), .Z(n14060) );
  XOR U13428 ( .A(p_input[1202]), .B(n14059), .Z(n14061) );
  XNOR U13429 ( .A(n14062), .B(n14063), .Z(n14059) );
  AND U13430 ( .A(n1500), .B(n14064), .Z(n14063) );
  XOR U13431 ( .A(n14065), .B(n14066), .Z(n14057) );
  AND U13432 ( .A(n1504), .B(n14067), .Z(n14066) );
  XOR U13433 ( .A(n14068), .B(n14069), .Z(n14054) );
  AND U13434 ( .A(n1508), .B(n14067), .Z(n14069) );
  XNOR U13435 ( .A(n14070), .B(n14068), .Z(n14067) );
  IV U13436 ( .A(n14065), .Z(n14070) );
  XOR U13437 ( .A(n14071), .B(n14072), .Z(n14065) );
  AND U13438 ( .A(n1511), .B(n14064), .Z(n14072) );
  XNOR U13439 ( .A(n14062), .B(n14071), .Z(n14064) );
  XNOR U13440 ( .A(n14073), .B(n14074), .Z(n14062) );
  AND U13441 ( .A(n1515), .B(n14075), .Z(n14074) );
  XOR U13442 ( .A(p_input[1218]), .B(n14073), .Z(n14075) );
  XNOR U13443 ( .A(n14076), .B(n14077), .Z(n14073) );
  AND U13444 ( .A(n1519), .B(n14078), .Z(n14077) );
  XOR U13445 ( .A(n14079), .B(n14080), .Z(n14071) );
  AND U13446 ( .A(n1523), .B(n14081), .Z(n14080) );
  XOR U13447 ( .A(n14082), .B(n14083), .Z(n14068) );
  AND U13448 ( .A(n1527), .B(n14081), .Z(n14083) );
  XNOR U13449 ( .A(n14084), .B(n14082), .Z(n14081) );
  IV U13450 ( .A(n14079), .Z(n14084) );
  XOR U13451 ( .A(n14085), .B(n14086), .Z(n14079) );
  AND U13452 ( .A(n1530), .B(n14078), .Z(n14086) );
  XNOR U13453 ( .A(n14076), .B(n14085), .Z(n14078) );
  XNOR U13454 ( .A(n14087), .B(n14088), .Z(n14076) );
  AND U13455 ( .A(n1534), .B(n14089), .Z(n14088) );
  XOR U13456 ( .A(p_input[1234]), .B(n14087), .Z(n14089) );
  XNOR U13457 ( .A(n14090), .B(n14091), .Z(n14087) );
  AND U13458 ( .A(n1538), .B(n14092), .Z(n14091) );
  XOR U13459 ( .A(n14093), .B(n14094), .Z(n14085) );
  AND U13460 ( .A(n1542), .B(n14095), .Z(n14094) );
  XOR U13461 ( .A(n14096), .B(n14097), .Z(n14082) );
  AND U13462 ( .A(n1546), .B(n14095), .Z(n14097) );
  XNOR U13463 ( .A(n14098), .B(n14096), .Z(n14095) );
  IV U13464 ( .A(n14093), .Z(n14098) );
  XOR U13465 ( .A(n14099), .B(n14100), .Z(n14093) );
  AND U13466 ( .A(n1549), .B(n14092), .Z(n14100) );
  XNOR U13467 ( .A(n14090), .B(n14099), .Z(n14092) );
  XNOR U13468 ( .A(n14101), .B(n14102), .Z(n14090) );
  AND U13469 ( .A(n1553), .B(n14103), .Z(n14102) );
  XOR U13470 ( .A(p_input[1250]), .B(n14101), .Z(n14103) );
  XNOR U13471 ( .A(n14104), .B(n14105), .Z(n14101) );
  AND U13472 ( .A(n1557), .B(n14106), .Z(n14105) );
  XOR U13473 ( .A(n14107), .B(n14108), .Z(n14099) );
  AND U13474 ( .A(n1561), .B(n14109), .Z(n14108) );
  XOR U13475 ( .A(n14110), .B(n14111), .Z(n14096) );
  AND U13476 ( .A(n1565), .B(n14109), .Z(n14111) );
  XNOR U13477 ( .A(n14112), .B(n14110), .Z(n14109) );
  IV U13478 ( .A(n14107), .Z(n14112) );
  XOR U13479 ( .A(n14113), .B(n14114), .Z(n14107) );
  AND U13480 ( .A(n1568), .B(n14106), .Z(n14114) );
  XNOR U13481 ( .A(n14104), .B(n14113), .Z(n14106) );
  XNOR U13482 ( .A(n14115), .B(n14116), .Z(n14104) );
  AND U13483 ( .A(n1572), .B(n14117), .Z(n14116) );
  XOR U13484 ( .A(p_input[1266]), .B(n14115), .Z(n14117) );
  XNOR U13485 ( .A(n14118), .B(n14119), .Z(n14115) );
  AND U13486 ( .A(n1576), .B(n14120), .Z(n14119) );
  XOR U13487 ( .A(n14121), .B(n14122), .Z(n14113) );
  AND U13488 ( .A(n1580), .B(n14123), .Z(n14122) );
  XOR U13489 ( .A(n14124), .B(n14125), .Z(n14110) );
  AND U13490 ( .A(n1584), .B(n14123), .Z(n14125) );
  XNOR U13491 ( .A(n14126), .B(n14124), .Z(n14123) );
  IV U13492 ( .A(n14121), .Z(n14126) );
  XOR U13493 ( .A(n14127), .B(n14128), .Z(n14121) );
  AND U13494 ( .A(n1587), .B(n14120), .Z(n14128) );
  XNOR U13495 ( .A(n14118), .B(n14127), .Z(n14120) );
  XNOR U13496 ( .A(n14129), .B(n14130), .Z(n14118) );
  AND U13497 ( .A(n1591), .B(n14131), .Z(n14130) );
  XOR U13498 ( .A(p_input[1282]), .B(n14129), .Z(n14131) );
  XNOR U13499 ( .A(n14132), .B(n14133), .Z(n14129) );
  AND U13500 ( .A(n1595), .B(n14134), .Z(n14133) );
  XOR U13501 ( .A(n14135), .B(n14136), .Z(n14127) );
  AND U13502 ( .A(n1599), .B(n14137), .Z(n14136) );
  XOR U13503 ( .A(n14138), .B(n14139), .Z(n14124) );
  AND U13504 ( .A(n1603), .B(n14137), .Z(n14139) );
  XNOR U13505 ( .A(n14140), .B(n14138), .Z(n14137) );
  IV U13506 ( .A(n14135), .Z(n14140) );
  XOR U13507 ( .A(n14141), .B(n14142), .Z(n14135) );
  AND U13508 ( .A(n1606), .B(n14134), .Z(n14142) );
  XNOR U13509 ( .A(n14132), .B(n14141), .Z(n14134) );
  XNOR U13510 ( .A(n14143), .B(n14144), .Z(n14132) );
  AND U13511 ( .A(n1610), .B(n14145), .Z(n14144) );
  XOR U13512 ( .A(p_input[1298]), .B(n14143), .Z(n14145) );
  XNOR U13513 ( .A(n14146), .B(n14147), .Z(n14143) );
  AND U13514 ( .A(n1614), .B(n14148), .Z(n14147) );
  XOR U13515 ( .A(n14149), .B(n14150), .Z(n14141) );
  AND U13516 ( .A(n1618), .B(n14151), .Z(n14150) );
  XOR U13517 ( .A(n14152), .B(n14153), .Z(n14138) );
  AND U13518 ( .A(n1622), .B(n14151), .Z(n14153) );
  XNOR U13519 ( .A(n14154), .B(n14152), .Z(n14151) );
  IV U13520 ( .A(n14149), .Z(n14154) );
  XOR U13521 ( .A(n14155), .B(n14156), .Z(n14149) );
  AND U13522 ( .A(n1625), .B(n14148), .Z(n14156) );
  XNOR U13523 ( .A(n14146), .B(n14155), .Z(n14148) );
  XNOR U13524 ( .A(n14157), .B(n14158), .Z(n14146) );
  AND U13525 ( .A(n1629), .B(n14159), .Z(n14158) );
  XOR U13526 ( .A(p_input[1314]), .B(n14157), .Z(n14159) );
  XNOR U13527 ( .A(n14160), .B(n14161), .Z(n14157) );
  AND U13528 ( .A(n1633), .B(n14162), .Z(n14161) );
  XOR U13529 ( .A(n14163), .B(n14164), .Z(n14155) );
  AND U13530 ( .A(n1637), .B(n14165), .Z(n14164) );
  XOR U13531 ( .A(n14166), .B(n14167), .Z(n14152) );
  AND U13532 ( .A(n1641), .B(n14165), .Z(n14167) );
  XNOR U13533 ( .A(n14168), .B(n14166), .Z(n14165) );
  IV U13534 ( .A(n14163), .Z(n14168) );
  XOR U13535 ( .A(n14169), .B(n14170), .Z(n14163) );
  AND U13536 ( .A(n1644), .B(n14162), .Z(n14170) );
  XNOR U13537 ( .A(n14160), .B(n14169), .Z(n14162) );
  XNOR U13538 ( .A(n14171), .B(n14172), .Z(n14160) );
  AND U13539 ( .A(n1648), .B(n14173), .Z(n14172) );
  XOR U13540 ( .A(p_input[1330]), .B(n14171), .Z(n14173) );
  XNOR U13541 ( .A(n14174), .B(n14175), .Z(n14171) );
  AND U13542 ( .A(n1652), .B(n14176), .Z(n14175) );
  XOR U13543 ( .A(n14177), .B(n14178), .Z(n14169) );
  AND U13544 ( .A(n1656), .B(n14179), .Z(n14178) );
  XOR U13545 ( .A(n14180), .B(n14181), .Z(n14166) );
  AND U13546 ( .A(n1660), .B(n14179), .Z(n14181) );
  XNOR U13547 ( .A(n14182), .B(n14180), .Z(n14179) );
  IV U13548 ( .A(n14177), .Z(n14182) );
  XOR U13549 ( .A(n14183), .B(n14184), .Z(n14177) );
  AND U13550 ( .A(n1663), .B(n14176), .Z(n14184) );
  XNOR U13551 ( .A(n14174), .B(n14183), .Z(n14176) );
  XNOR U13552 ( .A(n14185), .B(n14186), .Z(n14174) );
  AND U13553 ( .A(n1667), .B(n14187), .Z(n14186) );
  XOR U13554 ( .A(p_input[1346]), .B(n14185), .Z(n14187) );
  XNOR U13555 ( .A(n14188), .B(n14189), .Z(n14185) );
  AND U13556 ( .A(n1671), .B(n14190), .Z(n14189) );
  XOR U13557 ( .A(n14191), .B(n14192), .Z(n14183) );
  AND U13558 ( .A(n1675), .B(n14193), .Z(n14192) );
  XOR U13559 ( .A(n14194), .B(n14195), .Z(n14180) );
  AND U13560 ( .A(n1679), .B(n14193), .Z(n14195) );
  XNOR U13561 ( .A(n14196), .B(n14194), .Z(n14193) );
  IV U13562 ( .A(n14191), .Z(n14196) );
  XOR U13563 ( .A(n14197), .B(n14198), .Z(n14191) );
  AND U13564 ( .A(n1682), .B(n14190), .Z(n14198) );
  XNOR U13565 ( .A(n14188), .B(n14197), .Z(n14190) );
  XNOR U13566 ( .A(n14199), .B(n14200), .Z(n14188) );
  AND U13567 ( .A(n1686), .B(n14201), .Z(n14200) );
  XOR U13568 ( .A(p_input[1362]), .B(n14199), .Z(n14201) );
  XNOR U13569 ( .A(n14202), .B(n14203), .Z(n14199) );
  AND U13570 ( .A(n1690), .B(n14204), .Z(n14203) );
  XOR U13571 ( .A(n14205), .B(n14206), .Z(n14197) );
  AND U13572 ( .A(n1694), .B(n14207), .Z(n14206) );
  XOR U13573 ( .A(n14208), .B(n14209), .Z(n14194) );
  AND U13574 ( .A(n1698), .B(n14207), .Z(n14209) );
  XNOR U13575 ( .A(n14210), .B(n14208), .Z(n14207) );
  IV U13576 ( .A(n14205), .Z(n14210) );
  XOR U13577 ( .A(n14211), .B(n14212), .Z(n14205) );
  AND U13578 ( .A(n1701), .B(n14204), .Z(n14212) );
  XNOR U13579 ( .A(n14202), .B(n14211), .Z(n14204) );
  XNOR U13580 ( .A(n14213), .B(n14214), .Z(n14202) );
  AND U13581 ( .A(n1705), .B(n14215), .Z(n14214) );
  XOR U13582 ( .A(p_input[1378]), .B(n14213), .Z(n14215) );
  XNOR U13583 ( .A(n14216), .B(n14217), .Z(n14213) );
  AND U13584 ( .A(n1709), .B(n14218), .Z(n14217) );
  XOR U13585 ( .A(n14219), .B(n14220), .Z(n14211) );
  AND U13586 ( .A(n1713), .B(n14221), .Z(n14220) );
  XOR U13587 ( .A(n14222), .B(n14223), .Z(n14208) );
  AND U13588 ( .A(n1717), .B(n14221), .Z(n14223) );
  XNOR U13589 ( .A(n14224), .B(n14222), .Z(n14221) );
  IV U13590 ( .A(n14219), .Z(n14224) );
  XOR U13591 ( .A(n14225), .B(n14226), .Z(n14219) );
  AND U13592 ( .A(n1720), .B(n14218), .Z(n14226) );
  XNOR U13593 ( .A(n14216), .B(n14225), .Z(n14218) );
  XNOR U13594 ( .A(n14227), .B(n14228), .Z(n14216) );
  AND U13595 ( .A(n1724), .B(n14229), .Z(n14228) );
  XOR U13596 ( .A(p_input[1394]), .B(n14227), .Z(n14229) );
  XNOR U13597 ( .A(n14230), .B(n14231), .Z(n14227) );
  AND U13598 ( .A(n1728), .B(n14232), .Z(n14231) );
  XOR U13599 ( .A(n14233), .B(n14234), .Z(n14225) );
  AND U13600 ( .A(n1732), .B(n14235), .Z(n14234) );
  XOR U13601 ( .A(n14236), .B(n14237), .Z(n14222) );
  AND U13602 ( .A(n1736), .B(n14235), .Z(n14237) );
  XNOR U13603 ( .A(n14238), .B(n14236), .Z(n14235) );
  IV U13604 ( .A(n14233), .Z(n14238) );
  XOR U13605 ( .A(n14239), .B(n14240), .Z(n14233) );
  AND U13606 ( .A(n1739), .B(n14232), .Z(n14240) );
  XNOR U13607 ( .A(n14230), .B(n14239), .Z(n14232) );
  XNOR U13608 ( .A(n14241), .B(n14242), .Z(n14230) );
  AND U13609 ( .A(n1743), .B(n14243), .Z(n14242) );
  XOR U13610 ( .A(p_input[1410]), .B(n14241), .Z(n14243) );
  XNOR U13611 ( .A(n14244), .B(n14245), .Z(n14241) );
  AND U13612 ( .A(n1747), .B(n14246), .Z(n14245) );
  XOR U13613 ( .A(n14247), .B(n14248), .Z(n14239) );
  AND U13614 ( .A(n1751), .B(n14249), .Z(n14248) );
  XOR U13615 ( .A(n14250), .B(n14251), .Z(n14236) );
  AND U13616 ( .A(n1755), .B(n14249), .Z(n14251) );
  XNOR U13617 ( .A(n14252), .B(n14250), .Z(n14249) );
  IV U13618 ( .A(n14247), .Z(n14252) );
  XOR U13619 ( .A(n14253), .B(n14254), .Z(n14247) );
  AND U13620 ( .A(n1758), .B(n14246), .Z(n14254) );
  XNOR U13621 ( .A(n14244), .B(n14253), .Z(n14246) );
  XNOR U13622 ( .A(n14255), .B(n14256), .Z(n14244) );
  AND U13623 ( .A(n1762), .B(n14257), .Z(n14256) );
  XOR U13624 ( .A(p_input[1426]), .B(n14255), .Z(n14257) );
  XNOR U13625 ( .A(n14258), .B(n14259), .Z(n14255) );
  AND U13626 ( .A(n1766), .B(n14260), .Z(n14259) );
  XOR U13627 ( .A(n14261), .B(n14262), .Z(n14253) );
  AND U13628 ( .A(n1770), .B(n14263), .Z(n14262) );
  XOR U13629 ( .A(n14264), .B(n14265), .Z(n14250) );
  AND U13630 ( .A(n1774), .B(n14263), .Z(n14265) );
  XNOR U13631 ( .A(n14266), .B(n14264), .Z(n14263) );
  IV U13632 ( .A(n14261), .Z(n14266) );
  XOR U13633 ( .A(n14267), .B(n14268), .Z(n14261) );
  AND U13634 ( .A(n1777), .B(n14260), .Z(n14268) );
  XNOR U13635 ( .A(n14258), .B(n14267), .Z(n14260) );
  XNOR U13636 ( .A(n14269), .B(n14270), .Z(n14258) );
  AND U13637 ( .A(n1781), .B(n14271), .Z(n14270) );
  XOR U13638 ( .A(p_input[1442]), .B(n14269), .Z(n14271) );
  XNOR U13639 ( .A(n14272), .B(n14273), .Z(n14269) );
  AND U13640 ( .A(n1785), .B(n14274), .Z(n14273) );
  XOR U13641 ( .A(n14275), .B(n14276), .Z(n14267) );
  AND U13642 ( .A(n1789), .B(n14277), .Z(n14276) );
  XOR U13643 ( .A(n14278), .B(n14279), .Z(n14264) );
  AND U13644 ( .A(n1793), .B(n14277), .Z(n14279) );
  XNOR U13645 ( .A(n14280), .B(n14278), .Z(n14277) );
  IV U13646 ( .A(n14275), .Z(n14280) );
  XOR U13647 ( .A(n14281), .B(n14282), .Z(n14275) );
  AND U13648 ( .A(n1796), .B(n14274), .Z(n14282) );
  XNOR U13649 ( .A(n14272), .B(n14281), .Z(n14274) );
  XNOR U13650 ( .A(n14283), .B(n14284), .Z(n14272) );
  AND U13651 ( .A(n1800), .B(n14285), .Z(n14284) );
  XOR U13652 ( .A(p_input[1458]), .B(n14283), .Z(n14285) );
  XNOR U13653 ( .A(n14286), .B(n14287), .Z(n14283) );
  AND U13654 ( .A(n1804), .B(n14288), .Z(n14287) );
  XOR U13655 ( .A(n14289), .B(n14290), .Z(n14281) );
  AND U13656 ( .A(n1808), .B(n14291), .Z(n14290) );
  XOR U13657 ( .A(n14292), .B(n14293), .Z(n14278) );
  AND U13658 ( .A(n1812), .B(n14291), .Z(n14293) );
  XNOR U13659 ( .A(n14294), .B(n14292), .Z(n14291) );
  IV U13660 ( .A(n14289), .Z(n14294) );
  XOR U13661 ( .A(n14295), .B(n14296), .Z(n14289) );
  AND U13662 ( .A(n1815), .B(n14288), .Z(n14296) );
  XNOR U13663 ( .A(n14286), .B(n14295), .Z(n14288) );
  XNOR U13664 ( .A(n14297), .B(n14298), .Z(n14286) );
  AND U13665 ( .A(n1819), .B(n14299), .Z(n14298) );
  XOR U13666 ( .A(p_input[1474]), .B(n14297), .Z(n14299) );
  XNOR U13667 ( .A(n14300), .B(n14301), .Z(n14297) );
  AND U13668 ( .A(n1823), .B(n14302), .Z(n14301) );
  XOR U13669 ( .A(n14303), .B(n14304), .Z(n14295) );
  AND U13670 ( .A(n1827), .B(n14305), .Z(n14304) );
  XOR U13671 ( .A(n14306), .B(n14307), .Z(n14292) );
  AND U13672 ( .A(n1831), .B(n14305), .Z(n14307) );
  XNOR U13673 ( .A(n14308), .B(n14306), .Z(n14305) );
  IV U13674 ( .A(n14303), .Z(n14308) );
  XOR U13675 ( .A(n14309), .B(n14310), .Z(n14303) );
  AND U13676 ( .A(n1834), .B(n14302), .Z(n14310) );
  XNOR U13677 ( .A(n14300), .B(n14309), .Z(n14302) );
  XNOR U13678 ( .A(n14311), .B(n14312), .Z(n14300) );
  AND U13679 ( .A(n1838), .B(n14313), .Z(n14312) );
  XOR U13680 ( .A(p_input[1490]), .B(n14311), .Z(n14313) );
  XNOR U13681 ( .A(n14314), .B(n14315), .Z(n14311) );
  AND U13682 ( .A(n1842), .B(n14316), .Z(n14315) );
  XOR U13683 ( .A(n14317), .B(n14318), .Z(n14309) );
  AND U13684 ( .A(n1846), .B(n14319), .Z(n14318) );
  XOR U13685 ( .A(n14320), .B(n14321), .Z(n14306) );
  AND U13686 ( .A(n1850), .B(n14319), .Z(n14321) );
  XNOR U13687 ( .A(n14322), .B(n14320), .Z(n14319) );
  IV U13688 ( .A(n14317), .Z(n14322) );
  XOR U13689 ( .A(n14323), .B(n14324), .Z(n14317) );
  AND U13690 ( .A(n1853), .B(n14316), .Z(n14324) );
  XNOR U13691 ( .A(n14314), .B(n14323), .Z(n14316) );
  XNOR U13692 ( .A(n14325), .B(n14326), .Z(n14314) );
  AND U13693 ( .A(n1857), .B(n14327), .Z(n14326) );
  XOR U13694 ( .A(p_input[1506]), .B(n14325), .Z(n14327) );
  XNOR U13695 ( .A(n14328), .B(n14329), .Z(n14325) );
  AND U13696 ( .A(n1861), .B(n14330), .Z(n14329) );
  XOR U13697 ( .A(n14331), .B(n14332), .Z(n14323) );
  AND U13698 ( .A(n1865), .B(n14333), .Z(n14332) );
  XOR U13699 ( .A(n14334), .B(n14335), .Z(n14320) );
  AND U13700 ( .A(n1869), .B(n14333), .Z(n14335) );
  XNOR U13701 ( .A(n14336), .B(n14334), .Z(n14333) );
  IV U13702 ( .A(n14331), .Z(n14336) );
  XOR U13703 ( .A(n14337), .B(n14338), .Z(n14331) );
  AND U13704 ( .A(n1872), .B(n14330), .Z(n14338) );
  XNOR U13705 ( .A(n14328), .B(n14337), .Z(n14330) );
  XNOR U13706 ( .A(n14339), .B(n14340), .Z(n14328) );
  AND U13707 ( .A(n1876), .B(n14341), .Z(n14340) );
  XOR U13708 ( .A(p_input[1522]), .B(n14339), .Z(n14341) );
  XNOR U13709 ( .A(n14342), .B(n14343), .Z(n14339) );
  AND U13710 ( .A(n1880), .B(n14344), .Z(n14343) );
  XOR U13711 ( .A(n14345), .B(n14346), .Z(n14337) );
  AND U13712 ( .A(n1884), .B(n14347), .Z(n14346) );
  XOR U13713 ( .A(n14348), .B(n14349), .Z(n14334) );
  AND U13714 ( .A(n1888), .B(n14347), .Z(n14349) );
  XNOR U13715 ( .A(n14350), .B(n14348), .Z(n14347) );
  IV U13716 ( .A(n14345), .Z(n14350) );
  XOR U13717 ( .A(n14351), .B(n14352), .Z(n14345) );
  AND U13718 ( .A(n1891), .B(n14344), .Z(n14352) );
  XNOR U13719 ( .A(n14342), .B(n14351), .Z(n14344) );
  XNOR U13720 ( .A(n14353), .B(n14354), .Z(n14342) );
  AND U13721 ( .A(n1895), .B(n14355), .Z(n14354) );
  XOR U13722 ( .A(p_input[1538]), .B(n14353), .Z(n14355) );
  XNOR U13723 ( .A(n14356), .B(n14357), .Z(n14353) );
  AND U13724 ( .A(n1899), .B(n14358), .Z(n14357) );
  XOR U13725 ( .A(n14359), .B(n14360), .Z(n14351) );
  AND U13726 ( .A(n1903), .B(n14361), .Z(n14360) );
  XOR U13727 ( .A(n14362), .B(n14363), .Z(n14348) );
  AND U13728 ( .A(n1907), .B(n14361), .Z(n14363) );
  XNOR U13729 ( .A(n14364), .B(n14362), .Z(n14361) );
  IV U13730 ( .A(n14359), .Z(n14364) );
  XOR U13731 ( .A(n14365), .B(n14366), .Z(n14359) );
  AND U13732 ( .A(n1910), .B(n14358), .Z(n14366) );
  XNOR U13733 ( .A(n14356), .B(n14365), .Z(n14358) );
  XNOR U13734 ( .A(n14367), .B(n14368), .Z(n14356) );
  AND U13735 ( .A(n1914), .B(n14369), .Z(n14368) );
  XOR U13736 ( .A(p_input[1554]), .B(n14367), .Z(n14369) );
  XNOR U13737 ( .A(n14370), .B(n14371), .Z(n14367) );
  AND U13738 ( .A(n1918), .B(n14372), .Z(n14371) );
  XOR U13739 ( .A(n14373), .B(n14374), .Z(n14365) );
  AND U13740 ( .A(n1922), .B(n14375), .Z(n14374) );
  XOR U13741 ( .A(n14376), .B(n14377), .Z(n14362) );
  AND U13742 ( .A(n1926), .B(n14375), .Z(n14377) );
  XNOR U13743 ( .A(n14378), .B(n14376), .Z(n14375) );
  IV U13744 ( .A(n14373), .Z(n14378) );
  XOR U13745 ( .A(n14379), .B(n14380), .Z(n14373) );
  AND U13746 ( .A(n1929), .B(n14372), .Z(n14380) );
  XNOR U13747 ( .A(n14370), .B(n14379), .Z(n14372) );
  XNOR U13748 ( .A(n14381), .B(n14382), .Z(n14370) );
  AND U13749 ( .A(n1933), .B(n14383), .Z(n14382) );
  XOR U13750 ( .A(p_input[1570]), .B(n14381), .Z(n14383) );
  XNOR U13751 ( .A(n14384), .B(n14385), .Z(n14381) );
  AND U13752 ( .A(n1937), .B(n14386), .Z(n14385) );
  XOR U13753 ( .A(n14387), .B(n14388), .Z(n14379) );
  AND U13754 ( .A(n1941), .B(n14389), .Z(n14388) );
  XOR U13755 ( .A(n14390), .B(n14391), .Z(n14376) );
  AND U13756 ( .A(n1945), .B(n14389), .Z(n14391) );
  XNOR U13757 ( .A(n14392), .B(n14390), .Z(n14389) );
  IV U13758 ( .A(n14387), .Z(n14392) );
  XOR U13759 ( .A(n14393), .B(n14394), .Z(n14387) );
  AND U13760 ( .A(n1948), .B(n14386), .Z(n14394) );
  XNOR U13761 ( .A(n14384), .B(n14393), .Z(n14386) );
  XNOR U13762 ( .A(n14395), .B(n14396), .Z(n14384) );
  AND U13763 ( .A(n1952), .B(n14397), .Z(n14396) );
  XOR U13764 ( .A(p_input[1586]), .B(n14395), .Z(n14397) );
  XNOR U13765 ( .A(n14398), .B(n14399), .Z(n14395) );
  AND U13766 ( .A(n1956), .B(n14400), .Z(n14399) );
  XOR U13767 ( .A(n14401), .B(n14402), .Z(n14393) );
  AND U13768 ( .A(n1960), .B(n14403), .Z(n14402) );
  XOR U13769 ( .A(n14404), .B(n14405), .Z(n14390) );
  AND U13770 ( .A(n1964), .B(n14403), .Z(n14405) );
  XNOR U13771 ( .A(n14406), .B(n14404), .Z(n14403) );
  IV U13772 ( .A(n14401), .Z(n14406) );
  XOR U13773 ( .A(n14407), .B(n14408), .Z(n14401) );
  AND U13774 ( .A(n1967), .B(n14400), .Z(n14408) );
  XNOR U13775 ( .A(n14398), .B(n14407), .Z(n14400) );
  XNOR U13776 ( .A(n14409), .B(n14410), .Z(n14398) );
  AND U13777 ( .A(n1971), .B(n14411), .Z(n14410) );
  XOR U13778 ( .A(p_input[1602]), .B(n14409), .Z(n14411) );
  XNOR U13779 ( .A(n14412), .B(n14413), .Z(n14409) );
  AND U13780 ( .A(n1975), .B(n14414), .Z(n14413) );
  XOR U13781 ( .A(n14415), .B(n14416), .Z(n14407) );
  AND U13782 ( .A(n1979), .B(n14417), .Z(n14416) );
  XOR U13783 ( .A(n14418), .B(n14419), .Z(n14404) );
  AND U13784 ( .A(n1983), .B(n14417), .Z(n14419) );
  XNOR U13785 ( .A(n14420), .B(n14418), .Z(n14417) );
  IV U13786 ( .A(n14415), .Z(n14420) );
  XOR U13787 ( .A(n14421), .B(n14422), .Z(n14415) );
  AND U13788 ( .A(n1986), .B(n14414), .Z(n14422) );
  XNOR U13789 ( .A(n14412), .B(n14421), .Z(n14414) );
  XNOR U13790 ( .A(n14423), .B(n14424), .Z(n14412) );
  AND U13791 ( .A(n1990), .B(n14425), .Z(n14424) );
  XOR U13792 ( .A(p_input[1618]), .B(n14423), .Z(n14425) );
  XNOR U13793 ( .A(n14426), .B(n14427), .Z(n14423) );
  AND U13794 ( .A(n1994), .B(n14428), .Z(n14427) );
  XOR U13795 ( .A(n14429), .B(n14430), .Z(n14421) );
  AND U13796 ( .A(n1998), .B(n14431), .Z(n14430) );
  XOR U13797 ( .A(n14432), .B(n14433), .Z(n14418) );
  AND U13798 ( .A(n2002), .B(n14431), .Z(n14433) );
  XNOR U13799 ( .A(n14434), .B(n14432), .Z(n14431) );
  IV U13800 ( .A(n14429), .Z(n14434) );
  XOR U13801 ( .A(n14435), .B(n14436), .Z(n14429) );
  AND U13802 ( .A(n2005), .B(n14428), .Z(n14436) );
  XNOR U13803 ( .A(n14426), .B(n14435), .Z(n14428) );
  XNOR U13804 ( .A(n14437), .B(n14438), .Z(n14426) );
  AND U13805 ( .A(n2009), .B(n14439), .Z(n14438) );
  XOR U13806 ( .A(p_input[1634]), .B(n14437), .Z(n14439) );
  XNOR U13807 ( .A(n14440), .B(n14441), .Z(n14437) );
  AND U13808 ( .A(n2013), .B(n14442), .Z(n14441) );
  XOR U13809 ( .A(n14443), .B(n14444), .Z(n14435) );
  AND U13810 ( .A(n2017), .B(n14445), .Z(n14444) );
  XOR U13811 ( .A(n14446), .B(n14447), .Z(n14432) );
  AND U13812 ( .A(n2021), .B(n14445), .Z(n14447) );
  XNOR U13813 ( .A(n14448), .B(n14446), .Z(n14445) );
  IV U13814 ( .A(n14443), .Z(n14448) );
  XOR U13815 ( .A(n14449), .B(n14450), .Z(n14443) );
  AND U13816 ( .A(n2024), .B(n14442), .Z(n14450) );
  XNOR U13817 ( .A(n14440), .B(n14449), .Z(n14442) );
  XNOR U13818 ( .A(n14451), .B(n14452), .Z(n14440) );
  AND U13819 ( .A(n2028), .B(n14453), .Z(n14452) );
  XOR U13820 ( .A(p_input[1650]), .B(n14451), .Z(n14453) );
  XNOR U13821 ( .A(n14454), .B(n14455), .Z(n14451) );
  AND U13822 ( .A(n2032), .B(n14456), .Z(n14455) );
  XOR U13823 ( .A(n14457), .B(n14458), .Z(n14449) );
  AND U13824 ( .A(n2036), .B(n14459), .Z(n14458) );
  XOR U13825 ( .A(n14460), .B(n14461), .Z(n14446) );
  AND U13826 ( .A(n2040), .B(n14459), .Z(n14461) );
  XNOR U13827 ( .A(n14462), .B(n14460), .Z(n14459) );
  IV U13828 ( .A(n14457), .Z(n14462) );
  XOR U13829 ( .A(n14463), .B(n14464), .Z(n14457) );
  AND U13830 ( .A(n2043), .B(n14456), .Z(n14464) );
  XNOR U13831 ( .A(n14454), .B(n14463), .Z(n14456) );
  XNOR U13832 ( .A(n14465), .B(n14466), .Z(n14454) );
  AND U13833 ( .A(n2047), .B(n14467), .Z(n14466) );
  XOR U13834 ( .A(p_input[1666]), .B(n14465), .Z(n14467) );
  XNOR U13835 ( .A(n14468), .B(n14469), .Z(n14465) );
  AND U13836 ( .A(n2051), .B(n14470), .Z(n14469) );
  XOR U13837 ( .A(n14471), .B(n14472), .Z(n14463) );
  AND U13838 ( .A(n2055), .B(n14473), .Z(n14472) );
  XOR U13839 ( .A(n14474), .B(n14475), .Z(n14460) );
  AND U13840 ( .A(n2059), .B(n14473), .Z(n14475) );
  XNOR U13841 ( .A(n14476), .B(n14474), .Z(n14473) );
  IV U13842 ( .A(n14471), .Z(n14476) );
  XOR U13843 ( .A(n14477), .B(n14478), .Z(n14471) );
  AND U13844 ( .A(n2062), .B(n14470), .Z(n14478) );
  XNOR U13845 ( .A(n14468), .B(n14477), .Z(n14470) );
  XNOR U13846 ( .A(n14479), .B(n14480), .Z(n14468) );
  AND U13847 ( .A(n2066), .B(n14481), .Z(n14480) );
  XOR U13848 ( .A(p_input[1682]), .B(n14479), .Z(n14481) );
  XNOR U13849 ( .A(n14482), .B(n14483), .Z(n14479) );
  AND U13850 ( .A(n2070), .B(n14484), .Z(n14483) );
  XOR U13851 ( .A(n14485), .B(n14486), .Z(n14477) );
  AND U13852 ( .A(n2074), .B(n14487), .Z(n14486) );
  XOR U13853 ( .A(n14488), .B(n14489), .Z(n14474) );
  AND U13854 ( .A(n2078), .B(n14487), .Z(n14489) );
  XNOR U13855 ( .A(n14490), .B(n14488), .Z(n14487) );
  IV U13856 ( .A(n14485), .Z(n14490) );
  XOR U13857 ( .A(n14491), .B(n14492), .Z(n14485) );
  AND U13858 ( .A(n2081), .B(n14484), .Z(n14492) );
  XNOR U13859 ( .A(n14482), .B(n14491), .Z(n14484) );
  XNOR U13860 ( .A(n14493), .B(n14494), .Z(n14482) );
  AND U13861 ( .A(n2085), .B(n14495), .Z(n14494) );
  XOR U13862 ( .A(p_input[1698]), .B(n14493), .Z(n14495) );
  XNOR U13863 ( .A(n14496), .B(n14497), .Z(n14493) );
  AND U13864 ( .A(n2089), .B(n14498), .Z(n14497) );
  XOR U13865 ( .A(n14499), .B(n14500), .Z(n14491) );
  AND U13866 ( .A(n2093), .B(n14501), .Z(n14500) );
  XOR U13867 ( .A(n14502), .B(n14503), .Z(n14488) );
  AND U13868 ( .A(n2097), .B(n14501), .Z(n14503) );
  XNOR U13869 ( .A(n14504), .B(n14502), .Z(n14501) );
  IV U13870 ( .A(n14499), .Z(n14504) );
  XOR U13871 ( .A(n14505), .B(n14506), .Z(n14499) );
  AND U13872 ( .A(n2100), .B(n14498), .Z(n14506) );
  XNOR U13873 ( .A(n14496), .B(n14505), .Z(n14498) );
  XNOR U13874 ( .A(n14507), .B(n14508), .Z(n14496) );
  AND U13875 ( .A(n2104), .B(n14509), .Z(n14508) );
  XOR U13876 ( .A(p_input[1714]), .B(n14507), .Z(n14509) );
  XNOR U13877 ( .A(n14510), .B(n14511), .Z(n14507) );
  AND U13878 ( .A(n2108), .B(n14512), .Z(n14511) );
  XOR U13879 ( .A(n14513), .B(n14514), .Z(n14505) );
  AND U13880 ( .A(n2112), .B(n14515), .Z(n14514) );
  XOR U13881 ( .A(n14516), .B(n14517), .Z(n14502) );
  AND U13882 ( .A(n2116), .B(n14515), .Z(n14517) );
  XNOR U13883 ( .A(n14518), .B(n14516), .Z(n14515) );
  IV U13884 ( .A(n14513), .Z(n14518) );
  XOR U13885 ( .A(n14519), .B(n14520), .Z(n14513) );
  AND U13886 ( .A(n2119), .B(n14512), .Z(n14520) );
  XNOR U13887 ( .A(n14510), .B(n14519), .Z(n14512) );
  XNOR U13888 ( .A(n14521), .B(n14522), .Z(n14510) );
  AND U13889 ( .A(n2123), .B(n14523), .Z(n14522) );
  XOR U13890 ( .A(p_input[1730]), .B(n14521), .Z(n14523) );
  XNOR U13891 ( .A(n14524), .B(n14525), .Z(n14521) );
  AND U13892 ( .A(n2127), .B(n14526), .Z(n14525) );
  XOR U13893 ( .A(n14527), .B(n14528), .Z(n14519) );
  AND U13894 ( .A(n2131), .B(n14529), .Z(n14528) );
  XOR U13895 ( .A(n14530), .B(n14531), .Z(n14516) );
  AND U13896 ( .A(n2135), .B(n14529), .Z(n14531) );
  XNOR U13897 ( .A(n14532), .B(n14530), .Z(n14529) );
  IV U13898 ( .A(n14527), .Z(n14532) );
  XOR U13899 ( .A(n14533), .B(n14534), .Z(n14527) );
  AND U13900 ( .A(n2138), .B(n14526), .Z(n14534) );
  XNOR U13901 ( .A(n14524), .B(n14533), .Z(n14526) );
  XNOR U13902 ( .A(n14535), .B(n14536), .Z(n14524) );
  AND U13903 ( .A(n2142), .B(n14537), .Z(n14536) );
  XOR U13904 ( .A(p_input[1746]), .B(n14535), .Z(n14537) );
  XNOR U13905 ( .A(n14538), .B(n14539), .Z(n14535) );
  AND U13906 ( .A(n2146), .B(n14540), .Z(n14539) );
  XOR U13907 ( .A(n14541), .B(n14542), .Z(n14533) );
  AND U13908 ( .A(n2150), .B(n14543), .Z(n14542) );
  XOR U13909 ( .A(n14544), .B(n14545), .Z(n14530) );
  AND U13910 ( .A(n2154), .B(n14543), .Z(n14545) );
  XNOR U13911 ( .A(n14546), .B(n14544), .Z(n14543) );
  IV U13912 ( .A(n14541), .Z(n14546) );
  XOR U13913 ( .A(n14547), .B(n14548), .Z(n14541) );
  AND U13914 ( .A(n2157), .B(n14540), .Z(n14548) );
  XNOR U13915 ( .A(n14538), .B(n14547), .Z(n14540) );
  XNOR U13916 ( .A(n14549), .B(n14550), .Z(n14538) );
  AND U13917 ( .A(n2161), .B(n14551), .Z(n14550) );
  XOR U13918 ( .A(p_input[1762]), .B(n14549), .Z(n14551) );
  XNOR U13919 ( .A(n14552), .B(n14553), .Z(n14549) );
  AND U13920 ( .A(n2165), .B(n14554), .Z(n14553) );
  XOR U13921 ( .A(n14555), .B(n14556), .Z(n14547) );
  AND U13922 ( .A(n2169), .B(n14557), .Z(n14556) );
  XOR U13923 ( .A(n14558), .B(n14559), .Z(n14544) );
  AND U13924 ( .A(n2173), .B(n14557), .Z(n14559) );
  XNOR U13925 ( .A(n14560), .B(n14558), .Z(n14557) );
  IV U13926 ( .A(n14555), .Z(n14560) );
  XOR U13927 ( .A(n14561), .B(n14562), .Z(n14555) );
  AND U13928 ( .A(n2176), .B(n14554), .Z(n14562) );
  XNOR U13929 ( .A(n14552), .B(n14561), .Z(n14554) );
  XNOR U13930 ( .A(n14563), .B(n14564), .Z(n14552) );
  AND U13931 ( .A(n2180), .B(n14565), .Z(n14564) );
  XOR U13932 ( .A(p_input[1778]), .B(n14563), .Z(n14565) );
  XNOR U13933 ( .A(n14566), .B(n14567), .Z(n14563) );
  AND U13934 ( .A(n2184), .B(n14568), .Z(n14567) );
  XOR U13935 ( .A(n14569), .B(n14570), .Z(n14561) );
  AND U13936 ( .A(n2188), .B(n14571), .Z(n14570) );
  XOR U13937 ( .A(n14572), .B(n14573), .Z(n14558) );
  AND U13938 ( .A(n2192), .B(n14571), .Z(n14573) );
  XNOR U13939 ( .A(n14574), .B(n14572), .Z(n14571) );
  IV U13940 ( .A(n14569), .Z(n14574) );
  XOR U13941 ( .A(n14575), .B(n14576), .Z(n14569) );
  AND U13942 ( .A(n2195), .B(n14568), .Z(n14576) );
  XNOR U13943 ( .A(n14566), .B(n14575), .Z(n14568) );
  XNOR U13944 ( .A(n14577), .B(n14578), .Z(n14566) );
  AND U13945 ( .A(n2199), .B(n14579), .Z(n14578) );
  XOR U13946 ( .A(p_input[1794]), .B(n14577), .Z(n14579) );
  XNOR U13947 ( .A(n14580), .B(n14581), .Z(n14577) );
  AND U13948 ( .A(n2203), .B(n14582), .Z(n14581) );
  XOR U13949 ( .A(n14583), .B(n14584), .Z(n14575) );
  AND U13950 ( .A(n2207), .B(n14585), .Z(n14584) );
  XOR U13951 ( .A(n14586), .B(n14587), .Z(n14572) );
  AND U13952 ( .A(n2211), .B(n14585), .Z(n14587) );
  XNOR U13953 ( .A(n14588), .B(n14586), .Z(n14585) );
  IV U13954 ( .A(n14583), .Z(n14588) );
  XOR U13955 ( .A(n14589), .B(n14590), .Z(n14583) );
  AND U13956 ( .A(n2214), .B(n14582), .Z(n14590) );
  XNOR U13957 ( .A(n14580), .B(n14589), .Z(n14582) );
  XNOR U13958 ( .A(n14591), .B(n14592), .Z(n14580) );
  AND U13959 ( .A(n2218), .B(n14593), .Z(n14592) );
  XOR U13960 ( .A(p_input[1810]), .B(n14591), .Z(n14593) );
  XNOR U13961 ( .A(n14594), .B(n14595), .Z(n14591) );
  AND U13962 ( .A(n2222), .B(n14596), .Z(n14595) );
  XOR U13963 ( .A(n14597), .B(n14598), .Z(n14589) );
  AND U13964 ( .A(n2226), .B(n14599), .Z(n14598) );
  XOR U13965 ( .A(n14600), .B(n14601), .Z(n14586) );
  AND U13966 ( .A(n2230), .B(n14599), .Z(n14601) );
  XNOR U13967 ( .A(n14602), .B(n14600), .Z(n14599) );
  IV U13968 ( .A(n14597), .Z(n14602) );
  XOR U13969 ( .A(n14603), .B(n14604), .Z(n14597) );
  AND U13970 ( .A(n2233), .B(n14596), .Z(n14604) );
  XNOR U13971 ( .A(n14594), .B(n14603), .Z(n14596) );
  XNOR U13972 ( .A(n14605), .B(n14606), .Z(n14594) );
  AND U13973 ( .A(n2237), .B(n14607), .Z(n14606) );
  XOR U13974 ( .A(p_input[1826]), .B(n14605), .Z(n14607) );
  XNOR U13975 ( .A(n14608), .B(n14609), .Z(n14605) );
  AND U13976 ( .A(n2241), .B(n14610), .Z(n14609) );
  XOR U13977 ( .A(n14611), .B(n14612), .Z(n14603) );
  AND U13978 ( .A(n2245), .B(n14613), .Z(n14612) );
  XOR U13979 ( .A(n14614), .B(n14615), .Z(n14600) );
  AND U13980 ( .A(n2249), .B(n14613), .Z(n14615) );
  XNOR U13981 ( .A(n14616), .B(n14614), .Z(n14613) );
  IV U13982 ( .A(n14611), .Z(n14616) );
  XOR U13983 ( .A(n14617), .B(n14618), .Z(n14611) );
  AND U13984 ( .A(n2252), .B(n14610), .Z(n14618) );
  XNOR U13985 ( .A(n14608), .B(n14617), .Z(n14610) );
  XNOR U13986 ( .A(n14619), .B(n14620), .Z(n14608) );
  AND U13987 ( .A(n2256), .B(n14621), .Z(n14620) );
  XOR U13988 ( .A(p_input[1842]), .B(n14619), .Z(n14621) );
  XNOR U13989 ( .A(n14622), .B(n14623), .Z(n14619) );
  AND U13990 ( .A(n2260), .B(n14624), .Z(n14623) );
  XOR U13991 ( .A(n14625), .B(n14626), .Z(n14617) );
  AND U13992 ( .A(n2264), .B(n14627), .Z(n14626) );
  XOR U13993 ( .A(n14628), .B(n14629), .Z(n14614) );
  AND U13994 ( .A(n2268), .B(n14627), .Z(n14629) );
  XNOR U13995 ( .A(n14630), .B(n14628), .Z(n14627) );
  IV U13996 ( .A(n14625), .Z(n14630) );
  XOR U13997 ( .A(n14631), .B(n14632), .Z(n14625) );
  AND U13998 ( .A(n2271), .B(n14624), .Z(n14632) );
  XNOR U13999 ( .A(n14622), .B(n14631), .Z(n14624) );
  XNOR U14000 ( .A(n14633), .B(n14634), .Z(n14622) );
  AND U14001 ( .A(n2275), .B(n14635), .Z(n14634) );
  XOR U14002 ( .A(p_input[1858]), .B(n14633), .Z(n14635) );
  XNOR U14003 ( .A(n14636), .B(n14637), .Z(n14633) );
  AND U14004 ( .A(n2279), .B(n14638), .Z(n14637) );
  XOR U14005 ( .A(n14639), .B(n14640), .Z(n14631) );
  AND U14006 ( .A(n2283), .B(n14641), .Z(n14640) );
  XOR U14007 ( .A(n14642), .B(n14643), .Z(n14628) );
  AND U14008 ( .A(n2287), .B(n14641), .Z(n14643) );
  XNOR U14009 ( .A(n14644), .B(n14642), .Z(n14641) );
  IV U14010 ( .A(n14639), .Z(n14644) );
  XOR U14011 ( .A(n14645), .B(n14646), .Z(n14639) );
  AND U14012 ( .A(n2290), .B(n14638), .Z(n14646) );
  XNOR U14013 ( .A(n14636), .B(n14645), .Z(n14638) );
  XNOR U14014 ( .A(n14647), .B(n14648), .Z(n14636) );
  AND U14015 ( .A(n2294), .B(n14649), .Z(n14648) );
  XOR U14016 ( .A(p_input[1874]), .B(n14647), .Z(n14649) );
  XNOR U14017 ( .A(n14650), .B(n14651), .Z(n14647) );
  AND U14018 ( .A(n2298), .B(n14652), .Z(n14651) );
  XOR U14019 ( .A(n14653), .B(n14654), .Z(n14645) );
  AND U14020 ( .A(n2302), .B(n14655), .Z(n14654) );
  XOR U14021 ( .A(n14656), .B(n14657), .Z(n14642) );
  AND U14022 ( .A(n2306), .B(n14655), .Z(n14657) );
  XNOR U14023 ( .A(n14658), .B(n14656), .Z(n14655) );
  IV U14024 ( .A(n14653), .Z(n14658) );
  XOR U14025 ( .A(n14659), .B(n14660), .Z(n14653) );
  AND U14026 ( .A(n2309), .B(n14652), .Z(n14660) );
  XNOR U14027 ( .A(n14650), .B(n14659), .Z(n14652) );
  XNOR U14028 ( .A(n14661), .B(n14662), .Z(n14650) );
  AND U14029 ( .A(n2313), .B(n14663), .Z(n14662) );
  XOR U14030 ( .A(p_input[1890]), .B(n14661), .Z(n14663) );
  XNOR U14031 ( .A(n14664), .B(n14665), .Z(n14661) );
  AND U14032 ( .A(n2317), .B(n14666), .Z(n14665) );
  XOR U14033 ( .A(n14667), .B(n14668), .Z(n14659) );
  AND U14034 ( .A(n2321), .B(n14669), .Z(n14668) );
  XOR U14035 ( .A(n14670), .B(n14671), .Z(n14656) );
  AND U14036 ( .A(n2325), .B(n14669), .Z(n14671) );
  XNOR U14037 ( .A(n14672), .B(n14670), .Z(n14669) );
  IV U14038 ( .A(n14667), .Z(n14672) );
  XOR U14039 ( .A(n14673), .B(n14674), .Z(n14667) );
  AND U14040 ( .A(n2328), .B(n14666), .Z(n14674) );
  XNOR U14041 ( .A(n14664), .B(n14673), .Z(n14666) );
  XNOR U14042 ( .A(n14675), .B(n14676), .Z(n14664) );
  AND U14043 ( .A(n2332), .B(n14677), .Z(n14676) );
  XOR U14044 ( .A(p_input[1906]), .B(n14675), .Z(n14677) );
  XNOR U14045 ( .A(n14678), .B(n14679), .Z(n14675) );
  AND U14046 ( .A(n2336), .B(n14680), .Z(n14679) );
  XOR U14047 ( .A(n14681), .B(n14682), .Z(n14673) );
  AND U14048 ( .A(n2340), .B(n14683), .Z(n14682) );
  XOR U14049 ( .A(n14684), .B(n14685), .Z(n14670) );
  AND U14050 ( .A(n2344), .B(n14683), .Z(n14685) );
  XNOR U14051 ( .A(n14686), .B(n14684), .Z(n14683) );
  IV U14052 ( .A(n14681), .Z(n14686) );
  XOR U14053 ( .A(n14687), .B(n14688), .Z(n14681) );
  AND U14054 ( .A(n2347), .B(n14680), .Z(n14688) );
  XNOR U14055 ( .A(n14678), .B(n14687), .Z(n14680) );
  XNOR U14056 ( .A(n14689), .B(n14690), .Z(n14678) );
  AND U14057 ( .A(n2351), .B(n14691), .Z(n14690) );
  XOR U14058 ( .A(p_input[1922]), .B(n14689), .Z(n14691) );
  XNOR U14059 ( .A(n14692), .B(n14693), .Z(n14689) );
  AND U14060 ( .A(n2355), .B(n14694), .Z(n14693) );
  XOR U14061 ( .A(n14695), .B(n14696), .Z(n14687) );
  AND U14062 ( .A(n2359), .B(n14697), .Z(n14696) );
  XOR U14063 ( .A(n14698), .B(n14699), .Z(n14684) );
  AND U14064 ( .A(n2363), .B(n14697), .Z(n14699) );
  XNOR U14065 ( .A(n14700), .B(n14698), .Z(n14697) );
  IV U14066 ( .A(n14695), .Z(n14700) );
  XOR U14067 ( .A(n14701), .B(n14702), .Z(n14695) );
  AND U14068 ( .A(n2366), .B(n14694), .Z(n14702) );
  XNOR U14069 ( .A(n14692), .B(n14701), .Z(n14694) );
  XNOR U14070 ( .A(n14703), .B(n14704), .Z(n14692) );
  AND U14071 ( .A(n2370), .B(n14705), .Z(n14704) );
  XOR U14072 ( .A(p_input[1938]), .B(n14703), .Z(n14705) );
  XNOR U14073 ( .A(n14706), .B(n14707), .Z(n14703) );
  AND U14074 ( .A(n2374), .B(n14708), .Z(n14707) );
  XOR U14075 ( .A(n14709), .B(n14710), .Z(n14701) );
  AND U14076 ( .A(n2378), .B(n14711), .Z(n14710) );
  XOR U14077 ( .A(n14712), .B(n14713), .Z(n14698) );
  AND U14078 ( .A(n2382), .B(n14711), .Z(n14713) );
  XNOR U14079 ( .A(n14714), .B(n14712), .Z(n14711) );
  IV U14080 ( .A(n14709), .Z(n14714) );
  XOR U14081 ( .A(n14715), .B(n14716), .Z(n14709) );
  AND U14082 ( .A(n2385), .B(n14708), .Z(n14716) );
  XNOR U14083 ( .A(n14706), .B(n14715), .Z(n14708) );
  XNOR U14084 ( .A(n14717), .B(n14718), .Z(n14706) );
  AND U14085 ( .A(n2389), .B(n14719), .Z(n14718) );
  XOR U14086 ( .A(p_input[1954]), .B(n14717), .Z(n14719) );
  XNOR U14087 ( .A(n14720), .B(n14721), .Z(n14717) );
  AND U14088 ( .A(n2393), .B(n14722), .Z(n14721) );
  XOR U14089 ( .A(n14723), .B(n14724), .Z(n14715) );
  AND U14090 ( .A(n2397), .B(n14725), .Z(n14724) );
  XOR U14091 ( .A(n14726), .B(n14727), .Z(n14712) );
  AND U14092 ( .A(n2401), .B(n14725), .Z(n14727) );
  XNOR U14093 ( .A(n14728), .B(n14726), .Z(n14725) );
  IV U14094 ( .A(n14723), .Z(n14728) );
  XOR U14095 ( .A(n14729), .B(n14730), .Z(n14723) );
  AND U14096 ( .A(n2404), .B(n14722), .Z(n14730) );
  XNOR U14097 ( .A(n14720), .B(n14729), .Z(n14722) );
  XNOR U14098 ( .A(n14731), .B(n14732), .Z(n14720) );
  AND U14099 ( .A(n2408), .B(n14733), .Z(n14732) );
  XOR U14100 ( .A(p_input[1970]), .B(n14731), .Z(n14733) );
  XNOR U14101 ( .A(n14734), .B(n14735), .Z(n14731) );
  AND U14102 ( .A(n2412), .B(n14736), .Z(n14735) );
  XOR U14103 ( .A(n14737), .B(n14738), .Z(n14729) );
  AND U14104 ( .A(n2416), .B(n14739), .Z(n14738) );
  XOR U14105 ( .A(n14740), .B(n14741), .Z(n14726) );
  AND U14106 ( .A(n2420), .B(n14739), .Z(n14741) );
  XNOR U14107 ( .A(n14742), .B(n14740), .Z(n14739) );
  IV U14108 ( .A(n14737), .Z(n14742) );
  XOR U14109 ( .A(n14743), .B(n14744), .Z(n14737) );
  AND U14110 ( .A(n2423), .B(n14736), .Z(n14744) );
  XNOR U14111 ( .A(n14734), .B(n14743), .Z(n14736) );
  XNOR U14112 ( .A(n14745), .B(n14746), .Z(n14734) );
  AND U14113 ( .A(n2427), .B(n14747), .Z(n14746) );
  XOR U14114 ( .A(p_input[1986]), .B(n14745), .Z(n14747) );
  XOR U14115 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n14748), 
        .Z(n14745) );
  AND U14116 ( .A(n2430), .B(n14749), .Z(n14748) );
  XOR U14117 ( .A(n14750), .B(n14751), .Z(n14743) );
  AND U14118 ( .A(n2434), .B(n14752), .Z(n14751) );
  XOR U14119 ( .A(n14753), .B(n14754), .Z(n14740) );
  AND U14120 ( .A(n2438), .B(n14752), .Z(n14754) );
  XNOR U14121 ( .A(n14755), .B(n14753), .Z(n14752) );
  IV U14122 ( .A(n14750), .Z(n14755) );
  XOR U14123 ( .A(n14756), .B(n14757), .Z(n14750) );
  AND U14124 ( .A(n2441), .B(n14749), .Z(n14757) );
  XOR U14125 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n14756), 
        .Z(n14749) );
  XOR U14126 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n14758), 
        .Z(n14756) );
  AND U14127 ( .A(n2443), .B(n14759), .Z(n14758) );
  XOR U14128 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n14760), .Z(n14753) );
  AND U14129 ( .A(n2446), .B(n14759), .Z(n14760) );
  XOR U14130 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n14759) );
  XOR U14131 ( .A(n11244), .B(n14761), .Z(o[17]) );
  AND U14132 ( .A(n62), .B(n14762), .Z(n11244) );
  XOR U14133 ( .A(n11245), .B(n14761), .Z(n14762) );
  XOR U14134 ( .A(n14763), .B(n43), .Z(n14761) );
  AND U14135 ( .A(n65), .B(n14764), .Z(n43) );
  XOR U14136 ( .A(n44), .B(n14763), .Z(n14764) );
  XOR U14137 ( .A(n14765), .B(n14766), .Z(n44) );
  AND U14138 ( .A(n70), .B(n14767), .Z(n14766) );
  XOR U14139 ( .A(p_input[1]), .B(n14765), .Z(n14767) );
  XNOR U14140 ( .A(n14768), .B(n14769), .Z(n14765) );
  AND U14141 ( .A(n74), .B(n14770), .Z(n14769) );
  XOR U14142 ( .A(n14771), .B(n14772), .Z(n14763) );
  AND U14143 ( .A(n78), .B(n14773), .Z(n14772) );
  XOR U14144 ( .A(n14774), .B(n14775), .Z(n11245) );
  AND U14145 ( .A(n82), .B(n14773), .Z(n14775) );
  XNOR U14146 ( .A(n14776), .B(n14774), .Z(n14773) );
  IV U14147 ( .A(n14771), .Z(n14776) );
  XOR U14148 ( .A(n14777), .B(n14778), .Z(n14771) );
  AND U14149 ( .A(n86), .B(n14770), .Z(n14778) );
  XNOR U14150 ( .A(n14768), .B(n14777), .Z(n14770) );
  XNOR U14151 ( .A(n14779), .B(n14780), .Z(n14768) );
  AND U14152 ( .A(n90), .B(n14781), .Z(n14780) );
  XOR U14153 ( .A(p_input[17]), .B(n14779), .Z(n14781) );
  XNOR U14154 ( .A(n14782), .B(n14783), .Z(n14779) );
  AND U14155 ( .A(n94), .B(n14784), .Z(n14783) );
  XOR U14156 ( .A(n14785), .B(n14786), .Z(n14777) );
  AND U14157 ( .A(n98), .B(n14787), .Z(n14786) );
  XOR U14158 ( .A(n14788), .B(n14789), .Z(n14774) );
  AND U14159 ( .A(n102), .B(n14787), .Z(n14789) );
  XNOR U14160 ( .A(n14790), .B(n14788), .Z(n14787) );
  IV U14161 ( .A(n14785), .Z(n14790) );
  XOR U14162 ( .A(n14791), .B(n14792), .Z(n14785) );
  AND U14163 ( .A(n105), .B(n14784), .Z(n14792) );
  XNOR U14164 ( .A(n14782), .B(n14791), .Z(n14784) );
  XNOR U14165 ( .A(n14793), .B(n14794), .Z(n14782) );
  AND U14166 ( .A(n109), .B(n14795), .Z(n14794) );
  XOR U14167 ( .A(p_input[33]), .B(n14793), .Z(n14795) );
  XNOR U14168 ( .A(n14796), .B(n14797), .Z(n14793) );
  AND U14169 ( .A(n113), .B(n14798), .Z(n14797) );
  XOR U14170 ( .A(n14799), .B(n14800), .Z(n14791) );
  AND U14171 ( .A(n117), .B(n14801), .Z(n14800) );
  XOR U14172 ( .A(n14802), .B(n14803), .Z(n14788) );
  AND U14173 ( .A(n121), .B(n14801), .Z(n14803) );
  XNOR U14174 ( .A(n14804), .B(n14802), .Z(n14801) );
  IV U14175 ( .A(n14799), .Z(n14804) );
  XOR U14176 ( .A(n14805), .B(n14806), .Z(n14799) );
  AND U14177 ( .A(n124), .B(n14798), .Z(n14806) );
  XNOR U14178 ( .A(n14796), .B(n14805), .Z(n14798) );
  XNOR U14179 ( .A(n14807), .B(n14808), .Z(n14796) );
  AND U14180 ( .A(n128), .B(n14809), .Z(n14808) );
  XOR U14181 ( .A(p_input[49]), .B(n14807), .Z(n14809) );
  XNOR U14182 ( .A(n14810), .B(n14811), .Z(n14807) );
  AND U14183 ( .A(n132), .B(n14812), .Z(n14811) );
  XOR U14184 ( .A(n14813), .B(n14814), .Z(n14805) );
  AND U14185 ( .A(n136), .B(n14815), .Z(n14814) );
  XOR U14186 ( .A(n14816), .B(n14817), .Z(n14802) );
  AND U14187 ( .A(n140), .B(n14815), .Z(n14817) );
  XNOR U14188 ( .A(n14818), .B(n14816), .Z(n14815) );
  IV U14189 ( .A(n14813), .Z(n14818) );
  XOR U14190 ( .A(n14819), .B(n14820), .Z(n14813) );
  AND U14191 ( .A(n143), .B(n14812), .Z(n14820) );
  XNOR U14192 ( .A(n14810), .B(n14819), .Z(n14812) );
  XNOR U14193 ( .A(n14821), .B(n14822), .Z(n14810) );
  AND U14194 ( .A(n147), .B(n14823), .Z(n14822) );
  XOR U14195 ( .A(p_input[65]), .B(n14821), .Z(n14823) );
  XNOR U14196 ( .A(n14824), .B(n14825), .Z(n14821) );
  AND U14197 ( .A(n151), .B(n14826), .Z(n14825) );
  XOR U14198 ( .A(n14827), .B(n14828), .Z(n14819) );
  AND U14199 ( .A(n155), .B(n14829), .Z(n14828) );
  XOR U14200 ( .A(n14830), .B(n14831), .Z(n14816) );
  AND U14201 ( .A(n159), .B(n14829), .Z(n14831) );
  XNOR U14202 ( .A(n14832), .B(n14830), .Z(n14829) );
  IV U14203 ( .A(n14827), .Z(n14832) );
  XOR U14204 ( .A(n14833), .B(n14834), .Z(n14827) );
  AND U14205 ( .A(n162), .B(n14826), .Z(n14834) );
  XNOR U14206 ( .A(n14824), .B(n14833), .Z(n14826) );
  XNOR U14207 ( .A(n14835), .B(n14836), .Z(n14824) );
  AND U14208 ( .A(n166), .B(n14837), .Z(n14836) );
  XOR U14209 ( .A(p_input[81]), .B(n14835), .Z(n14837) );
  XNOR U14210 ( .A(n14838), .B(n14839), .Z(n14835) );
  AND U14211 ( .A(n170), .B(n14840), .Z(n14839) );
  XOR U14212 ( .A(n14841), .B(n14842), .Z(n14833) );
  AND U14213 ( .A(n174), .B(n14843), .Z(n14842) );
  XOR U14214 ( .A(n14844), .B(n14845), .Z(n14830) );
  AND U14215 ( .A(n178), .B(n14843), .Z(n14845) );
  XNOR U14216 ( .A(n14846), .B(n14844), .Z(n14843) );
  IV U14217 ( .A(n14841), .Z(n14846) );
  XOR U14218 ( .A(n14847), .B(n14848), .Z(n14841) );
  AND U14219 ( .A(n181), .B(n14840), .Z(n14848) );
  XNOR U14220 ( .A(n14838), .B(n14847), .Z(n14840) );
  XNOR U14221 ( .A(n14849), .B(n14850), .Z(n14838) );
  AND U14222 ( .A(n185), .B(n14851), .Z(n14850) );
  XOR U14223 ( .A(p_input[97]), .B(n14849), .Z(n14851) );
  XNOR U14224 ( .A(n14852), .B(n14853), .Z(n14849) );
  AND U14225 ( .A(n189), .B(n14854), .Z(n14853) );
  XOR U14226 ( .A(n14855), .B(n14856), .Z(n14847) );
  AND U14227 ( .A(n193), .B(n14857), .Z(n14856) );
  XOR U14228 ( .A(n14858), .B(n14859), .Z(n14844) );
  AND U14229 ( .A(n197), .B(n14857), .Z(n14859) );
  XNOR U14230 ( .A(n14860), .B(n14858), .Z(n14857) );
  IV U14231 ( .A(n14855), .Z(n14860) );
  XOR U14232 ( .A(n14861), .B(n14862), .Z(n14855) );
  AND U14233 ( .A(n200), .B(n14854), .Z(n14862) );
  XNOR U14234 ( .A(n14852), .B(n14861), .Z(n14854) );
  XNOR U14235 ( .A(n14863), .B(n14864), .Z(n14852) );
  AND U14236 ( .A(n204), .B(n14865), .Z(n14864) );
  XOR U14237 ( .A(p_input[113]), .B(n14863), .Z(n14865) );
  XNOR U14238 ( .A(n14866), .B(n14867), .Z(n14863) );
  AND U14239 ( .A(n208), .B(n14868), .Z(n14867) );
  XOR U14240 ( .A(n14869), .B(n14870), .Z(n14861) );
  AND U14241 ( .A(n212), .B(n14871), .Z(n14870) );
  XOR U14242 ( .A(n14872), .B(n14873), .Z(n14858) );
  AND U14243 ( .A(n216), .B(n14871), .Z(n14873) );
  XNOR U14244 ( .A(n14874), .B(n14872), .Z(n14871) );
  IV U14245 ( .A(n14869), .Z(n14874) );
  XOR U14246 ( .A(n14875), .B(n14876), .Z(n14869) );
  AND U14247 ( .A(n219), .B(n14868), .Z(n14876) );
  XNOR U14248 ( .A(n14866), .B(n14875), .Z(n14868) );
  XNOR U14249 ( .A(n14877), .B(n14878), .Z(n14866) );
  AND U14250 ( .A(n223), .B(n14879), .Z(n14878) );
  XOR U14251 ( .A(p_input[129]), .B(n14877), .Z(n14879) );
  XNOR U14252 ( .A(n14880), .B(n14881), .Z(n14877) );
  AND U14253 ( .A(n227), .B(n14882), .Z(n14881) );
  XOR U14254 ( .A(n14883), .B(n14884), .Z(n14875) );
  AND U14255 ( .A(n231), .B(n14885), .Z(n14884) );
  XOR U14256 ( .A(n14886), .B(n14887), .Z(n14872) );
  AND U14257 ( .A(n235), .B(n14885), .Z(n14887) );
  XNOR U14258 ( .A(n14888), .B(n14886), .Z(n14885) );
  IV U14259 ( .A(n14883), .Z(n14888) );
  XOR U14260 ( .A(n14889), .B(n14890), .Z(n14883) );
  AND U14261 ( .A(n238), .B(n14882), .Z(n14890) );
  XNOR U14262 ( .A(n14880), .B(n14889), .Z(n14882) );
  XNOR U14263 ( .A(n14891), .B(n14892), .Z(n14880) );
  AND U14264 ( .A(n242), .B(n14893), .Z(n14892) );
  XOR U14265 ( .A(p_input[145]), .B(n14891), .Z(n14893) );
  XNOR U14266 ( .A(n14894), .B(n14895), .Z(n14891) );
  AND U14267 ( .A(n246), .B(n14896), .Z(n14895) );
  XOR U14268 ( .A(n14897), .B(n14898), .Z(n14889) );
  AND U14269 ( .A(n250), .B(n14899), .Z(n14898) );
  XOR U14270 ( .A(n14900), .B(n14901), .Z(n14886) );
  AND U14271 ( .A(n254), .B(n14899), .Z(n14901) );
  XNOR U14272 ( .A(n14902), .B(n14900), .Z(n14899) );
  IV U14273 ( .A(n14897), .Z(n14902) );
  XOR U14274 ( .A(n14903), .B(n14904), .Z(n14897) );
  AND U14275 ( .A(n257), .B(n14896), .Z(n14904) );
  XNOR U14276 ( .A(n14894), .B(n14903), .Z(n14896) );
  XNOR U14277 ( .A(n14905), .B(n14906), .Z(n14894) );
  AND U14278 ( .A(n261), .B(n14907), .Z(n14906) );
  XOR U14279 ( .A(p_input[161]), .B(n14905), .Z(n14907) );
  XNOR U14280 ( .A(n14908), .B(n14909), .Z(n14905) );
  AND U14281 ( .A(n265), .B(n14910), .Z(n14909) );
  XOR U14282 ( .A(n14911), .B(n14912), .Z(n14903) );
  AND U14283 ( .A(n269), .B(n14913), .Z(n14912) );
  XOR U14284 ( .A(n14914), .B(n14915), .Z(n14900) );
  AND U14285 ( .A(n273), .B(n14913), .Z(n14915) );
  XNOR U14286 ( .A(n14916), .B(n14914), .Z(n14913) );
  IV U14287 ( .A(n14911), .Z(n14916) );
  XOR U14288 ( .A(n14917), .B(n14918), .Z(n14911) );
  AND U14289 ( .A(n276), .B(n14910), .Z(n14918) );
  XNOR U14290 ( .A(n14908), .B(n14917), .Z(n14910) );
  XNOR U14291 ( .A(n14919), .B(n14920), .Z(n14908) );
  AND U14292 ( .A(n280), .B(n14921), .Z(n14920) );
  XOR U14293 ( .A(p_input[177]), .B(n14919), .Z(n14921) );
  XNOR U14294 ( .A(n14922), .B(n14923), .Z(n14919) );
  AND U14295 ( .A(n284), .B(n14924), .Z(n14923) );
  XOR U14296 ( .A(n14925), .B(n14926), .Z(n14917) );
  AND U14297 ( .A(n288), .B(n14927), .Z(n14926) );
  XOR U14298 ( .A(n14928), .B(n14929), .Z(n14914) );
  AND U14299 ( .A(n292), .B(n14927), .Z(n14929) );
  XNOR U14300 ( .A(n14930), .B(n14928), .Z(n14927) );
  IV U14301 ( .A(n14925), .Z(n14930) );
  XOR U14302 ( .A(n14931), .B(n14932), .Z(n14925) );
  AND U14303 ( .A(n295), .B(n14924), .Z(n14932) );
  XNOR U14304 ( .A(n14922), .B(n14931), .Z(n14924) );
  XNOR U14305 ( .A(n14933), .B(n14934), .Z(n14922) );
  AND U14306 ( .A(n299), .B(n14935), .Z(n14934) );
  XOR U14307 ( .A(p_input[193]), .B(n14933), .Z(n14935) );
  XNOR U14308 ( .A(n14936), .B(n14937), .Z(n14933) );
  AND U14309 ( .A(n303), .B(n14938), .Z(n14937) );
  XOR U14310 ( .A(n14939), .B(n14940), .Z(n14931) );
  AND U14311 ( .A(n307), .B(n14941), .Z(n14940) );
  XOR U14312 ( .A(n14942), .B(n14943), .Z(n14928) );
  AND U14313 ( .A(n311), .B(n14941), .Z(n14943) );
  XNOR U14314 ( .A(n14944), .B(n14942), .Z(n14941) );
  IV U14315 ( .A(n14939), .Z(n14944) );
  XOR U14316 ( .A(n14945), .B(n14946), .Z(n14939) );
  AND U14317 ( .A(n314), .B(n14938), .Z(n14946) );
  XNOR U14318 ( .A(n14936), .B(n14945), .Z(n14938) );
  XNOR U14319 ( .A(n14947), .B(n14948), .Z(n14936) );
  AND U14320 ( .A(n318), .B(n14949), .Z(n14948) );
  XOR U14321 ( .A(p_input[209]), .B(n14947), .Z(n14949) );
  XNOR U14322 ( .A(n14950), .B(n14951), .Z(n14947) );
  AND U14323 ( .A(n322), .B(n14952), .Z(n14951) );
  XOR U14324 ( .A(n14953), .B(n14954), .Z(n14945) );
  AND U14325 ( .A(n326), .B(n14955), .Z(n14954) );
  XOR U14326 ( .A(n14956), .B(n14957), .Z(n14942) );
  AND U14327 ( .A(n330), .B(n14955), .Z(n14957) );
  XNOR U14328 ( .A(n14958), .B(n14956), .Z(n14955) );
  IV U14329 ( .A(n14953), .Z(n14958) );
  XOR U14330 ( .A(n14959), .B(n14960), .Z(n14953) );
  AND U14331 ( .A(n333), .B(n14952), .Z(n14960) );
  XNOR U14332 ( .A(n14950), .B(n14959), .Z(n14952) );
  XNOR U14333 ( .A(n14961), .B(n14962), .Z(n14950) );
  AND U14334 ( .A(n337), .B(n14963), .Z(n14962) );
  XOR U14335 ( .A(p_input[225]), .B(n14961), .Z(n14963) );
  XNOR U14336 ( .A(n14964), .B(n14965), .Z(n14961) );
  AND U14337 ( .A(n341), .B(n14966), .Z(n14965) );
  XOR U14338 ( .A(n14967), .B(n14968), .Z(n14959) );
  AND U14339 ( .A(n345), .B(n14969), .Z(n14968) );
  XOR U14340 ( .A(n14970), .B(n14971), .Z(n14956) );
  AND U14341 ( .A(n349), .B(n14969), .Z(n14971) );
  XNOR U14342 ( .A(n14972), .B(n14970), .Z(n14969) );
  IV U14343 ( .A(n14967), .Z(n14972) );
  XOR U14344 ( .A(n14973), .B(n14974), .Z(n14967) );
  AND U14345 ( .A(n352), .B(n14966), .Z(n14974) );
  XNOR U14346 ( .A(n14964), .B(n14973), .Z(n14966) );
  XNOR U14347 ( .A(n14975), .B(n14976), .Z(n14964) );
  AND U14348 ( .A(n356), .B(n14977), .Z(n14976) );
  XOR U14349 ( .A(p_input[241]), .B(n14975), .Z(n14977) );
  XNOR U14350 ( .A(n14978), .B(n14979), .Z(n14975) );
  AND U14351 ( .A(n360), .B(n14980), .Z(n14979) );
  XOR U14352 ( .A(n14981), .B(n14982), .Z(n14973) );
  AND U14353 ( .A(n364), .B(n14983), .Z(n14982) );
  XOR U14354 ( .A(n14984), .B(n14985), .Z(n14970) );
  AND U14355 ( .A(n368), .B(n14983), .Z(n14985) );
  XNOR U14356 ( .A(n14986), .B(n14984), .Z(n14983) );
  IV U14357 ( .A(n14981), .Z(n14986) );
  XOR U14358 ( .A(n14987), .B(n14988), .Z(n14981) );
  AND U14359 ( .A(n371), .B(n14980), .Z(n14988) );
  XNOR U14360 ( .A(n14978), .B(n14987), .Z(n14980) );
  XNOR U14361 ( .A(n14989), .B(n14990), .Z(n14978) );
  AND U14362 ( .A(n375), .B(n14991), .Z(n14990) );
  XOR U14363 ( .A(p_input[257]), .B(n14989), .Z(n14991) );
  XNOR U14364 ( .A(n14992), .B(n14993), .Z(n14989) );
  AND U14365 ( .A(n379), .B(n14994), .Z(n14993) );
  XOR U14366 ( .A(n14995), .B(n14996), .Z(n14987) );
  AND U14367 ( .A(n383), .B(n14997), .Z(n14996) );
  XOR U14368 ( .A(n14998), .B(n14999), .Z(n14984) );
  AND U14369 ( .A(n387), .B(n14997), .Z(n14999) );
  XNOR U14370 ( .A(n15000), .B(n14998), .Z(n14997) );
  IV U14371 ( .A(n14995), .Z(n15000) );
  XOR U14372 ( .A(n15001), .B(n15002), .Z(n14995) );
  AND U14373 ( .A(n390), .B(n14994), .Z(n15002) );
  XNOR U14374 ( .A(n14992), .B(n15001), .Z(n14994) );
  XNOR U14375 ( .A(n15003), .B(n15004), .Z(n14992) );
  AND U14376 ( .A(n394), .B(n15005), .Z(n15004) );
  XOR U14377 ( .A(p_input[273]), .B(n15003), .Z(n15005) );
  XNOR U14378 ( .A(n15006), .B(n15007), .Z(n15003) );
  AND U14379 ( .A(n398), .B(n15008), .Z(n15007) );
  XOR U14380 ( .A(n15009), .B(n15010), .Z(n15001) );
  AND U14381 ( .A(n402), .B(n15011), .Z(n15010) );
  XOR U14382 ( .A(n15012), .B(n15013), .Z(n14998) );
  AND U14383 ( .A(n406), .B(n15011), .Z(n15013) );
  XNOR U14384 ( .A(n15014), .B(n15012), .Z(n15011) );
  IV U14385 ( .A(n15009), .Z(n15014) );
  XOR U14386 ( .A(n15015), .B(n15016), .Z(n15009) );
  AND U14387 ( .A(n409), .B(n15008), .Z(n15016) );
  XNOR U14388 ( .A(n15006), .B(n15015), .Z(n15008) );
  XNOR U14389 ( .A(n15017), .B(n15018), .Z(n15006) );
  AND U14390 ( .A(n413), .B(n15019), .Z(n15018) );
  XOR U14391 ( .A(p_input[289]), .B(n15017), .Z(n15019) );
  XNOR U14392 ( .A(n15020), .B(n15021), .Z(n15017) );
  AND U14393 ( .A(n417), .B(n15022), .Z(n15021) );
  XOR U14394 ( .A(n15023), .B(n15024), .Z(n15015) );
  AND U14395 ( .A(n421), .B(n15025), .Z(n15024) );
  XOR U14396 ( .A(n15026), .B(n15027), .Z(n15012) );
  AND U14397 ( .A(n425), .B(n15025), .Z(n15027) );
  XNOR U14398 ( .A(n15028), .B(n15026), .Z(n15025) );
  IV U14399 ( .A(n15023), .Z(n15028) );
  XOR U14400 ( .A(n15029), .B(n15030), .Z(n15023) );
  AND U14401 ( .A(n428), .B(n15022), .Z(n15030) );
  XNOR U14402 ( .A(n15020), .B(n15029), .Z(n15022) );
  XNOR U14403 ( .A(n15031), .B(n15032), .Z(n15020) );
  AND U14404 ( .A(n432), .B(n15033), .Z(n15032) );
  XOR U14405 ( .A(p_input[305]), .B(n15031), .Z(n15033) );
  XNOR U14406 ( .A(n15034), .B(n15035), .Z(n15031) );
  AND U14407 ( .A(n436), .B(n15036), .Z(n15035) );
  XOR U14408 ( .A(n15037), .B(n15038), .Z(n15029) );
  AND U14409 ( .A(n440), .B(n15039), .Z(n15038) );
  XOR U14410 ( .A(n15040), .B(n15041), .Z(n15026) );
  AND U14411 ( .A(n444), .B(n15039), .Z(n15041) );
  XNOR U14412 ( .A(n15042), .B(n15040), .Z(n15039) );
  IV U14413 ( .A(n15037), .Z(n15042) );
  XOR U14414 ( .A(n15043), .B(n15044), .Z(n15037) );
  AND U14415 ( .A(n447), .B(n15036), .Z(n15044) );
  XNOR U14416 ( .A(n15034), .B(n15043), .Z(n15036) );
  XNOR U14417 ( .A(n15045), .B(n15046), .Z(n15034) );
  AND U14418 ( .A(n451), .B(n15047), .Z(n15046) );
  XOR U14419 ( .A(p_input[321]), .B(n15045), .Z(n15047) );
  XNOR U14420 ( .A(n15048), .B(n15049), .Z(n15045) );
  AND U14421 ( .A(n455), .B(n15050), .Z(n15049) );
  XOR U14422 ( .A(n15051), .B(n15052), .Z(n15043) );
  AND U14423 ( .A(n459), .B(n15053), .Z(n15052) );
  XOR U14424 ( .A(n15054), .B(n15055), .Z(n15040) );
  AND U14425 ( .A(n463), .B(n15053), .Z(n15055) );
  XNOR U14426 ( .A(n15056), .B(n15054), .Z(n15053) );
  IV U14427 ( .A(n15051), .Z(n15056) );
  XOR U14428 ( .A(n15057), .B(n15058), .Z(n15051) );
  AND U14429 ( .A(n466), .B(n15050), .Z(n15058) );
  XNOR U14430 ( .A(n15048), .B(n15057), .Z(n15050) );
  XNOR U14431 ( .A(n15059), .B(n15060), .Z(n15048) );
  AND U14432 ( .A(n470), .B(n15061), .Z(n15060) );
  XOR U14433 ( .A(p_input[337]), .B(n15059), .Z(n15061) );
  XNOR U14434 ( .A(n15062), .B(n15063), .Z(n15059) );
  AND U14435 ( .A(n474), .B(n15064), .Z(n15063) );
  XOR U14436 ( .A(n15065), .B(n15066), .Z(n15057) );
  AND U14437 ( .A(n478), .B(n15067), .Z(n15066) );
  XOR U14438 ( .A(n15068), .B(n15069), .Z(n15054) );
  AND U14439 ( .A(n482), .B(n15067), .Z(n15069) );
  XNOR U14440 ( .A(n15070), .B(n15068), .Z(n15067) );
  IV U14441 ( .A(n15065), .Z(n15070) );
  XOR U14442 ( .A(n15071), .B(n15072), .Z(n15065) );
  AND U14443 ( .A(n485), .B(n15064), .Z(n15072) );
  XNOR U14444 ( .A(n15062), .B(n15071), .Z(n15064) );
  XNOR U14445 ( .A(n15073), .B(n15074), .Z(n15062) );
  AND U14446 ( .A(n489), .B(n15075), .Z(n15074) );
  XOR U14447 ( .A(p_input[353]), .B(n15073), .Z(n15075) );
  XNOR U14448 ( .A(n15076), .B(n15077), .Z(n15073) );
  AND U14449 ( .A(n493), .B(n15078), .Z(n15077) );
  XOR U14450 ( .A(n15079), .B(n15080), .Z(n15071) );
  AND U14451 ( .A(n497), .B(n15081), .Z(n15080) );
  XOR U14452 ( .A(n15082), .B(n15083), .Z(n15068) );
  AND U14453 ( .A(n501), .B(n15081), .Z(n15083) );
  XNOR U14454 ( .A(n15084), .B(n15082), .Z(n15081) );
  IV U14455 ( .A(n15079), .Z(n15084) );
  XOR U14456 ( .A(n15085), .B(n15086), .Z(n15079) );
  AND U14457 ( .A(n504), .B(n15078), .Z(n15086) );
  XNOR U14458 ( .A(n15076), .B(n15085), .Z(n15078) );
  XNOR U14459 ( .A(n15087), .B(n15088), .Z(n15076) );
  AND U14460 ( .A(n508), .B(n15089), .Z(n15088) );
  XOR U14461 ( .A(p_input[369]), .B(n15087), .Z(n15089) );
  XNOR U14462 ( .A(n15090), .B(n15091), .Z(n15087) );
  AND U14463 ( .A(n512), .B(n15092), .Z(n15091) );
  XOR U14464 ( .A(n15093), .B(n15094), .Z(n15085) );
  AND U14465 ( .A(n516), .B(n15095), .Z(n15094) );
  XOR U14466 ( .A(n15096), .B(n15097), .Z(n15082) );
  AND U14467 ( .A(n520), .B(n15095), .Z(n15097) );
  XNOR U14468 ( .A(n15098), .B(n15096), .Z(n15095) );
  IV U14469 ( .A(n15093), .Z(n15098) );
  XOR U14470 ( .A(n15099), .B(n15100), .Z(n15093) );
  AND U14471 ( .A(n523), .B(n15092), .Z(n15100) );
  XNOR U14472 ( .A(n15090), .B(n15099), .Z(n15092) );
  XNOR U14473 ( .A(n15101), .B(n15102), .Z(n15090) );
  AND U14474 ( .A(n527), .B(n15103), .Z(n15102) );
  XOR U14475 ( .A(p_input[385]), .B(n15101), .Z(n15103) );
  XNOR U14476 ( .A(n15104), .B(n15105), .Z(n15101) );
  AND U14477 ( .A(n531), .B(n15106), .Z(n15105) );
  XOR U14478 ( .A(n15107), .B(n15108), .Z(n15099) );
  AND U14479 ( .A(n535), .B(n15109), .Z(n15108) );
  XOR U14480 ( .A(n15110), .B(n15111), .Z(n15096) );
  AND U14481 ( .A(n539), .B(n15109), .Z(n15111) );
  XNOR U14482 ( .A(n15112), .B(n15110), .Z(n15109) );
  IV U14483 ( .A(n15107), .Z(n15112) );
  XOR U14484 ( .A(n15113), .B(n15114), .Z(n15107) );
  AND U14485 ( .A(n542), .B(n15106), .Z(n15114) );
  XNOR U14486 ( .A(n15104), .B(n15113), .Z(n15106) );
  XNOR U14487 ( .A(n15115), .B(n15116), .Z(n15104) );
  AND U14488 ( .A(n546), .B(n15117), .Z(n15116) );
  XOR U14489 ( .A(p_input[401]), .B(n15115), .Z(n15117) );
  XNOR U14490 ( .A(n15118), .B(n15119), .Z(n15115) );
  AND U14491 ( .A(n550), .B(n15120), .Z(n15119) );
  XOR U14492 ( .A(n15121), .B(n15122), .Z(n15113) );
  AND U14493 ( .A(n554), .B(n15123), .Z(n15122) );
  XOR U14494 ( .A(n15124), .B(n15125), .Z(n15110) );
  AND U14495 ( .A(n558), .B(n15123), .Z(n15125) );
  XNOR U14496 ( .A(n15126), .B(n15124), .Z(n15123) );
  IV U14497 ( .A(n15121), .Z(n15126) );
  XOR U14498 ( .A(n15127), .B(n15128), .Z(n15121) );
  AND U14499 ( .A(n561), .B(n15120), .Z(n15128) );
  XNOR U14500 ( .A(n15118), .B(n15127), .Z(n15120) );
  XNOR U14501 ( .A(n15129), .B(n15130), .Z(n15118) );
  AND U14502 ( .A(n565), .B(n15131), .Z(n15130) );
  XOR U14503 ( .A(p_input[417]), .B(n15129), .Z(n15131) );
  XNOR U14504 ( .A(n15132), .B(n15133), .Z(n15129) );
  AND U14505 ( .A(n569), .B(n15134), .Z(n15133) );
  XOR U14506 ( .A(n15135), .B(n15136), .Z(n15127) );
  AND U14507 ( .A(n573), .B(n15137), .Z(n15136) );
  XOR U14508 ( .A(n15138), .B(n15139), .Z(n15124) );
  AND U14509 ( .A(n577), .B(n15137), .Z(n15139) );
  XNOR U14510 ( .A(n15140), .B(n15138), .Z(n15137) );
  IV U14511 ( .A(n15135), .Z(n15140) );
  XOR U14512 ( .A(n15141), .B(n15142), .Z(n15135) );
  AND U14513 ( .A(n580), .B(n15134), .Z(n15142) );
  XNOR U14514 ( .A(n15132), .B(n15141), .Z(n15134) );
  XNOR U14515 ( .A(n15143), .B(n15144), .Z(n15132) );
  AND U14516 ( .A(n584), .B(n15145), .Z(n15144) );
  XOR U14517 ( .A(p_input[433]), .B(n15143), .Z(n15145) );
  XNOR U14518 ( .A(n15146), .B(n15147), .Z(n15143) );
  AND U14519 ( .A(n588), .B(n15148), .Z(n15147) );
  XOR U14520 ( .A(n15149), .B(n15150), .Z(n15141) );
  AND U14521 ( .A(n592), .B(n15151), .Z(n15150) );
  XOR U14522 ( .A(n15152), .B(n15153), .Z(n15138) );
  AND U14523 ( .A(n596), .B(n15151), .Z(n15153) );
  XNOR U14524 ( .A(n15154), .B(n15152), .Z(n15151) );
  IV U14525 ( .A(n15149), .Z(n15154) );
  XOR U14526 ( .A(n15155), .B(n15156), .Z(n15149) );
  AND U14527 ( .A(n599), .B(n15148), .Z(n15156) );
  XNOR U14528 ( .A(n15146), .B(n15155), .Z(n15148) );
  XNOR U14529 ( .A(n15157), .B(n15158), .Z(n15146) );
  AND U14530 ( .A(n603), .B(n15159), .Z(n15158) );
  XOR U14531 ( .A(p_input[449]), .B(n15157), .Z(n15159) );
  XNOR U14532 ( .A(n15160), .B(n15161), .Z(n15157) );
  AND U14533 ( .A(n607), .B(n15162), .Z(n15161) );
  XOR U14534 ( .A(n15163), .B(n15164), .Z(n15155) );
  AND U14535 ( .A(n611), .B(n15165), .Z(n15164) );
  XOR U14536 ( .A(n15166), .B(n15167), .Z(n15152) );
  AND U14537 ( .A(n615), .B(n15165), .Z(n15167) );
  XNOR U14538 ( .A(n15168), .B(n15166), .Z(n15165) );
  IV U14539 ( .A(n15163), .Z(n15168) );
  XOR U14540 ( .A(n15169), .B(n15170), .Z(n15163) );
  AND U14541 ( .A(n618), .B(n15162), .Z(n15170) );
  XNOR U14542 ( .A(n15160), .B(n15169), .Z(n15162) );
  XNOR U14543 ( .A(n15171), .B(n15172), .Z(n15160) );
  AND U14544 ( .A(n622), .B(n15173), .Z(n15172) );
  XOR U14545 ( .A(p_input[465]), .B(n15171), .Z(n15173) );
  XNOR U14546 ( .A(n15174), .B(n15175), .Z(n15171) );
  AND U14547 ( .A(n626), .B(n15176), .Z(n15175) );
  XOR U14548 ( .A(n15177), .B(n15178), .Z(n15169) );
  AND U14549 ( .A(n630), .B(n15179), .Z(n15178) );
  XOR U14550 ( .A(n15180), .B(n15181), .Z(n15166) );
  AND U14551 ( .A(n634), .B(n15179), .Z(n15181) );
  XNOR U14552 ( .A(n15182), .B(n15180), .Z(n15179) );
  IV U14553 ( .A(n15177), .Z(n15182) );
  XOR U14554 ( .A(n15183), .B(n15184), .Z(n15177) );
  AND U14555 ( .A(n637), .B(n15176), .Z(n15184) );
  XNOR U14556 ( .A(n15174), .B(n15183), .Z(n15176) );
  XNOR U14557 ( .A(n15185), .B(n15186), .Z(n15174) );
  AND U14558 ( .A(n641), .B(n15187), .Z(n15186) );
  XOR U14559 ( .A(p_input[481]), .B(n15185), .Z(n15187) );
  XNOR U14560 ( .A(n15188), .B(n15189), .Z(n15185) );
  AND U14561 ( .A(n645), .B(n15190), .Z(n15189) );
  XOR U14562 ( .A(n15191), .B(n15192), .Z(n15183) );
  AND U14563 ( .A(n649), .B(n15193), .Z(n15192) );
  XOR U14564 ( .A(n15194), .B(n15195), .Z(n15180) );
  AND U14565 ( .A(n653), .B(n15193), .Z(n15195) );
  XNOR U14566 ( .A(n15196), .B(n15194), .Z(n15193) );
  IV U14567 ( .A(n15191), .Z(n15196) );
  XOR U14568 ( .A(n15197), .B(n15198), .Z(n15191) );
  AND U14569 ( .A(n656), .B(n15190), .Z(n15198) );
  XNOR U14570 ( .A(n15188), .B(n15197), .Z(n15190) );
  XNOR U14571 ( .A(n15199), .B(n15200), .Z(n15188) );
  AND U14572 ( .A(n660), .B(n15201), .Z(n15200) );
  XOR U14573 ( .A(p_input[497]), .B(n15199), .Z(n15201) );
  XNOR U14574 ( .A(n15202), .B(n15203), .Z(n15199) );
  AND U14575 ( .A(n664), .B(n15204), .Z(n15203) );
  XOR U14576 ( .A(n15205), .B(n15206), .Z(n15197) );
  AND U14577 ( .A(n668), .B(n15207), .Z(n15206) );
  XOR U14578 ( .A(n15208), .B(n15209), .Z(n15194) );
  AND U14579 ( .A(n672), .B(n15207), .Z(n15209) );
  XNOR U14580 ( .A(n15210), .B(n15208), .Z(n15207) );
  IV U14581 ( .A(n15205), .Z(n15210) );
  XOR U14582 ( .A(n15211), .B(n15212), .Z(n15205) );
  AND U14583 ( .A(n675), .B(n15204), .Z(n15212) );
  XNOR U14584 ( .A(n15202), .B(n15211), .Z(n15204) );
  XNOR U14585 ( .A(n15213), .B(n15214), .Z(n15202) );
  AND U14586 ( .A(n679), .B(n15215), .Z(n15214) );
  XOR U14587 ( .A(p_input[513]), .B(n15213), .Z(n15215) );
  XNOR U14588 ( .A(n15216), .B(n15217), .Z(n15213) );
  AND U14589 ( .A(n683), .B(n15218), .Z(n15217) );
  XOR U14590 ( .A(n15219), .B(n15220), .Z(n15211) );
  AND U14591 ( .A(n687), .B(n15221), .Z(n15220) );
  XOR U14592 ( .A(n15222), .B(n15223), .Z(n15208) );
  AND U14593 ( .A(n691), .B(n15221), .Z(n15223) );
  XNOR U14594 ( .A(n15224), .B(n15222), .Z(n15221) );
  IV U14595 ( .A(n15219), .Z(n15224) );
  XOR U14596 ( .A(n15225), .B(n15226), .Z(n15219) );
  AND U14597 ( .A(n694), .B(n15218), .Z(n15226) );
  XNOR U14598 ( .A(n15216), .B(n15225), .Z(n15218) );
  XNOR U14599 ( .A(n15227), .B(n15228), .Z(n15216) );
  AND U14600 ( .A(n698), .B(n15229), .Z(n15228) );
  XOR U14601 ( .A(p_input[529]), .B(n15227), .Z(n15229) );
  XNOR U14602 ( .A(n15230), .B(n15231), .Z(n15227) );
  AND U14603 ( .A(n702), .B(n15232), .Z(n15231) );
  XOR U14604 ( .A(n15233), .B(n15234), .Z(n15225) );
  AND U14605 ( .A(n706), .B(n15235), .Z(n15234) );
  XOR U14606 ( .A(n15236), .B(n15237), .Z(n15222) );
  AND U14607 ( .A(n710), .B(n15235), .Z(n15237) );
  XNOR U14608 ( .A(n15238), .B(n15236), .Z(n15235) );
  IV U14609 ( .A(n15233), .Z(n15238) );
  XOR U14610 ( .A(n15239), .B(n15240), .Z(n15233) );
  AND U14611 ( .A(n713), .B(n15232), .Z(n15240) );
  XNOR U14612 ( .A(n15230), .B(n15239), .Z(n15232) );
  XNOR U14613 ( .A(n15241), .B(n15242), .Z(n15230) );
  AND U14614 ( .A(n717), .B(n15243), .Z(n15242) );
  XOR U14615 ( .A(p_input[545]), .B(n15241), .Z(n15243) );
  XNOR U14616 ( .A(n15244), .B(n15245), .Z(n15241) );
  AND U14617 ( .A(n721), .B(n15246), .Z(n15245) );
  XOR U14618 ( .A(n15247), .B(n15248), .Z(n15239) );
  AND U14619 ( .A(n725), .B(n15249), .Z(n15248) );
  XOR U14620 ( .A(n15250), .B(n15251), .Z(n15236) );
  AND U14621 ( .A(n729), .B(n15249), .Z(n15251) );
  XNOR U14622 ( .A(n15252), .B(n15250), .Z(n15249) );
  IV U14623 ( .A(n15247), .Z(n15252) );
  XOR U14624 ( .A(n15253), .B(n15254), .Z(n15247) );
  AND U14625 ( .A(n732), .B(n15246), .Z(n15254) );
  XNOR U14626 ( .A(n15244), .B(n15253), .Z(n15246) );
  XNOR U14627 ( .A(n15255), .B(n15256), .Z(n15244) );
  AND U14628 ( .A(n736), .B(n15257), .Z(n15256) );
  XOR U14629 ( .A(p_input[561]), .B(n15255), .Z(n15257) );
  XNOR U14630 ( .A(n15258), .B(n15259), .Z(n15255) );
  AND U14631 ( .A(n740), .B(n15260), .Z(n15259) );
  XOR U14632 ( .A(n15261), .B(n15262), .Z(n15253) );
  AND U14633 ( .A(n744), .B(n15263), .Z(n15262) );
  XOR U14634 ( .A(n15264), .B(n15265), .Z(n15250) );
  AND U14635 ( .A(n748), .B(n15263), .Z(n15265) );
  XNOR U14636 ( .A(n15266), .B(n15264), .Z(n15263) );
  IV U14637 ( .A(n15261), .Z(n15266) );
  XOR U14638 ( .A(n15267), .B(n15268), .Z(n15261) );
  AND U14639 ( .A(n751), .B(n15260), .Z(n15268) );
  XNOR U14640 ( .A(n15258), .B(n15267), .Z(n15260) );
  XNOR U14641 ( .A(n15269), .B(n15270), .Z(n15258) );
  AND U14642 ( .A(n755), .B(n15271), .Z(n15270) );
  XOR U14643 ( .A(p_input[577]), .B(n15269), .Z(n15271) );
  XNOR U14644 ( .A(n15272), .B(n15273), .Z(n15269) );
  AND U14645 ( .A(n759), .B(n15274), .Z(n15273) );
  XOR U14646 ( .A(n15275), .B(n15276), .Z(n15267) );
  AND U14647 ( .A(n763), .B(n15277), .Z(n15276) );
  XOR U14648 ( .A(n15278), .B(n15279), .Z(n15264) );
  AND U14649 ( .A(n767), .B(n15277), .Z(n15279) );
  XNOR U14650 ( .A(n15280), .B(n15278), .Z(n15277) );
  IV U14651 ( .A(n15275), .Z(n15280) );
  XOR U14652 ( .A(n15281), .B(n15282), .Z(n15275) );
  AND U14653 ( .A(n770), .B(n15274), .Z(n15282) );
  XNOR U14654 ( .A(n15272), .B(n15281), .Z(n15274) );
  XNOR U14655 ( .A(n15283), .B(n15284), .Z(n15272) );
  AND U14656 ( .A(n774), .B(n15285), .Z(n15284) );
  XOR U14657 ( .A(p_input[593]), .B(n15283), .Z(n15285) );
  XNOR U14658 ( .A(n15286), .B(n15287), .Z(n15283) );
  AND U14659 ( .A(n778), .B(n15288), .Z(n15287) );
  XOR U14660 ( .A(n15289), .B(n15290), .Z(n15281) );
  AND U14661 ( .A(n782), .B(n15291), .Z(n15290) );
  XOR U14662 ( .A(n15292), .B(n15293), .Z(n15278) );
  AND U14663 ( .A(n786), .B(n15291), .Z(n15293) );
  XNOR U14664 ( .A(n15294), .B(n15292), .Z(n15291) );
  IV U14665 ( .A(n15289), .Z(n15294) );
  XOR U14666 ( .A(n15295), .B(n15296), .Z(n15289) );
  AND U14667 ( .A(n789), .B(n15288), .Z(n15296) );
  XNOR U14668 ( .A(n15286), .B(n15295), .Z(n15288) );
  XNOR U14669 ( .A(n15297), .B(n15298), .Z(n15286) );
  AND U14670 ( .A(n793), .B(n15299), .Z(n15298) );
  XOR U14671 ( .A(p_input[609]), .B(n15297), .Z(n15299) );
  XNOR U14672 ( .A(n15300), .B(n15301), .Z(n15297) );
  AND U14673 ( .A(n797), .B(n15302), .Z(n15301) );
  XOR U14674 ( .A(n15303), .B(n15304), .Z(n15295) );
  AND U14675 ( .A(n801), .B(n15305), .Z(n15304) );
  XOR U14676 ( .A(n15306), .B(n15307), .Z(n15292) );
  AND U14677 ( .A(n805), .B(n15305), .Z(n15307) );
  XNOR U14678 ( .A(n15308), .B(n15306), .Z(n15305) );
  IV U14679 ( .A(n15303), .Z(n15308) );
  XOR U14680 ( .A(n15309), .B(n15310), .Z(n15303) );
  AND U14681 ( .A(n808), .B(n15302), .Z(n15310) );
  XNOR U14682 ( .A(n15300), .B(n15309), .Z(n15302) );
  XNOR U14683 ( .A(n15311), .B(n15312), .Z(n15300) );
  AND U14684 ( .A(n812), .B(n15313), .Z(n15312) );
  XOR U14685 ( .A(p_input[625]), .B(n15311), .Z(n15313) );
  XNOR U14686 ( .A(n15314), .B(n15315), .Z(n15311) );
  AND U14687 ( .A(n816), .B(n15316), .Z(n15315) );
  XOR U14688 ( .A(n15317), .B(n15318), .Z(n15309) );
  AND U14689 ( .A(n820), .B(n15319), .Z(n15318) );
  XOR U14690 ( .A(n15320), .B(n15321), .Z(n15306) );
  AND U14691 ( .A(n824), .B(n15319), .Z(n15321) );
  XNOR U14692 ( .A(n15322), .B(n15320), .Z(n15319) );
  IV U14693 ( .A(n15317), .Z(n15322) );
  XOR U14694 ( .A(n15323), .B(n15324), .Z(n15317) );
  AND U14695 ( .A(n827), .B(n15316), .Z(n15324) );
  XNOR U14696 ( .A(n15314), .B(n15323), .Z(n15316) );
  XNOR U14697 ( .A(n15325), .B(n15326), .Z(n15314) );
  AND U14698 ( .A(n831), .B(n15327), .Z(n15326) );
  XOR U14699 ( .A(p_input[641]), .B(n15325), .Z(n15327) );
  XNOR U14700 ( .A(n15328), .B(n15329), .Z(n15325) );
  AND U14701 ( .A(n835), .B(n15330), .Z(n15329) );
  XOR U14702 ( .A(n15331), .B(n15332), .Z(n15323) );
  AND U14703 ( .A(n839), .B(n15333), .Z(n15332) );
  XOR U14704 ( .A(n15334), .B(n15335), .Z(n15320) );
  AND U14705 ( .A(n843), .B(n15333), .Z(n15335) );
  XNOR U14706 ( .A(n15336), .B(n15334), .Z(n15333) );
  IV U14707 ( .A(n15331), .Z(n15336) );
  XOR U14708 ( .A(n15337), .B(n15338), .Z(n15331) );
  AND U14709 ( .A(n846), .B(n15330), .Z(n15338) );
  XNOR U14710 ( .A(n15328), .B(n15337), .Z(n15330) );
  XNOR U14711 ( .A(n15339), .B(n15340), .Z(n15328) );
  AND U14712 ( .A(n850), .B(n15341), .Z(n15340) );
  XOR U14713 ( .A(p_input[657]), .B(n15339), .Z(n15341) );
  XNOR U14714 ( .A(n15342), .B(n15343), .Z(n15339) );
  AND U14715 ( .A(n854), .B(n15344), .Z(n15343) );
  XOR U14716 ( .A(n15345), .B(n15346), .Z(n15337) );
  AND U14717 ( .A(n858), .B(n15347), .Z(n15346) );
  XOR U14718 ( .A(n15348), .B(n15349), .Z(n15334) );
  AND U14719 ( .A(n862), .B(n15347), .Z(n15349) );
  XNOR U14720 ( .A(n15350), .B(n15348), .Z(n15347) );
  IV U14721 ( .A(n15345), .Z(n15350) );
  XOR U14722 ( .A(n15351), .B(n15352), .Z(n15345) );
  AND U14723 ( .A(n865), .B(n15344), .Z(n15352) );
  XNOR U14724 ( .A(n15342), .B(n15351), .Z(n15344) );
  XNOR U14725 ( .A(n15353), .B(n15354), .Z(n15342) );
  AND U14726 ( .A(n869), .B(n15355), .Z(n15354) );
  XOR U14727 ( .A(p_input[673]), .B(n15353), .Z(n15355) );
  XNOR U14728 ( .A(n15356), .B(n15357), .Z(n15353) );
  AND U14729 ( .A(n873), .B(n15358), .Z(n15357) );
  XOR U14730 ( .A(n15359), .B(n15360), .Z(n15351) );
  AND U14731 ( .A(n877), .B(n15361), .Z(n15360) );
  XOR U14732 ( .A(n15362), .B(n15363), .Z(n15348) );
  AND U14733 ( .A(n881), .B(n15361), .Z(n15363) );
  XNOR U14734 ( .A(n15364), .B(n15362), .Z(n15361) );
  IV U14735 ( .A(n15359), .Z(n15364) );
  XOR U14736 ( .A(n15365), .B(n15366), .Z(n15359) );
  AND U14737 ( .A(n884), .B(n15358), .Z(n15366) );
  XNOR U14738 ( .A(n15356), .B(n15365), .Z(n15358) );
  XNOR U14739 ( .A(n15367), .B(n15368), .Z(n15356) );
  AND U14740 ( .A(n888), .B(n15369), .Z(n15368) );
  XOR U14741 ( .A(p_input[689]), .B(n15367), .Z(n15369) );
  XNOR U14742 ( .A(n15370), .B(n15371), .Z(n15367) );
  AND U14743 ( .A(n892), .B(n15372), .Z(n15371) );
  XOR U14744 ( .A(n15373), .B(n15374), .Z(n15365) );
  AND U14745 ( .A(n896), .B(n15375), .Z(n15374) );
  XOR U14746 ( .A(n15376), .B(n15377), .Z(n15362) );
  AND U14747 ( .A(n900), .B(n15375), .Z(n15377) );
  XNOR U14748 ( .A(n15378), .B(n15376), .Z(n15375) );
  IV U14749 ( .A(n15373), .Z(n15378) );
  XOR U14750 ( .A(n15379), .B(n15380), .Z(n15373) );
  AND U14751 ( .A(n903), .B(n15372), .Z(n15380) );
  XNOR U14752 ( .A(n15370), .B(n15379), .Z(n15372) );
  XNOR U14753 ( .A(n15381), .B(n15382), .Z(n15370) );
  AND U14754 ( .A(n907), .B(n15383), .Z(n15382) );
  XOR U14755 ( .A(p_input[705]), .B(n15381), .Z(n15383) );
  XNOR U14756 ( .A(n15384), .B(n15385), .Z(n15381) );
  AND U14757 ( .A(n911), .B(n15386), .Z(n15385) );
  XOR U14758 ( .A(n15387), .B(n15388), .Z(n15379) );
  AND U14759 ( .A(n915), .B(n15389), .Z(n15388) );
  XOR U14760 ( .A(n15390), .B(n15391), .Z(n15376) );
  AND U14761 ( .A(n919), .B(n15389), .Z(n15391) );
  XNOR U14762 ( .A(n15392), .B(n15390), .Z(n15389) );
  IV U14763 ( .A(n15387), .Z(n15392) );
  XOR U14764 ( .A(n15393), .B(n15394), .Z(n15387) );
  AND U14765 ( .A(n922), .B(n15386), .Z(n15394) );
  XNOR U14766 ( .A(n15384), .B(n15393), .Z(n15386) );
  XNOR U14767 ( .A(n15395), .B(n15396), .Z(n15384) );
  AND U14768 ( .A(n926), .B(n15397), .Z(n15396) );
  XOR U14769 ( .A(p_input[721]), .B(n15395), .Z(n15397) );
  XNOR U14770 ( .A(n15398), .B(n15399), .Z(n15395) );
  AND U14771 ( .A(n930), .B(n15400), .Z(n15399) );
  XOR U14772 ( .A(n15401), .B(n15402), .Z(n15393) );
  AND U14773 ( .A(n934), .B(n15403), .Z(n15402) );
  XOR U14774 ( .A(n15404), .B(n15405), .Z(n15390) );
  AND U14775 ( .A(n938), .B(n15403), .Z(n15405) );
  XNOR U14776 ( .A(n15406), .B(n15404), .Z(n15403) );
  IV U14777 ( .A(n15401), .Z(n15406) );
  XOR U14778 ( .A(n15407), .B(n15408), .Z(n15401) );
  AND U14779 ( .A(n941), .B(n15400), .Z(n15408) );
  XNOR U14780 ( .A(n15398), .B(n15407), .Z(n15400) );
  XNOR U14781 ( .A(n15409), .B(n15410), .Z(n15398) );
  AND U14782 ( .A(n945), .B(n15411), .Z(n15410) );
  XOR U14783 ( .A(p_input[737]), .B(n15409), .Z(n15411) );
  XNOR U14784 ( .A(n15412), .B(n15413), .Z(n15409) );
  AND U14785 ( .A(n949), .B(n15414), .Z(n15413) );
  XOR U14786 ( .A(n15415), .B(n15416), .Z(n15407) );
  AND U14787 ( .A(n953), .B(n15417), .Z(n15416) );
  XOR U14788 ( .A(n15418), .B(n15419), .Z(n15404) );
  AND U14789 ( .A(n957), .B(n15417), .Z(n15419) );
  XNOR U14790 ( .A(n15420), .B(n15418), .Z(n15417) );
  IV U14791 ( .A(n15415), .Z(n15420) );
  XOR U14792 ( .A(n15421), .B(n15422), .Z(n15415) );
  AND U14793 ( .A(n960), .B(n15414), .Z(n15422) );
  XNOR U14794 ( .A(n15412), .B(n15421), .Z(n15414) );
  XNOR U14795 ( .A(n15423), .B(n15424), .Z(n15412) );
  AND U14796 ( .A(n964), .B(n15425), .Z(n15424) );
  XOR U14797 ( .A(p_input[753]), .B(n15423), .Z(n15425) );
  XNOR U14798 ( .A(n15426), .B(n15427), .Z(n15423) );
  AND U14799 ( .A(n968), .B(n15428), .Z(n15427) );
  XOR U14800 ( .A(n15429), .B(n15430), .Z(n15421) );
  AND U14801 ( .A(n972), .B(n15431), .Z(n15430) );
  XOR U14802 ( .A(n15432), .B(n15433), .Z(n15418) );
  AND U14803 ( .A(n976), .B(n15431), .Z(n15433) );
  XNOR U14804 ( .A(n15434), .B(n15432), .Z(n15431) );
  IV U14805 ( .A(n15429), .Z(n15434) );
  XOR U14806 ( .A(n15435), .B(n15436), .Z(n15429) );
  AND U14807 ( .A(n979), .B(n15428), .Z(n15436) );
  XNOR U14808 ( .A(n15426), .B(n15435), .Z(n15428) );
  XNOR U14809 ( .A(n15437), .B(n15438), .Z(n15426) );
  AND U14810 ( .A(n983), .B(n15439), .Z(n15438) );
  XOR U14811 ( .A(p_input[769]), .B(n15437), .Z(n15439) );
  XNOR U14812 ( .A(n15440), .B(n15441), .Z(n15437) );
  AND U14813 ( .A(n987), .B(n15442), .Z(n15441) );
  XOR U14814 ( .A(n15443), .B(n15444), .Z(n15435) );
  AND U14815 ( .A(n991), .B(n15445), .Z(n15444) );
  XOR U14816 ( .A(n15446), .B(n15447), .Z(n15432) );
  AND U14817 ( .A(n995), .B(n15445), .Z(n15447) );
  XNOR U14818 ( .A(n15448), .B(n15446), .Z(n15445) );
  IV U14819 ( .A(n15443), .Z(n15448) );
  XOR U14820 ( .A(n15449), .B(n15450), .Z(n15443) );
  AND U14821 ( .A(n998), .B(n15442), .Z(n15450) );
  XNOR U14822 ( .A(n15440), .B(n15449), .Z(n15442) );
  XNOR U14823 ( .A(n15451), .B(n15452), .Z(n15440) );
  AND U14824 ( .A(n1002), .B(n15453), .Z(n15452) );
  XOR U14825 ( .A(p_input[785]), .B(n15451), .Z(n15453) );
  XNOR U14826 ( .A(n15454), .B(n15455), .Z(n15451) );
  AND U14827 ( .A(n1006), .B(n15456), .Z(n15455) );
  XOR U14828 ( .A(n15457), .B(n15458), .Z(n15449) );
  AND U14829 ( .A(n1010), .B(n15459), .Z(n15458) );
  XOR U14830 ( .A(n15460), .B(n15461), .Z(n15446) );
  AND U14831 ( .A(n1014), .B(n15459), .Z(n15461) );
  XNOR U14832 ( .A(n15462), .B(n15460), .Z(n15459) );
  IV U14833 ( .A(n15457), .Z(n15462) );
  XOR U14834 ( .A(n15463), .B(n15464), .Z(n15457) );
  AND U14835 ( .A(n1017), .B(n15456), .Z(n15464) );
  XNOR U14836 ( .A(n15454), .B(n15463), .Z(n15456) );
  XNOR U14837 ( .A(n15465), .B(n15466), .Z(n15454) );
  AND U14838 ( .A(n1021), .B(n15467), .Z(n15466) );
  XOR U14839 ( .A(p_input[801]), .B(n15465), .Z(n15467) );
  XNOR U14840 ( .A(n15468), .B(n15469), .Z(n15465) );
  AND U14841 ( .A(n1025), .B(n15470), .Z(n15469) );
  XOR U14842 ( .A(n15471), .B(n15472), .Z(n15463) );
  AND U14843 ( .A(n1029), .B(n15473), .Z(n15472) );
  XOR U14844 ( .A(n15474), .B(n15475), .Z(n15460) );
  AND U14845 ( .A(n1033), .B(n15473), .Z(n15475) );
  XNOR U14846 ( .A(n15476), .B(n15474), .Z(n15473) );
  IV U14847 ( .A(n15471), .Z(n15476) );
  XOR U14848 ( .A(n15477), .B(n15478), .Z(n15471) );
  AND U14849 ( .A(n1036), .B(n15470), .Z(n15478) );
  XNOR U14850 ( .A(n15468), .B(n15477), .Z(n15470) );
  XNOR U14851 ( .A(n15479), .B(n15480), .Z(n15468) );
  AND U14852 ( .A(n1040), .B(n15481), .Z(n15480) );
  XOR U14853 ( .A(p_input[817]), .B(n15479), .Z(n15481) );
  XNOR U14854 ( .A(n15482), .B(n15483), .Z(n15479) );
  AND U14855 ( .A(n1044), .B(n15484), .Z(n15483) );
  XOR U14856 ( .A(n15485), .B(n15486), .Z(n15477) );
  AND U14857 ( .A(n1048), .B(n15487), .Z(n15486) );
  XOR U14858 ( .A(n15488), .B(n15489), .Z(n15474) );
  AND U14859 ( .A(n1052), .B(n15487), .Z(n15489) );
  XNOR U14860 ( .A(n15490), .B(n15488), .Z(n15487) );
  IV U14861 ( .A(n15485), .Z(n15490) );
  XOR U14862 ( .A(n15491), .B(n15492), .Z(n15485) );
  AND U14863 ( .A(n1055), .B(n15484), .Z(n15492) );
  XNOR U14864 ( .A(n15482), .B(n15491), .Z(n15484) );
  XNOR U14865 ( .A(n15493), .B(n15494), .Z(n15482) );
  AND U14866 ( .A(n1059), .B(n15495), .Z(n15494) );
  XOR U14867 ( .A(p_input[833]), .B(n15493), .Z(n15495) );
  XNOR U14868 ( .A(n15496), .B(n15497), .Z(n15493) );
  AND U14869 ( .A(n1063), .B(n15498), .Z(n15497) );
  XOR U14870 ( .A(n15499), .B(n15500), .Z(n15491) );
  AND U14871 ( .A(n1067), .B(n15501), .Z(n15500) );
  XOR U14872 ( .A(n15502), .B(n15503), .Z(n15488) );
  AND U14873 ( .A(n1071), .B(n15501), .Z(n15503) );
  XNOR U14874 ( .A(n15504), .B(n15502), .Z(n15501) );
  IV U14875 ( .A(n15499), .Z(n15504) );
  XOR U14876 ( .A(n15505), .B(n15506), .Z(n15499) );
  AND U14877 ( .A(n1074), .B(n15498), .Z(n15506) );
  XNOR U14878 ( .A(n15496), .B(n15505), .Z(n15498) );
  XNOR U14879 ( .A(n15507), .B(n15508), .Z(n15496) );
  AND U14880 ( .A(n1078), .B(n15509), .Z(n15508) );
  XOR U14881 ( .A(p_input[849]), .B(n15507), .Z(n15509) );
  XNOR U14882 ( .A(n15510), .B(n15511), .Z(n15507) );
  AND U14883 ( .A(n1082), .B(n15512), .Z(n15511) );
  XOR U14884 ( .A(n15513), .B(n15514), .Z(n15505) );
  AND U14885 ( .A(n1086), .B(n15515), .Z(n15514) );
  XOR U14886 ( .A(n15516), .B(n15517), .Z(n15502) );
  AND U14887 ( .A(n1090), .B(n15515), .Z(n15517) );
  XNOR U14888 ( .A(n15518), .B(n15516), .Z(n15515) );
  IV U14889 ( .A(n15513), .Z(n15518) );
  XOR U14890 ( .A(n15519), .B(n15520), .Z(n15513) );
  AND U14891 ( .A(n1093), .B(n15512), .Z(n15520) );
  XNOR U14892 ( .A(n15510), .B(n15519), .Z(n15512) );
  XNOR U14893 ( .A(n15521), .B(n15522), .Z(n15510) );
  AND U14894 ( .A(n1097), .B(n15523), .Z(n15522) );
  XOR U14895 ( .A(p_input[865]), .B(n15521), .Z(n15523) );
  XNOR U14896 ( .A(n15524), .B(n15525), .Z(n15521) );
  AND U14897 ( .A(n1101), .B(n15526), .Z(n15525) );
  XOR U14898 ( .A(n15527), .B(n15528), .Z(n15519) );
  AND U14899 ( .A(n1105), .B(n15529), .Z(n15528) );
  XOR U14900 ( .A(n15530), .B(n15531), .Z(n15516) );
  AND U14901 ( .A(n1109), .B(n15529), .Z(n15531) );
  XNOR U14902 ( .A(n15532), .B(n15530), .Z(n15529) );
  IV U14903 ( .A(n15527), .Z(n15532) );
  XOR U14904 ( .A(n15533), .B(n15534), .Z(n15527) );
  AND U14905 ( .A(n1112), .B(n15526), .Z(n15534) );
  XNOR U14906 ( .A(n15524), .B(n15533), .Z(n15526) );
  XNOR U14907 ( .A(n15535), .B(n15536), .Z(n15524) );
  AND U14908 ( .A(n1116), .B(n15537), .Z(n15536) );
  XOR U14909 ( .A(p_input[881]), .B(n15535), .Z(n15537) );
  XNOR U14910 ( .A(n15538), .B(n15539), .Z(n15535) );
  AND U14911 ( .A(n1120), .B(n15540), .Z(n15539) );
  XOR U14912 ( .A(n15541), .B(n15542), .Z(n15533) );
  AND U14913 ( .A(n1124), .B(n15543), .Z(n15542) );
  XOR U14914 ( .A(n15544), .B(n15545), .Z(n15530) );
  AND U14915 ( .A(n1128), .B(n15543), .Z(n15545) );
  XNOR U14916 ( .A(n15546), .B(n15544), .Z(n15543) );
  IV U14917 ( .A(n15541), .Z(n15546) );
  XOR U14918 ( .A(n15547), .B(n15548), .Z(n15541) );
  AND U14919 ( .A(n1131), .B(n15540), .Z(n15548) );
  XNOR U14920 ( .A(n15538), .B(n15547), .Z(n15540) );
  XNOR U14921 ( .A(n15549), .B(n15550), .Z(n15538) );
  AND U14922 ( .A(n1135), .B(n15551), .Z(n15550) );
  XOR U14923 ( .A(p_input[897]), .B(n15549), .Z(n15551) );
  XNOR U14924 ( .A(n15552), .B(n15553), .Z(n15549) );
  AND U14925 ( .A(n1139), .B(n15554), .Z(n15553) );
  XOR U14926 ( .A(n15555), .B(n15556), .Z(n15547) );
  AND U14927 ( .A(n1143), .B(n15557), .Z(n15556) );
  XOR U14928 ( .A(n15558), .B(n15559), .Z(n15544) );
  AND U14929 ( .A(n1147), .B(n15557), .Z(n15559) );
  XNOR U14930 ( .A(n15560), .B(n15558), .Z(n15557) );
  IV U14931 ( .A(n15555), .Z(n15560) );
  XOR U14932 ( .A(n15561), .B(n15562), .Z(n15555) );
  AND U14933 ( .A(n1150), .B(n15554), .Z(n15562) );
  XNOR U14934 ( .A(n15552), .B(n15561), .Z(n15554) );
  XNOR U14935 ( .A(n15563), .B(n15564), .Z(n15552) );
  AND U14936 ( .A(n1154), .B(n15565), .Z(n15564) );
  XOR U14937 ( .A(p_input[913]), .B(n15563), .Z(n15565) );
  XNOR U14938 ( .A(n15566), .B(n15567), .Z(n15563) );
  AND U14939 ( .A(n1158), .B(n15568), .Z(n15567) );
  XOR U14940 ( .A(n15569), .B(n15570), .Z(n15561) );
  AND U14941 ( .A(n1162), .B(n15571), .Z(n15570) );
  XOR U14942 ( .A(n15572), .B(n15573), .Z(n15558) );
  AND U14943 ( .A(n1166), .B(n15571), .Z(n15573) );
  XNOR U14944 ( .A(n15574), .B(n15572), .Z(n15571) );
  IV U14945 ( .A(n15569), .Z(n15574) );
  XOR U14946 ( .A(n15575), .B(n15576), .Z(n15569) );
  AND U14947 ( .A(n1169), .B(n15568), .Z(n15576) );
  XNOR U14948 ( .A(n15566), .B(n15575), .Z(n15568) );
  XNOR U14949 ( .A(n15577), .B(n15578), .Z(n15566) );
  AND U14950 ( .A(n1173), .B(n15579), .Z(n15578) );
  XOR U14951 ( .A(p_input[929]), .B(n15577), .Z(n15579) );
  XNOR U14952 ( .A(n15580), .B(n15581), .Z(n15577) );
  AND U14953 ( .A(n1177), .B(n15582), .Z(n15581) );
  XOR U14954 ( .A(n15583), .B(n15584), .Z(n15575) );
  AND U14955 ( .A(n1181), .B(n15585), .Z(n15584) );
  XOR U14956 ( .A(n15586), .B(n15587), .Z(n15572) );
  AND U14957 ( .A(n1185), .B(n15585), .Z(n15587) );
  XNOR U14958 ( .A(n15588), .B(n15586), .Z(n15585) );
  IV U14959 ( .A(n15583), .Z(n15588) );
  XOR U14960 ( .A(n15589), .B(n15590), .Z(n15583) );
  AND U14961 ( .A(n1188), .B(n15582), .Z(n15590) );
  XNOR U14962 ( .A(n15580), .B(n15589), .Z(n15582) );
  XNOR U14963 ( .A(n15591), .B(n15592), .Z(n15580) );
  AND U14964 ( .A(n1192), .B(n15593), .Z(n15592) );
  XOR U14965 ( .A(p_input[945]), .B(n15591), .Z(n15593) );
  XNOR U14966 ( .A(n15594), .B(n15595), .Z(n15591) );
  AND U14967 ( .A(n1196), .B(n15596), .Z(n15595) );
  XOR U14968 ( .A(n15597), .B(n15598), .Z(n15589) );
  AND U14969 ( .A(n1200), .B(n15599), .Z(n15598) );
  XOR U14970 ( .A(n15600), .B(n15601), .Z(n15586) );
  AND U14971 ( .A(n1204), .B(n15599), .Z(n15601) );
  XNOR U14972 ( .A(n15602), .B(n15600), .Z(n15599) );
  IV U14973 ( .A(n15597), .Z(n15602) );
  XOR U14974 ( .A(n15603), .B(n15604), .Z(n15597) );
  AND U14975 ( .A(n1207), .B(n15596), .Z(n15604) );
  XNOR U14976 ( .A(n15594), .B(n15603), .Z(n15596) );
  XNOR U14977 ( .A(n15605), .B(n15606), .Z(n15594) );
  AND U14978 ( .A(n1211), .B(n15607), .Z(n15606) );
  XOR U14979 ( .A(p_input[961]), .B(n15605), .Z(n15607) );
  XNOR U14980 ( .A(n15608), .B(n15609), .Z(n15605) );
  AND U14981 ( .A(n1215), .B(n15610), .Z(n15609) );
  XOR U14982 ( .A(n15611), .B(n15612), .Z(n15603) );
  AND U14983 ( .A(n1219), .B(n15613), .Z(n15612) );
  XOR U14984 ( .A(n15614), .B(n15615), .Z(n15600) );
  AND U14985 ( .A(n1223), .B(n15613), .Z(n15615) );
  XNOR U14986 ( .A(n15616), .B(n15614), .Z(n15613) );
  IV U14987 ( .A(n15611), .Z(n15616) );
  XOR U14988 ( .A(n15617), .B(n15618), .Z(n15611) );
  AND U14989 ( .A(n1226), .B(n15610), .Z(n15618) );
  XNOR U14990 ( .A(n15608), .B(n15617), .Z(n15610) );
  XNOR U14991 ( .A(n15619), .B(n15620), .Z(n15608) );
  AND U14992 ( .A(n1230), .B(n15621), .Z(n15620) );
  XOR U14993 ( .A(p_input[977]), .B(n15619), .Z(n15621) );
  XNOR U14994 ( .A(n15622), .B(n15623), .Z(n15619) );
  AND U14995 ( .A(n1234), .B(n15624), .Z(n15623) );
  XOR U14996 ( .A(n15625), .B(n15626), .Z(n15617) );
  AND U14997 ( .A(n1238), .B(n15627), .Z(n15626) );
  XOR U14998 ( .A(n15628), .B(n15629), .Z(n15614) );
  AND U14999 ( .A(n1242), .B(n15627), .Z(n15629) );
  XNOR U15000 ( .A(n15630), .B(n15628), .Z(n15627) );
  IV U15001 ( .A(n15625), .Z(n15630) );
  XOR U15002 ( .A(n15631), .B(n15632), .Z(n15625) );
  AND U15003 ( .A(n1245), .B(n15624), .Z(n15632) );
  XNOR U15004 ( .A(n15622), .B(n15631), .Z(n15624) );
  XNOR U15005 ( .A(n15633), .B(n15634), .Z(n15622) );
  AND U15006 ( .A(n1249), .B(n15635), .Z(n15634) );
  XOR U15007 ( .A(p_input[993]), .B(n15633), .Z(n15635) );
  XNOR U15008 ( .A(n15636), .B(n15637), .Z(n15633) );
  AND U15009 ( .A(n1253), .B(n15638), .Z(n15637) );
  XOR U15010 ( .A(n15639), .B(n15640), .Z(n15631) );
  AND U15011 ( .A(n1257), .B(n15641), .Z(n15640) );
  XOR U15012 ( .A(n15642), .B(n15643), .Z(n15628) );
  AND U15013 ( .A(n1261), .B(n15641), .Z(n15643) );
  XNOR U15014 ( .A(n15644), .B(n15642), .Z(n15641) );
  IV U15015 ( .A(n15639), .Z(n15644) );
  XOR U15016 ( .A(n15645), .B(n15646), .Z(n15639) );
  AND U15017 ( .A(n1264), .B(n15638), .Z(n15646) );
  XNOR U15018 ( .A(n15636), .B(n15645), .Z(n15638) );
  XNOR U15019 ( .A(n15647), .B(n15648), .Z(n15636) );
  AND U15020 ( .A(n1268), .B(n15649), .Z(n15648) );
  XOR U15021 ( .A(p_input[1009]), .B(n15647), .Z(n15649) );
  XNOR U15022 ( .A(n15650), .B(n15651), .Z(n15647) );
  AND U15023 ( .A(n1272), .B(n15652), .Z(n15651) );
  XOR U15024 ( .A(n15653), .B(n15654), .Z(n15645) );
  AND U15025 ( .A(n1276), .B(n15655), .Z(n15654) );
  XOR U15026 ( .A(n15656), .B(n15657), .Z(n15642) );
  AND U15027 ( .A(n1280), .B(n15655), .Z(n15657) );
  XNOR U15028 ( .A(n15658), .B(n15656), .Z(n15655) );
  IV U15029 ( .A(n15653), .Z(n15658) );
  XOR U15030 ( .A(n15659), .B(n15660), .Z(n15653) );
  AND U15031 ( .A(n1283), .B(n15652), .Z(n15660) );
  XNOR U15032 ( .A(n15650), .B(n15659), .Z(n15652) );
  XNOR U15033 ( .A(n15661), .B(n15662), .Z(n15650) );
  AND U15034 ( .A(n1287), .B(n15663), .Z(n15662) );
  XOR U15035 ( .A(p_input[1025]), .B(n15661), .Z(n15663) );
  XNOR U15036 ( .A(n15664), .B(n15665), .Z(n15661) );
  AND U15037 ( .A(n1291), .B(n15666), .Z(n15665) );
  XOR U15038 ( .A(n15667), .B(n15668), .Z(n15659) );
  AND U15039 ( .A(n1295), .B(n15669), .Z(n15668) );
  XOR U15040 ( .A(n15670), .B(n15671), .Z(n15656) );
  AND U15041 ( .A(n1299), .B(n15669), .Z(n15671) );
  XNOR U15042 ( .A(n15672), .B(n15670), .Z(n15669) );
  IV U15043 ( .A(n15667), .Z(n15672) );
  XOR U15044 ( .A(n15673), .B(n15674), .Z(n15667) );
  AND U15045 ( .A(n1302), .B(n15666), .Z(n15674) );
  XNOR U15046 ( .A(n15664), .B(n15673), .Z(n15666) );
  XNOR U15047 ( .A(n15675), .B(n15676), .Z(n15664) );
  AND U15048 ( .A(n1306), .B(n15677), .Z(n15676) );
  XOR U15049 ( .A(p_input[1041]), .B(n15675), .Z(n15677) );
  XNOR U15050 ( .A(n15678), .B(n15679), .Z(n15675) );
  AND U15051 ( .A(n1310), .B(n15680), .Z(n15679) );
  XOR U15052 ( .A(n15681), .B(n15682), .Z(n15673) );
  AND U15053 ( .A(n1314), .B(n15683), .Z(n15682) );
  XOR U15054 ( .A(n15684), .B(n15685), .Z(n15670) );
  AND U15055 ( .A(n1318), .B(n15683), .Z(n15685) );
  XNOR U15056 ( .A(n15686), .B(n15684), .Z(n15683) );
  IV U15057 ( .A(n15681), .Z(n15686) );
  XOR U15058 ( .A(n15687), .B(n15688), .Z(n15681) );
  AND U15059 ( .A(n1321), .B(n15680), .Z(n15688) );
  XNOR U15060 ( .A(n15678), .B(n15687), .Z(n15680) );
  XNOR U15061 ( .A(n15689), .B(n15690), .Z(n15678) );
  AND U15062 ( .A(n1325), .B(n15691), .Z(n15690) );
  XOR U15063 ( .A(p_input[1057]), .B(n15689), .Z(n15691) );
  XNOR U15064 ( .A(n15692), .B(n15693), .Z(n15689) );
  AND U15065 ( .A(n1329), .B(n15694), .Z(n15693) );
  XOR U15066 ( .A(n15695), .B(n15696), .Z(n15687) );
  AND U15067 ( .A(n1333), .B(n15697), .Z(n15696) );
  XOR U15068 ( .A(n15698), .B(n15699), .Z(n15684) );
  AND U15069 ( .A(n1337), .B(n15697), .Z(n15699) );
  XNOR U15070 ( .A(n15700), .B(n15698), .Z(n15697) );
  IV U15071 ( .A(n15695), .Z(n15700) );
  XOR U15072 ( .A(n15701), .B(n15702), .Z(n15695) );
  AND U15073 ( .A(n1340), .B(n15694), .Z(n15702) );
  XNOR U15074 ( .A(n15692), .B(n15701), .Z(n15694) );
  XNOR U15075 ( .A(n15703), .B(n15704), .Z(n15692) );
  AND U15076 ( .A(n1344), .B(n15705), .Z(n15704) );
  XOR U15077 ( .A(p_input[1073]), .B(n15703), .Z(n15705) );
  XNOR U15078 ( .A(n15706), .B(n15707), .Z(n15703) );
  AND U15079 ( .A(n1348), .B(n15708), .Z(n15707) );
  XOR U15080 ( .A(n15709), .B(n15710), .Z(n15701) );
  AND U15081 ( .A(n1352), .B(n15711), .Z(n15710) );
  XOR U15082 ( .A(n15712), .B(n15713), .Z(n15698) );
  AND U15083 ( .A(n1356), .B(n15711), .Z(n15713) );
  XNOR U15084 ( .A(n15714), .B(n15712), .Z(n15711) );
  IV U15085 ( .A(n15709), .Z(n15714) );
  XOR U15086 ( .A(n15715), .B(n15716), .Z(n15709) );
  AND U15087 ( .A(n1359), .B(n15708), .Z(n15716) );
  XNOR U15088 ( .A(n15706), .B(n15715), .Z(n15708) );
  XNOR U15089 ( .A(n15717), .B(n15718), .Z(n15706) );
  AND U15090 ( .A(n1363), .B(n15719), .Z(n15718) );
  XOR U15091 ( .A(p_input[1089]), .B(n15717), .Z(n15719) );
  XNOR U15092 ( .A(n15720), .B(n15721), .Z(n15717) );
  AND U15093 ( .A(n1367), .B(n15722), .Z(n15721) );
  XOR U15094 ( .A(n15723), .B(n15724), .Z(n15715) );
  AND U15095 ( .A(n1371), .B(n15725), .Z(n15724) );
  XOR U15096 ( .A(n15726), .B(n15727), .Z(n15712) );
  AND U15097 ( .A(n1375), .B(n15725), .Z(n15727) );
  XNOR U15098 ( .A(n15728), .B(n15726), .Z(n15725) );
  IV U15099 ( .A(n15723), .Z(n15728) );
  XOR U15100 ( .A(n15729), .B(n15730), .Z(n15723) );
  AND U15101 ( .A(n1378), .B(n15722), .Z(n15730) );
  XNOR U15102 ( .A(n15720), .B(n15729), .Z(n15722) );
  XNOR U15103 ( .A(n15731), .B(n15732), .Z(n15720) );
  AND U15104 ( .A(n1382), .B(n15733), .Z(n15732) );
  XOR U15105 ( .A(p_input[1105]), .B(n15731), .Z(n15733) );
  XNOR U15106 ( .A(n15734), .B(n15735), .Z(n15731) );
  AND U15107 ( .A(n1386), .B(n15736), .Z(n15735) );
  XOR U15108 ( .A(n15737), .B(n15738), .Z(n15729) );
  AND U15109 ( .A(n1390), .B(n15739), .Z(n15738) );
  XOR U15110 ( .A(n15740), .B(n15741), .Z(n15726) );
  AND U15111 ( .A(n1394), .B(n15739), .Z(n15741) );
  XNOR U15112 ( .A(n15742), .B(n15740), .Z(n15739) );
  IV U15113 ( .A(n15737), .Z(n15742) );
  XOR U15114 ( .A(n15743), .B(n15744), .Z(n15737) );
  AND U15115 ( .A(n1397), .B(n15736), .Z(n15744) );
  XNOR U15116 ( .A(n15734), .B(n15743), .Z(n15736) );
  XNOR U15117 ( .A(n15745), .B(n15746), .Z(n15734) );
  AND U15118 ( .A(n1401), .B(n15747), .Z(n15746) );
  XOR U15119 ( .A(p_input[1121]), .B(n15745), .Z(n15747) );
  XNOR U15120 ( .A(n15748), .B(n15749), .Z(n15745) );
  AND U15121 ( .A(n1405), .B(n15750), .Z(n15749) );
  XOR U15122 ( .A(n15751), .B(n15752), .Z(n15743) );
  AND U15123 ( .A(n1409), .B(n15753), .Z(n15752) );
  XOR U15124 ( .A(n15754), .B(n15755), .Z(n15740) );
  AND U15125 ( .A(n1413), .B(n15753), .Z(n15755) );
  XNOR U15126 ( .A(n15756), .B(n15754), .Z(n15753) );
  IV U15127 ( .A(n15751), .Z(n15756) );
  XOR U15128 ( .A(n15757), .B(n15758), .Z(n15751) );
  AND U15129 ( .A(n1416), .B(n15750), .Z(n15758) );
  XNOR U15130 ( .A(n15748), .B(n15757), .Z(n15750) );
  XNOR U15131 ( .A(n15759), .B(n15760), .Z(n15748) );
  AND U15132 ( .A(n1420), .B(n15761), .Z(n15760) );
  XOR U15133 ( .A(p_input[1137]), .B(n15759), .Z(n15761) );
  XNOR U15134 ( .A(n15762), .B(n15763), .Z(n15759) );
  AND U15135 ( .A(n1424), .B(n15764), .Z(n15763) );
  XOR U15136 ( .A(n15765), .B(n15766), .Z(n15757) );
  AND U15137 ( .A(n1428), .B(n15767), .Z(n15766) );
  XOR U15138 ( .A(n15768), .B(n15769), .Z(n15754) );
  AND U15139 ( .A(n1432), .B(n15767), .Z(n15769) );
  XNOR U15140 ( .A(n15770), .B(n15768), .Z(n15767) );
  IV U15141 ( .A(n15765), .Z(n15770) );
  XOR U15142 ( .A(n15771), .B(n15772), .Z(n15765) );
  AND U15143 ( .A(n1435), .B(n15764), .Z(n15772) );
  XNOR U15144 ( .A(n15762), .B(n15771), .Z(n15764) );
  XNOR U15145 ( .A(n15773), .B(n15774), .Z(n15762) );
  AND U15146 ( .A(n1439), .B(n15775), .Z(n15774) );
  XOR U15147 ( .A(p_input[1153]), .B(n15773), .Z(n15775) );
  XNOR U15148 ( .A(n15776), .B(n15777), .Z(n15773) );
  AND U15149 ( .A(n1443), .B(n15778), .Z(n15777) );
  XOR U15150 ( .A(n15779), .B(n15780), .Z(n15771) );
  AND U15151 ( .A(n1447), .B(n15781), .Z(n15780) );
  XOR U15152 ( .A(n15782), .B(n15783), .Z(n15768) );
  AND U15153 ( .A(n1451), .B(n15781), .Z(n15783) );
  XNOR U15154 ( .A(n15784), .B(n15782), .Z(n15781) );
  IV U15155 ( .A(n15779), .Z(n15784) );
  XOR U15156 ( .A(n15785), .B(n15786), .Z(n15779) );
  AND U15157 ( .A(n1454), .B(n15778), .Z(n15786) );
  XNOR U15158 ( .A(n15776), .B(n15785), .Z(n15778) );
  XNOR U15159 ( .A(n15787), .B(n15788), .Z(n15776) );
  AND U15160 ( .A(n1458), .B(n15789), .Z(n15788) );
  XOR U15161 ( .A(p_input[1169]), .B(n15787), .Z(n15789) );
  XNOR U15162 ( .A(n15790), .B(n15791), .Z(n15787) );
  AND U15163 ( .A(n1462), .B(n15792), .Z(n15791) );
  XOR U15164 ( .A(n15793), .B(n15794), .Z(n15785) );
  AND U15165 ( .A(n1466), .B(n15795), .Z(n15794) );
  XOR U15166 ( .A(n15796), .B(n15797), .Z(n15782) );
  AND U15167 ( .A(n1470), .B(n15795), .Z(n15797) );
  XNOR U15168 ( .A(n15798), .B(n15796), .Z(n15795) );
  IV U15169 ( .A(n15793), .Z(n15798) );
  XOR U15170 ( .A(n15799), .B(n15800), .Z(n15793) );
  AND U15171 ( .A(n1473), .B(n15792), .Z(n15800) );
  XNOR U15172 ( .A(n15790), .B(n15799), .Z(n15792) );
  XNOR U15173 ( .A(n15801), .B(n15802), .Z(n15790) );
  AND U15174 ( .A(n1477), .B(n15803), .Z(n15802) );
  XOR U15175 ( .A(p_input[1185]), .B(n15801), .Z(n15803) );
  XNOR U15176 ( .A(n15804), .B(n15805), .Z(n15801) );
  AND U15177 ( .A(n1481), .B(n15806), .Z(n15805) );
  XOR U15178 ( .A(n15807), .B(n15808), .Z(n15799) );
  AND U15179 ( .A(n1485), .B(n15809), .Z(n15808) );
  XOR U15180 ( .A(n15810), .B(n15811), .Z(n15796) );
  AND U15181 ( .A(n1489), .B(n15809), .Z(n15811) );
  XNOR U15182 ( .A(n15812), .B(n15810), .Z(n15809) );
  IV U15183 ( .A(n15807), .Z(n15812) );
  XOR U15184 ( .A(n15813), .B(n15814), .Z(n15807) );
  AND U15185 ( .A(n1492), .B(n15806), .Z(n15814) );
  XNOR U15186 ( .A(n15804), .B(n15813), .Z(n15806) );
  XNOR U15187 ( .A(n15815), .B(n15816), .Z(n15804) );
  AND U15188 ( .A(n1496), .B(n15817), .Z(n15816) );
  XOR U15189 ( .A(p_input[1201]), .B(n15815), .Z(n15817) );
  XNOR U15190 ( .A(n15818), .B(n15819), .Z(n15815) );
  AND U15191 ( .A(n1500), .B(n15820), .Z(n15819) );
  XOR U15192 ( .A(n15821), .B(n15822), .Z(n15813) );
  AND U15193 ( .A(n1504), .B(n15823), .Z(n15822) );
  XOR U15194 ( .A(n15824), .B(n15825), .Z(n15810) );
  AND U15195 ( .A(n1508), .B(n15823), .Z(n15825) );
  XNOR U15196 ( .A(n15826), .B(n15824), .Z(n15823) );
  IV U15197 ( .A(n15821), .Z(n15826) );
  XOR U15198 ( .A(n15827), .B(n15828), .Z(n15821) );
  AND U15199 ( .A(n1511), .B(n15820), .Z(n15828) );
  XNOR U15200 ( .A(n15818), .B(n15827), .Z(n15820) );
  XNOR U15201 ( .A(n15829), .B(n15830), .Z(n15818) );
  AND U15202 ( .A(n1515), .B(n15831), .Z(n15830) );
  XOR U15203 ( .A(p_input[1217]), .B(n15829), .Z(n15831) );
  XNOR U15204 ( .A(n15832), .B(n15833), .Z(n15829) );
  AND U15205 ( .A(n1519), .B(n15834), .Z(n15833) );
  XOR U15206 ( .A(n15835), .B(n15836), .Z(n15827) );
  AND U15207 ( .A(n1523), .B(n15837), .Z(n15836) );
  XOR U15208 ( .A(n15838), .B(n15839), .Z(n15824) );
  AND U15209 ( .A(n1527), .B(n15837), .Z(n15839) );
  XNOR U15210 ( .A(n15840), .B(n15838), .Z(n15837) );
  IV U15211 ( .A(n15835), .Z(n15840) );
  XOR U15212 ( .A(n15841), .B(n15842), .Z(n15835) );
  AND U15213 ( .A(n1530), .B(n15834), .Z(n15842) );
  XNOR U15214 ( .A(n15832), .B(n15841), .Z(n15834) );
  XNOR U15215 ( .A(n15843), .B(n15844), .Z(n15832) );
  AND U15216 ( .A(n1534), .B(n15845), .Z(n15844) );
  XOR U15217 ( .A(p_input[1233]), .B(n15843), .Z(n15845) );
  XNOR U15218 ( .A(n15846), .B(n15847), .Z(n15843) );
  AND U15219 ( .A(n1538), .B(n15848), .Z(n15847) );
  XOR U15220 ( .A(n15849), .B(n15850), .Z(n15841) );
  AND U15221 ( .A(n1542), .B(n15851), .Z(n15850) );
  XOR U15222 ( .A(n15852), .B(n15853), .Z(n15838) );
  AND U15223 ( .A(n1546), .B(n15851), .Z(n15853) );
  XNOR U15224 ( .A(n15854), .B(n15852), .Z(n15851) );
  IV U15225 ( .A(n15849), .Z(n15854) );
  XOR U15226 ( .A(n15855), .B(n15856), .Z(n15849) );
  AND U15227 ( .A(n1549), .B(n15848), .Z(n15856) );
  XNOR U15228 ( .A(n15846), .B(n15855), .Z(n15848) );
  XNOR U15229 ( .A(n15857), .B(n15858), .Z(n15846) );
  AND U15230 ( .A(n1553), .B(n15859), .Z(n15858) );
  XOR U15231 ( .A(p_input[1249]), .B(n15857), .Z(n15859) );
  XNOR U15232 ( .A(n15860), .B(n15861), .Z(n15857) );
  AND U15233 ( .A(n1557), .B(n15862), .Z(n15861) );
  XOR U15234 ( .A(n15863), .B(n15864), .Z(n15855) );
  AND U15235 ( .A(n1561), .B(n15865), .Z(n15864) );
  XOR U15236 ( .A(n15866), .B(n15867), .Z(n15852) );
  AND U15237 ( .A(n1565), .B(n15865), .Z(n15867) );
  XNOR U15238 ( .A(n15868), .B(n15866), .Z(n15865) );
  IV U15239 ( .A(n15863), .Z(n15868) );
  XOR U15240 ( .A(n15869), .B(n15870), .Z(n15863) );
  AND U15241 ( .A(n1568), .B(n15862), .Z(n15870) );
  XNOR U15242 ( .A(n15860), .B(n15869), .Z(n15862) );
  XNOR U15243 ( .A(n15871), .B(n15872), .Z(n15860) );
  AND U15244 ( .A(n1572), .B(n15873), .Z(n15872) );
  XOR U15245 ( .A(p_input[1265]), .B(n15871), .Z(n15873) );
  XNOR U15246 ( .A(n15874), .B(n15875), .Z(n15871) );
  AND U15247 ( .A(n1576), .B(n15876), .Z(n15875) );
  XOR U15248 ( .A(n15877), .B(n15878), .Z(n15869) );
  AND U15249 ( .A(n1580), .B(n15879), .Z(n15878) );
  XOR U15250 ( .A(n15880), .B(n15881), .Z(n15866) );
  AND U15251 ( .A(n1584), .B(n15879), .Z(n15881) );
  XNOR U15252 ( .A(n15882), .B(n15880), .Z(n15879) );
  IV U15253 ( .A(n15877), .Z(n15882) );
  XOR U15254 ( .A(n15883), .B(n15884), .Z(n15877) );
  AND U15255 ( .A(n1587), .B(n15876), .Z(n15884) );
  XNOR U15256 ( .A(n15874), .B(n15883), .Z(n15876) );
  XNOR U15257 ( .A(n15885), .B(n15886), .Z(n15874) );
  AND U15258 ( .A(n1591), .B(n15887), .Z(n15886) );
  XOR U15259 ( .A(p_input[1281]), .B(n15885), .Z(n15887) );
  XNOR U15260 ( .A(n15888), .B(n15889), .Z(n15885) );
  AND U15261 ( .A(n1595), .B(n15890), .Z(n15889) );
  XOR U15262 ( .A(n15891), .B(n15892), .Z(n15883) );
  AND U15263 ( .A(n1599), .B(n15893), .Z(n15892) );
  XOR U15264 ( .A(n15894), .B(n15895), .Z(n15880) );
  AND U15265 ( .A(n1603), .B(n15893), .Z(n15895) );
  XNOR U15266 ( .A(n15896), .B(n15894), .Z(n15893) );
  IV U15267 ( .A(n15891), .Z(n15896) );
  XOR U15268 ( .A(n15897), .B(n15898), .Z(n15891) );
  AND U15269 ( .A(n1606), .B(n15890), .Z(n15898) );
  XNOR U15270 ( .A(n15888), .B(n15897), .Z(n15890) );
  XNOR U15271 ( .A(n15899), .B(n15900), .Z(n15888) );
  AND U15272 ( .A(n1610), .B(n15901), .Z(n15900) );
  XOR U15273 ( .A(p_input[1297]), .B(n15899), .Z(n15901) );
  XNOR U15274 ( .A(n15902), .B(n15903), .Z(n15899) );
  AND U15275 ( .A(n1614), .B(n15904), .Z(n15903) );
  XOR U15276 ( .A(n15905), .B(n15906), .Z(n15897) );
  AND U15277 ( .A(n1618), .B(n15907), .Z(n15906) );
  XOR U15278 ( .A(n15908), .B(n15909), .Z(n15894) );
  AND U15279 ( .A(n1622), .B(n15907), .Z(n15909) );
  XNOR U15280 ( .A(n15910), .B(n15908), .Z(n15907) );
  IV U15281 ( .A(n15905), .Z(n15910) );
  XOR U15282 ( .A(n15911), .B(n15912), .Z(n15905) );
  AND U15283 ( .A(n1625), .B(n15904), .Z(n15912) );
  XNOR U15284 ( .A(n15902), .B(n15911), .Z(n15904) );
  XNOR U15285 ( .A(n15913), .B(n15914), .Z(n15902) );
  AND U15286 ( .A(n1629), .B(n15915), .Z(n15914) );
  XOR U15287 ( .A(p_input[1313]), .B(n15913), .Z(n15915) );
  XNOR U15288 ( .A(n15916), .B(n15917), .Z(n15913) );
  AND U15289 ( .A(n1633), .B(n15918), .Z(n15917) );
  XOR U15290 ( .A(n15919), .B(n15920), .Z(n15911) );
  AND U15291 ( .A(n1637), .B(n15921), .Z(n15920) );
  XOR U15292 ( .A(n15922), .B(n15923), .Z(n15908) );
  AND U15293 ( .A(n1641), .B(n15921), .Z(n15923) );
  XNOR U15294 ( .A(n15924), .B(n15922), .Z(n15921) );
  IV U15295 ( .A(n15919), .Z(n15924) );
  XOR U15296 ( .A(n15925), .B(n15926), .Z(n15919) );
  AND U15297 ( .A(n1644), .B(n15918), .Z(n15926) );
  XNOR U15298 ( .A(n15916), .B(n15925), .Z(n15918) );
  XNOR U15299 ( .A(n15927), .B(n15928), .Z(n15916) );
  AND U15300 ( .A(n1648), .B(n15929), .Z(n15928) );
  XOR U15301 ( .A(p_input[1329]), .B(n15927), .Z(n15929) );
  XNOR U15302 ( .A(n15930), .B(n15931), .Z(n15927) );
  AND U15303 ( .A(n1652), .B(n15932), .Z(n15931) );
  XOR U15304 ( .A(n15933), .B(n15934), .Z(n15925) );
  AND U15305 ( .A(n1656), .B(n15935), .Z(n15934) );
  XOR U15306 ( .A(n15936), .B(n15937), .Z(n15922) );
  AND U15307 ( .A(n1660), .B(n15935), .Z(n15937) );
  XNOR U15308 ( .A(n15938), .B(n15936), .Z(n15935) );
  IV U15309 ( .A(n15933), .Z(n15938) );
  XOR U15310 ( .A(n15939), .B(n15940), .Z(n15933) );
  AND U15311 ( .A(n1663), .B(n15932), .Z(n15940) );
  XNOR U15312 ( .A(n15930), .B(n15939), .Z(n15932) );
  XNOR U15313 ( .A(n15941), .B(n15942), .Z(n15930) );
  AND U15314 ( .A(n1667), .B(n15943), .Z(n15942) );
  XOR U15315 ( .A(p_input[1345]), .B(n15941), .Z(n15943) );
  XNOR U15316 ( .A(n15944), .B(n15945), .Z(n15941) );
  AND U15317 ( .A(n1671), .B(n15946), .Z(n15945) );
  XOR U15318 ( .A(n15947), .B(n15948), .Z(n15939) );
  AND U15319 ( .A(n1675), .B(n15949), .Z(n15948) );
  XOR U15320 ( .A(n15950), .B(n15951), .Z(n15936) );
  AND U15321 ( .A(n1679), .B(n15949), .Z(n15951) );
  XNOR U15322 ( .A(n15952), .B(n15950), .Z(n15949) );
  IV U15323 ( .A(n15947), .Z(n15952) );
  XOR U15324 ( .A(n15953), .B(n15954), .Z(n15947) );
  AND U15325 ( .A(n1682), .B(n15946), .Z(n15954) );
  XNOR U15326 ( .A(n15944), .B(n15953), .Z(n15946) );
  XNOR U15327 ( .A(n15955), .B(n15956), .Z(n15944) );
  AND U15328 ( .A(n1686), .B(n15957), .Z(n15956) );
  XOR U15329 ( .A(p_input[1361]), .B(n15955), .Z(n15957) );
  XNOR U15330 ( .A(n15958), .B(n15959), .Z(n15955) );
  AND U15331 ( .A(n1690), .B(n15960), .Z(n15959) );
  XOR U15332 ( .A(n15961), .B(n15962), .Z(n15953) );
  AND U15333 ( .A(n1694), .B(n15963), .Z(n15962) );
  XOR U15334 ( .A(n15964), .B(n15965), .Z(n15950) );
  AND U15335 ( .A(n1698), .B(n15963), .Z(n15965) );
  XNOR U15336 ( .A(n15966), .B(n15964), .Z(n15963) );
  IV U15337 ( .A(n15961), .Z(n15966) );
  XOR U15338 ( .A(n15967), .B(n15968), .Z(n15961) );
  AND U15339 ( .A(n1701), .B(n15960), .Z(n15968) );
  XNOR U15340 ( .A(n15958), .B(n15967), .Z(n15960) );
  XNOR U15341 ( .A(n15969), .B(n15970), .Z(n15958) );
  AND U15342 ( .A(n1705), .B(n15971), .Z(n15970) );
  XOR U15343 ( .A(p_input[1377]), .B(n15969), .Z(n15971) );
  XNOR U15344 ( .A(n15972), .B(n15973), .Z(n15969) );
  AND U15345 ( .A(n1709), .B(n15974), .Z(n15973) );
  XOR U15346 ( .A(n15975), .B(n15976), .Z(n15967) );
  AND U15347 ( .A(n1713), .B(n15977), .Z(n15976) );
  XOR U15348 ( .A(n15978), .B(n15979), .Z(n15964) );
  AND U15349 ( .A(n1717), .B(n15977), .Z(n15979) );
  XNOR U15350 ( .A(n15980), .B(n15978), .Z(n15977) );
  IV U15351 ( .A(n15975), .Z(n15980) );
  XOR U15352 ( .A(n15981), .B(n15982), .Z(n15975) );
  AND U15353 ( .A(n1720), .B(n15974), .Z(n15982) );
  XNOR U15354 ( .A(n15972), .B(n15981), .Z(n15974) );
  XNOR U15355 ( .A(n15983), .B(n15984), .Z(n15972) );
  AND U15356 ( .A(n1724), .B(n15985), .Z(n15984) );
  XOR U15357 ( .A(p_input[1393]), .B(n15983), .Z(n15985) );
  XNOR U15358 ( .A(n15986), .B(n15987), .Z(n15983) );
  AND U15359 ( .A(n1728), .B(n15988), .Z(n15987) );
  XOR U15360 ( .A(n15989), .B(n15990), .Z(n15981) );
  AND U15361 ( .A(n1732), .B(n15991), .Z(n15990) );
  XOR U15362 ( .A(n15992), .B(n15993), .Z(n15978) );
  AND U15363 ( .A(n1736), .B(n15991), .Z(n15993) );
  XNOR U15364 ( .A(n15994), .B(n15992), .Z(n15991) );
  IV U15365 ( .A(n15989), .Z(n15994) );
  XOR U15366 ( .A(n15995), .B(n15996), .Z(n15989) );
  AND U15367 ( .A(n1739), .B(n15988), .Z(n15996) );
  XNOR U15368 ( .A(n15986), .B(n15995), .Z(n15988) );
  XNOR U15369 ( .A(n15997), .B(n15998), .Z(n15986) );
  AND U15370 ( .A(n1743), .B(n15999), .Z(n15998) );
  XOR U15371 ( .A(p_input[1409]), .B(n15997), .Z(n15999) );
  XNOR U15372 ( .A(n16000), .B(n16001), .Z(n15997) );
  AND U15373 ( .A(n1747), .B(n16002), .Z(n16001) );
  XOR U15374 ( .A(n16003), .B(n16004), .Z(n15995) );
  AND U15375 ( .A(n1751), .B(n16005), .Z(n16004) );
  XOR U15376 ( .A(n16006), .B(n16007), .Z(n15992) );
  AND U15377 ( .A(n1755), .B(n16005), .Z(n16007) );
  XNOR U15378 ( .A(n16008), .B(n16006), .Z(n16005) );
  IV U15379 ( .A(n16003), .Z(n16008) );
  XOR U15380 ( .A(n16009), .B(n16010), .Z(n16003) );
  AND U15381 ( .A(n1758), .B(n16002), .Z(n16010) );
  XNOR U15382 ( .A(n16000), .B(n16009), .Z(n16002) );
  XNOR U15383 ( .A(n16011), .B(n16012), .Z(n16000) );
  AND U15384 ( .A(n1762), .B(n16013), .Z(n16012) );
  XOR U15385 ( .A(p_input[1425]), .B(n16011), .Z(n16013) );
  XNOR U15386 ( .A(n16014), .B(n16015), .Z(n16011) );
  AND U15387 ( .A(n1766), .B(n16016), .Z(n16015) );
  XOR U15388 ( .A(n16017), .B(n16018), .Z(n16009) );
  AND U15389 ( .A(n1770), .B(n16019), .Z(n16018) );
  XOR U15390 ( .A(n16020), .B(n16021), .Z(n16006) );
  AND U15391 ( .A(n1774), .B(n16019), .Z(n16021) );
  XNOR U15392 ( .A(n16022), .B(n16020), .Z(n16019) );
  IV U15393 ( .A(n16017), .Z(n16022) );
  XOR U15394 ( .A(n16023), .B(n16024), .Z(n16017) );
  AND U15395 ( .A(n1777), .B(n16016), .Z(n16024) );
  XNOR U15396 ( .A(n16014), .B(n16023), .Z(n16016) );
  XNOR U15397 ( .A(n16025), .B(n16026), .Z(n16014) );
  AND U15398 ( .A(n1781), .B(n16027), .Z(n16026) );
  XOR U15399 ( .A(p_input[1441]), .B(n16025), .Z(n16027) );
  XNOR U15400 ( .A(n16028), .B(n16029), .Z(n16025) );
  AND U15401 ( .A(n1785), .B(n16030), .Z(n16029) );
  XOR U15402 ( .A(n16031), .B(n16032), .Z(n16023) );
  AND U15403 ( .A(n1789), .B(n16033), .Z(n16032) );
  XOR U15404 ( .A(n16034), .B(n16035), .Z(n16020) );
  AND U15405 ( .A(n1793), .B(n16033), .Z(n16035) );
  XNOR U15406 ( .A(n16036), .B(n16034), .Z(n16033) );
  IV U15407 ( .A(n16031), .Z(n16036) );
  XOR U15408 ( .A(n16037), .B(n16038), .Z(n16031) );
  AND U15409 ( .A(n1796), .B(n16030), .Z(n16038) );
  XNOR U15410 ( .A(n16028), .B(n16037), .Z(n16030) );
  XNOR U15411 ( .A(n16039), .B(n16040), .Z(n16028) );
  AND U15412 ( .A(n1800), .B(n16041), .Z(n16040) );
  XOR U15413 ( .A(p_input[1457]), .B(n16039), .Z(n16041) );
  XNOR U15414 ( .A(n16042), .B(n16043), .Z(n16039) );
  AND U15415 ( .A(n1804), .B(n16044), .Z(n16043) );
  XOR U15416 ( .A(n16045), .B(n16046), .Z(n16037) );
  AND U15417 ( .A(n1808), .B(n16047), .Z(n16046) );
  XOR U15418 ( .A(n16048), .B(n16049), .Z(n16034) );
  AND U15419 ( .A(n1812), .B(n16047), .Z(n16049) );
  XNOR U15420 ( .A(n16050), .B(n16048), .Z(n16047) );
  IV U15421 ( .A(n16045), .Z(n16050) );
  XOR U15422 ( .A(n16051), .B(n16052), .Z(n16045) );
  AND U15423 ( .A(n1815), .B(n16044), .Z(n16052) );
  XNOR U15424 ( .A(n16042), .B(n16051), .Z(n16044) );
  XNOR U15425 ( .A(n16053), .B(n16054), .Z(n16042) );
  AND U15426 ( .A(n1819), .B(n16055), .Z(n16054) );
  XOR U15427 ( .A(p_input[1473]), .B(n16053), .Z(n16055) );
  XNOR U15428 ( .A(n16056), .B(n16057), .Z(n16053) );
  AND U15429 ( .A(n1823), .B(n16058), .Z(n16057) );
  XOR U15430 ( .A(n16059), .B(n16060), .Z(n16051) );
  AND U15431 ( .A(n1827), .B(n16061), .Z(n16060) );
  XOR U15432 ( .A(n16062), .B(n16063), .Z(n16048) );
  AND U15433 ( .A(n1831), .B(n16061), .Z(n16063) );
  XNOR U15434 ( .A(n16064), .B(n16062), .Z(n16061) );
  IV U15435 ( .A(n16059), .Z(n16064) );
  XOR U15436 ( .A(n16065), .B(n16066), .Z(n16059) );
  AND U15437 ( .A(n1834), .B(n16058), .Z(n16066) );
  XNOR U15438 ( .A(n16056), .B(n16065), .Z(n16058) );
  XNOR U15439 ( .A(n16067), .B(n16068), .Z(n16056) );
  AND U15440 ( .A(n1838), .B(n16069), .Z(n16068) );
  XOR U15441 ( .A(p_input[1489]), .B(n16067), .Z(n16069) );
  XNOR U15442 ( .A(n16070), .B(n16071), .Z(n16067) );
  AND U15443 ( .A(n1842), .B(n16072), .Z(n16071) );
  XOR U15444 ( .A(n16073), .B(n16074), .Z(n16065) );
  AND U15445 ( .A(n1846), .B(n16075), .Z(n16074) );
  XOR U15446 ( .A(n16076), .B(n16077), .Z(n16062) );
  AND U15447 ( .A(n1850), .B(n16075), .Z(n16077) );
  XNOR U15448 ( .A(n16078), .B(n16076), .Z(n16075) );
  IV U15449 ( .A(n16073), .Z(n16078) );
  XOR U15450 ( .A(n16079), .B(n16080), .Z(n16073) );
  AND U15451 ( .A(n1853), .B(n16072), .Z(n16080) );
  XNOR U15452 ( .A(n16070), .B(n16079), .Z(n16072) );
  XNOR U15453 ( .A(n16081), .B(n16082), .Z(n16070) );
  AND U15454 ( .A(n1857), .B(n16083), .Z(n16082) );
  XOR U15455 ( .A(p_input[1505]), .B(n16081), .Z(n16083) );
  XNOR U15456 ( .A(n16084), .B(n16085), .Z(n16081) );
  AND U15457 ( .A(n1861), .B(n16086), .Z(n16085) );
  XOR U15458 ( .A(n16087), .B(n16088), .Z(n16079) );
  AND U15459 ( .A(n1865), .B(n16089), .Z(n16088) );
  XOR U15460 ( .A(n16090), .B(n16091), .Z(n16076) );
  AND U15461 ( .A(n1869), .B(n16089), .Z(n16091) );
  XNOR U15462 ( .A(n16092), .B(n16090), .Z(n16089) );
  IV U15463 ( .A(n16087), .Z(n16092) );
  XOR U15464 ( .A(n16093), .B(n16094), .Z(n16087) );
  AND U15465 ( .A(n1872), .B(n16086), .Z(n16094) );
  XNOR U15466 ( .A(n16084), .B(n16093), .Z(n16086) );
  XNOR U15467 ( .A(n16095), .B(n16096), .Z(n16084) );
  AND U15468 ( .A(n1876), .B(n16097), .Z(n16096) );
  XOR U15469 ( .A(p_input[1521]), .B(n16095), .Z(n16097) );
  XNOR U15470 ( .A(n16098), .B(n16099), .Z(n16095) );
  AND U15471 ( .A(n1880), .B(n16100), .Z(n16099) );
  XOR U15472 ( .A(n16101), .B(n16102), .Z(n16093) );
  AND U15473 ( .A(n1884), .B(n16103), .Z(n16102) );
  XOR U15474 ( .A(n16104), .B(n16105), .Z(n16090) );
  AND U15475 ( .A(n1888), .B(n16103), .Z(n16105) );
  XNOR U15476 ( .A(n16106), .B(n16104), .Z(n16103) );
  IV U15477 ( .A(n16101), .Z(n16106) );
  XOR U15478 ( .A(n16107), .B(n16108), .Z(n16101) );
  AND U15479 ( .A(n1891), .B(n16100), .Z(n16108) );
  XNOR U15480 ( .A(n16098), .B(n16107), .Z(n16100) );
  XNOR U15481 ( .A(n16109), .B(n16110), .Z(n16098) );
  AND U15482 ( .A(n1895), .B(n16111), .Z(n16110) );
  XOR U15483 ( .A(p_input[1537]), .B(n16109), .Z(n16111) );
  XNOR U15484 ( .A(n16112), .B(n16113), .Z(n16109) );
  AND U15485 ( .A(n1899), .B(n16114), .Z(n16113) );
  XOR U15486 ( .A(n16115), .B(n16116), .Z(n16107) );
  AND U15487 ( .A(n1903), .B(n16117), .Z(n16116) );
  XOR U15488 ( .A(n16118), .B(n16119), .Z(n16104) );
  AND U15489 ( .A(n1907), .B(n16117), .Z(n16119) );
  XNOR U15490 ( .A(n16120), .B(n16118), .Z(n16117) );
  IV U15491 ( .A(n16115), .Z(n16120) );
  XOR U15492 ( .A(n16121), .B(n16122), .Z(n16115) );
  AND U15493 ( .A(n1910), .B(n16114), .Z(n16122) );
  XNOR U15494 ( .A(n16112), .B(n16121), .Z(n16114) );
  XNOR U15495 ( .A(n16123), .B(n16124), .Z(n16112) );
  AND U15496 ( .A(n1914), .B(n16125), .Z(n16124) );
  XOR U15497 ( .A(p_input[1553]), .B(n16123), .Z(n16125) );
  XNOR U15498 ( .A(n16126), .B(n16127), .Z(n16123) );
  AND U15499 ( .A(n1918), .B(n16128), .Z(n16127) );
  XOR U15500 ( .A(n16129), .B(n16130), .Z(n16121) );
  AND U15501 ( .A(n1922), .B(n16131), .Z(n16130) );
  XOR U15502 ( .A(n16132), .B(n16133), .Z(n16118) );
  AND U15503 ( .A(n1926), .B(n16131), .Z(n16133) );
  XNOR U15504 ( .A(n16134), .B(n16132), .Z(n16131) );
  IV U15505 ( .A(n16129), .Z(n16134) );
  XOR U15506 ( .A(n16135), .B(n16136), .Z(n16129) );
  AND U15507 ( .A(n1929), .B(n16128), .Z(n16136) );
  XNOR U15508 ( .A(n16126), .B(n16135), .Z(n16128) );
  XNOR U15509 ( .A(n16137), .B(n16138), .Z(n16126) );
  AND U15510 ( .A(n1933), .B(n16139), .Z(n16138) );
  XOR U15511 ( .A(p_input[1569]), .B(n16137), .Z(n16139) );
  XNOR U15512 ( .A(n16140), .B(n16141), .Z(n16137) );
  AND U15513 ( .A(n1937), .B(n16142), .Z(n16141) );
  XOR U15514 ( .A(n16143), .B(n16144), .Z(n16135) );
  AND U15515 ( .A(n1941), .B(n16145), .Z(n16144) );
  XOR U15516 ( .A(n16146), .B(n16147), .Z(n16132) );
  AND U15517 ( .A(n1945), .B(n16145), .Z(n16147) );
  XNOR U15518 ( .A(n16148), .B(n16146), .Z(n16145) );
  IV U15519 ( .A(n16143), .Z(n16148) );
  XOR U15520 ( .A(n16149), .B(n16150), .Z(n16143) );
  AND U15521 ( .A(n1948), .B(n16142), .Z(n16150) );
  XNOR U15522 ( .A(n16140), .B(n16149), .Z(n16142) );
  XNOR U15523 ( .A(n16151), .B(n16152), .Z(n16140) );
  AND U15524 ( .A(n1952), .B(n16153), .Z(n16152) );
  XOR U15525 ( .A(p_input[1585]), .B(n16151), .Z(n16153) );
  XNOR U15526 ( .A(n16154), .B(n16155), .Z(n16151) );
  AND U15527 ( .A(n1956), .B(n16156), .Z(n16155) );
  XOR U15528 ( .A(n16157), .B(n16158), .Z(n16149) );
  AND U15529 ( .A(n1960), .B(n16159), .Z(n16158) );
  XOR U15530 ( .A(n16160), .B(n16161), .Z(n16146) );
  AND U15531 ( .A(n1964), .B(n16159), .Z(n16161) );
  XNOR U15532 ( .A(n16162), .B(n16160), .Z(n16159) );
  IV U15533 ( .A(n16157), .Z(n16162) );
  XOR U15534 ( .A(n16163), .B(n16164), .Z(n16157) );
  AND U15535 ( .A(n1967), .B(n16156), .Z(n16164) );
  XNOR U15536 ( .A(n16154), .B(n16163), .Z(n16156) );
  XNOR U15537 ( .A(n16165), .B(n16166), .Z(n16154) );
  AND U15538 ( .A(n1971), .B(n16167), .Z(n16166) );
  XOR U15539 ( .A(p_input[1601]), .B(n16165), .Z(n16167) );
  XNOR U15540 ( .A(n16168), .B(n16169), .Z(n16165) );
  AND U15541 ( .A(n1975), .B(n16170), .Z(n16169) );
  XOR U15542 ( .A(n16171), .B(n16172), .Z(n16163) );
  AND U15543 ( .A(n1979), .B(n16173), .Z(n16172) );
  XOR U15544 ( .A(n16174), .B(n16175), .Z(n16160) );
  AND U15545 ( .A(n1983), .B(n16173), .Z(n16175) );
  XNOR U15546 ( .A(n16176), .B(n16174), .Z(n16173) );
  IV U15547 ( .A(n16171), .Z(n16176) );
  XOR U15548 ( .A(n16177), .B(n16178), .Z(n16171) );
  AND U15549 ( .A(n1986), .B(n16170), .Z(n16178) );
  XNOR U15550 ( .A(n16168), .B(n16177), .Z(n16170) );
  XNOR U15551 ( .A(n16179), .B(n16180), .Z(n16168) );
  AND U15552 ( .A(n1990), .B(n16181), .Z(n16180) );
  XOR U15553 ( .A(p_input[1617]), .B(n16179), .Z(n16181) );
  XNOR U15554 ( .A(n16182), .B(n16183), .Z(n16179) );
  AND U15555 ( .A(n1994), .B(n16184), .Z(n16183) );
  XOR U15556 ( .A(n16185), .B(n16186), .Z(n16177) );
  AND U15557 ( .A(n1998), .B(n16187), .Z(n16186) );
  XOR U15558 ( .A(n16188), .B(n16189), .Z(n16174) );
  AND U15559 ( .A(n2002), .B(n16187), .Z(n16189) );
  XNOR U15560 ( .A(n16190), .B(n16188), .Z(n16187) );
  IV U15561 ( .A(n16185), .Z(n16190) );
  XOR U15562 ( .A(n16191), .B(n16192), .Z(n16185) );
  AND U15563 ( .A(n2005), .B(n16184), .Z(n16192) );
  XNOR U15564 ( .A(n16182), .B(n16191), .Z(n16184) );
  XNOR U15565 ( .A(n16193), .B(n16194), .Z(n16182) );
  AND U15566 ( .A(n2009), .B(n16195), .Z(n16194) );
  XOR U15567 ( .A(p_input[1633]), .B(n16193), .Z(n16195) );
  XNOR U15568 ( .A(n16196), .B(n16197), .Z(n16193) );
  AND U15569 ( .A(n2013), .B(n16198), .Z(n16197) );
  XOR U15570 ( .A(n16199), .B(n16200), .Z(n16191) );
  AND U15571 ( .A(n2017), .B(n16201), .Z(n16200) );
  XOR U15572 ( .A(n16202), .B(n16203), .Z(n16188) );
  AND U15573 ( .A(n2021), .B(n16201), .Z(n16203) );
  XNOR U15574 ( .A(n16204), .B(n16202), .Z(n16201) );
  IV U15575 ( .A(n16199), .Z(n16204) );
  XOR U15576 ( .A(n16205), .B(n16206), .Z(n16199) );
  AND U15577 ( .A(n2024), .B(n16198), .Z(n16206) );
  XNOR U15578 ( .A(n16196), .B(n16205), .Z(n16198) );
  XNOR U15579 ( .A(n16207), .B(n16208), .Z(n16196) );
  AND U15580 ( .A(n2028), .B(n16209), .Z(n16208) );
  XOR U15581 ( .A(p_input[1649]), .B(n16207), .Z(n16209) );
  XNOR U15582 ( .A(n16210), .B(n16211), .Z(n16207) );
  AND U15583 ( .A(n2032), .B(n16212), .Z(n16211) );
  XOR U15584 ( .A(n16213), .B(n16214), .Z(n16205) );
  AND U15585 ( .A(n2036), .B(n16215), .Z(n16214) );
  XOR U15586 ( .A(n16216), .B(n16217), .Z(n16202) );
  AND U15587 ( .A(n2040), .B(n16215), .Z(n16217) );
  XNOR U15588 ( .A(n16218), .B(n16216), .Z(n16215) );
  IV U15589 ( .A(n16213), .Z(n16218) );
  XOR U15590 ( .A(n16219), .B(n16220), .Z(n16213) );
  AND U15591 ( .A(n2043), .B(n16212), .Z(n16220) );
  XNOR U15592 ( .A(n16210), .B(n16219), .Z(n16212) );
  XNOR U15593 ( .A(n16221), .B(n16222), .Z(n16210) );
  AND U15594 ( .A(n2047), .B(n16223), .Z(n16222) );
  XOR U15595 ( .A(p_input[1665]), .B(n16221), .Z(n16223) );
  XNOR U15596 ( .A(n16224), .B(n16225), .Z(n16221) );
  AND U15597 ( .A(n2051), .B(n16226), .Z(n16225) );
  XOR U15598 ( .A(n16227), .B(n16228), .Z(n16219) );
  AND U15599 ( .A(n2055), .B(n16229), .Z(n16228) );
  XOR U15600 ( .A(n16230), .B(n16231), .Z(n16216) );
  AND U15601 ( .A(n2059), .B(n16229), .Z(n16231) );
  XNOR U15602 ( .A(n16232), .B(n16230), .Z(n16229) );
  IV U15603 ( .A(n16227), .Z(n16232) );
  XOR U15604 ( .A(n16233), .B(n16234), .Z(n16227) );
  AND U15605 ( .A(n2062), .B(n16226), .Z(n16234) );
  XNOR U15606 ( .A(n16224), .B(n16233), .Z(n16226) );
  XNOR U15607 ( .A(n16235), .B(n16236), .Z(n16224) );
  AND U15608 ( .A(n2066), .B(n16237), .Z(n16236) );
  XOR U15609 ( .A(p_input[1681]), .B(n16235), .Z(n16237) );
  XNOR U15610 ( .A(n16238), .B(n16239), .Z(n16235) );
  AND U15611 ( .A(n2070), .B(n16240), .Z(n16239) );
  XOR U15612 ( .A(n16241), .B(n16242), .Z(n16233) );
  AND U15613 ( .A(n2074), .B(n16243), .Z(n16242) );
  XOR U15614 ( .A(n16244), .B(n16245), .Z(n16230) );
  AND U15615 ( .A(n2078), .B(n16243), .Z(n16245) );
  XNOR U15616 ( .A(n16246), .B(n16244), .Z(n16243) );
  IV U15617 ( .A(n16241), .Z(n16246) );
  XOR U15618 ( .A(n16247), .B(n16248), .Z(n16241) );
  AND U15619 ( .A(n2081), .B(n16240), .Z(n16248) );
  XNOR U15620 ( .A(n16238), .B(n16247), .Z(n16240) );
  XNOR U15621 ( .A(n16249), .B(n16250), .Z(n16238) );
  AND U15622 ( .A(n2085), .B(n16251), .Z(n16250) );
  XOR U15623 ( .A(p_input[1697]), .B(n16249), .Z(n16251) );
  XNOR U15624 ( .A(n16252), .B(n16253), .Z(n16249) );
  AND U15625 ( .A(n2089), .B(n16254), .Z(n16253) );
  XOR U15626 ( .A(n16255), .B(n16256), .Z(n16247) );
  AND U15627 ( .A(n2093), .B(n16257), .Z(n16256) );
  XOR U15628 ( .A(n16258), .B(n16259), .Z(n16244) );
  AND U15629 ( .A(n2097), .B(n16257), .Z(n16259) );
  XNOR U15630 ( .A(n16260), .B(n16258), .Z(n16257) );
  IV U15631 ( .A(n16255), .Z(n16260) );
  XOR U15632 ( .A(n16261), .B(n16262), .Z(n16255) );
  AND U15633 ( .A(n2100), .B(n16254), .Z(n16262) );
  XNOR U15634 ( .A(n16252), .B(n16261), .Z(n16254) );
  XNOR U15635 ( .A(n16263), .B(n16264), .Z(n16252) );
  AND U15636 ( .A(n2104), .B(n16265), .Z(n16264) );
  XOR U15637 ( .A(p_input[1713]), .B(n16263), .Z(n16265) );
  XNOR U15638 ( .A(n16266), .B(n16267), .Z(n16263) );
  AND U15639 ( .A(n2108), .B(n16268), .Z(n16267) );
  XOR U15640 ( .A(n16269), .B(n16270), .Z(n16261) );
  AND U15641 ( .A(n2112), .B(n16271), .Z(n16270) );
  XOR U15642 ( .A(n16272), .B(n16273), .Z(n16258) );
  AND U15643 ( .A(n2116), .B(n16271), .Z(n16273) );
  XNOR U15644 ( .A(n16274), .B(n16272), .Z(n16271) );
  IV U15645 ( .A(n16269), .Z(n16274) );
  XOR U15646 ( .A(n16275), .B(n16276), .Z(n16269) );
  AND U15647 ( .A(n2119), .B(n16268), .Z(n16276) );
  XNOR U15648 ( .A(n16266), .B(n16275), .Z(n16268) );
  XNOR U15649 ( .A(n16277), .B(n16278), .Z(n16266) );
  AND U15650 ( .A(n2123), .B(n16279), .Z(n16278) );
  XOR U15651 ( .A(p_input[1729]), .B(n16277), .Z(n16279) );
  XNOR U15652 ( .A(n16280), .B(n16281), .Z(n16277) );
  AND U15653 ( .A(n2127), .B(n16282), .Z(n16281) );
  XOR U15654 ( .A(n16283), .B(n16284), .Z(n16275) );
  AND U15655 ( .A(n2131), .B(n16285), .Z(n16284) );
  XOR U15656 ( .A(n16286), .B(n16287), .Z(n16272) );
  AND U15657 ( .A(n2135), .B(n16285), .Z(n16287) );
  XNOR U15658 ( .A(n16288), .B(n16286), .Z(n16285) );
  IV U15659 ( .A(n16283), .Z(n16288) );
  XOR U15660 ( .A(n16289), .B(n16290), .Z(n16283) );
  AND U15661 ( .A(n2138), .B(n16282), .Z(n16290) );
  XNOR U15662 ( .A(n16280), .B(n16289), .Z(n16282) );
  XNOR U15663 ( .A(n16291), .B(n16292), .Z(n16280) );
  AND U15664 ( .A(n2142), .B(n16293), .Z(n16292) );
  XOR U15665 ( .A(p_input[1745]), .B(n16291), .Z(n16293) );
  XNOR U15666 ( .A(n16294), .B(n16295), .Z(n16291) );
  AND U15667 ( .A(n2146), .B(n16296), .Z(n16295) );
  XOR U15668 ( .A(n16297), .B(n16298), .Z(n16289) );
  AND U15669 ( .A(n2150), .B(n16299), .Z(n16298) );
  XOR U15670 ( .A(n16300), .B(n16301), .Z(n16286) );
  AND U15671 ( .A(n2154), .B(n16299), .Z(n16301) );
  XNOR U15672 ( .A(n16302), .B(n16300), .Z(n16299) );
  IV U15673 ( .A(n16297), .Z(n16302) );
  XOR U15674 ( .A(n16303), .B(n16304), .Z(n16297) );
  AND U15675 ( .A(n2157), .B(n16296), .Z(n16304) );
  XNOR U15676 ( .A(n16294), .B(n16303), .Z(n16296) );
  XNOR U15677 ( .A(n16305), .B(n16306), .Z(n16294) );
  AND U15678 ( .A(n2161), .B(n16307), .Z(n16306) );
  XOR U15679 ( .A(p_input[1761]), .B(n16305), .Z(n16307) );
  XNOR U15680 ( .A(n16308), .B(n16309), .Z(n16305) );
  AND U15681 ( .A(n2165), .B(n16310), .Z(n16309) );
  XOR U15682 ( .A(n16311), .B(n16312), .Z(n16303) );
  AND U15683 ( .A(n2169), .B(n16313), .Z(n16312) );
  XOR U15684 ( .A(n16314), .B(n16315), .Z(n16300) );
  AND U15685 ( .A(n2173), .B(n16313), .Z(n16315) );
  XNOR U15686 ( .A(n16316), .B(n16314), .Z(n16313) );
  IV U15687 ( .A(n16311), .Z(n16316) );
  XOR U15688 ( .A(n16317), .B(n16318), .Z(n16311) );
  AND U15689 ( .A(n2176), .B(n16310), .Z(n16318) );
  XNOR U15690 ( .A(n16308), .B(n16317), .Z(n16310) );
  XNOR U15691 ( .A(n16319), .B(n16320), .Z(n16308) );
  AND U15692 ( .A(n2180), .B(n16321), .Z(n16320) );
  XOR U15693 ( .A(p_input[1777]), .B(n16319), .Z(n16321) );
  XNOR U15694 ( .A(n16322), .B(n16323), .Z(n16319) );
  AND U15695 ( .A(n2184), .B(n16324), .Z(n16323) );
  XOR U15696 ( .A(n16325), .B(n16326), .Z(n16317) );
  AND U15697 ( .A(n2188), .B(n16327), .Z(n16326) );
  XOR U15698 ( .A(n16328), .B(n16329), .Z(n16314) );
  AND U15699 ( .A(n2192), .B(n16327), .Z(n16329) );
  XNOR U15700 ( .A(n16330), .B(n16328), .Z(n16327) );
  IV U15701 ( .A(n16325), .Z(n16330) );
  XOR U15702 ( .A(n16331), .B(n16332), .Z(n16325) );
  AND U15703 ( .A(n2195), .B(n16324), .Z(n16332) );
  XNOR U15704 ( .A(n16322), .B(n16331), .Z(n16324) );
  XNOR U15705 ( .A(n16333), .B(n16334), .Z(n16322) );
  AND U15706 ( .A(n2199), .B(n16335), .Z(n16334) );
  XOR U15707 ( .A(p_input[1793]), .B(n16333), .Z(n16335) );
  XNOR U15708 ( .A(n16336), .B(n16337), .Z(n16333) );
  AND U15709 ( .A(n2203), .B(n16338), .Z(n16337) );
  XOR U15710 ( .A(n16339), .B(n16340), .Z(n16331) );
  AND U15711 ( .A(n2207), .B(n16341), .Z(n16340) );
  XOR U15712 ( .A(n16342), .B(n16343), .Z(n16328) );
  AND U15713 ( .A(n2211), .B(n16341), .Z(n16343) );
  XNOR U15714 ( .A(n16344), .B(n16342), .Z(n16341) );
  IV U15715 ( .A(n16339), .Z(n16344) );
  XOR U15716 ( .A(n16345), .B(n16346), .Z(n16339) );
  AND U15717 ( .A(n2214), .B(n16338), .Z(n16346) );
  XNOR U15718 ( .A(n16336), .B(n16345), .Z(n16338) );
  XNOR U15719 ( .A(n16347), .B(n16348), .Z(n16336) );
  AND U15720 ( .A(n2218), .B(n16349), .Z(n16348) );
  XOR U15721 ( .A(p_input[1809]), .B(n16347), .Z(n16349) );
  XNOR U15722 ( .A(n16350), .B(n16351), .Z(n16347) );
  AND U15723 ( .A(n2222), .B(n16352), .Z(n16351) );
  XOR U15724 ( .A(n16353), .B(n16354), .Z(n16345) );
  AND U15725 ( .A(n2226), .B(n16355), .Z(n16354) );
  XOR U15726 ( .A(n16356), .B(n16357), .Z(n16342) );
  AND U15727 ( .A(n2230), .B(n16355), .Z(n16357) );
  XNOR U15728 ( .A(n16358), .B(n16356), .Z(n16355) );
  IV U15729 ( .A(n16353), .Z(n16358) );
  XOR U15730 ( .A(n16359), .B(n16360), .Z(n16353) );
  AND U15731 ( .A(n2233), .B(n16352), .Z(n16360) );
  XNOR U15732 ( .A(n16350), .B(n16359), .Z(n16352) );
  XNOR U15733 ( .A(n16361), .B(n16362), .Z(n16350) );
  AND U15734 ( .A(n2237), .B(n16363), .Z(n16362) );
  XOR U15735 ( .A(p_input[1825]), .B(n16361), .Z(n16363) );
  XNOR U15736 ( .A(n16364), .B(n16365), .Z(n16361) );
  AND U15737 ( .A(n2241), .B(n16366), .Z(n16365) );
  XOR U15738 ( .A(n16367), .B(n16368), .Z(n16359) );
  AND U15739 ( .A(n2245), .B(n16369), .Z(n16368) );
  XOR U15740 ( .A(n16370), .B(n16371), .Z(n16356) );
  AND U15741 ( .A(n2249), .B(n16369), .Z(n16371) );
  XNOR U15742 ( .A(n16372), .B(n16370), .Z(n16369) );
  IV U15743 ( .A(n16367), .Z(n16372) );
  XOR U15744 ( .A(n16373), .B(n16374), .Z(n16367) );
  AND U15745 ( .A(n2252), .B(n16366), .Z(n16374) );
  XNOR U15746 ( .A(n16364), .B(n16373), .Z(n16366) );
  XNOR U15747 ( .A(n16375), .B(n16376), .Z(n16364) );
  AND U15748 ( .A(n2256), .B(n16377), .Z(n16376) );
  XOR U15749 ( .A(p_input[1841]), .B(n16375), .Z(n16377) );
  XNOR U15750 ( .A(n16378), .B(n16379), .Z(n16375) );
  AND U15751 ( .A(n2260), .B(n16380), .Z(n16379) );
  XOR U15752 ( .A(n16381), .B(n16382), .Z(n16373) );
  AND U15753 ( .A(n2264), .B(n16383), .Z(n16382) );
  XOR U15754 ( .A(n16384), .B(n16385), .Z(n16370) );
  AND U15755 ( .A(n2268), .B(n16383), .Z(n16385) );
  XNOR U15756 ( .A(n16386), .B(n16384), .Z(n16383) );
  IV U15757 ( .A(n16381), .Z(n16386) );
  XOR U15758 ( .A(n16387), .B(n16388), .Z(n16381) );
  AND U15759 ( .A(n2271), .B(n16380), .Z(n16388) );
  XNOR U15760 ( .A(n16378), .B(n16387), .Z(n16380) );
  XNOR U15761 ( .A(n16389), .B(n16390), .Z(n16378) );
  AND U15762 ( .A(n2275), .B(n16391), .Z(n16390) );
  XOR U15763 ( .A(p_input[1857]), .B(n16389), .Z(n16391) );
  XNOR U15764 ( .A(n16392), .B(n16393), .Z(n16389) );
  AND U15765 ( .A(n2279), .B(n16394), .Z(n16393) );
  XOR U15766 ( .A(n16395), .B(n16396), .Z(n16387) );
  AND U15767 ( .A(n2283), .B(n16397), .Z(n16396) );
  XOR U15768 ( .A(n16398), .B(n16399), .Z(n16384) );
  AND U15769 ( .A(n2287), .B(n16397), .Z(n16399) );
  XNOR U15770 ( .A(n16400), .B(n16398), .Z(n16397) );
  IV U15771 ( .A(n16395), .Z(n16400) );
  XOR U15772 ( .A(n16401), .B(n16402), .Z(n16395) );
  AND U15773 ( .A(n2290), .B(n16394), .Z(n16402) );
  XNOR U15774 ( .A(n16392), .B(n16401), .Z(n16394) );
  XNOR U15775 ( .A(n16403), .B(n16404), .Z(n16392) );
  AND U15776 ( .A(n2294), .B(n16405), .Z(n16404) );
  XOR U15777 ( .A(p_input[1873]), .B(n16403), .Z(n16405) );
  XNOR U15778 ( .A(n16406), .B(n16407), .Z(n16403) );
  AND U15779 ( .A(n2298), .B(n16408), .Z(n16407) );
  XOR U15780 ( .A(n16409), .B(n16410), .Z(n16401) );
  AND U15781 ( .A(n2302), .B(n16411), .Z(n16410) );
  XOR U15782 ( .A(n16412), .B(n16413), .Z(n16398) );
  AND U15783 ( .A(n2306), .B(n16411), .Z(n16413) );
  XNOR U15784 ( .A(n16414), .B(n16412), .Z(n16411) );
  IV U15785 ( .A(n16409), .Z(n16414) );
  XOR U15786 ( .A(n16415), .B(n16416), .Z(n16409) );
  AND U15787 ( .A(n2309), .B(n16408), .Z(n16416) );
  XNOR U15788 ( .A(n16406), .B(n16415), .Z(n16408) );
  XNOR U15789 ( .A(n16417), .B(n16418), .Z(n16406) );
  AND U15790 ( .A(n2313), .B(n16419), .Z(n16418) );
  XOR U15791 ( .A(p_input[1889]), .B(n16417), .Z(n16419) );
  XNOR U15792 ( .A(n16420), .B(n16421), .Z(n16417) );
  AND U15793 ( .A(n2317), .B(n16422), .Z(n16421) );
  XOR U15794 ( .A(n16423), .B(n16424), .Z(n16415) );
  AND U15795 ( .A(n2321), .B(n16425), .Z(n16424) );
  XOR U15796 ( .A(n16426), .B(n16427), .Z(n16412) );
  AND U15797 ( .A(n2325), .B(n16425), .Z(n16427) );
  XNOR U15798 ( .A(n16428), .B(n16426), .Z(n16425) );
  IV U15799 ( .A(n16423), .Z(n16428) );
  XOR U15800 ( .A(n16429), .B(n16430), .Z(n16423) );
  AND U15801 ( .A(n2328), .B(n16422), .Z(n16430) );
  XNOR U15802 ( .A(n16420), .B(n16429), .Z(n16422) );
  XNOR U15803 ( .A(n16431), .B(n16432), .Z(n16420) );
  AND U15804 ( .A(n2332), .B(n16433), .Z(n16432) );
  XOR U15805 ( .A(p_input[1905]), .B(n16431), .Z(n16433) );
  XNOR U15806 ( .A(n16434), .B(n16435), .Z(n16431) );
  AND U15807 ( .A(n2336), .B(n16436), .Z(n16435) );
  XOR U15808 ( .A(n16437), .B(n16438), .Z(n16429) );
  AND U15809 ( .A(n2340), .B(n16439), .Z(n16438) );
  XOR U15810 ( .A(n16440), .B(n16441), .Z(n16426) );
  AND U15811 ( .A(n2344), .B(n16439), .Z(n16441) );
  XNOR U15812 ( .A(n16442), .B(n16440), .Z(n16439) );
  IV U15813 ( .A(n16437), .Z(n16442) );
  XOR U15814 ( .A(n16443), .B(n16444), .Z(n16437) );
  AND U15815 ( .A(n2347), .B(n16436), .Z(n16444) );
  XNOR U15816 ( .A(n16434), .B(n16443), .Z(n16436) );
  XNOR U15817 ( .A(n16445), .B(n16446), .Z(n16434) );
  AND U15818 ( .A(n2351), .B(n16447), .Z(n16446) );
  XOR U15819 ( .A(p_input[1921]), .B(n16445), .Z(n16447) );
  XNOR U15820 ( .A(n16448), .B(n16449), .Z(n16445) );
  AND U15821 ( .A(n2355), .B(n16450), .Z(n16449) );
  XOR U15822 ( .A(n16451), .B(n16452), .Z(n16443) );
  AND U15823 ( .A(n2359), .B(n16453), .Z(n16452) );
  XOR U15824 ( .A(n16454), .B(n16455), .Z(n16440) );
  AND U15825 ( .A(n2363), .B(n16453), .Z(n16455) );
  XNOR U15826 ( .A(n16456), .B(n16454), .Z(n16453) );
  IV U15827 ( .A(n16451), .Z(n16456) );
  XOR U15828 ( .A(n16457), .B(n16458), .Z(n16451) );
  AND U15829 ( .A(n2366), .B(n16450), .Z(n16458) );
  XNOR U15830 ( .A(n16448), .B(n16457), .Z(n16450) );
  XNOR U15831 ( .A(n16459), .B(n16460), .Z(n16448) );
  AND U15832 ( .A(n2370), .B(n16461), .Z(n16460) );
  XOR U15833 ( .A(p_input[1937]), .B(n16459), .Z(n16461) );
  XNOR U15834 ( .A(n16462), .B(n16463), .Z(n16459) );
  AND U15835 ( .A(n2374), .B(n16464), .Z(n16463) );
  XOR U15836 ( .A(n16465), .B(n16466), .Z(n16457) );
  AND U15837 ( .A(n2378), .B(n16467), .Z(n16466) );
  XOR U15838 ( .A(n16468), .B(n16469), .Z(n16454) );
  AND U15839 ( .A(n2382), .B(n16467), .Z(n16469) );
  XNOR U15840 ( .A(n16470), .B(n16468), .Z(n16467) );
  IV U15841 ( .A(n16465), .Z(n16470) );
  XOR U15842 ( .A(n16471), .B(n16472), .Z(n16465) );
  AND U15843 ( .A(n2385), .B(n16464), .Z(n16472) );
  XNOR U15844 ( .A(n16462), .B(n16471), .Z(n16464) );
  XNOR U15845 ( .A(n16473), .B(n16474), .Z(n16462) );
  AND U15846 ( .A(n2389), .B(n16475), .Z(n16474) );
  XOR U15847 ( .A(p_input[1953]), .B(n16473), .Z(n16475) );
  XNOR U15848 ( .A(n16476), .B(n16477), .Z(n16473) );
  AND U15849 ( .A(n2393), .B(n16478), .Z(n16477) );
  XOR U15850 ( .A(n16479), .B(n16480), .Z(n16471) );
  AND U15851 ( .A(n2397), .B(n16481), .Z(n16480) );
  XOR U15852 ( .A(n16482), .B(n16483), .Z(n16468) );
  AND U15853 ( .A(n2401), .B(n16481), .Z(n16483) );
  XNOR U15854 ( .A(n16484), .B(n16482), .Z(n16481) );
  IV U15855 ( .A(n16479), .Z(n16484) );
  XOR U15856 ( .A(n16485), .B(n16486), .Z(n16479) );
  AND U15857 ( .A(n2404), .B(n16478), .Z(n16486) );
  XNOR U15858 ( .A(n16476), .B(n16485), .Z(n16478) );
  XNOR U15859 ( .A(n16487), .B(n16488), .Z(n16476) );
  AND U15860 ( .A(n2408), .B(n16489), .Z(n16488) );
  XOR U15861 ( .A(p_input[1969]), .B(n16487), .Z(n16489) );
  XNOR U15862 ( .A(n16490), .B(n16491), .Z(n16487) );
  AND U15863 ( .A(n2412), .B(n16492), .Z(n16491) );
  XOR U15864 ( .A(n16493), .B(n16494), .Z(n16485) );
  AND U15865 ( .A(n2416), .B(n16495), .Z(n16494) );
  XOR U15866 ( .A(n16496), .B(n16497), .Z(n16482) );
  AND U15867 ( .A(n2420), .B(n16495), .Z(n16497) );
  XNOR U15868 ( .A(n16498), .B(n16496), .Z(n16495) );
  IV U15869 ( .A(n16493), .Z(n16498) );
  XOR U15870 ( .A(n16499), .B(n16500), .Z(n16493) );
  AND U15871 ( .A(n2423), .B(n16492), .Z(n16500) );
  XNOR U15872 ( .A(n16490), .B(n16499), .Z(n16492) );
  XNOR U15873 ( .A(n16501), .B(n16502), .Z(n16490) );
  AND U15874 ( .A(n2427), .B(n16503), .Z(n16502) );
  XOR U15875 ( .A(p_input[1985]), .B(n16501), .Z(n16503) );
  XOR U15876 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n16504), 
        .Z(n16501) );
  AND U15877 ( .A(n2430), .B(n16505), .Z(n16504) );
  XOR U15878 ( .A(n16506), .B(n16507), .Z(n16499) );
  AND U15879 ( .A(n2434), .B(n16508), .Z(n16507) );
  XOR U15880 ( .A(n16509), .B(n16510), .Z(n16496) );
  AND U15881 ( .A(n2438), .B(n16508), .Z(n16510) );
  XNOR U15882 ( .A(n16511), .B(n16509), .Z(n16508) );
  IV U15883 ( .A(n16506), .Z(n16511) );
  XOR U15884 ( .A(n16512), .B(n16513), .Z(n16506) );
  AND U15885 ( .A(n2441), .B(n16505), .Z(n16513) );
  XOR U15886 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n16512), 
        .Z(n16505) );
  XOR U15887 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n16514), 
        .Z(n16512) );
  AND U15888 ( .A(n2443), .B(n16515), .Z(n16514) );
  XOR U15889 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n16516), .Z(n16509) );
  AND U15890 ( .A(n2446), .B(n16515), .Z(n16516) );
  XOR U15891 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n16515) );
  XOR U15892 ( .A(n16517), .B(n16518), .Z(o[16]) );
  XOR U15893 ( .A(n47), .B(n16519), .Z(o[15]) );
  AND U15894 ( .A(n62), .B(n16520), .Z(n47) );
  XOR U15895 ( .A(n48), .B(n16519), .Z(n16520) );
  XOR U15896 ( .A(n16521), .B(n16522), .Z(n16519) );
  AND U15897 ( .A(n82), .B(n16523), .Z(n16522) );
  XOR U15898 ( .A(n16524), .B(n13), .Z(n48) );
  AND U15899 ( .A(n65), .B(n16525), .Z(n13) );
  XOR U15900 ( .A(n14), .B(n16524), .Z(n16525) );
  XOR U15901 ( .A(n16526), .B(n16527), .Z(n14) );
  AND U15902 ( .A(n70), .B(n16528), .Z(n16527) );
  XOR U15903 ( .A(p_input[15]), .B(n16526), .Z(n16528) );
  XNOR U15904 ( .A(n16529), .B(n16530), .Z(n16526) );
  AND U15905 ( .A(n74), .B(n16531), .Z(n16530) );
  XOR U15906 ( .A(n16532), .B(n16533), .Z(n16524) );
  AND U15907 ( .A(n78), .B(n16523), .Z(n16533) );
  XNOR U15908 ( .A(n16534), .B(n16521), .Z(n16523) );
  XOR U15909 ( .A(n16535), .B(n16536), .Z(n16521) );
  AND U15910 ( .A(n102), .B(n16537), .Z(n16536) );
  IV U15911 ( .A(n16532), .Z(n16534) );
  XOR U15912 ( .A(n16538), .B(n16539), .Z(n16532) );
  AND U15913 ( .A(n86), .B(n16531), .Z(n16539) );
  XNOR U15914 ( .A(n16529), .B(n16538), .Z(n16531) );
  XNOR U15915 ( .A(n16540), .B(n16541), .Z(n16529) );
  AND U15916 ( .A(n90), .B(n16542), .Z(n16541) );
  XOR U15917 ( .A(p_input[31]), .B(n16540), .Z(n16542) );
  XNOR U15918 ( .A(n16543), .B(n16544), .Z(n16540) );
  AND U15919 ( .A(n94), .B(n16545), .Z(n16544) );
  XOR U15920 ( .A(n16546), .B(n16547), .Z(n16538) );
  AND U15921 ( .A(n98), .B(n16537), .Z(n16547) );
  XNOR U15922 ( .A(n16548), .B(n16535), .Z(n16537) );
  XOR U15923 ( .A(n16549), .B(n16550), .Z(n16535) );
  AND U15924 ( .A(n121), .B(n16551), .Z(n16550) );
  IV U15925 ( .A(n16546), .Z(n16548) );
  XOR U15926 ( .A(n16552), .B(n16553), .Z(n16546) );
  AND U15927 ( .A(n105), .B(n16545), .Z(n16553) );
  XNOR U15928 ( .A(n16543), .B(n16552), .Z(n16545) );
  XNOR U15929 ( .A(n16554), .B(n16555), .Z(n16543) );
  AND U15930 ( .A(n109), .B(n16556), .Z(n16555) );
  XOR U15931 ( .A(p_input[47]), .B(n16554), .Z(n16556) );
  XNOR U15932 ( .A(n16557), .B(n16558), .Z(n16554) );
  AND U15933 ( .A(n113), .B(n16559), .Z(n16558) );
  XOR U15934 ( .A(n16560), .B(n16561), .Z(n16552) );
  AND U15935 ( .A(n117), .B(n16551), .Z(n16561) );
  XNOR U15936 ( .A(n16562), .B(n16549), .Z(n16551) );
  XOR U15937 ( .A(n16563), .B(n16564), .Z(n16549) );
  AND U15938 ( .A(n140), .B(n16565), .Z(n16564) );
  IV U15939 ( .A(n16560), .Z(n16562) );
  XOR U15940 ( .A(n16566), .B(n16567), .Z(n16560) );
  AND U15941 ( .A(n124), .B(n16559), .Z(n16567) );
  XNOR U15942 ( .A(n16557), .B(n16566), .Z(n16559) );
  XNOR U15943 ( .A(n16568), .B(n16569), .Z(n16557) );
  AND U15944 ( .A(n128), .B(n16570), .Z(n16569) );
  XOR U15945 ( .A(p_input[63]), .B(n16568), .Z(n16570) );
  XNOR U15946 ( .A(n16571), .B(n16572), .Z(n16568) );
  AND U15947 ( .A(n132), .B(n16573), .Z(n16572) );
  XOR U15948 ( .A(n16574), .B(n16575), .Z(n16566) );
  AND U15949 ( .A(n136), .B(n16565), .Z(n16575) );
  XNOR U15950 ( .A(n16576), .B(n16563), .Z(n16565) );
  XOR U15951 ( .A(n16577), .B(n16578), .Z(n16563) );
  AND U15952 ( .A(n159), .B(n16579), .Z(n16578) );
  IV U15953 ( .A(n16574), .Z(n16576) );
  XOR U15954 ( .A(n16580), .B(n16581), .Z(n16574) );
  AND U15955 ( .A(n143), .B(n16573), .Z(n16581) );
  XNOR U15956 ( .A(n16571), .B(n16580), .Z(n16573) );
  XNOR U15957 ( .A(n16582), .B(n16583), .Z(n16571) );
  AND U15958 ( .A(n147), .B(n16584), .Z(n16583) );
  XOR U15959 ( .A(p_input[79]), .B(n16582), .Z(n16584) );
  XNOR U15960 ( .A(n16585), .B(n16586), .Z(n16582) );
  AND U15961 ( .A(n151), .B(n16587), .Z(n16586) );
  XOR U15962 ( .A(n16588), .B(n16589), .Z(n16580) );
  AND U15963 ( .A(n155), .B(n16579), .Z(n16589) );
  XNOR U15964 ( .A(n16590), .B(n16577), .Z(n16579) );
  XOR U15965 ( .A(n16591), .B(n16592), .Z(n16577) );
  AND U15966 ( .A(n178), .B(n16593), .Z(n16592) );
  IV U15967 ( .A(n16588), .Z(n16590) );
  XOR U15968 ( .A(n16594), .B(n16595), .Z(n16588) );
  AND U15969 ( .A(n162), .B(n16587), .Z(n16595) );
  XNOR U15970 ( .A(n16585), .B(n16594), .Z(n16587) );
  XNOR U15971 ( .A(n16596), .B(n16597), .Z(n16585) );
  AND U15972 ( .A(n166), .B(n16598), .Z(n16597) );
  XOR U15973 ( .A(p_input[95]), .B(n16596), .Z(n16598) );
  XNOR U15974 ( .A(n16599), .B(n16600), .Z(n16596) );
  AND U15975 ( .A(n170), .B(n16601), .Z(n16600) );
  XOR U15976 ( .A(n16602), .B(n16603), .Z(n16594) );
  AND U15977 ( .A(n174), .B(n16593), .Z(n16603) );
  XNOR U15978 ( .A(n16604), .B(n16591), .Z(n16593) );
  XOR U15979 ( .A(n16605), .B(n16606), .Z(n16591) );
  AND U15980 ( .A(n197), .B(n16607), .Z(n16606) );
  IV U15981 ( .A(n16602), .Z(n16604) );
  XOR U15982 ( .A(n16608), .B(n16609), .Z(n16602) );
  AND U15983 ( .A(n181), .B(n16601), .Z(n16609) );
  XNOR U15984 ( .A(n16599), .B(n16608), .Z(n16601) );
  XNOR U15985 ( .A(n16610), .B(n16611), .Z(n16599) );
  AND U15986 ( .A(n185), .B(n16612), .Z(n16611) );
  XOR U15987 ( .A(p_input[111]), .B(n16610), .Z(n16612) );
  XNOR U15988 ( .A(n16613), .B(n16614), .Z(n16610) );
  AND U15989 ( .A(n189), .B(n16615), .Z(n16614) );
  XOR U15990 ( .A(n16616), .B(n16617), .Z(n16608) );
  AND U15991 ( .A(n193), .B(n16607), .Z(n16617) );
  XNOR U15992 ( .A(n16618), .B(n16605), .Z(n16607) );
  XOR U15993 ( .A(n16619), .B(n16620), .Z(n16605) );
  AND U15994 ( .A(n216), .B(n16621), .Z(n16620) );
  IV U15995 ( .A(n16616), .Z(n16618) );
  XOR U15996 ( .A(n16622), .B(n16623), .Z(n16616) );
  AND U15997 ( .A(n200), .B(n16615), .Z(n16623) );
  XNOR U15998 ( .A(n16613), .B(n16622), .Z(n16615) );
  XNOR U15999 ( .A(n16624), .B(n16625), .Z(n16613) );
  AND U16000 ( .A(n204), .B(n16626), .Z(n16625) );
  XOR U16001 ( .A(p_input[127]), .B(n16624), .Z(n16626) );
  XNOR U16002 ( .A(n16627), .B(n16628), .Z(n16624) );
  AND U16003 ( .A(n208), .B(n16629), .Z(n16628) );
  XOR U16004 ( .A(n16630), .B(n16631), .Z(n16622) );
  AND U16005 ( .A(n212), .B(n16621), .Z(n16631) );
  XNOR U16006 ( .A(n16632), .B(n16619), .Z(n16621) );
  XOR U16007 ( .A(n16633), .B(n16634), .Z(n16619) );
  AND U16008 ( .A(n235), .B(n16635), .Z(n16634) );
  IV U16009 ( .A(n16630), .Z(n16632) );
  XOR U16010 ( .A(n16636), .B(n16637), .Z(n16630) );
  AND U16011 ( .A(n219), .B(n16629), .Z(n16637) );
  XNOR U16012 ( .A(n16627), .B(n16636), .Z(n16629) );
  XNOR U16013 ( .A(n16638), .B(n16639), .Z(n16627) );
  AND U16014 ( .A(n223), .B(n16640), .Z(n16639) );
  XOR U16015 ( .A(p_input[143]), .B(n16638), .Z(n16640) );
  XNOR U16016 ( .A(n16641), .B(n16642), .Z(n16638) );
  AND U16017 ( .A(n227), .B(n16643), .Z(n16642) );
  XOR U16018 ( .A(n16644), .B(n16645), .Z(n16636) );
  AND U16019 ( .A(n231), .B(n16635), .Z(n16645) );
  XNOR U16020 ( .A(n16646), .B(n16633), .Z(n16635) );
  XOR U16021 ( .A(n16647), .B(n16648), .Z(n16633) );
  AND U16022 ( .A(n254), .B(n16649), .Z(n16648) );
  IV U16023 ( .A(n16644), .Z(n16646) );
  XOR U16024 ( .A(n16650), .B(n16651), .Z(n16644) );
  AND U16025 ( .A(n238), .B(n16643), .Z(n16651) );
  XNOR U16026 ( .A(n16641), .B(n16650), .Z(n16643) );
  XNOR U16027 ( .A(n16652), .B(n16653), .Z(n16641) );
  AND U16028 ( .A(n242), .B(n16654), .Z(n16653) );
  XOR U16029 ( .A(p_input[159]), .B(n16652), .Z(n16654) );
  XNOR U16030 ( .A(n16655), .B(n16656), .Z(n16652) );
  AND U16031 ( .A(n246), .B(n16657), .Z(n16656) );
  XOR U16032 ( .A(n16658), .B(n16659), .Z(n16650) );
  AND U16033 ( .A(n250), .B(n16649), .Z(n16659) );
  XNOR U16034 ( .A(n16660), .B(n16647), .Z(n16649) );
  XOR U16035 ( .A(n16661), .B(n16662), .Z(n16647) );
  AND U16036 ( .A(n273), .B(n16663), .Z(n16662) );
  IV U16037 ( .A(n16658), .Z(n16660) );
  XOR U16038 ( .A(n16664), .B(n16665), .Z(n16658) );
  AND U16039 ( .A(n257), .B(n16657), .Z(n16665) );
  XNOR U16040 ( .A(n16655), .B(n16664), .Z(n16657) );
  XNOR U16041 ( .A(n16666), .B(n16667), .Z(n16655) );
  AND U16042 ( .A(n261), .B(n16668), .Z(n16667) );
  XOR U16043 ( .A(p_input[175]), .B(n16666), .Z(n16668) );
  XNOR U16044 ( .A(n16669), .B(n16670), .Z(n16666) );
  AND U16045 ( .A(n265), .B(n16671), .Z(n16670) );
  XOR U16046 ( .A(n16672), .B(n16673), .Z(n16664) );
  AND U16047 ( .A(n269), .B(n16663), .Z(n16673) );
  XNOR U16048 ( .A(n16674), .B(n16661), .Z(n16663) );
  XOR U16049 ( .A(n16675), .B(n16676), .Z(n16661) );
  AND U16050 ( .A(n292), .B(n16677), .Z(n16676) );
  IV U16051 ( .A(n16672), .Z(n16674) );
  XOR U16052 ( .A(n16678), .B(n16679), .Z(n16672) );
  AND U16053 ( .A(n276), .B(n16671), .Z(n16679) );
  XNOR U16054 ( .A(n16669), .B(n16678), .Z(n16671) );
  XNOR U16055 ( .A(n16680), .B(n16681), .Z(n16669) );
  AND U16056 ( .A(n280), .B(n16682), .Z(n16681) );
  XOR U16057 ( .A(p_input[191]), .B(n16680), .Z(n16682) );
  XNOR U16058 ( .A(n16683), .B(n16684), .Z(n16680) );
  AND U16059 ( .A(n284), .B(n16685), .Z(n16684) );
  XOR U16060 ( .A(n16686), .B(n16687), .Z(n16678) );
  AND U16061 ( .A(n288), .B(n16677), .Z(n16687) );
  XNOR U16062 ( .A(n16688), .B(n16675), .Z(n16677) );
  XOR U16063 ( .A(n16689), .B(n16690), .Z(n16675) );
  AND U16064 ( .A(n311), .B(n16691), .Z(n16690) );
  IV U16065 ( .A(n16686), .Z(n16688) );
  XOR U16066 ( .A(n16692), .B(n16693), .Z(n16686) );
  AND U16067 ( .A(n295), .B(n16685), .Z(n16693) );
  XNOR U16068 ( .A(n16683), .B(n16692), .Z(n16685) );
  XNOR U16069 ( .A(n16694), .B(n16695), .Z(n16683) );
  AND U16070 ( .A(n299), .B(n16696), .Z(n16695) );
  XOR U16071 ( .A(p_input[207]), .B(n16694), .Z(n16696) );
  XNOR U16072 ( .A(n16697), .B(n16698), .Z(n16694) );
  AND U16073 ( .A(n303), .B(n16699), .Z(n16698) );
  XOR U16074 ( .A(n16700), .B(n16701), .Z(n16692) );
  AND U16075 ( .A(n307), .B(n16691), .Z(n16701) );
  XNOR U16076 ( .A(n16702), .B(n16689), .Z(n16691) );
  XOR U16077 ( .A(n16703), .B(n16704), .Z(n16689) );
  AND U16078 ( .A(n330), .B(n16705), .Z(n16704) );
  IV U16079 ( .A(n16700), .Z(n16702) );
  XOR U16080 ( .A(n16706), .B(n16707), .Z(n16700) );
  AND U16081 ( .A(n314), .B(n16699), .Z(n16707) );
  XNOR U16082 ( .A(n16697), .B(n16706), .Z(n16699) );
  XNOR U16083 ( .A(n16708), .B(n16709), .Z(n16697) );
  AND U16084 ( .A(n318), .B(n16710), .Z(n16709) );
  XOR U16085 ( .A(p_input[223]), .B(n16708), .Z(n16710) );
  XNOR U16086 ( .A(n16711), .B(n16712), .Z(n16708) );
  AND U16087 ( .A(n322), .B(n16713), .Z(n16712) );
  XOR U16088 ( .A(n16714), .B(n16715), .Z(n16706) );
  AND U16089 ( .A(n326), .B(n16705), .Z(n16715) );
  XNOR U16090 ( .A(n16716), .B(n16703), .Z(n16705) );
  XOR U16091 ( .A(n16717), .B(n16718), .Z(n16703) );
  AND U16092 ( .A(n349), .B(n16719), .Z(n16718) );
  IV U16093 ( .A(n16714), .Z(n16716) );
  XOR U16094 ( .A(n16720), .B(n16721), .Z(n16714) );
  AND U16095 ( .A(n333), .B(n16713), .Z(n16721) );
  XNOR U16096 ( .A(n16711), .B(n16720), .Z(n16713) );
  XNOR U16097 ( .A(n16722), .B(n16723), .Z(n16711) );
  AND U16098 ( .A(n337), .B(n16724), .Z(n16723) );
  XOR U16099 ( .A(p_input[239]), .B(n16722), .Z(n16724) );
  XNOR U16100 ( .A(n16725), .B(n16726), .Z(n16722) );
  AND U16101 ( .A(n341), .B(n16727), .Z(n16726) );
  XOR U16102 ( .A(n16728), .B(n16729), .Z(n16720) );
  AND U16103 ( .A(n345), .B(n16719), .Z(n16729) );
  XNOR U16104 ( .A(n16730), .B(n16717), .Z(n16719) );
  XOR U16105 ( .A(n16731), .B(n16732), .Z(n16717) );
  AND U16106 ( .A(n368), .B(n16733), .Z(n16732) );
  IV U16107 ( .A(n16728), .Z(n16730) );
  XOR U16108 ( .A(n16734), .B(n16735), .Z(n16728) );
  AND U16109 ( .A(n352), .B(n16727), .Z(n16735) );
  XNOR U16110 ( .A(n16725), .B(n16734), .Z(n16727) );
  XNOR U16111 ( .A(n16736), .B(n16737), .Z(n16725) );
  AND U16112 ( .A(n356), .B(n16738), .Z(n16737) );
  XOR U16113 ( .A(p_input[255]), .B(n16736), .Z(n16738) );
  XNOR U16114 ( .A(n16739), .B(n16740), .Z(n16736) );
  AND U16115 ( .A(n360), .B(n16741), .Z(n16740) );
  XOR U16116 ( .A(n16742), .B(n16743), .Z(n16734) );
  AND U16117 ( .A(n364), .B(n16733), .Z(n16743) );
  XNOR U16118 ( .A(n16744), .B(n16731), .Z(n16733) );
  XOR U16119 ( .A(n16745), .B(n16746), .Z(n16731) );
  AND U16120 ( .A(n387), .B(n16747), .Z(n16746) );
  IV U16121 ( .A(n16742), .Z(n16744) );
  XOR U16122 ( .A(n16748), .B(n16749), .Z(n16742) );
  AND U16123 ( .A(n371), .B(n16741), .Z(n16749) );
  XNOR U16124 ( .A(n16739), .B(n16748), .Z(n16741) );
  XNOR U16125 ( .A(n16750), .B(n16751), .Z(n16739) );
  AND U16126 ( .A(n375), .B(n16752), .Z(n16751) );
  XOR U16127 ( .A(p_input[271]), .B(n16750), .Z(n16752) );
  XNOR U16128 ( .A(n16753), .B(n16754), .Z(n16750) );
  AND U16129 ( .A(n379), .B(n16755), .Z(n16754) );
  XOR U16130 ( .A(n16756), .B(n16757), .Z(n16748) );
  AND U16131 ( .A(n383), .B(n16747), .Z(n16757) );
  XNOR U16132 ( .A(n16758), .B(n16745), .Z(n16747) );
  XOR U16133 ( .A(n16759), .B(n16760), .Z(n16745) );
  AND U16134 ( .A(n406), .B(n16761), .Z(n16760) );
  IV U16135 ( .A(n16756), .Z(n16758) );
  XOR U16136 ( .A(n16762), .B(n16763), .Z(n16756) );
  AND U16137 ( .A(n390), .B(n16755), .Z(n16763) );
  XNOR U16138 ( .A(n16753), .B(n16762), .Z(n16755) );
  XNOR U16139 ( .A(n16764), .B(n16765), .Z(n16753) );
  AND U16140 ( .A(n394), .B(n16766), .Z(n16765) );
  XOR U16141 ( .A(p_input[287]), .B(n16764), .Z(n16766) );
  XNOR U16142 ( .A(n16767), .B(n16768), .Z(n16764) );
  AND U16143 ( .A(n398), .B(n16769), .Z(n16768) );
  XOR U16144 ( .A(n16770), .B(n16771), .Z(n16762) );
  AND U16145 ( .A(n402), .B(n16761), .Z(n16771) );
  XNOR U16146 ( .A(n16772), .B(n16759), .Z(n16761) );
  XOR U16147 ( .A(n16773), .B(n16774), .Z(n16759) );
  AND U16148 ( .A(n425), .B(n16775), .Z(n16774) );
  IV U16149 ( .A(n16770), .Z(n16772) );
  XOR U16150 ( .A(n16776), .B(n16777), .Z(n16770) );
  AND U16151 ( .A(n409), .B(n16769), .Z(n16777) );
  XNOR U16152 ( .A(n16767), .B(n16776), .Z(n16769) );
  XNOR U16153 ( .A(n16778), .B(n16779), .Z(n16767) );
  AND U16154 ( .A(n413), .B(n16780), .Z(n16779) );
  XOR U16155 ( .A(p_input[303]), .B(n16778), .Z(n16780) );
  XNOR U16156 ( .A(n16781), .B(n16782), .Z(n16778) );
  AND U16157 ( .A(n417), .B(n16783), .Z(n16782) );
  XOR U16158 ( .A(n16784), .B(n16785), .Z(n16776) );
  AND U16159 ( .A(n421), .B(n16775), .Z(n16785) );
  XNOR U16160 ( .A(n16786), .B(n16773), .Z(n16775) );
  XOR U16161 ( .A(n16787), .B(n16788), .Z(n16773) );
  AND U16162 ( .A(n444), .B(n16789), .Z(n16788) );
  IV U16163 ( .A(n16784), .Z(n16786) );
  XOR U16164 ( .A(n16790), .B(n16791), .Z(n16784) );
  AND U16165 ( .A(n428), .B(n16783), .Z(n16791) );
  XNOR U16166 ( .A(n16781), .B(n16790), .Z(n16783) );
  XNOR U16167 ( .A(n16792), .B(n16793), .Z(n16781) );
  AND U16168 ( .A(n432), .B(n16794), .Z(n16793) );
  XOR U16169 ( .A(p_input[319]), .B(n16792), .Z(n16794) );
  XNOR U16170 ( .A(n16795), .B(n16796), .Z(n16792) );
  AND U16171 ( .A(n436), .B(n16797), .Z(n16796) );
  XOR U16172 ( .A(n16798), .B(n16799), .Z(n16790) );
  AND U16173 ( .A(n440), .B(n16789), .Z(n16799) );
  XNOR U16174 ( .A(n16800), .B(n16787), .Z(n16789) );
  XOR U16175 ( .A(n16801), .B(n16802), .Z(n16787) );
  AND U16176 ( .A(n463), .B(n16803), .Z(n16802) );
  IV U16177 ( .A(n16798), .Z(n16800) );
  XOR U16178 ( .A(n16804), .B(n16805), .Z(n16798) );
  AND U16179 ( .A(n447), .B(n16797), .Z(n16805) );
  XNOR U16180 ( .A(n16795), .B(n16804), .Z(n16797) );
  XNOR U16181 ( .A(n16806), .B(n16807), .Z(n16795) );
  AND U16182 ( .A(n451), .B(n16808), .Z(n16807) );
  XOR U16183 ( .A(p_input[335]), .B(n16806), .Z(n16808) );
  XNOR U16184 ( .A(n16809), .B(n16810), .Z(n16806) );
  AND U16185 ( .A(n455), .B(n16811), .Z(n16810) );
  XOR U16186 ( .A(n16812), .B(n16813), .Z(n16804) );
  AND U16187 ( .A(n459), .B(n16803), .Z(n16813) );
  XNOR U16188 ( .A(n16814), .B(n16801), .Z(n16803) );
  XOR U16189 ( .A(n16815), .B(n16816), .Z(n16801) );
  AND U16190 ( .A(n482), .B(n16817), .Z(n16816) );
  IV U16191 ( .A(n16812), .Z(n16814) );
  XOR U16192 ( .A(n16818), .B(n16819), .Z(n16812) );
  AND U16193 ( .A(n466), .B(n16811), .Z(n16819) );
  XNOR U16194 ( .A(n16809), .B(n16818), .Z(n16811) );
  XNOR U16195 ( .A(n16820), .B(n16821), .Z(n16809) );
  AND U16196 ( .A(n470), .B(n16822), .Z(n16821) );
  XOR U16197 ( .A(p_input[351]), .B(n16820), .Z(n16822) );
  XNOR U16198 ( .A(n16823), .B(n16824), .Z(n16820) );
  AND U16199 ( .A(n474), .B(n16825), .Z(n16824) );
  XOR U16200 ( .A(n16826), .B(n16827), .Z(n16818) );
  AND U16201 ( .A(n478), .B(n16817), .Z(n16827) );
  XNOR U16202 ( .A(n16828), .B(n16815), .Z(n16817) );
  XOR U16203 ( .A(n16829), .B(n16830), .Z(n16815) );
  AND U16204 ( .A(n501), .B(n16831), .Z(n16830) );
  IV U16205 ( .A(n16826), .Z(n16828) );
  XOR U16206 ( .A(n16832), .B(n16833), .Z(n16826) );
  AND U16207 ( .A(n485), .B(n16825), .Z(n16833) );
  XNOR U16208 ( .A(n16823), .B(n16832), .Z(n16825) );
  XNOR U16209 ( .A(n16834), .B(n16835), .Z(n16823) );
  AND U16210 ( .A(n489), .B(n16836), .Z(n16835) );
  XOR U16211 ( .A(p_input[367]), .B(n16834), .Z(n16836) );
  XNOR U16212 ( .A(n16837), .B(n16838), .Z(n16834) );
  AND U16213 ( .A(n493), .B(n16839), .Z(n16838) );
  XOR U16214 ( .A(n16840), .B(n16841), .Z(n16832) );
  AND U16215 ( .A(n497), .B(n16831), .Z(n16841) );
  XNOR U16216 ( .A(n16842), .B(n16829), .Z(n16831) );
  XOR U16217 ( .A(n16843), .B(n16844), .Z(n16829) );
  AND U16218 ( .A(n520), .B(n16845), .Z(n16844) );
  IV U16219 ( .A(n16840), .Z(n16842) );
  XOR U16220 ( .A(n16846), .B(n16847), .Z(n16840) );
  AND U16221 ( .A(n504), .B(n16839), .Z(n16847) );
  XNOR U16222 ( .A(n16837), .B(n16846), .Z(n16839) );
  XNOR U16223 ( .A(n16848), .B(n16849), .Z(n16837) );
  AND U16224 ( .A(n508), .B(n16850), .Z(n16849) );
  XOR U16225 ( .A(p_input[383]), .B(n16848), .Z(n16850) );
  XNOR U16226 ( .A(n16851), .B(n16852), .Z(n16848) );
  AND U16227 ( .A(n512), .B(n16853), .Z(n16852) );
  XOR U16228 ( .A(n16854), .B(n16855), .Z(n16846) );
  AND U16229 ( .A(n516), .B(n16845), .Z(n16855) );
  XNOR U16230 ( .A(n16856), .B(n16843), .Z(n16845) );
  XOR U16231 ( .A(n16857), .B(n16858), .Z(n16843) );
  AND U16232 ( .A(n539), .B(n16859), .Z(n16858) );
  IV U16233 ( .A(n16854), .Z(n16856) );
  XOR U16234 ( .A(n16860), .B(n16861), .Z(n16854) );
  AND U16235 ( .A(n523), .B(n16853), .Z(n16861) );
  XNOR U16236 ( .A(n16851), .B(n16860), .Z(n16853) );
  XNOR U16237 ( .A(n16862), .B(n16863), .Z(n16851) );
  AND U16238 ( .A(n527), .B(n16864), .Z(n16863) );
  XOR U16239 ( .A(p_input[399]), .B(n16862), .Z(n16864) );
  XNOR U16240 ( .A(n16865), .B(n16866), .Z(n16862) );
  AND U16241 ( .A(n531), .B(n16867), .Z(n16866) );
  XOR U16242 ( .A(n16868), .B(n16869), .Z(n16860) );
  AND U16243 ( .A(n535), .B(n16859), .Z(n16869) );
  XNOR U16244 ( .A(n16870), .B(n16857), .Z(n16859) );
  XOR U16245 ( .A(n16871), .B(n16872), .Z(n16857) );
  AND U16246 ( .A(n558), .B(n16873), .Z(n16872) );
  IV U16247 ( .A(n16868), .Z(n16870) );
  XOR U16248 ( .A(n16874), .B(n16875), .Z(n16868) );
  AND U16249 ( .A(n542), .B(n16867), .Z(n16875) );
  XNOR U16250 ( .A(n16865), .B(n16874), .Z(n16867) );
  XNOR U16251 ( .A(n16876), .B(n16877), .Z(n16865) );
  AND U16252 ( .A(n546), .B(n16878), .Z(n16877) );
  XOR U16253 ( .A(p_input[415]), .B(n16876), .Z(n16878) );
  XNOR U16254 ( .A(n16879), .B(n16880), .Z(n16876) );
  AND U16255 ( .A(n550), .B(n16881), .Z(n16880) );
  XOR U16256 ( .A(n16882), .B(n16883), .Z(n16874) );
  AND U16257 ( .A(n554), .B(n16873), .Z(n16883) );
  XNOR U16258 ( .A(n16884), .B(n16871), .Z(n16873) );
  XOR U16259 ( .A(n16885), .B(n16886), .Z(n16871) );
  AND U16260 ( .A(n577), .B(n16887), .Z(n16886) );
  IV U16261 ( .A(n16882), .Z(n16884) );
  XOR U16262 ( .A(n16888), .B(n16889), .Z(n16882) );
  AND U16263 ( .A(n561), .B(n16881), .Z(n16889) );
  XNOR U16264 ( .A(n16879), .B(n16888), .Z(n16881) );
  XNOR U16265 ( .A(n16890), .B(n16891), .Z(n16879) );
  AND U16266 ( .A(n565), .B(n16892), .Z(n16891) );
  XOR U16267 ( .A(p_input[431]), .B(n16890), .Z(n16892) );
  XNOR U16268 ( .A(n16893), .B(n16894), .Z(n16890) );
  AND U16269 ( .A(n569), .B(n16895), .Z(n16894) );
  XOR U16270 ( .A(n16896), .B(n16897), .Z(n16888) );
  AND U16271 ( .A(n573), .B(n16887), .Z(n16897) );
  XNOR U16272 ( .A(n16898), .B(n16885), .Z(n16887) );
  XOR U16273 ( .A(n16899), .B(n16900), .Z(n16885) );
  AND U16274 ( .A(n596), .B(n16901), .Z(n16900) );
  IV U16275 ( .A(n16896), .Z(n16898) );
  XOR U16276 ( .A(n16902), .B(n16903), .Z(n16896) );
  AND U16277 ( .A(n580), .B(n16895), .Z(n16903) );
  XNOR U16278 ( .A(n16893), .B(n16902), .Z(n16895) );
  XNOR U16279 ( .A(n16904), .B(n16905), .Z(n16893) );
  AND U16280 ( .A(n584), .B(n16906), .Z(n16905) );
  XOR U16281 ( .A(p_input[447]), .B(n16904), .Z(n16906) );
  XNOR U16282 ( .A(n16907), .B(n16908), .Z(n16904) );
  AND U16283 ( .A(n588), .B(n16909), .Z(n16908) );
  XOR U16284 ( .A(n16910), .B(n16911), .Z(n16902) );
  AND U16285 ( .A(n592), .B(n16901), .Z(n16911) );
  XNOR U16286 ( .A(n16912), .B(n16899), .Z(n16901) );
  XOR U16287 ( .A(n16913), .B(n16914), .Z(n16899) );
  AND U16288 ( .A(n615), .B(n16915), .Z(n16914) );
  IV U16289 ( .A(n16910), .Z(n16912) );
  XOR U16290 ( .A(n16916), .B(n16917), .Z(n16910) );
  AND U16291 ( .A(n599), .B(n16909), .Z(n16917) );
  XNOR U16292 ( .A(n16907), .B(n16916), .Z(n16909) );
  XNOR U16293 ( .A(n16918), .B(n16919), .Z(n16907) );
  AND U16294 ( .A(n603), .B(n16920), .Z(n16919) );
  XOR U16295 ( .A(p_input[463]), .B(n16918), .Z(n16920) );
  XNOR U16296 ( .A(n16921), .B(n16922), .Z(n16918) );
  AND U16297 ( .A(n607), .B(n16923), .Z(n16922) );
  XOR U16298 ( .A(n16924), .B(n16925), .Z(n16916) );
  AND U16299 ( .A(n611), .B(n16915), .Z(n16925) );
  XNOR U16300 ( .A(n16926), .B(n16913), .Z(n16915) );
  XOR U16301 ( .A(n16927), .B(n16928), .Z(n16913) );
  AND U16302 ( .A(n634), .B(n16929), .Z(n16928) );
  IV U16303 ( .A(n16924), .Z(n16926) );
  XOR U16304 ( .A(n16930), .B(n16931), .Z(n16924) );
  AND U16305 ( .A(n618), .B(n16923), .Z(n16931) );
  XNOR U16306 ( .A(n16921), .B(n16930), .Z(n16923) );
  XNOR U16307 ( .A(n16932), .B(n16933), .Z(n16921) );
  AND U16308 ( .A(n622), .B(n16934), .Z(n16933) );
  XOR U16309 ( .A(p_input[479]), .B(n16932), .Z(n16934) );
  XNOR U16310 ( .A(n16935), .B(n16936), .Z(n16932) );
  AND U16311 ( .A(n626), .B(n16937), .Z(n16936) );
  XOR U16312 ( .A(n16938), .B(n16939), .Z(n16930) );
  AND U16313 ( .A(n630), .B(n16929), .Z(n16939) );
  XNOR U16314 ( .A(n16940), .B(n16927), .Z(n16929) );
  XOR U16315 ( .A(n16941), .B(n16942), .Z(n16927) );
  AND U16316 ( .A(n653), .B(n16943), .Z(n16942) );
  IV U16317 ( .A(n16938), .Z(n16940) );
  XOR U16318 ( .A(n16944), .B(n16945), .Z(n16938) );
  AND U16319 ( .A(n637), .B(n16937), .Z(n16945) );
  XNOR U16320 ( .A(n16935), .B(n16944), .Z(n16937) );
  XNOR U16321 ( .A(n16946), .B(n16947), .Z(n16935) );
  AND U16322 ( .A(n641), .B(n16948), .Z(n16947) );
  XOR U16323 ( .A(p_input[495]), .B(n16946), .Z(n16948) );
  XNOR U16324 ( .A(n16949), .B(n16950), .Z(n16946) );
  AND U16325 ( .A(n645), .B(n16951), .Z(n16950) );
  XOR U16326 ( .A(n16952), .B(n16953), .Z(n16944) );
  AND U16327 ( .A(n649), .B(n16943), .Z(n16953) );
  XNOR U16328 ( .A(n16954), .B(n16941), .Z(n16943) );
  XOR U16329 ( .A(n16955), .B(n16956), .Z(n16941) );
  AND U16330 ( .A(n672), .B(n16957), .Z(n16956) );
  IV U16331 ( .A(n16952), .Z(n16954) );
  XOR U16332 ( .A(n16958), .B(n16959), .Z(n16952) );
  AND U16333 ( .A(n656), .B(n16951), .Z(n16959) );
  XNOR U16334 ( .A(n16949), .B(n16958), .Z(n16951) );
  XNOR U16335 ( .A(n16960), .B(n16961), .Z(n16949) );
  AND U16336 ( .A(n660), .B(n16962), .Z(n16961) );
  XOR U16337 ( .A(p_input[511]), .B(n16960), .Z(n16962) );
  XNOR U16338 ( .A(n16963), .B(n16964), .Z(n16960) );
  AND U16339 ( .A(n664), .B(n16965), .Z(n16964) );
  XOR U16340 ( .A(n16966), .B(n16967), .Z(n16958) );
  AND U16341 ( .A(n668), .B(n16957), .Z(n16967) );
  XNOR U16342 ( .A(n16968), .B(n16955), .Z(n16957) );
  XOR U16343 ( .A(n16969), .B(n16970), .Z(n16955) );
  AND U16344 ( .A(n691), .B(n16971), .Z(n16970) );
  IV U16345 ( .A(n16966), .Z(n16968) );
  XOR U16346 ( .A(n16972), .B(n16973), .Z(n16966) );
  AND U16347 ( .A(n675), .B(n16965), .Z(n16973) );
  XNOR U16348 ( .A(n16963), .B(n16972), .Z(n16965) );
  XNOR U16349 ( .A(n16974), .B(n16975), .Z(n16963) );
  AND U16350 ( .A(n679), .B(n16976), .Z(n16975) );
  XOR U16351 ( .A(p_input[527]), .B(n16974), .Z(n16976) );
  XNOR U16352 ( .A(n16977), .B(n16978), .Z(n16974) );
  AND U16353 ( .A(n683), .B(n16979), .Z(n16978) );
  XOR U16354 ( .A(n16980), .B(n16981), .Z(n16972) );
  AND U16355 ( .A(n687), .B(n16971), .Z(n16981) );
  XNOR U16356 ( .A(n16982), .B(n16969), .Z(n16971) );
  XOR U16357 ( .A(n16983), .B(n16984), .Z(n16969) );
  AND U16358 ( .A(n710), .B(n16985), .Z(n16984) );
  IV U16359 ( .A(n16980), .Z(n16982) );
  XOR U16360 ( .A(n16986), .B(n16987), .Z(n16980) );
  AND U16361 ( .A(n694), .B(n16979), .Z(n16987) );
  XNOR U16362 ( .A(n16977), .B(n16986), .Z(n16979) );
  XNOR U16363 ( .A(n16988), .B(n16989), .Z(n16977) );
  AND U16364 ( .A(n698), .B(n16990), .Z(n16989) );
  XOR U16365 ( .A(p_input[543]), .B(n16988), .Z(n16990) );
  XNOR U16366 ( .A(n16991), .B(n16992), .Z(n16988) );
  AND U16367 ( .A(n702), .B(n16993), .Z(n16992) );
  XOR U16368 ( .A(n16994), .B(n16995), .Z(n16986) );
  AND U16369 ( .A(n706), .B(n16985), .Z(n16995) );
  XNOR U16370 ( .A(n16996), .B(n16983), .Z(n16985) );
  XOR U16371 ( .A(n16997), .B(n16998), .Z(n16983) );
  AND U16372 ( .A(n729), .B(n16999), .Z(n16998) );
  IV U16373 ( .A(n16994), .Z(n16996) );
  XOR U16374 ( .A(n17000), .B(n17001), .Z(n16994) );
  AND U16375 ( .A(n713), .B(n16993), .Z(n17001) );
  XNOR U16376 ( .A(n16991), .B(n17000), .Z(n16993) );
  XNOR U16377 ( .A(n17002), .B(n17003), .Z(n16991) );
  AND U16378 ( .A(n717), .B(n17004), .Z(n17003) );
  XOR U16379 ( .A(p_input[559]), .B(n17002), .Z(n17004) );
  XNOR U16380 ( .A(n17005), .B(n17006), .Z(n17002) );
  AND U16381 ( .A(n721), .B(n17007), .Z(n17006) );
  XOR U16382 ( .A(n17008), .B(n17009), .Z(n17000) );
  AND U16383 ( .A(n725), .B(n16999), .Z(n17009) );
  XNOR U16384 ( .A(n17010), .B(n16997), .Z(n16999) );
  XOR U16385 ( .A(n17011), .B(n17012), .Z(n16997) );
  AND U16386 ( .A(n748), .B(n17013), .Z(n17012) );
  IV U16387 ( .A(n17008), .Z(n17010) );
  XOR U16388 ( .A(n17014), .B(n17015), .Z(n17008) );
  AND U16389 ( .A(n732), .B(n17007), .Z(n17015) );
  XNOR U16390 ( .A(n17005), .B(n17014), .Z(n17007) );
  XNOR U16391 ( .A(n17016), .B(n17017), .Z(n17005) );
  AND U16392 ( .A(n736), .B(n17018), .Z(n17017) );
  XOR U16393 ( .A(p_input[575]), .B(n17016), .Z(n17018) );
  XNOR U16394 ( .A(n17019), .B(n17020), .Z(n17016) );
  AND U16395 ( .A(n740), .B(n17021), .Z(n17020) );
  XOR U16396 ( .A(n17022), .B(n17023), .Z(n17014) );
  AND U16397 ( .A(n744), .B(n17013), .Z(n17023) );
  XNOR U16398 ( .A(n17024), .B(n17011), .Z(n17013) );
  XOR U16399 ( .A(n17025), .B(n17026), .Z(n17011) );
  AND U16400 ( .A(n767), .B(n17027), .Z(n17026) );
  IV U16401 ( .A(n17022), .Z(n17024) );
  XOR U16402 ( .A(n17028), .B(n17029), .Z(n17022) );
  AND U16403 ( .A(n751), .B(n17021), .Z(n17029) );
  XNOR U16404 ( .A(n17019), .B(n17028), .Z(n17021) );
  XNOR U16405 ( .A(n17030), .B(n17031), .Z(n17019) );
  AND U16406 ( .A(n755), .B(n17032), .Z(n17031) );
  XOR U16407 ( .A(p_input[591]), .B(n17030), .Z(n17032) );
  XNOR U16408 ( .A(n17033), .B(n17034), .Z(n17030) );
  AND U16409 ( .A(n759), .B(n17035), .Z(n17034) );
  XOR U16410 ( .A(n17036), .B(n17037), .Z(n17028) );
  AND U16411 ( .A(n763), .B(n17027), .Z(n17037) );
  XNOR U16412 ( .A(n17038), .B(n17025), .Z(n17027) );
  XOR U16413 ( .A(n17039), .B(n17040), .Z(n17025) );
  AND U16414 ( .A(n786), .B(n17041), .Z(n17040) );
  IV U16415 ( .A(n17036), .Z(n17038) );
  XOR U16416 ( .A(n17042), .B(n17043), .Z(n17036) );
  AND U16417 ( .A(n770), .B(n17035), .Z(n17043) );
  XNOR U16418 ( .A(n17033), .B(n17042), .Z(n17035) );
  XNOR U16419 ( .A(n17044), .B(n17045), .Z(n17033) );
  AND U16420 ( .A(n774), .B(n17046), .Z(n17045) );
  XOR U16421 ( .A(p_input[607]), .B(n17044), .Z(n17046) );
  XNOR U16422 ( .A(n17047), .B(n17048), .Z(n17044) );
  AND U16423 ( .A(n778), .B(n17049), .Z(n17048) );
  XOR U16424 ( .A(n17050), .B(n17051), .Z(n17042) );
  AND U16425 ( .A(n782), .B(n17041), .Z(n17051) );
  XNOR U16426 ( .A(n17052), .B(n17039), .Z(n17041) );
  XOR U16427 ( .A(n17053), .B(n17054), .Z(n17039) );
  AND U16428 ( .A(n805), .B(n17055), .Z(n17054) );
  IV U16429 ( .A(n17050), .Z(n17052) );
  XOR U16430 ( .A(n17056), .B(n17057), .Z(n17050) );
  AND U16431 ( .A(n789), .B(n17049), .Z(n17057) );
  XNOR U16432 ( .A(n17047), .B(n17056), .Z(n17049) );
  XNOR U16433 ( .A(n17058), .B(n17059), .Z(n17047) );
  AND U16434 ( .A(n793), .B(n17060), .Z(n17059) );
  XOR U16435 ( .A(p_input[623]), .B(n17058), .Z(n17060) );
  XNOR U16436 ( .A(n17061), .B(n17062), .Z(n17058) );
  AND U16437 ( .A(n797), .B(n17063), .Z(n17062) );
  XOR U16438 ( .A(n17064), .B(n17065), .Z(n17056) );
  AND U16439 ( .A(n801), .B(n17055), .Z(n17065) );
  XNOR U16440 ( .A(n17066), .B(n17053), .Z(n17055) );
  XOR U16441 ( .A(n17067), .B(n17068), .Z(n17053) );
  AND U16442 ( .A(n824), .B(n17069), .Z(n17068) );
  IV U16443 ( .A(n17064), .Z(n17066) );
  XOR U16444 ( .A(n17070), .B(n17071), .Z(n17064) );
  AND U16445 ( .A(n808), .B(n17063), .Z(n17071) );
  XNOR U16446 ( .A(n17061), .B(n17070), .Z(n17063) );
  XNOR U16447 ( .A(n17072), .B(n17073), .Z(n17061) );
  AND U16448 ( .A(n812), .B(n17074), .Z(n17073) );
  XOR U16449 ( .A(p_input[639]), .B(n17072), .Z(n17074) );
  XNOR U16450 ( .A(n17075), .B(n17076), .Z(n17072) );
  AND U16451 ( .A(n816), .B(n17077), .Z(n17076) );
  XOR U16452 ( .A(n17078), .B(n17079), .Z(n17070) );
  AND U16453 ( .A(n820), .B(n17069), .Z(n17079) );
  XNOR U16454 ( .A(n17080), .B(n17067), .Z(n17069) );
  XOR U16455 ( .A(n17081), .B(n17082), .Z(n17067) );
  AND U16456 ( .A(n843), .B(n17083), .Z(n17082) );
  IV U16457 ( .A(n17078), .Z(n17080) );
  XOR U16458 ( .A(n17084), .B(n17085), .Z(n17078) );
  AND U16459 ( .A(n827), .B(n17077), .Z(n17085) );
  XNOR U16460 ( .A(n17075), .B(n17084), .Z(n17077) );
  XNOR U16461 ( .A(n17086), .B(n17087), .Z(n17075) );
  AND U16462 ( .A(n831), .B(n17088), .Z(n17087) );
  XOR U16463 ( .A(p_input[655]), .B(n17086), .Z(n17088) );
  XNOR U16464 ( .A(n17089), .B(n17090), .Z(n17086) );
  AND U16465 ( .A(n835), .B(n17091), .Z(n17090) );
  XOR U16466 ( .A(n17092), .B(n17093), .Z(n17084) );
  AND U16467 ( .A(n839), .B(n17083), .Z(n17093) );
  XNOR U16468 ( .A(n17094), .B(n17081), .Z(n17083) );
  XOR U16469 ( .A(n17095), .B(n17096), .Z(n17081) );
  AND U16470 ( .A(n862), .B(n17097), .Z(n17096) );
  IV U16471 ( .A(n17092), .Z(n17094) );
  XOR U16472 ( .A(n17098), .B(n17099), .Z(n17092) );
  AND U16473 ( .A(n846), .B(n17091), .Z(n17099) );
  XNOR U16474 ( .A(n17089), .B(n17098), .Z(n17091) );
  XNOR U16475 ( .A(n17100), .B(n17101), .Z(n17089) );
  AND U16476 ( .A(n850), .B(n17102), .Z(n17101) );
  XOR U16477 ( .A(p_input[671]), .B(n17100), .Z(n17102) );
  XNOR U16478 ( .A(n17103), .B(n17104), .Z(n17100) );
  AND U16479 ( .A(n854), .B(n17105), .Z(n17104) );
  XOR U16480 ( .A(n17106), .B(n17107), .Z(n17098) );
  AND U16481 ( .A(n858), .B(n17097), .Z(n17107) );
  XNOR U16482 ( .A(n17108), .B(n17095), .Z(n17097) );
  XOR U16483 ( .A(n17109), .B(n17110), .Z(n17095) );
  AND U16484 ( .A(n881), .B(n17111), .Z(n17110) );
  IV U16485 ( .A(n17106), .Z(n17108) );
  XOR U16486 ( .A(n17112), .B(n17113), .Z(n17106) );
  AND U16487 ( .A(n865), .B(n17105), .Z(n17113) );
  XNOR U16488 ( .A(n17103), .B(n17112), .Z(n17105) );
  XNOR U16489 ( .A(n17114), .B(n17115), .Z(n17103) );
  AND U16490 ( .A(n869), .B(n17116), .Z(n17115) );
  XOR U16491 ( .A(p_input[687]), .B(n17114), .Z(n17116) );
  XNOR U16492 ( .A(n17117), .B(n17118), .Z(n17114) );
  AND U16493 ( .A(n873), .B(n17119), .Z(n17118) );
  XOR U16494 ( .A(n17120), .B(n17121), .Z(n17112) );
  AND U16495 ( .A(n877), .B(n17111), .Z(n17121) );
  XNOR U16496 ( .A(n17122), .B(n17109), .Z(n17111) );
  XOR U16497 ( .A(n17123), .B(n17124), .Z(n17109) );
  AND U16498 ( .A(n900), .B(n17125), .Z(n17124) );
  IV U16499 ( .A(n17120), .Z(n17122) );
  XOR U16500 ( .A(n17126), .B(n17127), .Z(n17120) );
  AND U16501 ( .A(n884), .B(n17119), .Z(n17127) );
  XNOR U16502 ( .A(n17117), .B(n17126), .Z(n17119) );
  XNOR U16503 ( .A(n17128), .B(n17129), .Z(n17117) );
  AND U16504 ( .A(n888), .B(n17130), .Z(n17129) );
  XOR U16505 ( .A(p_input[703]), .B(n17128), .Z(n17130) );
  XNOR U16506 ( .A(n17131), .B(n17132), .Z(n17128) );
  AND U16507 ( .A(n892), .B(n17133), .Z(n17132) );
  XOR U16508 ( .A(n17134), .B(n17135), .Z(n17126) );
  AND U16509 ( .A(n896), .B(n17125), .Z(n17135) );
  XNOR U16510 ( .A(n17136), .B(n17123), .Z(n17125) );
  XOR U16511 ( .A(n17137), .B(n17138), .Z(n17123) );
  AND U16512 ( .A(n919), .B(n17139), .Z(n17138) );
  IV U16513 ( .A(n17134), .Z(n17136) );
  XOR U16514 ( .A(n17140), .B(n17141), .Z(n17134) );
  AND U16515 ( .A(n903), .B(n17133), .Z(n17141) );
  XNOR U16516 ( .A(n17131), .B(n17140), .Z(n17133) );
  XNOR U16517 ( .A(n17142), .B(n17143), .Z(n17131) );
  AND U16518 ( .A(n907), .B(n17144), .Z(n17143) );
  XOR U16519 ( .A(p_input[719]), .B(n17142), .Z(n17144) );
  XNOR U16520 ( .A(n17145), .B(n17146), .Z(n17142) );
  AND U16521 ( .A(n911), .B(n17147), .Z(n17146) );
  XOR U16522 ( .A(n17148), .B(n17149), .Z(n17140) );
  AND U16523 ( .A(n915), .B(n17139), .Z(n17149) );
  XNOR U16524 ( .A(n17150), .B(n17137), .Z(n17139) );
  XOR U16525 ( .A(n17151), .B(n17152), .Z(n17137) );
  AND U16526 ( .A(n938), .B(n17153), .Z(n17152) );
  IV U16527 ( .A(n17148), .Z(n17150) );
  XOR U16528 ( .A(n17154), .B(n17155), .Z(n17148) );
  AND U16529 ( .A(n922), .B(n17147), .Z(n17155) );
  XNOR U16530 ( .A(n17145), .B(n17154), .Z(n17147) );
  XNOR U16531 ( .A(n17156), .B(n17157), .Z(n17145) );
  AND U16532 ( .A(n926), .B(n17158), .Z(n17157) );
  XOR U16533 ( .A(p_input[735]), .B(n17156), .Z(n17158) );
  XNOR U16534 ( .A(n17159), .B(n17160), .Z(n17156) );
  AND U16535 ( .A(n930), .B(n17161), .Z(n17160) );
  XOR U16536 ( .A(n17162), .B(n17163), .Z(n17154) );
  AND U16537 ( .A(n934), .B(n17153), .Z(n17163) );
  XNOR U16538 ( .A(n17164), .B(n17151), .Z(n17153) );
  XOR U16539 ( .A(n17165), .B(n17166), .Z(n17151) );
  AND U16540 ( .A(n957), .B(n17167), .Z(n17166) );
  IV U16541 ( .A(n17162), .Z(n17164) );
  XOR U16542 ( .A(n17168), .B(n17169), .Z(n17162) );
  AND U16543 ( .A(n941), .B(n17161), .Z(n17169) );
  XNOR U16544 ( .A(n17159), .B(n17168), .Z(n17161) );
  XNOR U16545 ( .A(n17170), .B(n17171), .Z(n17159) );
  AND U16546 ( .A(n945), .B(n17172), .Z(n17171) );
  XOR U16547 ( .A(p_input[751]), .B(n17170), .Z(n17172) );
  XNOR U16548 ( .A(n17173), .B(n17174), .Z(n17170) );
  AND U16549 ( .A(n949), .B(n17175), .Z(n17174) );
  XOR U16550 ( .A(n17176), .B(n17177), .Z(n17168) );
  AND U16551 ( .A(n953), .B(n17167), .Z(n17177) );
  XNOR U16552 ( .A(n17178), .B(n17165), .Z(n17167) );
  XOR U16553 ( .A(n17179), .B(n17180), .Z(n17165) );
  AND U16554 ( .A(n976), .B(n17181), .Z(n17180) );
  IV U16555 ( .A(n17176), .Z(n17178) );
  XOR U16556 ( .A(n17182), .B(n17183), .Z(n17176) );
  AND U16557 ( .A(n960), .B(n17175), .Z(n17183) );
  XNOR U16558 ( .A(n17173), .B(n17182), .Z(n17175) );
  XNOR U16559 ( .A(n17184), .B(n17185), .Z(n17173) );
  AND U16560 ( .A(n964), .B(n17186), .Z(n17185) );
  XOR U16561 ( .A(p_input[767]), .B(n17184), .Z(n17186) );
  XNOR U16562 ( .A(n17187), .B(n17188), .Z(n17184) );
  AND U16563 ( .A(n968), .B(n17189), .Z(n17188) );
  XOR U16564 ( .A(n17190), .B(n17191), .Z(n17182) );
  AND U16565 ( .A(n972), .B(n17181), .Z(n17191) );
  XNOR U16566 ( .A(n17192), .B(n17179), .Z(n17181) );
  XOR U16567 ( .A(n17193), .B(n17194), .Z(n17179) );
  AND U16568 ( .A(n995), .B(n17195), .Z(n17194) );
  IV U16569 ( .A(n17190), .Z(n17192) );
  XOR U16570 ( .A(n17196), .B(n17197), .Z(n17190) );
  AND U16571 ( .A(n979), .B(n17189), .Z(n17197) );
  XNOR U16572 ( .A(n17187), .B(n17196), .Z(n17189) );
  XNOR U16573 ( .A(n17198), .B(n17199), .Z(n17187) );
  AND U16574 ( .A(n983), .B(n17200), .Z(n17199) );
  XOR U16575 ( .A(p_input[783]), .B(n17198), .Z(n17200) );
  XNOR U16576 ( .A(n17201), .B(n17202), .Z(n17198) );
  AND U16577 ( .A(n987), .B(n17203), .Z(n17202) );
  XOR U16578 ( .A(n17204), .B(n17205), .Z(n17196) );
  AND U16579 ( .A(n991), .B(n17195), .Z(n17205) );
  XNOR U16580 ( .A(n17206), .B(n17193), .Z(n17195) );
  XOR U16581 ( .A(n17207), .B(n17208), .Z(n17193) );
  AND U16582 ( .A(n1014), .B(n17209), .Z(n17208) );
  IV U16583 ( .A(n17204), .Z(n17206) );
  XOR U16584 ( .A(n17210), .B(n17211), .Z(n17204) );
  AND U16585 ( .A(n998), .B(n17203), .Z(n17211) );
  XNOR U16586 ( .A(n17201), .B(n17210), .Z(n17203) );
  XNOR U16587 ( .A(n17212), .B(n17213), .Z(n17201) );
  AND U16588 ( .A(n1002), .B(n17214), .Z(n17213) );
  XOR U16589 ( .A(p_input[799]), .B(n17212), .Z(n17214) );
  XNOR U16590 ( .A(n17215), .B(n17216), .Z(n17212) );
  AND U16591 ( .A(n1006), .B(n17217), .Z(n17216) );
  XOR U16592 ( .A(n17218), .B(n17219), .Z(n17210) );
  AND U16593 ( .A(n1010), .B(n17209), .Z(n17219) );
  XNOR U16594 ( .A(n17220), .B(n17207), .Z(n17209) );
  XOR U16595 ( .A(n17221), .B(n17222), .Z(n17207) );
  AND U16596 ( .A(n1033), .B(n17223), .Z(n17222) );
  IV U16597 ( .A(n17218), .Z(n17220) );
  XOR U16598 ( .A(n17224), .B(n17225), .Z(n17218) );
  AND U16599 ( .A(n1017), .B(n17217), .Z(n17225) );
  XNOR U16600 ( .A(n17215), .B(n17224), .Z(n17217) );
  XNOR U16601 ( .A(n17226), .B(n17227), .Z(n17215) );
  AND U16602 ( .A(n1021), .B(n17228), .Z(n17227) );
  XOR U16603 ( .A(p_input[815]), .B(n17226), .Z(n17228) );
  XNOR U16604 ( .A(n17229), .B(n17230), .Z(n17226) );
  AND U16605 ( .A(n1025), .B(n17231), .Z(n17230) );
  XOR U16606 ( .A(n17232), .B(n17233), .Z(n17224) );
  AND U16607 ( .A(n1029), .B(n17223), .Z(n17233) );
  XNOR U16608 ( .A(n17234), .B(n17221), .Z(n17223) );
  XOR U16609 ( .A(n17235), .B(n17236), .Z(n17221) );
  AND U16610 ( .A(n1052), .B(n17237), .Z(n17236) );
  IV U16611 ( .A(n17232), .Z(n17234) );
  XOR U16612 ( .A(n17238), .B(n17239), .Z(n17232) );
  AND U16613 ( .A(n1036), .B(n17231), .Z(n17239) );
  XNOR U16614 ( .A(n17229), .B(n17238), .Z(n17231) );
  XNOR U16615 ( .A(n17240), .B(n17241), .Z(n17229) );
  AND U16616 ( .A(n1040), .B(n17242), .Z(n17241) );
  XOR U16617 ( .A(p_input[831]), .B(n17240), .Z(n17242) );
  XNOR U16618 ( .A(n17243), .B(n17244), .Z(n17240) );
  AND U16619 ( .A(n1044), .B(n17245), .Z(n17244) );
  XOR U16620 ( .A(n17246), .B(n17247), .Z(n17238) );
  AND U16621 ( .A(n1048), .B(n17237), .Z(n17247) );
  XNOR U16622 ( .A(n17248), .B(n17235), .Z(n17237) );
  XOR U16623 ( .A(n17249), .B(n17250), .Z(n17235) );
  AND U16624 ( .A(n1071), .B(n17251), .Z(n17250) );
  IV U16625 ( .A(n17246), .Z(n17248) );
  XOR U16626 ( .A(n17252), .B(n17253), .Z(n17246) );
  AND U16627 ( .A(n1055), .B(n17245), .Z(n17253) );
  XNOR U16628 ( .A(n17243), .B(n17252), .Z(n17245) );
  XNOR U16629 ( .A(n17254), .B(n17255), .Z(n17243) );
  AND U16630 ( .A(n1059), .B(n17256), .Z(n17255) );
  XOR U16631 ( .A(p_input[847]), .B(n17254), .Z(n17256) );
  XNOR U16632 ( .A(n17257), .B(n17258), .Z(n17254) );
  AND U16633 ( .A(n1063), .B(n17259), .Z(n17258) );
  XOR U16634 ( .A(n17260), .B(n17261), .Z(n17252) );
  AND U16635 ( .A(n1067), .B(n17251), .Z(n17261) );
  XNOR U16636 ( .A(n17262), .B(n17249), .Z(n17251) );
  XOR U16637 ( .A(n17263), .B(n17264), .Z(n17249) );
  AND U16638 ( .A(n1090), .B(n17265), .Z(n17264) );
  IV U16639 ( .A(n17260), .Z(n17262) );
  XOR U16640 ( .A(n17266), .B(n17267), .Z(n17260) );
  AND U16641 ( .A(n1074), .B(n17259), .Z(n17267) );
  XNOR U16642 ( .A(n17257), .B(n17266), .Z(n17259) );
  XNOR U16643 ( .A(n17268), .B(n17269), .Z(n17257) );
  AND U16644 ( .A(n1078), .B(n17270), .Z(n17269) );
  XOR U16645 ( .A(p_input[863]), .B(n17268), .Z(n17270) );
  XNOR U16646 ( .A(n17271), .B(n17272), .Z(n17268) );
  AND U16647 ( .A(n1082), .B(n17273), .Z(n17272) );
  XOR U16648 ( .A(n17274), .B(n17275), .Z(n17266) );
  AND U16649 ( .A(n1086), .B(n17265), .Z(n17275) );
  XNOR U16650 ( .A(n17276), .B(n17263), .Z(n17265) );
  XOR U16651 ( .A(n17277), .B(n17278), .Z(n17263) );
  AND U16652 ( .A(n1109), .B(n17279), .Z(n17278) );
  IV U16653 ( .A(n17274), .Z(n17276) );
  XOR U16654 ( .A(n17280), .B(n17281), .Z(n17274) );
  AND U16655 ( .A(n1093), .B(n17273), .Z(n17281) );
  XNOR U16656 ( .A(n17271), .B(n17280), .Z(n17273) );
  XNOR U16657 ( .A(n17282), .B(n17283), .Z(n17271) );
  AND U16658 ( .A(n1097), .B(n17284), .Z(n17283) );
  XOR U16659 ( .A(p_input[879]), .B(n17282), .Z(n17284) );
  XNOR U16660 ( .A(n17285), .B(n17286), .Z(n17282) );
  AND U16661 ( .A(n1101), .B(n17287), .Z(n17286) );
  XOR U16662 ( .A(n17288), .B(n17289), .Z(n17280) );
  AND U16663 ( .A(n1105), .B(n17279), .Z(n17289) );
  XNOR U16664 ( .A(n17290), .B(n17277), .Z(n17279) );
  XOR U16665 ( .A(n17291), .B(n17292), .Z(n17277) );
  AND U16666 ( .A(n1128), .B(n17293), .Z(n17292) );
  IV U16667 ( .A(n17288), .Z(n17290) );
  XOR U16668 ( .A(n17294), .B(n17295), .Z(n17288) );
  AND U16669 ( .A(n1112), .B(n17287), .Z(n17295) );
  XNOR U16670 ( .A(n17285), .B(n17294), .Z(n17287) );
  XNOR U16671 ( .A(n17296), .B(n17297), .Z(n17285) );
  AND U16672 ( .A(n1116), .B(n17298), .Z(n17297) );
  XOR U16673 ( .A(p_input[895]), .B(n17296), .Z(n17298) );
  XNOR U16674 ( .A(n17299), .B(n17300), .Z(n17296) );
  AND U16675 ( .A(n1120), .B(n17301), .Z(n17300) );
  XOR U16676 ( .A(n17302), .B(n17303), .Z(n17294) );
  AND U16677 ( .A(n1124), .B(n17293), .Z(n17303) );
  XNOR U16678 ( .A(n17304), .B(n17291), .Z(n17293) );
  XOR U16679 ( .A(n17305), .B(n17306), .Z(n17291) );
  AND U16680 ( .A(n1147), .B(n17307), .Z(n17306) );
  IV U16681 ( .A(n17302), .Z(n17304) );
  XOR U16682 ( .A(n17308), .B(n17309), .Z(n17302) );
  AND U16683 ( .A(n1131), .B(n17301), .Z(n17309) );
  XNOR U16684 ( .A(n17299), .B(n17308), .Z(n17301) );
  XNOR U16685 ( .A(n17310), .B(n17311), .Z(n17299) );
  AND U16686 ( .A(n1135), .B(n17312), .Z(n17311) );
  XOR U16687 ( .A(p_input[911]), .B(n17310), .Z(n17312) );
  XNOR U16688 ( .A(n17313), .B(n17314), .Z(n17310) );
  AND U16689 ( .A(n1139), .B(n17315), .Z(n17314) );
  XOR U16690 ( .A(n17316), .B(n17317), .Z(n17308) );
  AND U16691 ( .A(n1143), .B(n17307), .Z(n17317) );
  XNOR U16692 ( .A(n17318), .B(n17305), .Z(n17307) );
  XOR U16693 ( .A(n17319), .B(n17320), .Z(n17305) );
  AND U16694 ( .A(n1166), .B(n17321), .Z(n17320) );
  IV U16695 ( .A(n17316), .Z(n17318) );
  XOR U16696 ( .A(n17322), .B(n17323), .Z(n17316) );
  AND U16697 ( .A(n1150), .B(n17315), .Z(n17323) );
  XNOR U16698 ( .A(n17313), .B(n17322), .Z(n17315) );
  XNOR U16699 ( .A(n17324), .B(n17325), .Z(n17313) );
  AND U16700 ( .A(n1154), .B(n17326), .Z(n17325) );
  XOR U16701 ( .A(p_input[927]), .B(n17324), .Z(n17326) );
  XNOR U16702 ( .A(n17327), .B(n17328), .Z(n17324) );
  AND U16703 ( .A(n1158), .B(n17329), .Z(n17328) );
  XOR U16704 ( .A(n17330), .B(n17331), .Z(n17322) );
  AND U16705 ( .A(n1162), .B(n17321), .Z(n17331) );
  XNOR U16706 ( .A(n17332), .B(n17319), .Z(n17321) );
  XOR U16707 ( .A(n17333), .B(n17334), .Z(n17319) );
  AND U16708 ( .A(n1185), .B(n17335), .Z(n17334) );
  IV U16709 ( .A(n17330), .Z(n17332) );
  XOR U16710 ( .A(n17336), .B(n17337), .Z(n17330) );
  AND U16711 ( .A(n1169), .B(n17329), .Z(n17337) );
  XNOR U16712 ( .A(n17327), .B(n17336), .Z(n17329) );
  XNOR U16713 ( .A(n17338), .B(n17339), .Z(n17327) );
  AND U16714 ( .A(n1173), .B(n17340), .Z(n17339) );
  XOR U16715 ( .A(p_input[943]), .B(n17338), .Z(n17340) );
  XNOR U16716 ( .A(n17341), .B(n17342), .Z(n17338) );
  AND U16717 ( .A(n1177), .B(n17343), .Z(n17342) );
  XOR U16718 ( .A(n17344), .B(n17345), .Z(n17336) );
  AND U16719 ( .A(n1181), .B(n17335), .Z(n17345) );
  XNOR U16720 ( .A(n17346), .B(n17333), .Z(n17335) );
  XOR U16721 ( .A(n17347), .B(n17348), .Z(n17333) );
  AND U16722 ( .A(n1204), .B(n17349), .Z(n17348) );
  IV U16723 ( .A(n17344), .Z(n17346) );
  XOR U16724 ( .A(n17350), .B(n17351), .Z(n17344) );
  AND U16725 ( .A(n1188), .B(n17343), .Z(n17351) );
  XNOR U16726 ( .A(n17341), .B(n17350), .Z(n17343) );
  XNOR U16727 ( .A(n17352), .B(n17353), .Z(n17341) );
  AND U16728 ( .A(n1192), .B(n17354), .Z(n17353) );
  XOR U16729 ( .A(p_input[959]), .B(n17352), .Z(n17354) );
  XNOR U16730 ( .A(n17355), .B(n17356), .Z(n17352) );
  AND U16731 ( .A(n1196), .B(n17357), .Z(n17356) );
  XOR U16732 ( .A(n17358), .B(n17359), .Z(n17350) );
  AND U16733 ( .A(n1200), .B(n17349), .Z(n17359) );
  XNOR U16734 ( .A(n17360), .B(n17347), .Z(n17349) );
  XOR U16735 ( .A(n17361), .B(n17362), .Z(n17347) );
  AND U16736 ( .A(n1223), .B(n17363), .Z(n17362) );
  IV U16737 ( .A(n17358), .Z(n17360) );
  XOR U16738 ( .A(n17364), .B(n17365), .Z(n17358) );
  AND U16739 ( .A(n1207), .B(n17357), .Z(n17365) );
  XNOR U16740 ( .A(n17355), .B(n17364), .Z(n17357) );
  XNOR U16741 ( .A(n17366), .B(n17367), .Z(n17355) );
  AND U16742 ( .A(n1211), .B(n17368), .Z(n17367) );
  XOR U16743 ( .A(p_input[975]), .B(n17366), .Z(n17368) );
  XNOR U16744 ( .A(n17369), .B(n17370), .Z(n17366) );
  AND U16745 ( .A(n1215), .B(n17371), .Z(n17370) );
  XOR U16746 ( .A(n17372), .B(n17373), .Z(n17364) );
  AND U16747 ( .A(n1219), .B(n17363), .Z(n17373) );
  XNOR U16748 ( .A(n17374), .B(n17361), .Z(n17363) );
  XOR U16749 ( .A(n17375), .B(n17376), .Z(n17361) );
  AND U16750 ( .A(n1242), .B(n17377), .Z(n17376) );
  IV U16751 ( .A(n17372), .Z(n17374) );
  XOR U16752 ( .A(n17378), .B(n17379), .Z(n17372) );
  AND U16753 ( .A(n1226), .B(n17371), .Z(n17379) );
  XNOR U16754 ( .A(n17369), .B(n17378), .Z(n17371) );
  XNOR U16755 ( .A(n17380), .B(n17381), .Z(n17369) );
  AND U16756 ( .A(n1230), .B(n17382), .Z(n17381) );
  XOR U16757 ( .A(p_input[991]), .B(n17380), .Z(n17382) );
  XNOR U16758 ( .A(n17383), .B(n17384), .Z(n17380) );
  AND U16759 ( .A(n1234), .B(n17385), .Z(n17384) );
  XOR U16760 ( .A(n17386), .B(n17387), .Z(n17378) );
  AND U16761 ( .A(n1238), .B(n17377), .Z(n17387) );
  XNOR U16762 ( .A(n17388), .B(n17375), .Z(n17377) );
  XOR U16763 ( .A(n17389), .B(n17390), .Z(n17375) );
  AND U16764 ( .A(n1261), .B(n17391), .Z(n17390) );
  IV U16765 ( .A(n17386), .Z(n17388) );
  XOR U16766 ( .A(n17392), .B(n17393), .Z(n17386) );
  AND U16767 ( .A(n1245), .B(n17385), .Z(n17393) );
  XNOR U16768 ( .A(n17383), .B(n17392), .Z(n17385) );
  XNOR U16769 ( .A(n17394), .B(n17395), .Z(n17383) );
  AND U16770 ( .A(n1249), .B(n17396), .Z(n17395) );
  XOR U16771 ( .A(p_input[1007]), .B(n17394), .Z(n17396) );
  XNOR U16772 ( .A(n17397), .B(n17398), .Z(n17394) );
  AND U16773 ( .A(n1253), .B(n17399), .Z(n17398) );
  XOR U16774 ( .A(n17400), .B(n17401), .Z(n17392) );
  AND U16775 ( .A(n1257), .B(n17391), .Z(n17401) );
  XNOR U16776 ( .A(n17402), .B(n17389), .Z(n17391) );
  XOR U16777 ( .A(n17403), .B(n17404), .Z(n17389) );
  AND U16778 ( .A(n1280), .B(n17405), .Z(n17404) );
  IV U16779 ( .A(n17400), .Z(n17402) );
  XOR U16780 ( .A(n17406), .B(n17407), .Z(n17400) );
  AND U16781 ( .A(n1264), .B(n17399), .Z(n17407) );
  XNOR U16782 ( .A(n17397), .B(n17406), .Z(n17399) );
  XNOR U16783 ( .A(n17408), .B(n17409), .Z(n17397) );
  AND U16784 ( .A(n1268), .B(n17410), .Z(n17409) );
  XOR U16785 ( .A(p_input[1023]), .B(n17408), .Z(n17410) );
  XNOR U16786 ( .A(n17411), .B(n17412), .Z(n17408) );
  AND U16787 ( .A(n1272), .B(n17413), .Z(n17412) );
  XOR U16788 ( .A(n17414), .B(n17415), .Z(n17406) );
  AND U16789 ( .A(n1276), .B(n17405), .Z(n17415) );
  XNOR U16790 ( .A(n17416), .B(n17403), .Z(n17405) );
  XOR U16791 ( .A(n17417), .B(n17418), .Z(n17403) );
  AND U16792 ( .A(n1299), .B(n17419), .Z(n17418) );
  IV U16793 ( .A(n17414), .Z(n17416) );
  XOR U16794 ( .A(n17420), .B(n17421), .Z(n17414) );
  AND U16795 ( .A(n1283), .B(n17413), .Z(n17421) );
  XNOR U16796 ( .A(n17411), .B(n17420), .Z(n17413) );
  XNOR U16797 ( .A(n17422), .B(n17423), .Z(n17411) );
  AND U16798 ( .A(n1287), .B(n17424), .Z(n17423) );
  XOR U16799 ( .A(p_input[1039]), .B(n17422), .Z(n17424) );
  XNOR U16800 ( .A(n17425), .B(n17426), .Z(n17422) );
  AND U16801 ( .A(n1291), .B(n17427), .Z(n17426) );
  XOR U16802 ( .A(n17428), .B(n17429), .Z(n17420) );
  AND U16803 ( .A(n1295), .B(n17419), .Z(n17429) );
  XNOR U16804 ( .A(n17430), .B(n17417), .Z(n17419) );
  XOR U16805 ( .A(n17431), .B(n17432), .Z(n17417) );
  AND U16806 ( .A(n1318), .B(n17433), .Z(n17432) );
  IV U16807 ( .A(n17428), .Z(n17430) );
  XOR U16808 ( .A(n17434), .B(n17435), .Z(n17428) );
  AND U16809 ( .A(n1302), .B(n17427), .Z(n17435) );
  XNOR U16810 ( .A(n17425), .B(n17434), .Z(n17427) );
  XNOR U16811 ( .A(n17436), .B(n17437), .Z(n17425) );
  AND U16812 ( .A(n1306), .B(n17438), .Z(n17437) );
  XOR U16813 ( .A(p_input[1055]), .B(n17436), .Z(n17438) );
  XNOR U16814 ( .A(n17439), .B(n17440), .Z(n17436) );
  AND U16815 ( .A(n1310), .B(n17441), .Z(n17440) );
  XOR U16816 ( .A(n17442), .B(n17443), .Z(n17434) );
  AND U16817 ( .A(n1314), .B(n17433), .Z(n17443) );
  XNOR U16818 ( .A(n17444), .B(n17431), .Z(n17433) );
  XOR U16819 ( .A(n17445), .B(n17446), .Z(n17431) );
  AND U16820 ( .A(n1337), .B(n17447), .Z(n17446) );
  IV U16821 ( .A(n17442), .Z(n17444) );
  XOR U16822 ( .A(n17448), .B(n17449), .Z(n17442) );
  AND U16823 ( .A(n1321), .B(n17441), .Z(n17449) );
  XNOR U16824 ( .A(n17439), .B(n17448), .Z(n17441) );
  XNOR U16825 ( .A(n17450), .B(n17451), .Z(n17439) );
  AND U16826 ( .A(n1325), .B(n17452), .Z(n17451) );
  XOR U16827 ( .A(p_input[1071]), .B(n17450), .Z(n17452) );
  XNOR U16828 ( .A(n17453), .B(n17454), .Z(n17450) );
  AND U16829 ( .A(n1329), .B(n17455), .Z(n17454) );
  XOR U16830 ( .A(n17456), .B(n17457), .Z(n17448) );
  AND U16831 ( .A(n1333), .B(n17447), .Z(n17457) );
  XNOR U16832 ( .A(n17458), .B(n17445), .Z(n17447) );
  XOR U16833 ( .A(n17459), .B(n17460), .Z(n17445) );
  AND U16834 ( .A(n1356), .B(n17461), .Z(n17460) );
  IV U16835 ( .A(n17456), .Z(n17458) );
  XOR U16836 ( .A(n17462), .B(n17463), .Z(n17456) );
  AND U16837 ( .A(n1340), .B(n17455), .Z(n17463) );
  XNOR U16838 ( .A(n17453), .B(n17462), .Z(n17455) );
  XNOR U16839 ( .A(n17464), .B(n17465), .Z(n17453) );
  AND U16840 ( .A(n1344), .B(n17466), .Z(n17465) );
  XOR U16841 ( .A(p_input[1087]), .B(n17464), .Z(n17466) );
  XNOR U16842 ( .A(n17467), .B(n17468), .Z(n17464) );
  AND U16843 ( .A(n1348), .B(n17469), .Z(n17468) );
  XOR U16844 ( .A(n17470), .B(n17471), .Z(n17462) );
  AND U16845 ( .A(n1352), .B(n17461), .Z(n17471) );
  XNOR U16846 ( .A(n17472), .B(n17459), .Z(n17461) );
  XOR U16847 ( .A(n17473), .B(n17474), .Z(n17459) );
  AND U16848 ( .A(n1375), .B(n17475), .Z(n17474) );
  IV U16849 ( .A(n17470), .Z(n17472) );
  XOR U16850 ( .A(n17476), .B(n17477), .Z(n17470) );
  AND U16851 ( .A(n1359), .B(n17469), .Z(n17477) );
  XNOR U16852 ( .A(n17467), .B(n17476), .Z(n17469) );
  XNOR U16853 ( .A(n17478), .B(n17479), .Z(n17467) );
  AND U16854 ( .A(n1363), .B(n17480), .Z(n17479) );
  XOR U16855 ( .A(p_input[1103]), .B(n17478), .Z(n17480) );
  XNOR U16856 ( .A(n17481), .B(n17482), .Z(n17478) );
  AND U16857 ( .A(n1367), .B(n17483), .Z(n17482) );
  XOR U16858 ( .A(n17484), .B(n17485), .Z(n17476) );
  AND U16859 ( .A(n1371), .B(n17475), .Z(n17485) );
  XNOR U16860 ( .A(n17486), .B(n17473), .Z(n17475) );
  XOR U16861 ( .A(n17487), .B(n17488), .Z(n17473) );
  AND U16862 ( .A(n1394), .B(n17489), .Z(n17488) );
  IV U16863 ( .A(n17484), .Z(n17486) );
  XOR U16864 ( .A(n17490), .B(n17491), .Z(n17484) );
  AND U16865 ( .A(n1378), .B(n17483), .Z(n17491) );
  XNOR U16866 ( .A(n17481), .B(n17490), .Z(n17483) );
  XNOR U16867 ( .A(n17492), .B(n17493), .Z(n17481) );
  AND U16868 ( .A(n1382), .B(n17494), .Z(n17493) );
  XOR U16869 ( .A(p_input[1119]), .B(n17492), .Z(n17494) );
  XNOR U16870 ( .A(n17495), .B(n17496), .Z(n17492) );
  AND U16871 ( .A(n1386), .B(n17497), .Z(n17496) );
  XOR U16872 ( .A(n17498), .B(n17499), .Z(n17490) );
  AND U16873 ( .A(n1390), .B(n17489), .Z(n17499) );
  XNOR U16874 ( .A(n17500), .B(n17487), .Z(n17489) );
  XOR U16875 ( .A(n17501), .B(n17502), .Z(n17487) );
  AND U16876 ( .A(n1413), .B(n17503), .Z(n17502) );
  IV U16877 ( .A(n17498), .Z(n17500) );
  XOR U16878 ( .A(n17504), .B(n17505), .Z(n17498) );
  AND U16879 ( .A(n1397), .B(n17497), .Z(n17505) );
  XNOR U16880 ( .A(n17495), .B(n17504), .Z(n17497) );
  XNOR U16881 ( .A(n17506), .B(n17507), .Z(n17495) );
  AND U16882 ( .A(n1401), .B(n17508), .Z(n17507) );
  XOR U16883 ( .A(p_input[1135]), .B(n17506), .Z(n17508) );
  XNOR U16884 ( .A(n17509), .B(n17510), .Z(n17506) );
  AND U16885 ( .A(n1405), .B(n17511), .Z(n17510) );
  XOR U16886 ( .A(n17512), .B(n17513), .Z(n17504) );
  AND U16887 ( .A(n1409), .B(n17503), .Z(n17513) );
  XNOR U16888 ( .A(n17514), .B(n17501), .Z(n17503) );
  XOR U16889 ( .A(n17515), .B(n17516), .Z(n17501) );
  AND U16890 ( .A(n1432), .B(n17517), .Z(n17516) );
  IV U16891 ( .A(n17512), .Z(n17514) );
  XOR U16892 ( .A(n17518), .B(n17519), .Z(n17512) );
  AND U16893 ( .A(n1416), .B(n17511), .Z(n17519) );
  XNOR U16894 ( .A(n17509), .B(n17518), .Z(n17511) );
  XNOR U16895 ( .A(n17520), .B(n17521), .Z(n17509) );
  AND U16896 ( .A(n1420), .B(n17522), .Z(n17521) );
  XOR U16897 ( .A(p_input[1151]), .B(n17520), .Z(n17522) );
  XNOR U16898 ( .A(n17523), .B(n17524), .Z(n17520) );
  AND U16899 ( .A(n1424), .B(n17525), .Z(n17524) );
  XOR U16900 ( .A(n17526), .B(n17527), .Z(n17518) );
  AND U16901 ( .A(n1428), .B(n17517), .Z(n17527) );
  XNOR U16902 ( .A(n17528), .B(n17515), .Z(n17517) );
  XOR U16903 ( .A(n17529), .B(n17530), .Z(n17515) );
  AND U16904 ( .A(n1451), .B(n17531), .Z(n17530) );
  IV U16905 ( .A(n17526), .Z(n17528) );
  XOR U16906 ( .A(n17532), .B(n17533), .Z(n17526) );
  AND U16907 ( .A(n1435), .B(n17525), .Z(n17533) );
  XNOR U16908 ( .A(n17523), .B(n17532), .Z(n17525) );
  XNOR U16909 ( .A(n17534), .B(n17535), .Z(n17523) );
  AND U16910 ( .A(n1439), .B(n17536), .Z(n17535) );
  XOR U16911 ( .A(p_input[1167]), .B(n17534), .Z(n17536) );
  XNOR U16912 ( .A(n17537), .B(n17538), .Z(n17534) );
  AND U16913 ( .A(n1443), .B(n17539), .Z(n17538) );
  XOR U16914 ( .A(n17540), .B(n17541), .Z(n17532) );
  AND U16915 ( .A(n1447), .B(n17531), .Z(n17541) );
  XNOR U16916 ( .A(n17542), .B(n17529), .Z(n17531) );
  XOR U16917 ( .A(n17543), .B(n17544), .Z(n17529) );
  AND U16918 ( .A(n1470), .B(n17545), .Z(n17544) );
  IV U16919 ( .A(n17540), .Z(n17542) );
  XOR U16920 ( .A(n17546), .B(n17547), .Z(n17540) );
  AND U16921 ( .A(n1454), .B(n17539), .Z(n17547) );
  XNOR U16922 ( .A(n17537), .B(n17546), .Z(n17539) );
  XNOR U16923 ( .A(n17548), .B(n17549), .Z(n17537) );
  AND U16924 ( .A(n1458), .B(n17550), .Z(n17549) );
  XOR U16925 ( .A(p_input[1183]), .B(n17548), .Z(n17550) );
  XNOR U16926 ( .A(n17551), .B(n17552), .Z(n17548) );
  AND U16927 ( .A(n1462), .B(n17553), .Z(n17552) );
  XOR U16928 ( .A(n17554), .B(n17555), .Z(n17546) );
  AND U16929 ( .A(n1466), .B(n17545), .Z(n17555) );
  XNOR U16930 ( .A(n17556), .B(n17543), .Z(n17545) );
  XOR U16931 ( .A(n17557), .B(n17558), .Z(n17543) );
  AND U16932 ( .A(n1489), .B(n17559), .Z(n17558) );
  IV U16933 ( .A(n17554), .Z(n17556) );
  XOR U16934 ( .A(n17560), .B(n17561), .Z(n17554) );
  AND U16935 ( .A(n1473), .B(n17553), .Z(n17561) );
  XNOR U16936 ( .A(n17551), .B(n17560), .Z(n17553) );
  XNOR U16937 ( .A(n17562), .B(n17563), .Z(n17551) );
  AND U16938 ( .A(n1477), .B(n17564), .Z(n17563) );
  XOR U16939 ( .A(p_input[1199]), .B(n17562), .Z(n17564) );
  XNOR U16940 ( .A(n17565), .B(n17566), .Z(n17562) );
  AND U16941 ( .A(n1481), .B(n17567), .Z(n17566) );
  XOR U16942 ( .A(n17568), .B(n17569), .Z(n17560) );
  AND U16943 ( .A(n1485), .B(n17559), .Z(n17569) );
  XNOR U16944 ( .A(n17570), .B(n17557), .Z(n17559) );
  XOR U16945 ( .A(n17571), .B(n17572), .Z(n17557) );
  AND U16946 ( .A(n1508), .B(n17573), .Z(n17572) );
  IV U16947 ( .A(n17568), .Z(n17570) );
  XOR U16948 ( .A(n17574), .B(n17575), .Z(n17568) );
  AND U16949 ( .A(n1492), .B(n17567), .Z(n17575) );
  XNOR U16950 ( .A(n17565), .B(n17574), .Z(n17567) );
  XNOR U16951 ( .A(n17576), .B(n17577), .Z(n17565) );
  AND U16952 ( .A(n1496), .B(n17578), .Z(n17577) );
  XOR U16953 ( .A(p_input[1215]), .B(n17576), .Z(n17578) );
  XNOR U16954 ( .A(n17579), .B(n17580), .Z(n17576) );
  AND U16955 ( .A(n1500), .B(n17581), .Z(n17580) );
  XOR U16956 ( .A(n17582), .B(n17583), .Z(n17574) );
  AND U16957 ( .A(n1504), .B(n17573), .Z(n17583) );
  XNOR U16958 ( .A(n17584), .B(n17571), .Z(n17573) );
  XOR U16959 ( .A(n17585), .B(n17586), .Z(n17571) );
  AND U16960 ( .A(n1527), .B(n17587), .Z(n17586) );
  IV U16961 ( .A(n17582), .Z(n17584) );
  XOR U16962 ( .A(n17588), .B(n17589), .Z(n17582) );
  AND U16963 ( .A(n1511), .B(n17581), .Z(n17589) );
  XNOR U16964 ( .A(n17579), .B(n17588), .Z(n17581) );
  XNOR U16965 ( .A(n17590), .B(n17591), .Z(n17579) );
  AND U16966 ( .A(n1515), .B(n17592), .Z(n17591) );
  XOR U16967 ( .A(p_input[1231]), .B(n17590), .Z(n17592) );
  XNOR U16968 ( .A(n17593), .B(n17594), .Z(n17590) );
  AND U16969 ( .A(n1519), .B(n17595), .Z(n17594) );
  XOR U16970 ( .A(n17596), .B(n17597), .Z(n17588) );
  AND U16971 ( .A(n1523), .B(n17587), .Z(n17597) );
  XNOR U16972 ( .A(n17598), .B(n17585), .Z(n17587) );
  XOR U16973 ( .A(n17599), .B(n17600), .Z(n17585) );
  AND U16974 ( .A(n1546), .B(n17601), .Z(n17600) );
  IV U16975 ( .A(n17596), .Z(n17598) );
  XOR U16976 ( .A(n17602), .B(n17603), .Z(n17596) );
  AND U16977 ( .A(n1530), .B(n17595), .Z(n17603) );
  XNOR U16978 ( .A(n17593), .B(n17602), .Z(n17595) );
  XNOR U16979 ( .A(n17604), .B(n17605), .Z(n17593) );
  AND U16980 ( .A(n1534), .B(n17606), .Z(n17605) );
  XOR U16981 ( .A(p_input[1247]), .B(n17604), .Z(n17606) );
  XNOR U16982 ( .A(n17607), .B(n17608), .Z(n17604) );
  AND U16983 ( .A(n1538), .B(n17609), .Z(n17608) );
  XOR U16984 ( .A(n17610), .B(n17611), .Z(n17602) );
  AND U16985 ( .A(n1542), .B(n17601), .Z(n17611) );
  XNOR U16986 ( .A(n17612), .B(n17599), .Z(n17601) );
  XOR U16987 ( .A(n17613), .B(n17614), .Z(n17599) );
  AND U16988 ( .A(n1565), .B(n17615), .Z(n17614) );
  IV U16989 ( .A(n17610), .Z(n17612) );
  XOR U16990 ( .A(n17616), .B(n17617), .Z(n17610) );
  AND U16991 ( .A(n1549), .B(n17609), .Z(n17617) );
  XNOR U16992 ( .A(n17607), .B(n17616), .Z(n17609) );
  XNOR U16993 ( .A(n17618), .B(n17619), .Z(n17607) );
  AND U16994 ( .A(n1553), .B(n17620), .Z(n17619) );
  XOR U16995 ( .A(p_input[1263]), .B(n17618), .Z(n17620) );
  XNOR U16996 ( .A(n17621), .B(n17622), .Z(n17618) );
  AND U16997 ( .A(n1557), .B(n17623), .Z(n17622) );
  XOR U16998 ( .A(n17624), .B(n17625), .Z(n17616) );
  AND U16999 ( .A(n1561), .B(n17615), .Z(n17625) );
  XNOR U17000 ( .A(n17626), .B(n17613), .Z(n17615) );
  XOR U17001 ( .A(n17627), .B(n17628), .Z(n17613) );
  AND U17002 ( .A(n1584), .B(n17629), .Z(n17628) );
  IV U17003 ( .A(n17624), .Z(n17626) );
  XOR U17004 ( .A(n17630), .B(n17631), .Z(n17624) );
  AND U17005 ( .A(n1568), .B(n17623), .Z(n17631) );
  XNOR U17006 ( .A(n17621), .B(n17630), .Z(n17623) );
  XNOR U17007 ( .A(n17632), .B(n17633), .Z(n17621) );
  AND U17008 ( .A(n1572), .B(n17634), .Z(n17633) );
  XOR U17009 ( .A(p_input[1279]), .B(n17632), .Z(n17634) );
  XNOR U17010 ( .A(n17635), .B(n17636), .Z(n17632) );
  AND U17011 ( .A(n1576), .B(n17637), .Z(n17636) );
  XOR U17012 ( .A(n17638), .B(n17639), .Z(n17630) );
  AND U17013 ( .A(n1580), .B(n17629), .Z(n17639) );
  XNOR U17014 ( .A(n17640), .B(n17627), .Z(n17629) );
  XOR U17015 ( .A(n17641), .B(n17642), .Z(n17627) );
  AND U17016 ( .A(n1603), .B(n17643), .Z(n17642) );
  IV U17017 ( .A(n17638), .Z(n17640) );
  XOR U17018 ( .A(n17644), .B(n17645), .Z(n17638) );
  AND U17019 ( .A(n1587), .B(n17637), .Z(n17645) );
  XNOR U17020 ( .A(n17635), .B(n17644), .Z(n17637) );
  XNOR U17021 ( .A(n17646), .B(n17647), .Z(n17635) );
  AND U17022 ( .A(n1591), .B(n17648), .Z(n17647) );
  XOR U17023 ( .A(p_input[1295]), .B(n17646), .Z(n17648) );
  XNOR U17024 ( .A(n17649), .B(n17650), .Z(n17646) );
  AND U17025 ( .A(n1595), .B(n17651), .Z(n17650) );
  XOR U17026 ( .A(n17652), .B(n17653), .Z(n17644) );
  AND U17027 ( .A(n1599), .B(n17643), .Z(n17653) );
  XNOR U17028 ( .A(n17654), .B(n17641), .Z(n17643) );
  XOR U17029 ( .A(n17655), .B(n17656), .Z(n17641) );
  AND U17030 ( .A(n1622), .B(n17657), .Z(n17656) );
  IV U17031 ( .A(n17652), .Z(n17654) );
  XOR U17032 ( .A(n17658), .B(n17659), .Z(n17652) );
  AND U17033 ( .A(n1606), .B(n17651), .Z(n17659) );
  XNOR U17034 ( .A(n17649), .B(n17658), .Z(n17651) );
  XNOR U17035 ( .A(n17660), .B(n17661), .Z(n17649) );
  AND U17036 ( .A(n1610), .B(n17662), .Z(n17661) );
  XOR U17037 ( .A(p_input[1311]), .B(n17660), .Z(n17662) );
  XNOR U17038 ( .A(n17663), .B(n17664), .Z(n17660) );
  AND U17039 ( .A(n1614), .B(n17665), .Z(n17664) );
  XOR U17040 ( .A(n17666), .B(n17667), .Z(n17658) );
  AND U17041 ( .A(n1618), .B(n17657), .Z(n17667) );
  XNOR U17042 ( .A(n17668), .B(n17655), .Z(n17657) );
  XOR U17043 ( .A(n17669), .B(n17670), .Z(n17655) );
  AND U17044 ( .A(n1641), .B(n17671), .Z(n17670) );
  IV U17045 ( .A(n17666), .Z(n17668) );
  XOR U17046 ( .A(n17672), .B(n17673), .Z(n17666) );
  AND U17047 ( .A(n1625), .B(n17665), .Z(n17673) );
  XNOR U17048 ( .A(n17663), .B(n17672), .Z(n17665) );
  XNOR U17049 ( .A(n17674), .B(n17675), .Z(n17663) );
  AND U17050 ( .A(n1629), .B(n17676), .Z(n17675) );
  XOR U17051 ( .A(p_input[1327]), .B(n17674), .Z(n17676) );
  XNOR U17052 ( .A(n17677), .B(n17678), .Z(n17674) );
  AND U17053 ( .A(n1633), .B(n17679), .Z(n17678) );
  XOR U17054 ( .A(n17680), .B(n17681), .Z(n17672) );
  AND U17055 ( .A(n1637), .B(n17671), .Z(n17681) );
  XNOR U17056 ( .A(n17682), .B(n17669), .Z(n17671) );
  XOR U17057 ( .A(n17683), .B(n17684), .Z(n17669) );
  AND U17058 ( .A(n1660), .B(n17685), .Z(n17684) );
  IV U17059 ( .A(n17680), .Z(n17682) );
  XOR U17060 ( .A(n17686), .B(n17687), .Z(n17680) );
  AND U17061 ( .A(n1644), .B(n17679), .Z(n17687) );
  XNOR U17062 ( .A(n17677), .B(n17686), .Z(n17679) );
  XNOR U17063 ( .A(n17688), .B(n17689), .Z(n17677) );
  AND U17064 ( .A(n1648), .B(n17690), .Z(n17689) );
  XOR U17065 ( .A(p_input[1343]), .B(n17688), .Z(n17690) );
  XNOR U17066 ( .A(n17691), .B(n17692), .Z(n17688) );
  AND U17067 ( .A(n1652), .B(n17693), .Z(n17692) );
  XOR U17068 ( .A(n17694), .B(n17695), .Z(n17686) );
  AND U17069 ( .A(n1656), .B(n17685), .Z(n17695) );
  XNOR U17070 ( .A(n17696), .B(n17683), .Z(n17685) );
  XOR U17071 ( .A(n17697), .B(n17698), .Z(n17683) );
  AND U17072 ( .A(n1679), .B(n17699), .Z(n17698) );
  IV U17073 ( .A(n17694), .Z(n17696) );
  XOR U17074 ( .A(n17700), .B(n17701), .Z(n17694) );
  AND U17075 ( .A(n1663), .B(n17693), .Z(n17701) );
  XNOR U17076 ( .A(n17691), .B(n17700), .Z(n17693) );
  XNOR U17077 ( .A(n17702), .B(n17703), .Z(n17691) );
  AND U17078 ( .A(n1667), .B(n17704), .Z(n17703) );
  XOR U17079 ( .A(p_input[1359]), .B(n17702), .Z(n17704) );
  XNOR U17080 ( .A(n17705), .B(n17706), .Z(n17702) );
  AND U17081 ( .A(n1671), .B(n17707), .Z(n17706) );
  XOR U17082 ( .A(n17708), .B(n17709), .Z(n17700) );
  AND U17083 ( .A(n1675), .B(n17699), .Z(n17709) );
  XNOR U17084 ( .A(n17710), .B(n17697), .Z(n17699) );
  XOR U17085 ( .A(n17711), .B(n17712), .Z(n17697) );
  AND U17086 ( .A(n1698), .B(n17713), .Z(n17712) );
  IV U17087 ( .A(n17708), .Z(n17710) );
  XOR U17088 ( .A(n17714), .B(n17715), .Z(n17708) );
  AND U17089 ( .A(n1682), .B(n17707), .Z(n17715) );
  XNOR U17090 ( .A(n17705), .B(n17714), .Z(n17707) );
  XNOR U17091 ( .A(n17716), .B(n17717), .Z(n17705) );
  AND U17092 ( .A(n1686), .B(n17718), .Z(n17717) );
  XOR U17093 ( .A(p_input[1375]), .B(n17716), .Z(n17718) );
  XNOR U17094 ( .A(n17719), .B(n17720), .Z(n17716) );
  AND U17095 ( .A(n1690), .B(n17721), .Z(n17720) );
  XOR U17096 ( .A(n17722), .B(n17723), .Z(n17714) );
  AND U17097 ( .A(n1694), .B(n17713), .Z(n17723) );
  XNOR U17098 ( .A(n17724), .B(n17711), .Z(n17713) );
  XOR U17099 ( .A(n17725), .B(n17726), .Z(n17711) );
  AND U17100 ( .A(n1717), .B(n17727), .Z(n17726) );
  IV U17101 ( .A(n17722), .Z(n17724) );
  XOR U17102 ( .A(n17728), .B(n17729), .Z(n17722) );
  AND U17103 ( .A(n1701), .B(n17721), .Z(n17729) );
  XNOR U17104 ( .A(n17719), .B(n17728), .Z(n17721) );
  XNOR U17105 ( .A(n17730), .B(n17731), .Z(n17719) );
  AND U17106 ( .A(n1705), .B(n17732), .Z(n17731) );
  XOR U17107 ( .A(p_input[1391]), .B(n17730), .Z(n17732) );
  XNOR U17108 ( .A(n17733), .B(n17734), .Z(n17730) );
  AND U17109 ( .A(n1709), .B(n17735), .Z(n17734) );
  XOR U17110 ( .A(n17736), .B(n17737), .Z(n17728) );
  AND U17111 ( .A(n1713), .B(n17727), .Z(n17737) );
  XNOR U17112 ( .A(n17738), .B(n17725), .Z(n17727) );
  XOR U17113 ( .A(n17739), .B(n17740), .Z(n17725) );
  AND U17114 ( .A(n1736), .B(n17741), .Z(n17740) );
  IV U17115 ( .A(n17736), .Z(n17738) );
  XOR U17116 ( .A(n17742), .B(n17743), .Z(n17736) );
  AND U17117 ( .A(n1720), .B(n17735), .Z(n17743) );
  XNOR U17118 ( .A(n17733), .B(n17742), .Z(n17735) );
  XNOR U17119 ( .A(n17744), .B(n17745), .Z(n17733) );
  AND U17120 ( .A(n1724), .B(n17746), .Z(n17745) );
  XOR U17121 ( .A(p_input[1407]), .B(n17744), .Z(n17746) );
  XNOR U17122 ( .A(n17747), .B(n17748), .Z(n17744) );
  AND U17123 ( .A(n1728), .B(n17749), .Z(n17748) );
  XOR U17124 ( .A(n17750), .B(n17751), .Z(n17742) );
  AND U17125 ( .A(n1732), .B(n17741), .Z(n17751) );
  XNOR U17126 ( .A(n17752), .B(n17739), .Z(n17741) );
  XOR U17127 ( .A(n17753), .B(n17754), .Z(n17739) );
  AND U17128 ( .A(n1755), .B(n17755), .Z(n17754) );
  IV U17129 ( .A(n17750), .Z(n17752) );
  XOR U17130 ( .A(n17756), .B(n17757), .Z(n17750) );
  AND U17131 ( .A(n1739), .B(n17749), .Z(n17757) );
  XNOR U17132 ( .A(n17747), .B(n17756), .Z(n17749) );
  XNOR U17133 ( .A(n17758), .B(n17759), .Z(n17747) );
  AND U17134 ( .A(n1743), .B(n17760), .Z(n17759) );
  XOR U17135 ( .A(p_input[1423]), .B(n17758), .Z(n17760) );
  XNOR U17136 ( .A(n17761), .B(n17762), .Z(n17758) );
  AND U17137 ( .A(n1747), .B(n17763), .Z(n17762) );
  XOR U17138 ( .A(n17764), .B(n17765), .Z(n17756) );
  AND U17139 ( .A(n1751), .B(n17755), .Z(n17765) );
  XNOR U17140 ( .A(n17766), .B(n17753), .Z(n17755) );
  XOR U17141 ( .A(n17767), .B(n17768), .Z(n17753) );
  AND U17142 ( .A(n1774), .B(n17769), .Z(n17768) );
  IV U17143 ( .A(n17764), .Z(n17766) );
  XOR U17144 ( .A(n17770), .B(n17771), .Z(n17764) );
  AND U17145 ( .A(n1758), .B(n17763), .Z(n17771) );
  XNOR U17146 ( .A(n17761), .B(n17770), .Z(n17763) );
  XNOR U17147 ( .A(n17772), .B(n17773), .Z(n17761) );
  AND U17148 ( .A(n1762), .B(n17774), .Z(n17773) );
  XOR U17149 ( .A(p_input[1439]), .B(n17772), .Z(n17774) );
  XNOR U17150 ( .A(n17775), .B(n17776), .Z(n17772) );
  AND U17151 ( .A(n1766), .B(n17777), .Z(n17776) );
  XOR U17152 ( .A(n17778), .B(n17779), .Z(n17770) );
  AND U17153 ( .A(n1770), .B(n17769), .Z(n17779) );
  XNOR U17154 ( .A(n17780), .B(n17767), .Z(n17769) );
  XOR U17155 ( .A(n17781), .B(n17782), .Z(n17767) );
  AND U17156 ( .A(n1793), .B(n17783), .Z(n17782) );
  IV U17157 ( .A(n17778), .Z(n17780) );
  XOR U17158 ( .A(n17784), .B(n17785), .Z(n17778) );
  AND U17159 ( .A(n1777), .B(n17777), .Z(n17785) );
  XNOR U17160 ( .A(n17775), .B(n17784), .Z(n17777) );
  XNOR U17161 ( .A(n17786), .B(n17787), .Z(n17775) );
  AND U17162 ( .A(n1781), .B(n17788), .Z(n17787) );
  XOR U17163 ( .A(p_input[1455]), .B(n17786), .Z(n17788) );
  XNOR U17164 ( .A(n17789), .B(n17790), .Z(n17786) );
  AND U17165 ( .A(n1785), .B(n17791), .Z(n17790) );
  XOR U17166 ( .A(n17792), .B(n17793), .Z(n17784) );
  AND U17167 ( .A(n1789), .B(n17783), .Z(n17793) );
  XNOR U17168 ( .A(n17794), .B(n17781), .Z(n17783) );
  XOR U17169 ( .A(n17795), .B(n17796), .Z(n17781) );
  AND U17170 ( .A(n1812), .B(n17797), .Z(n17796) );
  IV U17171 ( .A(n17792), .Z(n17794) );
  XOR U17172 ( .A(n17798), .B(n17799), .Z(n17792) );
  AND U17173 ( .A(n1796), .B(n17791), .Z(n17799) );
  XNOR U17174 ( .A(n17789), .B(n17798), .Z(n17791) );
  XNOR U17175 ( .A(n17800), .B(n17801), .Z(n17789) );
  AND U17176 ( .A(n1800), .B(n17802), .Z(n17801) );
  XOR U17177 ( .A(p_input[1471]), .B(n17800), .Z(n17802) );
  XNOR U17178 ( .A(n17803), .B(n17804), .Z(n17800) );
  AND U17179 ( .A(n1804), .B(n17805), .Z(n17804) );
  XOR U17180 ( .A(n17806), .B(n17807), .Z(n17798) );
  AND U17181 ( .A(n1808), .B(n17797), .Z(n17807) );
  XNOR U17182 ( .A(n17808), .B(n17795), .Z(n17797) );
  XOR U17183 ( .A(n17809), .B(n17810), .Z(n17795) );
  AND U17184 ( .A(n1831), .B(n17811), .Z(n17810) );
  IV U17185 ( .A(n17806), .Z(n17808) );
  XOR U17186 ( .A(n17812), .B(n17813), .Z(n17806) );
  AND U17187 ( .A(n1815), .B(n17805), .Z(n17813) );
  XNOR U17188 ( .A(n17803), .B(n17812), .Z(n17805) );
  XNOR U17189 ( .A(n17814), .B(n17815), .Z(n17803) );
  AND U17190 ( .A(n1819), .B(n17816), .Z(n17815) );
  XOR U17191 ( .A(p_input[1487]), .B(n17814), .Z(n17816) );
  XNOR U17192 ( .A(n17817), .B(n17818), .Z(n17814) );
  AND U17193 ( .A(n1823), .B(n17819), .Z(n17818) );
  XOR U17194 ( .A(n17820), .B(n17821), .Z(n17812) );
  AND U17195 ( .A(n1827), .B(n17811), .Z(n17821) );
  XNOR U17196 ( .A(n17822), .B(n17809), .Z(n17811) );
  XOR U17197 ( .A(n17823), .B(n17824), .Z(n17809) );
  AND U17198 ( .A(n1850), .B(n17825), .Z(n17824) );
  IV U17199 ( .A(n17820), .Z(n17822) );
  XOR U17200 ( .A(n17826), .B(n17827), .Z(n17820) );
  AND U17201 ( .A(n1834), .B(n17819), .Z(n17827) );
  XNOR U17202 ( .A(n17817), .B(n17826), .Z(n17819) );
  XNOR U17203 ( .A(n17828), .B(n17829), .Z(n17817) );
  AND U17204 ( .A(n1838), .B(n17830), .Z(n17829) );
  XOR U17205 ( .A(p_input[1503]), .B(n17828), .Z(n17830) );
  XNOR U17206 ( .A(n17831), .B(n17832), .Z(n17828) );
  AND U17207 ( .A(n1842), .B(n17833), .Z(n17832) );
  XOR U17208 ( .A(n17834), .B(n17835), .Z(n17826) );
  AND U17209 ( .A(n1846), .B(n17825), .Z(n17835) );
  XNOR U17210 ( .A(n17836), .B(n17823), .Z(n17825) );
  XOR U17211 ( .A(n17837), .B(n17838), .Z(n17823) );
  AND U17212 ( .A(n1869), .B(n17839), .Z(n17838) );
  IV U17213 ( .A(n17834), .Z(n17836) );
  XOR U17214 ( .A(n17840), .B(n17841), .Z(n17834) );
  AND U17215 ( .A(n1853), .B(n17833), .Z(n17841) );
  XNOR U17216 ( .A(n17831), .B(n17840), .Z(n17833) );
  XNOR U17217 ( .A(n17842), .B(n17843), .Z(n17831) );
  AND U17218 ( .A(n1857), .B(n17844), .Z(n17843) );
  XOR U17219 ( .A(p_input[1519]), .B(n17842), .Z(n17844) );
  XNOR U17220 ( .A(n17845), .B(n17846), .Z(n17842) );
  AND U17221 ( .A(n1861), .B(n17847), .Z(n17846) );
  XOR U17222 ( .A(n17848), .B(n17849), .Z(n17840) );
  AND U17223 ( .A(n1865), .B(n17839), .Z(n17849) );
  XNOR U17224 ( .A(n17850), .B(n17837), .Z(n17839) );
  XOR U17225 ( .A(n17851), .B(n17852), .Z(n17837) );
  AND U17226 ( .A(n1888), .B(n17853), .Z(n17852) );
  IV U17227 ( .A(n17848), .Z(n17850) );
  XOR U17228 ( .A(n17854), .B(n17855), .Z(n17848) );
  AND U17229 ( .A(n1872), .B(n17847), .Z(n17855) );
  XNOR U17230 ( .A(n17845), .B(n17854), .Z(n17847) );
  XNOR U17231 ( .A(n17856), .B(n17857), .Z(n17845) );
  AND U17232 ( .A(n1876), .B(n17858), .Z(n17857) );
  XOR U17233 ( .A(p_input[1535]), .B(n17856), .Z(n17858) );
  XNOR U17234 ( .A(n17859), .B(n17860), .Z(n17856) );
  AND U17235 ( .A(n1880), .B(n17861), .Z(n17860) );
  XOR U17236 ( .A(n17862), .B(n17863), .Z(n17854) );
  AND U17237 ( .A(n1884), .B(n17853), .Z(n17863) );
  XNOR U17238 ( .A(n17864), .B(n17851), .Z(n17853) );
  XOR U17239 ( .A(n17865), .B(n17866), .Z(n17851) );
  AND U17240 ( .A(n1907), .B(n17867), .Z(n17866) );
  IV U17241 ( .A(n17862), .Z(n17864) );
  XOR U17242 ( .A(n17868), .B(n17869), .Z(n17862) );
  AND U17243 ( .A(n1891), .B(n17861), .Z(n17869) );
  XNOR U17244 ( .A(n17859), .B(n17868), .Z(n17861) );
  XNOR U17245 ( .A(n17870), .B(n17871), .Z(n17859) );
  AND U17246 ( .A(n1895), .B(n17872), .Z(n17871) );
  XOR U17247 ( .A(p_input[1551]), .B(n17870), .Z(n17872) );
  XNOR U17248 ( .A(n17873), .B(n17874), .Z(n17870) );
  AND U17249 ( .A(n1899), .B(n17875), .Z(n17874) );
  XOR U17250 ( .A(n17876), .B(n17877), .Z(n17868) );
  AND U17251 ( .A(n1903), .B(n17867), .Z(n17877) );
  XNOR U17252 ( .A(n17878), .B(n17865), .Z(n17867) );
  XOR U17253 ( .A(n17879), .B(n17880), .Z(n17865) );
  AND U17254 ( .A(n1926), .B(n17881), .Z(n17880) );
  IV U17255 ( .A(n17876), .Z(n17878) );
  XOR U17256 ( .A(n17882), .B(n17883), .Z(n17876) );
  AND U17257 ( .A(n1910), .B(n17875), .Z(n17883) );
  XNOR U17258 ( .A(n17873), .B(n17882), .Z(n17875) );
  XNOR U17259 ( .A(n17884), .B(n17885), .Z(n17873) );
  AND U17260 ( .A(n1914), .B(n17886), .Z(n17885) );
  XOR U17261 ( .A(p_input[1567]), .B(n17884), .Z(n17886) );
  XNOR U17262 ( .A(n17887), .B(n17888), .Z(n17884) );
  AND U17263 ( .A(n1918), .B(n17889), .Z(n17888) );
  XOR U17264 ( .A(n17890), .B(n17891), .Z(n17882) );
  AND U17265 ( .A(n1922), .B(n17881), .Z(n17891) );
  XNOR U17266 ( .A(n17892), .B(n17879), .Z(n17881) );
  XOR U17267 ( .A(n17893), .B(n17894), .Z(n17879) );
  AND U17268 ( .A(n1945), .B(n17895), .Z(n17894) );
  IV U17269 ( .A(n17890), .Z(n17892) );
  XOR U17270 ( .A(n17896), .B(n17897), .Z(n17890) );
  AND U17271 ( .A(n1929), .B(n17889), .Z(n17897) );
  XNOR U17272 ( .A(n17887), .B(n17896), .Z(n17889) );
  XNOR U17273 ( .A(n17898), .B(n17899), .Z(n17887) );
  AND U17274 ( .A(n1933), .B(n17900), .Z(n17899) );
  XOR U17275 ( .A(p_input[1583]), .B(n17898), .Z(n17900) );
  XNOR U17276 ( .A(n17901), .B(n17902), .Z(n17898) );
  AND U17277 ( .A(n1937), .B(n17903), .Z(n17902) );
  XOR U17278 ( .A(n17904), .B(n17905), .Z(n17896) );
  AND U17279 ( .A(n1941), .B(n17895), .Z(n17905) );
  XNOR U17280 ( .A(n17906), .B(n17893), .Z(n17895) );
  XOR U17281 ( .A(n17907), .B(n17908), .Z(n17893) );
  AND U17282 ( .A(n1964), .B(n17909), .Z(n17908) );
  IV U17283 ( .A(n17904), .Z(n17906) );
  XOR U17284 ( .A(n17910), .B(n17911), .Z(n17904) );
  AND U17285 ( .A(n1948), .B(n17903), .Z(n17911) );
  XNOR U17286 ( .A(n17901), .B(n17910), .Z(n17903) );
  XNOR U17287 ( .A(n17912), .B(n17913), .Z(n17901) );
  AND U17288 ( .A(n1952), .B(n17914), .Z(n17913) );
  XOR U17289 ( .A(p_input[1599]), .B(n17912), .Z(n17914) );
  XNOR U17290 ( .A(n17915), .B(n17916), .Z(n17912) );
  AND U17291 ( .A(n1956), .B(n17917), .Z(n17916) );
  XOR U17292 ( .A(n17918), .B(n17919), .Z(n17910) );
  AND U17293 ( .A(n1960), .B(n17909), .Z(n17919) );
  XNOR U17294 ( .A(n17920), .B(n17907), .Z(n17909) );
  XOR U17295 ( .A(n17921), .B(n17922), .Z(n17907) );
  AND U17296 ( .A(n1983), .B(n17923), .Z(n17922) );
  IV U17297 ( .A(n17918), .Z(n17920) );
  XOR U17298 ( .A(n17924), .B(n17925), .Z(n17918) );
  AND U17299 ( .A(n1967), .B(n17917), .Z(n17925) );
  XNOR U17300 ( .A(n17915), .B(n17924), .Z(n17917) );
  XNOR U17301 ( .A(n17926), .B(n17927), .Z(n17915) );
  AND U17302 ( .A(n1971), .B(n17928), .Z(n17927) );
  XOR U17303 ( .A(p_input[1615]), .B(n17926), .Z(n17928) );
  XNOR U17304 ( .A(n17929), .B(n17930), .Z(n17926) );
  AND U17305 ( .A(n1975), .B(n17931), .Z(n17930) );
  XOR U17306 ( .A(n17932), .B(n17933), .Z(n17924) );
  AND U17307 ( .A(n1979), .B(n17923), .Z(n17933) );
  XNOR U17308 ( .A(n17934), .B(n17921), .Z(n17923) );
  XOR U17309 ( .A(n17935), .B(n17936), .Z(n17921) );
  AND U17310 ( .A(n2002), .B(n17937), .Z(n17936) );
  IV U17311 ( .A(n17932), .Z(n17934) );
  XOR U17312 ( .A(n17938), .B(n17939), .Z(n17932) );
  AND U17313 ( .A(n1986), .B(n17931), .Z(n17939) );
  XNOR U17314 ( .A(n17929), .B(n17938), .Z(n17931) );
  XNOR U17315 ( .A(n17940), .B(n17941), .Z(n17929) );
  AND U17316 ( .A(n1990), .B(n17942), .Z(n17941) );
  XOR U17317 ( .A(p_input[1631]), .B(n17940), .Z(n17942) );
  XNOR U17318 ( .A(n17943), .B(n17944), .Z(n17940) );
  AND U17319 ( .A(n1994), .B(n17945), .Z(n17944) );
  XOR U17320 ( .A(n17946), .B(n17947), .Z(n17938) );
  AND U17321 ( .A(n1998), .B(n17937), .Z(n17947) );
  XNOR U17322 ( .A(n17948), .B(n17935), .Z(n17937) );
  XOR U17323 ( .A(n17949), .B(n17950), .Z(n17935) );
  AND U17324 ( .A(n2021), .B(n17951), .Z(n17950) );
  IV U17325 ( .A(n17946), .Z(n17948) );
  XOR U17326 ( .A(n17952), .B(n17953), .Z(n17946) );
  AND U17327 ( .A(n2005), .B(n17945), .Z(n17953) );
  XNOR U17328 ( .A(n17943), .B(n17952), .Z(n17945) );
  XNOR U17329 ( .A(n17954), .B(n17955), .Z(n17943) );
  AND U17330 ( .A(n2009), .B(n17956), .Z(n17955) );
  XOR U17331 ( .A(p_input[1647]), .B(n17954), .Z(n17956) );
  XNOR U17332 ( .A(n17957), .B(n17958), .Z(n17954) );
  AND U17333 ( .A(n2013), .B(n17959), .Z(n17958) );
  XOR U17334 ( .A(n17960), .B(n17961), .Z(n17952) );
  AND U17335 ( .A(n2017), .B(n17951), .Z(n17961) );
  XNOR U17336 ( .A(n17962), .B(n17949), .Z(n17951) );
  XOR U17337 ( .A(n17963), .B(n17964), .Z(n17949) );
  AND U17338 ( .A(n2040), .B(n17965), .Z(n17964) );
  IV U17339 ( .A(n17960), .Z(n17962) );
  XOR U17340 ( .A(n17966), .B(n17967), .Z(n17960) );
  AND U17341 ( .A(n2024), .B(n17959), .Z(n17967) );
  XNOR U17342 ( .A(n17957), .B(n17966), .Z(n17959) );
  XNOR U17343 ( .A(n17968), .B(n17969), .Z(n17957) );
  AND U17344 ( .A(n2028), .B(n17970), .Z(n17969) );
  XOR U17345 ( .A(p_input[1663]), .B(n17968), .Z(n17970) );
  XNOR U17346 ( .A(n17971), .B(n17972), .Z(n17968) );
  AND U17347 ( .A(n2032), .B(n17973), .Z(n17972) );
  XOR U17348 ( .A(n17974), .B(n17975), .Z(n17966) );
  AND U17349 ( .A(n2036), .B(n17965), .Z(n17975) );
  XNOR U17350 ( .A(n17976), .B(n17963), .Z(n17965) );
  XOR U17351 ( .A(n17977), .B(n17978), .Z(n17963) );
  AND U17352 ( .A(n2059), .B(n17979), .Z(n17978) );
  IV U17353 ( .A(n17974), .Z(n17976) );
  XOR U17354 ( .A(n17980), .B(n17981), .Z(n17974) );
  AND U17355 ( .A(n2043), .B(n17973), .Z(n17981) );
  XNOR U17356 ( .A(n17971), .B(n17980), .Z(n17973) );
  XNOR U17357 ( .A(n17982), .B(n17983), .Z(n17971) );
  AND U17358 ( .A(n2047), .B(n17984), .Z(n17983) );
  XOR U17359 ( .A(p_input[1679]), .B(n17982), .Z(n17984) );
  XNOR U17360 ( .A(n17985), .B(n17986), .Z(n17982) );
  AND U17361 ( .A(n2051), .B(n17987), .Z(n17986) );
  XOR U17362 ( .A(n17988), .B(n17989), .Z(n17980) );
  AND U17363 ( .A(n2055), .B(n17979), .Z(n17989) );
  XNOR U17364 ( .A(n17990), .B(n17977), .Z(n17979) );
  XOR U17365 ( .A(n17991), .B(n17992), .Z(n17977) );
  AND U17366 ( .A(n2078), .B(n17993), .Z(n17992) );
  IV U17367 ( .A(n17988), .Z(n17990) );
  XOR U17368 ( .A(n17994), .B(n17995), .Z(n17988) );
  AND U17369 ( .A(n2062), .B(n17987), .Z(n17995) );
  XNOR U17370 ( .A(n17985), .B(n17994), .Z(n17987) );
  XNOR U17371 ( .A(n17996), .B(n17997), .Z(n17985) );
  AND U17372 ( .A(n2066), .B(n17998), .Z(n17997) );
  XOR U17373 ( .A(p_input[1695]), .B(n17996), .Z(n17998) );
  XNOR U17374 ( .A(n17999), .B(n18000), .Z(n17996) );
  AND U17375 ( .A(n2070), .B(n18001), .Z(n18000) );
  XOR U17376 ( .A(n18002), .B(n18003), .Z(n17994) );
  AND U17377 ( .A(n2074), .B(n17993), .Z(n18003) );
  XNOR U17378 ( .A(n18004), .B(n17991), .Z(n17993) );
  XOR U17379 ( .A(n18005), .B(n18006), .Z(n17991) );
  AND U17380 ( .A(n2097), .B(n18007), .Z(n18006) );
  IV U17381 ( .A(n18002), .Z(n18004) );
  XOR U17382 ( .A(n18008), .B(n18009), .Z(n18002) );
  AND U17383 ( .A(n2081), .B(n18001), .Z(n18009) );
  XNOR U17384 ( .A(n17999), .B(n18008), .Z(n18001) );
  XNOR U17385 ( .A(n18010), .B(n18011), .Z(n17999) );
  AND U17386 ( .A(n2085), .B(n18012), .Z(n18011) );
  XOR U17387 ( .A(p_input[1711]), .B(n18010), .Z(n18012) );
  XNOR U17388 ( .A(n18013), .B(n18014), .Z(n18010) );
  AND U17389 ( .A(n2089), .B(n18015), .Z(n18014) );
  XOR U17390 ( .A(n18016), .B(n18017), .Z(n18008) );
  AND U17391 ( .A(n2093), .B(n18007), .Z(n18017) );
  XNOR U17392 ( .A(n18018), .B(n18005), .Z(n18007) );
  XOR U17393 ( .A(n18019), .B(n18020), .Z(n18005) );
  AND U17394 ( .A(n2116), .B(n18021), .Z(n18020) );
  IV U17395 ( .A(n18016), .Z(n18018) );
  XOR U17396 ( .A(n18022), .B(n18023), .Z(n18016) );
  AND U17397 ( .A(n2100), .B(n18015), .Z(n18023) );
  XNOR U17398 ( .A(n18013), .B(n18022), .Z(n18015) );
  XNOR U17399 ( .A(n18024), .B(n18025), .Z(n18013) );
  AND U17400 ( .A(n2104), .B(n18026), .Z(n18025) );
  XOR U17401 ( .A(p_input[1727]), .B(n18024), .Z(n18026) );
  XNOR U17402 ( .A(n18027), .B(n18028), .Z(n18024) );
  AND U17403 ( .A(n2108), .B(n18029), .Z(n18028) );
  XOR U17404 ( .A(n18030), .B(n18031), .Z(n18022) );
  AND U17405 ( .A(n2112), .B(n18021), .Z(n18031) );
  XNOR U17406 ( .A(n18032), .B(n18019), .Z(n18021) );
  XOR U17407 ( .A(n18033), .B(n18034), .Z(n18019) );
  AND U17408 ( .A(n2135), .B(n18035), .Z(n18034) );
  IV U17409 ( .A(n18030), .Z(n18032) );
  XOR U17410 ( .A(n18036), .B(n18037), .Z(n18030) );
  AND U17411 ( .A(n2119), .B(n18029), .Z(n18037) );
  XNOR U17412 ( .A(n18027), .B(n18036), .Z(n18029) );
  XNOR U17413 ( .A(n18038), .B(n18039), .Z(n18027) );
  AND U17414 ( .A(n2123), .B(n18040), .Z(n18039) );
  XOR U17415 ( .A(p_input[1743]), .B(n18038), .Z(n18040) );
  XNOR U17416 ( .A(n18041), .B(n18042), .Z(n18038) );
  AND U17417 ( .A(n2127), .B(n18043), .Z(n18042) );
  XOR U17418 ( .A(n18044), .B(n18045), .Z(n18036) );
  AND U17419 ( .A(n2131), .B(n18035), .Z(n18045) );
  XNOR U17420 ( .A(n18046), .B(n18033), .Z(n18035) );
  XOR U17421 ( .A(n18047), .B(n18048), .Z(n18033) );
  AND U17422 ( .A(n2154), .B(n18049), .Z(n18048) );
  IV U17423 ( .A(n18044), .Z(n18046) );
  XOR U17424 ( .A(n18050), .B(n18051), .Z(n18044) );
  AND U17425 ( .A(n2138), .B(n18043), .Z(n18051) );
  XNOR U17426 ( .A(n18041), .B(n18050), .Z(n18043) );
  XNOR U17427 ( .A(n18052), .B(n18053), .Z(n18041) );
  AND U17428 ( .A(n2142), .B(n18054), .Z(n18053) );
  XOR U17429 ( .A(p_input[1759]), .B(n18052), .Z(n18054) );
  XNOR U17430 ( .A(n18055), .B(n18056), .Z(n18052) );
  AND U17431 ( .A(n2146), .B(n18057), .Z(n18056) );
  XOR U17432 ( .A(n18058), .B(n18059), .Z(n18050) );
  AND U17433 ( .A(n2150), .B(n18049), .Z(n18059) );
  XNOR U17434 ( .A(n18060), .B(n18047), .Z(n18049) );
  XOR U17435 ( .A(n18061), .B(n18062), .Z(n18047) );
  AND U17436 ( .A(n2173), .B(n18063), .Z(n18062) );
  IV U17437 ( .A(n18058), .Z(n18060) );
  XOR U17438 ( .A(n18064), .B(n18065), .Z(n18058) );
  AND U17439 ( .A(n2157), .B(n18057), .Z(n18065) );
  XNOR U17440 ( .A(n18055), .B(n18064), .Z(n18057) );
  XNOR U17441 ( .A(n18066), .B(n18067), .Z(n18055) );
  AND U17442 ( .A(n2161), .B(n18068), .Z(n18067) );
  XOR U17443 ( .A(p_input[1775]), .B(n18066), .Z(n18068) );
  XNOR U17444 ( .A(n18069), .B(n18070), .Z(n18066) );
  AND U17445 ( .A(n2165), .B(n18071), .Z(n18070) );
  XOR U17446 ( .A(n18072), .B(n18073), .Z(n18064) );
  AND U17447 ( .A(n2169), .B(n18063), .Z(n18073) );
  XNOR U17448 ( .A(n18074), .B(n18061), .Z(n18063) );
  XOR U17449 ( .A(n18075), .B(n18076), .Z(n18061) );
  AND U17450 ( .A(n2192), .B(n18077), .Z(n18076) );
  IV U17451 ( .A(n18072), .Z(n18074) );
  XOR U17452 ( .A(n18078), .B(n18079), .Z(n18072) );
  AND U17453 ( .A(n2176), .B(n18071), .Z(n18079) );
  XNOR U17454 ( .A(n18069), .B(n18078), .Z(n18071) );
  XNOR U17455 ( .A(n18080), .B(n18081), .Z(n18069) );
  AND U17456 ( .A(n2180), .B(n18082), .Z(n18081) );
  XOR U17457 ( .A(p_input[1791]), .B(n18080), .Z(n18082) );
  XNOR U17458 ( .A(n18083), .B(n18084), .Z(n18080) );
  AND U17459 ( .A(n2184), .B(n18085), .Z(n18084) );
  XOR U17460 ( .A(n18086), .B(n18087), .Z(n18078) );
  AND U17461 ( .A(n2188), .B(n18077), .Z(n18087) );
  XNOR U17462 ( .A(n18088), .B(n18075), .Z(n18077) );
  XOR U17463 ( .A(n18089), .B(n18090), .Z(n18075) );
  AND U17464 ( .A(n2211), .B(n18091), .Z(n18090) );
  IV U17465 ( .A(n18086), .Z(n18088) );
  XOR U17466 ( .A(n18092), .B(n18093), .Z(n18086) );
  AND U17467 ( .A(n2195), .B(n18085), .Z(n18093) );
  XNOR U17468 ( .A(n18083), .B(n18092), .Z(n18085) );
  XNOR U17469 ( .A(n18094), .B(n18095), .Z(n18083) );
  AND U17470 ( .A(n2199), .B(n18096), .Z(n18095) );
  XOR U17471 ( .A(p_input[1807]), .B(n18094), .Z(n18096) );
  XNOR U17472 ( .A(n18097), .B(n18098), .Z(n18094) );
  AND U17473 ( .A(n2203), .B(n18099), .Z(n18098) );
  XOR U17474 ( .A(n18100), .B(n18101), .Z(n18092) );
  AND U17475 ( .A(n2207), .B(n18091), .Z(n18101) );
  XNOR U17476 ( .A(n18102), .B(n18089), .Z(n18091) );
  XOR U17477 ( .A(n18103), .B(n18104), .Z(n18089) );
  AND U17478 ( .A(n2230), .B(n18105), .Z(n18104) );
  IV U17479 ( .A(n18100), .Z(n18102) );
  XOR U17480 ( .A(n18106), .B(n18107), .Z(n18100) );
  AND U17481 ( .A(n2214), .B(n18099), .Z(n18107) );
  XNOR U17482 ( .A(n18097), .B(n18106), .Z(n18099) );
  XNOR U17483 ( .A(n18108), .B(n18109), .Z(n18097) );
  AND U17484 ( .A(n2218), .B(n18110), .Z(n18109) );
  XOR U17485 ( .A(p_input[1823]), .B(n18108), .Z(n18110) );
  XNOR U17486 ( .A(n18111), .B(n18112), .Z(n18108) );
  AND U17487 ( .A(n2222), .B(n18113), .Z(n18112) );
  XOR U17488 ( .A(n18114), .B(n18115), .Z(n18106) );
  AND U17489 ( .A(n2226), .B(n18105), .Z(n18115) );
  XNOR U17490 ( .A(n18116), .B(n18103), .Z(n18105) );
  XOR U17491 ( .A(n18117), .B(n18118), .Z(n18103) );
  AND U17492 ( .A(n2249), .B(n18119), .Z(n18118) );
  IV U17493 ( .A(n18114), .Z(n18116) );
  XOR U17494 ( .A(n18120), .B(n18121), .Z(n18114) );
  AND U17495 ( .A(n2233), .B(n18113), .Z(n18121) );
  XNOR U17496 ( .A(n18111), .B(n18120), .Z(n18113) );
  XNOR U17497 ( .A(n18122), .B(n18123), .Z(n18111) );
  AND U17498 ( .A(n2237), .B(n18124), .Z(n18123) );
  XOR U17499 ( .A(p_input[1839]), .B(n18122), .Z(n18124) );
  XNOR U17500 ( .A(n18125), .B(n18126), .Z(n18122) );
  AND U17501 ( .A(n2241), .B(n18127), .Z(n18126) );
  XOR U17502 ( .A(n18128), .B(n18129), .Z(n18120) );
  AND U17503 ( .A(n2245), .B(n18119), .Z(n18129) );
  XNOR U17504 ( .A(n18130), .B(n18117), .Z(n18119) );
  XOR U17505 ( .A(n18131), .B(n18132), .Z(n18117) );
  AND U17506 ( .A(n2268), .B(n18133), .Z(n18132) );
  IV U17507 ( .A(n18128), .Z(n18130) );
  XOR U17508 ( .A(n18134), .B(n18135), .Z(n18128) );
  AND U17509 ( .A(n2252), .B(n18127), .Z(n18135) );
  XNOR U17510 ( .A(n18125), .B(n18134), .Z(n18127) );
  XNOR U17511 ( .A(n18136), .B(n18137), .Z(n18125) );
  AND U17512 ( .A(n2256), .B(n18138), .Z(n18137) );
  XOR U17513 ( .A(p_input[1855]), .B(n18136), .Z(n18138) );
  XNOR U17514 ( .A(n18139), .B(n18140), .Z(n18136) );
  AND U17515 ( .A(n2260), .B(n18141), .Z(n18140) );
  XOR U17516 ( .A(n18142), .B(n18143), .Z(n18134) );
  AND U17517 ( .A(n2264), .B(n18133), .Z(n18143) );
  XNOR U17518 ( .A(n18144), .B(n18131), .Z(n18133) );
  XOR U17519 ( .A(n18145), .B(n18146), .Z(n18131) );
  AND U17520 ( .A(n2287), .B(n18147), .Z(n18146) );
  IV U17521 ( .A(n18142), .Z(n18144) );
  XOR U17522 ( .A(n18148), .B(n18149), .Z(n18142) );
  AND U17523 ( .A(n2271), .B(n18141), .Z(n18149) );
  XNOR U17524 ( .A(n18139), .B(n18148), .Z(n18141) );
  XNOR U17525 ( .A(n18150), .B(n18151), .Z(n18139) );
  AND U17526 ( .A(n2275), .B(n18152), .Z(n18151) );
  XOR U17527 ( .A(p_input[1871]), .B(n18150), .Z(n18152) );
  XNOR U17528 ( .A(n18153), .B(n18154), .Z(n18150) );
  AND U17529 ( .A(n2279), .B(n18155), .Z(n18154) );
  XOR U17530 ( .A(n18156), .B(n18157), .Z(n18148) );
  AND U17531 ( .A(n2283), .B(n18147), .Z(n18157) );
  XNOR U17532 ( .A(n18158), .B(n18145), .Z(n18147) );
  XOR U17533 ( .A(n18159), .B(n18160), .Z(n18145) );
  AND U17534 ( .A(n2306), .B(n18161), .Z(n18160) );
  IV U17535 ( .A(n18156), .Z(n18158) );
  XOR U17536 ( .A(n18162), .B(n18163), .Z(n18156) );
  AND U17537 ( .A(n2290), .B(n18155), .Z(n18163) );
  XNOR U17538 ( .A(n18153), .B(n18162), .Z(n18155) );
  XNOR U17539 ( .A(n18164), .B(n18165), .Z(n18153) );
  AND U17540 ( .A(n2294), .B(n18166), .Z(n18165) );
  XOR U17541 ( .A(p_input[1887]), .B(n18164), .Z(n18166) );
  XNOR U17542 ( .A(n18167), .B(n18168), .Z(n18164) );
  AND U17543 ( .A(n2298), .B(n18169), .Z(n18168) );
  XOR U17544 ( .A(n18170), .B(n18171), .Z(n18162) );
  AND U17545 ( .A(n2302), .B(n18161), .Z(n18171) );
  XNOR U17546 ( .A(n18172), .B(n18159), .Z(n18161) );
  XOR U17547 ( .A(n18173), .B(n18174), .Z(n18159) );
  AND U17548 ( .A(n2325), .B(n18175), .Z(n18174) );
  IV U17549 ( .A(n18170), .Z(n18172) );
  XOR U17550 ( .A(n18176), .B(n18177), .Z(n18170) );
  AND U17551 ( .A(n2309), .B(n18169), .Z(n18177) );
  XNOR U17552 ( .A(n18167), .B(n18176), .Z(n18169) );
  XNOR U17553 ( .A(n18178), .B(n18179), .Z(n18167) );
  AND U17554 ( .A(n2313), .B(n18180), .Z(n18179) );
  XOR U17555 ( .A(p_input[1903]), .B(n18178), .Z(n18180) );
  XNOR U17556 ( .A(n18181), .B(n18182), .Z(n18178) );
  AND U17557 ( .A(n2317), .B(n18183), .Z(n18182) );
  XOR U17558 ( .A(n18184), .B(n18185), .Z(n18176) );
  AND U17559 ( .A(n2321), .B(n18175), .Z(n18185) );
  XNOR U17560 ( .A(n18186), .B(n18173), .Z(n18175) );
  XOR U17561 ( .A(n18187), .B(n18188), .Z(n18173) );
  AND U17562 ( .A(n2344), .B(n18189), .Z(n18188) );
  IV U17563 ( .A(n18184), .Z(n18186) );
  XOR U17564 ( .A(n18190), .B(n18191), .Z(n18184) );
  AND U17565 ( .A(n2328), .B(n18183), .Z(n18191) );
  XNOR U17566 ( .A(n18181), .B(n18190), .Z(n18183) );
  XNOR U17567 ( .A(n18192), .B(n18193), .Z(n18181) );
  AND U17568 ( .A(n2332), .B(n18194), .Z(n18193) );
  XOR U17569 ( .A(p_input[1919]), .B(n18192), .Z(n18194) );
  XNOR U17570 ( .A(n18195), .B(n18196), .Z(n18192) );
  AND U17571 ( .A(n2336), .B(n18197), .Z(n18196) );
  XOR U17572 ( .A(n18198), .B(n18199), .Z(n18190) );
  AND U17573 ( .A(n2340), .B(n18189), .Z(n18199) );
  XNOR U17574 ( .A(n18200), .B(n18187), .Z(n18189) );
  XOR U17575 ( .A(n18201), .B(n18202), .Z(n18187) );
  AND U17576 ( .A(n2363), .B(n18203), .Z(n18202) );
  IV U17577 ( .A(n18198), .Z(n18200) );
  XOR U17578 ( .A(n18204), .B(n18205), .Z(n18198) );
  AND U17579 ( .A(n2347), .B(n18197), .Z(n18205) );
  XNOR U17580 ( .A(n18195), .B(n18204), .Z(n18197) );
  XNOR U17581 ( .A(n18206), .B(n18207), .Z(n18195) );
  AND U17582 ( .A(n2351), .B(n18208), .Z(n18207) );
  XOR U17583 ( .A(p_input[1935]), .B(n18206), .Z(n18208) );
  XNOR U17584 ( .A(n18209), .B(n18210), .Z(n18206) );
  AND U17585 ( .A(n2355), .B(n18211), .Z(n18210) );
  XOR U17586 ( .A(n18212), .B(n18213), .Z(n18204) );
  AND U17587 ( .A(n2359), .B(n18203), .Z(n18213) );
  XNOR U17588 ( .A(n18214), .B(n18201), .Z(n18203) );
  XOR U17589 ( .A(n18215), .B(n18216), .Z(n18201) );
  AND U17590 ( .A(n2382), .B(n18217), .Z(n18216) );
  IV U17591 ( .A(n18212), .Z(n18214) );
  XOR U17592 ( .A(n18218), .B(n18219), .Z(n18212) );
  AND U17593 ( .A(n2366), .B(n18211), .Z(n18219) );
  XNOR U17594 ( .A(n18209), .B(n18218), .Z(n18211) );
  XNOR U17595 ( .A(n18220), .B(n18221), .Z(n18209) );
  AND U17596 ( .A(n2370), .B(n18222), .Z(n18221) );
  XOR U17597 ( .A(p_input[1951]), .B(n18220), .Z(n18222) );
  XNOR U17598 ( .A(n18223), .B(n18224), .Z(n18220) );
  AND U17599 ( .A(n2374), .B(n18225), .Z(n18224) );
  XOR U17600 ( .A(n18226), .B(n18227), .Z(n18218) );
  AND U17601 ( .A(n2378), .B(n18217), .Z(n18227) );
  XNOR U17602 ( .A(n18228), .B(n18215), .Z(n18217) );
  XOR U17603 ( .A(n18229), .B(n18230), .Z(n18215) );
  AND U17604 ( .A(n2401), .B(n18231), .Z(n18230) );
  IV U17605 ( .A(n18226), .Z(n18228) );
  XOR U17606 ( .A(n18232), .B(n18233), .Z(n18226) );
  AND U17607 ( .A(n2385), .B(n18225), .Z(n18233) );
  XNOR U17608 ( .A(n18223), .B(n18232), .Z(n18225) );
  XNOR U17609 ( .A(n18234), .B(n18235), .Z(n18223) );
  AND U17610 ( .A(n2389), .B(n18236), .Z(n18235) );
  XOR U17611 ( .A(p_input[1967]), .B(n18234), .Z(n18236) );
  XNOR U17612 ( .A(n18237), .B(n18238), .Z(n18234) );
  AND U17613 ( .A(n2393), .B(n18239), .Z(n18238) );
  XOR U17614 ( .A(n18240), .B(n18241), .Z(n18232) );
  AND U17615 ( .A(n2397), .B(n18231), .Z(n18241) );
  XNOR U17616 ( .A(n18242), .B(n18229), .Z(n18231) );
  XOR U17617 ( .A(n18243), .B(n18244), .Z(n18229) );
  AND U17618 ( .A(n2420), .B(n18245), .Z(n18244) );
  IV U17619 ( .A(n18240), .Z(n18242) );
  XOR U17620 ( .A(n18246), .B(n18247), .Z(n18240) );
  AND U17621 ( .A(n2404), .B(n18239), .Z(n18247) );
  XNOR U17622 ( .A(n18237), .B(n18246), .Z(n18239) );
  XNOR U17623 ( .A(n18248), .B(n18249), .Z(n18237) );
  AND U17624 ( .A(n2408), .B(n18250), .Z(n18249) );
  XOR U17625 ( .A(p_input[1983]), .B(n18248), .Z(n18250) );
  XNOR U17626 ( .A(n18251), .B(n18252), .Z(n18248) );
  AND U17627 ( .A(n2412), .B(n18253), .Z(n18252) );
  XOR U17628 ( .A(n18254), .B(n18255), .Z(n18246) );
  AND U17629 ( .A(n2416), .B(n18245), .Z(n18255) );
  XNOR U17630 ( .A(n18256), .B(n18243), .Z(n18245) );
  XOR U17631 ( .A(n18257), .B(n18258), .Z(n18243) );
  AND U17632 ( .A(n2438), .B(n18259), .Z(n18258) );
  IV U17633 ( .A(n18254), .Z(n18256) );
  XOR U17634 ( .A(n18260), .B(n18261), .Z(n18254) );
  AND U17635 ( .A(n2423), .B(n18253), .Z(n18261) );
  XNOR U17636 ( .A(n18251), .B(n18260), .Z(n18253) );
  XNOR U17637 ( .A(n18262), .B(n18263), .Z(n18251) );
  AND U17638 ( .A(n2427), .B(n18264), .Z(n18263) );
  XOR U17639 ( .A(p_input[1999]), .B(n18262), .Z(n18264) );
  XOR U17640 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n18265), 
        .Z(n18262) );
  AND U17641 ( .A(n2430), .B(n18266), .Z(n18265) );
  XOR U17642 ( .A(n18267), .B(n18268), .Z(n18260) );
  AND U17643 ( .A(n2434), .B(n18259), .Z(n18268) );
  XNOR U17644 ( .A(n18269), .B(n18257), .Z(n18259) );
  XOR U17645 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n18270), .Z(n18257) );
  AND U17646 ( .A(n2446), .B(n18271), .Z(n18270) );
  IV U17647 ( .A(n18267), .Z(n18269) );
  XOR U17648 ( .A(n18272), .B(n18273), .Z(n18267) );
  AND U17649 ( .A(n2441), .B(n18266), .Z(n18273) );
  XOR U17650 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n18272), 
        .Z(n18266) );
  XOR U17651 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n18274), 
        .Z(n18272) );
  AND U17652 ( .A(n2443), .B(n18271), .Z(n18274) );
  XOR U17653 ( .A(n18275), .B(n18276), .Z(n18271) );
  IV U17654 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n18276)
         );
  IV U17655 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n18275) );
  XOR U17656 ( .A(n49), .B(n18277), .Z(o[14]) );
  AND U17657 ( .A(n62), .B(n18278), .Z(n49) );
  XOR U17658 ( .A(n50), .B(n18277), .Z(n18278) );
  XOR U17659 ( .A(n18279), .B(n18280), .Z(n18277) );
  AND U17660 ( .A(n82), .B(n18281), .Z(n18280) );
  XOR U17661 ( .A(n18282), .B(n15), .Z(n50) );
  AND U17662 ( .A(n65), .B(n18283), .Z(n15) );
  XOR U17663 ( .A(n16), .B(n18282), .Z(n18283) );
  XOR U17664 ( .A(n18284), .B(n18285), .Z(n16) );
  AND U17665 ( .A(n70), .B(n18286), .Z(n18285) );
  XOR U17666 ( .A(p_input[14]), .B(n18284), .Z(n18286) );
  XNOR U17667 ( .A(n18287), .B(n18288), .Z(n18284) );
  AND U17668 ( .A(n74), .B(n18289), .Z(n18288) );
  XOR U17669 ( .A(n18290), .B(n18291), .Z(n18282) );
  AND U17670 ( .A(n78), .B(n18281), .Z(n18291) );
  XNOR U17671 ( .A(n18292), .B(n18279), .Z(n18281) );
  XOR U17672 ( .A(n18293), .B(n18294), .Z(n18279) );
  AND U17673 ( .A(n102), .B(n18295), .Z(n18294) );
  IV U17674 ( .A(n18290), .Z(n18292) );
  XOR U17675 ( .A(n18296), .B(n18297), .Z(n18290) );
  AND U17676 ( .A(n86), .B(n18289), .Z(n18297) );
  XNOR U17677 ( .A(n18287), .B(n18296), .Z(n18289) );
  XNOR U17678 ( .A(n18298), .B(n18299), .Z(n18287) );
  AND U17679 ( .A(n90), .B(n18300), .Z(n18299) );
  XOR U17680 ( .A(p_input[30]), .B(n18298), .Z(n18300) );
  XNOR U17681 ( .A(n18301), .B(n18302), .Z(n18298) );
  AND U17682 ( .A(n94), .B(n18303), .Z(n18302) );
  XOR U17683 ( .A(n18304), .B(n18305), .Z(n18296) );
  AND U17684 ( .A(n98), .B(n18295), .Z(n18305) );
  XNOR U17685 ( .A(n18306), .B(n18293), .Z(n18295) );
  XOR U17686 ( .A(n18307), .B(n18308), .Z(n18293) );
  AND U17687 ( .A(n121), .B(n18309), .Z(n18308) );
  IV U17688 ( .A(n18304), .Z(n18306) );
  XOR U17689 ( .A(n18310), .B(n18311), .Z(n18304) );
  AND U17690 ( .A(n105), .B(n18303), .Z(n18311) );
  XNOR U17691 ( .A(n18301), .B(n18310), .Z(n18303) );
  XNOR U17692 ( .A(n18312), .B(n18313), .Z(n18301) );
  AND U17693 ( .A(n109), .B(n18314), .Z(n18313) );
  XOR U17694 ( .A(p_input[46]), .B(n18312), .Z(n18314) );
  XNOR U17695 ( .A(n18315), .B(n18316), .Z(n18312) );
  AND U17696 ( .A(n113), .B(n18317), .Z(n18316) );
  XOR U17697 ( .A(n18318), .B(n18319), .Z(n18310) );
  AND U17698 ( .A(n117), .B(n18309), .Z(n18319) );
  XNOR U17699 ( .A(n18320), .B(n18307), .Z(n18309) );
  XOR U17700 ( .A(n18321), .B(n18322), .Z(n18307) );
  AND U17701 ( .A(n140), .B(n18323), .Z(n18322) );
  IV U17702 ( .A(n18318), .Z(n18320) );
  XOR U17703 ( .A(n18324), .B(n18325), .Z(n18318) );
  AND U17704 ( .A(n124), .B(n18317), .Z(n18325) );
  XNOR U17705 ( .A(n18315), .B(n18324), .Z(n18317) );
  XNOR U17706 ( .A(n18326), .B(n18327), .Z(n18315) );
  AND U17707 ( .A(n128), .B(n18328), .Z(n18327) );
  XOR U17708 ( .A(p_input[62]), .B(n18326), .Z(n18328) );
  XNOR U17709 ( .A(n18329), .B(n18330), .Z(n18326) );
  AND U17710 ( .A(n132), .B(n18331), .Z(n18330) );
  XOR U17711 ( .A(n18332), .B(n18333), .Z(n18324) );
  AND U17712 ( .A(n136), .B(n18323), .Z(n18333) );
  XNOR U17713 ( .A(n18334), .B(n18321), .Z(n18323) );
  XOR U17714 ( .A(n18335), .B(n18336), .Z(n18321) );
  AND U17715 ( .A(n159), .B(n18337), .Z(n18336) );
  IV U17716 ( .A(n18332), .Z(n18334) );
  XOR U17717 ( .A(n18338), .B(n18339), .Z(n18332) );
  AND U17718 ( .A(n143), .B(n18331), .Z(n18339) );
  XNOR U17719 ( .A(n18329), .B(n18338), .Z(n18331) );
  XNOR U17720 ( .A(n18340), .B(n18341), .Z(n18329) );
  AND U17721 ( .A(n147), .B(n18342), .Z(n18341) );
  XOR U17722 ( .A(p_input[78]), .B(n18340), .Z(n18342) );
  XNOR U17723 ( .A(n18343), .B(n18344), .Z(n18340) );
  AND U17724 ( .A(n151), .B(n18345), .Z(n18344) );
  XOR U17725 ( .A(n18346), .B(n18347), .Z(n18338) );
  AND U17726 ( .A(n155), .B(n18337), .Z(n18347) );
  XNOR U17727 ( .A(n18348), .B(n18335), .Z(n18337) );
  XOR U17728 ( .A(n18349), .B(n18350), .Z(n18335) );
  AND U17729 ( .A(n178), .B(n18351), .Z(n18350) );
  IV U17730 ( .A(n18346), .Z(n18348) );
  XOR U17731 ( .A(n18352), .B(n18353), .Z(n18346) );
  AND U17732 ( .A(n162), .B(n18345), .Z(n18353) );
  XNOR U17733 ( .A(n18343), .B(n18352), .Z(n18345) );
  XNOR U17734 ( .A(n18354), .B(n18355), .Z(n18343) );
  AND U17735 ( .A(n166), .B(n18356), .Z(n18355) );
  XOR U17736 ( .A(p_input[94]), .B(n18354), .Z(n18356) );
  XNOR U17737 ( .A(n18357), .B(n18358), .Z(n18354) );
  AND U17738 ( .A(n170), .B(n18359), .Z(n18358) );
  XOR U17739 ( .A(n18360), .B(n18361), .Z(n18352) );
  AND U17740 ( .A(n174), .B(n18351), .Z(n18361) );
  XNOR U17741 ( .A(n18362), .B(n18349), .Z(n18351) );
  XOR U17742 ( .A(n18363), .B(n18364), .Z(n18349) );
  AND U17743 ( .A(n197), .B(n18365), .Z(n18364) );
  IV U17744 ( .A(n18360), .Z(n18362) );
  XOR U17745 ( .A(n18366), .B(n18367), .Z(n18360) );
  AND U17746 ( .A(n181), .B(n18359), .Z(n18367) );
  XNOR U17747 ( .A(n18357), .B(n18366), .Z(n18359) );
  XNOR U17748 ( .A(n18368), .B(n18369), .Z(n18357) );
  AND U17749 ( .A(n185), .B(n18370), .Z(n18369) );
  XOR U17750 ( .A(p_input[110]), .B(n18368), .Z(n18370) );
  XNOR U17751 ( .A(n18371), .B(n18372), .Z(n18368) );
  AND U17752 ( .A(n189), .B(n18373), .Z(n18372) );
  XOR U17753 ( .A(n18374), .B(n18375), .Z(n18366) );
  AND U17754 ( .A(n193), .B(n18365), .Z(n18375) );
  XNOR U17755 ( .A(n18376), .B(n18363), .Z(n18365) );
  XOR U17756 ( .A(n18377), .B(n18378), .Z(n18363) );
  AND U17757 ( .A(n216), .B(n18379), .Z(n18378) );
  IV U17758 ( .A(n18374), .Z(n18376) );
  XOR U17759 ( .A(n18380), .B(n18381), .Z(n18374) );
  AND U17760 ( .A(n200), .B(n18373), .Z(n18381) );
  XNOR U17761 ( .A(n18371), .B(n18380), .Z(n18373) );
  XNOR U17762 ( .A(n18382), .B(n18383), .Z(n18371) );
  AND U17763 ( .A(n204), .B(n18384), .Z(n18383) );
  XOR U17764 ( .A(p_input[126]), .B(n18382), .Z(n18384) );
  XNOR U17765 ( .A(n18385), .B(n18386), .Z(n18382) );
  AND U17766 ( .A(n208), .B(n18387), .Z(n18386) );
  XOR U17767 ( .A(n18388), .B(n18389), .Z(n18380) );
  AND U17768 ( .A(n212), .B(n18379), .Z(n18389) );
  XNOR U17769 ( .A(n18390), .B(n18377), .Z(n18379) );
  XOR U17770 ( .A(n18391), .B(n18392), .Z(n18377) );
  AND U17771 ( .A(n235), .B(n18393), .Z(n18392) );
  IV U17772 ( .A(n18388), .Z(n18390) );
  XOR U17773 ( .A(n18394), .B(n18395), .Z(n18388) );
  AND U17774 ( .A(n219), .B(n18387), .Z(n18395) );
  XNOR U17775 ( .A(n18385), .B(n18394), .Z(n18387) );
  XNOR U17776 ( .A(n18396), .B(n18397), .Z(n18385) );
  AND U17777 ( .A(n223), .B(n18398), .Z(n18397) );
  XOR U17778 ( .A(p_input[142]), .B(n18396), .Z(n18398) );
  XNOR U17779 ( .A(n18399), .B(n18400), .Z(n18396) );
  AND U17780 ( .A(n227), .B(n18401), .Z(n18400) );
  XOR U17781 ( .A(n18402), .B(n18403), .Z(n18394) );
  AND U17782 ( .A(n231), .B(n18393), .Z(n18403) );
  XNOR U17783 ( .A(n18404), .B(n18391), .Z(n18393) );
  XOR U17784 ( .A(n18405), .B(n18406), .Z(n18391) );
  AND U17785 ( .A(n254), .B(n18407), .Z(n18406) );
  IV U17786 ( .A(n18402), .Z(n18404) );
  XOR U17787 ( .A(n18408), .B(n18409), .Z(n18402) );
  AND U17788 ( .A(n238), .B(n18401), .Z(n18409) );
  XNOR U17789 ( .A(n18399), .B(n18408), .Z(n18401) );
  XNOR U17790 ( .A(n18410), .B(n18411), .Z(n18399) );
  AND U17791 ( .A(n242), .B(n18412), .Z(n18411) );
  XOR U17792 ( .A(p_input[158]), .B(n18410), .Z(n18412) );
  XNOR U17793 ( .A(n18413), .B(n18414), .Z(n18410) );
  AND U17794 ( .A(n246), .B(n18415), .Z(n18414) );
  XOR U17795 ( .A(n18416), .B(n18417), .Z(n18408) );
  AND U17796 ( .A(n250), .B(n18407), .Z(n18417) );
  XNOR U17797 ( .A(n18418), .B(n18405), .Z(n18407) );
  XOR U17798 ( .A(n18419), .B(n18420), .Z(n18405) );
  AND U17799 ( .A(n273), .B(n18421), .Z(n18420) );
  IV U17800 ( .A(n18416), .Z(n18418) );
  XOR U17801 ( .A(n18422), .B(n18423), .Z(n18416) );
  AND U17802 ( .A(n257), .B(n18415), .Z(n18423) );
  XNOR U17803 ( .A(n18413), .B(n18422), .Z(n18415) );
  XNOR U17804 ( .A(n18424), .B(n18425), .Z(n18413) );
  AND U17805 ( .A(n261), .B(n18426), .Z(n18425) );
  XOR U17806 ( .A(p_input[174]), .B(n18424), .Z(n18426) );
  XNOR U17807 ( .A(n18427), .B(n18428), .Z(n18424) );
  AND U17808 ( .A(n265), .B(n18429), .Z(n18428) );
  XOR U17809 ( .A(n18430), .B(n18431), .Z(n18422) );
  AND U17810 ( .A(n269), .B(n18421), .Z(n18431) );
  XNOR U17811 ( .A(n18432), .B(n18419), .Z(n18421) );
  XOR U17812 ( .A(n18433), .B(n18434), .Z(n18419) );
  AND U17813 ( .A(n292), .B(n18435), .Z(n18434) );
  IV U17814 ( .A(n18430), .Z(n18432) );
  XOR U17815 ( .A(n18436), .B(n18437), .Z(n18430) );
  AND U17816 ( .A(n276), .B(n18429), .Z(n18437) );
  XNOR U17817 ( .A(n18427), .B(n18436), .Z(n18429) );
  XNOR U17818 ( .A(n18438), .B(n18439), .Z(n18427) );
  AND U17819 ( .A(n280), .B(n18440), .Z(n18439) );
  XOR U17820 ( .A(p_input[190]), .B(n18438), .Z(n18440) );
  XNOR U17821 ( .A(n18441), .B(n18442), .Z(n18438) );
  AND U17822 ( .A(n284), .B(n18443), .Z(n18442) );
  XOR U17823 ( .A(n18444), .B(n18445), .Z(n18436) );
  AND U17824 ( .A(n288), .B(n18435), .Z(n18445) );
  XNOR U17825 ( .A(n18446), .B(n18433), .Z(n18435) );
  XOR U17826 ( .A(n18447), .B(n18448), .Z(n18433) );
  AND U17827 ( .A(n311), .B(n18449), .Z(n18448) );
  IV U17828 ( .A(n18444), .Z(n18446) );
  XOR U17829 ( .A(n18450), .B(n18451), .Z(n18444) );
  AND U17830 ( .A(n295), .B(n18443), .Z(n18451) );
  XNOR U17831 ( .A(n18441), .B(n18450), .Z(n18443) );
  XNOR U17832 ( .A(n18452), .B(n18453), .Z(n18441) );
  AND U17833 ( .A(n299), .B(n18454), .Z(n18453) );
  XOR U17834 ( .A(p_input[206]), .B(n18452), .Z(n18454) );
  XNOR U17835 ( .A(n18455), .B(n18456), .Z(n18452) );
  AND U17836 ( .A(n303), .B(n18457), .Z(n18456) );
  XOR U17837 ( .A(n18458), .B(n18459), .Z(n18450) );
  AND U17838 ( .A(n307), .B(n18449), .Z(n18459) );
  XNOR U17839 ( .A(n18460), .B(n18447), .Z(n18449) );
  XOR U17840 ( .A(n18461), .B(n18462), .Z(n18447) );
  AND U17841 ( .A(n330), .B(n18463), .Z(n18462) );
  IV U17842 ( .A(n18458), .Z(n18460) );
  XOR U17843 ( .A(n18464), .B(n18465), .Z(n18458) );
  AND U17844 ( .A(n314), .B(n18457), .Z(n18465) );
  XNOR U17845 ( .A(n18455), .B(n18464), .Z(n18457) );
  XNOR U17846 ( .A(n18466), .B(n18467), .Z(n18455) );
  AND U17847 ( .A(n318), .B(n18468), .Z(n18467) );
  XOR U17848 ( .A(p_input[222]), .B(n18466), .Z(n18468) );
  XNOR U17849 ( .A(n18469), .B(n18470), .Z(n18466) );
  AND U17850 ( .A(n322), .B(n18471), .Z(n18470) );
  XOR U17851 ( .A(n18472), .B(n18473), .Z(n18464) );
  AND U17852 ( .A(n326), .B(n18463), .Z(n18473) );
  XNOR U17853 ( .A(n18474), .B(n18461), .Z(n18463) );
  XOR U17854 ( .A(n18475), .B(n18476), .Z(n18461) );
  AND U17855 ( .A(n349), .B(n18477), .Z(n18476) );
  IV U17856 ( .A(n18472), .Z(n18474) );
  XOR U17857 ( .A(n18478), .B(n18479), .Z(n18472) );
  AND U17858 ( .A(n333), .B(n18471), .Z(n18479) );
  XNOR U17859 ( .A(n18469), .B(n18478), .Z(n18471) );
  XNOR U17860 ( .A(n18480), .B(n18481), .Z(n18469) );
  AND U17861 ( .A(n337), .B(n18482), .Z(n18481) );
  XOR U17862 ( .A(p_input[238]), .B(n18480), .Z(n18482) );
  XNOR U17863 ( .A(n18483), .B(n18484), .Z(n18480) );
  AND U17864 ( .A(n341), .B(n18485), .Z(n18484) );
  XOR U17865 ( .A(n18486), .B(n18487), .Z(n18478) );
  AND U17866 ( .A(n345), .B(n18477), .Z(n18487) );
  XNOR U17867 ( .A(n18488), .B(n18475), .Z(n18477) );
  XOR U17868 ( .A(n18489), .B(n18490), .Z(n18475) );
  AND U17869 ( .A(n368), .B(n18491), .Z(n18490) );
  IV U17870 ( .A(n18486), .Z(n18488) );
  XOR U17871 ( .A(n18492), .B(n18493), .Z(n18486) );
  AND U17872 ( .A(n352), .B(n18485), .Z(n18493) );
  XNOR U17873 ( .A(n18483), .B(n18492), .Z(n18485) );
  XNOR U17874 ( .A(n18494), .B(n18495), .Z(n18483) );
  AND U17875 ( .A(n356), .B(n18496), .Z(n18495) );
  XOR U17876 ( .A(p_input[254]), .B(n18494), .Z(n18496) );
  XNOR U17877 ( .A(n18497), .B(n18498), .Z(n18494) );
  AND U17878 ( .A(n360), .B(n18499), .Z(n18498) );
  XOR U17879 ( .A(n18500), .B(n18501), .Z(n18492) );
  AND U17880 ( .A(n364), .B(n18491), .Z(n18501) );
  XNOR U17881 ( .A(n18502), .B(n18489), .Z(n18491) );
  XOR U17882 ( .A(n18503), .B(n18504), .Z(n18489) );
  AND U17883 ( .A(n387), .B(n18505), .Z(n18504) );
  IV U17884 ( .A(n18500), .Z(n18502) );
  XOR U17885 ( .A(n18506), .B(n18507), .Z(n18500) );
  AND U17886 ( .A(n371), .B(n18499), .Z(n18507) );
  XNOR U17887 ( .A(n18497), .B(n18506), .Z(n18499) );
  XNOR U17888 ( .A(n18508), .B(n18509), .Z(n18497) );
  AND U17889 ( .A(n375), .B(n18510), .Z(n18509) );
  XOR U17890 ( .A(p_input[270]), .B(n18508), .Z(n18510) );
  XNOR U17891 ( .A(n18511), .B(n18512), .Z(n18508) );
  AND U17892 ( .A(n379), .B(n18513), .Z(n18512) );
  XOR U17893 ( .A(n18514), .B(n18515), .Z(n18506) );
  AND U17894 ( .A(n383), .B(n18505), .Z(n18515) );
  XNOR U17895 ( .A(n18516), .B(n18503), .Z(n18505) );
  XOR U17896 ( .A(n18517), .B(n18518), .Z(n18503) );
  AND U17897 ( .A(n406), .B(n18519), .Z(n18518) );
  IV U17898 ( .A(n18514), .Z(n18516) );
  XOR U17899 ( .A(n18520), .B(n18521), .Z(n18514) );
  AND U17900 ( .A(n390), .B(n18513), .Z(n18521) );
  XNOR U17901 ( .A(n18511), .B(n18520), .Z(n18513) );
  XNOR U17902 ( .A(n18522), .B(n18523), .Z(n18511) );
  AND U17903 ( .A(n394), .B(n18524), .Z(n18523) );
  XOR U17904 ( .A(p_input[286]), .B(n18522), .Z(n18524) );
  XNOR U17905 ( .A(n18525), .B(n18526), .Z(n18522) );
  AND U17906 ( .A(n398), .B(n18527), .Z(n18526) );
  XOR U17907 ( .A(n18528), .B(n18529), .Z(n18520) );
  AND U17908 ( .A(n402), .B(n18519), .Z(n18529) );
  XNOR U17909 ( .A(n18530), .B(n18517), .Z(n18519) );
  XOR U17910 ( .A(n18531), .B(n18532), .Z(n18517) );
  AND U17911 ( .A(n425), .B(n18533), .Z(n18532) );
  IV U17912 ( .A(n18528), .Z(n18530) );
  XOR U17913 ( .A(n18534), .B(n18535), .Z(n18528) );
  AND U17914 ( .A(n409), .B(n18527), .Z(n18535) );
  XNOR U17915 ( .A(n18525), .B(n18534), .Z(n18527) );
  XNOR U17916 ( .A(n18536), .B(n18537), .Z(n18525) );
  AND U17917 ( .A(n413), .B(n18538), .Z(n18537) );
  XOR U17918 ( .A(p_input[302]), .B(n18536), .Z(n18538) );
  XNOR U17919 ( .A(n18539), .B(n18540), .Z(n18536) );
  AND U17920 ( .A(n417), .B(n18541), .Z(n18540) );
  XOR U17921 ( .A(n18542), .B(n18543), .Z(n18534) );
  AND U17922 ( .A(n421), .B(n18533), .Z(n18543) );
  XNOR U17923 ( .A(n18544), .B(n18531), .Z(n18533) );
  XOR U17924 ( .A(n18545), .B(n18546), .Z(n18531) );
  AND U17925 ( .A(n444), .B(n18547), .Z(n18546) );
  IV U17926 ( .A(n18542), .Z(n18544) );
  XOR U17927 ( .A(n18548), .B(n18549), .Z(n18542) );
  AND U17928 ( .A(n428), .B(n18541), .Z(n18549) );
  XNOR U17929 ( .A(n18539), .B(n18548), .Z(n18541) );
  XNOR U17930 ( .A(n18550), .B(n18551), .Z(n18539) );
  AND U17931 ( .A(n432), .B(n18552), .Z(n18551) );
  XOR U17932 ( .A(p_input[318]), .B(n18550), .Z(n18552) );
  XNOR U17933 ( .A(n18553), .B(n18554), .Z(n18550) );
  AND U17934 ( .A(n436), .B(n18555), .Z(n18554) );
  XOR U17935 ( .A(n18556), .B(n18557), .Z(n18548) );
  AND U17936 ( .A(n440), .B(n18547), .Z(n18557) );
  XNOR U17937 ( .A(n18558), .B(n18545), .Z(n18547) );
  XOR U17938 ( .A(n18559), .B(n18560), .Z(n18545) );
  AND U17939 ( .A(n463), .B(n18561), .Z(n18560) );
  IV U17940 ( .A(n18556), .Z(n18558) );
  XOR U17941 ( .A(n18562), .B(n18563), .Z(n18556) );
  AND U17942 ( .A(n447), .B(n18555), .Z(n18563) );
  XNOR U17943 ( .A(n18553), .B(n18562), .Z(n18555) );
  XNOR U17944 ( .A(n18564), .B(n18565), .Z(n18553) );
  AND U17945 ( .A(n451), .B(n18566), .Z(n18565) );
  XOR U17946 ( .A(p_input[334]), .B(n18564), .Z(n18566) );
  XNOR U17947 ( .A(n18567), .B(n18568), .Z(n18564) );
  AND U17948 ( .A(n455), .B(n18569), .Z(n18568) );
  XOR U17949 ( .A(n18570), .B(n18571), .Z(n18562) );
  AND U17950 ( .A(n459), .B(n18561), .Z(n18571) );
  XNOR U17951 ( .A(n18572), .B(n18559), .Z(n18561) );
  XOR U17952 ( .A(n18573), .B(n18574), .Z(n18559) );
  AND U17953 ( .A(n482), .B(n18575), .Z(n18574) );
  IV U17954 ( .A(n18570), .Z(n18572) );
  XOR U17955 ( .A(n18576), .B(n18577), .Z(n18570) );
  AND U17956 ( .A(n466), .B(n18569), .Z(n18577) );
  XNOR U17957 ( .A(n18567), .B(n18576), .Z(n18569) );
  XNOR U17958 ( .A(n18578), .B(n18579), .Z(n18567) );
  AND U17959 ( .A(n470), .B(n18580), .Z(n18579) );
  XOR U17960 ( .A(p_input[350]), .B(n18578), .Z(n18580) );
  XNOR U17961 ( .A(n18581), .B(n18582), .Z(n18578) );
  AND U17962 ( .A(n474), .B(n18583), .Z(n18582) );
  XOR U17963 ( .A(n18584), .B(n18585), .Z(n18576) );
  AND U17964 ( .A(n478), .B(n18575), .Z(n18585) );
  XNOR U17965 ( .A(n18586), .B(n18573), .Z(n18575) );
  XOR U17966 ( .A(n18587), .B(n18588), .Z(n18573) );
  AND U17967 ( .A(n501), .B(n18589), .Z(n18588) );
  IV U17968 ( .A(n18584), .Z(n18586) );
  XOR U17969 ( .A(n18590), .B(n18591), .Z(n18584) );
  AND U17970 ( .A(n485), .B(n18583), .Z(n18591) );
  XNOR U17971 ( .A(n18581), .B(n18590), .Z(n18583) );
  XNOR U17972 ( .A(n18592), .B(n18593), .Z(n18581) );
  AND U17973 ( .A(n489), .B(n18594), .Z(n18593) );
  XOR U17974 ( .A(p_input[366]), .B(n18592), .Z(n18594) );
  XNOR U17975 ( .A(n18595), .B(n18596), .Z(n18592) );
  AND U17976 ( .A(n493), .B(n18597), .Z(n18596) );
  XOR U17977 ( .A(n18598), .B(n18599), .Z(n18590) );
  AND U17978 ( .A(n497), .B(n18589), .Z(n18599) );
  XNOR U17979 ( .A(n18600), .B(n18587), .Z(n18589) );
  XOR U17980 ( .A(n18601), .B(n18602), .Z(n18587) );
  AND U17981 ( .A(n520), .B(n18603), .Z(n18602) );
  IV U17982 ( .A(n18598), .Z(n18600) );
  XOR U17983 ( .A(n18604), .B(n18605), .Z(n18598) );
  AND U17984 ( .A(n504), .B(n18597), .Z(n18605) );
  XNOR U17985 ( .A(n18595), .B(n18604), .Z(n18597) );
  XNOR U17986 ( .A(n18606), .B(n18607), .Z(n18595) );
  AND U17987 ( .A(n508), .B(n18608), .Z(n18607) );
  XOR U17988 ( .A(p_input[382]), .B(n18606), .Z(n18608) );
  XNOR U17989 ( .A(n18609), .B(n18610), .Z(n18606) );
  AND U17990 ( .A(n512), .B(n18611), .Z(n18610) );
  XOR U17991 ( .A(n18612), .B(n18613), .Z(n18604) );
  AND U17992 ( .A(n516), .B(n18603), .Z(n18613) );
  XNOR U17993 ( .A(n18614), .B(n18601), .Z(n18603) );
  XOR U17994 ( .A(n18615), .B(n18616), .Z(n18601) );
  AND U17995 ( .A(n539), .B(n18617), .Z(n18616) );
  IV U17996 ( .A(n18612), .Z(n18614) );
  XOR U17997 ( .A(n18618), .B(n18619), .Z(n18612) );
  AND U17998 ( .A(n523), .B(n18611), .Z(n18619) );
  XNOR U17999 ( .A(n18609), .B(n18618), .Z(n18611) );
  XNOR U18000 ( .A(n18620), .B(n18621), .Z(n18609) );
  AND U18001 ( .A(n527), .B(n18622), .Z(n18621) );
  XOR U18002 ( .A(p_input[398]), .B(n18620), .Z(n18622) );
  XNOR U18003 ( .A(n18623), .B(n18624), .Z(n18620) );
  AND U18004 ( .A(n531), .B(n18625), .Z(n18624) );
  XOR U18005 ( .A(n18626), .B(n18627), .Z(n18618) );
  AND U18006 ( .A(n535), .B(n18617), .Z(n18627) );
  XNOR U18007 ( .A(n18628), .B(n18615), .Z(n18617) );
  XOR U18008 ( .A(n18629), .B(n18630), .Z(n18615) );
  AND U18009 ( .A(n558), .B(n18631), .Z(n18630) );
  IV U18010 ( .A(n18626), .Z(n18628) );
  XOR U18011 ( .A(n18632), .B(n18633), .Z(n18626) );
  AND U18012 ( .A(n542), .B(n18625), .Z(n18633) );
  XNOR U18013 ( .A(n18623), .B(n18632), .Z(n18625) );
  XNOR U18014 ( .A(n18634), .B(n18635), .Z(n18623) );
  AND U18015 ( .A(n546), .B(n18636), .Z(n18635) );
  XOR U18016 ( .A(p_input[414]), .B(n18634), .Z(n18636) );
  XNOR U18017 ( .A(n18637), .B(n18638), .Z(n18634) );
  AND U18018 ( .A(n550), .B(n18639), .Z(n18638) );
  XOR U18019 ( .A(n18640), .B(n18641), .Z(n18632) );
  AND U18020 ( .A(n554), .B(n18631), .Z(n18641) );
  XNOR U18021 ( .A(n18642), .B(n18629), .Z(n18631) );
  XOR U18022 ( .A(n18643), .B(n18644), .Z(n18629) );
  AND U18023 ( .A(n577), .B(n18645), .Z(n18644) );
  IV U18024 ( .A(n18640), .Z(n18642) );
  XOR U18025 ( .A(n18646), .B(n18647), .Z(n18640) );
  AND U18026 ( .A(n561), .B(n18639), .Z(n18647) );
  XNOR U18027 ( .A(n18637), .B(n18646), .Z(n18639) );
  XNOR U18028 ( .A(n18648), .B(n18649), .Z(n18637) );
  AND U18029 ( .A(n565), .B(n18650), .Z(n18649) );
  XOR U18030 ( .A(p_input[430]), .B(n18648), .Z(n18650) );
  XNOR U18031 ( .A(n18651), .B(n18652), .Z(n18648) );
  AND U18032 ( .A(n569), .B(n18653), .Z(n18652) );
  XOR U18033 ( .A(n18654), .B(n18655), .Z(n18646) );
  AND U18034 ( .A(n573), .B(n18645), .Z(n18655) );
  XNOR U18035 ( .A(n18656), .B(n18643), .Z(n18645) );
  XOR U18036 ( .A(n18657), .B(n18658), .Z(n18643) );
  AND U18037 ( .A(n596), .B(n18659), .Z(n18658) );
  IV U18038 ( .A(n18654), .Z(n18656) );
  XOR U18039 ( .A(n18660), .B(n18661), .Z(n18654) );
  AND U18040 ( .A(n580), .B(n18653), .Z(n18661) );
  XNOR U18041 ( .A(n18651), .B(n18660), .Z(n18653) );
  XNOR U18042 ( .A(n18662), .B(n18663), .Z(n18651) );
  AND U18043 ( .A(n584), .B(n18664), .Z(n18663) );
  XOR U18044 ( .A(p_input[446]), .B(n18662), .Z(n18664) );
  XNOR U18045 ( .A(n18665), .B(n18666), .Z(n18662) );
  AND U18046 ( .A(n588), .B(n18667), .Z(n18666) );
  XOR U18047 ( .A(n18668), .B(n18669), .Z(n18660) );
  AND U18048 ( .A(n592), .B(n18659), .Z(n18669) );
  XNOR U18049 ( .A(n18670), .B(n18657), .Z(n18659) );
  XOR U18050 ( .A(n18671), .B(n18672), .Z(n18657) );
  AND U18051 ( .A(n615), .B(n18673), .Z(n18672) );
  IV U18052 ( .A(n18668), .Z(n18670) );
  XOR U18053 ( .A(n18674), .B(n18675), .Z(n18668) );
  AND U18054 ( .A(n599), .B(n18667), .Z(n18675) );
  XNOR U18055 ( .A(n18665), .B(n18674), .Z(n18667) );
  XNOR U18056 ( .A(n18676), .B(n18677), .Z(n18665) );
  AND U18057 ( .A(n603), .B(n18678), .Z(n18677) );
  XOR U18058 ( .A(p_input[462]), .B(n18676), .Z(n18678) );
  XNOR U18059 ( .A(n18679), .B(n18680), .Z(n18676) );
  AND U18060 ( .A(n607), .B(n18681), .Z(n18680) );
  XOR U18061 ( .A(n18682), .B(n18683), .Z(n18674) );
  AND U18062 ( .A(n611), .B(n18673), .Z(n18683) );
  XNOR U18063 ( .A(n18684), .B(n18671), .Z(n18673) );
  XOR U18064 ( .A(n18685), .B(n18686), .Z(n18671) );
  AND U18065 ( .A(n634), .B(n18687), .Z(n18686) );
  IV U18066 ( .A(n18682), .Z(n18684) );
  XOR U18067 ( .A(n18688), .B(n18689), .Z(n18682) );
  AND U18068 ( .A(n618), .B(n18681), .Z(n18689) );
  XNOR U18069 ( .A(n18679), .B(n18688), .Z(n18681) );
  XNOR U18070 ( .A(n18690), .B(n18691), .Z(n18679) );
  AND U18071 ( .A(n622), .B(n18692), .Z(n18691) );
  XOR U18072 ( .A(p_input[478]), .B(n18690), .Z(n18692) );
  XNOR U18073 ( .A(n18693), .B(n18694), .Z(n18690) );
  AND U18074 ( .A(n626), .B(n18695), .Z(n18694) );
  XOR U18075 ( .A(n18696), .B(n18697), .Z(n18688) );
  AND U18076 ( .A(n630), .B(n18687), .Z(n18697) );
  XNOR U18077 ( .A(n18698), .B(n18685), .Z(n18687) );
  XOR U18078 ( .A(n18699), .B(n18700), .Z(n18685) );
  AND U18079 ( .A(n653), .B(n18701), .Z(n18700) );
  IV U18080 ( .A(n18696), .Z(n18698) );
  XOR U18081 ( .A(n18702), .B(n18703), .Z(n18696) );
  AND U18082 ( .A(n637), .B(n18695), .Z(n18703) );
  XNOR U18083 ( .A(n18693), .B(n18702), .Z(n18695) );
  XNOR U18084 ( .A(n18704), .B(n18705), .Z(n18693) );
  AND U18085 ( .A(n641), .B(n18706), .Z(n18705) );
  XOR U18086 ( .A(p_input[494]), .B(n18704), .Z(n18706) );
  XNOR U18087 ( .A(n18707), .B(n18708), .Z(n18704) );
  AND U18088 ( .A(n645), .B(n18709), .Z(n18708) );
  XOR U18089 ( .A(n18710), .B(n18711), .Z(n18702) );
  AND U18090 ( .A(n649), .B(n18701), .Z(n18711) );
  XNOR U18091 ( .A(n18712), .B(n18699), .Z(n18701) );
  XOR U18092 ( .A(n18713), .B(n18714), .Z(n18699) );
  AND U18093 ( .A(n672), .B(n18715), .Z(n18714) );
  IV U18094 ( .A(n18710), .Z(n18712) );
  XOR U18095 ( .A(n18716), .B(n18717), .Z(n18710) );
  AND U18096 ( .A(n656), .B(n18709), .Z(n18717) );
  XNOR U18097 ( .A(n18707), .B(n18716), .Z(n18709) );
  XNOR U18098 ( .A(n18718), .B(n18719), .Z(n18707) );
  AND U18099 ( .A(n660), .B(n18720), .Z(n18719) );
  XOR U18100 ( .A(p_input[510]), .B(n18718), .Z(n18720) );
  XNOR U18101 ( .A(n18721), .B(n18722), .Z(n18718) );
  AND U18102 ( .A(n664), .B(n18723), .Z(n18722) );
  XOR U18103 ( .A(n18724), .B(n18725), .Z(n18716) );
  AND U18104 ( .A(n668), .B(n18715), .Z(n18725) );
  XNOR U18105 ( .A(n18726), .B(n18713), .Z(n18715) );
  XOR U18106 ( .A(n18727), .B(n18728), .Z(n18713) );
  AND U18107 ( .A(n691), .B(n18729), .Z(n18728) );
  IV U18108 ( .A(n18724), .Z(n18726) );
  XOR U18109 ( .A(n18730), .B(n18731), .Z(n18724) );
  AND U18110 ( .A(n675), .B(n18723), .Z(n18731) );
  XNOR U18111 ( .A(n18721), .B(n18730), .Z(n18723) );
  XNOR U18112 ( .A(n18732), .B(n18733), .Z(n18721) );
  AND U18113 ( .A(n679), .B(n18734), .Z(n18733) );
  XOR U18114 ( .A(p_input[526]), .B(n18732), .Z(n18734) );
  XNOR U18115 ( .A(n18735), .B(n18736), .Z(n18732) );
  AND U18116 ( .A(n683), .B(n18737), .Z(n18736) );
  XOR U18117 ( .A(n18738), .B(n18739), .Z(n18730) );
  AND U18118 ( .A(n687), .B(n18729), .Z(n18739) );
  XNOR U18119 ( .A(n18740), .B(n18727), .Z(n18729) );
  XOR U18120 ( .A(n18741), .B(n18742), .Z(n18727) );
  AND U18121 ( .A(n710), .B(n18743), .Z(n18742) );
  IV U18122 ( .A(n18738), .Z(n18740) );
  XOR U18123 ( .A(n18744), .B(n18745), .Z(n18738) );
  AND U18124 ( .A(n694), .B(n18737), .Z(n18745) );
  XNOR U18125 ( .A(n18735), .B(n18744), .Z(n18737) );
  XNOR U18126 ( .A(n18746), .B(n18747), .Z(n18735) );
  AND U18127 ( .A(n698), .B(n18748), .Z(n18747) );
  XOR U18128 ( .A(p_input[542]), .B(n18746), .Z(n18748) );
  XNOR U18129 ( .A(n18749), .B(n18750), .Z(n18746) );
  AND U18130 ( .A(n702), .B(n18751), .Z(n18750) );
  XOR U18131 ( .A(n18752), .B(n18753), .Z(n18744) );
  AND U18132 ( .A(n706), .B(n18743), .Z(n18753) );
  XNOR U18133 ( .A(n18754), .B(n18741), .Z(n18743) );
  XOR U18134 ( .A(n18755), .B(n18756), .Z(n18741) );
  AND U18135 ( .A(n729), .B(n18757), .Z(n18756) );
  IV U18136 ( .A(n18752), .Z(n18754) );
  XOR U18137 ( .A(n18758), .B(n18759), .Z(n18752) );
  AND U18138 ( .A(n713), .B(n18751), .Z(n18759) );
  XNOR U18139 ( .A(n18749), .B(n18758), .Z(n18751) );
  XNOR U18140 ( .A(n18760), .B(n18761), .Z(n18749) );
  AND U18141 ( .A(n717), .B(n18762), .Z(n18761) );
  XOR U18142 ( .A(p_input[558]), .B(n18760), .Z(n18762) );
  XNOR U18143 ( .A(n18763), .B(n18764), .Z(n18760) );
  AND U18144 ( .A(n721), .B(n18765), .Z(n18764) );
  XOR U18145 ( .A(n18766), .B(n18767), .Z(n18758) );
  AND U18146 ( .A(n725), .B(n18757), .Z(n18767) );
  XNOR U18147 ( .A(n18768), .B(n18755), .Z(n18757) );
  XOR U18148 ( .A(n18769), .B(n18770), .Z(n18755) );
  AND U18149 ( .A(n748), .B(n18771), .Z(n18770) );
  IV U18150 ( .A(n18766), .Z(n18768) );
  XOR U18151 ( .A(n18772), .B(n18773), .Z(n18766) );
  AND U18152 ( .A(n732), .B(n18765), .Z(n18773) );
  XNOR U18153 ( .A(n18763), .B(n18772), .Z(n18765) );
  XNOR U18154 ( .A(n18774), .B(n18775), .Z(n18763) );
  AND U18155 ( .A(n736), .B(n18776), .Z(n18775) );
  XOR U18156 ( .A(p_input[574]), .B(n18774), .Z(n18776) );
  XNOR U18157 ( .A(n18777), .B(n18778), .Z(n18774) );
  AND U18158 ( .A(n740), .B(n18779), .Z(n18778) );
  XOR U18159 ( .A(n18780), .B(n18781), .Z(n18772) );
  AND U18160 ( .A(n744), .B(n18771), .Z(n18781) );
  XNOR U18161 ( .A(n18782), .B(n18769), .Z(n18771) );
  XOR U18162 ( .A(n18783), .B(n18784), .Z(n18769) );
  AND U18163 ( .A(n767), .B(n18785), .Z(n18784) );
  IV U18164 ( .A(n18780), .Z(n18782) );
  XOR U18165 ( .A(n18786), .B(n18787), .Z(n18780) );
  AND U18166 ( .A(n751), .B(n18779), .Z(n18787) );
  XNOR U18167 ( .A(n18777), .B(n18786), .Z(n18779) );
  XNOR U18168 ( .A(n18788), .B(n18789), .Z(n18777) );
  AND U18169 ( .A(n755), .B(n18790), .Z(n18789) );
  XOR U18170 ( .A(p_input[590]), .B(n18788), .Z(n18790) );
  XNOR U18171 ( .A(n18791), .B(n18792), .Z(n18788) );
  AND U18172 ( .A(n759), .B(n18793), .Z(n18792) );
  XOR U18173 ( .A(n18794), .B(n18795), .Z(n18786) );
  AND U18174 ( .A(n763), .B(n18785), .Z(n18795) );
  XNOR U18175 ( .A(n18796), .B(n18783), .Z(n18785) );
  XOR U18176 ( .A(n18797), .B(n18798), .Z(n18783) );
  AND U18177 ( .A(n786), .B(n18799), .Z(n18798) );
  IV U18178 ( .A(n18794), .Z(n18796) );
  XOR U18179 ( .A(n18800), .B(n18801), .Z(n18794) );
  AND U18180 ( .A(n770), .B(n18793), .Z(n18801) );
  XNOR U18181 ( .A(n18791), .B(n18800), .Z(n18793) );
  XNOR U18182 ( .A(n18802), .B(n18803), .Z(n18791) );
  AND U18183 ( .A(n774), .B(n18804), .Z(n18803) );
  XOR U18184 ( .A(p_input[606]), .B(n18802), .Z(n18804) );
  XNOR U18185 ( .A(n18805), .B(n18806), .Z(n18802) );
  AND U18186 ( .A(n778), .B(n18807), .Z(n18806) );
  XOR U18187 ( .A(n18808), .B(n18809), .Z(n18800) );
  AND U18188 ( .A(n782), .B(n18799), .Z(n18809) );
  XNOR U18189 ( .A(n18810), .B(n18797), .Z(n18799) );
  XOR U18190 ( .A(n18811), .B(n18812), .Z(n18797) );
  AND U18191 ( .A(n805), .B(n18813), .Z(n18812) );
  IV U18192 ( .A(n18808), .Z(n18810) );
  XOR U18193 ( .A(n18814), .B(n18815), .Z(n18808) );
  AND U18194 ( .A(n789), .B(n18807), .Z(n18815) );
  XNOR U18195 ( .A(n18805), .B(n18814), .Z(n18807) );
  XNOR U18196 ( .A(n18816), .B(n18817), .Z(n18805) );
  AND U18197 ( .A(n793), .B(n18818), .Z(n18817) );
  XOR U18198 ( .A(p_input[622]), .B(n18816), .Z(n18818) );
  XNOR U18199 ( .A(n18819), .B(n18820), .Z(n18816) );
  AND U18200 ( .A(n797), .B(n18821), .Z(n18820) );
  XOR U18201 ( .A(n18822), .B(n18823), .Z(n18814) );
  AND U18202 ( .A(n801), .B(n18813), .Z(n18823) );
  XNOR U18203 ( .A(n18824), .B(n18811), .Z(n18813) );
  XOR U18204 ( .A(n18825), .B(n18826), .Z(n18811) );
  AND U18205 ( .A(n824), .B(n18827), .Z(n18826) );
  IV U18206 ( .A(n18822), .Z(n18824) );
  XOR U18207 ( .A(n18828), .B(n18829), .Z(n18822) );
  AND U18208 ( .A(n808), .B(n18821), .Z(n18829) );
  XNOR U18209 ( .A(n18819), .B(n18828), .Z(n18821) );
  XNOR U18210 ( .A(n18830), .B(n18831), .Z(n18819) );
  AND U18211 ( .A(n812), .B(n18832), .Z(n18831) );
  XOR U18212 ( .A(p_input[638]), .B(n18830), .Z(n18832) );
  XNOR U18213 ( .A(n18833), .B(n18834), .Z(n18830) );
  AND U18214 ( .A(n816), .B(n18835), .Z(n18834) );
  XOR U18215 ( .A(n18836), .B(n18837), .Z(n18828) );
  AND U18216 ( .A(n820), .B(n18827), .Z(n18837) );
  XNOR U18217 ( .A(n18838), .B(n18825), .Z(n18827) );
  XOR U18218 ( .A(n18839), .B(n18840), .Z(n18825) );
  AND U18219 ( .A(n843), .B(n18841), .Z(n18840) );
  IV U18220 ( .A(n18836), .Z(n18838) );
  XOR U18221 ( .A(n18842), .B(n18843), .Z(n18836) );
  AND U18222 ( .A(n827), .B(n18835), .Z(n18843) );
  XNOR U18223 ( .A(n18833), .B(n18842), .Z(n18835) );
  XNOR U18224 ( .A(n18844), .B(n18845), .Z(n18833) );
  AND U18225 ( .A(n831), .B(n18846), .Z(n18845) );
  XOR U18226 ( .A(p_input[654]), .B(n18844), .Z(n18846) );
  XNOR U18227 ( .A(n18847), .B(n18848), .Z(n18844) );
  AND U18228 ( .A(n835), .B(n18849), .Z(n18848) );
  XOR U18229 ( .A(n18850), .B(n18851), .Z(n18842) );
  AND U18230 ( .A(n839), .B(n18841), .Z(n18851) );
  XNOR U18231 ( .A(n18852), .B(n18839), .Z(n18841) );
  XOR U18232 ( .A(n18853), .B(n18854), .Z(n18839) );
  AND U18233 ( .A(n862), .B(n18855), .Z(n18854) );
  IV U18234 ( .A(n18850), .Z(n18852) );
  XOR U18235 ( .A(n18856), .B(n18857), .Z(n18850) );
  AND U18236 ( .A(n846), .B(n18849), .Z(n18857) );
  XNOR U18237 ( .A(n18847), .B(n18856), .Z(n18849) );
  XNOR U18238 ( .A(n18858), .B(n18859), .Z(n18847) );
  AND U18239 ( .A(n850), .B(n18860), .Z(n18859) );
  XOR U18240 ( .A(p_input[670]), .B(n18858), .Z(n18860) );
  XNOR U18241 ( .A(n18861), .B(n18862), .Z(n18858) );
  AND U18242 ( .A(n854), .B(n18863), .Z(n18862) );
  XOR U18243 ( .A(n18864), .B(n18865), .Z(n18856) );
  AND U18244 ( .A(n858), .B(n18855), .Z(n18865) );
  XNOR U18245 ( .A(n18866), .B(n18853), .Z(n18855) );
  XOR U18246 ( .A(n18867), .B(n18868), .Z(n18853) );
  AND U18247 ( .A(n881), .B(n18869), .Z(n18868) );
  IV U18248 ( .A(n18864), .Z(n18866) );
  XOR U18249 ( .A(n18870), .B(n18871), .Z(n18864) );
  AND U18250 ( .A(n865), .B(n18863), .Z(n18871) );
  XNOR U18251 ( .A(n18861), .B(n18870), .Z(n18863) );
  XNOR U18252 ( .A(n18872), .B(n18873), .Z(n18861) );
  AND U18253 ( .A(n869), .B(n18874), .Z(n18873) );
  XOR U18254 ( .A(p_input[686]), .B(n18872), .Z(n18874) );
  XNOR U18255 ( .A(n18875), .B(n18876), .Z(n18872) );
  AND U18256 ( .A(n873), .B(n18877), .Z(n18876) );
  XOR U18257 ( .A(n18878), .B(n18879), .Z(n18870) );
  AND U18258 ( .A(n877), .B(n18869), .Z(n18879) );
  XNOR U18259 ( .A(n18880), .B(n18867), .Z(n18869) );
  XOR U18260 ( .A(n18881), .B(n18882), .Z(n18867) );
  AND U18261 ( .A(n900), .B(n18883), .Z(n18882) );
  IV U18262 ( .A(n18878), .Z(n18880) );
  XOR U18263 ( .A(n18884), .B(n18885), .Z(n18878) );
  AND U18264 ( .A(n884), .B(n18877), .Z(n18885) );
  XNOR U18265 ( .A(n18875), .B(n18884), .Z(n18877) );
  XNOR U18266 ( .A(n18886), .B(n18887), .Z(n18875) );
  AND U18267 ( .A(n888), .B(n18888), .Z(n18887) );
  XOR U18268 ( .A(p_input[702]), .B(n18886), .Z(n18888) );
  XNOR U18269 ( .A(n18889), .B(n18890), .Z(n18886) );
  AND U18270 ( .A(n892), .B(n18891), .Z(n18890) );
  XOR U18271 ( .A(n18892), .B(n18893), .Z(n18884) );
  AND U18272 ( .A(n896), .B(n18883), .Z(n18893) );
  XNOR U18273 ( .A(n18894), .B(n18881), .Z(n18883) );
  XOR U18274 ( .A(n18895), .B(n18896), .Z(n18881) );
  AND U18275 ( .A(n919), .B(n18897), .Z(n18896) );
  IV U18276 ( .A(n18892), .Z(n18894) );
  XOR U18277 ( .A(n18898), .B(n18899), .Z(n18892) );
  AND U18278 ( .A(n903), .B(n18891), .Z(n18899) );
  XNOR U18279 ( .A(n18889), .B(n18898), .Z(n18891) );
  XNOR U18280 ( .A(n18900), .B(n18901), .Z(n18889) );
  AND U18281 ( .A(n907), .B(n18902), .Z(n18901) );
  XOR U18282 ( .A(p_input[718]), .B(n18900), .Z(n18902) );
  XNOR U18283 ( .A(n18903), .B(n18904), .Z(n18900) );
  AND U18284 ( .A(n911), .B(n18905), .Z(n18904) );
  XOR U18285 ( .A(n18906), .B(n18907), .Z(n18898) );
  AND U18286 ( .A(n915), .B(n18897), .Z(n18907) );
  XNOR U18287 ( .A(n18908), .B(n18895), .Z(n18897) );
  XOR U18288 ( .A(n18909), .B(n18910), .Z(n18895) );
  AND U18289 ( .A(n938), .B(n18911), .Z(n18910) );
  IV U18290 ( .A(n18906), .Z(n18908) );
  XOR U18291 ( .A(n18912), .B(n18913), .Z(n18906) );
  AND U18292 ( .A(n922), .B(n18905), .Z(n18913) );
  XNOR U18293 ( .A(n18903), .B(n18912), .Z(n18905) );
  XNOR U18294 ( .A(n18914), .B(n18915), .Z(n18903) );
  AND U18295 ( .A(n926), .B(n18916), .Z(n18915) );
  XOR U18296 ( .A(p_input[734]), .B(n18914), .Z(n18916) );
  XNOR U18297 ( .A(n18917), .B(n18918), .Z(n18914) );
  AND U18298 ( .A(n930), .B(n18919), .Z(n18918) );
  XOR U18299 ( .A(n18920), .B(n18921), .Z(n18912) );
  AND U18300 ( .A(n934), .B(n18911), .Z(n18921) );
  XNOR U18301 ( .A(n18922), .B(n18909), .Z(n18911) );
  XOR U18302 ( .A(n18923), .B(n18924), .Z(n18909) );
  AND U18303 ( .A(n957), .B(n18925), .Z(n18924) );
  IV U18304 ( .A(n18920), .Z(n18922) );
  XOR U18305 ( .A(n18926), .B(n18927), .Z(n18920) );
  AND U18306 ( .A(n941), .B(n18919), .Z(n18927) );
  XNOR U18307 ( .A(n18917), .B(n18926), .Z(n18919) );
  XNOR U18308 ( .A(n18928), .B(n18929), .Z(n18917) );
  AND U18309 ( .A(n945), .B(n18930), .Z(n18929) );
  XOR U18310 ( .A(p_input[750]), .B(n18928), .Z(n18930) );
  XNOR U18311 ( .A(n18931), .B(n18932), .Z(n18928) );
  AND U18312 ( .A(n949), .B(n18933), .Z(n18932) );
  XOR U18313 ( .A(n18934), .B(n18935), .Z(n18926) );
  AND U18314 ( .A(n953), .B(n18925), .Z(n18935) );
  XNOR U18315 ( .A(n18936), .B(n18923), .Z(n18925) );
  XOR U18316 ( .A(n18937), .B(n18938), .Z(n18923) );
  AND U18317 ( .A(n976), .B(n18939), .Z(n18938) );
  IV U18318 ( .A(n18934), .Z(n18936) );
  XOR U18319 ( .A(n18940), .B(n18941), .Z(n18934) );
  AND U18320 ( .A(n960), .B(n18933), .Z(n18941) );
  XNOR U18321 ( .A(n18931), .B(n18940), .Z(n18933) );
  XNOR U18322 ( .A(n18942), .B(n18943), .Z(n18931) );
  AND U18323 ( .A(n964), .B(n18944), .Z(n18943) );
  XOR U18324 ( .A(p_input[766]), .B(n18942), .Z(n18944) );
  XNOR U18325 ( .A(n18945), .B(n18946), .Z(n18942) );
  AND U18326 ( .A(n968), .B(n18947), .Z(n18946) );
  XOR U18327 ( .A(n18948), .B(n18949), .Z(n18940) );
  AND U18328 ( .A(n972), .B(n18939), .Z(n18949) );
  XNOR U18329 ( .A(n18950), .B(n18937), .Z(n18939) );
  XOR U18330 ( .A(n18951), .B(n18952), .Z(n18937) );
  AND U18331 ( .A(n995), .B(n18953), .Z(n18952) );
  IV U18332 ( .A(n18948), .Z(n18950) );
  XOR U18333 ( .A(n18954), .B(n18955), .Z(n18948) );
  AND U18334 ( .A(n979), .B(n18947), .Z(n18955) );
  XNOR U18335 ( .A(n18945), .B(n18954), .Z(n18947) );
  XNOR U18336 ( .A(n18956), .B(n18957), .Z(n18945) );
  AND U18337 ( .A(n983), .B(n18958), .Z(n18957) );
  XOR U18338 ( .A(p_input[782]), .B(n18956), .Z(n18958) );
  XNOR U18339 ( .A(n18959), .B(n18960), .Z(n18956) );
  AND U18340 ( .A(n987), .B(n18961), .Z(n18960) );
  XOR U18341 ( .A(n18962), .B(n18963), .Z(n18954) );
  AND U18342 ( .A(n991), .B(n18953), .Z(n18963) );
  XNOR U18343 ( .A(n18964), .B(n18951), .Z(n18953) );
  XOR U18344 ( .A(n18965), .B(n18966), .Z(n18951) );
  AND U18345 ( .A(n1014), .B(n18967), .Z(n18966) );
  IV U18346 ( .A(n18962), .Z(n18964) );
  XOR U18347 ( .A(n18968), .B(n18969), .Z(n18962) );
  AND U18348 ( .A(n998), .B(n18961), .Z(n18969) );
  XNOR U18349 ( .A(n18959), .B(n18968), .Z(n18961) );
  XNOR U18350 ( .A(n18970), .B(n18971), .Z(n18959) );
  AND U18351 ( .A(n1002), .B(n18972), .Z(n18971) );
  XOR U18352 ( .A(p_input[798]), .B(n18970), .Z(n18972) );
  XNOR U18353 ( .A(n18973), .B(n18974), .Z(n18970) );
  AND U18354 ( .A(n1006), .B(n18975), .Z(n18974) );
  XOR U18355 ( .A(n18976), .B(n18977), .Z(n18968) );
  AND U18356 ( .A(n1010), .B(n18967), .Z(n18977) );
  XNOR U18357 ( .A(n18978), .B(n18965), .Z(n18967) );
  XOR U18358 ( .A(n18979), .B(n18980), .Z(n18965) );
  AND U18359 ( .A(n1033), .B(n18981), .Z(n18980) );
  IV U18360 ( .A(n18976), .Z(n18978) );
  XOR U18361 ( .A(n18982), .B(n18983), .Z(n18976) );
  AND U18362 ( .A(n1017), .B(n18975), .Z(n18983) );
  XNOR U18363 ( .A(n18973), .B(n18982), .Z(n18975) );
  XNOR U18364 ( .A(n18984), .B(n18985), .Z(n18973) );
  AND U18365 ( .A(n1021), .B(n18986), .Z(n18985) );
  XOR U18366 ( .A(p_input[814]), .B(n18984), .Z(n18986) );
  XNOR U18367 ( .A(n18987), .B(n18988), .Z(n18984) );
  AND U18368 ( .A(n1025), .B(n18989), .Z(n18988) );
  XOR U18369 ( .A(n18990), .B(n18991), .Z(n18982) );
  AND U18370 ( .A(n1029), .B(n18981), .Z(n18991) );
  XNOR U18371 ( .A(n18992), .B(n18979), .Z(n18981) );
  XOR U18372 ( .A(n18993), .B(n18994), .Z(n18979) );
  AND U18373 ( .A(n1052), .B(n18995), .Z(n18994) );
  IV U18374 ( .A(n18990), .Z(n18992) );
  XOR U18375 ( .A(n18996), .B(n18997), .Z(n18990) );
  AND U18376 ( .A(n1036), .B(n18989), .Z(n18997) );
  XNOR U18377 ( .A(n18987), .B(n18996), .Z(n18989) );
  XNOR U18378 ( .A(n18998), .B(n18999), .Z(n18987) );
  AND U18379 ( .A(n1040), .B(n19000), .Z(n18999) );
  XOR U18380 ( .A(p_input[830]), .B(n18998), .Z(n19000) );
  XNOR U18381 ( .A(n19001), .B(n19002), .Z(n18998) );
  AND U18382 ( .A(n1044), .B(n19003), .Z(n19002) );
  XOR U18383 ( .A(n19004), .B(n19005), .Z(n18996) );
  AND U18384 ( .A(n1048), .B(n18995), .Z(n19005) );
  XNOR U18385 ( .A(n19006), .B(n18993), .Z(n18995) );
  XOR U18386 ( .A(n19007), .B(n19008), .Z(n18993) );
  AND U18387 ( .A(n1071), .B(n19009), .Z(n19008) );
  IV U18388 ( .A(n19004), .Z(n19006) );
  XOR U18389 ( .A(n19010), .B(n19011), .Z(n19004) );
  AND U18390 ( .A(n1055), .B(n19003), .Z(n19011) );
  XNOR U18391 ( .A(n19001), .B(n19010), .Z(n19003) );
  XNOR U18392 ( .A(n19012), .B(n19013), .Z(n19001) );
  AND U18393 ( .A(n1059), .B(n19014), .Z(n19013) );
  XOR U18394 ( .A(p_input[846]), .B(n19012), .Z(n19014) );
  XNOR U18395 ( .A(n19015), .B(n19016), .Z(n19012) );
  AND U18396 ( .A(n1063), .B(n19017), .Z(n19016) );
  XOR U18397 ( .A(n19018), .B(n19019), .Z(n19010) );
  AND U18398 ( .A(n1067), .B(n19009), .Z(n19019) );
  XNOR U18399 ( .A(n19020), .B(n19007), .Z(n19009) );
  XOR U18400 ( .A(n19021), .B(n19022), .Z(n19007) );
  AND U18401 ( .A(n1090), .B(n19023), .Z(n19022) );
  IV U18402 ( .A(n19018), .Z(n19020) );
  XOR U18403 ( .A(n19024), .B(n19025), .Z(n19018) );
  AND U18404 ( .A(n1074), .B(n19017), .Z(n19025) );
  XNOR U18405 ( .A(n19015), .B(n19024), .Z(n19017) );
  XNOR U18406 ( .A(n19026), .B(n19027), .Z(n19015) );
  AND U18407 ( .A(n1078), .B(n19028), .Z(n19027) );
  XOR U18408 ( .A(p_input[862]), .B(n19026), .Z(n19028) );
  XNOR U18409 ( .A(n19029), .B(n19030), .Z(n19026) );
  AND U18410 ( .A(n1082), .B(n19031), .Z(n19030) );
  XOR U18411 ( .A(n19032), .B(n19033), .Z(n19024) );
  AND U18412 ( .A(n1086), .B(n19023), .Z(n19033) );
  XNOR U18413 ( .A(n19034), .B(n19021), .Z(n19023) );
  XOR U18414 ( .A(n19035), .B(n19036), .Z(n19021) );
  AND U18415 ( .A(n1109), .B(n19037), .Z(n19036) );
  IV U18416 ( .A(n19032), .Z(n19034) );
  XOR U18417 ( .A(n19038), .B(n19039), .Z(n19032) );
  AND U18418 ( .A(n1093), .B(n19031), .Z(n19039) );
  XNOR U18419 ( .A(n19029), .B(n19038), .Z(n19031) );
  XNOR U18420 ( .A(n19040), .B(n19041), .Z(n19029) );
  AND U18421 ( .A(n1097), .B(n19042), .Z(n19041) );
  XOR U18422 ( .A(p_input[878]), .B(n19040), .Z(n19042) );
  XNOR U18423 ( .A(n19043), .B(n19044), .Z(n19040) );
  AND U18424 ( .A(n1101), .B(n19045), .Z(n19044) );
  XOR U18425 ( .A(n19046), .B(n19047), .Z(n19038) );
  AND U18426 ( .A(n1105), .B(n19037), .Z(n19047) );
  XNOR U18427 ( .A(n19048), .B(n19035), .Z(n19037) );
  XOR U18428 ( .A(n19049), .B(n19050), .Z(n19035) );
  AND U18429 ( .A(n1128), .B(n19051), .Z(n19050) );
  IV U18430 ( .A(n19046), .Z(n19048) );
  XOR U18431 ( .A(n19052), .B(n19053), .Z(n19046) );
  AND U18432 ( .A(n1112), .B(n19045), .Z(n19053) );
  XNOR U18433 ( .A(n19043), .B(n19052), .Z(n19045) );
  XNOR U18434 ( .A(n19054), .B(n19055), .Z(n19043) );
  AND U18435 ( .A(n1116), .B(n19056), .Z(n19055) );
  XOR U18436 ( .A(p_input[894]), .B(n19054), .Z(n19056) );
  XNOR U18437 ( .A(n19057), .B(n19058), .Z(n19054) );
  AND U18438 ( .A(n1120), .B(n19059), .Z(n19058) );
  XOR U18439 ( .A(n19060), .B(n19061), .Z(n19052) );
  AND U18440 ( .A(n1124), .B(n19051), .Z(n19061) );
  XNOR U18441 ( .A(n19062), .B(n19049), .Z(n19051) );
  XOR U18442 ( .A(n19063), .B(n19064), .Z(n19049) );
  AND U18443 ( .A(n1147), .B(n19065), .Z(n19064) );
  IV U18444 ( .A(n19060), .Z(n19062) );
  XOR U18445 ( .A(n19066), .B(n19067), .Z(n19060) );
  AND U18446 ( .A(n1131), .B(n19059), .Z(n19067) );
  XNOR U18447 ( .A(n19057), .B(n19066), .Z(n19059) );
  XNOR U18448 ( .A(n19068), .B(n19069), .Z(n19057) );
  AND U18449 ( .A(n1135), .B(n19070), .Z(n19069) );
  XOR U18450 ( .A(p_input[910]), .B(n19068), .Z(n19070) );
  XNOR U18451 ( .A(n19071), .B(n19072), .Z(n19068) );
  AND U18452 ( .A(n1139), .B(n19073), .Z(n19072) );
  XOR U18453 ( .A(n19074), .B(n19075), .Z(n19066) );
  AND U18454 ( .A(n1143), .B(n19065), .Z(n19075) );
  XNOR U18455 ( .A(n19076), .B(n19063), .Z(n19065) );
  XOR U18456 ( .A(n19077), .B(n19078), .Z(n19063) );
  AND U18457 ( .A(n1166), .B(n19079), .Z(n19078) );
  IV U18458 ( .A(n19074), .Z(n19076) );
  XOR U18459 ( .A(n19080), .B(n19081), .Z(n19074) );
  AND U18460 ( .A(n1150), .B(n19073), .Z(n19081) );
  XNOR U18461 ( .A(n19071), .B(n19080), .Z(n19073) );
  XNOR U18462 ( .A(n19082), .B(n19083), .Z(n19071) );
  AND U18463 ( .A(n1154), .B(n19084), .Z(n19083) );
  XOR U18464 ( .A(p_input[926]), .B(n19082), .Z(n19084) );
  XNOR U18465 ( .A(n19085), .B(n19086), .Z(n19082) );
  AND U18466 ( .A(n1158), .B(n19087), .Z(n19086) );
  XOR U18467 ( .A(n19088), .B(n19089), .Z(n19080) );
  AND U18468 ( .A(n1162), .B(n19079), .Z(n19089) );
  XNOR U18469 ( .A(n19090), .B(n19077), .Z(n19079) );
  XOR U18470 ( .A(n19091), .B(n19092), .Z(n19077) );
  AND U18471 ( .A(n1185), .B(n19093), .Z(n19092) );
  IV U18472 ( .A(n19088), .Z(n19090) );
  XOR U18473 ( .A(n19094), .B(n19095), .Z(n19088) );
  AND U18474 ( .A(n1169), .B(n19087), .Z(n19095) );
  XNOR U18475 ( .A(n19085), .B(n19094), .Z(n19087) );
  XNOR U18476 ( .A(n19096), .B(n19097), .Z(n19085) );
  AND U18477 ( .A(n1173), .B(n19098), .Z(n19097) );
  XOR U18478 ( .A(p_input[942]), .B(n19096), .Z(n19098) );
  XNOR U18479 ( .A(n19099), .B(n19100), .Z(n19096) );
  AND U18480 ( .A(n1177), .B(n19101), .Z(n19100) );
  XOR U18481 ( .A(n19102), .B(n19103), .Z(n19094) );
  AND U18482 ( .A(n1181), .B(n19093), .Z(n19103) );
  XNOR U18483 ( .A(n19104), .B(n19091), .Z(n19093) );
  XOR U18484 ( .A(n19105), .B(n19106), .Z(n19091) );
  AND U18485 ( .A(n1204), .B(n19107), .Z(n19106) );
  IV U18486 ( .A(n19102), .Z(n19104) );
  XOR U18487 ( .A(n19108), .B(n19109), .Z(n19102) );
  AND U18488 ( .A(n1188), .B(n19101), .Z(n19109) );
  XNOR U18489 ( .A(n19099), .B(n19108), .Z(n19101) );
  XNOR U18490 ( .A(n19110), .B(n19111), .Z(n19099) );
  AND U18491 ( .A(n1192), .B(n19112), .Z(n19111) );
  XOR U18492 ( .A(p_input[958]), .B(n19110), .Z(n19112) );
  XNOR U18493 ( .A(n19113), .B(n19114), .Z(n19110) );
  AND U18494 ( .A(n1196), .B(n19115), .Z(n19114) );
  XOR U18495 ( .A(n19116), .B(n19117), .Z(n19108) );
  AND U18496 ( .A(n1200), .B(n19107), .Z(n19117) );
  XNOR U18497 ( .A(n19118), .B(n19105), .Z(n19107) );
  XOR U18498 ( .A(n19119), .B(n19120), .Z(n19105) );
  AND U18499 ( .A(n1223), .B(n19121), .Z(n19120) );
  IV U18500 ( .A(n19116), .Z(n19118) );
  XOR U18501 ( .A(n19122), .B(n19123), .Z(n19116) );
  AND U18502 ( .A(n1207), .B(n19115), .Z(n19123) );
  XNOR U18503 ( .A(n19113), .B(n19122), .Z(n19115) );
  XNOR U18504 ( .A(n19124), .B(n19125), .Z(n19113) );
  AND U18505 ( .A(n1211), .B(n19126), .Z(n19125) );
  XOR U18506 ( .A(p_input[974]), .B(n19124), .Z(n19126) );
  XNOR U18507 ( .A(n19127), .B(n19128), .Z(n19124) );
  AND U18508 ( .A(n1215), .B(n19129), .Z(n19128) );
  XOR U18509 ( .A(n19130), .B(n19131), .Z(n19122) );
  AND U18510 ( .A(n1219), .B(n19121), .Z(n19131) );
  XNOR U18511 ( .A(n19132), .B(n19119), .Z(n19121) );
  XOR U18512 ( .A(n19133), .B(n19134), .Z(n19119) );
  AND U18513 ( .A(n1242), .B(n19135), .Z(n19134) );
  IV U18514 ( .A(n19130), .Z(n19132) );
  XOR U18515 ( .A(n19136), .B(n19137), .Z(n19130) );
  AND U18516 ( .A(n1226), .B(n19129), .Z(n19137) );
  XNOR U18517 ( .A(n19127), .B(n19136), .Z(n19129) );
  XNOR U18518 ( .A(n19138), .B(n19139), .Z(n19127) );
  AND U18519 ( .A(n1230), .B(n19140), .Z(n19139) );
  XOR U18520 ( .A(p_input[990]), .B(n19138), .Z(n19140) );
  XNOR U18521 ( .A(n19141), .B(n19142), .Z(n19138) );
  AND U18522 ( .A(n1234), .B(n19143), .Z(n19142) );
  XOR U18523 ( .A(n19144), .B(n19145), .Z(n19136) );
  AND U18524 ( .A(n1238), .B(n19135), .Z(n19145) );
  XNOR U18525 ( .A(n19146), .B(n19133), .Z(n19135) );
  XOR U18526 ( .A(n19147), .B(n19148), .Z(n19133) );
  AND U18527 ( .A(n1261), .B(n19149), .Z(n19148) );
  IV U18528 ( .A(n19144), .Z(n19146) );
  XOR U18529 ( .A(n19150), .B(n19151), .Z(n19144) );
  AND U18530 ( .A(n1245), .B(n19143), .Z(n19151) );
  XNOR U18531 ( .A(n19141), .B(n19150), .Z(n19143) );
  XNOR U18532 ( .A(n19152), .B(n19153), .Z(n19141) );
  AND U18533 ( .A(n1249), .B(n19154), .Z(n19153) );
  XOR U18534 ( .A(p_input[1006]), .B(n19152), .Z(n19154) );
  XNOR U18535 ( .A(n19155), .B(n19156), .Z(n19152) );
  AND U18536 ( .A(n1253), .B(n19157), .Z(n19156) );
  XOR U18537 ( .A(n19158), .B(n19159), .Z(n19150) );
  AND U18538 ( .A(n1257), .B(n19149), .Z(n19159) );
  XNOR U18539 ( .A(n19160), .B(n19147), .Z(n19149) );
  XOR U18540 ( .A(n19161), .B(n19162), .Z(n19147) );
  AND U18541 ( .A(n1280), .B(n19163), .Z(n19162) );
  IV U18542 ( .A(n19158), .Z(n19160) );
  XOR U18543 ( .A(n19164), .B(n19165), .Z(n19158) );
  AND U18544 ( .A(n1264), .B(n19157), .Z(n19165) );
  XNOR U18545 ( .A(n19155), .B(n19164), .Z(n19157) );
  XNOR U18546 ( .A(n19166), .B(n19167), .Z(n19155) );
  AND U18547 ( .A(n1268), .B(n19168), .Z(n19167) );
  XOR U18548 ( .A(p_input[1022]), .B(n19166), .Z(n19168) );
  XNOR U18549 ( .A(n19169), .B(n19170), .Z(n19166) );
  AND U18550 ( .A(n1272), .B(n19171), .Z(n19170) );
  XOR U18551 ( .A(n19172), .B(n19173), .Z(n19164) );
  AND U18552 ( .A(n1276), .B(n19163), .Z(n19173) );
  XNOR U18553 ( .A(n19174), .B(n19161), .Z(n19163) );
  XOR U18554 ( .A(n19175), .B(n19176), .Z(n19161) );
  AND U18555 ( .A(n1299), .B(n19177), .Z(n19176) );
  IV U18556 ( .A(n19172), .Z(n19174) );
  XOR U18557 ( .A(n19178), .B(n19179), .Z(n19172) );
  AND U18558 ( .A(n1283), .B(n19171), .Z(n19179) );
  XNOR U18559 ( .A(n19169), .B(n19178), .Z(n19171) );
  XNOR U18560 ( .A(n19180), .B(n19181), .Z(n19169) );
  AND U18561 ( .A(n1287), .B(n19182), .Z(n19181) );
  XOR U18562 ( .A(p_input[1038]), .B(n19180), .Z(n19182) );
  XNOR U18563 ( .A(n19183), .B(n19184), .Z(n19180) );
  AND U18564 ( .A(n1291), .B(n19185), .Z(n19184) );
  XOR U18565 ( .A(n19186), .B(n19187), .Z(n19178) );
  AND U18566 ( .A(n1295), .B(n19177), .Z(n19187) );
  XNOR U18567 ( .A(n19188), .B(n19175), .Z(n19177) );
  XOR U18568 ( .A(n19189), .B(n19190), .Z(n19175) );
  AND U18569 ( .A(n1318), .B(n19191), .Z(n19190) );
  IV U18570 ( .A(n19186), .Z(n19188) );
  XOR U18571 ( .A(n19192), .B(n19193), .Z(n19186) );
  AND U18572 ( .A(n1302), .B(n19185), .Z(n19193) );
  XNOR U18573 ( .A(n19183), .B(n19192), .Z(n19185) );
  XNOR U18574 ( .A(n19194), .B(n19195), .Z(n19183) );
  AND U18575 ( .A(n1306), .B(n19196), .Z(n19195) );
  XOR U18576 ( .A(p_input[1054]), .B(n19194), .Z(n19196) );
  XNOR U18577 ( .A(n19197), .B(n19198), .Z(n19194) );
  AND U18578 ( .A(n1310), .B(n19199), .Z(n19198) );
  XOR U18579 ( .A(n19200), .B(n19201), .Z(n19192) );
  AND U18580 ( .A(n1314), .B(n19191), .Z(n19201) );
  XNOR U18581 ( .A(n19202), .B(n19189), .Z(n19191) );
  XOR U18582 ( .A(n19203), .B(n19204), .Z(n19189) );
  AND U18583 ( .A(n1337), .B(n19205), .Z(n19204) );
  IV U18584 ( .A(n19200), .Z(n19202) );
  XOR U18585 ( .A(n19206), .B(n19207), .Z(n19200) );
  AND U18586 ( .A(n1321), .B(n19199), .Z(n19207) );
  XNOR U18587 ( .A(n19197), .B(n19206), .Z(n19199) );
  XNOR U18588 ( .A(n19208), .B(n19209), .Z(n19197) );
  AND U18589 ( .A(n1325), .B(n19210), .Z(n19209) );
  XOR U18590 ( .A(p_input[1070]), .B(n19208), .Z(n19210) );
  XNOR U18591 ( .A(n19211), .B(n19212), .Z(n19208) );
  AND U18592 ( .A(n1329), .B(n19213), .Z(n19212) );
  XOR U18593 ( .A(n19214), .B(n19215), .Z(n19206) );
  AND U18594 ( .A(n1333), .B(n19205), .Z(n19215) );
  XNOR U18595 ( .A(n19216), .B(n19203), .Z(n19205) );
  XOR U18596 ( .A(n19217), .B(n19218), .Z(n19203) );
  AND U18597 ( .A(n1356), .B(n19219), .Z(n19218) );
  IV U18598 ( .A(n19214), .Z(n19216) );
  XOR U18599 ( .A(n19220), .B(n19221), .Z(n19214) );
  AND U18600 ( .A(n1340), .B(n19213), .Z(n19221) );
  XNOR U18601 ( .A(n19211), .B(n19220), .Z(n19213) );
  XNOR U18602 ( .A(n19222), .B(n19223), .Z(n19211) );
  AND U18603 ( .A(n1344), .B(n19224), .Z(n19223) );
  XOR U18604 ( .A(p_input[1086]), .B(n19222), .Z(n19224) );
  XNOR U18605 ( .A(n19225), .B(n19226), .Z(n19222) );
  AND U18606 ( .A(n1348), .B(n19227), .Z(n19226) );
  XOR U18607 ( .A(n19228), .B(n19229), .Z(n19220) );
  AND U18608 ( .A(n1352), .B(n19219), .Z(n19229) );
  XNOR U18609 ( .A(n19230), .B(n19217), .Z(n19219) );
  XOR U18610 ( .A(n19231), .B(n19232), .Z(n19217) );
  AND U18611 ( .A(n1375), .B(n19233), .Z(n19232) );
  IV U18612 ( .A(n19228), .Z(n19230) );
  XOR U18613 ( .A(n19234), .B(n19235), .Z(n19228) );
  AND U18614 ( .A(n1359), .B(n19227), .Z(n19235) );
  XNOR U18615 ( .A(n19225), .B(n19234), .Z(n19227) );
  XNOR U18616 ( .A(n19236), .B(n19237), .Z(n19225) );
  AND U18617 ( .A(n1363), .B(n19238), .Z(n19237) );
  XOR U18618 ( .A(p_input[1102]), .B(n19236), .Z(n19238) );
  XNOR U18619 ( .A(n19239), .B(n19240), .Z(n19236) );
  AND U18620 ( .A(n1367), .B(n19241), .Z(n19240) );
  XOR U18621 ( .A(n19242), .B(n19243), .Z(n19234) );
  AND U18622 ( .A(n1371), .B(n19233), .Z(n19243) );
  XNOR U18623 ( .A(n19244), .B(n19231), .Z(n19233) );
  XOR U18624 ( .A(n19245), .B(n19246), .Z(n19231) );
  AND U18625 ( .A(n1394), .B(n19247), .Z(n19246) );
  IV U18626 ( .A(n19242), .Z(n19244) );
  XOR U18627 ( .A(n19248), .B(n19249), .Z(n19242) );
  AND U18628 ( .A(n1378), .B(n19241), .Z(n19249) );
  XNOR U18629 ( .A(n19239), .B(n19248), .Z(n19241) );
  XNOR U18630 ( .A(n19250), .B(n19251), .Z(n19239) );
  AND U18631 ( .A(n1382), .B(n19252), .Z(n19251) );
  XOR U18632 ( .A(p_input[1118]), .B(n19250), .Z(n19252) );
  XNOR U18633 ( .A(n19253), .B(n19254), .Z(n19250) );
  AND U18634 ( .A(n1386), .B(n19255), .Z(n19254) );
  XOR U18635 ( .A(n19256), .B(n19257), .Z(n19248) );
  AND U18636 ( .A(n1390), .B(n19247), .Z(n19257) );
  XNOR U18637 ( .A(n19258), .B(n19245), .Z(n19247) );
  XOR U18638 ( .A(n19259), .B(n19260), .Z(n19245) );
  AND U18639 ( .A(n1413), .B(n19261), .Z(n19260) );
  IV U18640 ( .A(n19256), .Z(n19258) );
  XOR U18641 ( .A(n19262), .B(n19263), .Z(n19256) );
  AND U18642 ( .A(n1397), .B(n19255), .Z(n19263) );
  XNOR U18643 ( .A(n19253), .B(n19262), .Z(n19255) );
  XNOR U18644 ( .A(n19264), .B(n19265), .Z(n19253) );
  AND U18645 ( .A(n1401), .B(n19266), .Z(n19265) );
  XOR U18646 ( .A(p_input[1134]), .B(n19264), .Z(n19266) );
  XNOR U18647 ( .A(n19267), .B(n19268), .Z(n19264) );
  AND U18648 ( .A(n1405), .B(n19269), .Z(n19268) );
  XOR U18649 ( .A(n19270), .B(n19271), .Z(n19262) );
  AND U18650 ( .A(n1409), .B(n19261), .Z(n19271) );
  XNOR U18651 ( .A(n19272), .B(n19259), .Z(n19261) );
  XOR U18652 ( .A(n19273), .B(n19274), .Z(n19259) );
  AND U18653 ( .A(n1432), .B(n19275), .Z(n19274) );
  IV U18654 ( .A(n19270), .Z(n19272) );
  XOR U18655 ( .A(n19276), .B(n19277), .Z(n19270) );
  AND U18656 ( .A(n1416), .B(n19269), .Z(n19277) );
  XNOR U18657 ( .A(n19267), .B(n19276), .Z(n19269) );
  XNOR U18658 ( .A(n19278), .B(n19279), .Z(n19267) );
  AND U18659 ( .A(n1420), .B(n19280), .Z(n19279) );
  XOR U18660 ( .A(p_input[1150]), .B(n19278), .Z(n19280) );
  XNOR U18661 ( .A(n19281), .B(n19282), .Z(n19278) );
  AND U18662 ( .A(n1424), .B(n19283), .Z(n19282) );
  XOR U18663 ( .A(n19284), .B(n19285), .Z(n19276) );
  AND U18664 ( .A(n1428), .B(n19275), .Z(n19285) );
  XNOR U18665 ( .A(n19286), .B(n19273), .Z(n19275) );
  XOR U18666 ( .A(n19287), .B(n19288), .Z(n19273) );
  AND U18667 ( .A(n1451), .B(n19289), .Z(n19288) );
  IV U18668 ( .A(n19284), .Z(n19286) );
  XOR U18669 ( .A(n19290), .B(n19291), .Z(n19284) );
  AND U18670 ( .A(n1435), .B(n19283), .Z(n19291) );
  XNOR U18671 ( .A(n19281), .B(n19290), .Z(n19283) );
  XNOR U18672 ( .A(n19292), .B(n19293), .Z(n19281) );
  AND U18673 ( .A(n1439), .B(n19294), .Z(n19293) );
  XOR U18674 ( .A(p_input[1166]), .B(n19292), .Z(n19294) );
  XNOR U18675 ( .A(n19295), .B(n19296), .Z(n19292) );
  AND U18676 ( .A(n1443), .B(n19297), .Z(n19296) );
  XOR U18677 ( .A(n19298), .B(n19299), .Z(n19290) );
  AND U18678 ( .A(n1447), .B(n19289), .Z(n19299) );
  XNOR U18679 ( .A(n19300), .B(n19287), .Z(n19289) );
  XOR U18680 ( .A(n19301), .B(n19302), .Z(n19287) );
  AND U18681 ( .A(n1470), .B(n19303), .Z(n19302) );
  IV U18682 ( .A(n19298), .Z(n19300) );
  XOR U18683 ( .A(n19304), .B(n19305), .Z(n19298) );
  AND U18684 ( .A(n1454), .B(n19297), .Z(n19305) );
  XNOR U18685 ( .A(n19295), .B(n19304), .Z(n19297) );
  XNOR U18686 ( .A(n19306), .B(n19307), .Z(n19295) );
  AND U18687 ( .A(n1458), .B(n19308), .Z(n19307) );
  XOR U18688 ( .A(p_input[1182]), .B(n19306), .Z(n19308) );
  XNOR U18689 ( .A(n19309), .B(n19310), .Z(n19306) );
  AND U18690 ( .A(n1462), .B(n19311), .Z(n19310) );
  XOR U18691 ( .A(n19312), .B(n19313), .Z(n19304) );
  AND U18692 ( .A(n1466), .B(n19303), .Z(n19313) );
  XNOR U18693 ( .A(n19314), .B(n19301), .Z(n19303) );
  XOR U18694 ( .A(n19315), .B(n19316), .Z(n19301) );
  AND U18695 ( .A(n1489), .B(n19317), .Z(n19316) );
  IV U18696 ( .A(n19312), .Z(n19314) );
  XOR U18697 ( .A(n19318), .B(n19319), .Z(n19312) );
  AND U18698 ( .A(n1473), .B(n19311), .Z(n19319) );
  XNOR U18699 ( .A(n19309), .B(n19318), .Z(n19311) );
  XNOR U18700 ( .A(n19320), .B(n19321), .Z(n19309) );
  AND U18701 ( .A(n1477), .B(n19322), .Z(n19321) );
  XOR U18702 ( .A(p_input[1198]), .B(n19320), .Z(n19322) );
  XNOR U18703 ( .A(n19323), .B(n19324), .Z(n19320) );
  AND U18704 ( .A(n1481), .B(n19325), .Z(n19324) );
  XOR U18705 ( .A(n19326), .B(n19327), .Z(n19318) );
  AND U18706 ( .A(n1485), .B(n19317), .Z(n19327) );
  XNOR U18707 ( .A(n19328), .B(n19315), .Z(n19317) );
  XOR U18708 ( .A(n19329), .B(n19330), .Z(n19315) );
  AND U18709 ( .A(n1508), .B(n19331), .Z(n19330) );
  IV U18710 ( .A(n19326), .Z(n19328) );
  XOR U18711 ( .A(n19332), .B(n19333), .Z(n19326) );
  AND U18712 ( .A(n1492), .B(n19325), .Z(n19333) );
  XNOR U18713 ( .A(n19323), .B(n19332), .Z(n19325) );
  XNOR U18714 ( .A(n19334), .B(n19335), .Z(n19323) );
  AND U18715 ( .A(n1496), .B(n19336), .Z(n19335) );
  XOR U18716 ( .A(p_input[1214]), .B(n19334), .Z(n19336) );
  XNOR U18717 ( .A(n19337), .B(n19338), .Z(n19334) );
  AND U18718 ( .A(n1500), .B(n19339), .Z(n19338) );
  XOR U18719 ( .A(n19340), .B(n19341), .Z(n19332) );
  AND U18720 ( .A(n1504), .B(n19331), .Z(n19341) );
  XNOR U18721 ( .A(n19342), .B(n19329), .Z(n19331) );
  XOR U18722 ( .A(n19343), .B(n19344), .Z(n19329) );
  AND U18723 ( .A(n1527), .B(n19345), .Z(n19344) );
  IV U18724 ( .A(n19340), .Z(n19342) );
  XOR U18725 ( .A(n19346), .B(n19347), .Z(n19340) );
  AND U18726 ( .A(n1511), .B(n19339), .Z(n19347) );
  XNOR U18727 ( .A(n19337), .B(n19346), .Z(n19339) );
  XNOR U18728 ( .A(n19348), .B(n19349), .Z(n19337) );
  AND U18729 ( .A(n1515), .B(n19350), .Z(n19349) );
  XOR U18730 ( .A(p_input[1230]), .B(n19348), .Z(n19350) );
  XNOR U18731 ( .A(n19351), .B(n19352), .Z(n19348) );
  AND U18732 ( .A(n1519), .B(n19353), .Z(n19352) );
  XOR U18733 ( .A(n19354), .B(n19355), .Z(n19346) );
  AND U18734 ( .A(n1523), .B(n19345), .Z(n19355) );
  XNOR U18735 ( .A(n19356), .B(n19343), .Z(n19345) );
  XOR U18736 ( .A(n19357), .B(n19358), .Z(n19343) );
  AND U18737 ( .A(n1546), .B(n19359), .Z(n19358) );
  IV U18738 ( .A(n19354), .Z(n19356) );
  XOR U18739 ( .A(n19360), .B(n19361), .Z(n19354) );
  AND U18740 ( .A(n1530), .B(n19353), .Z(n19361) );
  XNOR U18741 ( .A(n19351), .B(n19360), .Z(n19353) );
  XNOR U18742 ( .A(n19362), .B(n19363), .Z(n19351) );
  AND U18743 ( .A(n1534), .B(n19364), .Z(n19363) );
  XOR U18744 ( .A(p_input[1246]), .B(n19362), .Z(n19364) );
  XNOR U18745 ( .A(n19365), .B(n19366), .Z(n19362) );
  AND U18746 ( .A(n1538), .B(n19367), .Z(n19366) );
  XOR U18747 ( .A(n19368), .B(n19369), .Z(n19360) );
  AND U18748 ( .A(n1542), .B(n19359), .Z(n19369) );
  XNOR U18749 ( .A(n19370), .B(n19357), .Z(n19359) );
  XOR U18750 ( .A(n19371), .B(n19372), .Z(n19357) );
  AND U18751 ( .A(n1565), .B(n19373), .Z(n19372) );
  IV U18752 ( .A(n19368), .Z(n19370) );
  XOR U18753 ( .A(n19374), .B(n19375), .Z(n19368) );
  AND U18754 ( .A(n1549), .B(n19367), .Z(n19375) );
  XNOR U18755 ( .A(n19365), .B(n19374), .Z(n19367) );
  XNOR U18756 ( .A(n19376), .B(n19377), .Z(n19365) );
  AND U18757 ( .A(n1553), .B(n19378), .Z(n19377) );
  XOR U18758 ( .A(p_input[1262]), .B(n19376), .Z(n19378) );
  XNOR U18759 ( .A(n19379), .B(n19380), .Z(n19376) );
  AND U18760 ( .A(n1557), .B(n19381), .Z(n19380) );
  XOR U18761 ( .A(n19382), .B(n19383), .Z(n19374) );
  AND U18762 ( .A(n1561), .B(n19373), .Z(n19383) );
  XNOR U18763 ( .A(n19384), .B(n19371), .Z(n19373) );
  XOR U18764 ( .A(n19385), .B(n19386), .Z(n19371) );
  AND U18765 ( .A(n1584), .B(n19387), .Z(n19386) );
  IV U18766 ( .A(n19382), .Z(n19384) );
  XOR U18767 ( .A(n19388), .B(n19389), .Z(n19382) );
  AND U18768 ( .A(n1568), .B(n19381), .Z(n19389) );
  XNOR U18769 ( .A(n19379), .B(n19388), .Z(n19381) );
  XNOR U18770 ( .A(n19390), .B(n19391), .Z(n19379) );
  AND U18771 ( .A(n1572), .B(n19392), .Z(n19391) );
  XOR U18772 ( .A(p_input[1278]), .B(n19390), .Z(n19392) );
  XNOR U18773 ( .A(n19393), .B(n19394), .Z(n19390) );
  AND U18774 ( .A(n1576), .B(n19395), .Z(n19394) );
  XOR U18775 ( .A(n19396), .B(n19397), .Z(n19388) );
  AND U18776 ( .A(n1580), .B(n19387), .Z(n19397) );
  XNOR U18777 ( .A(n19398), .B(n19385), .Z(n19387) );
  XOR U18778 ( .A(n19399), .B(n19400), .Z(n19385) );
  AND U18779 ( .A(n1603), .B(n19401), .Z(n19400) );
  IV U18780 ( .A(n19396), .Z(n19398) );
  XOR U18781 ( .A(n19402), .B(n19403), .Z(n19396) );
  AND U18782 ( .A(n1587), .B(n19395), .Z(n19403) );
  XNOR U18783 ( .A(n19393), .B(n19402), .Z(n19395) );
  XNOR U18784 ( .A(n19404), .B(n19405), .Z(n19393) );
  AND U18785 ( .A(n1591), .B(n19406), .Z(n19405) );
  XOR U18786 ( .A(p_input[1294]), .B(n19404), .Z(n19406) );
  XNOR U18787 ( .A(n19407), .B(n19408), .Z(n19404) );
  AND U18788 ( .A(n1595), .B(n19409), .Z(n19408) );
  XOR U18789 ( .A(n19410), .B(n19411), .Z(n19402) );
  AND U18790 ( .A(n1599), .B(n19401), .Z(n19411) );
  XNOR U18791 ( .A(n19412), .B(n19399), .Z(n19401) );
  XOR U18792 ( .A(n19413), .B(n19414), .Z(n19399) );
  AND U18793 ( .A(n1622), .B(n19415), .Z(n19414) );
  IV U18794 ( .A(n19410), .Z(n19412) );
  XOR U18795 ( .A(n19416), .B(n19417), .Z(n19410) );
  AND U18796 ( .A(n1606), .B(n19409), .Z(n19417) );
  XNOR U18797 ( .A(n19407), .B(n19416), .Z(n19409) );
  XNOR U18798 ( .A(n19418), .B(n19419), .Z(n19407) );
  AND U18799 ( .A(n1610), .B(n19420), .Z(n19419) );
  XOR U18800 ( .A(p_input[1310]), .B(n19418), .Z(n19420) );
  XNOR U18801 ( .A(n19421), .B(n19422), .Z(n19418) );
  AND U18802 ( .A(n1614), .B(n19423), .Z(n19422) );
  XOR U18803 ( .A(n19424), .B(n19425), .Z(n19416) );
  AND U18804 ( .A(n1618), .B(n19415), .Z(n19425) );
  XNOR U18805 ( .A(n19426), .B(n19413), .Z(n19415) );
  XOR U18806 ( .A(n19427), .B(n19428), .Z(n19413) );
  AND U18807 ( .A(n1641), .B(n19429), .Z(n19428) );
  IV U18808 ( .A(n19424), .Z(n19426) );
  XOR U18809 ( .A(n19430), .B(n19431), .Z(n19424) );
  AND U18810 ( .A(n1625), .B(n19423), .Z(n19431) );
  XNOR U18811 ( .A(n19421), .B(n19430), .Z(n19423) );
  XNOR U18812 ( .A(n19432), .B(n19433), .Z(n19421) );
  AND U18813 ( .A(n1629), .B(n19434), .Z(n19433) );
  XOR U18814 ( .A(p_input[1326]), .B(n19432), .Z(n19434) );
  XNOR U18815 ( .A(n19435), .B(n19436), .Z(n19432) );
  AND U18816 ( .A(n1633), .B(n19437), .Z(n19436) );
  XOR U18817 ( .A(n19438), .B(n19439), .Z(n19430) );
  AND U18818 ( .A(n1637), .B(n19429), .Z(n19439) );
  XNOR U18819 ( .A(n19440), .B(n19427), .Z(n19429) );
  XOR U18820 ( .A(n19441), .B(n19442), .Z(n19427) );
  AND U18821 ( .A(n1660), .B(n19443), .Z(n19442) );
  IV U18822 ( .A(n19438), .Z(n19440) );
  XOR U18823 ( .A(n19444), .B(n19445), .Z(n19438) );
  AND U18824 ( .A(n1644), .B(n19437), .Z(n19445) );
  XNOR U18825 ( .A(n19435), .B(n19444), .Z(n19437) );
  XNOR U18826 ( .A(n19446), .B(n19447), .Z(n19435) );
  AND U18827 ( .A(n1648), .B(n19448), .Z(n19447) );
  XOR U18828 ( .A(p_input[1342]), .B(n19446), .Z(n19448) );
  XNOR U18829 ( .A(n19449), .B(n19450), .Z(n19446) );
  AND U18830 ( .A(n1652), .B(n19451), .Z(n19450) );
  XOR U18831 ( .A(n19452), .B(n19453), .Z(n19444) );
  AND U18832 ( .A(n1656), .B(n19443), .Z(n19453) );
  XNOR U18833 ( .A(n19454), .B(n19441), .Z(n19443) );
  XOR U18834 ( .A(n19455), .B(n19456), .Z(n19441) );
  AND U18835 ( .A(n1679), .B(n19457), .Z(n19456) );
  IV U18836 ( .A(n19452), .Z(n19454) );
  XOR U18837 ( .A(n19458), .B(n19459), .Z(n19452) );
  AND U18838 ( .A(n1663), .B(n19451), .Z(n19459) );
  XNOR U18839 ( .A(n19449), .B(n19458), .Z(n19451) );
  XNOR U18840 ( .A(n19460), .B(n19461), .Z(n19449) );
  AND U18841 ( .A(n1667), .B(n19462), .Z(n19461) );
  XOR U18842 ( .A(p_input[1358]), .B(n19460), .Z(n19462) );
  XNOR U18843 ( .A(n19463), .B(n19464), .Z(n19460) );
  AND U18844 ( .A(n1671), .B(n19465), .Z(n19464) );
  XOR U18845 ( .A(n19466), .B(n19467), .Z(n19458) );
  AND U18846 ( .A(n1675), .B(n19457), .Z(n19467) );
  XNOR U18847 ( .A(n19468), .B(n19455), .Z(n19457) );
  XOR U18848 ( .A(n19469), .B(n19470), .Z(n19455) );
  AND U18849 ( .A(n1698), .B(n19471), .Z(n19470) );
  IV U18850 ( .A(n19466), .Z(n19468) );
  XOR U18851 ( .A(n19472), .B(n19473), .Z(n19466) );
  AND U18852 ( .A(n1682), .B(n19465), .Z(n19473) );
  XNOR U18853 ( .A(n19463), .B(n19472), .Z(n19465) );
  XNOR U18854 ( .A(n19474), .B(n19475), .Z(n19463) );
  AND U18855 ( .A(n1686), .B(n19476), .Z(n19475) );
  XOR U18856 ( .A(p_input[1374]), .B(n19474), .Z(n19476) );
  XNOR U18857 ( .A(n19477), .B(n19478), .Z(n19474) );
  AND U18858 ( .A(n1690), .B(n19479), .Z(n19478) );
  XOR U18859 ( .A(n19480), .B(n19481), .Z(n19472) );
  AND U18860 ( .A(n1694), .B(n19471), .Z(n19481) );
  XNOR U18861 ( .A(n19482), .B(n19469), .Z(n19471) );
  XOR U18862 ( .A(n19483), .B(n19484), .Z(n19469) );
  AND U18863 ( .A(n1717), .B(n19485), .Z(n19484) );
  IV U18864 ( .A(n19480), .Z(n19482) );
  XOR U18865 ( .A(n19486), .B(n19487), .Z(n19480) );
  AND U18866 ( .A(n1701), .B(n19479), .Z(n19487) );
  XNOR U18867 ( .A(n19477), .B(n19486), .Z(n19479) );
  XNOR U18868 ( .A(n19488), .B(n19489), .Z(n19477) );
  AND U18869 ( .A(n1705), .B(n19490), .Z(n19489) );
  XOR U18870 ( .A(p_input[1390]), .B(n19488), .Z(n19490) );
  XNOR U18871 ( .A(n19491), .B(n19492), .Z(n19488) );
  AND U18872 ( .A(n1709), .B(n19493), .Z(n19492) );
  XOR U18873 ( .A(n19494), .B(n19495), .Z(n19486) );
  AND U18874 ( .A(n1713), .B(n19485), .Z(n19495) );
  XNOR U18875 ( .A(n19496), .B(n19483), .Z(n19485) );
  XOR U18876 ( .A(n19497), .B(n19498), .Z(n19483) );
  AND U18877 ( .A(n1736), .B(n19499), .Z(n19498) );
  IV U18878 ( .A(n19494), .Z(n19496) );
  XOR U18879 ( .A(n19500), .B(n19501), .Z(n19494) );
  AND U18880 ( .A(n1720), .B(n19493), .Z(n19501) );
  XNOR U18881 ( .A(n19491), .B(n19500), .Z(n19493) );
  XNOR U18882 ( .A(n19502), .B(n19503), .Z(n19491) );
  AND U18883 ( .A(n1724), .B(n19504), .Z(n19503) );
  XOR U18884 ( .A(p_input[1406]), .B(n19502), .Z(n19504) );
  XNOR U18885 ( .A(n19505), .B(n19506), .Z(n19502) );
  AND U18886 ( .A(n1728), .B(n19507), .Z(n19506) );
  XOR U18887 ( .A(n19508), .B(n19509), .Z(n19500) );
  AND U18888 ( .A(n1732), .B(n19499), .Z(n19509) );
  XNOR U18889 ( .A(n19510), .B(n19497), .Z(n19499) );
  XOR U18890 ( .A(n19511), .B(n19512), .Z(n19497) );
  AND U18891 ( .A(n1755), .B(n19513), .Z(n19512) );
  IV U18892 ( .A(n19508), .Z(n19510) );
  XOR U18893 ( .A(n19514), .B(n19515), .Z(n19508) );
  AND U18894 ( .A(n1739), .B(n19507), .Z(n19515) );
  XNOR U18895 ( .A(n19505), .B(n19514), .Z(n19507) );
  XNOR U18896 ( .A(n19516), .B(n19517), .Z(n19505) );
  AND U18897 ( .A(n1743), .B(n19518), .Z(n19517) );
  XOR U18898 ( .A(p_input[1422]), .B(n19516), .Z(n19518) );
  XNOR U18899 ( .A(n19519), .B(n19520), .Z(n19516) );
  AND U18900 ( .A(n1747), .B(n19521), .Z(n19520) );
  XOR U18901 ( .A(n19522), .B(n19523), .Z(n19514) );
  AND U18902 ( .A(n1751), .B(n19513), .Z(n19523) );
  XNOR U18903 ( .A(n19524), .B(n19511), .Z(n19513) );
  XOR U18904 ( .A(n19525), .B(n19526), .Z(n19511) );
  AND U18905 ( .A(n1774), .B(n19527), .Z(n19526) );
  IV U18906 ( .A(n19522), .Z(n19524) );
  XOR U18907 ( .A(n19528), .B(n19529), .Z(n19522) );
  AND U18908 ( .A(n1758), .B(n19521), .Z(n19529) );
  XNOR U18909 ( .A(n19519), .B(n19528), .Z(n19521) );
  XNOR U18910 ( .A(n19530), .B(n19531), .Z(n19519) );
  AND U18911 ( .A(n1762), .B(n19532), .Z(n19531) );
  XOR U18912 ( .A(p_input[1438]), .B(n19530), .Z(n19532) );
  XNOR U18913 ( .A(n19533), .B(n19534), .Z(n19530) );
  AND U18914 ( .A(n1766), .B(n19535), .Z(n19534) );
  XOR U18915 ( .A(n19536), .B(n19537), .Z(n19528) );
  AND U18916 ( .A(n1770), .B(n19527), .Z(n19537) );
  XNOR U18917 ( .A(n19538), .B(n19525), .Z(n19527) );
  XOR U18918 ( .A(n19539), .B(n19540), .Z(n19525) );
  AND U18919 ( .A(n1793), .B(n19541), .Z(n19540) );
  IV U18920 ( .A(n19536), .Z(n19538) );
  XOR U18921 ( .A(n19542), .B(n19543), .Z(n19536) );
  AND U18922 ( .A(n1777), .B(n19535), .Z(n19543) );
  XNOR U18923 ( .A(n19533), .B(n19542), .Z(n19535) );
  XNOR U18924 ( .A(n19544), .B(n19545), .Z(n19533) );
  AND U18925 ( .A(n1781), .B(n19546), .Z(n19545) );
  XOR U18926 ( .A(p_input[1454]), .B(n19544), .Z(n19546) );
  XNOR U18927 ( .A(n19547), .B(n19548), .Z(n19544) );
  AND U18928 ( .A(n1785), .B(n19549), .Z(n19548) );
  XOR U18929 ( .A(n19550), .B(n19551), .Z(n19542) );
  AND U18930 ( .A(n1789), .B(n19541), .Z(n19551) );
  XNOR U18931 ( .A(n19552), .B(n19539), .Z(n19541) );
  XOR U18932 ( .A(n19553), .B(n19554), .Z(n19539) );
  AND U18933 ( .A(n1812), .B(n19555), .Z(n19554) );
  IV U18934 ( .A(n19550), .Z(n19552) );
  XOR U18935 ( .A(n19556), .B(n19557), .Z(n19550) );
  AND U18936 ( .A(n1796), .B(n19549), .Z(n19557) );
  XNOR U18937 ( .A(n19547), .B(n19556), .Z(n19549) );
  XNOR U18938 ( .A(n19558), .B(n19559), .Z(n19547) );
  AND U18939 ( .A(n1800), .B(n19560), .Z(n19559) );
  XOR U18940 ( .A(p_input[1470]), .B(n19558), .Z(n19560) );
  XNOR U18941 ( .A(n19561), .B(n19562), .Z(n19558) );
  AND U18942 ( .A(n1804), .B(n19563), .Z(n19562) );
  XOR U18943 ( .A(n19564), .B(n19565), .Z(n19556) );
  AND U18944 ( .A(n1808), .B(n19555), .Z(n19565) );
  XNOR U18945 ( .A(n19566), .B(n19553), .Z(n19555) );
  XOR U18946 ( .A(n19567), .B(n19568), .Z(n19553) );
  AND U18947 ( .A(n1831), .B(n19569), .Z(n19568) );
  IV U18948 ( .A(n19564), .Z(n19566) );
  XOR U18949 ( .A(n19570), .B(n19571), .Z(n19564) );
  AND U18950 ( .A(n1815), .B(n19563), .Z(n19571) );
  XNOR U18951 ( .A(n19561), .B(n19570), .Z(n19563) );
  XNOR U18952 ( .A(n19572), .B(n19573), .Z(n19561) );
  AND U18953 ( .A(n1819), .B(n19574), .Z(n19573) );
  XOR U18954 ( .A(p_input[1486]), .B(n19572), .Z(n19574) );
  XNOR U18955 ( .A(n19575), .B(n19576), .Z(n19572) );
  AND U18956 ( .A(n1823), .B(n19577), .Z(n19576) );
  XOR U18957 ( .A(n19578), .B(n19579), .Z(n19570) );
  AND U18958 ( .A(n1827), .B(n19569), .Z(n19579) );
  XNOR U18959 ( .A(n19580), .B(n19567), .Z(n19569) );
  XOR U18960 ( .A(n19581), .B(n19582), .Z(n19567) );
  AND U18961 ( .A(n1850), .B(n19583), .Z(n19582) );
  IV U18962 ( .A(n19578), .Z(n19580) );
  XOR U18963 ( .A(n19584), .B(n19585), .Z(n19578) );
  AND U18964 ( .A(n1834), .B(n19577), .Z(n19585) );
  XNOR U18965 ( .A(n19575), .B(n19584), .Z(n19577) );
  XNOR U18966 ( .A(n19586), .B(n19587), .Z(n19575) );
  AND U18967 ( .A(n1838), .B(n19588), .Z(n19587) );
  XOR U18968 ( .A(p_input[1502]), .B(n19586), .Z(n19588) );
  XNOR U18969 ( .A(n19589), .B(n19590), .Z(n19586) );
  AND U18970 ( .A(n1842), .B(n19591), .Z(n19590) );
  XOR U18971 ( .A(n19592), .B(n19593), .Z(n19584) );
  AND U18972 ( .A(n1846), .B(n19583), .Z(n19593) );
  XNOR U18973 ( .A(n19594), .B(n19581), .Z(n19583) );
  XOR U18974 ( .A(n19595), .B(n19596), .Z(n19581) );
  AND U18975 ( .A(n1869), .B(n19597), .Z(n19596) );
  IV U18976 ( .A(n19592), .Z(n19594) );
  XOR U18977 ( .A(n19598), .B(n19599), .Z(n19592) );
  AND U18978 ( .A(n1853), .B(n19591), .Z(n19599) );
  XNOR U18979 ( .A(n19589), .B(n19598), .Z(n19591) );
  XNOR U18980 ( .A(n19600), .B(n19601), .Z(n19589) );
  AND U18981 ( .A(n1857), .B(n19602), .Z(n19601) );
  XOR U18982 ( .A(p_input[1518]), .B(n19600), .Z(n19602) );
  XNOR U18983 ( .A(n19603), .B(n19604), .Z(n19600) );
  AND U18984 ( .A(n1861), .B(n19605), .Z(n19604) );
  XOR U18985 ( .A(n19606), .B(n19607), .Z(n19598) );
  AND U18986 ( .A(n1865), .B(n19597), .Z(n19607) );
  XNOR U18987 ( .A(n19608), .B(n19595), .Z(n19597) );
  XOR U18988 ( .A(n19609), .B(n19610), .Z(n19595) );
  AND U18989 ( .A(n1888), .B(n19611), .Z(n19610) );
  IV U18990 ( .A(n19606), .Z(n19608) );
  XOR U18991 ( .A(n19612), .B(n19613), .Z(n19606) );
  AND U18992 ( .A(n1872), .B(n19605), .Z(n19613) );
  XNOR U18993 ( .A(n19603), .B(n19612), .Z(n19605) );
  XNOR U18994 ( .A(n19614), .B(n19615), .Z(n19603) );
  AND U18995 ( .A(n1876), .B(n19616), .Z(n19615) );
  XOR U18996 ( .A(p_input[1534]), .B(n19614), .Z(n19616) );
  XNOR U18997 ( .A(n19617), .B(n19618), .Z(n19614) );
  AND U18998 ( .A(n1880), .B(n19619), .Z(n19618) );
  XOR U18999 ( .A(n19620), .B(n19621), .Z(n19612) );
  AND U19000 ( .A(n1884), .B(n19611), .Z(n19621) );
  XNOR U19001 ( .A(n19622), .B(n19609), .Z(n19611) );
  XOR U19002 ( .A(n19623), .B(n19624), .Z(n19609) );
  AND U19003 ( .A(n1907), .B(n19625), .Z(n19624) );
  IV U19004 ( .A(n19620), .Z(n19622) );
  XOR U19005 ( .A(n19626), .B(n19627), .Z(n19620) );
  AND U19006 ( .A(n1891), .B(n19619), .Z(n19627) );
  XNOR U19007 ( .A(n19617), .B(n19626), .Z(n19619) );
  XNOR U19008 ( .A(n19628), .B(n19629), .Z(n19617) );
  AND U19009 ( .A(n1895), .B(n19630), .Z(n19629) );
  XOR U19010 ( .A(p_input[1550]), .B(n19628), .Z(n19630) );
  XNOR U19011 ( .A(n19631), .B(n19632), .Z(n19628) );
  AND U19012 ( .A(n1899), .B(n19633), .Z(n19632) );
  XOR U19013 ( .A(n19634), .B(n19635), .Z(n19626) );
  AND U19014 ( .A(n1903), .B(n19625), .Z(n19635) );
  XNOR U19015 ( .A(n19636), .B(n19623), .Z(n19625) );
  XOR U19016 ( .A(n19637), .B(n19638), .Z(n19623) );
  AND U19017 ( .A(n1926), .B(n19639), .Z(n19638) );
  IV U19018 ( .A(n19634), .Z(n19636) );
  XOR U19019 ( .A(n19640), .B(n19641), .Z(n19634) );
  AND U19020 ( .A(n1910), .B(n19633), .Z(n19641) );
  XNOR U19021 ( .A(n19631), .B(n19640), .Z(n19633) );
  XNOR U19022 ( .A(n19642), .B(n19643), .Z(n19631) );
  AND U19023 ( .A(n1914), .B(n19644), .Z(n19643) );
  XOR U19024 ( .A(p_input[1566]), .B(n19642), .Z(n19644) );
  XNOR U19025 ( .A(n19645), .B(n19646), .Z(n19642) );
  AND U19026 ( .A(n1918), .B(n19647), .Z(n19646) );
  XOR U19027 ( .A(n19648), .B(n19649), .Z(n19640) );
  AND U19028 ( .A(n1922), .B(n19639), .Z(n19649) );
  XNOR U19029 ( .A(n19650), .B(n19637), .Z(n19639) );
  XOR U19030 ( .A(n19651), .B(n19652), .Z(n19637) );
  AND U19031 ( .A(n1945), .B(n19653), .Z(n19652) );
  IV U19032 ( .A(n19648), .Z(n19650) );
  XOR U19033 ( .A(n19654), .B(n19655), .Z(n19648) );
  AND U19034 ( .A(n1929), .B(n19647), .Z(n19655) );
  XNOR U19035 ( .A(n19645), .B(n19654), .Z(n19647) );
  XNOR U19036 ( .A(n19656), .B(n19657), .Z(n19645) );
  AND U19037 ( .A(n1933), .B(n19658), .Z(n19657) );
  XOR U19038 ( .A(p_input[1582]), .B(n19656), .Z(n19658) );
  XNOR U19039 ( .A(n19659), .B(n19660), .Z(n19656) );
  AND U19040 ( .A(n1937), .B(n19661), .Z(n19660) );
  XOR U19041 ( .A(n19662), .B(n19663), .Z(n19654) );
  AND U19042 ( .A(n1941), .B(n19653), .Z(n19663) );
  XNOR U19043 ( .A(n19664), .B(n19651), .Z(n19653) );
  XOR U19044 ( .A(n19665), .B(n19666), .Z(n19651) );
  AND U19045 ( .A(n1964), .B(n19667), .Z(n19666) );
  IV U19046 ( .A(n19662), .Z(n19664) );
  XOR U19047 ( .A(n19668), .B(n19669), .Z(n19662) );
  AND U19048 ( .A(n1948), .B(n19661), .Z(n19669) );
  XNOR U19049 ( .A(n19659), .B(n19668), .Z(n19661) );
  XNOR U19050 ( .A(n19670), .B(n19671), .Z(n19659) );
  AND U19051 ( .A(n1952), .B(n19672), .Z(n19671) );
  XOR U19052 ( .A(p_input[1598]), .B(n19670), .Z(n19672) );
  XNOR U19053 ( .A(n19673), .B(n19674), .Z(n19670) );
  AND U19054 ( .A(n1956), .B(n19675), .Z(n19674) );
  XOR U19055 ( .A(n19676), .B(n19677), .Z(n19668) );
  AND U19056 ( .A(n1960), .B(n19667), .Z(n19677) );
  XNOR U19057 ( .A(n19678), .B(n19665), .Z(n19667) );
  XOR U19058 ( .A(n19679), .B(n19680), .Z(n19665) );
  AND U19059 ( .A(n1983), .B(n19681), .Z(n19680) );
  IV U19060 ( .A(n19676), .Z(n19678) );
  XOR U19061 ( .A(n19682), .B(n19683), .Z(n19676) );
  AND U19062 ( .A(n1967), .B(n19675), .Z(n19683) );
  XNOR U19063 ( .A(n19673), .B(n19682), .Z(n19675) );
  XNOR U19064 ( .A(n19684), .B(n19685), .Z(n19673) );
  AND U19065 ( .A(n1971), .B(n19686), .Z(n19685) );
  XOR U19066 ( .A(p_input[1614]), .B(n19684), .Z(n19686) );
  XNOR U19067 ( .A(n19687), .B(n19688), .Z(n19684) );
  AND U19068 ( .A(n1975), .B(n19689), .Z(n19688) );
  XOR U19069 ( .A(n19690), .B(n19691), .Z(n19682) );
  AND U19070 ( .A(n1979), .B(n19681), .Z(n19691) );
  XNOR U19071 ( .A(n19692), .B(n19679), .Z(n19681) );
  XOR U19072 ( .A(n19693), .B(n19694), .Z(n19679) );
  AND U19073 ( .A(n2002), .B(n19695), .Z(n19694) );
  IV U19074 ( .A(n19690), .Z(n19692) );
  XOR U19075 ( .A(n19696), .B(n19697), .Z(n19690) );
  AND U19076 ( .A(n1986), .B(n19689), .Z(n19697) );
  XNOR U19077 ( .A(n19687), .B(n19696), .Z(n19689) );
  XNOR U19078 ( .A(n19698), .B(n19699), .Z(n19687) );
  AND U19079 ( .A(n1990), .B(n19700), .Z(n19699) );
  XOR U19080 ( .A(p_input[1630]), .B(n19698), .Z(n19700) );
  XNOR U19081 ( .A(n19701), .B(n19702), .Z(n19698) );
  AND U19082 ( .A(n1994), .B(n19703), .Z(n19702) );
  XOR U19083 ( .A(n19704), .B(n19705), .Z(n19696) );
  AND U19084 ( .A(n1998), .B(n19695), .Z(n19705) );
  XNOR U19085 ( .A(n19706), .B(n19693), .Z(n19695) );
  XOR U19086 ( .A(n19707), .B(n19708), .Z(n19693) );
  AND U19087 ( .A(n2021), .B(n19709), .Z(n19708) );
  IV U19088 ( .A(n19704), .Z(n19706) );
  XOR U19089 ( .A(n19710), .B(n19711), .Z(n19704) );
  AND U19090 ( .A(n2005), .B(n19703), .Z(n19711) );
  XNOR U19091 ( .A(n19701), .B(n19710), .Z(n19703) );
  XNOR U19092 ( .A(n19712), .B(n19713), .Z(n19701) );
  AND U19093 ( .A(n2009), .B(n19714), .Z(n19713) );
  XOR U19094 ( .A(p_input[1646]), .B(n19712), .Z(n19714) );
  XNOR U19095 ( .A(n19715), .B(n19716), .Z(n19712) );
  AND U19096 ( .A(n2013), .B(n19717), .Z(n19716) );
  XOR U19097 ( .A(n19718), .B(n19719), .Z(n19710) );
  AND U19098 ( .A(n2017), .B(n19709), .Z(n19719) );
  XNOR U19099 ( .A(n19720), .B(n19707), .Z(n19709) );
  XOR U19100 ( .A(n19721), .B(n19722), .Z(n19707) );
  AND U19101 ( .A(n2040), .B(n19723), .Z(n19722) );
  IV U19102 ( .A(n19718), .Z(n19720) );
  XOR U19103 ( .A(n19724), .B(n19725), .Z(n19718) );
  AND U19104 ( .A(n2024), .B(n19717), .Z(n19725) );
  XNOR U19105 ( .A(n19715), .B(n19724), .Z(n19717) );
  XNOR U19106 ( .A(n19726), .B(n19727), .Z(n19715) );
  AND U19107 ( .A(n2028), .B(n19728), .Z(n19727) );
  XOR U19108 ( .A(p_input[1662]), .B(n19726), .Z(n19728) );
  XNOR U19109 ( .A(n19729), .B(n19730), .Z(n19726) );
  AND U19110 ( .A(n2032), .B(n19731), .Z(n19730) );
  XOR U19111 ( .A(n19732), .B(n19733), .Z(n19724) );
  AND U19112 ( .A(n2036), .B(n19723), .Z(n19733) );
  XNOR U19113 ( .A(n19734), .B(n19721), .Z(n19723) );
  XOR U19114 ( .A(n19735), .B(n19736), .Z(n19721) );
  AND U19115 ( .A(n2059), .B(n19737), .Z(n19736) );
  IV U19116 ( .A(n19732), .Z(n19734) );
  XOR U19117 ( .A(n19738), .B(n19739), .Z(n19732) );
  AND U19118 ( .A(n2043), .B(n19731), .Z(n19739) );
  XNOR U19119 ( .A(n19729), .B(n19738), .Z(n19731) );
  XNOR U19120 ( .A(n19740), .B(n19741), .Z(n19729) );
  AND U19121 ( .A(n2047), .B(n19742), .Z(n19741) );
  XOR U19122 ( .A(p_input[1678]), .B(n19740), .Z(n19742) );
  XNOR U19123 ( .A(n19743), .B(n19744), .Z(n19740) );
  AND U19124 ( .A(n2051), .B(n19745), .Z(n19744) );
  XOR U19125 ( .A(n19746), .B(n19747), .Z(n19738) );
  AND U19126 ( .A(n2055), .B(n19737), .Z(n19747) );
  XNOR U19127 ( .A(n19748), .B(n19735), .Z(n19737) );
  XOR U19128 ( .A(n19749), .B(n19750), .Z(n19735) );
  AND U19129 ( .A(n2078), .B(n19751), .Z(n19750) );
  IV U19130 ( .A(n19746), .Z(n19748) );
  XOR U19131 ( .A(n19752), .B(n19753), .Z(n19746) );
  AND U19132 ( .A(n2062), .B(n19745), .Z(n19753) );
  XNOR U19133 ( .A(n19743), .B(n19752), .Z(n19745) );
  XNOR U19134 ( .A(n19754), .B(n19755), .Z(n19743) );
  AND U19135 ( .A(n2066), .B(n19756), .Z(n19755) );
  XOR U19136 ( .A(p_input[1694]), .B(n19754), .Z(n19756) );
  XNOR U19137 ( .A(n19757), .B(n19758), .Z(n19754) );
  AND U19138 ( .A(n2070), .B(n19759), .Z(n19758) );
  XOR U19139 ( .A(n19760), .B(n19761), .Z(n19752) );
  AND U19140 ( .A(n2074), .B(n19751), .Z(n19761) );
  XNOR U19141 ( .A(n19762), .B(n19749), .Z(n19751) );
  XOR U19142 ( .A(n19763), .B(n19764), .Z(n19749) );
  AND U19143 ( .A(n2097), .B(n19765), .Z(n19764) );
  IV U19144 ( .A(n19760), .Z(n19762) );
  XOR U19145 ( .A(n19766), .B(n19767), .Z(n19760) );
  AND U19146 ( .A(n2081), .B(n19759), .Z(n19767) );
  XNOR U19147 ( .A(n19757), .B(n19766), .Z(n19759) );
  XNOR U19148 ( .A(n19768), .B(n19769), .Z(n19757) );
  AND U19149 ( .A(n2085), .B(n19770), .Z(n19769) );
  XOR U19150 ( .A(p_input[1710]), .B(n19768), .Z(n19770) );
  XNOR U19151 ( .A(n19771), .B(n19772), .Z(n19768) );
  AND U19152 ( .A(n2089), .B(n19773), .Z(n19772) );
  XOR U19153 ( .A(n19774), .B(n19775), .Z(n19766) );
  AND U19154 ( .A(n2093), .B(n19765), .Z(n19775) );
  XNOR U19155 ( .A(n19776), .B(n19763), .Z(n19765) );
  XOR U19156 ( .A(n19777), .B(n19778), .Z(n19763) );
  AND U19157 ( .A(n2116), .B(n19779), .Z(n19778) );
  IV U19158 ( .A(n19774), .Z(n19776) );
  XOR U19159 ( .A(n19780), .B(n19781), .Z(n19774) );
  AND U19160 ( .A(n2100), .B(n19773), .Z(n19781) );
  XNOR U19161 ( .A(n19771), .B(n19780), .Z(n19773) );
  XNOR U19162 ( .A(n19782), .B(n19783), .Z(n19771) );
  AND U19163 ( .A(n2104), .B(n19784), .Z(n19783) );
  XOR U19164 ( .A(p_input[1726]), .B(n19782), .Z(n19784) );
  XNOR U19165 ( .A(n19785), .B(n19786), .Z(n19782) );
  AND U19166 ( .A(n2108), .B(n19787), .Z(n19786) );
  XOR U19167 ( .A(n19788), .B(n19789), .Z(n19780) );
  AND U19168 ( .A(n2112), .B(n19779), .Z(n19789) );
  XNOR U19169 ( .A(n19790), .B(n19777), .Z(n19779) );
  XOR U19170 ( .A(n19791), .B(n19792), .Z(n19777) );
  AND U19171 ( .A(n2135), .B(n19793), .Z(n19792) );
  IV U19172 ( .A(n19788), .Z(n19790) );
  XOR U19173 ( .A(n19794), .B(n19795), .Z(n19788) );
  AND U19174 ( .A(n2119), .B(n19787), .Z(n19795) );
  XNOR U19175 ( .A(n19785), .B(n19794), .Z(n19787) );
  XNOR U19176 ( .A(n19796), .B(n19797), .Z(n19785) );
  AND U19177 ( .A(n2123), .B(n19798), .Z(n19797) );
  XOR U19178 ( .A(p_input[1742]), .B(n19796), .Z(n19798) );
  XNOR U19179 ( .A(n19799), .B(n19800), .Z(n19796) );
  AND U19180 ( .A(n2127), .B(n19801), .Z(n19800) );
  XOR U19181 ( .A(n19802), .B(n19803), .Z(n19794) );
  AND U19182 ( .A(n2131), .B(n19793), .Z(n19803) );
  XNOR U19183 ( .A(n19804), .B(n19791), .Z(n19793) );
  XOR U19184 ( .A(n19805), .B(n19806), .Z(n19791) );
  AND U19185 ( .A(n2154), .B(n19807), .Z(n19806) );
  IV U19186 ( .A(n19802), .Z(n19804) );
  XOR U19187 ( .A(n19808), .B(n19809), .Z(n19802) );
  AND U19188 ( .A(n2138), .B(n19801), .Z(n19809) );
  XNOR U19189 ( .A(n19799), .B(n19808), .Z(n19801) );
  XNOR U19190 ( .A(n19810), .B(n19811), .Z(n19799) );
  AND U19191 ( .A(n2142), .B(n19812), .Z(n19811) );
  XOR U19192 ( .A(p_input[1758]), .B(n19810), .Z(n19812) );
  XNOR U19193 ( .A(n19813), .B(n19814), .Z(n19810) );
  AND U19194 ( .A(n2146), .B(n19815), .Z(n19814) );
  XOR U19195 ( .A(n19816), .B(n19817), .Z(n19808) );
  AND U19196 ( .A(n2150), .B(n19807), .Z(n19817) );
  XNOR U19197 ( .A(n19818), .B(n19805), .Z(n19807) );
  XOR U19198 ( .A(n19819), .B(n19820), .Z(n19805) );
  AND U19199 ( .A(n2173), .B(n19821), .Z(n19820) );
  IV U19200 ( .A(n19816), .Z(n19818) );
  XOR U19201 ( .A(n19822), .B(n19823), .Z(n19816) );
  AND U19202 ( .A(n2157), .B(n19815), .Z(n19823) );
  XNOR U19203 ( .A(n19813), .B(n19822), .Z(n19815) );
  XNOR U19204 ( .A(n19824), .B(n19825), .Z(n19813) );
  AND U19205 ( .A(n2161), .B(n19826), .Z(n19825) );
  XOR U19206 ( .A(p_input[1774]), .B(n19824), .Z(n19826) );
  XNOR U19207 ( .A(n19827), .B(n19828), .Z(n19824) );
  AND U19208 ( .A(n2165), .B(n19829), .Z(n19828) );
  XOR U19209 ( .A(n19830), .B(n19831), .Z(n19822) );
  AND U19210 ( .A(n2169), .B(n19821), .Z(n19831) );
  XNOR U19211 ( .A(n19832), .B(n19819), .Z(n19821) );
  XOR U19212 ( .A(n19833), .B(n19834), .Z(n19819) );
  AND U19213 ( .A(n2192), .B(n19835), .Z(n19834) );
  IV U19214 ( .A(n19830), .Z(n19832) );
  XOR U19215 ( .A(n19836), .B(n19837), .Z(n19830) );
  AND U19216 ( .A(n2176), .B(n19829), .Z(n19837) );
  XNOR U19217 ( .A(n19827), .B(n19836), .Z(n19829) );
  XNOR U19218 ( .A(n19838), .B(n19839), .Z(n19827) );
  AND U19219 ( .A(n2180), .B(n19840), .Z(n19839) );
  XOR U19220 ( .A(p_input[1790]), .B(n19838), .Z(n19840) );
  XNOR U19221 ( .A(n19841), .B(n19842), .Z(n19838) );
  AND U19222 ( .A(n2184), .B(n19843), .Z(n19842) );
  XOR U19223 ( .A(n19844), .B(n19845), .Z(n19836) );
  AND U19224 ( .A(n2188), .B(n19835), .Z(n19845) );
  XNOR U19225 ( .A(n19846), .B(n19833), .Z(n19835) );
  XOR U19226 ( .A(n19847), .B(n19848), .Z(n19833) );
  AND U19227 ( .A(n2211), .B(n19849), .Z(n19848) );
  IV U19228 ( .A(n19844), .Z(n19846) );
  XOR U19229 ( .A(n19850), .B(n19851), .Z(n19844) );
  AND U19230 ( .A(n2195), .B(n19843), .Z(n19851) );
  XNOR U19231 ( .A(n19841), .B(n19850), .Z(n19843) );
  XNOR U19232 ( .A(n19852), .B(n19853), .Z(n19841) );
  AND U19233 ( .A(n2199), .B(n19854), .Z(n19853) );
  XOR U19234 ( .A(p_input[1806]), .B(n19852), .Z(n19854) );
  XNOR U19235 ( .A(n19855), .B(n19856), .Z(n19852) );
  AND U19236 ( .A(n2203), .B(n19857), .Z(n19856) );
  XOR U19237 ( .A(n19858), .B(n19859), .Z(n19850) );
  AND U19238 ( .A(n2207), .B(n19849), .Z(n19859) );
  XNOR U19239 ( .A(n19860), .B(n19847), .Z(n19849) );
  XOR U19240 ( .A(n19861), .B(n19862), .Z(n19847) );
  AND U19241 ( .A(n2230), .B(n19863), .Z(n19862) );
  IV U19242 ( .A(n19858), .Z(n19860) );
  XOR U19243 ( .A(n19864), .B(n19865), .Z(n19858) );
  AND U19244 ( .A(n2214), .B(n19857), .Z(n19865) );
  XNOR U19245 ( .A(n19855), .B(n19864), .Z(n19857) );
  XNOR U19246 ( .A(n19866), .B(n19867), .Z(n19855) );
  AND U19247 ( .A(n2218), .B(n19868), .Z(n19867) );
  XOR U19248 ( .A(p_input[1822]), .B(n19866), .Z(n19868) );
  XNOR U19249 ( .A(n19869), .B(n19870), .Z(n19866) );
  AND U19250 ( .A(n2222), .B(n19871), .Z(n19870) );
  XOR U19251 ( .A(n19872), .B(n19873), .Z(n19864) );
  AND U19252 ( .A(n2226), .B(n19863), .Z(n19873) );
  XNOR U19253 ( .A(n19874), .B(n19861), .Z(n19863) );
  XOR U19254 ( .A(n19875), .B(n19876), .Z(n19861) );
  AND U19255 ( .A(n2249), .B(n19877), .Z(n19876) );
  IV U19256 ( .A(n19872), .Z(n19874) );
  XOR U19257 ( .A(n19878), .B(n19879), .Z(n19872) );
  AND U19258 ( .A(n2233), .B(n19871), .Z(n19879) );
  XNOR U19259 ( .A(n19869), .B(n19878), .Z(n19871) );
  XNOR U19260 ( .A(n19880), .B(n19881), .Z(n19869) );
  AND U19261 ( .A(n2237), .B(n19882), .Z(n19881) );
  XOR U19262 ( .A(p_input[1838]), .B(n19880), .Z(n19882) );
  XNOR U19263 ( .A(n19883), .B(n19884), .Z(n19880) );
  AND U19264 ( .A(n2241), .B(n19885), .Z(n19884) );
  XOR U19265 ( .A(n19886), .B(n19887), .Z(n19878) );
  AND U19266 ( .A(n2245), .B(n19877), .Z(n19887) );
  XNOR U19267 ( .A(n19888), .B(n19875), .Z(n19877) );
  XOR U19268 ( .A(n19889), .B(n19890), .Z(n19875) );
  AND U19269 ( .A(n2268), .B(n19891), .Z(n19890) );
  IV U19270 ( .A(n19886), .Z(n19888) );
  XOR U19271 ( .A(n19892), .B(n19893), .Z(n19886) );
  AND U19272 ( .A(n2252), .B(n19885), .Z(n19893) );
  XNOR U19273 ( .A(n19883), .B(n19892), .Z(n19885) );
  XNOR U19274 ( .A(n19894), .B(n19895), .Z(n19883) );
  AND U19275 ( .A(n2256), .B(n19896), .Z(n19895) );
  XOR U19276 ( .A(p_input[1854]), .B(n19894), .Z(n19896) );
  XNOR U19277 ( .A(n19897), .B(n19898), .Z(n19894) );
  AND U19278 ( .A(n2260), .B(n19899), .Z(n19898) );
  XOR U19279 ( .A(n19900), .B(n19901), .Z(n19892) );
  AND U19280 ( .A(n2264), .B(n19891), .Z(n19901) );
  XNOR U19281 ( .A(n19902), .B(n19889), .Z(n19891) );
  XOR U19282 ( .A(n19903), .B(n19904), .Z(n19889) );
  AND U19283 ( .A(n2287), .B(n19905), .Z(n19904) );
  IV U19284 ( .A(n19900), .Z(n19902) );
  XOR U19285 ( .A(n19906), .B(n19907), .Z(n19900) );
  AND U19286 ( .A(n2271), .B(n19899), .Z(n19907) );
  XNOR U19287 ( .A(n19897), .B(n19906), .Z(n19899) );
  XNOR U19288 ( .A(n19908), .B(n19909), .Z(n19897) );
  AND U19289 ( .A(n2275), .B(n19910), .Z(n19909) );
  XOR U19290 ( .A(p_input[1870]), .B(n19908), .Z(n19910) );
  XNOR U19291 ( .A(n19911), .B(n19912), .Z(n19908) );
  AND U19292 ( .A(n2279), .B(n19913), .Z(n19912) );
  XOR U19293 ( .A(n19914), .B(n19915), .Z(n19906) );
  AND U19294 ( .A(n2283), .B(n19905), .Z(n19915) );
  XNOR U19295 ( .A(n19916), .B(n19903), .Z(n19905) );
  XOR U19296 ( .A(n19917), .B(n19918), .Z(n19903) );
  AND U19297 ( .A(n2306), .B(n19919), .Z(n19918) );
  IV U19298 ( .A(n19914), .Z(n19916) );
  XOR U19299 ( .A(n19920), .B(n19921), .Z(n19914) );
  AND U19300 ( .A(n2290), .B(n19913), .Z(n19921) );
  XNOR U19301 ( .A(n19911), .B(n19920), .Z(n19913) );
  XNOR U19302 ( .A(n19922), .B(n19923), .Z(n19911) );
  AND U19303 ( .A(n2294), .B(n19924), .Z(n19923) );
  XOR U19304 ( .A(p_input[1886]), .B(n19922), .Z(n19924) );
  XNOR U19305 ( .A(n19925), .B(n19926), .Z(n19922) );
  AND U19306 ( .A(n2298), .B(n19927), .Z(n19926) );
  XOR U19307 ( .A(n19928), .B(n19929), .Z(n19920) );
  AND U19308 ( .A(n2302), .B(n19919), .Z(n19929) );
  XNOR U19309 ( .A(n19930), .B(n19917), .Z(n19919) );
  XOR U19310 ( .A(n19931), .B(n19932), .Z(n19917) );
  AND U19311 ( .A(n2325), .B(n19933), .Z(n19932) );
  IV U19312 ( .A(n19928), .Z(n19930) );
  XOR U19313 ( .A(n19934), .B(n19935), .Z(n19928) );
  AND U19314 ( .A(n2309), .B(n19927), .Z(n19935) );
  XNOR U19315 ( .A(n19925), .B(n19934), .Z(n19927) );
  XNOR U19316 ( .A(n19936), .B(n19937), .Z(n19925) );
  AND U19317 ( .A(n2313), .B(n19938), .Z(n19937) );
  XOR U19318 ( .A(p_input[1902]), .B(n19936), .Z(n19938) );
  XNOR U19319 ( .A(n19939), .B(n19940), .Z(n19936) );
  AND U19320 ( .A(n2317), .B(n19941), .Z(n19940) );
  XOR U19321 ( .A(n19942), .B(n19943), .Z(n19934) );
  AND U19322 ( .A(n2321), .B(n19933), .Z(n19943) );
  XNOR U19323 ( .A(n19944), .B(n19931), .Z(n19933) );
  XOR U19324 ( .A(n19945), .B(n19946), .Z(n19931) );
  AND U19325 ( .A(n2344), .B(n19947), .Z(n19946) );
  IV U19326 ( .A(n19942), .Z(n19944) );
  XOR U19327 ( .A(n19948), .B(n19949), .Z(n19942) );
  AND U19328 ( .A(n2328), .B(n19941), .Z(n19949) );
  XNOR U19329 ( .A(n19939), .B(n19948), .Z(n19941) );
  XNOR U19330 ( .A(n19950), .B(n19951), .Z(n19939) );
  AND U19331 ( .A(n2332), .B(n19952), .Z(n19951) );
  XOR U19332 ( .A(p_input[1918]), .B(n19950), .Z(n19952) );
  XNOR U19333 ( .A(n19953), .B(n19954), .Z(n19950) );
  AND U19334 ( .A(n2336), .B(n19955), .Z(n19954) );
  XOR U19335 ( .A(n19956), .B(n19957), .Z(n19948) );
  AND U19336 ( .A(n2340), .B(n19947), .Z(n19957) );
  XNOR U19337 ( .A(n19958), .B(n19945), .Z(n19947) );
  XOR U19338 ( .A(n19959), .B(n19960), .Z(n19945) );
  AND U19339 ( .A(n2363), .B(n19961), .Z(n19960) );
  IV U19340 ( .A(n19956), .Z(n19958) );
  XOR U19341 ( .A(n19962), .B(n19963), .Z(n19956) );
  AND U19342 ( .A(n2347), .B(n19955), .Z(n19963) );
  XNOR U19343 ( .A(n19953), .B(n19962), .Z(n19955) );
  XNOR U19344 ( .A(n19964), .B(n19965), .Z(n19953) );
  AND U19345 ( .A(n2351), .B(n19966), .Z(n19965) );
  XOR U19346 ( .A(p_input[1934]), .B(n19964), .Z(n19966) );
  XNOR U19347 ( .A(n19967), .B(n19968), .Z(n19964) );
  AND U19348 ( .A(n2355), .B(n19969), .Z(n19968) );
  XOR U19349 ( .A(n19970), .B(n19971), .Z(n19962) );
  AND U19350 ( .A(n2359), .B(n19961), .Z(n19971) );
  XNOR U19351 ( .A(n19972), .B(n19959), .Z(n19961) );
  XOR U19352 ( .A(n19973), .B(n19974), .Z(n19959) );
  AND U19353 ( .A(n2382), .B(n19975), .Z(n19974) );
  IV U19354 ( .A(n19970), .Z(n19972) );
  XOR U19355 ( .A(n19976), .B(n19977), .Z(n19970) );
  AND U19356 ( .A(n2366), .B(n19969), .Z(n19977) );
  XNOR U19357 ( .A(n19967), .B(n19976), .Z(n19969) );
  XNOR U19358 ( .A(n19978), .B(n19979), .Z(n19967) );
  AND U19359 ( .A(n2370), .B(n19980), .Z(n19979) );
  XOR U19360 ( .A(p_input[1950]), .B(n19978), .Z(n19980) );
  XNOR U19361 ( .A(n19981), .B(n19982), .Z(n19978) );
  AND U19362 ( .A(n2374), .B(n19983), .Z(n19982) );
  XOR U19363 ( .A(n19984), .B(n19985), .Z(n19976) );
  AND U19364 ( .A(n2378), .B(n19975), .Z(n19985) );
  XNOR U19365 ( .A(n19986), .B(n19973), .Z(n19975) );
  XOR U19366 ( .A(n19987), .B(n19988), .Z(n19973) );
  AND U19367 ( .A(n2401), .B(n19989), .Z(n19988) );
  IV U19368 ( .A(n19984), .Z(n19986) );
  XOR U19369 ( .A(n19990), .B(n19991), .Z(n19984) );
  AND U19370 ( .A(n2385), .B(n19983), .Z(n19991) );
  XNOR U19371 ( .A(n19981), .B(n19990), .Z(n19983) );
  XNOR U19372 ( .A(n19992), .B(n19993), .Z(n19981) );
  AND U19373 ( .A(n2389), .B(n19994), .Z(n19993) );
  XOR U19374 ( .A(p_input[1966]), .B(n19992), .Z(n19994) );
  XNOR U19375 ( .A(n19995), .B(n19996), .Z(n19992) );
  AND U19376 ( .A(n2393), .B(n19997), .Z(n19996) );
  XOR U19377 ( .A(n19998), .B(n19999), .Z(n19990) );
  AND U19378 ( .A(n2397), .B(n19989), .Z(n19999) );
  XNOR U19379 ( .A(n20000), .B(n19987), .Z(n19989) );
  XOR U19380 ( .A(n20001), .B(n20002), .Z(n19987) );
  AND U19381 ( .A(n2420), .B(n20003), .Z(n20002) );
  IV U19382 ( .A(n19998), .Z(n20000) );
  XOR U19383 ( .A(n20004), .B(n20005), .Z(n19998) );
  AND U19384 ( .A(n2404), .B(n19997), .Z(n20005) );
  XNOR U19385 ( .A(n19995), .B(n20004), .Z(n19997) );
  XNOR U19386 ( .A(n20006), .B(n20007), .Z(n19995) );
  AND U19387 ( .A(n2408), .B(n20008), .Z(n20007) );
  XOR U19388 ( .A(p_input[1982]), .B(n20006), .Z(n20008) );
  XNOR U19389 ( .A(n20009), .B(n20010), .Z(n20006) );
  AND U19390 ( .A(n2412), .B(n20011), .Z(n20010) );
  XOR U19391 ( .A(n20012), .B(n20013), .Z(n20004) );
  AND U19392 ( .A(n2416), .B(n20003), .Z(n20013) );
  XNOR U19393 ( .A(n20014), .B(n20001), .Z(n20003) );
  XOR U19394 ( .A(n20015), .B(n20016), .Z(n20001) );
  AND U19395 ( .A(n2438), .B(n20017), .Z(n20016) );
  IV U19396 ( .A(n20012), .Z(n20014) );
  XOR U19397 ( .A(n20018), .B(n20019), .Z(n20012) );
  AND U19398 ( .A(n2423), .B(n20011), .Z(n20019) );
  XNOR U19399 ( .A(n20009), .B(n20018), .Z(n20011) );
  XNOR U19400 ( .A(n20020), .B(n20021), .Z(n20009) );
  AND U19401 ( .A(n2427), .B(n20022), .Z(n20021) );
  XOR U19402 ( .A(p_input[1998]), .B(n20020), .Z(n20022) );
  XOR U19403 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n20023), 
        .Z(n20020) );
  AND U19404 ( .A(n2430), .B(n20024), .Z(n20023) );
  XOR U19405 ( .A(n20025), .B(n20026), .Z(n20018) );
  AND U19406 ( .A(n2434), .B(n20017), .Z(n20026) );
  XNOR U19407 ( .A(n20027), .B(n20015), .Z(n20017) );
  XOR U19408 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n20028), .Z(n20015) );
  AND U19409 ( .A(n2446), .B(n20029), .Z(n20028) );
  IV U19410 ( .A(n20025), .Z(n20027) );
  XOR U19411 ( .A(n20030), .B(n20031), .Z(n20025) );
  AND U19412 ( .A(n2441), .B(n20024), .Z(n20031) );
  XOR U19413 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n20030), 
        .Z(n20024) );
  XOR U19414 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n20032), 
        .Z(n20030) );
  AND U19415 ( .A(n2443), .B(n20029), .Z(n20032) );
  XOR U19416 ( .A(n20033), .B(n20034), .Z(n20029) );
  IV U19417 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n20034)
         );
  IV U19418 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n20033) );
  XOR U19419 ( .A(n53), .B(n20035), .Z(o[13]) );
  AND U19420 ( .A(n62), .B(n20036), .Z(n53) );
  XOR U19421 ( .A(n54), .B(n20035), .Z(n20036) );
  XOR U19422 ( .A(n20037), .B(n20038), .Z(n20035) );
  AND U19423 ( .A(n82), .B(n20039), .Z(n20038) );
  XOR U19424 ( .A(n20040), .B(n17), .Z(n54) );
  AND U19425 ( .A(n65), .B(n20041), .Z(n17) );
  XOR U19426 ( .A(n18), .B(n20040), .Z(n20041) );
  XOR U19427 ( .A(n20042), .B(n20043), .Z(n18) );
  AND U19428 ( .A(n70), .B(n20044), .Z(n20043) );
  XOR U19429 ( .A(p_input[13]), .B(n20042), .Z(n20044) );
  XNOR U19430 ( .A(n20045), .B(n20046), .Z(n20042) );
  AND U19431 ( .A(n74), .B(n20047), .Z(n20046) );
  XOR U19432 ( .A(n20048), .B(n20049), .Z(n20040) );
  AND U19433 ( .A(n78), .B(n20039), .Z(n20049) );
  XNOR U19434 ( .A(n20050), .B(n20037), .Z(n20039) );
  XOR U19435 ( .A(n20051), .B(n20052), .Z(n20037) );
  AND U19436 ( .A(n102), .B(n20053), .Z(n20052) );
  IV U19437 ( .A(n20048), .Z(n20050) );
  XOR U19438 ( .A(n20054), .B(n20055), .Z(n20048) );
  AND U19439 ( .A(n86), .B(n20047), .Z(n20055) );
  XNOR U19440 ( .A(n20045), .B(n20054), .Z(n20047) );
  XNOR U19441 ( .A(n20056), .B(n20057), .Z(n20045) );
  AND U19442 ( .A(n90), .B(n20058), .Z(n20057) );
  XOR U19443 ( .A(p_input[29]), .B(n20056), .Z(n20058) );
  XNOR U19444 ( .A(n20059), .B(n20060), .Z(n20056) );
  AND U19445 ( .A(n94), .B(n20061), .Z(n20060) );
  XOR U19446 ( .A(n20062), .B(n20063), .Z(n20054) );
  AND U19447 ( .A(n98), .B(n20053), .Z(n20063) );
  XNOR U19448 ( .A(n20064), .B(n20051), .Z(n20053) );
  XOR U19449 ( .A(n20065), .B(n20066), .Z(n20051) );
  AND U19450 ( .A(n121), .B(n20067), .Z(n20066) );
  IV U19451 ( .A(n20062), .Z(n20064) );
  XOR U19452 ( .A(n20068), .B(n20069), .Z(n20062) );
  AND U19453 ( .A(n105), .B(n20061), .Z(n20069) );
  XNOR U19454 ( .A(n20059), .B(n20068), .Z(n20061) );
  XNOR U19455 ( .A(n20070), .B(n20071), .Z(n20059) );
  AND U19456 ( .A(n109), .B(n20072), .Z(n20071) );
  XOR U19457 ( .A(p_input[45]), .B(n20070), .Z(n20072) );
  XNOR U19458 ( .A(n20073), .B(n20074), .Z(n20070) );
  AND U19459 ( .A(n113), .B(n20075), .Z(n20074) );
  XOR U19460 ( .A(n20076), .B(n20077), .Z(n20068) );
  AND U19461 ( .A(n117), .B(n20067), .Z(n20077) );
  XNOR U19462 ( .A(n20078), .B(n20065), .Z(n20067) );
  XOR U19463 ( .A(n20079), .B(n20080), .Z(n20065) );
  AND U19464 ( .A(n140), .B(n20081), .Z(n20080) );
  IV U19465 ( .A(n20076), .Z(n20078) );
  XOR U19466 ( .A(n20082), .B(n20083), .Z(n20076) );
  AND U19467 ( .A(n124), .B(n20075), .Z(n20083) );
  XNOR U19468 ( .A(n20073), .B(n20082), .Z(n20075) );
  XNOR U19469 ( .A(n20084), .B(n20085), .Z(n20073) );
  AND U19470 ( .A(n128), .B(n20086), .Z(n20085) );
  XOR U19471 ( .A(p_input[61]), .B(n20084), .Z(n20086) );
  XNOR U19472 ( .A(n20087), .B(n20088), .Z(n20084) );
  AND U19473 ( .A(n132), .B(n20089), .Z(n20088) );
  XOR U19474 ( .A(n20090), .B(n20091), .Z(n20082) );
  AND U19475 ( .A(n136), .B(n20081), .Z(n20091) );
  XNOR U19476 ( .A(n20092), .B(n20079), .Z(n20081) );
  XOR U19477 ( .A(n20093), .B(n20094), .Z(n20079) );
  AND U19478 ( .A(n159), .B(n20095), .Z(n20094) );
  IV U19479 ( .A(n20090), .Z(n20092) );
  XOR U19480 ( .A(n20096), .B(n20097), .Z(n20090) );
  AND U19481 ( .A(n143), .B(n20089), .Z(n20097) );
  XNOR U19482 ( .A(n20087), .B(n20096), .Z(n20089) );
  XNOR U19483 ( .A(n20098), .B(n20099), .Z(n20087) );
  AND U19484 ( .A(n147), .B(n20100), .Z(n20099) );
  XOR U19485 ( .A(p_input[77]), .B(n20098), .Z(n20100) );
  XNOR U19486 ( .A(n20101), .B(n20102), .Z(n20098) );
  AND U19487 ( .A(n151), .B(n20103), .Z(n20102) );
  XOR U19488 ( .A(n20104), .B(n20105), .Z(n20096) );
  AND U19489 ( .A(n155), .B(n20095), .Z(n20105) );
  XNOR U19490 ( .A(n20106), .B(n20093), .Z(n20095) );
  XOR U19491 ( .A(n20107), .B(n20108), .Z(n20093) );
  AND U19492 ( .A(n178), .B(n20109), .Z(n20108) );
  IV U19493 ( .A(n20104), .Z(n20106) );
  XOR U19494 ( .A(n20110), .B(n20111), .Z(n20104) );
  AND U19495 ( .A(n162), .B(n20103), .Z(n20111) );
  XNOR U19496 ( .A(n20101), .B(n20110), .Z(n20103) );
  XNOR U19497 ( .A(n20112), .B(n20113), .Z(n20101) );
  AND U19498 ( .A(n166), .B(n20114), .Z(n20113) );
  XOR U19499 ( .A(p_input[93]), .B(n20112), .Z(n20114) );
  XNOR U19500 ( .A(n20115), .B(n20116), .Z(n20112) );
  AND U19501 ( .A(n170), .B(n20117), .Z(n20116) );
  XOR U19502 ( .A(n20118), .B(n20119), .Z(n20110) );
  AND U19503 ( .A(n174), .B(n20109), .Z(n20119) );
  XNOR U19504 ( .A(n20120), .B(n20107), .Z(n20109) );
  XOR U19505 ( .A(n20121), .B(n20122), .Z(n20107) );
  AND U19506 ( .A(n197), .B(n20123), .Z(n20122) );
  IV U19507 ( .A(n20118), .Z(n20120) );
  XOR U19508 ( .A(n20124), .B(n20125), .Z(n20118) );
  AND U19509 ( .A(n181), .B(n20117), .Z(n20125) );
  XNOR U19510 ( .A(n20115), .B(n20124), .Z(n20117) );
  XNOR U19511 ( .A(n20126), .B(n20127), .Z(n20115) );
  AND U19512 ( .A(n185), .B(n20128), .Z(n20127) );
  XOR U19513 ( .A(p_input[109]), .B(n20126), .Z(n20128) );
  XNOR U19514 ( .A(n20129), .B(n20130), .Z(n20126) );
  AND U19515 ( .A(n189), .B(n20131), .Z(n20130) );
  XOR U19516 ( .A(n20132), .B(n20133), .Z(n20124) );
  AND U19517 ( .A(n193), .B(n20123), .Z(n20133) );
  XNOR U19518 ( .A(n20134), .B(n20121), .Z(n20123) );
  XOR U19519 ( .A(n20135), .B(n20136), .Z(n20121) );
  AND U19520 ( .A(n216), .B(n20137), .Z(n20136) );
  IV U19521 ( .A(n20132), .Z(n20134) );
  XOR U19522 ( .A(n20138), .B(n20139), .Z(n20132) );
  AND U19523 ( .A(n200), .B(n20131), .Z(n20139) );
  XNOR U19524 ( .A(n20129), .B(n20138), .Z(n20131) );
  XNOR U19525 ( .A(n20140), .B(n20141), .Z(n20129) );
  AND U19526 ( .A(n204), .B(n20142), .Z(n20141) );
  XOR U19527 ( .A(p_input[125]), .B(n20140), .Z(n20142) );
  XNOR U19528 ( .A(n20143), .B(n20144), .Z(n20140) );
  AND U19529 ( .A(n208), .B(n20145), .Z(n20144) );
  XOR U19530 ( .A(n20146), .B(n20147), .Z(n20138) );
  AND U19531 ( .A(n212), .B(n20137), .Z(n20147) );
  XNOR U19532 ( .A(n20148), .B(n20135), .Z(n20137) );
  XOR U19533 ( .A(n20149), .B(n20150), .Z(n20135) );
  AND U19534 ( .A(n235), .B(n20151), .Z(n20150) );
  IV U19535 ( .A(n20146), .Z(n20148) );
  XOR U19536 ( .A(n20152), .B(n20153), .Z(n20146) );
  AND U19537 ( .A(n219), .B(n20145), .Z(n20153) );
  XNOR U19538 ( .A(n20143), .B(n20152), .Z(n20145) );
  XNOR U19539 ( .A(n20154), .B(n20155), .Z(n20143) );
  AND U19540 ( .A(n223), .B(n20156), .Z(n20155) );
  XOR U19541 ( .A(p_input[141]), .B(n20154), .Z(n20156) );
  XNOR U19542 ( .A(n20157), .B(n20158), .Z(n20154) );
  AND U19543 ( .A(n227), .B(n20159), .Z(n20158) );
  XOR U19544 ( .A(n20160), .B(n20161), .Z(n20152) );
  AND U19545 ( .A(n231), .B(n20151), .Z(n20161) );
  XNOR U19546 ( .A(n20162), .B(n20149), .Z(n20151) );
  XOR U19547 ( .A(n20163), .B(n20164), .Z(n20149) );
  AND U19548 ( .A(n254), .B(n20165), .Z(n20164) );
  IV U19549 ( .A(n20160), .Z(n20162) );
  XOR U19550 ( .A(n20166), .B(n20167), .Z(n20160) );
  AND U19551 ( .A(n238), .B(n20159), .Z(n20167) );
  XNOR U19552 ( .A(n20157), .B(n20166), .Z(n20159) );
  XNOR U19553 ( .A(n20168), .B(n20169), .Z(n20157) );
  AND U19554 ( .A(n242), .B(n20170), .Z(n20169) );
  XOR U19555 ( .A(p_input[157]), .B(n20168), .Z(n20170) );
  XNOR U19556 ( .A(n20171), .B(n20172), .Z(n20168) );
  AND U19557 ( .A(n246), .B(n20173), .Z(n20172) );
  XOR U19558 ( .A(n20174), .B(n20175), .Z(n20166) );
  AND U19559 ( .A(n250), .B(n20165), .Z(n20175) );
  XNOR U19560 ( .A(n20176), .B(n20163), .Z(n20165) );
  XOR U19561 ( .A(n20177), .B(n20178), .Z(n20163) );
  AND U19562 ( .A(n273), .B(n20179), .Z(n20178) );
  IV U19563 ( .A(n20174), .Z(n20176) );
  XOR U19564 ( .A(n20180), .B(n20181), .Z(n20174) );
  AND U19565 ( .A(n257), .B(n20173), .Z(n20181) );
  XNOR U19566 ( .A(n20171), .B(n20180), .Z(n20173) );
  XNOR U19567 ( .A(n20182), .B(n20183), .Z(n20171) );
  AND U19568 ( .A(n261), .B(n20184), .Z(n20183) );
  XOR U19569 ( .A(p_input[173]), .B(n20182), .Z(n20184) );
  XNOR U19570 ( .A(n20185), .B(n20186), .Z(n20182) );
  AND U19571 ( .A(n265), .B(n20187), .Z(n20186) );
  XOR U19572 ( .A(n20188), .B(n20189), .Z(n20180) );
  AND U19573 ( .A(n269), .B(n20179), .Z(n20189) );
  XNOR U19574 ( .A(n20190), .B(n20177), .Z(n20179) );
  XOR U19575 ( .A(n20191), .B(n20192), .Z(n20177) );
  AND U19576 ( .A(n292), .B(n20193), .Z(n20192) );
  IV U19577 ( .A(n20188), .Z(n20190) );
  XOR U19578 ( .A(n20194), .B(n20195), .Z(n20188) );
  AND U19579 ( .A(n276), .B(n20187), .Z(n20195) );
  XNOR U19580 ( .A(n20185), .B(n20194), .Z(n20187) );
  XNOR U19581 ( .A(n20196), .B(n20197), .Z(n20185) );
  AND U19582 ( .A(n280), .B(n20198), .Z(n20197) );
  XOR U19583 ( .A(p_input[189]), .B(n20196), .Z(n20198) );
  XNOR U19584 ( .A(n20199), .B(n20200), .Z(n20196) );
  AND U19585 ( .A(n284), .B(n20201), .Z(n20200) );
  XOR U19586 ( .A(n20202), .B(n20203), .Z(n20194) );
  AND U19587 ( .A(n288), .B(n20193), .Z(n20203) );
  XNOR U19588 ( .A(n20204), .B(n20191), .Z(n20193) );
  XOR U19589 ( .A(n20205), .B(n20206), .Z(n20191) );
  AND U19590 ( .A(n311), .B(n20207), .Z(n20206) );
  IV U19591 ( .A(n20202), .Z(n20204) );
  XOR U19592 ( .A(n20208), .B(n20209), .Z(n20202) );
  AND U19593 ( .A(n295), .B(n20201), .Z(n20209) );
  XNOR U19594 ( .A(n20199), .B(n20208), .Z(n20201) );
  XNOR U19595 ( .A(n20210), .B(n20211), .Z(n20199) );
  AND U19596 ( .A(n299), .B(n20212), .Z(n20211) );
  XOR U19597 ( .A(p_input[205]), .B(n20210), .Z(n20212) );
  XNOR U19598 ( .A(n20213), .B(n20214), .Z(n20210) );
  AND U19599 ( .A(n303), .B(n20215), .Z(n20214) );
  XOR U19600 ( .A(n20216), .B(n20217), .Z(n20208) );
  AND U19601 ( .A(n307), .B(n20207), .Z(n20217) );
  XNOR U19602 ( .A(n20218), .B(n20205), .Z(n20207) );
  XOR U19603 ( .A(n20219), .B(n20220), .Z(n20205) );
  AND U19604 ( .A(n330), .B(n20221), .Z(n20220) );
  IV U19605 ( .A(n20216), .Z(n20218) );
  XOR U19606 ( .A(n20222), .B(n20223), .Z(n20216) );
  AND U19607 ( .A(n314), .B(n20215), .Z(n20223) );
  XNOR U19608 ( .A(n20213), .B(n20222), .Z(n20215) );
  XNOR U19609 ( .A(n20224), .B(n20225), .Z(n20213) );
  AND U19610 ( .A(n318), .B(n20226), .Z(n20225) );
  XOR U19611 ( .A(p_input[221]), .B(n20224), .Z(n20226) );
  XNOR U19612 ( .A(n20227), .B(n20228), .Z(n20224) );
  AND U19613 ( .A(n322), .B(n20229), .Z(n20228) );
  XOR U19614 ( .A(n20230), .B(n20231), .Z(n20222) );
  AND U19615 ( .A(n326), .B(n20221), .Z(n20231) );
  XNOR U19616 ( .A(n20232), .B(n20219), .Z(n20221) );
  XOR U19617 ( .A(n20233), .B(n20234), .Z(n20219) );
  AND U19618 ( .A(n349), .B(n20235), .Z(n20234) );
  IV U19619 ( .A(n20230), .Z(n20232) );
  XOR U19620 ( .A(n20236), .B(n20237), .Z(n20230) );
  AND U19621 ( .A(n333), .B(n20229), .Z(n20237) );
  XNOR U19622 ( .A(n20227), .B(n20236), .Z(n20229) );
  XNOR U19623 ( .A(n20238), .B(n20239), .Z(n20227) );
  AND U19624 ( .A(n337), .B(n20240), .Z(n20239) );
  XOR U19625 ( .A(p_input[237]), .B(n20238), .Z(n20240) );
  XNOR U19626 ( .A(n20241), .B(n20242), .Z(n20238) );
  AND U19627 ( .A(n341), .B(n20243), .Z(n20242) );
  XOR U19628 ( .A(n20244), .B(n20245), .Z(n20236) );
  AND U19629 ( .A(n345), .B(n20235), .Z(n20245) );
  XNOR U19630 ( .A(n20246), .B(n20233), .Z(n20235) );
  XOR U19631 ( .A(n20247), .B(n20248), .Z(n20233) );
  AND U19632 ( .A(n368), .B(n20249), .Z(n20248) );
  IV U19633 ( .A(n20244), .Z(n20246) );
  XOR U19634 ( .A(n20250), .B(n20251), .Z(n20244) );
  AND U19635 ( .A(n352), .B(n20243), .Z(n20251) );
  XNOR U19636 ( .A(n20241), .B(n20250), .Z(n20243) );
  XNOR U19637 ( .A(n20252), .B(n20253), .Z(n20241) );
  AND U19638 ( .A(n356), .B(n20254), .Z(n20253) );
  XOR U19639 ( .A(p_input[253]), .B(n20252), .Z(n20254) );
  XNOR U19640 ( .A(n20255), .B(n20256), .Z(n20252) );
  AND U19641 ( .A(n360), .B(n20257), .Z(n20256) );
  XOR U19642 ( .A(n20258), .B(n20259), .Z(n20250) );
  AND U19643 ( .A(n364), .B(n20249), .Z(n20259) );
  XNOR U19644 ( .A(n20260), .B(n20247), .Z(n20249) );
  XOR U19645 ( .A(n20261), .B(n20262), .Z(n20247) );
  AND U19646 ( .A(n387), .B(n20263), .Z(n20262) );
  IV U19647 ( .A(n20258), .Z(n20260) );
  XOR U19648 ( .A(n20264), .B(n20265), .Z(n20258) );
  AND U19649 ( .A(n371), .B(n20257), .Z(n20265) );
  XNOR U19650 ( .A(n20255), .B(n20264), .Z(n20257) );
  XNOR U19651 ( .A(n20266), .B(n20267), .Z(n20255) );
  AND U19652 ( .A(n375), .B(n20268), .Z(n20267) );
  XOR U19653 ( .A(p_input[269]), .B(n20266), .Z(n20268) );
  XNOR U19654 ( .A(n20269), .B(n20270), .Z(n20266) );
  AND U19655 ( .A(n379), .B(n20271), .Z(n20270) );
  XOR U19656 ( .A(n20272), .B(n20273), .Z(n20264) );
  AND U19657 ( .A(n383), .B(n20263), .Z(n20273) );
  XNOR U19658 ( .A(n20274), .B(n20261), .Z(n20263) );
  XOR U19659 ( .A(n20275), .B(n20276), .Z(n20261) );
  AND U19660 ( .A(n406), .B(n20277), .Z(n20276) );
  IV U19661 ( .A(n20272), .Z(n20274) );
  XOR U19662 ( .A(n20278), .B(n20279), .Z(n20272) );
  AND U19663 ( .A(n390), .B(n20271), .Z(n20279) );
  XNOR U19664 ( .A(n20269), .B(n20278), .Z(n20271) );
  XNOR U19665 ( .A(n20280), .B(n20281), .Z(n20269) );
  AND U19666 ( .A(n394), .B(n20282), .Z(n20281) );
  XOR U19667 ( .A(p_input[285]), .B(n20280), .Z(n20282) );
  XNOR U19668 ( .A(n20283), .B(n20284), .Z(n20280) );
  AND U19669 ( .A(n398), .B(n20285), .Z(n20284) );
  XOR U19670 ( .A(n20286), .B(n20287), .Z(n20278) );
  AND U19671 ( .A(n402), .B(n20277), .Z(n20287) );
  XNOR U19672 ( .A(n20288), .B(n20275), .Z(n20277) );
  XOR U19673 ( .A(n20289), .B(n20290), .Z(n20275) );
  AND U19674 ( .A(n425), .B(n20291), .Z(n20290) );
  IV U19675 ( .A(n20286), .Z(n20288) );
  XOR U19676 ( .A(n20292), .B(n20293), .Z(n20286) );
  AND U19677 ( .A(n409), .B(n20285), .Z(n20293) );
  XNOR U19678 ( .A(n20283), .B(n20292), .Z(n20285) );
  XNOR U19679 ( .A(n20294), .B(n20295), .Z(n20283) );
  AND U19680 ( .A(n413), .B(n20296), .Z(n20295) );
  XOR U19681 ( .A(p_input[301]), .B(n20294), .Z(n20296) );
  XNOR U19682 ( .A(n20297), .B(n20298), .Z(n20294) );
  AND U19683 ( .A(n417), .B(n20299), .Z(n20298) );
  XOR U19684 ( .A(n20300), .B(n20301), .Z(n20292) );
  AND U19685 ( .A(n421), .B(n20291), .Z(n20301) );
  XNOR U19686 ( .A(n20302), .B(n20289), .Z(n20291) );
  XOR U19687 ( .A(n20303), .B(n20304), .Z(n20289) );
  AND U19688 ( .A(n444), .B(n20305), .Z(n20304) );
  IV U19689 ( .A(n20300), .Z(n20302) );
  XOR U19690 ( .A(n20306), .B(n20307), .Z(n20300) );
  AND U19691 ( .A(n428), .B(n20299), .Z(n20307) );
  XNOR U19692 ( .A(n20297), .B(n20306), .Z(n20299) );
  XNOR U19693 ( .A(n20308), .B(n20309), .Z(n20297) );
  AND U19694 ( .A(n432), .B(n20310), .Z(n20309) );
  XOR U19695 ( .A(p_input[317]), .B(n20308), .Z(n20310) );
  XNOR U19696 ( .A(n20311), .B(n20312), .Z(n20308) );
  AND U19697 ( .A(n436), .B(n20313), .Z(n20312) );
  XOR U19698 ( .A(n20314), .B(n20315), .Z(n20306) );
  AND U19699 ( .A(n440), .B(n20305), .Z(n20315) );
  XNOR U19700 ( .A(n20316), .B(n20303), .Z(n20305) );
  XOR U19701 ( .A(n20317), .B(n20318), .Z(n20303) );
  AND U19702 ( .A(n463), .B(n20319), .Z(n20318) );
  IV U19703 ( .A(n20314), .Z(n20316) );
  XOR U19704 ( .A(n20320), .B(n20321), .Z(n20314) );
  AND U19705 ( .A(n447), .B(n20313), .Z(n20321) );
  XNOR U19706 ( .A(n20311), .B(n20320), .Z(n20313) );
  XNOR U19707 ( .A(n20322), .B(n20323), .Z(n20311) );
  AND U19708 ( .A(n451), .B(n20324), .Z(n20323) );
  XOR U19709 ( .A(p_input[333]), .B(n20322), .Z(n20324) );
  XNOR U19710 ( .A(n20325), .B(n20326), .Z(n20322) );
  AND U19711 ( .A(n455), .B(n20327), .Z(n20326) );
  XOR U19712 ( .A(n20328), .B(n20329), .Z(n20320) );
  AND U19713 ( .A(n459), .B(n20319), .Z(n20329) );
  XNOR U19714 ( .A(n20330), .B(n20317), .Z(n20319) );
  XOR U19715 ( .A(n20331), .B(n20332), .Z(n20317) );
  AND U19716 ( .A(n482), .B(n20333), .Z(n20332) );
  IV U19717 ( .A(n20328), .Z(n20330) );
  XOR U19718 ( .A(n20334), .B(n20335), .Z(n20328) );
  AND U19719 ( .A(n466), .B(n20327), .Z(n20335) );
  XNOR U19720 ( .A(n20325), .B(n20334), .Z(n20327) );
  XNOR U19721 ( .A(n20336), .B(n20337), .Z(n20325) );
  AND U19722 ( .A(n470), .B(n20338), .Z(n20337) );
  XOR U19723 ( .A(p_input[349]), .B(n20336), .Z(n20338) );
  XNOR U19724 ( .A(n20339), .B(n20340), .Z(n20336) );
  AND U19725 ( .A(n474), .B(n20341), .Z(n20340) );
  XOR U19726 ( .A(n20342), .B(n20343), .Z(n20334) );
  AND U19727 ( .A(n478), .B(n20333), .Z(n20343) );
  XNOR U19728 ( .A(n20344), .B(n20331), .Z(n20333) );
  XOR U19729 ( .A(n20345), .B(n20346), .Z(n20331) );
  AND U19730 ( .A(n501), .B(n20347), .Z(n20346) );
  IV U19731 ( .A(n20342), .Z(n20344) );
  XOR U19732 ( .A(n20348), .B(n20349), .Z(n20342) );
  AND U19733 ( .A(n485), .B(n20341), .Z(n20349) );
  XNOR U19734 ( .A(n20339), .B(n20348), .Z(n20341) );
  XNOR U19735 ( .A(n20350), .B(n20351), .Z(n20339) );
  AND U19736 ( .A(n489), .B(n20352), .Z(n20351) );
  XOR U19737 ( .A(p_input[365]), .B(n20350), .Z(n20352) );
  XNOR U19738 ( .A(n20353), .B(n20354), .Z(n20350) );
  AND U19739 ( .A(n493), .B(n20355), .Z(n20354) );
  XOR U19740 ( .A(n20356), .B(n20357), .Z(n20348) );
  AND U19741 ( .A(n497), .B(n20347), .Z(n20357) );
  XNOR U19742 ( .A(n20358), .B(n20345), .Z(n20347) );
  XOR U19743 ( .A(n20359), .B(n20360), .Z(n20345) );
  AND U19744 ( .A(n520), .B(n20361), .Z(n20360) );
  IV U19745 ( .A(n20356), .Z(n20358) );
  XOR U19746 ( .A(n20362), .B(n20363), .Z(n20356) );
  AND U19747 ( .A(n504), .B(n20355), .Z(n20363) );
  XNOR U19748 ( .A(n20353), .B(n20362), .Z(n20355) );
  XNOR U19749 ( .A(n20364), .B(n20365), .Z(n20353) );
  AND U19750 ( .A(n508), .B(n20366), .Z(n20365) );
  XOR U19751 ( .A(p_input[381]), .B(n20364), .Z(n20366) );
  XNOR U19752 ( .A(n20367), .B(n20368), .Z(n20364) );
  AND U19753 ( .A(n512), .B(n20369), .Z(n20368) );
  XOR U19754 ( .A(n20370), .B(n20371), .Z(n20362) );
  AND U19755 ( .A(n516), .B(n20361), .Z(n20371) );
  XNOR U19756 ( .A(n20372), .B(n20359), .Z(n20361) );
  XOR U19757 ( .A(n20373), .B(n20374), .Z(n20359) );
  AND U19758 ( .A(n539), .B(n20375), .Z(n20374) );
  IV U19759 ( .A(n20370), .Z(n20372) );
  XOR U19760 ( .A(n20376), .B(n20377), .Z(n20370) );
  AND U19761 ( .A(n523), .B(n20369), .Z(n20377) );
  XNOR U19762 ( .A(n20367), .B(n20376), .Z(n20369) );
  XNOR U19763 ( .A(n20378), .B(n20379), .Z(n20367) );
  AND U19764 ( .A(n527), .B(n20380), .Z(n20379) );
  XOR U19765 ( .A(p_input[397]), .B(n20378), .Z(n20380) );
  XNOR U19766 ( .A(n20381), .B(n20382), .Z(n20378) );
  AND U19767 ( .A(n531), .B(n20383), .Z(n20382) );
  XOR U19768 ( .A(n20384), .B(n20385), .Z(n20376) );
  AND U19769 ( .A(n535), .B(n20375), .Z(n20385) );
  XNOR U19770 ( .A(n20386), .B(n20373), .Z(n20375) );
  XOR U19771 ( .A(n20387), .B(n20388), .Z(n20373) );
  AND U19772 ( .A(n558), .B(n20389), .Z(n20388) );
  IV U19773 ( .A(n20384), .Z(n20386) );
  XOR U19774 ( .A(n20390), .B(n20391), .Z(n20384) );
  AND U19775 ( .A(n542), .B(n20383), .Z(n20391) );
  XNOR U19776 ( .A(n20381), .B(n20390), .Z(n20383) );
  XNOR U19777 ( .A(n20392), .B(n20393), .Z(n20381) );
  AND U19778 ( .A(n546), .B(n20394), .Z(n20393) );
  XOR U19779 ( .A(p_input[413]), .B(n20392), .Z(n20394) );
  XNOR U19780 ( .A(n20395), .B(n20396), .Z(n20392) );
  AND U19781 ( .A(n550), .B(n20397), .Z(n20396) );
  XOR U19782 ( .A(n20398), .B(n20399), .Z(n20390) );
  AND U19783 ( .A(n554), .B(n20389), .Z(n20399) );
  XNOR U19784 ( .A(n20400), .B(n20387), .Z(n20389) );
  XOR U19785 ( .A(n20401), .B(n20402), .Z(n20387) );
  AND U19786 ( .A(n577), .B(n20403), .Z(n20402) );
  IV U19787 ( .A(n20398), .Z(n20400) );
  XOR U19788 ( .A(n20404), .B(n20405), .Z(n20398) );
  AND U19789 ( .A(n561), .B(n20397), .Z(n20405) );
  XNOR U19790 ( .A(n20395), .B(n20404), .Z(n20397) );
  XNOR U19791 ( .A(n20406), .B(n20407), .Z(n20395) );
  AND U19792 ( .A(n565), .B(n20408), .Z(n20407) );
  XOR U19793 ( .A(p_input[429]), .B(n20406), .Z(n20408) );
  XNOR U19794 ( .A(n20409), .B(n20410), .Z(n20406) );
  AND U19795 ( .A(n569), .B(n20411), .Z(n20410) );
  XOR U19796 ( .A(n20412), .B(n20413), .Z(n20404) );
  AND U19797 ( .A(n573), .B(n20403), .Z(n20413) );
  XNOR U19798 ( .A(n20414), .B(n20401), .Z(n20403) );
  XOR U19799 ( .A(n20415), .B(n20416), .Z(n20401) );
  AND U19800 ( .A(n596), .B(n20417), .Z(n20416) );
  IV U19801 ( .A(n20412), .Z(n20414) );
  XOR U19802 ( .A(n20418), .B(n20419), .Z(n20412) );
  AND U19803 ( .A(n580), .B(n20411), .Z(n20419) );
  XNOR U19804 ( .A(n20409), .B(n20418), .Z(n20411) );
  XNOR U19805 ( .A(n20420), .B(n20421), .Z(n20409) );
  AND U19806 ( .A(n584), .B(n20422), .Z(n20421) );
  XOR U19807 ( .A(p_input[445]), .B(n20420), .Z(n20422) );
  XNOR U19808 ( .A(n20423), .B(n20424), .Z(n20420) );
  AND U19809 ( .A(n588), .B(n20425), .Z(n20424) );
  XOR U19810 ( .A(n20426), .B(n20427), .Z(n20418) );
  AND U19811 ( .A(n592), .B(n20417), .Z(n20427) );
  XNOR U19812 ( .A(n20428), .B(n20415), .Z(n20417) );
  XOR U19813 ( .A(n20429), .B(n20430), .Z(n20415) );
  AND U19814 ( .A(n615), .B(n20431), .Z(n20430) );
  IV U19815 ( .A(n20426), .Z(n20428) );
  XOR U19816 ( .A(n20432), .B(n20433), .Z(n20426) );
  AND U19817 ( .A(n599), .B(n20425), .Z(n20433) );
  XNOR U19818 ( .A(n20423), .B(n20432), .Z(n20425) );
  XNOR U19819 ( .A(n20434), .B(n20435), .Z(n20423) );
  AND U19820 ( .A(n603), .B(n20436), .Z(n20435) );
  XOR U19821 ( .A(p_input[461]), .B(n20434), .Z(n20436) );
  XNOR U19822 ( .A(n20437), .B(n20438), .Z(n20434) );
  AND U19823 ( .A(n607), .B(n20439), .Z(n20438) );
  XOR U19824 ( .A(n20440), .B(n20441), .Z(n20432) );
  AND U19825 ( .A(n611), .B(n20431), .Z(n20441) );
  XNOR U19826 ( .A(n20442), .B(n20429), .Z(n20431) );
  XOR U19827 ( .A(n20443), .B(n20444), .Z(n20429) );
  AND U19828 ( .A(n634), .B(n20445), .Z(n20444) );
  IV U19829 ( .A(n20440), .Z(n20442) );
  XOR U19830 ( .A(n20446), .B(n20447), .Z(n20440) );
  AND U19831 ( .A(n618), .B(n20439), .Z(n20447) );
  XNOR U19832 ( .A(n20437), .B(n20446), .Z(n20439) );
  XNOR U19833 ( .A(n20448), .B(n20449), .Z(n20437) );
  AND U19834 ( .A(n622), .B(n20450), .Z(n20449) );
  XOR U19835 ( .A(p_input[477]), .B(n20448), .Z(n20450) );
  XNOR U19836 ( .A(n20451), .B(n20452), .Z(n20448) );
  AND U19837 ( .A(n626), .B(n20453), .Z(n20452) );
  XOR U19838 ( .A(n20454), .B(n20455), .Z(n20446) );
  AND U19839 ( .A(n630), .B(n20445), .Z(n20455) );
  XNOR U19840 ( .A(n20456), .B(n20443), .Z(n20445) );
  XOR U19841 ( .A(n20457), .B(n20458), .Z(n20443) );
  AND U19842 ( .A(n653), .B(n20459), .Z(n20458) );
  IV U19843 ( .A(n20454), .Z(n20456) );
  XOR U19844 ( .A(n20460), .B(n20461), .Z(n20454) );
  AND U19845 ( .A(n637), .B(n20453), .Z(n20461) );
  XNOR U19846 ( .A(n20451), .B(n20460), .Z(n20453) );
  XNOR U19847 ( .A(n20462), .B(n20463), .Z(n20451) );
  AND U19848 ( .A(n641), .B(n20464), .Z(n20463) );
  XOR U19849 ( .A(p_input[493]), .B(n20462), .Z(n20464) );
  XNOR U19850 ( .A(n20465), .B(n20466), .Z(n20462) );
  AND U19851 ( .A(n645), .B(n20467), .Z(n20466) );
  XOR U19852 ( .A(n20468), .B(n20469), .Z(n20460) );
  AND U19853 ( .A(n649), .B(n20459), .Z(n20469) );
  XNOR U19854 ( .A(n20470), .B(n20457), .Z(n20459) );
  XOR U19855 ( .A(n20471), .B(n20472), .Z(n20457) );
  AND U19856 ( .A(n672), .B(n20473), .Z(n20472) );
  IV U19857 ( .A(n20468), .Z(n20470) );
  XOR U19858 ( .A(n20474), .B(n20475), .Z(n20468) );
  AND U19859 ( .A(n656), .B(n20467), .Z(n20475) );
  XNOR U19860 ( .A(n20465), .B(n20474), .Z(n20467) );
  XNOR U19861 ( .A(n20476), .B(n20477), .Z(n20465) );
  AND U19862 ( .A(n660), .B(n20478), .Z(n20477) );
  XOR U19863 ( .A(p_input[509]), .B(n20476), .Z(n20478) );
  XNOR U19864 ( .A(n20479), .B(n20480), .Z(n20476) );
  AND U19865 ( .A(n664), .B(n20481), .Z(n20480) );
  XOR U19866 ( .A(n20482), .B(n20483), .Z(n20474) );
  AND U19867 ( .A(n668), .B(n20473), .Z(n20483) );
  XNOR U19868 ( .A(n20484), .B(n20471), .Z(n20473) );
  XOR U19869 ( .A(n20485), .B(n20486), .Z(n20471) );
  AND U19870 ( .A(n691), .B(n20487), .Z(n20486) );
  IV U19871 ( .A(n20482), .Z(n20484) );
  XOR U19872 ( .A(n20488), .B(n20489), .Z(n20482) );
  AND U19873 ( .A(n675), .B(n20481), .Z(n20489) );
  XNOR U19874 ( .A(n20479), .B(n20488), .Z(n20481) );
  XNOR U19875 ( .A(n20490), .B(n20491), .Z(n20479) );
  AND U19876 ( .A(n679), .B(n20492), .Z(n20491) );
  XOR U19877 ( .A(p_input[525]), .B(n20490), .Z(n20492) );
  XNOR U19878 ( .A(n20493), .B(n20494), .Z(n20490) );
  AND U19879 ( .A(n683), .B(n20495), .Z(n20494) );
  XOR U19880 ( .A(n20496), .B(n20497), .Z(n20488) );
  AND U19881 ( .A(n687), .B(n20487), .Z(n20497) );
  XNOR U19882 ( .A(n20498), .B(n20485), .Z(n20487) );
  XOR U19883 ( .A(n20499), .B(n20500), .Z(n20485) );
  AND U19884 ( .A(n710), .B(n20501), .Z(n20500) );
  IV U19885 ( .A(n20496), .Z(n20498) );
  XOR U19886 ( .A(n20502), .B(n20503), .Z(n20496) );
  AND U19887 ( .A(n694), .B(n20495), .Z(n20503) );
  XNOR U19888 ( .A(n20493), .B(n20502), .Z(n20495) );
  XNOR U19889 ( .A(n20504), .B(n20505), .Z(n20493) );
  AND U19890 ( .A(n698), .B(n20506), .Z(n20505) );
  XOR U19891 ( .A(p_input[541]), .B(n20504), .Z(n20506) );
  XNOR U19892 ( .A(n20507), .B(n20508), .Z(n20504) );
  AND U19893 ( .A(n702), .B(n20509), .Z(n20508) );
  XOR U19894 ( .A(n20510), .B(n20511), .Z(n20502) );
  AND U19895 ( .A(n706), .B(n20501), .Z(n20511) );
  XNOR U19896 ( .A(n20512), .B(n20499), .Z(n20501) );
  XOR U19897 ( .A(n20513), .B(n20514), .Z(n20499) );
  AND U19898 ( .A(n729), .B(n20515), .Z(n20514) );
  IV U19899 ( .A(n20510), .Z(n20512) );
  XOR U19900 ( .A(n20516), .B(n20517), .Z(n20510) );
  AND U19901 ( .A(n713), .B(n20509), .Z(n20517) );
  XNOR U19902 ( .A(n20507), .B(n20516), .Z(n20509) );
  XNOR U19903 ( .A(n20518), .B(n20519), .Z(n20507) );
  AND U19904 ( .A(n717), .B(n20520), .Z(n20519) );
  XOR U19905 ( .A(p_input[557]), .B(n20518), .Z(n20520) );
  XNOR U19906 ( .A(n20521), .B(n20522), .Z(n20518) );
  AND U19907 ( .A(n721), .B(n20523), .Z(n20522) );
  XOR U19908 ( .A(n20524), .B(n20525), .Z(n20516) );
  AND U19909 ( .A(n725), .B(n20515), .Z(n20525) );
  XNOR U19910 ( .A(n20526), .B(n20513), .Z(n20515) );
  XOR U19911 ( .A(n20527), .B(n20528), .Z(n20513) );
  AND U19912 ( .A(n748), .B(n20529), .Z(n20528) );
  IV U19913 ( .A(n20524), .Z(n20526) );
  XOR U19914 ( .A(n20530), .B(n20531), .Z(n20524) );
  AND U19915 ( .A(n732), .B(n20523), .Z(n20531) );
  XNOR U19916 ( .A(n20521), .B(n20530), .Z(n20523) );
  XNOR U19917 ( .A(n20532), .B(n20533), .Z(n20521) );
  AND U19918 ( .A(n736), .B(n20534), .Z(n20533) );
  XOR U19919 ( .A(p_input[573]), .B(n20532), .Z(n20534) );
  XNOR U19920 ( .A(n20535), .B(n20536), .Z(n20532) );
  AND U19921 ( .A(n740), .B(n20537), .Z(n20536) );
  XOR U19922 ( .A(n20538), .B(n20539), .Z(n20530) );
  AND U19923 ( .A(n744), .B(n20529), .Z(n20539) );
  XNOR U19924 ( .A(n20540), .B(n20527), .Z(n20529) );
  XOR U19925 ( .A(n20541), .B(n20542), .Z(n20527) );
  AND U19926 ( .A(n767), .B(n20543), .Z(n20542) );
  IV U19927 ( .A(n20538), .Z(n20540) );
  XOR U19928 ( .A(n20544), .B(n20545), .Z(n20538) );
  AND U19929 ( .A(n751), .B(n20537), .Z(n20545) );
  XNOR U19930 ( .A(n20535), .B(n20544), .Z(n20537) );
  XNOR U19931 ( .A(n20546), .B(n20547), .Z(n20535) );
  AND U19932 ( .A(n755), .B(n20548), .Z(n20547) );
  XOR U19933 ( .A(p_input[589]), .B(n20546), .Z(n20548) );
  XNOR U19934 ( .A(n20549), .B(n20550), .Z(n20546) );
  AND U19935 ( .A(n759), .B(n20551), .Z(n20550) );
  XOR U19936 ( .A(n20552), .B(n20553), .Z(n20544) );
  AND U19937 ( .A(n763), .B(n20543), .Z(n20553) );
  XNOR U19938 ( .A(n20554), .B(n20541), .Z(n20543) );
  XOR U19939 ( .A(n20555), .B(n20556), .Z(n20541) );
  AND U19940 ( .A(n786), .B(n20557), .Z(n20556) );
  IV U19941 ( .A(n20552), .Z(n20554) );
  XOR U19942 ( .A(n20558), .B(n20559), .Z(n20552) );
  AND U19943 ( .A(n770), .B(n20551), .Z(n20559) );
  XNOR U19944 ( .A(n20549), .B(n20558), .Z(n20551) );
  XNOR U19945 ( .A(n20560), .B(n20561), .Z(n20549) );
  AND U19946 ( .A(n774), .B(n20562), .Z(n20561) );
  XOR U19947 ( .A(p_input[605]), .B(n20560), .Z(n20562) );
  XNOR U19948 ( .A(n20563), .B(n20564), .Z(n20560) );
  AND U19949 ( .A(n778), .B(n20565), .Z(n20564) );
  XOR U19950 ( .A(n20566), .B(n20567), .Z(n20558) );
  AND U19951 ( .A(n782), .B(n20557), .Z(n20567) );
  XNOR U19952 ( .A(n20568), .B(n20555), .Z(n20557) );
  XOR U19953 ( .A(n20569), .B(n20570), .Z(n20555) );
  AND U19954 ( .A(n805), .B(n20571), .Z(n20570) );
  IV U19955 ( .A(n20566), .Z(n20568) );
  XOR U19956 ( .A(n20572), .B(n20573), .Z(n20566) );
  AND U19957 ( .A(n789), .B(n20565), .Z(n20573) );
  XNOR U19958 ( .A(n20563), .B(n20572), .Z(n20565) );
  XNOR U19959 ( .A(n20574), .B(n20575), .Z(n20563) );
  AND U19960 ( .A(n793), .B(n20576), .Z(n20575) );
  XOR U19961 ( .A(p_input[621]), .B(n20574), .Z(n20576) );
  XNOR U19962 ( .A(n20577), .B(n20578), .Z(n20574) );
  AND U19963 ( .A(n797), .B(n20579), .Z(n20578) );
  XOR U19964 ( .A(n20580), .B(n20581), .Z(n20572) );
  AND U19965 ( .A(n801), .B(n20571), .Z(n20581) );
  XNOR U19966 ( .A(n20582), .B(n20569), .Z(n20571) );
  XOR U19967 ( .A(n20583), .B(n20584), .Z(n20569) );
  AND U19968 ( .A(n824), .B(n20585), .Z(n20584) );
  IV U19969 ( .A(n20580), .Z(n20582) );
  XOR U19970 ( .A(n20586), .B(n20587), .Z(n20580) );
  AND U19971 ( .A(n808), .B(n20579), .Z(n20587) );
  XNOR U19972 ( .A(n20577), .B(n20586), .Z(n20579) );
  XNOR U19973 ( .A(n20588), .B(n20589), .Z(n20577) );
  AND U19974 ( .A(n812), .B(n20590), .Z(n20589) );
  XOR U19975 ( .A(p_input[637]), .B(n20588), .Z(n20590) );
  XNOR U19976 ( .A(n20591), .B(n20592), .Z(n20588) );
  AND U19977 ( .A(n816), .B(n20593), .Z(n20592) );
  XOR U19978 ( .A(n20594), .B(n20595), .Z(n20586) );
  AND U19979 ( .A(n820), .B(n20585), .Z(n20595) );
  XNOR U19980 ( .A(n20596), .B(n20583), .Z(n20585) );
  XOR U19981 ( .A(n20597), .B(n20598), .Z(n20583) );
  AND U19982 ( .A(n843), .B(n20599), .Z(n20598) );
  IV U19983 ( .A(n20594), .Z(n20596) );
  XOR U19984 ( .A(n20600), .B(n20601), .Z(n20594) );
  AND U19985 ( .A(n827), .B(n20593), .Z(n20601) );
  XNOR U19986 ( .A(n20591), .B(n20600), .Z(n20593) );
  XNOR U19987 ( .A(n20602), .B(n20603), .Z(n20591) );
  AND U19988 ( .A(n831), .B(n20604), .Z(n20603) );
  XOR U19989 ( .A(p_input[653]), .B(n20602), .Z(n20604) );
  XNOR U19990 ( .A(n20605), .B(n20606), .Z(n20602) );
  AND U19991 ( .A(n835), .B(n20607), .Z(n20606) );
  XOR U19992 ( .A(n20608), .B(n20609), .Z(n20600) );
  AND U19993 ( .A(n839), .B(n20599), .Z(n20609) );
  XNOR U19994 ( .A(n20610), .B(n20597), .Z(n20599) );
  XOR U19995 ( .A(n20611), .B(n20612), .Z(n20597) );
  AND U19996 ( .A(n862), .B(n20613), .Z(n20612) );
  IV U19997 ( .A(n20608), .Z(n20610) );
  XOR U19998 ( .A(n20614), .B(n20615), .Z(n20608) );
  AND U19999 ( .A(n846), .B(n20607), .Z(n20615) );
  XNOR U20000 ( .A(n20605), .B(n20614), .Z(n20607) );
  XNOR U20001 ( .A(n20616), .B(n20617), .Z(n20605) );
  AND U20002 ( .A(n850), .B(n20618), .Z(n20617) );
  XOR U20003 ( .A(p_input[669]), .B(n20616), .Z(n20618) );
  XNOR U20004 ( .A(n20619), .B(n20620), .Z(n20616) );
  AND U20005 ( .A(n854), .B(n20621), .Z(n20620) );
  XOR U20006 ( .A(n20622), .B(n20623), .Z(n20614) );
  AND U20007 ( .A(n858), .B(n20613), .Z(n20623) );
  XNOR U20008 ( .A(n20624), .B(n20611), .Z(n20613) );
  XOR U20009 ( .A(n20625), .B(n20626), .Z(n20611) );
  AND U20010 ( .A(n881), .B(n20627), .Z(n20626) );
  IV U20011 ( .A(n20622), .Z(n20624) );
  XOR U20012 ( .A(n20628), .B(n20629), .Z(n20622) );
  AND U20013 ( .A(n865), .B(n20621), .Z(n20629) );
  XNOR U20014 ( .A(n20619), .B(n20628), .Z(n20621) );
  XNOR U20015 ( .A(n20630), .B(n20631), .Z(n20619) );
  AND U20016 ( .A(n869), .B(n20632), .Z(n20631) );
  XOR U20017 ( .A(p_input[685]), .B(n20630), .Z(n20632) );
  XNOR U20018 ( .A(n20633), .B(n20634), .Z(n20630) );
  AND U20019 ( .A(n873), .B(n20635), .Z(n20634) );
  XOR U20020 ( .A(n20636), .B(n20637), .Z(n20628) );
  AND U20021 ( .A(n877), .B(n20627), .Z(n20637) );
  XNOR U20022 ( .A(n20638), .B(n20625), .Z(n20627) );
  XOR U20023 ( .A(n20639), .B(n20640), .Z(n20625) );
  AND U20024 ( .A(n900), .B(n20641), .Z(n20640) );
  IV U20025 ( .A(n20636), .Z(n20638) );
  XOR U20026 ( .A(n20642), .B(n20643), .Z(n20636) );
  AND U20027 ( .A(n884), .B(n20635), .Z(n20643) );
  XNOR U20028 ( .A(n20633), .B(n20642), .Z(n20635) );
  XNOR U20029 ( .A(n20644), .B(n20645), .Z(n20633) );
  AND U20030 ( .A(n888), .B(n20646), .Z(n20645) );
  XOR U20031 ( .A(p_input[701]), .B(n20644), .Z(n20646) );
  XNOR U20032 ( .A(n20647), .B(n20648), .Z(n20644) );
  AND U20033 ( .A(n892), .B(n20649), .Z(n20648) );
  XOR U20034 ( .A(n20650), .B(n20651), .Z(n20642) );
  AND U20035 ( .A(n896), .B(n20641), .Z(n20651) );
  XNOR U20036 ( .A(n20652), .B(n20639), .Z(n20641) );
  XOR U20037 ( .A(n20653), .B(n20654), .Z(n20639) );
  AND U20038 ( .A(n919), .B(n20655), .Z(n20654) );
  IV U20039 ( .A(n20650), .Z(n20652) );
  XOR U20040 ( .A(n20656), .B(n20657), .Z(n20650) );
  AND U20041 ( .A(n903), .B(n20649), .Z(n20657) );
  XNOR U20042 ( .A(n20647), .B(n20656), .Z(n20649) );
  XNOR U20043 ( .A(n20658), .B(n20659), .Z(n20647) );
  AND U20044 ( .A(n907), .B(n20660), .Z(n20659) );
  XOR U20045 ( .A(p_input[717]), .B(n20658), .Z(n20660) );
  XNOR U20046 ( .A(n20661), .B(n20662), .Z(n20658) );
  AND U20047 ( .A(n911), .B(n20663), .Z(n20662) );
  XOR U20048 ( .A(n20664), .B(n20665), .Z(n20656) );
  AND U20049 ( .A(n915), .B(n20655), .Z(n20665) );
  XNOR U20050 ( .A(n20666), .B(n20653), .Z(n20655) );
  XOR U20051 ( .A(n20667), .B(n20668), .Z(n20653) );
  AND U20052 ( .A(n938), .B(n20669), .Z(n20668) );
  IV U20053 ( .A(n20664), .Z(n20666) );
  XOR U20054 ( .A(n20670), .B(n20671), .Z(n20664) );
  AND U20055 ( .A(n922), .B(n20663), .Z(n20671) );
  XNOR U20056 ( .A(n20661), .B(n20670), .Z(n20663) );
  XNOR U20057 ( .A(n20672), .B(n20673), .Z(n20661) );
  AND U20058 ( .A(n926), .B(n20674), .Z(n20673) );
  XOR U20059 ( .A(p_input[733]), .B(n20672), .Z(n20674) );
  XNOR U20060 ( .A(n20675), .B(n20676), .Z(n20672) );
  AND U20061 ( .A(n930), .B(n20677), .Z(n20676) );
  XOR U20062 ( .A(n20678), .B(n20679), .Z(n20670) );
  AND U20063 ( .A(n934), .B(n20669), .Z(n20679) );
  XNOR U20064 ( .A(n20680), .B(n20667), .Z(n20669) );
  XOR U20065 ( .A(n20681), .B(n20682), .Z(n20667) );
  AND U20066 ( .A(n957), .B(n20683), .Z(n20682) );
  IV U20067 ( .A(n20678), .Z(n20680) );
  XOR U20068 ( .A(n20684), .B(n20685), .Z(n20678) );
  AND U20069 ( .A(n941), .B(n20677), .Z(n20685) );
  XNOR U20070 ( .A(n20675), .B(n20684), .Z(n20677) );
  XNOR U20071 ( .A(n20686), .B(n20687), .Z(n20675) );
  AND U20072 ( .A(n945), .B(n20688), .Z(n20687) );
  XOR U20073 ( .A(p_input[749]), .B(n20686), .Z(n20688) );
  XNOR U20074 ( .A(n20689), .B(n20690), .Z(n20686) );
  AND U20075 ( .A(n949), .B(n20691), .Z(n20690) );
  XOR U20076 ( .A(n20692), .B(n20693), .Z(n20684) );
  AND U20077 ( .A(n953), .B(n20683), .Z(n20693) );
  XNOR U20078 ( .A(n20694), .B(n20681), .Z(n20683) );
  XOR U20079 ( .A(n20695), .B(n20696), .Z(n20681) );
  AND U20080 ( .A(n976), .B(n20697), .Z(n20696) );
  IV U20081 ( .A(n20692), .Z(n20694) );
  XOR U20082 ( .A(n20698), .B(n20699), .Z(n20692) );
  AND U20083 ( .A(n960), .B(n20691), .Z(n20699) );
  XNOR U20084 ( .A(n20689), .B(n20698), .Z(n20691) );
  XNOR U20085 ( .A(n20700), .B(n20701), .Z(n20689) );
  AND U20086 ( .A(n964), .B(n20702), .Z(n20701) );
  XOR U20087 ( .A(p_input[765]), .B(n20700), .Z(n20702) );
  XNOR U20088 ( .A(n20703), .B(n20704), .Z(n20700) );
  AND U20089 ( .A(n968), .B(n20705), .Z(n20704) );
  XOR U20090 ( .A(n20706), .B(n20707), .Z(n20698) );
  AND U20091 ( .A(n972), .B(n20697), .Z(n20707) );
  XNOR U20092 ( .A(n20708), .B(n20695), .Z(n20697) );
  XOR U20093 ( .A(n20709), .B(n20710), .Z(n20695) );
  AND U20094 ( .A(n995), .B(n20711), .Z(n20710) );
  IV U20095 ( .A(n20706), .Z(n20708) );
  XOR U20096 ( .A(n20712), .B(n20713), .Z(n20706) );
  AND U20097 ( .A(n979), .B(n20705), .Z(n20713) );
  XNOR U20098 ( .A(n20703), .B(n20712), .Z(n20705) );
  XNOR U20099 ( .A(n20714), .B(n20715), .Z(n20703) );
  AND U20100 ( .A(n983), .B(n20716), .Z(n20715) );
  XOR U20101 ( .A(p_input[781]), .B(n20714), .Z(n20716) );
  XNOR U20102 ( .A(n20717), .B(n20718), .Z(n20714) );
  AND U20103 ( .A(n987), .B(n20719), .Z(n20718) );
  XOR U20104 ( .A(n20720), .B(n20721), .Z(n20712) );
  AND U20105 ( .A(n991), .B(n20711), .Z(n20721) );
  XNOR U20106 ( .A(n20722), .B(n20709), .Z(n20711) );
  XOR U20107 ( .A(n20723), .B(n20724), .Z(n20709) );
  AND U20108 ( .A(n1014), .B(n20725), .Z(n20724) );
  IV U20109 ( .A(n20720), .Z(n20722) );
  XOR U20110 ( .A(n20726), .B(n20727), .Z(n20720) );
  AND U20111 ( .A(n998), .B(n20719), .Z(n20727) );
  XNOR U20112 ( .A(n20717), .B(n20726), .Z(n20719) );
  XNOR U20113 ( .A(n20728), .B(n20729), .Z(n20717) );
  AND U20114 ( .A(n1002), .B(n20730), .Z(n20729) );
  XOR U20115 ( .A(p_input[797]), .B(n20728), .Z(n20730) );
  XNOR U20116 ( .A(n20731), .B(n20732), .Z(n20728) );
  AND U20117 ( .A(n1006), .B(n20733), .Z(n20732) );
  XOR U20118 ( .A(n20734), .B(n20735), .Z(n20726) );
  AND U20119 ( .A(n1010), .B(n20725), .Z(n20735) );
  XNOR U20120 ( .A(n20736), .B(n20723), .Z(n20725) );
  XOR U20121 ( .A(n20737), .B(n20738), .Z(n20723) );
  AND U20122 ( .A(n1033), .B(n20739), .Z(n20738) );
  IV U20123 ( .A(n20734), .Z(n20736) );
  XOR U20124 ( .A(n20740), .B(n20741), .Z(n20734) );
  AND U20125 ( .A(n1017), .B(n20733), .Z(n20741) );
  XNOR U20126 ( .A(n20731), .B(n20740), .Z(n20733) );
  XNOR U20127 ( .A(n20742), .B(n20743), .Z(n20731) );
  AND U20128 ( .A(n1021), .B(n20744), .Z(n20743) );
  XOR U20129 ( .A(p_input[813]), .B(n20742), .Z(n20744) );
  XNOR U20130 ( .A(n20745), .B(n20746), .Z(n20742) );
  AND U20131 ( .A(n1025), .B(n20747), .Z(n20746) );
  XOR U20132 ( .A(n20748), .B(n20749), .Z(n20740) );
  AND U20133 ( .A(n1029), .B(n20739), .Z(n20749) );
  XNOR U20134 ( .A(n20750), .B(n20737), .Z(n20739) );
  XOR U20135 ( .A(n20751), .B(n20752), .Z(n20737) );
  AND U20136 ( .A(n1052), .B(n20753), .Z(n20752) );
  IV U20137 ( .A(n20748), .Z(n20750) );
  XOR U20138 ( .A(n20754), .B(n20755), .Z(n20748) );
  AND U20139 ( .A(n1036), .B(n20747), .Z(n20755) );
  XNOR U20140 ( .A(n20745), .B(n20754), .Z(n20747) );
  XNOR U20141 ( .A(n20756), .B(n20757), .Z(n20745) );
  AND U20142 ( .A(n1040), .B(n20758), .Z(n20757) );
  XOR U20143 ( .A(p_input[829]), .B(n20756), .Z(n20758) );
  XNOR U20144 ( .A(n20759), .B(n20760), .Z(n20756) );
  AND U20145 ( .A(n1044), .B(n20761), .Z(n20760) );
  XOR U20146 ( .A(n20762), .B(n20763), .Z(n20754) );
  AND U20147 ( .A(n1048), .B(n20753), .Z(n20763) );
  XNOR U20148 ( .A(n20764), .B(n20751), .Z(n20753) );
  XOR U20149 ( .A(n20765), .B(n20766), .Z(n20751) );
  AND U20150 ( .A(n1071), .B(n20767), .Z(n20766) );
  IV U20151 ( .A(n20762), .Z(n20764) );
  XOR U20152 ( .A(n20768), .B(n20769), .Z(n20762) );
  AND U20153 ( .A(n1055), .B(n20761), .Z(n20769) );
  XNOR U20154 ( .A(n20759), .B(n20768), .Z(n20761) );
  XNOR U20155 ( .A(n20770), .B(n20771), .Z(n20759) );
  AND U20156 ( .A(n1059), .B(n20772), .Z(n20771) );
  XOR U20157 ( .A(p_input[845]), .B(n20770), .Z(n20772) );
  XNOR U20158 ( .A(n20773), .B(n20774), .Z(n20770) );
  AND U20159 ( .A(n1063), .B(n20775), .Z(n20774) );
  XOR U20160 ( .A(n20776), .B(n20777), .Z(n20768) );
  AND U20161 ( .A(n1067), .B(n20767), .Z(n20777) );
  XNOR U20162 ( .A(n20778), .B(n20765), .Z(n20767) );
  XOR U20163 ( .A(n20779), .B(n20780), .Z(n20765) );
  AND U20164 ( .A(n1090), .B(n20781), .Z(n20780) );
  IV U20165 ( .A(n20776), .Z(n20778) );
  XOR U20166 ( .A(n20782), .B(n20783), .Z(n20776) );
  AND U20167 ( .A(n1074), .B(n20775), .Z(n20783) );
  XNOR U20168 ( .A(n20773), .B(n20782), .Z(n20775) );
  XNOR U20169 ( .A(n20784), .B(n20785), .Z(n20773) );
  AND U20170 ( .A(n1078), .B(n20786), .Z(n20785) );
  XOR U20171 ( .A(p_input[861]), .B(n20784), .Z(n20786) );
  XNOR U20172 ( .A(n20787), .B(n20788), .Z(n20784) );
  AND U20173 ( .A(n1082), .B(n20789), .Z(n20788) );
  XOR U20174 ( .A(n20790), .B(n20791), .Z(n20782) );
  AND U20175 ( .A(n1086), .B(n20781), .Z(n20791) );
  XNOR U20176 ( .A(n20792), .B(n20779), .Z(n20781) );
  XOR U20177 ( .A(n20793), .B(n20794), .Z(n20779) );
  AND U20178 ( .A(n1109), .B(n20795), .Z(n20794) );
  IV U20179 ( .A(n20790), .Z(n20792) );
  XOR U20180 ( .A(n20796), .B(n20797), .Z(n20790) );
  AND U20181 ( .A(n1093), .B(n20789), .Z(n20797) );
  XNOR U20182 ( .A(n20787), .B(n20796), .Z(n20789) );
  XNOR U20183 ( .A(n20798), .B(n20799), .Z(n20787) );
  AND U20184 ( .A(n1097), .B(n20800), .Z(n20799) );
  XOR U20185 ( .A(p_input[877]), .B(n20798), .Z(n20800) );
  XNOR U20186 ( .A(n20801), .B(n20802), .Z(n20798) );
  AND U20187 ( .A(n1101), .B(n20803), .Z(n20802) );
  XOR U20188 ( .A(n20804), .B(n20805), .Z(n20796) );
  AND U20189 ( .A(n1105), .B(n20795), .Z(n20805) );
  XNOR U20190 ( .A(n20806), .B(n20793), .Z(n20795) );
  XOR U20191 ( .A(n20807), .B(n20808), .Z(n20793) );
  AND U20192 ( .A(n1128), .B(n20809), .Z(n20808) );
  IV U20193 ( .A(n20804), .Z(n20806) );
  XOR U20194 ( .A(n20810), .B(n20811), .Z(n20804) );
  AND U20195 ( .A(n1112), .B(n20803), .Z(n20811) );
  XNOR U20196 ( .A(n20801), .B(n20810), .Z(n20803) );
  XNOR U20197 ( .A(n20812), .B(n20813), .Z(n20801) );
  AND U20198 ( .A(n1116), .B(n20814), .Z(n20813) );
  XOR U20199 ( .A(p_input[893]), .B(n20812), .Z(n20814) );
  XNOR U20200 ( .A(n20815), .B(n20816), .Z(n20812) );
  AND U20201 ( .A(n1120), .B(n20817), .Z(n20816) );
  XOR U20202 ( .A(n20818), .B(n20819), .Z(n20810) );
  AND U20203 ( .A(n1124), .B(n20809), .Z(n20819) );
  XNOR U20204 ( .A(n20820), .B(n20807), .Z(n20809) );
  XOR U20205 ( .A(n20821), .B(n20822), .Z(n20807) );
  AND U20206 ( .A(n1147), .B(n20823), .Z(n20822) );
  IV U20207 ( .A(n20818), .Z(n20820) );
  XOR U20208 ( .A(n20824), .B(n20825), .Z(n20818) );
  AND U20209 ( .A(n1131), .B(n20817), .Z(n20825) );
  XNOR U20210 ( .A(n20815), .B(n20824), .Z(n20817) );
  XNOR U20211 ( .A(n20826), .B(n20827), .Z(n20815) );
  AND U20212 ( .A(n1135), .B(n20828), .Z(n20827) );
  XOR U20213 ( .A(p_input[909]), .B(n20826), .Z(n20828) );
  XNOR U20214 ( .A(n20829), .B(n20830), .Z(n20826) );
  AND U20215 ( .A(n1139), .B(n20831), .Z(n20830) );
  XOR U20216 ( .A(n20832), .B(n20833), .Z(n20824) );
  AND U20217 ( .A(n1143), .B(n20823), .Z(n20833) );
  XNOR U20218 ( .A(n20834), .B(n20821), .Z(n20823) );
  XOR U20219 ( .A(n20835), .B(n20836), .Z(n20821) );
  AND U20220 ( .A(n1166), .B(n20837), .Z(n20836) );
  IV U20221 ( .A(n20832), .Z(n20834) );
  XOR U20222 ( .A(n20838), .B(n20839), .Z(n20832) );
  AND U20223 ( .A(n1150), .B(n20831), .Z(n20839) );
  XNOR U20224 ( .A(n20829), .B(n20838), .Z(n20831) );
  XNOR U20225 ( .A(n20840), .B(n20841), .Z(n20829) );
  AND U20226 ( .A(n1154), .B(n20842), .Z(n20841) );
  XOR U20227 ( .A(p_input[925]), .B(n20840), .Z(n20842) );
  XNOR U20228 ( .A(n20843), .B(n20844), .Z(n20840) );
  AND U20229 ( .A(n1158), .B(n20845), .Z(n20844) );
  XOR U20230 ( .A(n20846), .B(n20847), .Z(n20838) );
  AND U20231 ( .A(n1162), .B(n20837), .Z(n20847) );
  XNOR U20232 ( .A(n20848), .B(n20835), .Z(n20837) );
  XOR U20233 ( .A(n20849), .B(n20850), .Z(n20835) );
  AND U20234 ( .A(n1185), .B(n20851), .Z(n20850) );
  IV U20235 ( .A(n20846), .Z(n20848) );
  XOR U20236 ( .A(n20852), .B(n20853), .Z(n20846) );
  AND U20237 ( .A(n1169), .B(n20845), .Z(n20853) );
  XNOR U20238 ( .A(n20843), .B(n20852), .Z(n20845) );
  XNOR U20239 ( .A(n20854), .B(n20855), .Z(n20843) );
  AND U20240 ( .A(n1173), .B(n20856), .Z(n20855) );
  XOR U20241 ( .A(p_input[941]), .B(n20854), .Z(n20856) );
  XNOR U20242 ( .A(n20857), .B(n20858), .Z(n20854) );
  AND U20243 ( .A(n1177), .B(n20859), .Z(n20858) );
  XOR U20244 ( .A(n20860), .B(n20861), .Z(n20852) );
  AND U20245 ( .A(n1181), .B(n20851), .Z(n20861) );
  XNOR U20246 ( .A(n20862), .B(n20849), .Z(n20851) );
  XOR U20247 ( .A(n20863), .B(n20864), .Z(n20849) );
  AND U20248 ( .A(n1204), .B(n20865), .Z(n20864) );
  IV U20249 ( .A(n20860), .Z(n20862) );
  XOR U20250 ( .A(n20866), .B(n20867), .Z(n20860) );
  AND U20251 ( .A(n1188), .B(n20859), .Z(n20867) );
  XNOR U20252 ( .A(n20857), .B(n20866), .Z(n20859) );
  XNOR U20253 ( .A(n20868), .B(n20869), .Z(n20857) );
  AND U20254 ( .A(n1192), .B(n20870), .Z(n20869) );
  XOR U20255 ( .A(p_input[957]), .B(n20868), .Z(n20870) );
  XNOR U20256 ( .A(n20871), .B(n20872), .Z(n20868) );
  AND U20257 ( .A(n1196), .B(n20873), .Z(n20872) );
  XOR U20258 ( .A(n20874), .B(n20875), .Z(n20866) );
  AND U20259 ( .A(n1200), .B(n20865), .Z(n20875) );
  XNOR U20260 ( .A(n20876), .B(n20863), .Z(n20865) );
  XOR U20261 ( .A(n20877), .B(n20878), .Z(n20863) );
  AND U20262 ( .A(n1223), .B(n20879), .Z(n20878) );
  IV U20263 ( .A(n20874), .Z(n20876) );
  XOR U20264 ( .A(n20880), .B(n20881), .Z(n20874) );
  AND U20265 ( .A(n1207), .B(n20873), .Z(n20881) );
  XNOR U20266 ( .A(n20871), .B(n20880), .Z(n20873) );
  XNOR U20267 ( .A(n20882), .B(n20883), .Z(n20871) );
  AND U20268 ( .A(n1211), .B(n20884), .Z(n20883) );
  XOR U20269 ( .A(p_input[973]), .B(n20882), .Z(n20884) );
  XNOR U20270 ( .A(n20885), .B(n20886), .Z(n20882) );
  AND U20271 ( .A(n1215), .B(n20887), .Z(n20886) );
  XOR U20272 ( .A(n20888), .B(n20889), .Z(n20880) );
  AND U20273 ( .A(n1219), .B(n20879), .Z(n20889) );
  XNOR U20274 ( .A(n20890), .B(n20877), .Z(n20879) );
  XOR U20275 ( .A(n20891), .B(n20892), .Z(n20877) );
  AND U20276 ( .A(n1242), .B(n20893), .Z(n20892) );
  IV U20277 ( .A(n20888), .Z(n20890) );
  XOR U20278 ( .A(n20894), .B(n20895), .Z(n20888) );
  AND U20279 ( .A(n1226), .B(n20887), .Z(n20895) );
  XNOR U20280 ( .A(n20885), .B(n20894), .Z(n20887) );
  XNOR U20281 ( .A(n20896), .B(n20897), .Z(n20885) );
  AND U20282 ( .A(n1230), .B(n20898), .Z(n20897) );
  XOR U20283 ( .A(p_input[989]), .B(n20896), .Z(n20898) );
  XNOR U20284 ( .A(n20899), .B(n20900), .Z(n20896) );
  AND U20285 ( .A(n1234), .B(n20901), .Z(n20900) );
  XOR U20286 ( .A(n20902), .B(n20903), .Z(n20894) );
  AND U20287 ( .A(n1238), .B(n20893), .Z(n20903) );
  XNOR U20288 ( .A(n20904), .B(n20891), .Z(n20893) );
  XOR U20289 ( .A(n20905), .B(n20906), .Z(n20891) );
  AND U20290 ( .A(n1261), .B(n20907), .Z(n20906) );
  IV U20291 ( .A(n20902), .Z(n20904) );
  XOR U20292 ( .A(n20908), .B(n20909), .Z(n20902) );
  AND U20293 ( .A(n1245), .B(n20901), .Z(n20909) );
  XNOR U20294 ( .A(n20899), .B(n20908), .Z(n20901) );
  XNOR U20295 ( .A(n20910), .B(n20911), .Z(n20899) );
  AND U20296 ( .A(n1249), .B(n20912), .Z(n20911) );
  XOR U20297 ( .A(p_input[1005]), .B(n20910), .Z(n20912) );
  XNOR U20298 ( .A(n20913), .B(n20914), .Z(n20910) );
  AND U20299 ( .A(n1253), .B(n20915), .Z(n20914) );
  XOR U20300 ( .A(n20916), .B(n20917), .Z(n20908) );
  AND U20301 ( .A(n1257), .B(n20907), .Z(n20917) );
  XNOR U20302 ( .A(n20918), .B(n20905), .Z(n20907) );
  XOR U20303 ( .A(n20919), .B(n20920), .Z(n20905) );
  AND U20304 ( .A(n1280), .B(n20921), .Z(n20920) );
  IV U20305 ( .A(n20916), .Z(n20918) );
  XOR U20306 ( .A(n20922), .B(n20923), .Z(n20916) );
  AND U20307 ( .A(n1264), .B(n20915), .Z(n20923) );
  XNOR U20308 ( .A(n20913), .B(n20922), .Z(n20915) );
  XNOR U20309 ( .A(n20924), .B(n20925), .Z(n20913) );
  AND U20310 ( .A(n1268), .B(n20926), .Z(n20925) );
  XOR U20311 ( .A(p_input[1021]), .B(n20924), .Z(n20926) );
  XNOR U20312 ( .A(n20927), .B(n20928), .Z(n20924) );
  AND U20313 ( .A(n1272), .B(n20929), .Z(n20928) );
  XOR U20314 ( .A(n20930), .B(n20931), .Z(n20922) );
  AND U20315 ( .A(n1276), .B(n20921), .Z(n20931) );
  XNOR U20316 ( .A(n20932), .B(n20919), .Z(n20921) );
  XOR U20317 ( .A(n20933), .B(n20934), .Z(n20919) );
  AND U20318 ( .A(n1299), .B(n20935), .Z(n20934) );
  IV U20319 ( .A(n20930), .Z(n20932) );
  XOR U20320 ( .A(n20936), .B(n20937), .Z(n20930) );
  AND U20321 ( .A(n1283), .B(n20929), .Z(n20937) );
  XNOR U20322 ( .A(n20927), .B(n20936), .Z(n20929) );
  XNOR U20323 ( .A(n20938), .B(n20939), .Z(n20927) );
  AND U20324 ( .A(n1287), .B(n20940), .Z(n20939) );
  XOR U20325 ( .A(p_input[1037]), .B(n20938), .Z(n20940) );
  XNOR U20326 ( .A(n20941), .B(n20942), .Z(n20938) );
  AND U20327 ( .A(n1291), .B(n20943), .Z(n20942) );
  XOR U20328 ( .A(n20944), .B(n20945), .Z(n20936) );
  AND U20329 ( .A(n1295), .B(n20935), .Z(n20945) );
  XNOR U20330 ( .A(n20946), .B(n20933), .Z(n20935) );
  XOR U20331 ( .A(n20947), .B(n20948), .Z(n20933) );
  AND U20332 ( .A(n1318), .B(n20949), .Z(n20948) );
  IV U20333 ( .A(n20944), .Z(n20946) );
  XOR U20334 ( .A(n20950), .B(n20951), .Z(n20944) );
  AND U20335 ( .A(n1302), .B(n20943), .Z(n20951) );
  XNOR U20336 ( .A(n20941), .B(n20950), .Z(n20943) );
  XNOR U20337 ( .A(n20952), .B(n20953), .Z(n20941) );
  AND U20338 ( .A(n1306), .B(n20954), .Z(n20953) );
  XOR U20339 ( .A(p_input[1053]), .B(n20952), .Z(n20954) );
  XNOR U20340 ( .A(n20955), .B(n20956), .Z(n20952) );
  AND U20341 ( .A(n1310), .B(n20957), .Z(n20956) );
  XOR U20342 ( .A(n20958), .B(n20959), .Z(n20950) );
  AND U20343 ( .A(n1314), .B(n20949), .Z(n20959) );
  XNOR U20344 ( .A(n20960), .B(n20947), .Z(n20949) );
  XOR U20345 ( .A(n20961), .B(n20962), .Z(n20947) );
  AND U20346 ( .A(n1337), .B(n20963), .Z(n20962) );
  IV U20347 ( .A(n20958), .Z(n20960) );
  XOR U20348 ( .A(n20964), .B(n20965), .Z(n20958) );
  AND U20349 ( .A(n1321), .B(n20957), .Z(n20965) );
  XNOR U20350 ( .A(n20955), .B(n20964), .Z(n20957) );
  XNOR U20351 ( .A(n20966), .B(n20967), .Z(n20955) );
  AND U20352 ( .A(n1325), .B(n20968), .Z(n20967) );
  XOR U20353 ( .A(p_input[1069]), .B(n20966), .Z(n20968) );
  XNOR U20354 ( .A(n20969), .B(n20970), .Z(n20966) );
  AND U20355 ( .A(n1329), .B(n20971), .Z(n20970) );
  XOR U20356 ( .A(n20972), .B(n20973), .Z(n20964) );
  AND U20357 ( .A(n1333), .B(n20963), .Z(n20973) );
  XNOR U20358 ( .A(n20974), .B(n20961), .Z(n20963) );
  XOR U20359 ( .A(n20975), .B(n20976), .Z(n20961) );
  AND U20360 ( .A(n1356), .B(n20977), .Z(n20976) );
  IV U20361 ( .A(n20972), .Z(n20974) );
  XOR U20362 ( .A(n20978), .B(n20979), .Z(n20972) );
  AND U20363 ( .A(n1340), .B(n20971), .Z(n20979) );
  XNOR U20364 ( .A(n20969), .B(n20978), .Z(n20971) );
  XNOR U20365 ( .A(n20980), .B(n20981), .Z(n20969) );
  AND U20366 ( .A(n1344), .B(n20982), .Z(n20981) );
  XOR U20367 ( .A(p_input[1085]), .B(n20980), .Z(n20982) );
  XNOR U20368 ( .A(n20983), .B(n20984), .Z(n20980) );
  AND U20369 ( .A(n1348), .B(n20985), .Z(n20984) );
  XOR U20370 ( .A(n20986), .B(n20987), .Z(n20978) );
  AND U20371 ( .A(n1352), .B(n20977), .Z(n20987) );
  XNOR U20372 ( .A(n20988), .B(n20975), .Z(n20977) );
  XOR U20373 ( .A(n20989), .B(n20990), .Z(n20975) );
  AND U20374 ( .A(n1375), .B(n20991), .Z(n20990) );
  IV U20375 ( .A(n20986), .Z(n20988) );
  XOR U20376 ( .A(n20992), .B(n20993), .Z(n20986) );
  AND U20377 ( .A(n1359), .B(n20985), .Z(n20993) );
  XNOR U20378 ( .A(n20983), .B(n20992), .Z(n20985) );
  XNOR U20379 ( .A(n20994), .B(n20995), .Z(n20983) );
  AND U20380 ( .A(n1363), .B(n20996), .Z(n20995) );
  XOR U20381 ( .A(p_input[1101]), .B(n20994), .Z(n20996) );
  XNOR U20382 ( .A(n20997), .B(n20998), .Z(n20994) );
  AND U20383 ( .A(n1367), .B(n20999), .Z(n20998) );
  XOR U20384 ( .A(n21000), .B(n21001), .Z(n20992) );
  AND U20385 ( .A(n1371), .B(n20991), .Z(n21001) );
  XNOR U20386 ( .A(n21002), .B(n20989), .Z(n20991) );
  XOR U20387 ( .A(n21003), .B(n21004), .Z(n20989) );
  AND U20388 ( .A(n1394), .B(n21005), .Z(n21004) );
  IV U20389 ( .A(n21000), .Z(n21002) );
  XOR U20390 ( .A(n21006), .B(n21007), .Z(n21000) );
  AND U20391 ( .A(n1378), .B(n20999), .Z(n21007) );
  XNOR U20392 ( .A(n20997), .B(n21006), .Z(n20999) );
  XNOR U20393 ( .A(n21008), .B(n21009), .Z(n20997) );
  AND U20394 ( .A(n1382), .B(n21010), .Z(n21009) );
  XOR U20395 ( .A(p_input[1117]), .B(n21008), .Z(n21010) );
  XNOR U20396 ( .A(n21011), .B(n21012), .Z(n21008) );
  AND U20397 ( .A(n1386), .B(n21013), .Z(n21012) );
  XOR U20398 ( .A(n21014), .B(n21015), .Z(n21006) );
  AND U20399 ( .A(n1390), .B(n21005), .Z(n21015) );
  XNOR U20400 ( .A(n21016), .B(n21003), .Z(n21005) );
  XOR U20401 ( .A(n21017), .B(n21018), .Z(n21003) );
  AND U20402 ( .A(n1413), .B(n21019), .Z(n21018) );
  IV U20403 ( .A(n21014), .Z(n21016) );
  XOR U20404 ( .A(n21020), .B(n21021), .Z(n21014) );
  AND U20405 ( .A(n1397), .B(n21013), .Z(n21021) );
  XNOR U20406 ( .A(n21011), .B(n21020), .Z(n21013) );
  XNOR U20407 ( .A(n21022), .B(n21023), .Z(n21011) );
  AND U20408 ( .A(n1401), .B(n21024), .Z(n21023) );
  XOR U20409 ( .A(p_input[1133]), .B(n21022), .Z(n21024) );
  XNOR U20410 ( .A(n21025), .B(n21026), .Z(n21022) );
  AND U20411 ( .A(n1405), .B(n21027), .Z(n21026) );
  XOR U20412 ( .A(n21028), .B(n21029), .Z(n21020) );
  AND U20413 ( .A(n1409), .B(n21019), .Z(n21029) );
  XNOR U20414 ( .A(n21030), .B(n21017), .Z(n21019) );
  XOR U20415 ( .A(n21031), .B(n21032), .Z(n21017) );
  AND U20416 ( .A(n1432), .B(n21033), .Z(n21032) );
  IV U20417 ( .A(n21028), .Z(n21030) );
  XOR U20418 ( .A(n21034), .B(n21035), .Z(n21028) );
  AND U20419 ( .A(n1416), .B(n21027), .Z(n21035) );
  XNOR U20420 ( .A(n21025), .B(n21034), .Z(n21027) );
  XNOR U20421 ( .A(n21036), .B(n21037), .Z(n21025) );
  AND U20422 ( .A(n1420), .B(n21038), .Z(n21037) );
  XOR U20423 ( .A(p_input[1149]), .B(n21036), .Z(n21038) );
  XNOR U20424 ( .A(n21039), .B(n21040), .Z(n21036) );
  AND U20425 ( .A(n1424), .B(n21041), .Z(n21040) );
  XOR U20426 ( .A(n21042), .B(n21043), .Z(n21034) );
  AND U20427 ( .A(n1428), .B(n21033), .Z(n21043) );
  XNOR U20428 ( .A(n21044), .B(n21031), .Z(n21033) );
  XOR U20429 ( .A(n21045), .B(n21046), .Z(n21031) );
  AND U20430 ( .A(n1451), .B(n21047), .Z(n21046) );
  IV U20431 ( .A(n21042), .Z(n21044) );
  XOR U20432 ( .A(n21048), .B(n21049), .Z(n21042) );
  AND U20433 ( .A(n1435), .B(n21041), .Z(n21049) );
  XNOR U20434 ( .A(n21039), .B(n21048), .Z(n21041) );
  XNOR U20435 ( .A(n21050), .B(n21051), .Z(n21039) );
  AND U20436 ( .A(n1439), .B(n21052), .Z(n21051) );
  XOR U20437 ( .A(p_input[1165]), .B(n21050), .Z(n21052) );
  XNOR U20438 ( .A(n21053), .B(n21054), .Z(n21050) );
  AND U20439 ( .A(n1443), .B(n21055), .Z(n21054) );
  XOR U20440 ( .A(n21056), .B(n21057), .Z(n21048) );
  AND U20441 ( .A(n1447), .B(n21047), .Z(n21057) );
  XNOR U20442 ( .A(n21058), .B(n21045), .Z(n21047) );
  XOR U20443 ( .A(n21059), .B(n21060), .Z(n21045) );
  AND U20444 ( .A(n1470), .B(n21061), .Z(n21060) );
  IV U20445 ( .A(n21056), .Z(n21058) );
  XOR U20446 ( .A(n21062), .B(n21063), .Z(n21056) );
  AND U20447 ( .A(n1454), .B(n21055), .Z(n21063) );
  XNOR U20448 ( .A(n21053), .B(n21062), .Z(n21055) );
  XNOR U20449 ( .A(n21064), .B(n21065), .Z(n21053) );
  AND U20450 ( .A(n1458), .B(n21066), .Z(n21065) );
  XOR U20451 ( .A(p_input[1181]), .B(n21064), .Z(n21066) );
  XNOR U20452 ( .A(n21067), .B(n21068), .Z(n21064) );
  AND U20453 ( .A(n1462), .B(n21069), .Z(n21068) );
  XOR U20454 ( .A(n21070), .B(n21071), .Z(n21062) );
  AND U20455 ( .A(n1466), .B(n21061), .Z(n21071) );
  XNOR U20456 ( .A(n21072), .B(n21059), .Z(n21061) );
  XOR U20457 ( .A(n21073), .B(n21074), .Z(n21059) );
  AND U20458 ( .A(n1489), .B(n21075), .Z(n21074) );
  IV U20459 ( .A(n21070), .Z(n21072) );
  XOR U20460 ( .A(n21076), .B(n21077), .Z(n21070) );
  AND U20461 ( .A(n1473), .B(n21069), .Z(n21077) );
  XNOR U20462 ( .A(n21067), .B(n21076), .Z(n21069) );
  XNOR U20463 ( .A(n21078), .B(n21079), .Z(n21067) );
  AND U20464 ( .A(n1477), .B(n21080), .Z(n21079) );
  XOR U20465 ( .A(p_input[1197]), .B(n21078), .Z(n21080) );
  XNOR U20466 ( .A(n21081), .B(n21082), .Z(n21078) );
  AND U20467 ( .A(n1481), .B(n21083), .Z(n21082) );
  XOR U20468 ( .A(n21084), .B(n21085), .Z(n21076) );
  AND U20469 ( .A(n1485), .B(n21075), .Z(n21085) );
  XNOR U20470 ( .A(n21086), .B(n21073), .Z(n21075) );
  XOR U20471 ( .A(n21087), .B(n21088), .Z(n21073) );
  AND U20472 ( .A(n1508), .B(n21089), .Z(n21088) );
  IV U20473 ( .A(n21084), .Z(n21086) );
  XOR U20474 ( .A(n21090), .B(n21091), .Z(n21084) );
  AND U20475 ( .A(n1492), .B(n21083), .Z(n21091) );
  XNOR U20476 ( .A(n21081), .B(n21090), .Z(n21083) );
  XNOR U20477 ( .A(n21092), .B(n21093), .Z(n21081) );
  AND U20478 ( .A(n1496), .B(n21094), .Z(n21093) );
  XOR U20479 ( .A(p_input[1213]), .B(n21092), .Z(n21094) );
  XNOR U20480 ( .A(n21095), .B(n21096), .Z(n21092) );
  AND U20481 ( .A(n1500), .B(n21097), .Z(n21096) );
  XOR U20482 ( .A(n21098), .B(n21099), .Z(n21090) );
  AND U20483 ( .A(n1504), .B(n21089), .Z(n21099) );
  XNOR U20484 ( .A(n21100), .B(n21087), .Z(n21089) );
  XOR U20485 ( .A(n21101), .B(n21102), .Z(n21087) );
  AND U20486 ( .A(n1527), .B(n21103), .Z(n21102) );
  IV U20487 ( .A(n21098), .Z(n21100) );
  XOR U20488 ( .A(n21104), .B(n21105), .Z(n21098) );
  AND U20489 ( .A(n1511), .B(n21097), .Z(n21105) );
  XNOR U20490 ( .A(n21095), .B(n21104), .Z(n21097) );
  XNOR U20491 ( .A(n21106), .B(n21107), .Z(n21095) );
  AND U20492 ( .A(n1515), .B(n21108), .Z(n21107) );
  XOR U20493 ( .A(p_input[1229]), .B(n21106), .Z(n21108) );
  XNOR U20494 ( .A(n21109), .B(n21110), .Z(n21106) );
  AND U20495 ( .A(n1519), .B(n21111), .Z(n21110) );
  XOR U20496 ( .A(n21112), .B(n21113), .Z(n21104) );
  AND U20497 ( .A(n1523), .B(n21103), .Z(n21113) );
  XNOR U20498 ( .A(n21114), .B(n21101), .Z(n21103) );
  XOR U20499 ( .A(n21115), .B(n21116), .Z(n21101) );
  AND U20500 ( .A(n1546), .B(n21117), .Z(n21116) );
  IV U20501 ( .A(n21112), .Z(n21114) );
  XOR U20502 ( .A(n21118), .B(n21119), .Z(n21112) );
  AND U20503 ( .A(n1530), .B(n21111), .Z(n21119) );
  XNOR U20504 ( .A(n21109), .B(n21118), .Z(n21111) );
  XNOR U20505 ( .A(n21120), .B(n21121), .Z(n21109) );
  AND U20506 ( .A(n1534), .B(n21122), .Z(n21121) );
  XOR U20507 ( .A(p_input[1245]), .B(n21120), .Z(n21122) );
  XNOR U20508 ( .A(n21123), .B(n21124), .Z(n21120) );
  AND U20509 ( .A(n1538), .B(n21125), .Z(n21124) );
  XOR U20510 ( .A(n21126), .B(n21127), .Z(n21118) );
  AND U20511 ( .A(n1542), .B(n21117), .Z(n21127) );
  XNOR U20512 ( .A(n21128), .B(n21115), .Z(n21117) );
  XOR U20513 ( .A(n21129), .B(n21130), .Z(n21115) );
  AND U20514 ( .A(n1565), .B(n21131), .Z(n21130) );
  IV U20515 ( .A(n21126), .Z(n21128) );
  XOR U20516 ( .A(n21132), .B(n21133), .Z(n21126) );
  AND U20517 ( .A(n1549), .B(n21125), .Z(n21133) );
  XNOR U20518 ( .A(n21123), .B(n21132), .Z(n21125) );
  XNOR U20519 ( .A(n21134), .B(n21135), .Z(n21123) );
  AND U20520 ( .A(n1553), .B(n21136), .Z(n21135) );
  XOR U20521 ( .A(p_input[1261]), .B(n21134), .Z(n21136) );
  XNOR U20522 ( .A(n21137), .B(n21138), .Z(n21134) );
  AND U20523 ( .A(n1557), .B(n21139), .Z(n21138) );
  XOR U20524 ( .A(n21140), .B(n21141), .Z(n21132) );
  AND U20525 ( .A(n1561), .B(n21131), .Z(n21141) );
  XNOR U20526 ( .A(n21142), .B(n21129), .Z(n21131) );
  XOR U20527 ( .A(n21143), .B(n21144), .Z(n21129) );
  AND U20528 ( .A(n1584), .B(n21145), .Z(n21144) );
  IV U20529 ( .A(n21140), .Z(n21142) );
  XOR U20530 ( .A(n21146), .B(n21147), .Z(n21140) );
  AND U20531 ( .A(n1568), .B(n21139), .Z(n21147) );
  XNOR U20532 ( .A(n21137), .B(n21146), .Z(n21139) );
  XNOR U20533 ( .A(n21148), .B(n21149), .Z(n21137) );
  AND U20534 ( .A(n1572), .B(n21150), .Z(n21149) );
  XOR U20535 ( .A(p_input[1277]), .B(n21148), .Z(n21150) );
  XNOR U20536 ( .A(n21151), .B(n21152), .Z(n21148) );
  AND U20537 ( .A(n1576), .B(n21153), .Z(n21152) );
  XOR U20538 ( .A(n21154), .B(n21155), .Z(n21146) );
  AND U20539 ( .A(n1580), .B(n21145), .Z(n21155) );
  XNOR U20540 ( .A(n21156), .B(n21143), .Z(n21145) );
  XOR U20541 ( .A(n21157), .B(n21158), .Z(n21143) );
  AND U20542 ( .A(n1603), .B(n21159), .Z(n21158) );
  IV U20543 ( .A(n21154), .Z(n21156) );
  XOR U20544 ( .A(n21160), .B(n21161), .Z(n21154) );
  AND U20545 ( .A(n1587), .B(n21153), .Z(n21161) );
  XNOR U20546 ( .A(n21151), .B(n21160), .Z(n21153) );
  XNOR U20547 ( .A(n21162), .B(n21163), .Z(n21151) );
  AND U20548 ( .A(n1591), .B(n21164), .Z(n21163) );
  XOR U20549 ( .A(p_input[1293]), .B(n21162), .Z(n21164) );
  XNOR U20550 ( .A(n21165), .B(n21166), .Z(n21162) );
  AND U20551 ( .A(n1595), .B(n21167), .Z(n21166) );
  XOR U20552 ( .A(n21168), .B(n21169), .Z(n21160) );
  AND U20553 ( .A(n1599), .B(n21159), .Z(n21169) );
  XNOR U20554 ( .A(n21170), .B(n21157), .Z(n21159) );
  XOR U20555 ( .A(n21171), .B(n21172), .Z(n21157) );
  AND U20556 ( .A(n1622), .B(n21173), .Z(n21172) );
  IV U20557 ( .A(n21168), .Z(n21170) );
  XOR U20558 ( .A(n21174), .B(n21175), .Z(n21168) );
  AND U20559 ( .A(n1606), .B(n21167), .Z(n21175) );
  XNOR U20560 ( .A(n21165), .B(n21174), .Z(n21167) );
  XNOR U20561 ( .A(n21176), .B(n21177), .Z(n21165) );
  AND U20562 ( .A(n1610), .B(n21178), .Z(n21177) );
  XOR U20563 ( .A(p_input[1309]), .B(n21176), .Z(n21178) );
  XNOR U20564 ( .A(n21179), .B(n21180), .Z(n21176) );
  AND U20565 ( .A(n1614), .B(n21181), .Z(n21180) );
  XOR U20566 ( .A(n21182), .B(n21183), .Z(n21174) );
  AND U20567 ( .A(n1618), .B(n21173), .Z(n21183) );
  XNOR U20568 ( .A(n21184), .B(n21171), .Z(n21173) );
  XOR U20569 ( .A(n21185), .B(n21186), .Z(n21171) );
  AND U20570 ( .A(n1641), .B(n21187), .Z(n21186) );
  IV U20571 ( .A(n21182), .Z(n21184) );
  XOR U20572 ( .A(n21188), .B(n21189), .Z(n21182) );
  AND U20573 ( .A(n1625), .B(n21181), .Z(n21189) );
  XNOR U20574 ( .A(n21179), .B(n21188), .Z(n21181) );
  XNOR U20575 ( .A(n21190), .B(n21191), .Z(n21179) );
  AND U20576 ( .A(n1629), .B(n21192), .Z(n21191) );
  XOR U20577 ( .A(p_input[1325]), .B(n21190), .Z(n21192) );
  XNOR U20578 ( .A(n21193), .B(n21194), .Z(n21190) );
  AND U20579 ( .A(n1633), .B(n21195), .Z(n21194) );
  XOR U20580 ( .A(n21196), .B(n21197), .Z(n21188) );
  AND U20581 ( .A(n1637), .B(n21187), .Z(n21197) );
  XNOR U20582 ( .A(n21198), .B(n21185), .Z(n21187) );
  XOR U20583 ( .A(n21199), .B(n21200), .Z(n21185) );
  AND U20584 ( .A(n1660), .B(n21201), .Z(n21200) );
  IV U20585 ( .A(n21196), .Z(n21198) );
  XOR U20586 ( .A(n21202), .B(n21203), .Z(n21196) );
  AND U20587 ( .A(n1644), .B(n21195), .Z(n21203) );
  XNOR U20588 ( .A(n21193), .B(n21202), .Z(n21195) );
  XNOR U20589 ( .A(n21204), .B(n21205), .Z(n21193) );
  AND U20590 ( .A(n1648), .B(n21206), .Z(n21205) );
  XOR U20591 ( .A(p_input[1341]), .B(n21204), .Z(n21206) );
  XNOR U20592 ( .A(n21207), .B(n21208), .Z(n21204) );
  AND U20593 ( .A(n1652), .B(n21209), .Z(n21208) );
  XOR U20594 ( .A(n21210), .B(n21211), .Z(n21202) );
  AND U20595 ( .A(n1656), .B(n21201), .Z(n21211) );
  XNOR U20596 ( .A(n21212), .B(n21199), .Z(n21201) );
  XOR U20597 ( .A(n21213), .B(n21214), .Z(n21199) );
  AND U20598 ( .A(n1679), .B(n21215), .Z(n21214) );
  IV U20599 ( .A(n21210), .Z(n21212) );
  XOR U20600 ( .A(n21216), .B(n21217), .Z(n21210) );
  AND U20601 ( .A(n1663), .B(n21209), .Z(n21217) );
  XNOR U20602 ( .A(n21207), .B(n21216), .Z(n21209) );
  XNOR U20603 ( .A(n21218), .B(n21219), .Z(n21207) );
  AND U20604 ( .A(n1667), .B(n21220), .Z(n21219) );
  XOR U20605 ( .A(p_input[1357]), .B(n21218), .Z(n21220) );
  XNOR U20606 ( .A(n21221), .B(n21222), .Z(n21218) );
  AND U20607 ( .A(n1671), .B(n21223), .Z(n21222) );
  XOR U20608 ( .A(n21224), .B(n21225), .Z(n21216) );
  AND U20609 ( .A(n1675), .B(n21215), .Z(n21225) );
  XNOR U20610 ( .A(n21226), .B(n21213), .Z(n21215) );
  XOR U20611 ( .A(n21227), .B(n21228), .Z(n21213) );
  AND U20612 ( .A(n1698), .B(n21229), .Z(n21228) );
  IV U20613 ( .A(n21224), .Z(n21226) );
  XOR U20614 ( .A(n21230), .B(n21231), .Z(n21224) );
  AND U20615 ( .A(n1682), .B(n21223), .Z(n21231) );
  XNOR U20616 ( .A(n21221), .B(n21230), .Z(n21223) );
  XNOR U20617 ( .A(n21232), .B(n21233), .Z(n21221) );
  AND U20618 ( .A(n1686), .B(n21234), .Z(n21233) );
  XOR U20619 ( .A(p_input[1373]), .B(n21232), .Z(n21234) );
  XNOR U20620 ( .A(n21235), .B(n21236), .Z(n21232) );
  AND U20621 ( .A(n1690), .B(n21237), .Z(n21236) );
  XOR U20622 ( .A(n21238), .B(n21239), .Z(n21230) );
  AND U20623 ( .A(n1694), .B(n21229), .Z(n21239) );
  XNOR U20624 ( .A(n21240), .B(n21227), .Z(n21229) );
  XOR U20625 ( .A(n21241), .B(n21242), .Z(n21227) );
  AND U20626 ( .A(n1717), .B(n21243), .Z(n21242) );
  IV U20627 ( .A(n21238), .Z(n21240) );
  XOR U20628 ( .A(n21244), .B(n21245), .Z(n21238) );
  AND U20629 ( .A(n1701), .B(n21237), .Z(n21245) );
  XNOR U20630 ( .A(n21235), .B(n21244), .Z(n21237) );
  XNOR U20631 ( .A(n21246), .B(n21247), .Z(n21235) );
  AND U20632 ( .A(n1705), .B(n21248), .Z(n21247) );
  XOR U20633 ( .A(p_input[1389]), .B(n21246), .Z(n21248) );
  XNOR U20634 ( .A(n21249), .B(n21250), .Z(n21246) );
  AND U20635 ( .A(n1709), .B(n21251), .Z(n21250) );
  XOR U20636 ( .A(n21252), .B(n21253), .Z(n21244) );
  AND U20637 ( .A(n1713), .B(n21243), .Z(n21253) );
  XNOR U20638 ( .A(n21254), .B(n21241), .Z(n21243) );
  XOR U20639 ( .A(n21255), .B(n21256), .Z(n21241) );
  AND U20640 ( .A(n1736), .B(n21257), .Z(n21256) );
  IV U20641 ( .A(n21252), .Z(n21254) );
  XOR U20642 ( .A(n21258), .B(n21259), .Z(n21252) );
  AND U20643 ( .A(n1720), .B(n21251), .Z(n21259) );
  XNOR U20644 ( .A(n21249), .B(n21258), .Z(n21251) );
  XNOR U20645 ( .A(n21260), .B(n21261), .Z(n21249) );
  AND U20646 ( .A(n1724), .B(n21262), .Z(n21261) );
  XOR U20647 ( .A(p_input[1405]), .B(n21260), .Z(n21262) );
  XNOR U20648 ( .A(n21263), .B(n21264), .Z(n21260) );
  AND U20649 ( .A(n1728), .B(n21265), .Z(n21264) );
  XOR U20650 ( .A(n21266), .B(n21267), .Z(n21258) );
  AND U20651 ( .A(n1732), .B(n21257), .Z(n21267) );
  XNOR U20652 ( .A(n21268), .B(n21255), .Z(n21257) );
  XOR U20653 ( .A(n21269), .B(n21270), .Z(n21255) );
  AND U20654 ( .A(n1755), .B(n21271), .Z(n21270) );
  IV U20655 ( .A(n21266), .Z(n21268) );
  XOR U20656 ( .A(n21272), .B(n21273), .Z(n21266) );
  AND U20657 ( .A(n1739), .B(n21265), .Z(n21273) );
  XNOR U20658 ( .A(n21263), .B(n21272), .Z(n21265) );
  XNOR U20659 ( .A(n21274), .B(n21275), .Z(n21263) );
  AND U20660 ( .A(n1743), .B(n21276), .Z(n21275) );
  XOR U20661 ( .A(p_input[1421]), .B(n21274), .Z(n21276) );
  XNOR U20662 ( .A(n21277), .B(n21278), .Z(n21274) );
  AND U20663 ( .A(n1747), .B(n21279), .Z(n21278) );
  XOR U20664 ( .A(n21280), .B(n21281), .Z(n21272) );
  AND U20665 ( .A(n1751), .B(n21271), .Z(n21281) );
  XNOR U20666 ( .A(n21282), .B(n21269), .Z(n21271) );
  XOR U20667 ( .A(n21283), .B(n21284), .Z(n21269) );
  AND U20668 ( .A(n1774), .B(n21285), .Z(n21284) );
  IV U20669 ( .A(n21280), .Z(n21282) );
  XOR U20670 ( .A(n21286), .B(n21287), .Z(n21280) );
  AND U20671 ( .A(n1758), .B(n21279), .Z(n21287) );
  XNOR U20672 ( .A(n21277), .B(n21286), .Z(n21279) );
  XNOR U20673 ( .A(n21288), .B(n21289), .Z(n21277) );
  AND U20674 ( .A(n1762), .B(n21290), .Z(n21289) );
  XOR U20675 ( .A(p_input[1437]), .B(n21288), .Z(n21290) );
  XNOR U20676 ( .A(n21291), .B(n21292), .Z(n21288) );
  AND U20677 ( .A(n1766), .B(n21293), .Z(n21292) );
  XOR U20678 ( .A(n21294), .B(n21295), .Z(n21286) );
  AND U20679 ( .A(n1770), .B(n21285), .Z(n21295) );
  XNOR U20680 ( .A(n21296), .B(n21283), .Z(n21285) );
  XOR U20681 ( .A(n21297), .B(n21298), .Z(n21283) );
  AND U20682 ( .A(n1793), .B(n21299), .Z(n21298) );
  IV U20683 ( .A(n21294), .Z(n21296) );
  XOR U20684 ( .A(n21300), .B(n21301), .Z(n21294) );
  AND U20685 ( .A(n1777), .B(n21293), .Z(n21301) );
  XNOR U20686 ( .A(n21291), .B(n21300), .Z(n21293) );
  XNOR U20687 ( .A(n21302), .B(n21303), .Z(n21291) );
  AND U20688 ( .A(n1781), .B(n21304), .Z(n21303) );
  XOR U20689 ( .A(p_input[1453]), .B(n21302), .Z(n21304) );
  XNOR U20690 ( .A(n21305), .B(n21306), .Z(n21302) );
  AND U20691 ( .A(n1785), .B(n21307), .Z(n21306) );
  XOR U20692 ( .A(n21308), .B(n21309), .Z(n21300) );
  AND U20693 ( .A(n1789), .B(n21299), .Z(n21309) );
  XNOR U20694 ( .A(n21310), .B(n21297), .Z(n21299) );
  XOR U20695 ( .A(n21311), .B(n21312), .Z(n21297) );
  AND U20696 ( .A(n1812), .B(n21313), .Z(n21312) );
  IV U20697 ( .A(n21308), .Z(n21310) );
  XOR U20698 ( .A(n21314), .B(n21315), .Z(n21308) );
  AND U20699 ( .A(n1796), .B(n21307), .Z(n21315) );
  XNOR U20700 ( .A(n21305), .B(n21314), .Z(n21307) );
  XNOR U20701 ( .A(n21316), .B(n21317), .Z(n21305) );
  AND U20702 ( .A(n1800), .B(n21318), .Z(n21317) );
  XOR U20703 ( .A(p_input[1469]), .B(n21316), .Z(n21318) );
  XNOR U20704 ( .A(n21319), .B(n21320), .Z(n21316) );
  AND U20705 ( .A(n1804), .B(n21321), .Z(n21320) );
  XOR U20706 ( .A(n21322), .B(n21323), .Z(n21314) );
  AND U20707 ( .A(n1808), .B(n21313), .Z(n21323) );
  XNOR U20708 ( .A(n21324), .B(n21311), .Z(n21313) );
  XOR U20709 ( .A(n21325), .B(n21326), .Z(n21311) );
  AND U20710 ( .A(n1831), .B(n21327), .Z(n21326) );
  IV U20711 ( .A(n21322), .Z(n21324) );
  XOR U20712 ( .A(n21328), .B(n21329), .Z(n21322) );
  AND U20713 ( .A(n1815), .B(n21321), .Z(n21329) );
  XNOR U20714 ( .A(n21319), .B(n21328), .Z(n21321) );
  XNOR U20715 ( .A(n21330), .B(n21331), .Z(n21319) );
  AND U20716 ( .A(n1819), .B(n21332), .Z(n21331) );
  XOR U20717 ( .A(p_input[1485]), .B(n21330), .Z(n21332) );
  XNOR U20718 ( .A(n21333), .B(n21334), .Z(n21330) );
  AND U20719 ( .A(n1823), .B(n21335), .Z(n21334) );
  XOR U20720 ( .A(n21336), .B(n21337), .Z(n21328) );
  AND U20721 ( .A(n1827), .B(n21327), .Z(n21337) );
  XNOR U20722 ( .A(n21338), .B(n21325), .Z(n21327) );
  XOR U20723 ( .A(n21339), .B(n21340), .Z(n21325) );
  AND U20724 ( .A(n1850), .B(n21341), .Z(n21340) );
  IV U20725 ( .A(n21336), .Z(n21338) );
  XOR U20726 ( .A(n21342), .B(n21343), .Z(n21336) );
  AND U20727 ( .A(n1834), .B(n21335), .Z(n21343) );
  XNOR U20728 ( .A(n21333), .B(n21342), .Z(n21335) );
  XNOR U20729 ( .A(n21344), .B(n21345), .Z(n21333) );
  AND U20730 ( .A(n1838), .B(n21346), .Z(n21345) );
  XOR U20731 ( .A(p_input[1501]), .B(n21344), .Z(n21346) );
  XNOR U20732 ( .A(n21347), .B(n21348), .Z(n21344) );
  AND U20733 ( .A(n1842), .B(n21349), .Z(n21348) );
  XOR U20734 ( .A(n21350), .B(n21351), .Z(n21342) );
  AND U20735 ( .A(n1846), .B(n21341), .Z(n21351) );
  XNOR U20736 ( .A(n21352), .B(n21339), .Z(n21341) );
  XOR U20737 ( .A(n21353), .B(n21354), .Z(n21339) );
  AND U20738 ( .A(n1869), .B(n21355), .Z(n21354) );
  IV U20739 ( .A(n21350), .Z(n21352) );
  XOR U20740 ( .A(n21356), .B(n21357), .Z(n21350) );
  AND U20741 ( .A(n1853), .B(n21349), .Z(n21357) );
  XNOR U20742 ( .A(n21347), .B(n21356), .Z(n21349) );
  XNOR U20743 ( .A(n21358), .B(n21359), .Z(n21347) );
  AND U20744 ( .A(n1857), .B(n21360), .Z(n21359) );
  XOR U20745 ( .A(p_input[1517]), .B(n21358), .Z(n21360) );
  XNOR U20746 ( .A(n21361), .B(n21362), .Z(n21358) );
  AND U20747 ( .A(n1861), .B(n21363), .Z(n21362) );
  XOR U20748 ( .A(n21364), .B(n21365), .Z(n21356) );
  AND U20749 ( .A(n1865), .B(n21355), .Z(n21365) );
  XNOR U20750 ( .A(n21366), .B(n21353), .Z(n21355) );
  XOR U20751 ( .A(n21367), .B(n21368), .Z(n21353) );
  AND U20752 ( .A(n1888), .B(n21369), .Z(n21368) );
  IV U20753 ( .A(n21364), .Z(n21366) );
  XOR U20754 ( .A(n21370), .B(n21371), .Z(n21364) );
  AND U20755 ( .A(n1872), .B(n21363), .Z(n21371) );
  XNOR U20756 ( .A(n21361), .B(n21370), .Z(n21363) );
  XNOR U20757 ( .A(n21372), .B(n21373), .Z(n21361) );
  AND U20758 ( .A(n1876), .B(n21374), .Z(n21373) );
  XOR U20759 ( .A(p_input[1533]), .B(n21372), .Z(n21374) );
  XNOR U20760 ( .A(n21375), .B(n21376), .Z(n21372) );
  AND U20761 ( .A(n1880), .B(n21377), .Z(n21376) );
  XOR U20762 ( .A(n21378), .B(n21379), .Z(n21370) );
  AND U20763 ( .A(n1884), .B(n21369), .Z(n21379) );
  XNOR U20764 ( .A(n21380), .B(n21367), .Z(n21369) );
  XOR U20765 ( .A(n21381), .B(n21382), .Z(n21367) );
  AND U20766 ( .A(n1907), .B(n21383), .Z(n21382) );
  IV U20767 ( .A(n21378), .Z(n21380) );
  XOR U20768 ( .A(n21384), .B(n21385), .Z(n21378) );
  AND U20769 ( .A(n1891), .B(n21377), .Z(n21385) );
  XNOR U20770 ( .A(n21375), .B(n21384), .Z(n21377) );
  XNOR U20771 ( .A(n21386), .B(n21387), .Z(n21375) );
  AND U20772 ( .A(n1895), .B(n21388), .Z(n21387) );
  XOR U20773 ( .A(p_input[1549]), .B(n21386), .Z(n21388) );
  XNOR U20774 ( .A(n21389), .B(n21390), .Z(n21386) );
  AND U20775 ( .A(n1899), .B(n21391), .Z(n21390) );
  XOR U20776 ( .A(n21392), .B(n21393), .Z(n21384) );
  AND U20777 ( .A(n1903), .B(n21383), .Z(n21393) );
  XNOR U20778 ( .A(n21394), .B(n21381), .Z(n21383) );
  XOR U20779 ( .A(n21395), .B(n21396), .Z(n21381) );
  AND U20780 ( .A(n1926), .B(n21397), .Z(n21396) );
  IV U20781 ( .A(n21392), .Z(n21394) );
  XOR U20782 ( .A(n21398), .B(n21399), .Z(n21392) );
  AND U20783 ( .A(n1910), .B(n21391), .Z(n21399) );
  XNOR U20784 ( .A(n21389), .B(n21398), .Z(n21391) );
  XNOR U20785 ( .A(n21400), .B(n21401), .Z(n21389) );
  AND U20786 ( .A(n1914), .B(n21402), .Z(n21401) );
  XOR U20787 ( .A(p_input[1565]), .B(n21400), .Z(n21402) );
  XNOR U20788 ( .A(n21403), .B(n21404), .Z(n21400) );
  AND U20789 ( .A(n1918), .B(n21405), .Z(n21404) );
  XOR U20790 ( .A(n21406), .B(n21407), .Z(n21398) );
  AND U20791 ( .A(n1922), .B(n21397), .Z(n21407) );
  XNOR U20792 ( .A(n21408), .B(n21395), .Z(n21397) );
  XOR U20793 ( .A(n21409), .B(n21410), .Z(n21395) );
  AND U20794 ( .A(n1945), .B(n21411), .Z(n21410) );
  IV U20795 ( .A(n21406), .Z(n21408) );
  XOR U20796 ( .A(n21412), .B(n21413), .Z(n21406) );
  AND U20797 ( .A(n1929), .B(n21405), .Z(n21413) );
  XNOR U20798 ( .A(n21403), .B(n21412), .Z(n21405) );
  XNOR U20799 ( .A(n21414), .B(n21415), .Z(n21403) );
  AND U20800 ( .A(n1933), .B(n21416), .Z(n21415) );
  XOR U20801 ( .A(p_input[1581]), .B(n21414), .Z(n21416) );
  XNOR U20802 ( .A(n21417), .B(n21418), .Z(n21414) );
  AND U20803 ( .A(n1937), .B(n21419), .Z(n21418) );
  XOR U20804 ( .A(n21420), .B(n21421), .Z(n21412) );
  AND U20805 ( .A(n1941), .B(n21411), .Z(n21421) );
  XNOR U20806 ( .A(n21422), .B(n21409), .Z(n21411) );
  XOR U20807 ( .A(n21423), .B(n21424), .Z(n21409) );
  AND U20808 ( .A(n1964), .B(n21425), .Z(n21424) );
  IV U20809 ( .A(n21420), .Z(n21422) );
  XOR U20810 ( .A(n21426), .B(n21427), .Z(n21420) );
  AND U20811 ( .A(n1948), .B(n21419), .Z(n21427) );
  XNOR U20812 ( .A(n21417), .B(n21426), .Z(n21419) );
  XNOR U20813 ( .A(n21428), .B(n21429), .Z(n21417) );
  AND U20814 ( .A(n1952), .B(n21430), .Z(n21429) );
  XOR U20815 ( .A(p_input[1597]), .B(n21428), .Z(n21430) );
  XNOR U20816 ( .A(n21431), .B(n21432), .Z(n21428) );
  AND U20817 ( .A(n1956), .B(n21433), .Z(n21432) );
  XOR U20818 ( .A(n21434), .B(n21435), .Z(n21426) );
  AND U20819 ( .A(n1960), .B(n21425), .Z(n21435) );
  XNOR U20820 ( .A(n21436), .B(n21423), .Z(n21425) );
  XOR U20821 ( .A(n21437), .B(n21438), .Z(n21423) );
  AND U20822 ( .A(n1983), .B(n21439), .Z(n21438) );
  IV U20823 ( .A(n21434), .Z(n21436) );
  XOR U20824 ( .A(n21440), .B(n21441), .Z(n21434) );
  AND U20825 ( .A(n1967), .B(n21433), .Z(n21441) );
  XNOR U20826 ( .A(n21431), .B(n21440), .Z(n21433) );
  XNOR U20827 ( .A(n21442), .B(n21443), .Z(n21431) );
  AND U20828 ( .A(n1971), .B(n21444), .Z(n21443) );
  XOR U20829 ( .A(p_input[1613]), .B(n21442), .Z(n21444) );
  XNOR U20830 ( .A(n21445), .B(n21446), .Z(n21442) );
  AND U20831 ( .A(n1975), .B(n21447), .Z(n21446) );
  XOR U20832 ( .A(n21448), .B(n21449), .Z(n21440) );
  AND U20833 ( .A(n1979), .B(n21439), .Z(n21449) );
  XNOR U20834 ( .A(n21450), .B(n21437), .Z(n21439) );
  XOR U20835 ( .A(n21451), .B(n21452), .Z(n21437) );
  AND U20836 ( .A(n2002), .B(n21453), .Z(n21452) );
  IV U20837 ( .A(n21448), .Z(n21450) );
  XOR U20838 ( .A(n21454), .B(n21455), .Z(n21448) );
  AND U20839 ( .A(n1986), .B(n21447), .Z(n21455) );
  XNOR U20840 ( .A(n21445), .B(n21454), .Z(n21447) );
  XNOR U20841 ( .A(n21456), .B(n21457), .Z(n21445) );
  AND U20842 ( .A(n1990), .B(n21458), .Z(n21457) );
  XOR U20843 ( .A(p_input[1629]), .B(n21456), .Z(n21458) );
  XNOR U20844 ( .A(n21459), .B(n21460), .Z(n21456) );
  AND U20845 ( .A(n1994), .B(n21461), .Z(n21460) );
  XOR U20846 ( .A(n21462), .B(n21463), .Z(n21454) );
  AND U20847 ( .A(n1998), .B(n21453), .Z(n21463) );
  XNOR U20848 ( .A(n21464), .B(n21451), .Z(n21453) );
  XOR U20849 ( .A(n21465), .B(n21466), .Z(n21451) );
  AND U20850 ( .A(n2021), .B(n21467), .Z(n21466) );
  IV U20851 ( .A(n21462), .Z(n21464) );
  XOR U20852 ( .A(n21468), .B(n21469), .Z(n21462) );
  AND U20853 ( .A(n2005), .B(n21461), .Z(n21469) );
  XNOR U20854 ( .A(n21459), .B(n21468), .Z(n21461) );
  XNOR U20855 ( .A(n21470), .B(n21471), .Z(n21459) );
  AND U20856 ( .A(n2009), .B(n21472), .Z(n21471) );
  XOR U20857 ( .A(p_input[1645]), .B(n21470), .Z(n21472) );
  XNOR U20858 ( .A(n21473), .B(n21474), .Z(n21470) );
  AND U20859 ( .A(n2013), .B(n21475), .Z(n21474) );
  XOR U20860 ( .A(n21476), .B(n21477), .Z(n21468) );
  AND U20861 ( .A(n2017), .B(n21467), .Z(n21477) );
  XNOR U20862 ( .A(n21478), .B(n21465), .Z(n21467) );
  XOR U20863 ( .A(n21479), .B(n21480), .Z(n21465) );
  AND U20864 ( .A(n2040), .B(n21481), .Z(n21480) );
  IV U20865 ( .A(n21476), .Z(n21478) );
  XOR U20866 ( .A(n21482), .B(n21483), .Z(n21476) );
  AND U20867 ( .A(n2024), .B(n21475), .Z(n21483) );
  XNOR U20868 ( .A(n21473), .B(n21482), .Z(n21475) );
  XNOR U20869 ( .A(n21484), .B(n21485), .Z(n21473) );
  AND U20870 ( .A(n2028), .B(n21486), .Z(n21485) );
  XOR U20871 ( .A(p_input[1661]), .B(n21484), .Z(n21486) );
  XNOR U20872 ( .A(n21487), .B(n21488), .Z(n21484) );
  AND U20873 ( .A(n2032), .B(n21489), .Z(n21488) );
  XOR U20874 ( .A(n21490), .B(n21491), .Z(n21482) );
  AND U20875 ( .A(n2036), .B(n21481), .Z(n21491) );
  XNOR U20876 ( .A(n21492), .B(n21479), .Z(n21481) );
  XOR U20877 ( .A(n21493), .B(n21494), .Z(n21479) );
  AND U20878 ( .A(n2059), .B(n21495), .Z(n21494) );
  IV U20879 ( .A(n21490), .Z(n21492) );
  XOR U20880 ( .A(n21496), .B(n21497), .Z(n21490) );
  AND U20881 ( .A(n2043), .B(n21489), .Z(n21497) );
  XNOR U20882 ( .A(n21487), .B(n21496), .Z(n21489) );
  XNOR U20883 ( .A(n21498), .B(n21499), .Z(n21487) );
  AND U20884 ( .A(n2047), .B(n21500), .Z(n21499) );
  XOR U20885 ( .A(p_input[1677]), .B(n21498), .Z(n21500) );
  XNOR U20886 ( .A(n21501), .B(n21502), .Z(n21498) );
  AND U20887 ( .A(n2051), .B(n21503), .Z(n21502) );
  XOR U20888 ( .A(n21504), .B(n21505), .Z(n21496) );
  AND U20889 ( .A(n2055), .B(n21495), .Z(n21505) );
  XNOR U20890 ( .A(n21506), .B(n21493), .Z(n21495) );
  XOR U20891 ( .A(n21507), .B(n21508), .Z(n21493) );
  AND U20892 ( .A(n2078), .B(n21509), .Z(n21508) );
  IV U20893 ( .A(n21504), .Z(n21506) );
  XOR U20894 ( .A(n21510), .B(n21511), .Z(n21504) );
  AND U20895 ( .A(n2062), .B(n21503), .Z(n21511) );
  XNOR U20896 ( .A(n21501), .B(n21510), .Z(n21503) );
  XNOR U20897 ( .A(n21512), .B(n21513), .Z(n21501) );
  AND U20898 ( .A(n2066), .B(n21514), .Z(n21513) );
  XOR U20899 ( .A(p_input[1693]), .B(n21512), .Z(n21514) );
  XNOR U20900 ( .A(n21515), .B(n21516), .Z(n21512) );
  AND U20901 ( .A(n2070), .B(n21517), .Z(n21516) );
  XOR U20902 ( .A(n21518), .B(n21519), .Z(n21510) );
  AND U20903 ( .A(n2074), .B(n21509), .Z(n21519) );
  XNOR U20904 ( .A(n21520), .B(n21507), .Z(n21509) );
  XOR U20905 ( .A(n21521), .B(n21522), .Z(n21507) );
  AND U20906 ( .A(n2097), .B(n21523), .Z(n21522) );
  IV U20907 ( .A(n21518), .Z(n21520) );
  XOR U20908 ( .A(n21524), .B(n21525), .Z(n21518) );
  AND U20909 ( .A(n2081), .B(n21517), .Z(n21525) );
  XNOR U20910 ( .A(n21515), .B(n21524), .Z(n21517) );
  XNOR U20911 ( .A(n21526), .B(n21527), .Z(n21515) );
  AND U20912 ( .A(n2085), .B(n21528), .Z(n21527) );
  XOR U20913 ( .A(p_input[1709]), .B(n21526), .Z(n21528) );
  XNOR U20914 ( .A(n21529), .B(n21530), .Z(n21526) );
  AND U20915 ( .A(n2089), .B(n21531), .Z(n21530) );
  XOR U20916 ( .A(n21532), .B(n21533), .Z(n21524) );
  AND U20917 ( .A(n2093), .B(n21523), .Z(n21533) );
  XNOR U20918 ( .A(n21534), .B(n21521), .Z(n21523) );
  XOR U20919 ( .A(n21535), .B(n21536), .Z(n21521) );
  AND U20920 ( .A(n2116), .B(n21537), .Z(n21536) );
  IV U20921 ( .A(n21532), .Z(n21534) );
  XOR U20922 ( .A(n21538), .B(n21539), .Z(n21532) );
  AND U20923 ( .A(n2100), .B(n21531), .Z(n21539) );
  XNOR U20924 ( .A(n21529), .B(n21538), .Z(n21531) );
  XNOR U20925 ( .A(n21540), .B(n21541), .Z(n21529) );
  AND U20926 ( .A(n2104), .B(n21542), .Z(n21541) );
  XOR U20927 ( .A(p_input[1725]), .B(n21540), .Z(n21542) );
  XNOR U20928 ( .A(n21543), .B(n21544), .Z(n21540) );
  AND U20929 ( .A(n2108), .B(n21545), .Z(n21544) );
  XOR U20930 ( .A(n21546), .B(n21547), .Z(n21538) );
  AND U20931 ( .A(n2112), .B(n21537), .Z(n21547) );
  XNOR U20932 ( .A(n21548), .B(n21535), .Z(n21537) );
  XOR U20933 ( .A(n21549), .B(n21550), .Z(n21535) );
  AND U20934 ( .A(n2135), .B(n21551), .Z(n21550) );
  IV U20935 ( .A(n21546), .Z(n21548) );
  XOR U20936 ( .A(n21552), .B(n21553), .Z(n21546) );
  AND U20937 ( .A(n2119), .B(n21545), .Z(n21553) );
  XNOR U20938 ( .A(n21543), .B(n21552), .Z(n21545) );
  XNOR U20939 ( .A(n21554), .B(n21555), .Z(n21543) );
  AND U20940 ( .A(n2123), .B(n21556), .Z(n21555) );
  XOR U20941 ( .A(p_input[1741]), .B(n21554), .Z(n21556) );
  XNOR U20942 ( .A(n21557), .B(n21558), .Z(n21554) );
  AND U20943 ( .A(n2127), .B(n21559), .Z(n21558) );
  XOR U20944 ( .A(n21560), .B(n21561), .Z(n21552) );
  AND U20945 ( .A(n2131), .B(n21551), .Z(n21561) );
  XNOR U20946 ( .A(n21562), .B(n21549), .Z(n21551) );
  XOR U20947 ( .A(n21563), .B(n21564), .Z(n21549) );
  AND U20948 ( .A(n2154), .B(n21565), .Z(n21564) );
  IV U20949 ( .A(n21560), .Z(n21562) );
  XOR U20950 ( .A(n21566), .B(n21567), .Z(n21560) );
  AND U20951 ( .A(n2138), .B(n21559), .Z(n21567) );
  XNOR U20952 ( .A(n21557), .B(n21566), .Z(n21559) );
  XNOR U20953 ( .A(n21568), .B(n21569), .Z(n21557) );
  AND U20954 ( .A(n2142), .B(n21570), .Z(n21569) );
  XOR U20955 ( .A(p_input[1757]), .B(n21568), .Z(n21570) );
  XNOR U20956 ( .A(n21571), .B(n21572), .Z(n21568) );
  AND U20957 ( .A(n2146), .B(n21573), .Z(n21572) );
  XOR U20958 ( .A(n21574), .B(n21575), .Z(n21566) );
  AND U20959 ( .A(n2150), .B(n21565), .Z(n21575) );
  XNOR U20960 ( .A(n21576), .B(n21563), .Z(n21565) );
  XOR U20961 ( .A(n21577), .B(n21578), .Z(n21563) );
  AND U20962 ( .A(n2173), .B(n21579), .Z(n21578) );
  IV U20963 ( .A(n21574), .Z(n21576) );
  XOR U20964 ( .A(n21580), .B(n21581), .Z(n21574) );
  AND U20965 ( .A(n2157), .B(n21573), .Z(n21581) );
  XNOR U20966 ( .A(n21571), .B(n21580), .Z(n21573) );
  XNOR U20967 ( .A(n21582), .B(n21583), .Z(n21571) );
  AND U20968 ( .A(n2161), .B(n21584), .Z(n21583) );
  XOR U20969 ( .A(p_input[1773]), .B(n21582), .Z(n21584) );
  XNOR U20970 ( .A(n21585), .B(n21586), .Z(n21582) );
  AND U20971 ( .A(n2165), .B(n21587), .Z(n21586) );
  XOR U20972 ( .A(n21588), .B(n21589), .Z(n21580) );
  AND U20973 ( .A(n2169), .B(n21579), .Z(n21589) );
  XNOR U20974 ( .A(n21590), .B(n21577), .Z(n21579) );
  XOR U20975 ( .A(n21591), .B(n21592), .Z(n21577) );
  AND U20976 ( .A(n2192), .B(n21593), .Z(n21592) );
  IV U20977 ( .A(n21588), .Z(n21590) );
  XOR U20978 ( .A(n21594), .B(n21595), .Z(n21588) );
  AND U20979 ( .A(n2176), .B(n21587), .Z(n21595) );
  XNOR U20980 ( .A(n21585), .B(n21594), .Z(n21587) );
  XNOR U20981 ( .A(n21596), .B(n21597), .Z(n21585) );
  AND U20982 ( .A(n2180), .B(n21598), .Z(n21597) );
  XOR U20983 ( .A(p_input[1789]), .B(n21596), .Z(n21598) );
  XNOR U20984 ( .A(n21599), .B(n21600), .Z(n21596) );
  AND U20985 ( .A(n2184), .B(n21601), .Z(n21600) );
  XOR U20986 ( .A(n21602), .B(n21603), .Z(n21594) );
  AND U20987 ( .A(n2188), .B(n21593), .Z(n21603) );
  XNOR U20988 ( .A(n21604), .B(n21591), .Z(n21593) );
  XOR U20989 ( .A(n21605), .B(n21606), .Z(n21591) );
  AND U20990 ( .A(n2211), .B(n21607), .Z(n21606) );
  IV U20991 ( .A(n21602), .Z(n21604) );
  XOR U20992 ( .A(n21608), .B(n21609), .Z(n21602) );
  AND U20993 ( .A(n2195), .B(n21601), .Z(n21609) );
  XNOR U20994 ( .A(n21599), .B(n21608), .Z(n21601) );
  XNOR U20995 ( .A(n21610), .B(n21611), .Z(n21599) );
  AND U20996 ( .A(n2199), .B(n21612), .Z(n21611) );
  XOR U20997 ( .A(p_input[1805]), .B(n21610), .Z(n21612) );
  XNOR U20998 ( .A(n21613), .B(n21614), .Z(n21610) );
  AND U20999 ( .A(n2203), .B(n21615), .Z(n21614) );
  XOR U21000 ( .A(n21616), .B(n21617), .Z(n21608) );
  AND U21001 ( .A(n2207), .B(n21607), .Z(n21617) );
  XNOR U21002 ( .A(n21618), .B(n21605), .Z(n21607) );
  XOR U21003 ( .A(n21619), .B(n21620), .Z(n21605) );
  AND U21004 ( .A(n2230), .B(n21621), .Z(n21620) );
  IV U21005 ( .A(n21616), .Z(n21618) );
  XOR U21006 ( .A(n21622), .B(n21623), .Z(n21616) );
  AND U21007 ( .A(n2214), .B(n21615), .Z(n21623) );
  XNOR U21008 ( .A(n21613), .B(n21622), .Z(n21615) );
  XNOR U21009 ( .A(n21624), .B(n21625), .Z(n21613) );
  AND U21010 ( .A(n2218), .B(n21626), .Z(n21625) );
  XOR U21011 ( .A(p_input[1821]), .B(n21624), .Z(n21626) );
  XNOR U21012 ( .A(n21627), .B(n21628), .Z(n21624) );
  AND U21013 ( .A(n2222), .B(n21629), .Z(n21628) );
  XOR U21014 ( .A(n21630), .B(n21631), .Z(n21622) );
  AND U21015 ( .A(n2226), .B(n21621), .Z(n21631) );
  XNOR U21016 ( .A(n21632), .B(n21619), .Z(n21621) );
  XOR U21017 ( .A(n21633), .B(n21634), .Z(n21619) );
  AND U21018 ( .A(n2249), .B(n21635), .Z(n21634) );
  IV U21019 ( .A(n21630), .Z(n21632) );
  XOR U21020 ( .A(n21636), .B(n21637), .Z(n21630) );
  AND U21021 ( .A(n2233), .B(n21629), .Z(n21637) );
  XNOR U21022 ( .A(n21627), .B(n21636), .Z(n21629) );
  XNOR U21023 ( .A(n21638), .B(n21639), .Z(n21627) );
  AND U21024 ( .A(n2237), .B(n21640), .Z(n21639) );
  XOR U21025 ( .A(p_input[1837]), .B(n21638), .Z(n21640) );
  XNOR U21026 ( .A(n21641), .B(n21642), .Z(n21638) );
  AND U21027 ( .A(n2241), .B(n21643), .Z(n21642) );
  XOR U21028 ( .A(n21644), .B(n21645), .Z(n21636) );
  AND U21029 ( .A(n2245), .B(n21635), .Z(n21645) );
  XNOR U21030 ( .A(n21646), .B(n21633), .Z(n21635) );
  XOR U21031 ( .A(n21647), .B(n21648), .Z(n21633) );
  AND U21032 ( .A(n2268), .B(n21649), .Z(n21648) );
  IV U21033 ( .A(n21644), .Z(n21646) );
  XOR U21034 ( .A(n21650), .B(n21651), .Z(n21644) );
  AND U21035 ( .A(n2252), .B(n21643), .Z(n21651) );
  XNOR U21036 ( .A(n21641), .B(n21650), .Z(n21643) );
  XNOR U21037 ( .A(n21652), .B(n21653), .Z(n21641) );
  AND U21038 ( .A(n2256), .B(n21654), .Z(n21653) );
  XOR U21039 ( .A(p_input[1853]), .B(n21652), .Z(n21654) );
  XNOR U21040 ( .A(n21655), .B(n21656), .Z(n21652) );
  AND U21041 ( .A(n2260), .B(n21657), .Z(n21656) );
  XOR U21042 ( .A(n21658), .B(n21659), .Z(n21650) );
  AND U21043 ( .A(n2264), .B(n21649), .Z(n21659) );
  XNOR U21044 ( .A(n21660), .B(n21647), .Z(n21649) );
  XOR U21045 ( .A(n21661), .B(n21662), .Z(n21647) );
  AND U21046 ( .A(n2287), .B(n21663), .Z(n21662) );
  IV U21047 ( .A(n21658), .Z(n21660) );
  XOR U21048 ( .A(n21664), .B(n21665), .Z(n21658) );
  AND U21049 ( .A(n2271), .B(n21657), .Z(n21665) );
  XNOR U21050 ( .A(n21655), .B(n21664), .Z(n21657) );
  XNOR U21051 ( .A(n21666), .B(n21667), .Z(n21655) );
  AND U21052 ( .A(n2275), .B(n21668), .Z(n21667) );
  XOR U21053 ( .A(p_input[1869]), .B(n21666), .Z(n21668) );
  XNOR U21054 ( .A(n21669), .B(n21670), .Z(n21666) );
  AND U21055 ( .A(n2279), .B(n21671), .Z(n21670) );
  XOR U21056 ( .A(n21672), .B(n21673), .Z(n21664) );
  AND U21057 ( .A(n2283), .B(n21663), .Z(n21673) );
  XNOR U21058 ( .A(n21674), .B(n21661), .Z(n21663) );
  XOR U21059 ( .A(n21675), .B(n21676), .Z(n21661) );
  AND U21060 ( .A(n2306), .B(n21677), .Z(n21676) );
  IV U21061 ( .A(n21672), .Z(n21674) );
  XOR U21062 ( .A(n21678), .B(n21679), .Z(n21672) );
  AND U21063 ( .A(n2290), .B(n21671), .Z(n21679) );
  XNOR U21064 ( .A(n21669), .B(n21678), .Z(n21671) );
  XNOR U21065 ( .A(n21680), .B(n21681), .Z(n21669) );
  AND U21066 ( .A(n2294), .B(n21682), .Z(n21681) );
  XOR U21067 ( .A(p_input[1885]), .B(n21680), .Z(n21682) );
  XNOR U21068 ( .A(n21683), .B(n21684), .Z(n21680) );
  AND U21069 ( .A(n2298), .B(n21685), .Z(n21684) );
  XOR U21070 ( .A(n21686), .B(n21687), .Z(n21678) );
  AND U21071 ( .A(n2302), .B(n21677), .Z(n21687) );
  XNOR U21072 ( .A(n21688), .B(n21675), .Z(n21677) );
  XOR U21073 ( .A(n21689), .B(n21690), .Z(n21675) );
  AND U21074 ( .A(n2325), .B(n21691), .Z(n21690) );
  IV U21075 ( .A(n21686), .Z(n21688) );
  XOR U21076 ( .A(n21692), .B(n21693), .Z(n21686) );
  AND U21077 ( .A(n2309), .B(n21685), .Z(n21693) );
  XNOR U21078 ( .A(n21683), .B(n21692), .Z(n21685) );
  XNOR U21079 ( .A(n21694), .B(n21695), .Z(n21683) );
  AND U21080 ( .A(n2313), .B(n21696), .Z(n21695) );
  XOR U21081 ( .A(p_input[1901]), .B(n21694), .Z(n21696) );
  XNOR U21082 ( .A(n21697), .B(n21698), .Z(n21694) );
  AND U21083 ( .A(n2317), .B(n21699), .Z(n21698) );
  XOR U21084 ( .A(n21700), .B(n21701), .Z(n21692) );
  AND U21085 ( .A(n2321), .B(n21691), .Z(n21701) );
  XNOR U21086 ( .A(n21702), .B(n21689), .Z(n21691) );
  XOR U21087 ( .A(n21703), .B(n21704), .Z(n21689) );
  AND U21088 ( .A(n2344), .B(n21705), .Z(n21704) );
  IV U21089 ( .A(n21700), .Z(n21702) );
  XOR U21090 ( .A(n21706), .B(n21707), .Z(n21700) );
  AND U21091 ( .A(n2328), .B(n21699), .Z(n21707) );
  XNOR U21092 ( .A(n21697), .B(n21706), .Z(n21699) );
  XNOR U21093 ( .A(n21708), .B(n21709), .Z(n21697) );
  AND U21094 ( .A(n2332), .B(n21710), .Z(n21709) );
  XOR U21095 ( .A(p_input[1917]), .B(n21708), .Z(n21710) );
  XNOR U21096 ( .A(n21711), .B(n21712), .Z(n21708) );
  AND U21097 ( .A(n2336), .B(n21713), .Z(n21712) );
  XOR U21098 ( .A(n21714), .B(n21715), .Z(n21706) );
  AND U21099 ( .A(n2340), .B(n21705), .Z(n21715) );
  XNOR U21100 ( .A(n21716), .B(n21703), .Z(n21705) );
  XOR U21101 ( .A(n21717), .B(n21718), .Z(n21703) );
  AND U21102 ( .A(n2363), .B(n21719), .Z(n21718) );
  IV U21103 ( .A(n21714), .Z(n21716) );
  XOR U21104 ( .A(n21720), .B(n21721), .Z(n21714) );
  AND U21105 ( .A(n2347), .B(n21713), .Z(n21721) );
  XNOR U21106 ( .A(n21711), .B(n21720), .Z(n21713) );
  XNOR U21107 ( .A(n21722), .B(n21723), .Z(n21711) );
  AND U21108 ( .A(n2351), .B(n21724), .Z(n21723) );
  XOR U21109 ( .A(p_input[1933]), .B(n21722), .Z(n21724) );
  XNOR U21110 ( .A(n21725), .B(n21726), .Z(n21722) );
  AND U21111 ( .A(n2355), .B(n21727), .Z(n21726) );
  XOR U21112 ( .A(n21728), .B(n21729), .Z(n21720) );
  AND U21113 ( .A(n2359), .B(n21719), .Z(n21729) );
  XNOR U21114 ( .A(n21730), .B(n21717), .Z(n21719) );
  XOR U21115 ( .A(n21731), .B(n21732), .Z(n21717) );
  AND U21116 ( .A(n2382), .B(n21733), .Z(n21732) );
  IV U21117 ( .A(n21728), .Z(n21730) );
  XOR U21118 ( .A(n21734), .B(n21735), .Z(n21728) );
  AND U21119 ( .A(n2366), .B(n21727), .Z(n21735) );
  XNOR U21120 ( .A(n21725), .B(n21734), .Z(n21727) );
  XNOR U21121 ( .A(n21736), .B(n21737), .Z(n21725) );
  AND U21122 ( .A(n2370), .B(n21738), .Z(n21737) );
  XOR U21123 ( .A(p_input[1949]), .B(n21736), .Z(n21738) );
  XNOR U21124 ( .A(n21739), .B(n21740), .Z(n21736) );
  AND U21125 ( .A(n2374), .B(n21741), .Z(n21740) );
  XOR U21126 ( .A(n21742), .B(n21743), .Z(n21734) );
  AND U21127 ( .A(n2378), .B(n21733), .Z(n21743) );
  XNOR U21128 ( .A(n21744), .B(n21731), .Z(n21733) );
  XOR U21129 ( .A(n21745), .B(n21746), .Z(n21731) );
  AND U21130 ( .A(n2401), .B(n21747), .Z(n21746) );
  IV U21131 ( .A(n21742), .Z(n21744) );
  XOR U21132 ( .A(n21748), .B(n21749), .Z(n21742) );
  AND U21133 ( .A(n2385), .B(n21741), .Z(n21749) );
  XNOR U21134 ( .A(n21739), .B(n21748), .Z(n21741) );
  XNOR U21135 ( .A(n21750), .B(n21751), .Z(n21739) );
  AND U21136 ( .A(n2389), .B(n21752), .Z(n21751) );
  XOR U21137 ( .A(p_input[1965]), .B(n21750), .Z(n21752) );
  XNOR U21138 ( .A(n21753), .B(n21754), .Z(n21750) );
  AND U21139 ( .A(n2393), .B(n21755), .Z(n21754) );
  XOR U21140 ( .A(n21756), .B(n21757), .Z(n21748) );
  AND U21141 ( .A(n2397), .B(n21747), .Z(n21757) );
  XNOR U21142 ( .A(n21758), .B(n21745), .Z(n21747) );
  XOR U21143 ( .A(n21759), .B(n21760), .Z(n21745) );
  AND U21144 ( .A(n2420), .B(n21761), .Z(n21760) );
  IV U21145 ( .A(n21756), .Z(n21758) );
  XOR U21146 ( .A(n21762), .B(n21763), .Z(n21756) );
  AND U21147 ( .A(n2404), .B(n21755), .Z(n21763) );
  XNOR U21148 ( .A(n21753), .B(n21762), .Z(n21755) );
  XNOR U21149 ( .A(n21764), .B(n21765), .Z(n21753) );
  AND U21150 ( .A(n2408), .B(n21766), .Z(n21765) );
  XOR U21151 ( .A(p_input[1981]), .B(n21764), .Z(n21766) );
  XNOR U21152 ( .A(n21767), .B(n21768), .Z(n21764) );
  AND U21153 ( .A(n2412), .B(n21769), .Z(n21768) );
  XOR U21154 ( .A(n21770), .B(n21771), .Z(n21762) );
  AND U21155 ( .A(n2416), .B(n21761), .Z(n21771) );
  XNOR U21156 ( .A(n21772), .B(n21759), .Z(n21761) );
  XOR U21157 ( .A(n21773), .B(n21774), .Z(n21759) );
  AND U21158 ( .A(n2438), .B(n21775), .Z(n21774) );
  IV U21159 ( .A(n21770), .Z(n21772) );
  XOR U21160 ( .A(n21776), .B(n21777), .Z(n21770) );
  AND U21161 ( .A(n2423), .B(n21769), .Z(n21777) );
  XNOR U21162 ( .A(n21767), .B(n21776), .Z(n21769) );
  XNOR U21163 ( .A(n21778), .B(n21779), .Z(n21767) );
  AND U21164 ( .A(n2427), .B(n21780), .Z(n21779) );
  XOR U21165 ( .A(p_input[1997]), .B(n21778), .Z(n21780) );
  XOR U21166 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n21781), 
        .Z(n21778) );
  AND U21167 ( .A(n2430), .B(n21782), .Z(n21781) );
  XOR U21168 ( .A(n21783), .B(n21784), .Z(n21776) );
  AND U21169 ( .A(n2434), .B(n21775), .Z(n21784) );
  XNOR U21170 ( .A(n21785), .B(n21773), .Z(n21775) );
  XOR U21171 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n21786), .Z(n21773) );
  AND U21172 ( .A(n2446), .B(n21787), .Z(n21786) );
  IV U21173 ( .A(n21783), .Z(n21785) );
  XOR U21174 ( .A(n21788), .B(n21789), .Z(n21783) );
  AND U21175 ( .A(n2441), .B(n21782), .Z(n21789) );
  XOR U21176 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n21788), 
        .Z(n21782) );
  XOR U21177 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n21790), 
        .Z(n21788) );
  AND U21178 ( .A(n2443), .B(n21787), .Z(n21790) );
  XOR U21179 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n21787) );
  XOR U21180 ( .A(n55), .B(n21791), .Z(o[12]) );
  AND U21181 ( .A(n62), .B(n21792), .Z(n55) );
  XOR U21182 ( .A(n56), .B(n21791), .Z(n21792) );
  XOR U21183 ( .A(n21793), .B(n21794), .Z(n21791) );
  AND U21184 ( .A(n82), .B(n21795), .Z(n21794) );
  XOR U21185 ( .A(n21796), .B(n19), .Z(n56) );
  AND U21186 ( .A(n65), .B(n21797), .Z(n19) );
  XOR U21187 ( .A(n20), .B(n21796), .Z(n21797) );
  XOR U21188 ( .A(n21798), .B(n21799), .Z(n20) );
  AND U21189 ( .A(n70), .B(n21800), .Z(n21799) );
  XOR U21190 ( .A(p_input[12]), .B(n21798), .Z(n21800) );
  XNOR U21191 ( .A(n21801), .B(n21802), .Z(n21798) );
  AND U21192 ( .A(n74), .B(n21803), .Z(n21802) );
  XOR U21193 ( .A(n21804), .B(n21805), .Z(n21796) );
  AND U21194 ( .A(n78), .B(n21795), .Z(n21805) );
  XNOR U21195 ( .A(n21806), .B(n21793), .Z(n21795) );
  XOR U21196 ( .A(n21807), .B(n21808), .Z(n21793) );
  AND U21197 ( .A(n102), .B(n21809), .Z(n21808) );
  IV U21198 ( .A(n21804), .Z(n21806) );
  XOR U21199 ( .A(n21810), .B(n21811), .Z(n21804) );
  AND U21200 ( .A(n86), .B(n21803), .Z(n21811) );
  XNOR U21201 ( .A(n21801), .B(n21810), .Z(n21803) );
  XNOR U21202 ( .A(n21812), .B(n21813), .Z(n21801) );
  AND U21203 ( .A(n90), .B(n21814), .Z(n21813) );
  XOR U21204 ( .A(p_input[28]), .B(n21812), .Z(n21814) );
  XNOR U21205 ( .A(n21815), .B(n21816), .Z(n21812) );
  AND U21206 ( .A(n94), .B(n21817), .Z(n21816) );
  XOR U21207 ( .A(n21818), .B(n21819), .Z(n21810) );
  AND U21208 ( .A(n98), .B(n21809), .Z(n21819) );
  XNOR U21209 ( .A(n21820), .B(n21807), .Z(n21809) );
  XOR U21210 ( .A(n21821), .B(n21822), .Z(n21807) );
  AND U21211 ( .A(n121), .B(n21823), .Z(n21822) );
  IV U21212 ( .A(n21818), .Z(n21820) );
  XOR U21213 ( .A(n21824), .B(n21825), .Z(n21818) );
  AND U21214 ( .A(n105), .B(n21817), .Z(n21825) );
  XNOR U21215 ( .A(n21815), .B(n21824), .Z(n21817) );
  XNOR U21216 ( .A(n21826), .B(n21827), .Z(n21815) );
  AND U21217 ( .A(n109), .B(n21828), .Z(n21827) );
  XOR U21218 ( .A(p_input[44]), .B(n21826), .Z(n21828) );
  XNOR U21219 ( .A(n21829), .B(n21830), .Z(n21826) );
  AND U21220 ( .A(n113), .B(n21831), .Z(n21830) );
  XOR U21221 ( .A(n21832), .B(n21833), .Z(n21824) );
  AND U21222 ( .A(n117), .B(n21823), .Z(n21833) );
  XNOR U21223 ( .A(n21834), .B(n21821), .Z(n21823) );
  XOR U21224 ( .A(n21835), .B(n21836), .Z(n21821) );
  AND U21225 ( .A(n140), .B(n21837), .Z(n21836) );
  IV U21226 ( .A(n21832), .Z(n21834) );
  XOR U21227 ( .A(n21838), .B(n21839), .Z(n21832) );
  AND U21228 ( .A(n124), .B(n21831), .Z(n21839) );
  XNOR U21229 ( .A(n21829), .B(n21838), .Z(n21831) );
  XNOR U21230 ( .A(n21840), .B(n21841), .Z(n21829) );
  AND U21231 ( .A(n128), .B(n21842), .Z(n21841) );
  XOR U21232 ( .A(p_input[60]), .B(n21840), .Z(n21842) );
  XNOR U21233 ( .A(n21843), .B(n21844), .Z(n21840) );
  AND U21234 ( .A(n132), .B(n21845), .Z(n21844) );
  XOR U21235 ( .A(n21846), .B(n21847), .Z(n21838) );
  AND U21236 ( .A(n136), .B(n21837), .Z(n21847) );
  XNOR U21237 ( .A(n21848), .B(n21835), .Z(n21837) );
  XOR U21238 ( .A(n21849), .B(n21850), .Z(n21835) );
  AND U21239 ( .A(n159), .B(n21851), .Z(n21850) );
  IV U21240 ( .A(n21846), .Z(n21848) );
  XOR U21241 ( .A(n21852), .B(n21853), .Z(n21846) );
  AND U21242 ( .A(n143), .B(n21845), .Z(n21853) );
  XNOR U21243 ( .A(n21843), .B(n21852), .Z(n21845) );
  XNOR U21244 ( .A(n21854), .B(n21855), .Z(n21843) );
  AND U21245 ( .A(n147), .B(n21856), .Z(n21855) );
  XOR U21246 ( .A(p_input[76]), .B(n21854), .Z(n21856) );
  XNOR U21247 ( .A(n21857), .B(n21858), .Z(n21854) );
  AND U21248 ( .A(n151), .B(n21859), .Z(n21858) );
  XOR U21249 ( .A(n21860), .B(n21861), .Z(n21852) );
  AND U21250 ( .A(n155), .B(n21851), .Z(n21861) );
  XNOR U21251 ( .A(n21862), .B(n21849), .Z(n21851) );
  XOR U21252 ( .A(n21863), .B(n21864), .Z(n21849) );
  AND U21253 ( .A(n178), .B(n21865), .Z(n21864) );
  IV U21254 ( .A(n21860), .Z(n21862) );
  XOR U21255 ( .A(n21866), .B(n21867), .Z(n21860) );
  AND U21256 ( .A(n162), .B(n21859), .Z(n21867) );
  XNOR U21257 ( .A(n21857), .B(n21866), .Z(n21859) );
  XNOR U21258 ( .A(n21868), .B(n21869), .Z(n21857) );
  AND U21259 ( .A(n166), .B(n21870), .Z(n21869) );
  XOR U21260 ( .A(p_input[92]), .B(n21868), .Z(n21870) );
  XNOR U21261 ( .A(n21871), .B(n21872), .Z(n21868) );
  AND U21262 ( .A(n170), .B(n21873), .Z(n21872) );
  XOR U21263 ( .A(n21874), .B(n21875), .Z(n21866) );
  AND U21264 ( .A(n174), .B(n21865), .Z(n21875) );
  XNOR U21265 ( .A(n21876), .B(n21863), .Z(n21865) );
  XOR U21266 ( .A(n21877), .B(n21878), .Z(n21863) );
  AND U21267 ( .A(n197), .B(n21879), .Z(n21878) );
  IV U21268 ( .A(n21874), .Z(n21876) );
  XOR U21269 ( .A(n21880), .B(n21881), .Z(n21874) );
  AND U21270 ( .A(n181), .B(n21873), .Z(n21881) );
  XNOR U21271 ( .A(n21871), .B(n21880), .Z(n21873) );
  XNOR U21272 ( .A(n21882), .B(n21883), .Z(n21871) );
  AND U21273 ( .A(n185), .B(n21884), .Z(n21883) );
  XOR U21274 ( .A(p_input[108]), .B(n21882), .Z(n21884) );
  XNOR U21275 ( .A(n21885), .B(n21886), .Z(n21882) );
  AND U21276 ( .A(n189), .B(n21887), .Z(n21886) );
  XOR U21277 ( .A(n21888), .B(n21889), .Z(n21880) );
  AND U21278 ( .A(n193), .B(n21879), .Z(n21889) );
  XNOR U21279 ( .A(n21890), .B(n21877), .Z(n21879) );
  XOR U21280 ( .A(n21891), .B(n21892), .Z(n21877) );
  AND U21281 ( .A(n216), .B(n21893), .Z(n21892) );
  IV U21282 ( .A(n21888), .Z(n21890) );
  XOR U21283 ( .A(n21894), .B(n21895), .Z(n21888) );
  AND U21284 ( .A(n200), .B(n21887), .Z(n21895) );
  XNOR U21285 ( .A(n21885), .B(n21894), .Z(n21887) );
  XNOR U21286 ( .A(n21896), .B(n21897), .Z(n21885) );
  AND U21287 ( .A(n204), .B(n21898), .Z(n21897) );
  XOR U21288 ( .A(p_input[124]), .B(n21896), .Z(n21898) );
  XNOR U21289 ( .A(n21899), .B(n21900), .Z(n21896) );
  AND U21290 ( .A(n208), .B(n21901), .Z(n21900) );
  XOR U21291 ( .A(n21902), .B(n21903), .Z(n21894) );
  AND U21292 ( .A(n212), .B(n21893), .Z(n21903) );
  XNOR U21293 ( .A(n21904), .B(n21891), .Z(n21893) );
  XOR U21294 ( .A(n21905), .B(n21906), .Z(n21891) );
  AND U21295 ( .A(n235), .B(n21907), .Z(n21906) );
  IV U21296 ( .A(n21902), .Z(n21904) );
  XOR U21297 ( .A(n21908), .B(n21909), .Z(n21902) );
  AND U21298 ( .A(n219), .B(n21901), .Z(n21909) );
  XNOR U21299 ( .A(n21899), .B(n21908), .Z(n21901) );
  XNOR U21300 ( .A(n21910), .B(n21911), .Z(n21899) );
  AND U21301 ( .A(n223), .B(n21912), .Z(n21911) );
  XOR U21302 ( .A(p_input[140]), .B(n21910), .Z(n21912) );
  XNOR U21303 ( .A(n21913), .B(n21914), .Z(n21910) );
  AND U21304 ( .A(n227), .B(n21915), .Z(n21914) );
  XOR U21305 ( .A(n21916), .B(n21917), .Z(n21908) );
  AND U21306 ( .A(n231), .B(n21907), .Z(n21917) );
  XNOR U21307 ( .A(n21918), .B(n21905), .Z(n21907) );
  XOR U21308 ( .A(n21919), .B(n21920), .Z(n21905) );
  AND U21309 ( .A(n254), .B(n21921), .Z(n21920) );
  IV U21310 ( .A(n21916), .Z(n21918) );
  XOR U21311 ( .A(n21922), .B(n21923), .Z(n21916) );
  AND U21312 ( .A(n238), .B(n21915), .Z(n21923) );
  XNOR U21313 ( .A(n21913), .B(n21922), .Z(n21915) );
  XNOR U21314 ( .A(n21924), .B(n21925), .Z(n21913) );
  AND U21315 ( .A(n242), .B(n21926), .Z(n21925) );
  XOR U21316 ( .A(p_input[156]), .B(n21924), .Z(n21926) );
  XNOR U21317 ( .A(n21927), .B(n21928), .Z(n21924) );
  AND U21318 ( .A(n246), .B(n21929), .Z(n21928) );
  XOR U21319 ( .A(n21930), .B(n21931), .Z(n21922) );
  AND U21320 ( .A(n250), .B(n21921), .Z(n21931) );
  XNOR U21321 ( .A(n21932), .B(n21919), .Z(n21921) );
  XOR U21322 ( .A(n21933), .B(n21934), .Z(n21919) );
  AND U21323 ( .A(n273), .B(n21935), .Z(n21934) );
  IV U21324 ( .A(n21930), .Z(n21932) );
  XOR U21325 ( .A(n21936), .B(n21937), .Z(n21930) );
  AND U21326 ( .A(n257), .B(n21929), .Z(n21937) );
  XNOR U21327 ( .A(n21927), .B(n21936), .Z(n21929) );
  XNOR U21328 ( .A(n21938), .B(n21939), .Z(n21927) );
  AND U21329 ( .A(n261), .B(n21940), .Z(n21939) );
  XOR U21330 ( .A(p_input[172]), .B(n21938), .Z(n21940) );
  XNOR U21331 ( .A(n21941), .B(n21942), .Z(n21938) );
  AND U21332 ( .A(n265), .B(n21943), .Z(n21942) );
  XOR U21333 ( .A(n21944), .B(n21945), .Z(n21936) );
  AND U21334 ( .A(n269), .B(n21935), .Z(n21945) );
  XNOR U21335 ( .A(n21946), .B(n21933), .Z(n21935) );
  XOR U21336 ( .A(n21947), .B(n21948), .Z(n21933) );
  AND U21337 ( .A(n292), .B(n21949), .Z(n21948) );
  IV U21338 ( .A(n21944), .Z(n21946) );
  XOR U21339 ( .A(n21950), .B(n21951), .Z(n21944) );
  AND U21340 ( .A(n276), .B(n21943), .Z(n21951) );
  XNOR U21341 ( .A(n21941), .B(n21950), .Z(n21943) );
  XNOR U21342 ( .A(n21952), .B(n21953), .Z(n21941) );
  AND U21343 ( .A(n280), .B(n21954), .Z(n21953) );
  XOR U21344 ( .A(p_input[188]), .B(n21952), .Z(n21954) );
  XNOR U21345 ( .A(n21955), .B(n21956), .Z(n21952) );
  AND U21346 ( .A(n284), .B(n21957), .Z(n21956) );
  XOR U21347 ( .A(n21958), .B(n21959), .Z(n21950) );
  AND U21348 ( .A(n288), .B(n21949), .Z(n21959) );
  XNOR U21349 ( .A(n21960), .B(n21947), .Z(n21949) );
  XOR U21350 ( .A(n21961), .B(n21962), .Z(n21947) );
  AND U21351 ( .A(n311), .B(n21963), .Z(n21962) );
  IV U21352 ( .A(n21958), .Z(n21960) );
  XOR U21353 ( .A(n21964), .B(n21965), .Z(n21958) );
  AND U21354 ( .A(n295), .B(n21957), .Z(n21965) );
  XNOR U21355 ( .A(n21955), .B(n21964), .Z(n21957) );
  XNOR U21356 ( .A(n21966), .B(n21967), .Z(n21955) );
  AND U21357 ( .A(n299), .B(n21968), .Z(n21967) );
  XOR U21358 ( .A(p_input[204]), .B(n21966), .Z(n21968) );
  XNOR U21359 ( .A(n21969), .B(n21970), .Z(n21966) );
  AND U21360 ( .A(n303), .B(n21971), .Z(n21970) );
  XOR U21361 ( .A(n21972), .B(n21973), .Z(n21964) );
  AND U21362 ( .A(n307), .B(n21963), .Z(n21973) );
  XNOR U21363 ( .A(n21974), .B(n21961), .Z(n21963) );
  XOR U21364 ( .A(n21975), .B(n21976), .Z(n21961) );
  AND U21365 ( .A(n330), .B(n21977), .Z(n21976) );
  IV U21366 ( .A(n21972), .Z(n21974) );
  XOR U21367 ( .A(n21978), .B(n21979), .Z(n21972) );
  AND U21368 ( .A(n314), .B(n21971), .Z(n21979) );
  XNOR U21369 ( .A(n21969), .B(n21978), .Z(n21971) );
  XNOR U21370 ( .A(n21980), .B(n21981), .Z(n21969) );
  AND U21371 ( .A(n318), .B(n21982), .Z(n21981) );
  XOR U21372 ( .A(p_input[220]), .B(n21980), .Z(n21982) );
  XNOR U21373 ( .A(n21983), .B(n21984), .Z(n21980) );
  AND U21374 ( .A(n322), .B(n21985), .Z(n21984) );
  XOR U21375 ( .A(n21986), .B(n21987), .Z(n21978) );
  AND U21376 ( .A(n326), .B(n21977), .Z(n21987) );
  XNOR U21377 ( .A(n21988), .B(n21975), .Z(n21977) );
  XOR U21378 ( .A(n21989), .B(n21990), .Z(n21975) );
  AND U21379 ( .A(n349), .B(n21991), .Z(n21990) );
  IV U21380 ( .A(n21986), .Z(n21988) );
  XOR U21381 ( .A(n21992), .B(n21993), .Z(n21986) );
  AND U21382 ( .A(n333), .B(n21985), .Z(n21993) );
  XNOR U21383 ( .A(n21983), .B(n21992), .Z(n21985) );
  XNOR U21384 ( .A(n21994), .B(n21995), .Z(n21983) );
  AND U21385 ( .A(n337), .B(n21996), .Z(n21995) );
  XOR U21386 ( .A(p_input[236]), .B(n21994), .Z(n21996) );
  XNOR U21387 ( .A(n21997), .B(n21998), .Z(n21994) );
  AND U21388 ( .A(n341), .B(n21999), .Z(n21998) );
  XOR U21389 ( .A(n22000), .B(n22001), .Z(n21992) );
  AND U21390 ( .A(n345), .B(n21991), .Z(n22001) );
  XNOR U21391 ( .A(n22002), .B(n21989), .Z(n21991) );
  XOR U21392 ( .A(n22003), .B(n22004), .Z(n21989) );
  AND U21393 ( .A(n368), .B(n22005), .Z(n22004) );
  IV U21394 ( .A(n22000), .Z(n22002) );
  XOR U21395 ( .A(n22006), .B(n22007), .Z(n22000) );
  AND U21396 ( .A(n352), .B(n21999), .Z(n22007) );
  XNOR U21397 ( .A(n21997), .B(n22006), .Z(n21999) );
  XNOR U21398 ( .A(n22008), .B(n22009), .Z(n21997) );
  AND U21399 ( .A(n356), .B(n22010), .Z(n22009) );
  XOR U21400 ( .A(p_input[252]), .B(n22008), .Z(n22010) );
  XNOR U21401 ( .A(n22011), .B(n22012), .Z(n22008) );
  AND U21402 ( .A(n360), .B(n22013), .Z(n22012) );
  XOR U21403 ( .A(n22014), .B(n22015), .Z(n22006) );
  AND U21404 ( .A(n364), .B(n22005), .Z(n22015) );
  XNOR U21405 ( .A(n22016), .B(n22003), .Z(n22005) );
  XOR U21406 ( .A(n22017), .B(n22018), .Z(n22003) );
  AND U21407 ( .A(n387), .B(n22019), .Z(n22018) );
  IV U21408 ( .A(n22014), .Z(n22016) );
  XOR U21409 ( .A(n22020), .B(n22021), .Z(n22014) );
  AND U21410 ( .A(n371), .B(n22013), .Z(n22021) );
  XNOR U21411 ( .A(n22011), .B(n22020), .Z(n22013) );
  XNOR U21412 ( .A(n22022), .B(n22023), .Z(n22011) );
  AND U21413 ( .A(n375), .B(n22024), .Z(n22023) );
  XOR U21414 ( .A(p_input[268]), .B(n22022), .Z(n22024) );
  XNOR U21415 ( .A(n22025), .B(n22026), .Z(n22022) );
  AND U21416 ( .A(n379), .B(n22027), .Z(n22026) );
  XOR U21417 ( .A(n22028), .B(n22029), .Z(n22020) );
  AND U21418 ( .A(n383), .B(n22019), .Z(n22029) );
  XNOR U21419 ( .A(n22030), .B(n22017), .Z(n22019) );
  XOR U21420 ( .A(n22031), .B(n22032), .Z(n22017) );
  AND U21421 ( .A(n406), .B(n22033), .Z(n22032) );
  IV U21422 ( .A(n22028), .Z(n22030) );
  XOR U21423 ( .A(n22034), .B(n22035), .Z(n22028) );
  AND U21424 ( .A(n390), .B(n22027), .Z(n22035) );
  XNOR U21425 ( .A(n22025), .B(n22034), .Z(n22027) );
  XNOR U21426 ( .A(n22036), .B(n22037), .Z(n22025) );
  AND U21427 ( .A(n394), .B(n22038), .Z(n22037) );
  XOR U21428 ( .A(p_input[284]), .B(n22036), .Z(n22038) );
  XNOR U21429 ( .A(n22039), .B(n22040), .Z(n22036) );
  AND U21430 ( .A(n398), .B(n22041), .Z(n22040) );
  XOR U21431 ( .A(n22042), .B(n22043), .Z(n22034) );
  AND U21432 ( .A(n402), .B(n22033), .Z(n22043) );
  XNOR U21433 ( .A(n22044), .B(n22031), .Z(n22033) );
  XOR U21434 ( .A(n22045), .B(n22046), .Z(n22031) );
  AND U21435 ( .A(n425), .B(n22047), .Z(n22046) );
  IV U21436 ( .A(n22042), .Z(n22044) );
  XOR U21437 ( .A(n22048), .B(n22049), .Z(n22042) );
  AND U21438 ( .A(n409), .B(n22041), .Z(n22049) );
  XNOR U21439 ( .A(n22039), .B(n22048), .Z(n22041) );
  XNOR U21440 ( .A(n22050), .B(n22051), .Z(n22039) );
  AND U21441 ( .A(n413), .B(n22052), .Z(n22051) );
  XOR U21442 ( .A(p_input[300]), .B(n22050), .Z(n22052) );
  XNOR U21443 ( .A(n22053), .B(n22054), .Z(n22050) );
  AND U21444 ( .A(n417), .B(n22055), .Z(n22054) );
  XOR U21445 ( .A(n22056), .B(n22057), .Z(n22048) );
  AND U21446 ( .A(n421), .B(n22047), .Z(n22057) );
  XNOR U21447 ( .A(n22058), .B(n22045), .Z(n22047) );
  XOR U21448 ( .A(n22059), .B(n22060), .Z(n22045) );
  AND U21449 ( .A(n444), .B(n22061), .Z(n22060) );
  IV U21450 ( .A(n22056), .Z(n22058) );
  XOR U21451 ( .A(n22062), .B(n22063), .Z(n22056) );
  AND U21452 ( .A(n428), .B(n22055), .Z(n22063) );
  XNOR U21453 ( .A(n22053), .B(n22062), .Z(n22055) );
  XNOR U21454 ( .A(n22064), .B(n22065), .Z(n22053) );
  AND U21455 ( .A(n432), .B(n22066), .Z(n22065) );
  XOR U21456 ( .A(p_input[316]), .B(n22064), .Z(n22066) );
  XNOR U21457 ( .A(n22067), .B(n22068), .Z(n22064) );
  AND U21458 ( .A(n436), .B(n22069), .Z(n22068) );
  XOR U21459 ( .A(n22070), .B(n22071), .Z(n22062) );
  AND U21460 ( .A(n440), .B(n22061), .Z(n22071) );
  XNOR U21461 ( .A(n22072), .B(n22059), .Z(n22061) );
  XOR U21462 ( .A(n22073), .B(n22074), .Z(n22059) );
  AND U21463 ( .A(n463), .B(n22075), .Z(n22074) );
  IV U21464 ( .A(n22070), .Z(n22072) );
  XOR U21465 ( .A(n22076), .B(n22077), .Z(n22070) );
  AND U21466 ( .A(n447), .B(n22069), .Z(n22077) );
  XNOR U21467 ( .A(n22067), .B(n22076), .Z(n22069) );
  XNOR U21468 ( .A(n22078), .B(n22079), .Z(n22067) );
  AND U21469 ( .A(n451), .B(n22080), .Z(n22079) );
  XOR U21470 ( .A(p_input[332]), .B(n22078), .Z(n22080) );
  XNOR U21471 ( .A(n22081), .B(n22082), .Z(n22078) );
  AND U21472 ( .A(n455), .B(n22083), .Z(n22082) );
  XOR U21473 ( .A(n22084), .B(n22085), .Z(n22076) );
  AND U21474 ( .A(n459), .B(n22075), .Z(n22085) );
  XNOR U21475 ( .A(n22086), .B(n22073), .Z(n22075) );
  XOR U21476 ( .A(n22087), .B(n22088), .Z(n22073) );
  AND U21477 ( .A(n482), .B(n22089), .Z(n22088) );
  IV U21478 ( .A(n22084), .Z(n22086) );
  XOR U21479 ( .A(n22090), .B(n22091), .Z(n22084) );
  AND U21480 ( .A(n466), .B(n22083), .Z(n22091) );
  XNOR U21481 ( .A(n22081), .B(n22090), .Z(n22083) );
  XNOR U21482 ( .A(n22092), .B(n22093), .Z(n22081) );
  AND U21483 ( .A(n470), .B(n22094), .Z(n22093) );
  XOR U21484 ( .A(p_input[348]), .B(n22092), .Z(n22094) );
  XNOR U21485 ( .A(n22095), .B(n22096), .Z(n22092) );
  AND U21486 ( .A(n474), .B(n22097), .Z(n22096) );
  XOR U21487 ( .A(n22098), .B(n22099), .Z(n22090) );
  AND U21488 ( .A(n478), .B(n22089), .Z(n22099) );
  XNOR U21489 ( .A(n22100), .B(n22087), .Z(n22089) );
  XOR U21490 ( .A(n22101), .B(n22102), .Z(n22087) );
  AND U21491 ( .A(n501), .B(n22103), .Z(n22102) );
  IV U21492 ( .A(n22098), .Z(n22100) );
  XOR U21493 ( .A(n22104), .B(n22105), .Z(n22098) );
  AND U21494 ( .A(n485), .B(n22097), .Z(n22105) );
  XNOR U21495 ( .A(n22095), .B(n22104), .Z(n22097) );
  XNOR U21496 ( .A(n22106), .B(n22107), .Z(n22095) );
  AND U21497 ( .A(n489), .B(n22108), .Z(n22107) );
  XOR U21498 ( .A(p_input[364]), .B(n22106), .Z(n22108) );
  XNOR U21499 ( .A(n22109), .B(n22110), .Z(n22106) );
  AND U21500 ( .A(n493), .B(n22111), .Z(n22110) );
  XOR U21501 ( .A(n22112), .B(n22113), .Z(n22104) );
  AND U21502 ( .A(n497), .B(n22103), .Z(n22113) );
  XNOR U21503 ( .A(n22114), .B(n22101), .Z(n22103) );
  XOR U21504 ( .A(n22115), .B(n22116), .Z(n22101) );
  AND U21505 ( .A(n520), .B(n22117), .Z(n22116) );
  IV U21506 ( .A(n22112), .Z(n22114) );
  XOR U21507 ( .A(n22118), .B(n22119), .Z(n22112) );
  AND U21508 ( .A(n504), .B(n22111), .Z(n22119) );
  XNOR U21509 ( .A(n22109), .B(n22118), .Z(n22111) );
  XNOR U21510 ( .A(n22120), .B(n22121), .Z(n22109) );
  AND U21511 ( .A(n508), .B(n22122), .Z(n22121) );
  XOR U21512 ( .A(p_input[380]), .B(n22120), .Z(n22122) );
  XNOR U21513 ( .A(n22123), .B(n22124), .Z(n22120) );
  AND U21514 ( .A(n512), .B(n22125), .Z(n22124) );
  XOR U21515 ( .A(n22126), .B(n22127), .Z(n22118) );
  AND U21516 ( .A(n516), .B(n22117), .Z(n22127) );
  XNOR U21517 ( .A(n22128), .B(n22115), .Z(n22117) );
  XOR U21518 ( .A(n22129), .B(n22130), .Z(n22115) );
  AND U21519 ( .A(n539), .B(n22131), .Z(n22130) );
  IV U21520 ( .A(n22126), .Z(n22128) );
  XOR U21521 ( .A(n22132), .B(n22133), .Z(n22126) );
  AND U21522 ( .A(n523), .B(n22125), .Z(n22133) );
  XNOR U21523 ( .A(n22123), .B(n22132), .Z(n22125) );
  XNOR U21524 ( .A(n22134), .B(n22135), .Z(n22123) );
  AND U21525 ( .A(n527), .B(n22136), .Z(n22135) );
  XOR U21526 ( .A(p_input[396]), .B(n22134), .Z(n22136) );
  XNOR U21527 ( .A(n22137), .B(n22138), .Z(n22134) );
  AND U21528 ( .A(n531), .B(n22139), .Z(n22138) );
  XOR U21529 ( .A(n22140), .B(n22141), .Z(n22132) );
  AND U21530 ( .A(n535), .B(n22131), .Z(n22141) );
  XNOR U21531 ( .A(n22142), .B(n22129), .Z(n22131) );
  XOR U21532 ( .A(n22143), .B(n22144), .Z(n22129) );
  AND U21533 ( .A(n558), .B(n22145), .Z(n22144) );
  IV U21534 ( .A(n22140), .Z(n22142) );
  XOR U21535 ( .A(n22146), .B(n22147), .Z(n22140) );
  AND U21536 ( .A(n542), .B(n22139), .Z(n22147) );
  XNOR U21537 ( .A(n22137), .B(n22146), .Z(n22139) );
  XNOR U21538 ( .A(n22148), .B(n22149), .Z(n22137) );
  AND U21539 ( .A(n546), .B(n22150), .Z(n22149) );
  XOR U21540 ( .A(p_input[412]), .B(n22148), .Z(n22150) );
  XNOR U21541 ( .A(n22151), .B(n22152), .Z(n22148) );
  AND U21542 ( .A(n550), .B(n22153), .Z(n22152) );
  XOR U21543 ( .A(n22154), .B(n22155), .Z(n22146) );
  AND U21544 ( .A(n554), .B(n22145), .Z(n22155) );
  XNOR U21545 ( .A(n22156), .B(n22143), .Z(n22145) );
  XOR U21546 ( .A(n22157), .B(n22158), .Z(n22143) );
  AND U21547 ( .A(n577), .B(n22159), .Z(n22158) );
  IV U21548 ( .A(n22154), .Z(n22156) );
  XOR U21549 ( .A(n22160), .B(n22161), .Z(n22154) );
  AND U21550 ( .A(n561), .B(n22153), .Z(n22161) );
  XNOR U21551 ( .A(n22151), .B(n22160), .Z(n22153) );
  XNOR U21552 ( .A(n22162), .B(n22163), .Z(n22151) );
  AND U21553 ( .A(n565), .B(n22164), .Z(n22163) );
  XOR U21554 ( .A(p_input[428]), .B(n22162), .Z(n22164) );
  XNOR U21555 ( .A(n22165), .B(n22166), .Z(n22162) );
  AND U21556 ( .A(n569), .B(n22167), .Z(n22166) );
  XOR U21557 ( .A(n22168), .B(n22169), .Z(n22160) );
  AND U21558 ( .A(n573), .B(n22159), .Z(n22169) );
  XNOR U21559 ( .A(n22170), .B(n22157), .Z(n22159) );
  XOR U21560 ( .A(n22171), .B(n22172), .Z(n22157) );
  AND U21561 ( .A(n596), .B(n22173), .Z(n22172) );
  IV U21562 ( .A(n22168), .Z(n22170) );
  XOR U21563 ( .A(n22174), .B(n22175), .Z(n22168) );
  AND U21564 ( .A(n580), .B(n22167), .Z(n22175) );
  XNOR U21565 ( .A(n22165), .B(n22174), .Z(n22167) );
  XNOR U21566 ( .A(n22176), .B(n22177), .Z(n22165) );
  AND U21567 ( .A(n584), .B(n22178), .Z(n22177) );
  XOR U21568 ( .A(p_input[444]), .B(n22176), .Z(n22178) );
  XNOR U21569 ( .A(n22179), .B(n22180), .Z(n22176) );
  AND U21570 ( .A(n588), .B(n22181), .Z(n22180) );
  XOR U21571 ( .A(n22182), .B(n22183), .Z(n22174) );
  AND U21572 ( .A(n592), .B(n22173), .Z(n22183) );
  XNOR U21573 ( .A(n22184), .B(n22171), .Z(n22173) );
  XOR U21574 ( .A(n22185), .B(n22186), .Z(n22171) );
  AND U21575 ( .A(n615), .B(n22187), .Z(n22186) );
  IV U21576 ( .A(n22182), .Z(n22184) );
  XOR U21577 ( .A(n22188), .B(n22189), .Z(n22182) );
  AND U21578 ( .A(n599), .B(n22181), .Z(n22189) );
  XNOR U21579 ( .A(n22179), .B(n22188), .Z(n22181) );
  XNOR U21580 ( .A(n22190), .B(n22191), .Z(n22179) );
  AND U21581 ( .A(n603), .B(n22192), .Z(n22191) );
  XOR U21582 ( .A(p_input[460]), .B(n22190), .Z(n22192) );
  XNOR U21583 ( .A(n22193), .B(n22194), .Z(n22190) );
  AND U21584 ( .A(n607), .B(n22195), .Z(n22194) );
  XOR U21585 ( .A(n22196), .B(n22197), .Z(n22188) );
  AND U21586 ( .A(n611), .B(n22187), .Z(n22197) );
  XNOR U21587 ( .A(n22198), .B(n22185), .Z(n22187) );
  XOR U21588 ( .A(n22199), .B(n22200), .Z(n22185) );
  AND U21589 ( .A(n634), .B(n22201), .Z(n22200) );
  IV U21590 ( .A(n22196), .Z(n22198) );
  XOR U21591 ( .A(n22202), .B(n22203), .Z(n22196) );
  AND U21592 ( .A(n618), .B(n22195), .Z(n22203) );
  XNOR U21593 ( .A(n22193), .B(n22202), .Z(n22195) );
  XNOR U21594 ( .A(n22204), .B(n22205), .Z(n22193) );
  AND U21595 ( .A(n622), .B(n22206), .Z(n22205) );
  XOR U21596 ( .A(p_input[476]), .B(n22204), .Z(n22206) );
  XNOR U21597 ( .A(n22207), .B(n22208), .Z(n22204) );
  AND U21598 ( .A(n626), .B(n22209), .Z(n22208) );
  XOR U21599 ( .A(n22210), .B(n22211), .Z(n22202) );
  AND U21600 ( .A(n630), .B(n22201), .Z(n22211) );
  XNOR U21601 ( .A(n22212), .B(n22199), .Z(n22201) );
  XOR U21602 ( .A(n22213), .B(n22214), .Z(n22199) );
  AND U21603 ( .A(n653), .B(n22215), .Z(n22214) );
  IV U21604 ( .A(n22210), .Z(n22212) );
  XOR U21605 ( .A(n22216), .B(n22217), .Z(n22210) );
  AND U21606 ( .A(n637), .B(n22209), .Z(n22217) );
  XNOR U21607 ( .A(n22207), .B(n22216), .Z(n22209) );
  XNOR U21608 ( .A(n22218), .B(n22219), .Z(n22207) );
  AND U21609 ( .A(n641), .B(n22220), .Z(n22219) );
  XOR U21610 ( .A(p_input[492]), .B(n22218), .Z(n22220) );
  XNOR U21611 ( .A(n22221), .B(n22222), .Z(n22218) );
  AND U21612 ( .A(n645), .B(n22223), .Z(n22222) );
  XOR U21613 ( .A(n22224), .B(n22225), .Z(n22216) );
  AND U21614 ( .A(n649), .B(n22215), .Z(n22225) );
  XNOR U21615 ( .A(n22226), .B(n22213), .Z(n22215) );
  XOR U21616 ( .A(n22227), .B(n22228), .Z(n22213) );
  AND U21617 ( .A(n672), .B(n22229), .Z(n22228) );
  IV U21618 ( .A(n22224), .Z(n22226) );
  XOR U21619 ( .A(n22230), .B(n22231), .Z(n22224) );
  AND U21620 ( .A(n656), .B(n22223), .Z(n22231) );
  XNOR U21621 ( .A(n22221), .B(n22230), .Z(n22223) );
  XNOR U21622 ( .A(n22232), .B(n22233), .Z(n22221) );
  AND U21623 ( .A(n660), .B(n22234), .Z(n22233) );
  XOR U21624 ( .A(p_input[508]), .B(n22232), .Z(n22234) );
  XNOR U21625 ( .A(n22235), .B(n22236), .Z(n22232) );
  AND U21626 ( .A(n664), .B(n22237), .Z(n22236) );
  XOR U21627 ( .A(n22238), .B(n22239), .Z(n22230) );
  AND U21628 ( .A(n668), .B(n22229), .Z(n22239) );
  XNOR U21629 ( .A(n22240), .B(n22227), .Z(n22229) );
  XOR U21630 ( .A(n22241), .B(n22242), .Z(n22227) );
  AND U21631 ( .A(n691), .B(n22243), .Z(n22242) );
  IV U21632 ( .A(n22238), .Z(n22240) );
  XOR U21633 ( .A(n22244), .B(n22245), .Z(n22238) );
  AND U21634 ( .A(n675), .B(n22237), .Z(n22245) );
  XNOR U21635 ( .A(n22235), .B(n22244), .Z(n22237) );
  XNOR U21636 ( .A(n22246), .B(n22247), .Z(n22235) );
  AND U21637 ( .A(n679), .B(n22248), .Z(n22247) );
  XOR U21638 ( .A(p_input[524]), .B(n22246), .Z(n22248) );
  XNOR U21639 ( .A(n22249), .B(n22250), .Z(n22246) );
  AND U21640 ( .A(n683), .B(n22251), .Z(n22250) );
  XOR U21641 ( .A(n22252), .B(n22253), .Z(n22244) );
  AND U21642 ( .A(n687), .B(n22243), .Z(n22253) );
  XNOR U21643 ( .A(n22254), .B(n22241), .Z(n22243) );
  XOR U21644 ( .A(n22255), .B(n22256), .Z(n22241) );
  AND U21645 ( .A(n710), .B(n22257), .Z(n22256) );
  IV U21646 ( .A(n22252), .Z(n22254) );
  XOR U21647 ( .A(n22258), .B(n22259), .Z(n22252) );
  AND U21648 ( .A(n694), .B(n22251), .Z(n22259) );
  XNOR U21649 ( .A(n22249), .B(n22258), .Z(n22251) );
  XNOR U21650 ( .A(n22260), .B(n22261), .Z(n22249) );
  AND U21651 ( .A(n698), .B(n22262), .Z(n22261) );
  XOR U21652 ( .A(p_input[540]), .B(n22260), .Z(n22262) );
  XNOR U21653 ( .A(n22263), .B(n22264), .Z(n22260) );
  AND U21654 ( .A(n702), .B(n22265), .Z(n22264) );
  XOR U21655 ( .A(n22266), .B(n22267), .Z(n22258) );
  AND U21656 ( .A(n706), .B(n22257), .Z(n22267) );
  XNOR U21657 ( .A(n22268), .B(n22255), .Z(n22257) );
  XOR U21658 ( .A(n22269), .B(n22270), .Z(n22255) );
  AND U21659 ( .A(n729), .B(n22271), .Z(n22270) );
  IV U21660 ( .A(n22266), .Z(n22268) );
  XOR U21661 ( .A(n22272), .B(n22273), .Z(n22266) );
  AND U21662 ( .A(n713), .B(n22265), .Z(n22273) );
  XNOR U21663 ( .A(n22263), .B(n22272), .Z(n22265) );
  XNOR U21664 ( .A(n22274), .B(n22275), .Z(n22263) );
  AND U21665 ( .A(n717), .B(n22276), .Z(n22275) );
  XOR U21666 ( .A(p_input[556]), .B(n22274), .Z(n22276) );
  XNOR U21667 ( .A(n22277), .B(n22278), .Z(n22274) );
  AND U21668 ( .A(n721), .B(n22279), .Z(n22278) );
  XOR U21669 ( .A(n22280), .B(n22281), .Z(n22272) );
  AND U21670 ( .A(n725), .B(n22271), .Z(n22281) );
  XNOR U21671 ( .A(n22282), .B(n22269), .Z(n22271) );
  XOR U21672 ( .A(n22283), .B(n22284), .Z(n22269) );
  AND U21673 ( .A(n748), .B(n22285), .Z(n22284) );
  IV U21674 ( .A(n22280), .Z(n22282) );
  XOR U21675 ( .A(n22286), .B(n22287), .Z(n22280) );
  AND U21676 ( .A(n732), .B(n22279), .Z(n22287) );
  XNOR U21677 ( .A(n22277), .B(n22286), .Z(n22279) );
  XNOR U21678 ( .A(n22288), .B(n22289), .Z(n22277) );
  AND U21679 ( .A(n736), .B(n22290), .Z(n22289) );
  XOR U21680 ( .A(p_input[572]), .B(n22288), .Z(n22290) );
  XNOR U21681 ( .A(n22291), .B(n22292), .Z(n22288) );
  AND U21682 ( .A(n740), .B(n22293), .Z(n22292) );
  XOR U21683 ( .A(n22294), .B(n22295), .Z(n22286) );
  AND U21684 ( .A(n744), .B(n22285), .Z(n22295) );
  XNOR U21685 ( .A(n22296), .B(n22283), .Z(n22285) );
  XOR U21686 ( .A(n22297), .B(n22298), .Z(n22283) );
  AND U21687 ( .A(n767), .B(n22299), .Z(n22298) );
  IV U21688 ( .A(n22294), .Z(n22296) );
  XOR U21689 ( .A(n22300), .B(n22301), .Z(n22294) );
  AND U21690 ( .A(n751), .B(n22293), .Z(n22301) );
  XNOR U21691 ( .A(n22291), .B(n22300), .Z(n22293) );
  XNOR U21692 ( .A(n22302), .B(n22303), .Z(n22291) );
  AND U21693 ( .A(n755), .B(n22304), .Z(n22303) );
  XOR U21694 ( .A(p_input[588]), .B(n22302), .Z(n22304) );
  XNOR U21695 ( .A(n22305), .B(n22306), .Z(n22302) );
  AND U21696 ( .A(n759), .B(n22307), .Z(n22306) );
  XOR U21697 ( .A(n22308), .B(n22309), .Z(n22300) );
  AND U21698 ( .A(n763), .B(n22299), .Z(n22309) );
  XNOR U21699 ( .A(n22310), .B(n22297), .Z(n22299) );
  XOR U21700 ( .A(n22311), .B(n22312), .Z(n22297) );
  AND U21701 ( .A(n786), .B(n22313), .Z(n22312) );
  IV U21702 ( .A(n22308), .Z(n22310) );
  XOR U21703 ( .A(n22314), .B(n22315), .Z(n22308) );
  AND U21704 ( .A(n770), .B(n22307), .Z(n22315) );
  XNOR U21705 ( .A(n22305), .B(n22314), .Z(n22307) );
  XNOR U21706 ( .A(n22316), .B(n22317), .Z(n22305) );
  AND U21707 ( .A(n774), .B(n22318), .Z(n22317) );
  XOR U21708 ( .A(p_input[604]), .B(n22316), .Z(n22318) );
  XNOR U21709 ( .A(n22319), .B(n22320), .Z(n22316) );
  AND U21710 ( .A(n778), .B(n22321), .Z(n22320) );
  XOR U21711 ( .A(n22322), .B(n22323), .Z(n22314) );
  AND U21712 ( .A(n782), .B(n22313), .Z(n22323) );
  XNOR U21713 ( .A(n22324), .B(n22311), .Z(n22313) );
  XOR U21714 ( .A(n22325), .B(n22326), .Z(n22311) );
  AND U21715 ( .A(n805), .B(n22327), .Z(n22326) );
  IV U21716 ( .A(n22322), .Z(n22324) );
  XOR U21717 ( .A(n22328), .B(n22329), .Z(n22322) );
  AND U21718 ( .A(n789), .B(n22321), .Z(n22329) );
  XNOR U21719 ( .A(n22319), .B(n22328), .Z(n22321) );
  XNOR U21720 ( .A(n22330), .B(n22331), .Z(n22319) );
  AND U21721 ( .A(n793), .B(n22332), .Z(n22331) );
  XOR U21722 ( .A(p_input[620]), .B(n22330), .Z(n22332) );
  XNOR U21723 ( .A(n22333), .B(n22334), .Z(n22330) );
  AND U21724 ( .A(n797), .B(n22335), .Z(n22334) );
  XOR U21725 ( .A(n22336), .B(n22337), .Z(n22328) );
  AND U21726 ( .A(n801), .B(n22327), .Z(n22337) );
  XNOR U21727 ( .A(n22338), .B(n22325), .Z(n22327) );
  XOR U21728 ( .A(n22339), .B(n22340), .Z(n22325) );
  AND U21729 ( .A(n824), .B(n22341), .Z(n22340) );
  IV U21730 ( .A(n22336), .Z(n22338) );
  XOR U21731 ( .A(n22342), .B(n22343), .Z(n22336) );
  AND U21732 ( .A(n808), .B(n22335), .Z(n22343) );
  XNOR U21733 ( .A(n22333), .B(n22342), .Z(n22335) );
  XNOR U21734 ( .A(n22344), .B(n22345), .Z(n22333) );
  AND U21735 ( .A(n812), .B(n22346), .Z(n22345) );
  XOR U21736 ( .A(p_input[636]), .B(n22344), .Z(n22346) );
  XNOR U21737 ( .A(n22347), .B(n22348), .Z(n22344) );
  AND U21738 ( .A(n816), .B(n22349), .Z(n22348) );
  XOR U21739 ( .A(n22350), .B(n22351), .Z(n22342) );
  AND U21740 ( .A(n820), .B(n22341), .Z(n22351) );
  XNOR U21741 ( .A(n22352), .B(n22339), .Z(n22341) );
  XOR U21742 ( .A(n22353), .B(n22354), .Z(n22339) );
  AND U21743 ( .A(n843), .B(n22355), .Z(n22354) );
  IV U21744 ( .A(n22350), .Z(n22352) );
  XOR U21745 ( .A(n22356), .B(n22357), .Z(n22350) );
  AND U21746 ( .A(n827), .B(n22349), .Z(n22357) );
  XNOR U21747 ( .A(n22347), .B(n22356), .Z(n22349) );
  XNOR U21748 ( .A(n22358), .B(n22359), .Z(n22347) );
  AND U21749 ( .A(n831), .B(n22360), .Z(n22359) );
  XOR U21750 ( .A(p_input[652]), .B(n22358), .Z(n22360) );
  XNOR U21751 ( .A(n22361), .B(n22362), .Z(n22358) );
  AND U21752 ( .A(n835), .B(n22363), .Z(n22362) );
  XOR U21753 ( .A(n22364), .B(n22365), .Z(n22356) );
  AND U21754 ( .A(n839), .B(n22355), .Z(n22365) );
  XNOR U21755 ( .A(n22366), .B(n22353), .Z(n22355) );
  XOR U21756 ( .A(n22367), .B(n22368), .Z(n22353) );
  AND U21757 ( .A(n862), .B(n22369), .Z(n22368) );
  IV U21758 ( .A(n22364), .Z(n22366) );
  XOR U21759 ( .A(n22370), .B(n22371), .Z(n22364) );
  AND U21760 ( .A(n846), .B(n22363), .Z(n22371) );
  XNOR U21761 ( .A(n22361), .B(n22370), .Z(n22363) );
  XNOR U21762 ( .A(n22372), .B(n22373), .Z(n22361) );
  AND U21763 ( .A(n850), .B(n22374), .Z(n22373) );
  XOR U21764 ( .A(p_input[668]), .B(n22372), .Z(n22374) );
  XNOR U21765 ( .A(n22375), .B(n22376), .Z(n22372) );
  AND U21766 ( .A(n854), .B(n22377), .Z(n22376) );
  XOR U21767 ( .A(n22378), .B(n22379), .Z(n22370) );
  AND U21768 ( .A(n858), .B(n22369), .Z(n22379) );
  XNOR U21769 ( .A(n22380), .B(n22367), .Z(n22369) );
  XOR U21770 ( .A(n22381), .B(n22382), .Z(n22367) );
  AND U21771 ( .A(n881), .B(n22383), .Z(n22382) );
  IV U21772 ( .A(n22378), .Z(n22380) );
  XOR U21773 ( .A(n22384), .B(n22385), .Z(n22378) );
  AND U21774 ( .A(n865), .B(n22377), .Z(n22385) );
  XNOR U21775 ( .A(n22375), .B(n22384), .Z(n22377) );
  XNOR U21776 ( .A(n22386), .B(n22387), .Z(n22375) );
  AND U21777 ( .A(n869), .B(n22388), .Z(n22387) );
  XOR U21778 ( .A(p_input[684]), .B(n22386), .Z(n22388) );
  XNOR U21779 ( .A(n22389), .B(n22390), .Z(n22386) );
  AND U21780 ( .A(n873), .B(n22391), .Z(n22390) );
  XOR U21781 ( .A(n22392), .B(n22393), .Z(n22384) );
  AND U21782 ( .A(n877), .B(n22383), .Z(n22393) );
  XNOR U21783 ( .A(n22394), .B(n22381), .Z(n22383) );
  XOR U21784 ( .A(n22395), .B(n22396), .Z(n22381) );
  AND U21785 ( .A(n900), .B(n22397), .Z(n22396) );
  IV U21786 ( .A(n22392), .Z(n22394) );
  XOR U21787 ( .A(n22398), .B(n22399), .Z(n22392) );
  AND U21788 ( .A(n884), .B(n22391), .Z(n22399) );
  XNOR U21789 ( .A(n22389), .B(n22398), .Z(n22391) );
  XNOR U21790 ( .A(n22400), .B(n22401), .Z(n22389) );
  AND U21791 ( .A(n888), .B(n22402), .Z(n22401) );
  XOR U21792 ( .A(p_input[700]), .B(n22400), .Z(n22402) );
  XNOR U21793 ( .A(n22403), .B(n22404), .Z(n22400) );
  AND U21794 ( .A(n892), .B(n22405), .Z(n22404) );
  XOR U21795 ( .A(n22406), .B(n22407), .Z(n22398) );
  AND U21796 ( .A(n896), .B(n22397), .Z(n22407) );
  XNOR U21797 ( .A(n22408), .B(n22395), .Z(n22397) );
  XOR U21798 ( .A(n22409), .B(n22410), .Z(n22395) );
  AND U21799 ( .A(n919), .B(n22411), .Z(n22410) );
  IV U21800 ( .A(n22406), .Z(n22408) );
  XOR U21801 ( .A(n22412), .B(n22413), .Z(n22406) );
  AND U21802 ( .A(n903), .B(n22405), .Z(n22413) );
  XNOR U21803 ( .A(n22403), .B(n22412), .Z(n22405) );
  XNOR U21804 ( .A(n22414), .B(n22415), .Z(n22403) );
  AND U21805 ( .A(n907), .B(n22416), .Z(n22415) );
  XOR U21806 ( .A(p_input[716]), .B(n22414), .Z(n22416) );
  XNOR U21807 ( .A(n22417), .B(n22418), .Z(n22414) );
  AND U21808 ( .A(n911), .B(n22419), .Z(n22418) );
  XOR U21809 ( .A(n22420), .B(n22421), .Z(n22412) );
  AND U21810 ( .A(n915), .B(n22411), .Z(n22421) );
  XNOR U21811 ( .A(n22422), .B(n22409), .Z(n22411) );
  XOR U21812 ( .A(n22423), .B(n22424), .Z(n22409) );
  AND U21813 ( .A(n938), .B(n22425), .Z(n22424) );
  IV U21814 ( .A(n22420), .Z(n22422) );
  XOR U21815 ( .A(n22426), .B(n22427), .Z(n22420) );
  AND U21816 ( .A(n922), .B(n22419), .Z(n22427) );
  XNOR U21817 ( .A(n22417), .B(n22426), .Z(n22419) );
  XNOR U21818 ( .A(n22428), .B(n22429), .Z(n22417) );
  AND U21819 ( .A(n926), .B(n22430), .Z(n22429) );
  XOR U21820 ( .A(p_input[732]), .B(n22428), .Z(n22430) );
  XNOR U21821 ( .A(n22431), .B(n22432), .Z(n22428) );
  AND U21822 ( .A(n930), .B(n22433), .Z(n22432) );
  XOR U21823 ( .A(n22434), .B(n22435), .Z(n22426) );
  AND U21824 ( .A(n934), .B(n22425), .Z(n22435) );
  XNOR U21825 ( .A(n22436), .B(n22423), .Z(n22425) );
  XOR U21826 ( .A(n22437), .B(n22438), .Z(n22423) );
  AND U21827 ( .A(n957), .B(n22439), .Z(n22438) );
  IV U21828 ( .A(n22434), .Z(n22436) );
  XOR U21829 ( .A(n22440), .B(n22441), .Z(n22434) );
  AND U21830 ( .A(n941), .B(n22433), .Z(n22441) );
  XNOR U21831 ( .A(n22431), .B(n22440), .Z(n22433) );
  XNOR U21832 ( .A(n22442), .B(n22443), .Z(n22431) );
  AND U21833 ( .A(n945), .B(n22444), .Z(n22443) );
  XOR U21834 ( .A(p_input[748]), .B(n22442), .Z(n22444) );
  XNOR U21835 ( .A(n22445), .B(n22446), .Z(n22442) );
  AND U21836 ( .A(n949), .B(n22447), .Z(n22446) );
  XOR U21837 ( .A(n22448), .B(n22449), .Z(n22440) );
  AND U21838 ( .A(n953), .B(n22439), .Z(n22449) );
  XNOR U21839 ( .A(n22450), .B(n22437), .Z(n22439) );
  XOR U21840 ( .A(n22451), .B(n22452), .Z(n22437) );
  AND U21841 ( .A(n976), .B(n22453), .Z(n22452) );
  IV U21842 ( .A(n22448), .Z(n22450) );
  XOR U21843 ( .A(n22454), .B(n22455), .Z(n22448) );
  AND U21844 ( .A(n960), .B(n22447), .Z(n22455) );
  XNOR U21845 ( .A(n22445), .B(n22454), .Z(n22447) );
  XNOR U21846 ( .A(n22456), .B(n22457), .Z(n22445) );
  AND U21847 ( .A(n964), .B(n22458), .Z(n22457) );
  XOR U21848 ( .A(p_input[764]), .B(n22456), .Z(n22458) );
  XNOR U21849 ( .A(n22459), .B(n22460), .Z(n22456) );
  AND U21850 ( .A(n968), .B(n22461), .Z(n22460) );
  XOR U21851 ( .A(n22462), .B(n22463), .Z(n22454) );
  AND U21852 ( .A(n972), .B(n22453), .Z(n22463) );
  XNOR U21853 ( .A(n22464), .B(n22451), .Z(n22453) );
  XOR U21854 ( .A(n22465), .B(n22466), .Z(n22451) );
  AND U21855 ( .A(n995), .B(n22467), .Z(n22466) );
  IV U21856 ( .A(n22462), .Z(n22464) );
  XOR U21857 ( .A(n22468), .B(n22469), .Z(n22462) );
  AND U21858 ( .A(n979), .B(n22461), .Z(n22469) );
  XNOR U21859 ( .A(n22459), .B(n22468), .Z(n22461) );
  XNOR U21860 ( .A(n22470), .B(n22471), .Z(n22459) );
  AND U21861 ( .A(n983), .B(n22472), .Z(n22471) );
  XOR U21862 ( .A(p_input[780]), .B(n22470), .Z(n22472) );
  XNOR U21863 ( .A(n22473), .B(n22474), .Z(n22470) );
  AND U21864 ( .A(n987), .B(n22475), .Z(n22474) );
  XOR U21865 ( .A(n22476), .B(n22477), .Z(n22468) );
  AND U21866 ( .A(n991), .B(n22467), .Z(n22477) );
  XNOR U21867 ( .A(n22478), .B(n22465), .Z(n22467) );
  XOR U21868 ( .A(n22479), .B(n22480), .Z(n22465) );
  AND U21869 ( .A(n1014), .B(n22481), .Z(n22480) );
  IV U21870 ( .A(n22476), .Z(n22478) );
  XOR U21871 ( .A(n22482), .B(n22483), .Z(n22476) );
  AND U21872 ( .A(n998), .B(n22475), .Z(n22483) );
  XNOR U21873 ( .A(n22473), .B(n22482), .Z(n22475) );
  XNOR U21874 ( .A(n22484), .B(n22485), .Z(n22473) );
  AND U21875 ( .A(n1002), .B(n22486), .Z(n22485) );
  XOR U21876 ( .A(p_input[796]), .B(n22484), .Z(n22486) );
  XNOR U21877 ( .A(n22487), .B(n22488), .Z(n22484) );
  AND U21878 ( .A(n1006), .B(n22489), .Z(n22488) );
  XOR U21879 ( .A(n22490), .B(n22491), .Z(n22482) );
  AND U21880 ( .A(n1010), .B(n22481), .Z(n22491) );
  XNOR U21881 ( .A(n22492), .B(n22479), .Z(n22481) );
  XOR U21882 ( .A(n22493), .B(n22494), .Z(n22479) );
  AND U21883 ( .A(n1033), .B(n22495), .Z(n22494) );
  IV U21884 ( .A(n22490), .Z(n22492) );
  XOR U21885 ( .A(n22496), .B(n22497), .Z(n22490) );
  AND U21886 ( .A(n1017), .B(n22489), .Z(n22497) );
  XNOR U21887 ( .A(n22487), .B(n22496), .Z(n22489) );
  XNOR U21888 ( .A(n22498), .B(n22499), .Z(n22487) );
  AND U21889 ( .A(n1021), .B(n22500), .Z(n22499) );
  XOR U21890 ( .A(p_input[812]), .B(n22498), .Z(n22500) );
  XNOR U21891 ( .A(n22501), .B(n22502), .Z(n22498) );
  AND U21892 ( .A(n1025), .B(n22503), .Z(n22502) );
  XOR U21893 ( .A(n22504), .B(n22505), .Z(n22496) );
  AND U21894 ( .A(n1029), .B(n22495), .Z(n22505) );
  XNOR U21895 ( .A(n22506), .B(n22493), .Z(n22495) );
  XOR U21896 ( .A(n22507), .B(n22508), .Z(n22493) );
  AND U21897 ( .A(n1052), .B(n22509), .Z(n22508) );
  IV U21898 ( .A(n22504), .Z(n22506) );
  XOR U21899 ( .A(n22510), .B(n22511), .Z(n22504) );
  AND U21900 ( .A(n1036), .B(n22503), .Z(n22511) );
  XNOR U21901 ( .A(n22501), .B(n22510), .Z(n22503) );
  XNOR U21902 ( .A(n22512), .B(n22513), .Z(n22501) );
  AND U21903 ( .A(n1040), .B(n22514), .Z(n22513) );
  XOR U21904 ( .A(p_input[828]), .B(n22512), .Z(n22514) );
  XNOR U21905 ( .A(n22515), .B(n22516), .Z(n22512) );
  AND U21906 ( .A(n1044), .B(n22517), .Z(n22516) );
  XOR U21907 ( .A(n22518), .B(n22519), .Z(n22510) );
  AND U21908 ( .A(n1048), .B(n22509), .Z(n22519) );
  XNOR U21909 ( .A(n22520), .B(n22507), .Z(n22509) );
  XOR U21910 ( .A(n22521), .B(n22522), .Z(n22507) );
  AND U21911 ( .A(n1071), .B(n22523), .Z(n22522) );
  IV U21912 ( .A(n22518), .Z(n22520) );
  XOR U21913 ( .A(n22524), .B(n22525), .Z(n22518) );
  AND U21914 ( .A(n1055), .B(n22517), .Z(n22525) );
  XNOR U21915 ( .A(n22515), .B(n22524), .Z(n22517) );
  XNOR U21916 ( .A(n22526), .B(n22527), .Z(n22515) );
  AND U21917 ( .A(n1059), .B(n22528), .Z(n22527) );
  XOR U21918 ( .A(p_input[844]), .B(n22526), .Z(n22528) );
  XNOR U21919 ( .A(n22529), .B(n22530), .Z(n22526) );
  AND U21920 ( .A(n1063), .B(n22531), .Z(n22530) );
  XOR U21921 ( .A(n22532), .B(n22533), .Z(n22524) );
  AND U21922 ( .A(n1067), .B(n22523), .Z(n22533) );
  XNOR U21923 ( .A(n22534), .B(n22521), .Z(n22523) );
  XOR U21924 ( .A(n22535), .B(n22536), .Z(n22521) );
  AND U21925 ( .A(n1090), .B(n22537), .Z(n22536) );
  IV U21926 ( .A(n22532), .Z(n22534) );
  XOR U21927 ( .A(n22538), .B(n22539), .Z(n22532) );
  AND U21928 ( .A(n1074), .B(n22531), .Z(n22539) );
  XNOR U21929 ( .A(n22529), .B(n22538), .Z(n22531) );
  XNOR U21930 ( .A(n22540), .B(n22541), .Z(n22529) );
  AND U21931 ( .A(n1078), .B(n22542), .Z(n22541) );
  XOR U21932 ( .A(p_input[860]), .B(n22540), .Z(n22542) );
  XNOR U21933 ( .A(n22543), .B(n22544), .Z(n22540) );
  AND U21934 ( .A(n1082), .B(n22545), .Z(n22544) );
  XOR U21935 ( .A(n22546), .B(n22547), .Z(n22538) );
  AND U21936 ( .A(n1086), .B(n22537), .Z(n22547) );
  XNOR U21937 ( .A(n22548), .B(n22535), .Z(n22537) );
  XOR U21938 ( .A(n22549), .B(n22550), .Z(n22535) );
  AND U21939 ( .A(n1109), .B(n22551), .Z(n22550) );
  IV U21940 ( .A(n22546), .Z(n22548) );
  XOR U21941 ( .A(n22552), .B(n22553), .Z(n22546) );
  AND U21942 ( .A(n1093), .B(n22545), .Z(n22553) );
  XNOR U21943 ( .A(n22543), .B(n22552), .Z(n22545) );
  XNOR U21944 ( .A(n22554), .B(n22555), .Z(n22543) );
  AND U21945 ( .A(n1097), .B(n22556), .Z(n22555) );
  XOR U21946 ( .A(p_input[876]), .B(n22554), .Z(n22556) );
  XNOR U21947 ( .A(n22557), .B(n22558), .Z(n22554) );
  AND U21948 ( .A(n1101), .B(n22559), .Z(n22558) );
  XOR U21949 ( .A(n22560), .B(n22561), .Z(n22552) );
  AND U21950 ( .A(n1105), .B(n22551), .Z(n22561) );
  XNOR U21951 ( .A(n22562), .B(n22549), .Z(n22551) );
  XOR U21952 ( .A(n22563), .B(n22564), .Z(n22549) );
  AND U21953 ( .A(n1128), .B(n22565), .Z(n22564) );
  IV U21954 ( .A(n22560), .Z(n22562) );
  XOR U21955 ( .A(n22566), .B(n22567), .Z(n22560) );
  AND U21956 ( .A(n1112), .B(n22559), .Z(n22567) );
  XNOR U21957 ( .A(n22557), .B(n22566), .Z(n22559) );
  XNOR U21958 ( .A(n22568), .B(n22569), .Z(n22557) );
  AND U21959 ( .A(n1116), .B(n22570), .Z(n22569) );
  XOR U21960 ( .A(p_input[892]), .B(n22568), .Z(n22570) );
  XNOR U21961 ( .A(n22571), .B(n22572), .Z(n22568) );
  AND U21962 ( .A(n1120), .B(n22573), .Z(n22572) );
  XOR U21963 ( .A(n22574), .B(n22575), .Z(n22566) );
  AND U21964 ( .A(n1124), .B(n22565), .Z(n22575) );
  XNOR U21965 ( .A(n22576), .B(n22563), .Z(n22565) );
  XOR U21966 ( .A(n22577), .B(n22578), .Z(n22563) );
  AND U21967 ( .A(n1147), .B(n22579), .Z(n22578) );
  IV U21968 ( .A(n22574), .Z(n22576) );
  XOR U21969 ( .A(n22580), .B(n22581), .Z(n22574) );
  AND U21970 ( .A(n1131), .B(n22573), .Z(n22581) );
  XNOR U21971 ( .A(n22571), .B(n22580), .Z(n22573) );
  XNOR U21972 ( .A(n22582), .B(n22583), .Z(n22571) );
  AND U21973 ( .A(n1135), .B(n22584), .Z(n22583) );
  XOR U21974 ( .A(p_input[908]), .B(n22582), .Z(n22584) );
  XNOR U21975 ( .A(n22585), .B(n22586), .Z(n22582) );
  AND U21976 ( .A(n1139), .B(n22587), .Z(n22586) );
  XOR U21977 ( .A(n22588), .B(n22589), .Z(n22580) );
  AND U21978 ( .A(n1143), .B(n22579), .Z(n22589) );
  XNOR U21979 ( .A(n22590), .B(n22577), .Z(n22579) );
  XOR U21980 ( .A(n22591), .B(n22592), .Z(n22577) );
  AND U21981 ( .A(n1166), .B(n22593), .Z(n22592) );
  IV U21982 ( .A(n22588), .Z(n22590) );
  XOR U21983 ( .A(n22594), .B(n22595), .Z(n22588) );
  AND U21984 ( .A(n1150), .B(n22587), .Z(n22595) );
  XNOR U21985 ( .A(n22585), .B(n22594), .Z(n22587) );
  XNOR U21986 ( .A(n22596), .B(n22597), .Z(n22585) );
  AND U21987 ( .A(n1154), .B(n22598), .Z(n22597) );
  XOR U21988 ( .A(p_input[924]), .B(n22596), .Z(n22598) );
  XNOR U21989 ( .A(n22599), .B(n22600), .Z(n22596) );
  AND U21990 ( .A(n1158), .B(n22601), .Z(n22600) );
  XOR U21991 ( .A(n22602), .B(n22603), .Z(n22594) );
  AND U21992 ( .A(n1162), .B(n22593), .Z(n22603) );
  XNOR U21993 ( .A(n22604), .B(n22591), .Z(n22593) );
  XOR U21994 ( .A(n22605), .B(n22606), .Z(n22591) );
  AND U21995 ( .A(n1185), .B(n22607), .Z(n22606) );
  IV U21996 ( .A(n22602), .Z(n22604) );
  XOR U21997 ( .A(n22608), .B(n22609), .Z(n22602) );
  AND U21998 ( .A(n1169), .B(n22601), .Z(n22609) );
  XNOR U21999 ( .A(n22599), .B(n22608), .Z(n22601) );
  XNOR U22000 ( .A(n22610), .B(n22611), .Z(n22599) );
  AND U22001 ( .A(n1173), .B(n22612), .Z(n22611) );
  XOR U22002 ( .A(p_input[940]), .B(n22610), .Z(n22612) );
  XNOR U22003 ( .A(n22613), .B(n22614), .Z(n22610) );
  AND U22004 ( .A(n1177), .B(n22615), .Z(n22614) );
  XOR U22005 ( .A(n22616), .B(n22617), .Z(n22608) );
  AND U22006 ( .A(n1181), .B(n22607), .Z(n22617) );
  XNOR U22007 ( .A(n22618), .B(n22605), .Z(n22607) );
  XOR U22008 ( .A(n22619), .B(n22620), .Z(n22605) );
  AND U22009 ( .A(n1204), .B(n22621), .Z(n22620) );
  IV U22010 ( .A(n22616), .Z(n22618) );
  XOR U22011 ( .A(n22622), .B(n22623), .Z(n22616) );
  AND U22012 ( .A(n1188), .B(n22615), .Z(n22623) );
  XNOR U22013 ( .A(n22613), .B(n22622), .Z(n22615) );
  XNOR U22014 ( .A(n22624), .B(n22625), .Z(n22613) );
  AND U22015 ( .A(n1192), .B(n22626), .Z(n22625) );
  XOR U22016 ( .A(p_input[956]), .B(n22624), .Z(n22626) );
  XNOR U22017 ( .A(n22627), .B(n22628), .Z(n22624) );
  AND U22018 ( .A(n1196), .B(n22629), .Z(n22628) );
  XOR U22019 ( .A(n22630), .B(n22631), .Z(n22622) );
  AND U22020 ( .A(n1200), .B(n22621), .Z(n22631) );
  XNOR U22021 ( .A(n22632), .B(n22619), .Z(n22621) );
  XOR U22022 ( .A(n22633), .B(n22634), .Z(n22619) );
  AND U22023 ( .A(n1223), .B(n22635), .Z(n22634) );
  IV U22024 ( .A(n22630), .Z(n22632) );
  XOR U22025 ( .A(n22636), .B(n22637), .Z(n22630) );
  AND U22026 ( .A(n1207), .B(n22629), .Z(n22637) );
  XNOR U22027 ( .A(n22627), .B(n22636), .Z(n22629) );
  XNOR U22028 ( .A(n22638), .B(n22639), .Z(n22627) );
  AND U22029 ( .A(n1211), .B(n22640), .Z(n22639) );
  XOR U22030 ( .A(p_input[972]), .B(n22638), .Z(n22640) );
  XNOR U22031 ( .A(n22641), .B(n22642), .Z(n22638) );
  AND U22032 ( .A(n1215), .B(n22643), .Z(n22642) );
  XOR U22033 ( .A(n22644), .B(n22645), .Z(n22636) );
  AND U22034 ( .A(n1219), .B(n22635), .Z(n22645) );
  XNOR U22035 ( .A(n22646), .B(n22633), .Z(n22635) );
  XOR U22036 ( .A(n22647), .B(n22648), .Z(n22633) );
  AND U22037 ( .A(n1242), .B(n22649), .Z(n22648) );
  IV U22038 ( .A(n22644), .Z(n22646) );
  XOR U22039 ( .A(n22650), .B(n22651), .Z(n22644) );
  AND U22040 ( .A(n1226), .B(n22643), .Z(n22651) );
  XNOR U22041 ( .A(n22641), .B(n22650), .Z(n22643) );
  XNOR U22042 ( .A(n22652), .B(n22653), .Z(n22641) );
  AND U22043 ( .A(n1230), .B(n22654), .Z(n22653) );
  XOR U22044 ( .A(p_input[988]), .B(n22652), .Z(n22654) );
  XNOR U22045 ( .A(n22655), .B(n22656), .Z(n22652) );
  AND U22046 ( .A(n1234), .B(n22657), .Z(n22656) );
  XOR U22047 ( .A(n22658), .B(n22659), .Z(n22650) );
  AND U22048 ( .A(n1238), .B(n22649), .Z(n22659) );
  XNOR U22049 ( .A(n22660), .B(n22647), .Z(n22649) );
  XOR U22050 ( .A(n22661), .B(n22662), .Z(n22647) );
  AND U22051 ( .A(n1261), .B(n22663), .Z(n22662) );
  IV U22052 ( .A(n22658), .Z(n22660) );
  XOR U22053 ( .A(n22664), .B(n22665), .Z(n22658) );
  AND U22054 ( .A(n1245), .B(n22657), .Z(n22665) );
  XNOR U22055 ( .A(n22655), .B(n22664), .Z(n22657) );
  XNOR U22056 ( .A(n22666), .B(n22667), .Z(n22655) );
  AND U22057 ( .A(n1249), .B(n22668), .Z(n22667) );
  XOR U22058 ( .A(p_input[1004]), .B(n22666), .Z(n22668) );
  XNOR U22059 ( .A(n22669), .B(n22670), .Z(n22666) );
  AND U22060 ( .A(n1253), .B(n22671), .Z(n22670) );
  XOR U22061 ( .A(n22672), .B(n22673), .Z(n22664) );
  AND U22062 ( .A(n1257), .B(n22663), .Z(n22673) );
  XNOR U22063 ( .A(n22674), .B(n22661), .Z(n22663) );
  XOR U22064 ( .A(n22675), .B(n22676), .Z(n22661) );
  AND U22065 ( .A(n1280), .B(n22677), .Z(n22676) );
  IV U22066 ( .A(n22672), .Z(n22674) );
  XOR U22067 ( .A(n22678), .B(n22679), .Z(n22672) );
  AND U22068 ( .A(n1264), .B(n22671), .Z(n22679) );
  XNOR U22069 ( .A(n22669), .B(n22678), .Z(n22671) );
  XNOR U22070 ( .A(n22680), .B(n22681), .Z(n22669) );
  AND U22071 ( .A(n1268), .B(n22682), .Z(n22681) );
  XOR U22072 ( .A(p_input[1020]), .B(n22680), .Z(n22682) );
  XNOR U22073 ( .A(n22683), .B(n22684), .Z(n22680) );
  AND U22074 ( .A(n1272), .B(n22685), .Z(n22684) );
  XOR U22075 ( .A(n22686), .B(n22687), .Z(n22678) );
  AND U22076 ( .A(n1276), .B(n22677), .Z(n22687) );
  XNOR U22077 ( .A(n22688), .B(n22675), .Z(n22677) );
  XOR U22078 ( .A(n22689), .B(n22690), .Z(n22675) );
  AND U22079 ( .A(n1299), .B(n22691), .Z(n22690) );
  IV U22080 ( .A(n22686), .Z(n22688) );
  XOR U22081 ( .A(n22692), .B(n22693), .Z(n22686) );
  AND U22082 ( .A(n1283), .B(n22685), .Z(n22693) );
  XNOR U22083 ( .A(n22683), .B(n22692), .Z(n22685) );
  XNOR U22084 ( .A(n22694), .B(n22695), .Z(n22683) );
  AND U22085 ( .A(n1287), .B(n22696), .Z(n22695) );
  XOR U22086 ( .A(p_input[1036]), .B(n22694), .Z(n22696) );
  XNOR U22087 ( .A(n22697), .B(n22698), .Z(n22694) );
  AND U22088 ( .A(n1291), .B(n22699), .Z(n22698) );
  XOR U22089 ( .A(n22700), .B(n22701), .Z(n22692) );
  AND U22090 ( .A(n1295), .B(n22691), .Z(n22701) );
  XNOR U22091 ( .A(n22702), .B(n22689), .Z(n22691) );
  XOR U22092 ( .A(n22703), .B(n22704), .Z(n22689) );
  AND U22093 ( .A(n1318), .B(n22705), .Z(n22704) );
  IV U22094 ( .A(n22700), .Z(n22702) );
  XOR U22095 ( .A(n22706), .B(n22707), .Z(n22700) );
  AND U22096 ( .A(n1302), .B(n22699), .Z(n22707) );
  XNOR U22097 ( .A(n22697), .B(n22706), .Z(n22699) );
  XNOR U22098 ( .A(n22708), .B(n22709), .Z(n22697) );
  AND U22099 ( .A(n1306), .B(n22710), .Z(n22709) );
  XOR U22100 ( .A(p_input[1052]), .B(n22708), .Z(n22710) );
  XNOR U22101 ( .A(n22711), .B(n22712), .Z(n22708) );
  AND U22102 ( .A(n1310), .B(n22713), .Z(n22712) );
  XOR U22103 ( .A(n22714), .B(n22715), .Z(n22706) );
  AND U22104 ( .A(n1314), .B(n22705), .Z(n22715) );
  XNOR U22105 ( .A(n22716), .B(n22703), .Z(n22705) );
  XOR U22106 ( .A(n22717), .B(n22718), .Z(n22703) );
  AND U22107 ( .A(n1337), .B(n22719), .Z(n22718) );
  IV U22108 ( .A(n22714), .Z(n22716) );
  XOR U22109 ( .A(n22720), .B(n22721), .Z(n22714) );
  AND U22110 ( .A(n1321), .B(n22713), .Z(n22721) );
  XNOR U22111 ( .A(n22711), .B(n22720), .Z(n22713) );
  XNOR U22112 ( .A(n22722), .B(n22723), .Z(n22711) );
  AND U22113 ( .A(n1325), .B(n22724), .Z(n22723) );
  XOR U22114 ( .A(p_input[1068]), .B(n22722), .Z(n22724) );
  XNOR U22115 ( .A(n22725), .B(n22726), .Z(n22722) );
  AND U22116 ( .A(n1329), .B(n22727), .Z(n22726) );
  XOR U22117 ( .A(n22728), .B(n22729), .Z(n22720) );
  AND U22118 ( .A(n1333), .B(n22719), .Z(n22729) );
  XNOR U22119 ( .A(n22730), .B(n22717), .Z(n22719) );
  XOR U22120 ( .A(n22731), .B(n22732), .Z(n22717) );
  AND U22121 ( .A(n1356), .B(n22733), .Z(n22732) );
  IV U22122 ( .A(n22728), .Z(n22730) );
  XOR U22123 ( .A(n22734), .B(n22735), .Z(n22728) );
  AND U22124 ( .A(n1340), .B(n22727), .Z(n22735) );
  XNOR U22125 ( .A(n22725), .B(n22734), .Z(n22727) );
  XNOR U22126 ( .A(n22736), .B(n22737), .Z(n22725) );
  AND U22127 ( .A(n1344), .B(n22738), .Z(n22737) );
  XOR U22128 ( .A(p_input[1084]), .B(n22736), .Z(n22738) );
  XNOR U22129 ( .A(n22739), .B(n22740), .Z(n22736) );
  AND U22130 ( .A(n1348), .B(n22741), .Z(n22740) );
  XOR U22131 ( .A(n22742), .B(n22743), .Z(n22734) );
  AND U22132 ( .A(n1352), .B(n22733), .Z(n22743) );
  XNOR U22133 ( .A(n22744), .B(n22731), .Z(n22733) );
  XOR U22134 ( .A(n22745), .B(n22746), .Z(n22731) );
  AND U22135 ( .A(n1375), .B(n22747), .Z(n22746) );
  IV U22136 ( .A(n22742), .Z(n22744) );
  XOR U22137 ( .A(n22748), .B(n22749), .Z(n22742) );
  AND U22138 ( .A(n1359), .B(n22741), .Z(n22749) );
  XNOR U22139 ( .A(n22739), .B(n22748), .Z(n22741) );
  XNOR U22140 ( .A(n22750), .B(n22751), .Z(n22739) );
  AND U22141 ( .A(n1363), .B(n22752), .Z(n22751) );
  XOR U22142 ( .A(p_input[1100]), .B(n22750), .Z(n22752) );
  XNOR U22143 ( .A(n22753), .B(n22754), .Z(n22750) );
  AND U22144 ( .A(n1367), .B(n22755), .Z(n22754) );
  XOR U22145 ( .A(n22756), .B(n22757), .Z(n22748) );
  AND U22146 ( .A(n1371), .B(n22747), .Z(n22757) );
  XNOR U22147 ( .A(n22758), .B(n22745), .Z(n22747) );
  XOR U22148 ( .A(n22759), .B(n22760), .Z(n22745) );
  AND U22149 ( .A(n1394), .B(n22761), .Z(n22760) );
  IV U22150 ( .A(n22756), .Z(n22758) );
  XOR U22151 ( .A(n22762), .B(n22763), .Z(n22756) );
  AND U22152 ( .A(n1378), .B(n22755), .Z(n22763) );
  XNOR U22153 ( .A(n22753), .B(n22762), .Z(n22755) );
  XNOR U22154 ( .A(n22764), .B(n22765), .Z(n22753) );
  AND U22155 ( .A(n1382), .B(n22766), .Z(n22765) );
  XOR U22156 ( .A(p_input[1116]), .B(n22764), .Z(n22766) );
  XNOR U22157 ( .A(n22767), .B(n22768), .Z(n22764) );
  AND U22158 ( .A(n1386), .B(n22769), .Z(n22768) );
  XOR U22159 ( .A(n22770), .B(n22771), .Z(n22762) );
  AND U22160 ( .A(n1390), .B(n22761), .Z(n22771) );
  XNOR U22161 ( .A(n22772), .B(n22759), .Z(n22761) );
  XOR U22162 ( .A(n22773), .B(n22774), .Z(n22759) );
  AND U22163 ( .A(n1413), .B(n22775), .Z(n22774) );
  IV U22164 ( .A(n22770), .Z(n22772) );
  XOR U22165 ( .A(n22776), .B(n22777), .Z(n22770) );
  AND U22166 ( .A(n1397), .B(n22769), .Z(n22777) );
  XNOR U22167 ( .A(n22767), .B(n22776), .Z(n22769) );
  XNOR U22168 ( .A(n22778), .B(n22779), .Z(n22767) );
  AND U22169 ( .A(n1401), .B(n22780), .Z(n22779) );
  XOR U22170 ( .A(p_input[1132]), .B(n22778), .Z(n22780) );
  XNOR U22171 ( .A(n22781), .B(n22782), .Z(n22778) );
  AND U22172 ( .A(n1405), .B(n22783), .Z(n22782) );
  XOR U22173 ( .A(n22784), .B(n22785), .Z(n22776) );
  AND U22174 ( .A(n1409), .B(n22775), .Z(n22785) );
  XNOR U22175 ( .A(n22786), .B(n22773), .Z(n22775) );
  XOR U22176 ( .A(n22787), .B(n22788), .Z(n22773) );
  AND U22177 ( .A(n1432), .B(n22789), .Z(n22788) );
  IV U22178 ( .A(n22784), .Z(n22786) );
  XOR U22179 ( .A(n22790), .B(n22791), .Z(n22784) );
  AND U22180 ( .A(n1416), .B(n22783), .Z(n22791) );
  XNOR U22181 ( .A(n22781), .B(n22790), .Z(n22783) );
  XNOR U22182 ( .A(n22792), .B(n22793), .Z(n22781) );
  AND U22183 ( .A(n1420), .B(n22794), .Z(n22793) );
  XOR U22184 ( .A(p_input[1148]), .B(n22792), .Z(n22794) );
  XNOR U22185 ( .A(n22795), .B(n22796), .Z(n22792) );
  AND U22186 ( .A(n1424), .B(n22797), .Z(n22796) );
  XOR U22187 ( .A(n22798), .B(n22799), .Z(n22790) );
  AND U22188 ( .A(n1428), .B(n22789), .Z(n22799) );
  XNOR U22189 ( .A(n22800), .B(n22787), .Z(n22789) );
  XOR U22190 ( .A(n22801), .B(n22802), .Z(n22787) );
  AND U22191 ( .A(n1451), .B(n22803), .Z(n22802) );
  IV U22192 ( .A(n22798), .Z(n22800) );
  XOR U22193 ( .A(n22804), .B(n22805), .Z(n22798) );
  AND U22194 ( .A(n1435), .B(n22797), .Z(n22805) );
  XNOR U22195 ( .A(n22795), .B(n22804), .Z(n22797) );
  XNOR U22196 ( .A(n22806), .B(n22807), .Z(n22795) );
  AND U22197 ( .A(n1439), .B(n22808), .Z(n22807) );
  XOR U22198 ( .A(p_input[1164]), .B(n22806), .Z(n22808) );
  XNOR U22199 ( .A(n22809), .B(n22810), .Z(n22806) );
  AND U22200 ( .A(n1443), .B(n22811), .Z(n22810) );
  XOR U22201 ( .A(n22812), .B(n22813), .Z(n22804) );
  AND U22202 ( .A(n1447), .B(n22803), .Z(n22813) );
  XNOR U22203 ( .A(n22814), .B(n22801), .Z(n22803) );
  XOR U22204 ( .A(n22815), .B(n22816), .Z(n22801) );
  AND U22205 ( .A(n1470), .B(n22817), .Z(n22816) );
  IV U22206 ( .A(n22812), .Z(n22814) );
  XOR U22207 ( .A(n22818), .B(n22819), .Z(n22812) );
  AND U22208 ( .A(n1454), .B(n22811), .Z(n22819) );
  XNOR U22209 ( .A(n22809), .B(n22818), .Z(n22811) );
  XNOR U22210 ( .A(n22820), .B(n22821), .Z(n22809) );
  AND U22211 ( .A(n1458), .B(n22822), .Z(n22821) );
  XOR U22212 ( .A(p_input[1180]), .B(n22820), .Z(n22822) );
  XNOR U22213 ( .A(n22823), .B(n22824), .Z(n22820) );
  AND U22214 ( .A(n1462), .B(n22825), .Z(n22824) );
  XOR U22215 ( .A(n22826), .B(n22827), .Z(n22818) );
  AND U22216 ( .A(n1466), .B(n22817), .Z(n22827) );
  XNOR U22217 ( .A(n22828), .B(n22815), .Z(n22817) );
  XOR U22218 ( .A(n22829), .B(n22830), .Z(n22815) );
  AND U22219 ( .A(n1489), .B(n22831), .Z(n22830) );
  IV U22220 ( .A(n22826), .Z(n22828) );
  XOR U22221 ( .A(n22832), .B(n22833), .Z(n22826) );
  AND U22222 ( .A(n1473), .B(n22825), .Z(n22833) );
  XNOR U22223 ( .A(n22823), .B(n22832), .Z(n22825) );
  XNOR U22224 ( .A(n22834), .B(n22835), .Z(n22823) );
  AND U22225 ( .A(n1477), .B(n22836), .Z(n22835) );
  XOR U22226 ( .A(p_input[1196]), .B(n22834), .Z(n22836) );
  XNOR U22227 ( .A(n22837), .B(n22838), .Z(n22834) );
  AND U22228 ( .A(n1481), .B(n22839), .Z(n22838) );
  XOR U22229 ( .A(n22840), .B(n22841), .Z(n22832) );
  AND U22230 ( .A(n1485), .B(n22831), .Z(n22841) );
  XNOR U22231 ( .A(n22842), .B(n22829), .Z(n22831) );
  XOR U22232 ( .A(n22843), .B(n22844), .Z(n22829) );
  AND U22233 ( .A(n1508), .B(n22845), .Z(n22844) );
  IV U22234 ( .A(n22840), .Z(n22842) );
  XOR U22235 ( .A(n22846), .B(n22847), .Z(n22840) );
  AND U22236 ( .A(n1492), .B(n22839), .Z(n22847) );
  XNOR U22237 ( .A(n22837), .B(n22846), .Z(n22839) );
  XNOR U22238 ( .A(n22848), .B(n22849), .Z(n22837) );
  AND U22239 ( .A(n1496), .B(n22850), .Z(n22849) );
  XOR U22240 ( .A(p_input[1212]), .B(n22848), .Z(n22850) );
  XNOR U22241 ( .A(n22851), .B(n22852), .Z(n22848) );
  AND U22242 ( .A(n1500), .B(n22853), .Z(n22852) );
  XOR U22243 ( .A(n22854), .B(n22855), .Z(n22846) );
  AND U22244 ( .A(n1504), .B(n22845), .Z(n22855) );
  XNOR U22245 ( .A(n22856), .B(n22843), .Z(n22845) );
  XOR U22246 ( .A(n22857), .B(n22858), .Z(n22843) );
  AND U22247 ( .A(n1527), .B(n22859), .Z(n22858) );
  IV U22248 ( .A(n22854), .Z(n22856) );
  XOR U22249 ( .A(n22860), .B(n22861), .Z(n22854) );
  AND U22250 ( .A(n1511), .B(n22853), .Z(n22861) );
  XNOR U22251 ( .A(n22851), .B(n22860), .Z(n22853) );
  XNOR U22252 ( .A(n22862), .B(n22863), .Z(n22851) );
  AND U22253 ( .A(n1515), .B(n22864), .Z(n22863) );
  XOR U22254 ( .A(p_input[1228]), .B(n22862), .Z(n22864) );
  XNOR U22255 ( .A(n22865), .B(n22866), .Z(n22862) );
  AND U22256 ( .A(n1519), .B(n22867), .Z(n22866) );
  XOR U22257 ( .A(n22868), .B(n22869), .Z(n22860) );
  AND U22258 ( .A(n1523), .B(n22859), .Z(n22869) );
  XNOR U22259 ( .A(n22870), .B(n22857), .Z(n22859) );
  XOR U22260 ( .A(n22871), .B(n22872), .Z(n22857) );
  AND U22261 ( .A(n1546), .B(n22873), .Z(n22872) );
  IV U22262 ( .A(n22868), .Z(n22870) );
  XOR U22263 ( .A(n22874), .B(n22875), .Z(n22868) );
  AND U22264 ( .A(n1530), .B(n22867), .Z(n22875) );
  XNOR U22265 ( .A(n22865), .B(n22874), .Z(n22867) );
  XNOR U22266 ( .A(n22876), .B(n22877), .Z(n22865) );
  AND U22267 ( .A(n1534), .B(n22878), .Z(n22877) );
  XOR U22268 ( .A(p_input[1244]), .B(n22876), .Z(n22878) );
  XNOR U22269 ( .A(n22879), .B(n22880), .Z(n22876) );
  AND U22270 ( .A(n1538), .B(n22881), .Z(n22880) );
  XOR U22271 ( .A(n22882), .B(n22883), .Z(n22874) );
  AND U22272 ( .A(n1542), .B(n22873), .Z(n22883) );
  XNOR U22273 ( .A(n22884), .B(n22871), .Z(n22873) );
  XOR U22274 ( .A(n22885), .B(n22886), .Z(n22871) );
  AND U22275 ( .A(n1565), .B(n22887), .Z(n22886) );
  IV U22276 ( .A(n22882), .Z(n22884) );
  XOR U22277 ( .A(n22888), .B(n22889), .Z(n22882) );
  AND U22278 ( .A(n1549), .B(n22881), .Z(n22889) );
  XNOR U22279 ( .A(n22879), .B(n22888), .Z(n22881) );
  XNOR U22280 ( .A(n22890), .B(n22891), .Z(n22879) );
  AND U22281 ( .A(n1553), .B(n22892), .Z(n22891) );
  XOR U22282 ( .A(p_input[1260]), .B(n22890), .Z(n22892) );
  XNOR U22283 ( .A(n22893), .B(n22894), .Z(n22890) );
  AND U22284 ( .A(n1557), .B(n22895), .Z(n22894) );
  XOR U22285 ( .A(n22896), .B(n22897), .Z(n22888) );
  AND U22286 ( .A(n1561), .B(n22887), .Z(n22897) );
  XNOR U22287 ( .A(n22898), .B(n22885), .Z(n22887) );
  XOR U22288 ( .A(n22899), .B(n22900), .Z(n22885) );
  AND U22289 ( .A(n1584), .B(n22901), .Z(n22900) );
  IV U22290 ( .A(n22896), .Z(n22898) );
  XOR U22291 ( .A(n22902), .B(n22903), .Z(n22896) );
  AND U22292 ( .A(n1568), .B(n22895), .Z(n22903) );
  XNOR U22293 ( .A(n22893), .B(n22902), .Z(n22895) );
  XNOR U22294 ( .A(n22904), .B(n22905), .Z(n22893) );
  AND U22295 ( .A(n1572), .B(n22906), .Z(n22905) );
  XOR U22296 ( .A(p_input[1276]), .B(n22904), .Z(n22906) );
  XNOR U22297 ( .A(n22907), .B(n22908), .Z(n22904) );
  AND U22298 ( .A(n1576), .B(n22909), .Z(n22908) );
  XOR U22299 ( .A(n22910), .B(n22911), .Z(n22902) );
  AND U22300 ( .A(n1580), .B(n22901), .Z(n22911) );
  XNOR U22301 ( .A(n22912), .B(n22899), .Z(n22901) );
  XOR U22302 ( .A(n22913), .B(n22914), .Z(n22899) );
  AND U22303 ( .A(n1603), .B(n22915), .Z(n22914) );
  IV U22304 ( .A(n22910), .Z(n22912) );
  XOR U22305 ( .A(n22916), .B(n22917), .Z(n22910) );
  AND U22306 ( .A(n1587), .B(n22909), .Z(n22917) );
  XNOR U22307 ( .A(n22907), .B(n22916), .Z(n22909) );
  XNOR U22308 ( .A(n22918), .B(n22919), .Z(n22907) );
  AND U22309 ( .A(n1591), .B(n22920), .Z(n22919) );
  XOR U22310 ( .A(p_input[1292]), .B(n22918), .Z(n22920) );
  XNOR U22311 ( .A(n22921), .B(n22922), .Z(n22918) );
  AND U22312 ( .A(n1595), .B(n22923), .Z(n22922) );
  XOR U22313 ( .A(n22924), .B(n22925), .Z(n22916) );
  AND U22314 ( .A(n1599), .B(n22915), .Z(n22925) );
  XNOR U22315 ( .A(n22926), .B(n22913), .Z(n22915) );
  XOR U22316 ( .A(n22927), .B(n22928), .Z(n22913) );
  AND U22317 ( .A(n1622), .B(n22929), .Z(n22928) );
  IV U22318 ( .A(n22924), .Z(n22926) );
  XOR U22319 ( .A(n22930), .B(n22931), .Z(n22924) );
  AND U22320 ( .A(n1606), .B(n22923), .Z(n22931) );
  XNOR U22321 ( .A(n22921), .B(n22930), .Z(n22923) );
  XNOR U22322 ( .A(n22932), .B(n22933), .Z(n22921) );
  AND U22323 ( .A(n1610), .B(n22934), .Z(n22933) );
  XOR U22324 ( .A(p_input[1308]), .B(n22932), .Z(n22934) );
  XNOR U22325 ( .A(n22935), .B(n22936), .Z(n22932) );
  AND U22326 ( .A(n1614), .B(n22937), .Z(n22936) );
  XOR U22327 ( .A(n22938), .B(n22939), .Z(n22930) );
  AND U22328 ( .A(n1618), .B(n22929), .Z(n22939) );
  XNOR U22329 ( .A(n22940), .B(n22927), .Z(n22929) );
  XOR U22330 ( .A(n22941), .B(n22942), .Z(n22927) );
  AND U22331 ( .A(n1641), .B(n22943), .Z(n22942) );
  IV U22332 ( .A(n22938), .Z(n22940) );
  XOR U22333 ( .A(n22944), .B(n22945), .Z(n22938) );
  AND U22334 ( .A(n1625), .B(n22937), .Z(n22945) );
  XNOR U22335 ( .A(n22935), .B(n22944), .Z(n22937) );
  XNOR U22336 ( .A(n22946), .B(n22947), .Z(n22935) );
  AND U22337 ( .A(n1629), .B(n22948), .Z(n22947) );
  XOR U22338 ( .A(p_input[1324]), .B(n22946), .Z(n22948) );
  XNOR U22339 ( .A(n22949), .B(n22950), .Z(n22946) );
  AND U22340 ( .A(n1633), .B(n22951), .Z(n22950) );
  XOR U22341 ( .A(n22952), .B(n22953), .Z(n22944) );
  AND U22342 ( .A(n1637), .B(n22943), .Z(n22953) );
  XNOR U22343 ( .A(n22954), .B(n22941), .Z(n22943) );
  XOR U22344 ( .A(n22955), .B(n22956), .Z(n22941) );
  AND U22345 ( .A(n1660), .B(n22957), .Z(n22956) );
  IV U22346 ( .A(n22952), .Z(n22954) );
  XOR U22347 ( .A(n22958), .B(n22959), .Z(n22952) );
  AND U22348 ( .A(n1644), .B(n22951), .Z(n22959) );
  XNOR U22349 ( .A(n22949), .B(n22958), .Z(n22951) );
  XNOR U22350 ( .A(n22960), .B(n22961), .Z(n22949) );
  AND U22351 ( .A(n1648), .B(n22962), .Z(n22961) );
  XOR U22352 ( .A(p_input[1340]), .B(n22960), .Z(n22962) );
  XNOR U22353 ( .A(n22963), .B(n22964), .Z(n22960) );
  AND U22354 ( .A(n1652), .B(n22965), .Z(n22964) );
  XOR U22355 ( .A(n22966), .B(n22967), .Z(n22958) );
  AND U22356 ( .A(n1656), .B(n22957), .Z(n22967) );
  XNOR U22357 ( .A(n22968), .B(n22955), .Z(n22957) );
  XOR U22358 ( .A(n22969), .B(n22970), .Z(n22955) );
  AND U22359 ( .A(n1679), .B(n22971), .Z(n22970) );
  IV U22360 ( .A(n22966), .Z(n22968) );
  XOR U22361 ( .A(n22972), .B(n22973), .Z(n22966) );
  AND U22362 ( .A(n1663), .B(n22965), .Z(n22973) );
  XNOR U22363 ( .A(n22963), .B(n22972), .Z(n22965) );
  XNOR U22364 ( .A(n22974), .B(n22975), .Z(n22963) );
  AND U22365 ( .A(n1667), .B(n22976), .Z(n22975) );
  XOR U22366 ( .A(p_input[1356]), .B(n22974), .Z(n22976) );
  XNOR U22367 ( .A(n22977), .B(n22978), .Z(n22974) );
  AND U22368 ( .A(n1671), .B(n22979), .Z(n22978) );
  XOR U22369 ( .A(n22980), .B(n22981), .Z(n22972) );
  AND U22370 ( .A(n1675), .B(n22971), .Z(n22981) );
  XNOR U22371 ( .A(n22982), .B(n22969), .Z(n22971) );
  XOR U22372 ( .A(n22983), .B(n22984), .Z(n22969) );
  AND U22373 ( .A(n1698), .B(n22985), .Z(n22984) );
  IV U22374 ( .A(n22980), .Z(n22982) );
  XOR U22375 ( .A(n22986), .B(n22987), .Z(n22980) );
  AND U22376 ( .A(n1682), .B(n22979), .Z(n22987) );
  XNOR U22377 ( .A(n22977), .B(n22986), .Z(n22979) );
  XNOR U22378 ( .A(n22988), .B(n22989), .Z(n22977) );
  AND U22379 ( .A(n1686), .B(n22990), .Z(n22989) );
  XOR U22380 ( .A(p_input[1372]), .B(n22988), .Z(n22990) );
  XNOR U22381 ( .A(n22991), .B(n22992), .Z(n22988) );
  AND U22382 ( .A(n1690), .B(n22993), .Z(n22992) );
  XOR U22383 ( .A(n22994), .B(n22995), .Z(n22986) );
  AND U22384 ( .A(n1694), .B(n22985), .Z(n22995) );
  XNOR U22385 ( .A(n22996), .B(n22983), .Z(n22985) );
  XOR U22386 ( .A(n22997), .B(n22998), .Z(n22983) );
  AND U22387 ( .A(n1717), .B(n22999), .Z(n22998) );
  IV U22388 ( .A(n22994), .Z(n22996) );
  XOR U22389 ( .A(n23000), .B(n23001), .Z(n22994) );
  AND U22390 ( .A(n1701), .B(n22993), .Z(n23001) );
  XNOR U22391 ( .A(n22991), .B(n23000), .Z(n22993) );
  XNOR U22392 ( .A(n23002), .B(n23003), .Z(n22991) );
  AND U22393 ( .A(n1705), .B(n23004), .Z(n23003) );
  XOR U22394 ( .A(p_input[1388]), .B(n23002), .Z(n23004) );
  XNOR U22395 ( .A(n23005), .B(n23006), .Z(n23002) );
  AND U22396 ( .A(n1709), .B(n23007), .Z(n23006) );
  XOR U22397 ( .A(n23008), .B(n23009), .Z(n23000) );
  AND U22398 ( .A(n1713), .B(n22999), .Z(n23009) );
  XNOR U22399 ( .A(n23010), .B(n22997), .Z(n22999) );
  XOR U22400 ( .A(n23011), .B(n23012), .Z(n22997) );
  AND U22401 ( .A(n1736), .B(n23013), .Z(n23012) );
  IV U22402 ( .A(n23008), .Z(n23010) );
  XOR U22403 ( .A(n23014), .B(n23015), .Z(n23008) );
  AND U22404 ( .A(n1720), .B(n23007), .Z(n23015) );
  XNOR U22405 ( .A(n23005), .B(n23014), .Z(n23007) );
  XNOR U22406 ( .A(n23016), .B(n23017), .Z(n23005) );
  AND U22407 ( .A(n1724), .B(n23018), .Z(n23017) );
  XOR U22408 ( .A(p_input[1404]), .B(n23016), .Z(n23018) );
  XNOR U22409 ( .A(n23019), .B(n23020), .Z(n23016) );
  AND U22410 ( .A(n1728), .B(n23021), .Z(n23020) );
  XOR U22411 ( .A(n23022), .B(n23023), .Z(n23014) );
  AND U22412 ( .A(n1732), .B(n23013), .Z(n23023) );
  XNOR U22413 ( .A(n23024), .B(n23011), .Z(n23013) );
  XOR U22414 ( .A(n23025), .B(n23026), .Z(n23011) );
  AND U22415 ( .A(n1755), .B(n23027), .Z(n23026) );
  IV U22416 ( .A(n23022), .Z(n23024) );
  XOR U22417 ( .A(n23028), .B(n23029), .Z(n23022) );
  AND U22418 ( .A(n1739), .B(n23021), .Z(n23029) );
  XNOR U22419 ( .A(n23019), .B(n23028), .Z(n23021) );
  XNOR U22420 ( .A(n23030), .B(n23031), .Z(n23019) );
  AND U22421 ( .A(n1743), .B(n23032), .Z(n23031) );
  XOR U22422 ( .A(p_input[1420]), .B(n23030), .Z(n23032) );
  XNOR U22423 ( .A(n23033), .B(n23034), .Z(n23030) );
  AND U22424 ( .A(n1747), .B(n23035), .Z(n23034) );
  XOR U22425 ( .A(n23036), .B(n23037), .Z(n23028) );
  AND U22426 ( .A(n1751), .B(n23027), .Z(n23037) );
  XNOR U22427 ( .A(n23038), .B(n23025), .Z(n23027) );
  XOR U22428 ( .A(n23039), .B(n23040), .Z(n23025) );
  AND U22429 ( .A(n1774), .B(n23041), .Z(n23040) );
  IV U22430 ( .A(n23036), .Z(n23038) );
  XOR U22431 ( .A(n23042), .B(n23043), .Z(n23036) );
  AND U22432 ( .A(n1758), .B(n23035), .Z(n23043) );
  XNOR U22433 ( .A(n23033), .B(n23042), .Z(n23035) );
  XNOR U22434 ( .A(n23044), .B(n23045), .Z(n23033) );
  AND U22435 ( .A(n1762), .B(n23046), .Z(n23045) );
  XOR U22436 ( .A(p_input[1436]), .B(n23044), .Z(n23046) );
  XNOR U22437 ( .A(n23047), .B(n23048), .Z(n23044) );
  AND U22438 ( .A(n1766), .B(n23049), .Z(n23048) );
  XOR U22439 ( .A(n23050), .B(n23051), .Z(n23042) );
  AND U22440 ( .A(n1770), .B(n23041), .Z(n23051) );
  XNOR U22441 ( .A(n23052), .B(n23039), .Z(n23041) );
  XOR U22442 ( .A(n23053), .B(n23054), .Z(n23039) );
  AND U22443 ( .A(n1793), .B(n23055), .Z(n23054) );
  IV U22444 ( .A(n23050), .Z(n23052) );
  XOR U22445 ( .A(n23056), .B(n23057), .Z(n23050) );
  AND U22446 ( .A(n1777), .B(n23049), .Z(n23057) );
  XNOR U22447 ( .A(n23047), .B(n23056), .Z(n23049) );
  XNOR U22448 ( .A(n23058), .B(n23059), .Z(n23047) );
  AND U22449 ( .A(n1781), .B(n23060), .Z(n23059) );
  XOR U22450 ( .A(p_input[1452]), .B(n23058), .Z(n23060) );
  XNOR U22451 ( .A(n23061), .B(n23062), .Z(n23058) );
  AND U22452 ( .A(n1785), .B(n23063), .Z(n23062) );
  XOR U22453 ( .A(n23064), .B(n23065), .Z(n23056) );
  AND U22454 ( .A(n1789), .B(n23055), .Z(n23065) );
  XNOR U22455 ( .A(n23066), .B(n23053), .Z(n23055) );
  XOR U22456 ( .A(n23067), .B(n23068), .Z(n23053) );
  AND U22457 ( .A(n1812), .B(n23069), .Z(n23068) );
  IV U22458 ( .A(n23064), .Z(n23066) );
  XOR U22459 ( .A(n23070), .B(n23071), .Z(n23064) );
  AND U22460 ( .A(n1796), .B(n23063), .Z(n23071) );
  XNOR U22461 ( .A(n23061), .B(n23070), .Z(n23063) );
  XNOR U22462 ( .A(n23072), .B(n23073), .Z(n23061) );
  AND U22463 ( .A(n1800), .B(n23074), .Z(n23073) );
  XOR U22464 ( .A(p_input[1468]), .B(n23072), .Z(n23074) );
  XNOR U22465 ( .A(n23075), .B(n23076), .Z(n23072) );
  AND U22466 ( .A(n1804), .B(n23077), .Z(n23076) );
  XOR U22467 ( .A(n23078), .B(n23079), .Z(n23070) );
  AND U22468 ( .A(n1808), .B(n23069), .Z(n23079) );
  XNOR U22469 ( .A(n23080), .B(n23067), .Z(n23069) );
  XOR U22470 ( .A(n23081), .B(n23082), .Z(n23067) );
  AND U22471 ( .A(n1831), .B(n23083), .Z(n23082) );
  IV U22472 ( .A(n23078), .Z(n23080) );
  XOR U22473 ( .A(n23084), .B(n23085), .Z(n23078) );
  AND U22474 ( .A(n1815), .B(n23077), .Z(n23085) );
  XNOR U22475 ( .A(n23075), .B(n23084), .Z(n23077) );
  XNOR U22476 ( .A(n23086), .B(n23087), .Z(n23075) );
  AND U22477 ( .A(n1819), .B(n23088), .Z(n23087) );
  XOR U22478 ( .A(p_input[1484]), .B(n23086), .Z(n23088) );
  XNOR U22479 ( .A(n23089), .B(n23090), .Z(n23086) );
  AND U22480 ( .A(n1823), .B(n23091), .Z(n23090) );
  XOR U22481 ( .A(n23092), .B(n23093), .Z(n23084) );
  AND U22482 ( .A(n1827), .B(n23083), .Z(n23093) );
  XNOR U22483 ( .A(n23094), .B(n23081), .Z(n23083) );
  XOR U22484 ( .A(n23095), .B(n23096), .Z(n23081) );
  AND U22485 ( .A(n1850), .B(n23097), .Z(n23096) );
  IV U22486 ( .A(n23092), .Z(n23094) );
  XOR U22487 ( .A(n23098), .B(n23099), .Z(n23092) );
  AND U22488 ( .A(n1834), .B(n23091), .Z(n23099) );
  XNOR U22489 ( .A(n23089), .B(n23098), .Z(n23091) );
  XNOR U22490 ( .A(n23100), .B(n23101), .Z(n23089) );
  AND U22491 ( .A(n1838), .B(n23102), .Z(n23101) );
  XOR U22492 ( .A(p_input[1500]), .B(n23100), .Z(n23102) );
  XNOR U22493 ( .A(n23103), .B(n23104), .Z(n23100) );
  AND U22494 ( .A(n1842), .B(n23105), .Z(n23104) );
  XOR U22495 ( .A(n23106), .B(n23107), .Z(n23098) );
  AND U22496 ( .A(n1846), .B(n23097), .Z(n23107) );
  XNOR U22497 ( .A(n23108), .B(n23095), .Z(n23097) );
  XOR U22498 ( .A(n23109), .B(n23110), .Z(n23095) );
  AND U22499 ( .A(n1869), .B(n23111), .Z(n23110) );
  IV U22500 ( .A(n23106), .Z(n23108) );
  XOR U22501 ( .A(n23112), .B(n23113), .Z(n23106) );
  AND U22502 ( .A(n1853), .B(n23105), .Z(n23113) );
  XNOR U22503 ( .A(n23103), .B(n23112), .Z(n23105) );
  XNOR U22504 ( .A(n23114), .B(n23115), .Z(n23103) );
  AND U22505 ( .A(n1857), .B(n23116), .Z(n23115) );
  XOR U22506 ( .A(p_input[1516]), .B(n23114), .Z(n23116) );
  XNOR U22507 ( .A(n23117), .B(n23118), .Z(n23114) );
  AND U22508 ( .A(n1861), .B(n23119), .Z(n23118) );
  XOR U22509 ( .A(n23120), .B(n23121), .Z(n23112) );
  AND U22510 ( .A(n1865), .B(n23111), .Z(n23121) );
  XNOR U22511 ( .A(n23122), .B(n23109), .Z(n23111) );
  XOR U22512 ( .A(n23123), .B(n23124), .Z(n23109) );
  AND U22513 ( .A(n1888), .B(n23125), .Z(n23124) );
  IV U22514 ( .A(n23120), .Z(n23122) );
  XOR U22515 ( .A(n23126), .B(n23127), .Z(n23120) );
  AND U22516 ( .A(n1872), .B(n23119), .Z(n23127) );
  XNOR U22517 ( .A(n23117), .B(n23126), .Z(n23119) );
  XNOR U22518 ( .A(n23128), .B(n23129), .Z(n23117) );
  AND U22519 ( .A(n1876), .B(n23130), .Z(n23129) );
  XOR U22520 ( .A(p_input[1532]), .B(n23128), .Z(n23130) );
  XNOR U22521 ( .A(n23131), .B(n23132), .Z(n23128) );
  AND U22522 ( .A(n1880), .B(n23133), .Z(n23132) );
  XOR U22523 ( .A(n23134), .B(n23135), .Z(n23126) );
  AND U22524 ( .A(n1884), .B(n23125), .Z(n23135) );
  XNOR U22525 ( .A(n23136), .B(n23123), .Z(n23125) );
  XOR U22526 ( .A(n23137), .B(n23138), .Z(n23123) );
  AND U22527 ( .A(n1907), .B(n23139), .Z(n23138) );
  IV U22528 ( .A(n23134), .Z(n23136) );
  XOR U22529 ( .A(n23140), .B(n23141), .Z(n23134) );
  AND U22530 ( .A(n1891), .B(n23133), .Z(n23141) );
  XNOR U22531 ( .A(n23131), .B(n23140), .Z(n23133) );
  XNOR U22532 ( .A(n23142), .B(n23143), .Z(n23131) );
  AND U22533 ( .A(n1895), .B(n23144), .Z(n23143) );
  XOR U22534 ( .A(p_input[1548]), .B(n23142), .Z(n23144) );
  XNOR U22535 ( .A(n23145), .B(n23146), .Z(n23142) );
  AND U22536 ( .A(n1899), .B(n23147), .Z(n23146) );
  XOR U22537 ( .A(n23148), .B(n23149), .Z(n23140) );
  AND U22538 ( .A(n1903), .B(n23139), .Z(n23149) );
  XNOR U22539 ( .A(n23150), .B(n23137), .Z(n23139) );
  XOR U22540 ( .A(n23151), .B(n23152), .Z(n23137) );
  AND U22541 ( .A(n1926), .B(n23153), .Z(n23152) );
  IV U22542 ( .A(n23148), .Z(n23150) );
  XOR U22543 ( .A(n23154), .B(n23155), .Z(n23148) );
  AND U22544 ( .A(n1910), .B(n23147), .Z(n23155) );
  XNOR U22545 ( .A(n23145), .B(n23154), .Z(n23147) );
  XNOR U22546 ( .A(n23156), .B(n23157), .Z(n23145) );
  AND U22547 ( .A(n1914), .B(n23158), .Z(n23157) );
  XOR U22548 ( .A(p_input[1564]), .B(n23156), .Z(n23158) );
  XNOR U22549 ( .A(n23159), .B(n23160), .Z(n23156) );
  AND U22550 ( .A(n1918), .B(n23161), .Z(n23160) );
  XOR U22551 ( .A(n23162), .B(n23163), .Z(n23154) );
  AND U22552 ( .A(n1922), .B(n23153), .Z(n23163) );
  XNOR U22553 ( .A(n23164), .B(n23151), .Z(n23153) );
  XOR U22554 ( .A(n23165), .B(n23166), .Z(n23151) );
  AND U22555 ( .A(n1945), .B(n23167), .Z(n23166) );
  IV U22556 ( .A(n23162), .Z(n23164) );
  XOR U22557 ( .A(n23168), .B(n23169), .Z(n23162) );
  AND U22558 ( .A(n1929), .B(n23161), .Z(n23169) );
  XNOR U22559 ( .A(n23159), .B(n23168), .Z(n23161) );
  XNOR U22560 ( .A(n23170), .B(n23171), .Z(n23159) );
  AND U22561 ( .A(n1933), .B(n23172), .Z(n23171) );
  XOR U22562 ( .A(p_input[1580]), .B(n23170), .Z(n23172) );
  XNOR U22563 ( .A(n23173), .B(n23174), .Z(n23170) );
  AND U22564 ( .A(n1937), .B(n23175), .Z(n23174) );
  XOR U22565 ( .A(n23176), .B(n23177), .Z(n23168) );
  AND U22566 ( .A(n1941), .B(n23167), .Z(n23177) );
  XNOR U22567 ( .A(n23178), .B(n23165), .Z(n23167) );
  XOR U22568 ( .A(n23179), .B(n23180), .Z(n23165) );
  AND U22569 ( .A(n1964), .B(n23181), .Z(n23180) );
  IV U22570 ( .A(n23176), .Z(n23178) );
  XOR U22571 ( .A(n23182), .B(n23183), .Z(n23176) );
  AND U22572 ( .A(n1948), .B(n23175), .Z(n23183) );
  XNOR U22573 ( .A(n23173), .B(n23182), .Z(n23175) );
  XNOR U22574 ( .A(n23184), .B(n23185), .Z(n23173) );
  AND U22575 ( .A(n1952), .B(n23186), .Z(n23185) );
  XOR U22576 ( .A(p_input[1596]), .B(n23184), .Z(n23186) );
  XNOR U22577 ( .A(n23187), .B(n23188), .Z(n23184) );
  AND U22578 ( .A(n1956), .B(n23189), .Z(n23188) );
  XOR U22579 ( .A(n23190), .B(n23191), .Z(n23182) );
  AND U22580 ( .A(n1960), .B(n23181), .Z(n23191) );
  XNOR U22581 ( .A(n23192), .B(n23179), .Z(n23181) );
  XOR U22582 ( .A(n23193), .B(n23194), .Z(n23179) );
  AND U22583 ( .A(n1983), .B(n23195), .Z(n23194) );
  IV U22584 ( .A(n23190), .Z(n23192) );
  XOR U22585 ( .A(n23196), .B(n23197), .Z(n23190) );
  AND U22586 ( .A(n1967), .B(n23189), .Z(n23197) );
  XNOR U22587 ( .A(n23187), .B(n23196), .Z(n23189) );
  XNOR U22588 ( .A(n23198), .B(n23199), .Z(n23187) );
  AND U22589 ( .A(n1971), .B(n23200), .Z(n23199) );
  XOR U22590 ( .A(p_input[1612]), .B(n23198), .Z(n23200) );
  XNOR U22591 ( .A(n23201), .B(n23202), .Z(n23198) );
  AND U22592 ( .A(n1975), .B(n23203), .Z(n23202) );
  XOR U22593 ( .A(n23204), .B(n23205), .Z(n23196) );
  AND U22594 ( .A(n1979), .B(n23195), .Z(n23205) );
  XNOR U22595 ( .A(n23206), .B(n23193), .Z(n23195) );
  XOR U22596 ( .A(n23207), .B(n23208), .Z(n23193) );
  AND U22597 ( .A(n2002), .B(n23209), .Z(n23208) );
  IV U22598 ( .A(n23204), .Z(n23206) );
  XOR U22599 ( .A(n23210), .B(n23211), .Z(n23204) );
  AND U22600 ( .A(n1986), .B(n23203), .Z(n23211) );
  XNOR U22601 ( .A(n23201), .B(n23210), .Z(n23203) );
  XNOR U22602 ( .A(n23212), .B(n23213), .Z(n23201) );
  AND U22603 ( .A(n1990), .B(n23214), .Z(n23213) );
  XOR U22604 ( .A(p_input[1628]), .B(n23212), .Z(n23214) );
  XNOR U22605 ( .A(n23215), .B(n23216), .Z(n23212) );
  AND U22606 ( .A(n1994), .B(n23217), .Z(n23216) );
  XOR U22607 ( .A(n23218), .B(n23219), .Z(n23210) );
  AND U22608 ( .A(n1998), .B(n23209), .Z(n23219) );
  XNOR U22609 ( .A(n23220), .B(n23207), .Z(n23209) );
  XOR U22610 ( .A(n23221), .B(n23222), .Z(n23207) );
  AND U22611 ( .A(n2021), .B(n23223), .Z(n23222) );
  IV U22612 ( .A(n23218), .Z(n23220) );
  XOR U22613 ( .A(n23224), .B(n23225), .Z(n23218) );
  AND U22614 ( .A(n2005), .B(n23217), .Z(n23225) );
  XNOR U22615 ( .A(n23215), .B(n23224), .Z(n23217) );
  XNOR U22616 ( .A(n23226), .B(n23227), .Z(n23215) );
  AND U22617 ( .A(n2009), .B(n23228), .Z(n23227) );
  XOR U22618 ( .A(p_input[1644]), .B(n23226), .Z(n23228) );
  XNOR U22619 ( .A(n23229), .B(n23230), .Z(n23226) );
  AND U22620 ( .A(n2013), .B(n23231), .Z(n23230) );
  XOR U22621 ( .A(n23232), .B(n23233), .Z(n23224) );
  AND U22622 ( .A(n2017), .B(n23223), .Z(n23233) );
  XNOR U22623 ( .A(n23234), .B(n23221), .Z(n23223) );
  XOR U22624 ( .A(n23235), .B(n23236), .Z(n23221) );
  AND U22625 ( .A(n2040), .B(n23237), .Z(n23236) );
  IV U22626 ( .A(n23232), .Z(n23234) );
  XOR U22627 ( .A(n23238), .B(n23239), .Z(n23232) );
  AND U22628 ( .A(n2024), .B(n23231), .Z(n23239) );
  XNOR U22629 ( .A(n23229), .B(n23238), .Z(n23231) );
  XNOR U22630 ( .A(n23240), .B(n23241), .Z(n23229) );
  AND U22631 ( .A(n2028), .B(n23242), .Z(n23241) );
  XOR U22632 ( .A(p_input[1660]), .B(n23240), .Z(n23242) );
  XNOR U22633 ( .A(n23243), .B(n23244), .Z(n23240) );
  AND U22634 ( .A(n2032), .B(n23245), .Z(n23244) );
  XOR U22635 ( .A(n23246), .B(n23247), .Z(n23238) );
  AND U22636 ( .A(n2036), .B(n23237), .Z(n23247) );
  XNOR U22637 ( .A(n23248), .B(n23235), .Z(n23237) );
  XOR U22638 ( .A(n23249), .B(n23250), .Z(n23235) );
  AND U22639 ( .A(n2059), .B(n23251), .Z(n23250) );
  IV U22640 ( .A(n23246), .Z(n23248) );
  XOR U22641 ( .A(n23252), .B(n23253), .Z(n23246) );
  AND U22642 ( .A(n2043), .B(n23245), .Z(n23253) );
  XNOR U22643 ( .A(n23243), .B(n23252), .Z(n23245) );
  XNOR U22644 ( .A(n23254), .B(n23255), .Z(n23243) );
  AND U22645 ( .A(n2047), .B(n23256), .Z(n23255) );
  XOR U22646 ( .A(p_input[1676]), .B(n23254), .Z(n23256) );
  XNOR U22647 ( .A(n23257), .B(n23258), .Z(n23254) );
  AND U22648 ( .A(n2051), .B(n23259), .Z(n23258) );
  XOR U22649 ( .A(n23260), .B(n23261), .Z(n23252) );
  AND U22650 ( .A(n2055), .B(n23251), .Z(n23261) );
  XNOR U22651 ( .A(n23262), .B(n23249), .Z(n23251) );
  XOR U22652 ( .A(n23263), .B(n23264), .Z(n23249) );
  AND U22653 ( .A(n2078), .B(n23265), .Z(n23264) );
  IV U22654 ( .A(n23260), .Z(n23262) );
  XOR U22655 ( .A(n23266), .B(n23267), .Z(n23260) );
  AND U22656 ( .A(n2062), .B(n23259), .Z(n23267) );
  XNOR U22657 ( .A(n23257), .B(n23266), .Z(n23259) );
  XNOR U22658 ( .A(n23268), .B(n23269), .Z(n23257) );
  AND U22659 ( .A(n2066), .B(n23270), .Z(n23269) );
  XOR U22660 ( .A(p_input[1692]), .B(n23268), .Z(n23270) );
  XNOR U22661 ( .A(n23271), .B(n23272), .Z(n23268) );
  AND U22662 ( .A(n2070), .B(n23273), .Z(n23272) );
  XOR U22663 ( .A(n23274), .B(n23275), .Z(n23266) );
  AND U22664 ( .A(n2074), .B(n23265), .Z(n23275) );
  XNOR U22665 ( .A(n23276), .B(n23263), .Z(n23265) );
  XOR U22666 ( .A(n23277), .B(n23278), .Z(n23263) );
  AND U22667 ( .A(n2097), .B(n23279), .Z(n23278) );
  IV U22668 ( .A(n23274), .Z(n23276) );
  XOR U22669 ( .A(n23280), .B(n23281), .Z(n23274) );
  AND U22670 ( .A(n2081), .B(n23273), .Z(n23281) );
  XNOR U22671 ( .A(n23271), .B(n23280), .Z(n23273) );
  XNOR U22672 ( .A(n23282), .B(n23283), .Z(n23271) );
  AND U22673 ( .A(n2085), .B(n23284), .Z(n23283) );
  XOR U22674 ( .A(p_input[1708]), .B(n23282), .Z(n23284) );
  XNOR U22675 ( .A(n23285), .B(n23286), .Z(n23282) );
  AND U22676 ( .A(n2089), .B(n23287), .Z(n23286) );
  XOR U22677 ( .A(n23288), .B(n23289), .Z(n23280) );
  AND U22678 ( .A(n2093), .B(n23279), .Z(n23289) );
  XNOR U22679 ( .A(n23290), .B(n23277), .Z(n23279) );
  XOR U22680 ( .A(n23291), .B(n23292), .Z(n23277) );
  AND U22681 ( .A(n2116), .B(n23293), .Z(n23292) );
  IV U22682 ( .A(n23288), .Z(n23290) );
  XOR U22683 ( .A(n23294), .B(n23295), .Z(n23288) );
  AND U22684 ( .A(n2100), .B(n23287), .Z(n23295) );
  XNOR U22685 ( .A(n23285), .B(n23294), .Z(n23287) );
  XNOR U22686 ( .A(n23296), .B(n23297), .Z(n23285) );
  AND U22687 ( .A(n2104), .B(n23298), .Z(n23297) );
  XOR U22688 ( .A(p_input[1724]), .B(n23296), .Z(n23298) );
  XNOR U22689 ( .A(n23299), .B(n23300), .Z(n23296) );
  AND U22690 ( .A(n2108), .B(n23301), .Z(n23300) );
  XOR U22691 ( .A(n23302), .B(n23303), .Z(n23294) );
  AND U22692 ( .A(n2112), .B(n23293), .Z(n23303) );
  XNOR U22693 ( .A(n23304), .B(n23291), .Z(n23293) );
  XOR U22694 ( .A(n23305), .B(n23306), .Z(n23291) );
  AND U22695 ( .A(n2135), .B(n23307), .Z(n23306) );
  IV U22696 ( .A(n23302), .Z(n23304) );
  XOR U22697 ( .A(n23308), .B(n23309), .Z(n23302) );
  AND U22698 ( .A(n2119), .B(n23301), .Z(n23309) );
  XNOR U22699 ( .A(n23299), .B(n23308), .Z(n23301) );
  XNOR U22700 ( .A(n23310), .B(n23311), .Z(n23299) );
  AND U22701 ( .A(n2123), .B(n23312), .Z(n23311) );
  XOR U22702 ( .A(p_input[1740]), .B(n23310), .Z(n23312) );
  XNOR U22703 ( .A(n23313), .B(n23314), .Z(n23310) );
  AND U22704 ( .A(n2127), .B(n23315), .Z(n23314) );
  XOR U22705 ( .A(n23316), .B(n23317), .Z(n23308) );
  AND U22706 ( .A(n2131), .B(n23307), .Z(n23317) );
  XNOR U22707 ( .A(n23318), .B(n23305), .Z(n23307) );
  XOR U22708 ( .A(n23319), .B(n23320), .Z(n23305) );
  AND U22709 ( .A(n2154), .B(n23321), .Z(n23320) );
  IV U22710 ( .A(n23316), .Z(n23318) );
  XOR U22711 ( .A(n23322), .B(n23323), .Z(n23316) );
  AND U22712 ( .A(n2138), .B(n23315), .Z(n23323) );
  XNOR U22713 ( .A(n23313), .B(n23322), .Z(n23315) );
  XNOR U22714 ( .A(n23324), .B(n23325), .Z(n23313) );
  AND U22715 ( .A(n2142), .B(n23326), .Z(n23325) );
  XOR U22716 ( .A(p_input[1756]), .B(n23324), .Z(n23326) );
  XNOR U22717 ( .A(n23327), .B(n23328), .Z(n23324) );
  AND U22718 ( .A(n2146), .B(n23329), .Z(n23328) );
  XOR U22719 ( .A(n23330), .B(n23331), .Z(n23322) );
  AND U22720 ( .A(n2150), .B(n23321), .Z(n23331) );
  XNOR U22721 ( .A(n23332), .B(n23319), .Z(n23321) );
  XOR U22722 ( .A(n23333), .B(n23334), .Z(n23319) );
  AND U22723 ( .A(n2173), .B(n23335), .Z(n23334) );
  IV U22724 ( .A(n23330), .Z(n23332) );
  XOR U22725 ( .A(n23336), .B(n23337), .Z(n23330) );
  AND U22726 ( .A(n2157), .B(n23329), .Z(n23337) );
  XNOR U22727 ( .A(n23327), .B(n23336), .Z(n23329) );
  XNOR U22728 ( .A(n23338), .B(n23339), .Z(n23327) );
  AND U22729 ( .A(n2161), .B(n23340), .Z(n23339) );
  XOR U22730 ( .A(p_input[1772]), .B(n23338), .Z(n23340) );
  XNOR U22731 ( .A(n23341), .B(n23342), .Z(n23338) );
  AND U22732 ( .A(n2165), .B(n23343), .Z(n23342) );
  XOR U22733 ( .A(n23344), .B(n23345), .Z(n23336) );
  AND U22734 ( .A(n2169), .B(n23335), .Z(n23345) );
  XNOR U22735 ( .A(n23346), .B(n23333), .Z(n23335) );
  XOR U22736 ( .A(n23347), .B(n23348), .Z(n23333) );
  AND U22737 ( .A(n2192), .B(n23349), .Z(n23348) );
  IV U22738 ( .A(n23344), .Z(n23346) );
  XOR U22739 ( .A(n23350), .B(n23351), .Z(n23344) );
  AND U22740 ( .A(n2176), .B(n23343), .Z(n23351) );
  XNOR U22741 ( .A(n23341), .B(n23350), .Z(n23343) );
  XNOR U22742 ( .A(n23352), .B(n23353), .Z(n23341) );
  AND U22743 ( .A(n2180), .B(n23354), .Z(n23353) );
  XOR U22744 ( .A(p_input[1788]), .B(n23352), .Z(n23354) );
  XNOR U22745 ( .A(n23355), .B(n23356), .Z(n23352) );
  AND U22746 ( .A(n2184), .B(n23357), .Z(n23356) );
  XOR U22747 ( .A(n23358), .B(n23359), .Z(n23350) );
  AND U22748 ( .A(n2188), .B(n23349), .Z(n23359) );
  XNOR U22749 ( .A(n23360), .B(n23347), .Z(n23349) );
  XOR U22750 ( .A(n23361), .B(n23362), .Z(n23347) );
  AND U22751 ( .A(n2211), .B(n23363), .Z(n23362) );
  IV U22752 ( .A(n23358), .Z(n23360) );
  XOR U22753 ( .A(n23364), .B(n23365), .Z(n23358) );
  AND U22754 ( .A(n2195), .B(n23357), .Z(n23365) );
  XNOR U22755 ( .A(n23355), .B(n23364), .Z(n23357) );
  XNOR U22756 ( .A(n23366), .B(n23367), .Z(n23355) );
  AND U22757 ( .A(n2199), .B(n23368), .Z(n23367) );
  XOR U22758 ( .A(p_input[1804]), .B(n23366), .Z(n23368) );
  XNOR U22759 ( .A(n23369), .B(n23370), .Z(n23366) );
  AND U22760 ( .A(n2203), .B(n23371), .Z(n23370) );
  XOR U22761 ( .A(n23372), .B(n23373), .Z(n23364) );
  AND U22762 ( .A(n2207), .B(n23363), .Z(n23373) );
  XNOR U22763 ( .A(n23374), .B(n23361), .Z(n23363) );
  XOR U22764 ( .A(n23375), .B(n23376), .Z(n23361) );
  AND U22765 ( .A(n2230), .B(n23377), .Z(n23376) );
  IV U22766 ( .A(n23372), .Z(n23374) );
  XOR U22767 ( .A(n23378), .B(n23379), .Z(n23372) );
  AND U22768 ( .A(n2214), .B(n23371), .Z(n23379) );
  XNOR U22769 ( .A(n23369), .B(n23378), .Z(n23371) );
  XNOR U22770 ( .A(n23380), .B(n23381), .Z(n23369) );
  AND U22771 ( .A(n2218), .B(n23382), .Z(n23381) );
  XOR U22772 ( .A(p_input[1820]), .B(n23380), .Z(n23382) );
  XNOR U22773 ( .A(n23383), .B(n23384), .Z(n23380) );
  AND U22774 ( .A(n2222), .B(n23385), .Z(n23384) );
  XOR U22775 ( .A(n23386), .B(n23387), .Z(n23378) );
  AND U22776 ( .A(n2226), .B(n23377), .Z(n23387) );
  XNOR U22777 ( .A(n23388), .B(n23375), .Z(n23377) );
  XOR U22778 ( .A(n23389), .B(n23390), .Z(n23375) );
  AND U22779 ( .A(n2249), .B(n23391), .Z(n23390) );
  IV U22780 ( .A(n23386), .Z(n23388) );
  XOR U22781 ( .A(n23392), .B(n23393), .Z(n23386) );
  AND U22782 ( .A(n2233), .B(n23385), .Z(n23393) );
  XNOR U22783 ( .A(n23383), .B(n23392), .Z(n23385) );
  XNOR U22784 ( .A(n23394), .B(n23395), .Z(n23383) );
  AND U22785 ( .A(n2237), .B(n23396), .Z(n23395) );
  XOR U22786 ( .A(p_input[1836]), .B(n23394), .Z(n23396) );
  XNOR U22787 ( .A(n23397), .B(n23398), .Z(n23394) );
  AND U22788 ( .A(n2241), .B(n23399), .Z(n23398) );
  XOR U22789 ( .A(n23400), .B(n23401), .Z(n23392) );
  AND U22790 ( .A(n2245), .B(n23391), .Z(n23401) );
  XNOR U22791 ( .A(n23402), .B(n23389), .Z(n23391) );
  XOR U22792 ( .A(n23403), .B(n23404), .Z(n23389) );
  AND U22793 ( .A(n2268), .B(n23405), .Z(n23404) );
  IV U22794 ( .A(n23400), .Z(n23402) );
  XOR U22795 ( .A(n23406), .B(n23407), .Z(n23400) );
  AND U22796 ( .A(n2252), .B(n23399), .Z(n23407) );
  XNOR U22797 ( .A(n23397), .B(n23406), .Z(n23399) );
  XNOR U22798 ( .A(n23408), .B(n23409), .Z(n23397) );
  AND U22799 ( .A(n2256), .B(n23410), .Z(n23409) );
  XOR U22800 ( .A(p_input[1852]), .B(n23408), .Z(n23410) );
  XNOR U22801 ( .A(n23411), .B(n23412), .Z(n23408) );
  AND U22802 ( .A(n2260), .B(n23413), .Z(n23412) );
  XOR U22803 ( .A(n23414), .B(n23415), .Z(n23406) );
  AND U22804 ( .A(n2264), .B(n23405), .Z(n23415) );
  XNOR U22805 ( .A(n23416), .B(n23403), .Z(n23405) );
  XOR U22806 ( .A(n23417), .B(n23418), .Z(n23403) );
  AND U22807 ( .A(n2287), .B(n23419), .Z(n23418) );
  IV U22808 ( .A(n23414), .Z(n23416) );
  XOR U22809 ( .A(n23420), .B(n23421), .Z(n23414) );
  AND U22810 ( .A(n2271), .B(n23413), .Z(n23421) );
  XNOR U22811 ( .A(n23411), .B(n23420), .Z(n23413) );
  XNOR U22812 ( .A(n23422), .B(n23423), .Z(n23411) );
  AND U22813 ( .A(n2275), .B(n23424), .Z(n23423) );
  XOR U22814 ( .A(p_input[1868]), .B(n23422), .Z(n23424) );
  XNOR U22815 ( .A(n23425), .B(n23426), .Z(n23422) );
  AND U22816 ( .A(n2279), .B(n23427), .Z(n23426) );
  XOR U22817 ( .A(n23428), .B(n23429), .Z(n23420) );
  AND U22818 ( .A(n2283), .B(n23419), .Z(n23429) );
  XNOR U22819 ( .A(n23430), .B(n23417), .Z(n23419) );
  XOR U22820 ( .A(n23431), .B(n23432), .Z(n23417) );
  AND U22821 ( .A(n2306), .B(n23433), .Z(n23432) );
  IV U22822 ( .A(n23428), .Z(n23430) );
  XOR U22823 ( .A(n23434), .B(n23435), .Z(n23428) );
  AND U22824 ( .A(n2290), .B(n23427), .Z(n23435) );
  XNOR U22825 ( .A(n23425), .B(n23434), .Z(n23427) );
  XNOR U22826 ( .A(n23436), .B(n23437), .Z(n23425) );
  AND U22827 ( .A(n2294), .B(n23438), .Z(n23437) );
  XOR U22828 ( .A(p_input[1884]), .B(n23436), .Z(n23438) );
  XNOR U22829 ( .A(n23439), .B(n23440), .Z(n23436) );
  AND U22830 ( .A(n2298), .B(n23441), .Z(n23440) );
  XOR U22831 ( .A(n23442), .B(n23443), .Z(n23434) );
  AND U22832 ( .A(n2302), .B(n23433), .Z(n23443) );
  XNOR U22833 ( .A(n23444), .B(n23431), .Z(n23433) );
  XOR U22834 ( .A(n23445), .B(n23446), .Z(n23431) );
  AND U22835 ( .A(n2325), .B(n23447), .Z(n23446) );
  IV U22836 ( .A(n23442), .Z(n23444) );
  XOR U22837 ( .A(n23448), .B(n23449), .Z(n23442) );
  AND U22838 ( .A(n2309), .B(n23441), .Z(n23449) );
  XNOR U22839 ( .A(n23439), .B(n23448), .Z(n23441) );
  XNOR U22840 ( .A(n23450), .B(n23451), .Z(n23439) );
  AND U22841 ( .A(n2313), .B(n23452), .Z(n23451) );
  XOR U22842 ( .A(p_input[1900]), .B(n23450), .Z(n23452) );
  XNOR U22843 ( .A(n23453), .B(n23454), .Z(n23450) );
  AND U22844 ( .A(n2317), .B(n23455), .Z(n23454) );
  XOR U22845 ( .A(n23456), .B(n23457), .Z(n23448) );
  AND U22846 ( .A(n2321), .B(n23447), .Z(n23457) );
  XNOR U22847 ( .A(n23458), .B(n23445), .Z(n23447) );
  XOR U22848 ( .A(n23459), .B(n23460), .Z(n23445) );
  AND U22849 ( .A(n2344), .B(n23461), .Z(n23460) );
  IV U22850 ( .A(n23456), .Z(n23458) );
  XOR U22851 ( .A(n23462), .B(n23463), .Z(n23456) );
  AND U22852 ( .A(n2328), .B(n23455), .Z(n23463) );
  XNOR U22853 ( .A(n23453), .B(n23462), .Z(n23455) );
  XNOR U22854 ( .A(n23464), .B(n23465), .Z(n23453) );
  AND U22855 ( .A(n2332), .B(n23466), .Z(n23465) );
  XOR U22856 ( .A(p_input[1916]), .B(n23464), .Z(n23466) );
  XNOR U22857 ( .A(n23467), .B(n23468), .Z(n23464) );
  AND U22858 ( .A(n2336), .B(n23469), .Z(n23468) );
  XOR U22859 ( .A(n23470), .B(n23471), .Z(n23462) );
  AND U22860 ( .A(n2340), .B(n23461), .Z(n23471) );
  XNOR U22861 ( .A(n23472), .B(n23459), .Z(n23461) );
  XOR U22862 ( .A(n23473), .B(n23474), .Z(n23459) );
  AND U22863 ( .A(n2363), .B(n23475), .Z(n23474) );
  IV U22864 ( .A(n23470), .Z(n23472) );
  XOR U22865 ( .A(n23476), .B(n23477), .Z(n23470) );
  AND U22866 ( .A(n2347), .B(n23469), .Z(n23477) );
  XNOR U22867 ( .A(n23467), .B(n23476), .Z(n23469) );
  XNOR U22868 ( .A(n23478), .B(n23479), .Z(n23467) );
  AND U22869 ( .A(n2351), .B(n23480), .Z(n23479) );
  XOR U22870 ( .A(p_input[1932]), .B(n23478), .Z(n23480) );
  XNOR U22871 ( .A(n23481), .B(n23482), .Z(n23478) );
  AND U22872 ( .A(n2355), .B(n23483), .Z(n23482) );
  XOR U22873 ( .A(n23484), .B(n23485), .Z(n23476) );
  AND U22874 ( .A(n2359), .B(n23475), .Z(n23485) );
  XNOR U22875 ( .A(n23486), .B(n23473), .Z(n23475) );
  XOR U22876 ( .A(n23487), .B(n23488), .Z(n23473) );
  AND U22877 ( .A(n2382), .B(n23489), .Z(n23488) );
  IV U22878 ( .A(n23484), .Z(n23486) );
  XOR U22879 ( .A(n23490), .B(n23491), .Z(n23484) );
  AND U22880 ( .A(n2366), .B(n23483), .Z(n23491) );
  XNOR U22881 ( .A(n23481), .B(n23490), .Z(n23483) );
  XNOR U22882 ( .A(n23492), .B(n23493), .Z(n23481) );
  AND U22883 ( .A(n2370), .B(n23494), .Z(n23493) );
  XOR U22884 ( .A(p_input[1948]), .B(n23492), .Z(n23494) );
  XNOR U22885 ( .A(n23495), .B(n23496), .Z(n23492) );
  AND U22886 ( .A(n2374), .B(n23497), .Z(n23496) );
  XOR U22887 ( .A(n23498), .B(n23499), .Z(n23490) );
  AND U22888 ( .A(n2378), .B(n23489), .Z(n23499) );
  XNOR U22889 ( .A(n23500), .B(n23487), .Z(n23489) );
  XOR U22890 ( .A(n23501), .B(n23502), .Z(n23487) );
  AND U22891 ( .A(n2401), .B(n23503), .Z(n23502) );
  IV U22892 ( .A(n23498), .Z(n23500) );
  XOR U22893 ( .A(n23504), .B(n23505), .Z(n23498) );
  AND U22894 ( .A(n2385), .B(n23497), .Z(n23505) );
  XNOR U22895 ( .A(n23495), .B(n23504), .Z(n23497) );
  XNOR U22896 ( .A(n23506), .B(n23507), .Z(n23495) );
  AND U22897 ( .A(n2389), .B(n23508), .Z(n23507) );
  XOR U22898 ( .A(p_input[1964]), .B(n23506), .Z(n23508) );
  XNOR U22899 ( .A(n23509), .B(n23510), .Z(n23506) );
  AND U22900 ( .A(n2393), .B(n23511), .Z(n23510) );
  XOR U22901 ( .A(n23512), .B(n23513), .Z(n23504) );
  AND U22902 ( .A(n2397), .B(n23503), .Z(n23513) );
  XNOR U22903 ( .A(n23514), .B(n23501), .Z(n23503) );
  XOR U22904 ( .A(n23515), .B(n23516), .Z(n23501) );
  AND U22905 ( .A(n2420), .B(n23517), .Z(n23516) );
  IV U22906 ( .A(n23512), .Z(n23514) );
  XOR U22907 ( .A(n23518), .B(n23519), .Z(n23512) );
  AND U22908 ( .A(n2404), .B(n23511), .Z(n23519) );
  XNOR U22909 ( .A(n23509), .B(n23518), .Z(n23511) );
  XNOR U22910 ( .A(n23520), .B(n23521), .Z(n23509) );
  AND U22911 ( .A(n2408), .B(n23522), .Z(n23521) );
  XOR U22912 ( .A(p_input[1980]), .B(n23520), .Z(n23522) );
  XNOR U22913 ( .A(n23523), .B(n23524), .Z(n23520) );
  AND U22914 ( .A(n2412), .B(n23525), .Z(n23524) );
  XOR U22915 ( .A(n23526), .B(n23527), .Z(n23518) );
  AND U22916 ( .A(n2416), .B(n23517), .Z(n23527) );
  XNOR U22917 ( .A(n23528), .B(n23515), .Z(n23517) );
  XOR U22918 ( .A(n23529), .B(n23530), .Z(n23515) );
  AND U22919 ( .A(n2438), .B(n23531), .Z(n23530) );
  IV U22920 ( .A(n23526), .Z(n23528) );
  XOR U22921 ( .A(n23532), .B(n23533), .Z(n23526) );
  AND U22922 ( .A(n2423), .B(n23525), .Z(n23533) );
  XNOR U22923 ( .A(n23523), .B(n23532), .Z(n23525) );
  XNOR U22924 ( .A(n23534), .B(n23535), .Z(n23523) );
  AND U22925 ( .A(n2427), .B(n23536), .Z(n23535) );
  XOR U22926 ( .A(p_input[1996]), .B(n23534), .Z(n23536) );
  XOR U22927 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n23537), 
        .Z(n23534) );
  AND U22928 ( .A(n2430), .B(n23538), .Z(n23537) );
  XOR U22929 ( .A(n23539), .B(n23540), .Z(n23532) );
  AND U22930 ( .A(n2434), .B(n23531), .Z(n23540) );
  XNOR U22931 ( .A(n23541), .B(n23529), .Z(n23531) );
  XOR U22932 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n23542), .Z(n23529) );
  AND U22933 ( .A(n2446), .B(n23543), .Z(n23542) );
  IV U22934 ( .A(n23539), .Z(n23541) );
  XOR U22935 ( .A(n23544), .B(n23545), .Z(n23539) );
  AND U22936 ( .A(n2441), .B(n23538), .Z(n23545) );
  XOR U22937 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n23544), 
        .Z(n23538) );
  XOR U22938 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n23546), 
        .Z(n23544) );
  AND U22939 ( .A(n2443), .B(n23543), .Z(n23546) );
  XOR U22940 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n23543) );
  XOR U22941 ( .A(n57), .B(n23547), .Z(o[11]) );
  AND U22942 ( .A(n62), .B(n23548), .Z(n57) );
  XOR U22943 ( .A(n58), .B(n23547), .Z(n23548) );
  XOR U22944 ( .A(n23549), .B(n23550), .Z(n23547) );
  AND U22945 ( .A(n82), .B(n23551), .Z(n23550) );
  XOR U22946 ( .A(n23552), .B(n21), .Z(n58) );
  AND U22947 ( .A(n65), .B(n23553), .Z(n21) );
  XOR U22948 ( .A(n22), .B(n23552), .Z(n23553) );
  XOR U22949 ( .A(n23554), .B(n23555), .Z(n22) );
  AND U22950 ( .A(n70), .B(n23556), .Z(n23555) );
  XOR U22951 ( .A(p_input[11]), .B(n23554), .Z(n23556) );
  XNOR U22952 ( .A(n23557), .B(n23558), .Z(n23554) );
  AND U22953 ( .A(n74), .B(n23559), .Z(n23558) );
  XOR U22954 ( .A(n23560), .B(n23561), .Z(n23552) );
  AND U22955 ( .A(n78), .B(n23551), .Z(n23561) );
  XNOR U22956 ( .A(n23562), .B(n23549), .Z(n23551) );
  XOR U22957 ( .A(n23563), .B(n23564), .Z(n23549) );
  AND U22958 ( .A(n102), .B(n23565), .Z(n23564) );
  IV U22959 ( .A(n23560), .Z(n23562) );
  XOR U22960 ( .A(n23566), .B(n23567), .Z(n23560) );
  AND U22961 ( .A(n86), .B(n23559), .Z(n23567) );
  XNOR U22962 ( .A(n23557), .B(n23566), .Z(n23559) );
  XNOR U22963 ( .A(n23568), .B(n23569), .Z(n23557) );
  AND U22964 ( .A(n90), .B(n23570), .Z(n23569) );
  XOR U22965 ( .A(p_input[27]), .B(n23568), .Z(n23570) );
  XNOR U22966 ( .A(n23571), .B(n23572), .Z(n23568) );
  AND U22967 ( .A(n94), .B(n23573), .Z(n23572) );
  XOR U22968 ( .A(n23574), .B(n23575), .Z(n23566) );
  AND U22969 ( .A(n98), .B(n23565), .Z(n23575) );
  XNOR U22970 ( .A(n23576), .B(n23563), .Z(n23565) );
  XOR U22971 ( .A(n23577), .B(n23578), .Z(n23563) );
  AND U22972 ( .A(n121), .B(n23579), .Z(n23578) );
  IV U22973 ( .A(n23574), .Z(n23576) );
  XOR U22974 ( .A(n23580), .B(n23581), .Z(n23574) );
  AND U22975 ( .A(n105), .B(n23573), .Z(n23581) );
  XNOR U22976 ( .A(n23571), .B(n23580), .Z(n23573) );
  XNOR U22977 ( .A(n23582), .B(n23583), .Z(n23571) );
  AND U22978 ( .A(n109), .B(n23584), .Z(n23583) );
  XOR U22979 ( .A(p_input[43]), .B(n23582), .Z(n23584) );
  XNOR U22980 ( .A(n23585), .B(n23586), .Z(n23582) );
  AND U22981 ( .A(n113), .B(n23587), .Z(n23586) );
  XOR U22982 ( .A(n23588), .B(n23589), .Z(n23580) );
  AND U22983 ( .A(n117), .B(n23579), .Z(n23589) );
  XNOR U22984 ( .A(n23590), .B(n23577), .Z(n23579) );
  XOR U22985 ( .A(n23591), .B(n23592), .Z(n23577) );
  AND U22986 ( .A(n140), .B(n23593), .Z(n23592) );
  IV U22987 ( .A(n23588), .Z(n23590) );
  XOR U22988 ( .A(n23594), .B(n23595), .Z(n23588) );
  AND U22989 ( .A(n124), .B(n23587), .Z(n23595) );
  XNOR U22990 ( .A(n23585), .B(n23594), .Z(n23587) );
  XNOR U22991 ( .A(n23596), .B(n23597), .Z(n23585) );
  AND U22992 ( .A(n128), .B(n23598), .Z(n23597) );
  XOR U22993 ( .A(p_input[59]), .B(n23596), .Z(n23598) );
  XNOR U22994 ( .A(n23599), .B(n23600), .Z(n23596) );
  AND U22995 ( .A(n132), .B(n23601), .Z(n23600) );
  XOR U22996 ( .A(n23602), .B(n23603), .Z(n23594) );
  AND U22997 ( .A(n136), .B(n23593), .Z(n23603) );
  XNOR U22998 ( .A(n23604), .B(n23591), .Z(n23593) );
  XOR U22999 ( .A(n23605), .B(n23606), .Z(n23591) );
  AND U23000 ( .A(n159), .B(n23607), .Z(n23606) );
  IV U23001 ( .A(n23602), .Z(n23604) );
  XOR U23002 ( .A(n23608), .B(n23609), .Z(n23602) );
  AND U23003 ( .A(n143), .B(n23601), .Z(n23609) );
  XNOR U23004 ( .A(n23599), .B(n23608), .Z(n23601) );
  XNOR U23005 ( .A(n23610), .B(n23611), .Z(n23599) );
  AND U23006 ( .A(n147), .B(n23612), .Z(n23611) );
  XOR U23007 ( .A(p_input[75]), .B(n23610), .Z(n23612) );
  XNOR U23008 ( .A(n23613), .B(n23614), .Z(n23610) );
  AND U23009 ( .A(n151), .B(n23615), .Z(n23614) );
  XOR U23010 ( .A(n23616), .B(n23617), .Z(n23608) );
  AND U23011 ( .A(n155), .B(n23607), .Z(n23617) );
  XNOR U23012 ( .A(n23618), .B(n23605), .Z(n23607) );
  XOR U23013 ( .A(n23619), .B(n23620), .Z(n23605) );
  AND U23014 ( .A(n178), .B(n23621), .Z(n23620) );
  IV U23015 ( .A(n23616), .Z(n23618) );
  XOR U23016 ( .A(n23622), .B(n23623), .Z(n23616) );
  AND U23017 ( .A(n162), .B(n23615), .Z(n23623) );
  XNOR U23018 ( .A(n23613), .B(n23622), .Z(n23615) );
  XNOR U23019 ( .A(n23624), .B(n23625), .Z(n23613) );
  AND U23020 ( .A(n166), .B(n23626), .Z(n23625) );
  XOR U23021 ( .A(p_input[91]), .B(n23624), .Z(n23626) );
  XNOR U23022 ( .A(n23627), .B(n23628), .Z(n23624) );
  AND U23023 ( .A(n170), .B(n23629), .Z(n23628) );
  XOR U23024 ( .A(n23630), .B(n23631), .Z(n23622) );
  AND U23025 ( .A(n174), .B(n23621), .Z(n23631) );
  XNOR U23026 ( .A(n23632), .B(n23619), .Z(n23621) );
  XOR U23027 ( .A(n23633), .B(n23634), .Z(n23619) );
  AND U23028 ( .A(n197), .B(n23635), .Z(n23634) );
  IV U23029 ( .A(n23630), .Z(n23632) );
  XOR U23030 ( .A(n23636), .B(n23637), .Z(n23630) );
  AND U23031 ( .A(n181), .B(n23629), .Z(n23637) );
  XNOR U23032 ( .A(n23627), .B(n23636), .Z(n23629) );
  XNOR U23033 ( .A(n23638), .B(n23639), .Z(n23627) );
  AND U23034 ( .A(n185), .B(n23640), .Z(n23639) );
  XOR U23035 ( .A(p_input[107]), .B(n23638), .Z(n23640) );
  XNOR U23036 ( .A(n23641), .B(n23642), .Z(n23638) );
  AND U23037 ( .A(n189), .B(n23643), .Z(n23642) );
  XOR U23038 ( .A(n23644), .B(n23645), .Z(n23636) );
  AND U23039 ( .A(n193), .B(n23635), .Z(n23645) );
  XNOR U23040 ( .A(n23646), .B(n23633), .Z(n23635) );
  XOR U23041 ( .A(n23647), .B(n23648), .Z(n23633) );
  AND U23042 ( .A(n216), .B(n23649), .Z(n23648) );
  IV U23043 ( .A(n23644), .Z(n23646) );
  XOR U23044 ( .A(n23650), .B(n23651), .Z(n23644) );
  AND U23045 ( .A(n200), .B(n23643), .Z(n23651) );
  XNOR U23046 ( .A(n23641), .B(n23650), .Z(n23643) );
  XNOR U23047 ( .A(n23652), .B(n23653), .Z(n23641) );
  AND U23048 ( .A(n204), .B(n23654), .Z(n23653) );
  XOR U23049 ( .A(p_input[123]), .B(n23652), .Z(n23654) );
  XNOR U23050 ( .A(n23655), .B(n23656), .Z(n23652) );
  AND U23051 ( .A(n208), .B(n23657), .Z(n23656) );
  XOR U23052 ( .A(n23658), .B(n23659), .Z(n23650) );
  AND U23053 ( .A(n212), .B(n23649), .Z(n23659) );
  XNOR U23054 ( .A(n23660), .B(n23647), .Z(n23649) );
  XOR U23055 ( .A(n23661), .B(n23662), .Z(n23647) );
  AND U23056 ( .A(n235), .B(n23663), .Z(n23662) );
  IV U23057 ( .A(n23658), .Z(n23660) );
  XOR U23058 ( .A(n23664), .B(n23665), .Z(n23658) );
  AND U23059 ( .A(n219), .B(n23657), .Z(n23665) );
  XNOR U23060 ( .A(n23655), .B(n23664), .Z(n23657) );
  XNOR U23061 ( .A(n23666), .B(n23667), .Z(n23655) );
  AND U23062 ( .A(n223), .B(n23668), .Z(n23667) );
  XOR U23063 ( .A(p_input[139]), .B(n23666), .Z(n23668) );
  XNOR U23064 ( .A(n23669), .B(n23670), .Z(n23666) );
  AND U23065 ( .A(n227), .B(n23671), .Z(n23670) );
  XOR U23066 ( .A(n23672), .B(n23673), .Z(n23664) );
  AND U23067 ( .A(n231), .B(n23663), .Z(n23673) );
  XNOR U23068 ( .A(n23674), .B(n23661), .Z(n23663) );
  XOR U23069 ( .A(n23675), .B(n23676), .Z(n23661) );
  AND U23070 ( .A(n254), .B(n23677), .Z(n23676) );
  IV U23071 ( .A(n23672), .Z(n23674) );
  XOR U23072 ( .A(n23678), .B(n23679), .Z(n23672) );
  AND U23073 ( .A(n238), .B(n23671), .Z(n23679) );
  XNOR U23074 ( .A(n23669), .B(n23678), .Z(n23671) );
  XNOR U23075 ( .A(n23680), .B(n23681), .Z(n23669) );
  AND U23076 ( .A(n242), .B(n23682), .Z(n23681) );
  XOR U23077 ( .A(p_input[155]), .B(n23680), .Z(n23682) );
  XNOR U23078 ( .A(n23683), .B(n23684), .Z(n23680) );
  AND U23079 ( .A(n246), .B(n23685), .Z(n23684) );
  XOR U23080 ( .A(n23686), .B(n23687), .Z(n23678) );
  AND U23081 ( .A(n250), .B(n23677), .Z(n23687) );
  XNOR U23082 ( .A(n23688), .B(n23675), .Z(n23677) );
  XOR U23083 ( .A(n23689), .B(n23690), .Z(n23675) );
  AND U23084 ( .A(n273), .B(n23691), .Z(n23690) );
  IV U23085 ( .A(n23686), .Z(n23688) );
  XOR U23086 ( .A(n23692), .B(n23693), .Z(n23686) );
  AND U23087 ( .A(n257), .B(n23685), .Z(n23693) );
  XNOR U23088 ( .A(n23683), .B(n23692), .Z(n23685) );
  XNOR U23089 ( .A(n23694), .B(n23695), .Z(n23683) );
  AND U23090 ( .A(n261), .B(n23696), .Z(n23695) );
  XOR U23091 ( .A(p_input[171]), .B(n23694), .Z(n23696) );
  XNOR U23092 ( .A(n23697), .B(n23698), .Z(n23694) );
  AND U23093 ( .A(n265), .B(n23699), .Z(n23698) );
  XOR U23094 ( .A(n23700), .B(n23701), .Z(n23692) );
  AND U23095 ( .A(n269), .B(n23691), .Z(n23701) );
  XNOR U23096 ( .A(n23702), .B(n23689), .Z(n23691) );
  XOR U23097 ( .A(n23703), .B(n23704), .Z(n23689) );
  AND U23098 ( .A(n292), .B(n23705), .Z(n23704) );
  IV U23099 ( .A(n23700), .Z(n23702) );
  XOR U23100 ( .A(n23706), .B(n23707), .Z(n23700) );
  AND U23101 ( .A(n276), .B(n23699), .Z(n23707) );
  XNOR U23102 ( .A(n23697), .B(n23706), .Z(n23699) );
  XNOR U23103 ( .A(n23708), .B(n23709), .Z(n23697) );
  AND U23104 ( .A(n280), .B(n23710), .Z(n23709) );
  XOR U23105 ( .A(p_input[187]), .B(n23708), .Z(n23710) );
  XNOR U23106 ( .A(n23711), .B(n23712), .Z(n23708) );
  AND U23107 ( .A(n284), .B(n23713), .Z(n23712) );
  XOR U23108 ( .A(n23714), .B(n23715), .Z(n23706) );
  AND U23109 ( .A(n288), .B(n23705), .Z(n23715) );
  XNOR U23110 ( .A(n23716), .B(n23703), .Z(n23705) );
  XOR U23111 ( .A(n23717), .B(n23718), .Z(n23703) );
  AND U23112 ( .A(n311), .B(n23719), .Z(n23718) );
  IV U23113 ( .A(n23714), .Z(n23716) );
  XOR U23114 ( .A(n23720), .B(n23721), .Z(n23714) );
  AND U23115 ( .A(n295), .B(n23713), .Z(n23721) );
  XNOR U23116 ( .A(n23711), .B(n23720), .Z(n23713) );
  XNOR U23117 ( .A(n23722), .B(n23723), .Z(n23711) );
  AND U23118 ( .A(n299), .B(n23724), .Z(n23723) );
  XOR U23119 ( .A(p_input[203]), .B(n23722), .Z(n23724) );
  XNOR U23120 ( .A(n23725), .B(n23726), .Z(n23722) );
  AND U23121 ( .A(n303), .B(n23727), .Z(n23726) );
  XOR U23122 ( .A(n23728), .B(n23729), .Z(n23720) );
  AND U23123 ( .A(n307), .B(n23719), .Z(n23729) );
  XNOR U23124 ( .A(n23730), .B(n23717), .Z(n23719) );
  XOR U23125 ( .A(n23731), .B(n23732), .Z(n23717) );
  AND U23126 ( .A(n330), .B(n23733), .Z(n23732) );
  IV U23127 ( .A(n23728), .Z(n23730) );
  XOR U23128 ( .A(n23734), .B(n23735), .Z(n23728) );
  AND U23129 ( .A(n314), .B(n23727), .Z(n23735) );
  XNOR U23130 ( .A(n23725), .B(n23734), .Z(n23727) );
  XNOR U23131 ( .A(n23736), .B(n23737), .Z(n23725) );
  AND U23132 ( .A(n318), .B(n23738), .Z(n23737) );
  XOR U23133 ( .A(p_input[219]), .B(n23736), .Z(n23738) );
  XNOR U23134 ( .A(n23739), .B(n23740), .Z(n23736) );
  AND U23135 ( .A(n322), .B(n23741), .Z(n23740) );
  XOR U23136 ( .A(n23742), .B(n23743), .Z(n23734) );
  AND U23137 ( .A(n326), .B(n23733), .Z(n23743) );
  XNOR U23138 ( .A(n23744), .B(n23731), .Z(n23733) );
  XOR U23139 ( .A(n23745), .B(n23746), .Z(n23731) );
  AND U23140 ( .A(n349), .B(n23747), .Z(n23746) );
  IV U23141 ( .A(n23742), .Z(n23744) );
  XOR U23142 ( .A(n23748), .B(n23749), .Z(n23742) );
  AND U23143 ( .A(n333), .B(n23741), .Z(n23749) );
  XNOR U23144 ( .A(n23739), .B(n23748), .Z(n23741) );
  XNOR U23145 ( .A(n23750), .B(n23751), .Z(n23739) );
  AND U23146 ( .A(n337), .B(n23752), .Z(n23751) );
  XOR U23147 ( .A(p_input[235]), .B(n23750), .Z(n23752) );
  XNOR U23148 ( .A(n23753), .B(n23754), .Z(n23750) );
  AND U23149 ( .A(n341), .B(n23755), .Z(n23754) );
  XOR U23150 ( .A(n23756), .B(n23757), .Z(n23748) );
  AND U23151 ( .A(n345), .B(n23747), .Z(n23757) );
  XNOR U23152 ( .A(n23758), .B(n23745), .Z(n23747) );
  XOR U23153 ( .A(n23759), .B(n23760), .Z(n23745) );
  AND U23154 ( .A(n368), .B(n23761), .Z(n23760) );
  IV U23155 ( .A(n23756), .Z(n23758) );
  XOR U23156 ( .A(n23762), .B(n23763), .Z(n23756) );
  AND U23157 ( .A(n352), .B(n23755), .Z(n23763) );
  XNOR U23158 ( .A(n23753), .B(n23762), .Z(n23755) );
  XNOR U23159 ( .A(n23764), .B(n23765), .Z(n23753) );
  AND U23160 ( .A(n356), .B(n23766), .Z(n23765) );
  XOR U23161 ( .A(p_input[251]), .B(n23764), .Z(n23766) );
  XNOR U23162 ( .A(n23767), .B(n23768), .Z(n23764) );
  AND U23163 ( .A(n360), .B(n23769), .Z(n23768) );
  XOR U23164 ( .A(n23770), .B(n23771), .Z(n23762) );
  AND U23165 ( .A(n364), .B(n23761), .Z(n23771) );
  XNOR U23166 ( .A(n23772), .B(n23759), .Z(n23761) );
  XOR U23167 ( .A(n23773), .B(n23774), .Z(n23759) );
  AND U23168 ( .A(n387), .B(n23775), .Z(n23774) );
  IV U23169 ( .A(n23770), .Z(n23772) );
  XOR U23170 ( .A(n23776), .B(n23777), .Z(n23770) );
  AND U23171 ( .A(n371), .B(n23769), .Z(n23777) );
  XNOR U23172 ( .A(n23767), .B(n23776), .Z(n23769) );
  XNOR U23173 ( .A(n23778), .B(n23779), .Z(n23767) );
  AND U23174 ( .A(n375), .B(n23780), .Z(n23779) );
  XOR U23175 ( .A(p_input[267]), .B(n23778), .Z(n23780) );
  XNOR U23176 ( .A(n23781), .B(n23782), .Z(n23778) );
  AND U23177 ( .A(n379), .B(n23783), .Z(n23782) );
  XOR U23178 ( .A(n23784), .B(n23785), .Z(n23776) );
  AND U23179 ( .A(n383), .B(n23775), .Z(n23785) );
  XNOR U23180 ( .A(n23786), .B(n23773), .Z(n23775) );
  XOR U23181 ( .A(n23787), .B(n23788), .Z(n23773) );
  AND U23182 ( .A(n406), .B(n23789), .Z(n23788) );
  IV U23183 ( .A(n23784), .Z(n23786) );
  XOR U23184 ( .A(n23790), .B(n23791), .Z(n23784) );
  AND U23185 ( .A(n390), .B(n23783), .Z(n23791) );
  XNOR U23186 ( .A(n23781), .B(n23790), .Z(n23783) );
  XNOR U23187 ( .A(n23792), .B(n23793), .Z(n23781) );
  AND U23188 ( .A(n394), .B(n23794), .Z(n23793) );
  XOR U23189 ( .A(p_input[283]), .B(n23792), .Z(n23794) );
  XNOR U23190 ( .A(n23795), .B(n23796), .Z(n23792) );
  AND U23191 ( .A(n398), .B(n23797), .Z(n23796) );
  XOR U23192 ( .A(n23798), .B(n23799), .Z(n23790) );
  AND U23193 ( .A(n402), .B(n23789), .Z(n23799) );
  XNOR U23194 ( .A(n23800), .B(n23787), .Z(n23789) );
  XOR U23195 ( .A(n23801), .B(n23802), .Z(n23787) );
  AND U23196 ( .A(n425), .B(n23803), .Z(n23802) );
  IV U23197 ( .A(n23798), .Z(n23800) );
  XOR U23198 ( .A(n23804), .B(n23805), .Z(n23798) );
  AND U23199 ( .A(n409), .B(n23797), .Z(n23805) );
  XNOR U23200 ( .A(n23795), .B(n23804), .Z(n23797) );
  XNOR U23201 ( .A(n23806), .B(n23807), .Z(n23795) );
  AND U23202 ( .A(n413), .B(n23808), .Z(n23807) );
  XOR U23203 ( .A(p_input[299]), .B(n23806), .Z(n23808) );
  XNOR U23204 ( .A(n23809), .B(n23810), .Z(n23806) );
  AND U23205 ( .A(n417), .B(n23811), .Z(n23810) );
  XOR U23206 ( .A(n23812), .B(n23813), .Z(n23804) );
  AND U23207 ( .A(n421), .B(n23803), .Z(n23813) );
  XNOR U23208 ( .A(n23814), .B(n23801), .Z(n23803) );
  XOR U23209 ( .A(n23815), .B(n23816), .Z(n23801) );
  AND U23210 ( .A(n444), .B(n23817), .Z(n23816) );
  IV U23211 ( .A(n23812), .Z(n23814) );
  XOR U23212 ( .A(n23818), .B(n23819), .Z(n23812) );
  AND U23213 ( .A(n428), .B(n23811), .Z(n23819) );
  XNOR U23214 ( .A(n23809), .B(n23818), .Z(n23811) );
  XNOR U23215 ( .A(n23820), .B(n23821), .Z(n23809) );
  AND U23216 ( .A(n432), .B(n23822), .Z(n23821) );
  XOR U23217 ( .A(p_input[315]), .B(n23820), .Z(n23822) );
  XNOR U23218 ( .A(n23823), .B(n23824), .Z(n23820) );
  AND U23219 ( .A(n436), .B(n23825), .Z(n23824) );
  XOR U23220 ( .A(n23826), .B(n23827), .Z(n23818) );
  AND U23221 ( .A(n440), .B(n23817), .Z(n23827) );
  XNOR U23222 ( .A(n23828), .B(n23815), .Z(n23817) );
  XOR U23223 ( .A(n23829), .B(n23830), .Z(n23815) );
  AND U23224 ( .A(n463), .B(n23831), .Z(n23830) );
  IV U23225 ( .A(n23826), .Z(n23828) );
  XOR U23226 ( .A(n23832), .B(n23833), .Z(n23826) );
  AND U23227 ( .A(n447), .B(n23825), .Z(n23833) );
  XNOR U23228 ( .A(n23823), .B(n23832), .Z(n23825) );
  XNOR U23229 ( .A(n23834), .B(n23835), .Z(n23823) );
  AND U23230 ( .A(n451), .B(n23836), .Z(n23835) );
  XOR U23231 ( .A(p_input[331]), .B(n23834), .Z(n23836) );
  XNOR U23232 ( .A(n23837), .B(n23838), .Z(n23834) );
  AND U23233 ( .A(n455), .B(n23839), .Z(n23838) );
  XOR U23234 ( .A(n23840), .B(n23841), .Z(n23832) );
  AND U23235 ( .A(n459), .B(n23831), .Z(n23841) );
  XNOR U23236 ( .A(n23842), .B(n23829), .Z(n23831) );
  XOR U23237 ( .A(n23843), .B(n23844), .Z(n23829) );
  AND U23238 ( .A(n482), .B(n23845), .Z(n23844) );
  IV U23239 ( .A(n23840), .Z(n23842) );
  XOR U23240 ( .A(n23846), .B(n23847), .Z(n23840) );
  AND U23241 ( .A(n466), .B(n23839), .Z(n23847) );
  XNOR U23242 ( .A(n23837), .B(n23846), .Z(n23839) );
  XNOR U23243 ( .A(n23848), .B(n23849), .Z(n23837) );
  AND U23244 ( .A(n470), .B(n23850), .Z(n23849) );
  XOR U23245 ( .A(p_input[347]), .B(n23848), .Z(n23850) );
  XNOR U23246 ( .A(n23851), .B(n23852), .Z(n23848) );
  AND U23247 ( .A(n474), .B(n23853), .Z(n23852) );
  XOR U23248 ( .A(n23854), .B(n23855), .Z(n23846) );
  AND U23249 ( .A(n478), .B(n23845), .Z(n23855) );
  XNOR U23250 ( .A(n23856), .B(n23843), .Z(n23845) );
  XOR U23251 ( .A(n23857), .B(n23858), .Z(n23843) );
  AND U23252 ( .A(n501), .B(n23859), .Z(n23858) );
  IV U23253 ( .A(n23854), .Z(n23856) );
  XOR U23254 ( .A(n23860), .B(n23861), .Z(n23854) );
  AND U23255 ( .A(n485), .B(n23853), .Z(n23861) );
  XNOR U23256 ( .A(n23851), .B(n23860), .Z(n23853) );
  XNOR U23257 ( .A(n23862), .B(n23863), .Z(n23851) );
  AND U23258 ( .A(n489), .B(n23864), .Z(n23863) );
  XOR U23259 ( .A(p_input[363]), .B(n23862), .Z(n23864) );
  XNOR U23260 ( .A(n23865), .B(n23866), .Z(n23862) );
  AND U23261 ( .A(n493), .B(n23867), .Z(n23866) );
  XOR U23262 ( .A(n23868), .B(n23869), .Z(n23860) );
  AND U23263 ( .A(n497), .B(n23859), .Z(n23869) );
  XNOR U23264 ( .A(n23870), .B(n23857), .Z(n23859) );
  XOR U23265 ( .A(n23871), .B(n23872), .Z(n23857) );
  AND U23266 ( .A(n520), .B(n23873), .Z(n23872) );
  IV U23267 ( .A(n23868), .Z(n23870) );
  XOR U23268 ( .A(n23874), .B(n23875), .Z(n23868) );
  AND U23269 ( .A(n504), .B(n23867), .Z(n23875) );
  XNOR U23270 ( .A(n23865), .B(n23874), .Z(n23867) );
  XNOR U23271 ( .A(n23876), .B(n23877), .Z(n23865) );
  AND U23272 ( .A(n508), .B(n23878), .Z(n23877) );
  XOR U23273 ( .A(p_input[379]), .B(n23876), .Z(n23878) );
  XNOR U23274 ( .A(n23879), .B(n23880), .Z(n23876) );
  AND U23275 ( .A(n512), .B(n23881), .Z(n23880) );
  XOR U23276 ( .A(n23882), .B(n23883), .Z(n23874) );
  AND U23277 ( .A(n516), .B(n23873), .Z(n23883) );
  XNOR U23278 ( .A(n23884), .B(n23871), .Z(n23873) );
  XOR U23279 ( .A(n23885), .B(n23886), .Z(n23871) );
  AND U23280 ( .A(n539), .B(n23887), .Z(n23886) );
  IV U23281 ( .A(n23882), .Z(n23884) );
  XOR U23282 ( .A(n23888), .B(n23889), .Z(n23882) );
  AND U23283 ( .A(n523), .B(n23881), .Z(n23889) );
  XNOR U23284 ( .A(n23879), .B(n23888), .Z(n23881) );
  XNOR U23285 ( .A(n23890), .B(n23891), .Z(n23879) );
  AND U23286 ( .A(n527), .B(n23892), .Z(n23891) );
  XOR U23287 ( .A(p_input[395]), .B(n23890), .Z(n23892) );
  XNOR U23288 ( .A(n23893), .B(n23894), .Z(n23890) );
  AND U23289 ( .A(n531), .B(n23895), .Z(n23894) );
  XOR U23290 ( .A(n23896), .B(n23897), .Z(n23888) );
  AND U23291 ( .A(n535), .B(n23887), .Z(n23897) );
  XNOR U23292 ( .A(n23898), .B(n23885), .Z(n23887) );
  XOR U23293 ( .A(n23899), .B(n23900), .Z(n23885) );
  AND U23294 ( .A(n558), .B(n23901), .Z(n23900) );
  IV U23295 ( .A(n23896), .Z(n23898) );
  XOR U23296 ( .A(n23902), .B(n23903), .Z(n23896) );
  AND U23297 ( .A(n542), .B(n23895), .Z(n23903) );
  XNOR U23298 ( .A(n23893), .B(n23902), .Z(n23895) );
  XNOR U23299 ( .A(n23904), .B(n23905), .Z(n23893) );
  AND U23300 ( .A(n546), .B(n23906), .Z(n23905) );
  XOR U23301 ( .A(p_input[411]), .B(n23904), .Z(n23906) );
  XNOR U23302 ( .A(n23907), .B(n23908), .Z(n23904) );
  AND U23303 ( .A(n550), .B(n23909), .Z(n23908) );
  XOR U23304 ( .A(n23910), .B(n23911), .Z(n23902) );
  AND U23305 ( .A(n554), .B(n23901), .Z(n23911) );
  XNOR U23306 ( .A(n23912), .B(n23899), .Z(n23901) );
  XOR U23307 ( .A(n23913), .B(n23914), .Z(n23899) );
  AND U23308 ( .A(n577), .B(n23915), .Z(n23914) );
  IV U23309 ( .A(n23910), .Z(n23912) );
  XOR U23310 ( .A(n23916), .B(n23917), .Z(n23910) );
  AND U23311 ( .A(n561), .B(n23909), .Z(n23917) );
  XNOR U23312 ( .A(n23907), .B(n23916), .Z(n23909) );
  XNOR U23313 ( .A(n23918), .B(n23919), .Z(n23907) );
  AND U23314 ( .A(n565), .B(n23920), .Z(n23919) );
  XOR U23315 ( .A(p_input[427]), .B(n23918), .Z(n23920) );
  XNOR U23316 ( .A(n23921), .B(n23922), .Z(n23918) );
  AND U23317 ( .A(n569), .B(n23923), .Z(n23922) );
  XOR U23318 ( .A(n23924), .B(n23925), .Z(n23916) );
  AND U23319 ( .A(n573), .B(n23915), .Z(n23925) );
  XNOR U23320 ( .A(n23926), .B(n23913), .Z(n23915) );
  XOR U23321 ( .A(n23927), .B(n23928), .Z(n23913) );
  AND U23322 ( .A(n596), .B(n23929), .Z(n23928) );
  IV U23323 ( .A(n23924), .Z(n23926) );
  XOR U23324 ( .A(n23930), .B(n23931), .Z(n23924) );
  AND U23325 ( .A(n580), .B(n23923), .Z(n23931) );
  XNOR U23326 ( .A(n23921), .B(n23930), .Z(n23923) );
  XNOR U23327 ( .A(n23932), .B(n23933), .Z(n23921) );
  AND U23328 ( .A(n584), .B(n23934), .Z(n23933) );
  XOR U23329 ( .A(p_input[443]), .B(n23932), .Z(n23934) );
  XNOR U23330 ( .A(n23935), .B(n23936), .Z(n23932) );
  AND U23331 ( .A(n588), .B(n23937), .Z(n23936) );
  XOR U23332 ( .A(n23938), .B(n23939), .Z(n23930) );
  AND U23333 ( .A(n592), .B(n23929), .Z(n23939) );
  XNOR U23334 ( .A(n23940), .B(n23927), .Z(n23929) );
  XOR U23335 ( .A(n23941), .B(n23942), .Z(n23927) );
  AND U23336 ( .A(n615), .B(n23943), .Z(n23942) );
  IV U23337 ( .A(n23938), .Z(n23940) );
  XOR U23338 ( .A(n23944), .B(n23945), .Z(n23938) );
  AND U23339 ( .A(n599), .B(n23937), .Z(n23945) );
  XNOR U23340 ( .A(n23935), .B(n23944), .Z(n23937) );
  XNOR U23341 ( .A(n23946), .B(n23947), .Z(n23935) );
  AND U23342 ( .A(n603), .B(n23948), .Z(n23947) );
  XOR U23343 ( .A(p_input[459]), .B(n23946), .Z(n23948) );
  XNOR U23344 ( .A(n23949), .B(n23950), .Z(n23946) );
  AND U23345 ( .A(n607), .B(n23951), .Z(n23950) );
  XOR U23346 ( .A(n23952), .B(n23953), .Z(n23944) );
  AND U23347 ( .A(n611), .B(n23943), .Z(n23953) );
  XNOR U23348 ( .A(n23954), .B(n23941), .Z(n23943) );
  XOR U23349 ( .A(n23955), .B(n23956), .Z(n23941) );
  AND U23350 ( .A(n634), .B(n23957), .Z(n23956) );
  IV U23351 ( .A(n23952), .Z(n23954) );
  XOR U23352 ( .A(n23958), .B(n23959), .Z(n23952) );
  AND U23353 ( .A(n618), .B(n23951), .Z(n23959) );
  XNOR U23354 ( .A(n23949), .B(n23958), .Z(n23951) );
  XNOR U23355 ( .A(n23960), .B(n23961), .Z(n23949) );
  AND U23356 ( .A(n622), .B(n23962), .Z(n23961) );
  XOR U23357 ( .A(p_input[475]), .B(n23960), .Z(n23962) );
  XNOR U23358 ( .A(n23963), .B(n23964), .Z(n23960) );
  AND U23359 ( .A(n626), .B(n23965), .Z(n23964) );
  XOR U23360 ( .A(n23966), .B(n23967), .Z(n23958) );
  AND U23361 ( .A(n630), .B(n23957), .Z(n23967) );
  XNOR U23362 ( .A(n23968), .B(n23955), .Z(n23957) );
  XOR U23363 ( .A(n23969), .B(n23970), .Z(n23955) );
  AND U23364 ( .A(n653), .B(n23971), .Z(n23970) );
  IV U23365 ( .A(n23966), .Z(n23968) );
  XOR U23366 ( .A(n23972), .B(n23973), .Z(n23966) );
  AND U23367 ( .A(n637), .B(n23965), .Z(n23973) );
  XNOR U23368 ( .A(n23963), .B(n23972), .Z(n23965) );
  XNOR U23369 ( .A(n23974), .B(n23975), .Z(n23963) );
  AND U23370 ( .A(n641), .B(n23976), .Z(n23975) );
  XOR U23371 ( .A(p_input[491]), .B(n23974), .Z(n23976) );
  XNOR U23372 ( .A(n23977), .B(n23978), .Z(n23974) );
  AND U23373 ( .A(n645), .B(n23979), .Z(n23978) );
  XOR U23374 ( .A(n23980), .B(n23981), .Z(n23972) );
  AND U23375 ( .A(n649), .B(n23971), .Z(n23981) );
  XNOR U23376 ( .A(n23982), .B(n23969), .Z(n23971) );
  XOR U23377 ( .A(n23983), .B(n23984), .Z(n23969) );
  AND U23378 ( .A(n672), .B(n23985), .Z(n23984) );
  IV U23379 ( .A(n23980), .Z(n23982) );
  XOR U23380 ( .A(n23986), .B(n23987), .Z(n23980) );
  AND U23381 ( .A(n656), .B(n23979), .Z(n23987) );
  XNOR U23382 ( .A(n23977), .B(n23986), .Z(n23979) );
  XNOR U23383 ( .A(n23988), .B(n23989), .Z(n23977) );
  AND U23384 ( .A(n660), .B(n23990), .Z(n23989) );
  XOR U23385 ( .A(p_input[507]), .B(n23988), .Z(n23990) );
  XNOR U23386 ( .A(n23991), .B(n23992), .Z(n23988) );
  AND U23387 ( .A(n664), .B(n23993), .Z(n23992) );
  XOR U23388 ( .A(n23994), .B(n23995), .Z(n23986) );
  AND U23389 ( .A(n668), .B(n23985), .Z(n23995) );
  XNOR U23390 ( .A(n23996), .B(n23983), .Z(n23985) );
  XOR U23391 ( .A(n23997), .B(n23998), .Z(n23983) );
  AND U23392 ( .A(n691), .B(n23999), .Z(n23998) );
  IV U23393 ( .A(n23994), .Z(n23996) );
  XOR U23394 ( .A(n24000), .B(n24001), .Z(n23994) );
  AND U23395 ( .A(n675), .B(n23993), .Z(n24001) );
  XNOR U23396 ( .A(n23991), .B(n24000), .Z(n23993) );
  XNOR U23397 ( .A(n24002), .B(n24003), .Z(n23991) );
  AND U23398 ( .A(n679), .B(n24004), .Z(n24003) );
  XOR U23399 ( .A(p_input[523]), .B(n24002), .Z(n24004) );
  XNOR U23400 ( .A(n24005), .B(n24006), .Z(n24002) );
  AND U23401 ( .A(n683), .B(n24007), .Z(n24006) );
  XOR U23402 ( .A(n24008), .B(n24009), .Z(n24000) );
  AND U23403 ( .A(n687), .B(n23999), .Z(n24009) );
  XNOR U23404 ( .A(n24010), .B(n23997), .Z(n23999) );
  XOR U23405 ( .A(n24011), .B(n24012), .Z(n23997) );
  AND U23406 ( .A(n710), .B(n24013), .Z(n24012) );
  IV U23407 ( .A(n24008), .Z(n24010) );
  XOR U23408 ( .A(n24014), .B(n24015), .Z(n24008) );
  AND U23409 ( .A(n694), .B(n24007), .Z(n24015) );
  XNOR U23410 ( .A(n24005), .B(n24014), .Z(n24007) );
  XNOR U23411 ( .A(n24016), .B(n24017), .Z(n24005) );
  AND U23412 ( .A(n698), .B(n24018), .Z(n24017) );
  XOR U23413 ( .A(p_input[539]), .B(n24016), .Z(n24018) );
  XNOR U23414 ( .A(n24019), .B(n24020), .Z(n24016) );
  AND U23415 ( .A(n702), .B(n24021), .Z(n24020) );
  XOR U23416 ( .A(n24022), .B(n24023), .Z(n24014) );
  AND U23417 ( .A(n706), .B(n24013), .Z(n24023) );
  XNOR U23418 ( .A(n24024), .B(n24011), .Z(n24013) );
  XOR U23419 ( .A(n24025), .B(n24026), .Z(n24011) );
  AND U23420 ( .A(n729), .B(n24027), .Z(n24026) );
  IV U23421 ( .A(n24022), .Z(n24024) );
  XOR U23422 ( .A(n24028), .B(n24029), .Z(n24022) );
  AND U23423 ( .A(n713), .B(n24021), .Z(n24029) );
  XNOR U23424 ( .A(n24019), .B(n24028), .Z(n24021) );
  XNOR U23425 ( .A(n24030), .B(n24031), .Z(n24019) );
  AND U23426 ( .A(n717), .B(n24032), .Z(n24031) );
  XOR U23427 ( .A(p_input[555]), .B(n24030), .Z(n24032) );
  XNOR U23428 ( .A(n24033), .B(n24034), .Z(n24030) );
  AND U23429 ( .A(n721), .B(n24035), .Z(n24034) );
  XOR U23430 ( .A(n24036), .B(n24037), .Z(n24028) );
  AND U23431 ( .A(n725), .B(n24027), .Z(n24037) );
  XNOR U23432 ( .A(n24038), .B(n24025), .Z(n24027) );
  XOR U23433 ( .A(n24039), .B(n24040), .Z(n24025) );
  AND U23434 ( .A(n748), .B(n24041), .Z(n24040) );
  IV U23435 ( .A(n24036), .Z(n24038) );
  XOR U23436 ( .A(n24042), .B(n24043), .Z(n24036) );
  AND U23437 ( .A(n732), .B(n24035), .Z(n24043) );
  XNOR U23438 ( .A(n24033), .B(n24042), .Z(n24035) );
  XNOR U23439 ( .A(n24044), .B(n24045), .Z(n24033) );
  AND U23440 ( .A(n736), .B(n24046), .Z(n24045) );
  XOR U23441 ( .A(p_input[571]), .B(n24044), .Z(n24046) );
  XNOR U23442 ( .A(n24047), .B(n24048), .Z(n24044) );
  AND U23443 ( .A(n740), .B(n24049), .Z(n24048) );
  XOR U23444 ( .A(n24050), .B(n24051), .Z(n24042) );
  AND U23445 ( .A(n744), .B(n24041), .Z(n24051) );
  XNOR U23446 ( .A(n24052), .B(n24039), .Z(n24041) );
  XOR U23447 ( .A(n24053), .B(n24054), .Z(n24039) );
  AND U23448 ( .A(n767), .B(n24055), .Z(n24054) );
  IV U23449 ( .A(n24050), .Z(n24052) );
  XOR U23450 ( .A(n24056), .B(n24057), .Z(n24050) );
  AND U23451 ( .A(n751), .B(n24049), .Z(n24057) );
  XNOR U23452 ( .A(n24047), .B(n24056), .Z(n24049) );
  XNOR U23453 ( .A(n24058), .B(n24059), .Z(n24047) );
  AND U23454 ( .A(n755), .B(n24060), .Z(n24059) );
  XOR U23455 ( .A(p_input[587]), .B(n24058), .Z(n24060) );
  XNOR U23456 ( .A(n24061), .B(n24062), .Z(n24058) );
  AND U23457 ( .A(n759), .B(n24063), .Z(n24062) );
  XOR U23458 ( .A(n24064), .B(n24065), .Z(n24056) );
  AND U23459 ( .A(n763), .B(n24055), .Z(n24065) );
  XNOR U23460 ( .A(n24066), .B(n24053), .Z(n24055) );
  XOR U23461 ( .A(n24067), .B(n24068), .Z(n24053) );
  AND U23462 ( .A(n786), .B(n24069), .Z(n24068) );
  IV U23463 ( .A(n24064), .Z(n24066) );
  XOR U23464 ( .A(n24070), .B(n24071), .Z(n24064) );
  AND U23465 ( .A(n770), .B(n24063), .Z(n24071) );
  XNOR U23466 ( .A(n24061), .B(n24070), .Z(n24063) );
  XNOR U23467 ( .A(n24072), .B(n24073), .Z(n24061) );
  AND U23468 ( .A(n774), .B(n24074), .Z(n24073) );
  XOR U23469 ( .A(p_input[603]), .B(n24072), .Z(n24074) );
  XNOR U23470 ( .A(n24075), .B(n24076), .Z(n24072) );
  AND U23471 ( .A(n778), .B(n24077), .Z(n24076) );
  XOR U23472 ( .A(n24078), .B(n24079), .Z(n24070) );
  AND U23473 ( .A(n782), .B(n24069), .Z(n24079) );
  XNOR U23474 ( .A(n24080), .B(n24067), .Z(n24069) );
  XOR U23475 ( .A(n24081), .B(n24082), .Z(n24067) );
  AND U23476 ( .A(n805), .B(n24083), .Z(n24082) );
  IV U23477 ( .A(n24078), .Z(n24080) );
  XOR U23478 ( .A(n24084), .B(n24085), .Z(n24078) );
  AND U23479 ( .A(n789), .B(n24077), .Z(n24085) );
  XNOR U23480 ( .A(n24075), .B(n24084), .Z(n24077) );
  XNOR U23481 ( .A(n24086), .B(n24087), .Z(n24075) );
  AND U23482 ( .A(n793), .B(n24088), .Z(n24087) );
  XOR U23483 ( .A(p_input[619]), .B(n24086), .Z(n24088) );
  XNOR U23484 ( .A(n24089), .B(n24090), .Z(n24086) );
  AND U23485 ( .A(n797), .B(n24091), .Z(n24090) );
  XOR U23486 ( .A(n24092), .B(n24093), .Z(n24084) );
  AND U23487 ( .A(n801), .B(n24083), .Z(n24093) );
  XNOR U23488 ( .A(n24094), .B(n24081), .Z(n24083) );
  XOR U23489 ( .A(n24095), .B(n24096), .Z(n24081) );
  AND U23490 ( .A(n824), .B(n24097), .Z(n24096) );
  IV U23491 ( .A(n24092), .Z(n24094) );
  XOR U23492 ( .A(n24098), .B(n24099), .Z(n24092) );
  AND U23493 ( .A(n808), .B(n24091), .Z(n24099) );
  XNOR U23494 ( .A(n24089), .B(n24098), .Z(n24091) );
  XNOR U23495 ( .A(n24100), .B(n24101), .Z(n24089) );
  AND U23496 ( .A(n812), .B(n24102), .Z(n24101) );
  XOR U23497 ( .A(p_input[635]), .B(n24100), .Z(n24102) );
  XNOR U23498 ( .A(n24103), .B(n24104), .Z(n24100) );
  AND U23499 ( .A(n816), .B(n24105), .Z(n24104) );
  XOR U23500 ( .A(n24106), .B(n24107), .Z(n24098) );
  AND U23501 ( .A(n820), .B(n24097), .Z(n24107) );
  XNOR U23502 ( .A(n24108), .B(n24095), .Z(n24097) );
  XOR U23503 ( .A(n24109), .B(n24110), .Z(n24095) );
  AND U23504 ( .A(n843), .B(n24111), .Z(n24110) );
  IV U23505 ( .A(n24106), .Z(n24108) );
  XOR U23506 ( .A(n24112), .B(n24113), .Z(n24106) );
  AND U23507 ( .A(n827), .B(n24105), .Z(n24113) );
  XNOR U23508 ( .A(n24103), .B(n24112), .Z(n24105) );
  XNOR U23509 ( .A(n24114), .B(n24115), .Z(n24103) );
  AND U23510 ( .A(n831), .B(n24116), .Z(n24115) );
  XOR U23511 ( .A(p_input[651]), .B(n24114), .Z(n24116) );
  XNOR U23512 ( .A(n24117), .B(n24118), .Z(n24114) );
  AND U23513 ( .A(n835), .B(n24119), .Z(n24118) );
  XOR U23514 ( .A(n24120), .B(n24121), .Z(n24112) );
  AND U23515 ( .A(n839), .B(n24111), .Z(n24121) );
  XNOR U23516 ( .A(n24122), .B(n24109), .Z(n24111) );
  XOR U23517 ( .A(n24123), .B(n24124), .Z(n24109) );
  AND U23518 ( .A(n862), .B(n24125), .Z(n24124) );
  IV U23519 ( .A(n24120), .Z(n24122) );
  XOR U23520 ( .A(n24126), .B(n24127), .Z(n24120) );
  AND U23521 ( .A(n846), .B(n24119), .Z(n24127) );
  XNOR U23522 ( .A(n24117), .B(n24126), .Z(n24119) );
  XNOR U23523 ( .A(n24128), .B(n24129), .Z(n24117) );
  AND U23524 ( .A(n850), .B(n24130), .Z(n24129) );
  XOR U23525 ( .A(p_input[667]), .B(n24128), .Z(n24130) );
  XNOR U23526 ( .A(n24131), .B(n24132), .Z(n24128) );
  AND U23527 ( .A(n854), .B(n24133), .Z(n24132) );
  XOR U23528 ( .A(n24134), .B(n24135), .Z(n24126) );
  AND U23529 ( .A(n858), .B(n24125), .Z(n24135) );
  XNOR U23530 ( .A(n24136), .B(n24123), .Z(n24125) );
  XOR U23531 ( .A(n24137), .B(n24138), .Z(n24123) );
  AND U23532 ( .A(n881), .B(n24139), .Z(n24138) );
  IV U23533 ( .A(n24134), .Z(n24136) );
  XOR U23534 ( .A(n24140), .B(n24141), .Z(n24134) );
  AND U23535 ( .A(n865), .B(n24133), .Z(n24141) );
  XNOR U23536 ( .A(n24131), .B(n24140), .Z(n24133) );
  XNOR U23537 ( .A(n24142), .B(n24143), .Z(n24131) );
  AND U23538 ( .A(n869), .B(n24144), .Z(n24143) );
  XOR U23539 ( .A(p_input[683]), .B(n24142), .Z(n24144) );
  XNOR U23540 ( .A(n24145), .B(n24146), .Z(n24142) );
  AND U23541 ( .A(n873), .B(n24147), .Z(n24146) );
  XOR U23542 ( .A(n24148), .B(n24149), .Z(n24140) );
  AND U23543 ( .A(n877), .B(n24139), .Z(n24149) );
  XNOR U23544 ( .A(n24150), .B(n24137), .Z(n24139) );
  XOR U23545 ( .A(n24151), .B(n24152), .Z(n24137) );
  AND U23546 ( .A(n900), .B(n24153), .Z(n24152) );
  IV U23547 ( .A(n24148), .Z(n24150) );
  XOR U23548 ( .A(n24154), .B(n24155), .Z(n24148) );
  AND U23549 ( .A(n884), .B(n24147), .Z(n24155) );
  XNOR U23550 ( .A(n24145), .B(n24154), .Z(n24147) );
  XNOR U23551 ( .A(n24156), .B(n24157), .Z(n24145) );
  AND U23552 ( .A(n888), .B(n24158), .Z(n24157) );
  XOR U23553 ( .A(p_input[699]), .B(n24156), .Z(n24158) );
  XNOR U23554 ( .A(n24159), .B(n24160), .Z(n24156) );
  AND U23555 ( .A(n892), .B(n24161), .Z(n24160) );
  XOR U23556 ( .A(n24162), .B(n24163), .Z(n24154) );
  AND U23557 ( .A(n896), .B(n24153), .Z(n24163) );
  XNOR U23558 ( .A(n24164), .B(n24151), .Z(n24153) );
  XOR U23559 ( .A(n24165), .B(n24166), .Z(n24151) );
  AND U23560 ( .A(n919), .B(n24167), .Z(n24166) );
  IV U23561 ( .A(n24162), .Z(n24164) );
  XOR U23562 ( .A(n24168), .B(n24169), .Z(n24162) );
  AND U23563 ( .A(n903), .B(n24161), .Z(n24169) );
  XNOR U23564 ( .A(n24159), .B(n24168), .Z(n24161) );
  XNOR U23565 ( .A(n24170), .B(n24171), .Z(n24159) );
  AND U23566 ( .A(n907), .B(n24172), .Z(n24171) );
  XOR U23567 ( .A(p_input[715]), .B(n24170), .Z(n24172) );
  XNOR U23568 ( .A(n24173), .B(n24174), .Z(n24170) );
  AND U23569 ( .A(n911), .B(n24175), .Z(n24174) );
  XOR U23570 ( .A(n24176), .B(n24177), .Z(n24168) );
  AND U23571 ( .A(n915), .B(n24167), .Z(n24177) );
  XNOR U23572 ( .A(n24178), .B(n24165), .Z(n24167) );
  XOR U23573 ( .A(n24179), .B(n24180), .Z(n24165) );
  AND U23574 ( .A(n938), .B(n24181), .Z(n24180) );
  IV U23575 ( .A(n24176), .Z(n24178) );
  XOR U23576 ( .A(n24182), .B(n24183), .Z(n24176) );
  AND U23577 ( .A(n922), .B(n24175), .Z(n24183) );
  XNOR U23578 ( .A(n24173), .B(n24182), .Z(n24175) );
  XNOR U23579 ( .A(n24184), .B(n24185), .Z(n24173) );
  AND U23580 ( .A(n926), .B(n24186), .Z(n24185) );
  XOR U23581 ( .A(p_input[731]), .B(n24184), .Z(n24186) );
  XNOR U23582 ( .A(n24187), .B(n24188), .Z(n24184) );
  AND U23583 ( .A(n930), .B(n24189), .Z(n24188) );
  XOR U23584 ( .A(n24190), .B(n24191), .Z(n24182) );
  AND U23585 ( .A(n934), .B(n24181), .Z(n24191) );
  XNOR U23586 ( .A(n24192), .B(n24179), .Z(n24181) );
  XOR U23587 ( .A(n24193), .B(n24194), .Z(n24179) );
  AND U23588 ( .A(n957), .B(n24195), .Z(n24194) );
  IV U23589 ( .A(n24190), .Z(n24192) );
  XOR U23590 ( .A(n24196), .B(n24197), .Z(n24190) );
  AND U23591 ( .A(n941), .B(n24189), .Z(n24197) );
  XNOR U23592 ( .A(n24187), .B(n24196), .Z(n24189) );
  XNOR U23593 ( .A(n24198), .B(n24199), .Z(n24187) );
  AND U23594 ( .A(n945), .B(n24200), .Z(n24199) );
  XOR U23595 ( .A(p_input[747]), .B(n24198), .Z(n24200) );
  XNOR U23596 ( .A(n24201), .B(n24202), .Z(n24198) );
  AND U23597 ( .A(n949), .B(n24203), .Z(n24202) );
  XOR U23598 ( .A(n24204), .B(n24205), .Z(n24196) );
  AND U23599 ( .A(n953), .B(n24195), .Z(n24205) );
  XNOR U23600 ( .A(n24206), .B(n24193), .Z(n24195) );
  XOR U23601 ( .A(n24207), .B(n24208), .Z(n24193) );
  AND U23602 ( .A(n976), .B(n24209), .Z(n24208) );
  IV U23603 ( .A(n24204), .Z(n24206) );
  XOR U23604 ( .A(n24210), .B(n24211), .Z(n24204) );
  AND U23605 ( .A(n960), .B(n24203), .Z(n24211) );
  XNOR U23606 ( .A(n24201), .B(n24210), .Z(n24203) );
  XNOR U23607 ( .A(n24212), .B(n24213), .Z(n24201) );
  AND U23608 ( .A(n964), .B(n24214), .Z(n24213) );
  XOR U23609 ( .A(p_input[763]), .B(n24212), .Z(n24214) );
  XNOR U23610 ( .A(n24215), .B(n24216), .Z(n24212) );
  AND U23611 ( .A(n968), .B(n24217), .Z(n24216) );
  XOR U23612 ( .A(n24218), .B(n24219), .Z(n24210) );
  AND U23613 ( .A(n972), .B(n24209), .Z(n24219) );
  XNOR U23614 ( .A(n24220), .B(n24207), .Z(n24209) );
  XOR U23615 ( .A(n24221), .B(n24222), .Z(n24207) );
  AND U23616 ( .A(n995), .B(n24223), .Z(n24222) );
  IV U23617 ( .A(n24218), .Z(n24220) );
  XOR U23618 ( .A(n24224), .B(n24225), .Z(n24218) );
  AND U23619 ( .A(n979), .B(n24217), .Z(n24225) );
  XNOR U23620 ( .A(n24215), .B(n24224), .Z(n24217) );
  XNOR U23621 ( .A(n24226), .B(n24227), .Z(n24215) );
  AND U23622 ( .A(n983), .B(n24228), .Z(n24227) );
  XOR U23623 ( .A(p_input[779]), .B(n24226), .Z(n24228) );
  XNOR U23624 ( .A(n24229), .B(n24230), .Z(n24226) );
  AND U23625 ( .A(n987), .B(n24231), .Z(n24230) );
  XOR U23626 ( .A(n24232), .B(n24233), .Z(n24224) );
  AND U23627 ( .A(n991), .B(n24223), .Z(n24233) );
  XNOR U23628 ( .A(n24234), .B(n24221), .Z(n24223) );
  XOR U23629 ( .A(n24235), .B(n24236), .Z(n24221) );
  AND U23630 ( .A(n1014), .B(n24237), .Z(n24236) );
  IV U23631 ( .A(n24232), .Z(n24234) );
  XOR U23632 ( .A(n24238), .B(n24239), .Z(n24232) );
  AND U23633 ( .A(n998), .B(n24231), .Z(n24239) );
  XNOR U23634 ( .A(n24229), .B(n24238), .Z(n24231) );
  XNOR U23635 ( .A(n24240), .B(n24241), .Z(n24229) );
  AND U23636 ( .A(n1002), .B(n24242), .Z(n24241) );
  XOR U23637 ( .A(p_input[795]), .B(n24240), .Z(n24242) );
  XNOR U23638 ( .A(n24243), .B(n24244), .Z(n24240) );
  AND U23639 ( .A(n1006), .B(n24245), .Z(n24244) );
  XOR U23640 ( .A(n24246), .B(n24247), .Z(n24238) );
  AND U23641 ( .A(n1010), .B(n24237), .Z(n24247) );
  XNOR U23642 ( .A(n24248), .B(n24235), .Z(n24237) );
  XOR U23643 ( .A(n24249), .B(n24250), .Z(n24235) );
  AND U23644 ( .A(n1033), .B(n24251), .Z(n24250) );
  IV U23645 ( .A(n24246), .Z(n24248) );
  XOR U23646 ( .A(n24252), .B(n24253), .Z(n24246) );
  AND U23647 ( .A(n1017), .B(n24245), .Z(n24253) );
  XNOR U23648 ( .A(n24243), .B(n24252), .Z(n24245) );
  XNOR U23649 ( .A(n24254), .B(n24255), .Z(n24243) );
  AND U23650 ( .A(n1021), .B(n24256), .Z(n24255) );
  XOR U23651 ( .A(p_input[811]), .B(n24254), .Z(n24256) );
  XNOR U23652 ( .A(n24257), .B(n24258), .Z(n24254) );
  AND U23653 ( .A(n1025), .B(n24259), .Z(n24258) );
  XOR U23654 ( .A(n24260), .B(n24261), .Z(n24252) );
  AND U23655 ( .A(n1029), .B(n24251), .Z(n24261) );
  XNOR U23656 ( .A(n24262), .B(n24249), .Z(n24251) );
  XOR U23657 ( .A(n24263), .B(n24264), .Z(n24249) );
  AND U23658 ( .A(n1052), .B(n24265), .Z(n24264) );
  IV U23659 ( .A(n24260), .Z(n24262) );
  XOR U23660 ( .A(n24266), .B(n24267), .Z(n24260) );
  AND U23661 ( .A(n1036), .B(n24259), .Z(n24267) );
  XNOR U23662 ( .A(n24257), .B(n24266), .Z(n24259) );
  XNOR U23663 ( .A(n24268), .B(n24269), .Z(n24257) );
  AND U23664 ( .A(n1040), .B(n24270), .Z(n24269) );
  XOR U23665 ( .A(p_input[827]), .B(n24268), .Z(n24270) );
  XNOR U23666 ( .A(n24271), .B(n24272), .Z(n24268) );
  AND U23667 ( .A(n1044), .B(n24273), .Z(n24272) );
  XOR U23668 ( .A(n24274), .B(n24275), .Z(n24266) );
  AND U23669 ( .A(n1048), .B(n24265), .Z(n24275) );
  XNOR U23670 ( .A(n24276), .B(n24263), .Z(n24265) );
  XOR U23671 ( .A(n24277), .B(n24278), .Z(n24263) );
  AND U23672 ( .A(n1071), .B(n24279), .Z(n24278) );
  IV U23673 ( .A(n24274), .Z(n24276) );
  XOR U23674 ( .A(n24280), .B(n24281), .Z(n24274) );
  AND U23675 ( .A(n1055), .B(n24273), .Z(n24281) );
  XNOR U23676 ( .A(n24271), .B(n24280), .Z(n24273) );
  XNOR U23677 ( .A(n24282), .B(n24283), .Z(n24271) );
  AND U23678 ( .A(n1059), .B(n24284), .Z(n24283) );
  XOR U23679 ( .A(p_input[843]), .B(n24282), .Z(n24284) );
  XNOR U23680 ( .A(n24285), .B(n24286), .Z(n24282) );
  AND U23681 ( .A(n1063), .B(n24287), .Z(n24286) );
  XOR U23682 ( .A(n24288), .B(n24289), .Z(n24280) );
  AND U23683 ( .A(n1067), .B(n24279), .Z(n24289) );
  XNOR U23684 ( .A(n24290), .B(n24277), .Z(n24279) );
  XOR U23685 ( .A(n24291), .B(n24292), .Z(n24277) );
  AND U23686 ( .A(n1090), .B(n24293), .Z(n24292) );
  IV U23687 ( .A(n24288), .Z(n24290) );
  XOR U23688 ( .A(n24294), .B(n24295), .Z(n24288) );
  AND U23689 ( .A(n1074), .B(n24287), .Z(n24295) );
  XNOR U23690 ( .A(n24285), .B(n24294), .Z(n24287) );
  XNOR U23691 ( .A(n24296), .B(n24297), .Z(n24285) );
  AND U23692 ( .A(n1078), .B(n24298), .Z(n24297) );
  XOR U23693 ( .A(p_input[859]), .B(n24296), .Z(n24298) );
  XNOR U23694 ( .A(n24299), .B(n24300), .Z(n24296) );
  AND U23695 ( .A(n1082), .B(n24301), .Z(n24300) );
  XOR U23696 ( .A(n24302), .B(n24303), .Z(n24294) );
  AND U23697 ( .A(n1086), .B(n24293), .Z(n24303) );
  XNOR U23698 ( .A(n24304), .B(n24291), .Z(n24293) );
  XOR U23699 ( .A(n24305), .B(n24306), .Z(n24291) );
  AND U23700 ( .A(n1109), .B(n24307), .Z(n24306) );
  IV U23701 ( .A(n24302), .Z(n24304) );
  XOR U23702 ( .A(n24308), .B(n24309), .Z(n24302) );
  AND U23703 ( .A(n1093), .B(n24301), .Z(n24309) );
  XNOR U23704 ( .A(n24299), .B(n24308), .Z(n24301) );
  XNOR U23705 ( .A(n24310), .B(n24311), .Z(n24299) );
  AND U23706 ( .A(n1097), .B(n24312), .Z(n24311) );
  XOR U23707 ( .A(p_input[875]), .B(n24310), .Z(n24312) );
  XNOR U23708 ( .A(n24313), .B(n24314), .Z(n24310) );
  AND U23709 ( .A(n1101), .B(n24315), .Z(n24314) );
  XOR U23710 ( .A(n24316), .B(n24317), .Z(n24308) );
  AND U23711 ( .A(n1105), .B(n24307), .Z(n24317) );
  XNOR U23712 ( .A(n24318), .B(n24305), .Z(n24307) );
  XOR U23713 ( .A(n24319), .B(n24320), .Z(n24305) );
  AND U23714 ( .A(n1128), .B(n24321), .Z(n24320) );
  IV U23715 ( .A(n24316), .Z(n24318) );
  XOR U23716 ( .A(n24322), .B(n24323), .Z(n24316) );
  AND U23717 ( .A(n1112), .B(n24315), .Z(n24323) );
  XNOR U23718 ( .A(n24313), .B(n24322), .Z(n24315) );
  XNOR U23719 ( .A(n24324), .B(n24325), .Z(n24313) );
  AND U23720 ( .A(n1116), .B(n24326), .Z(n24325) );
  XOR U23721 ( .A(p_input[891]), .B(n24324), .Z(n24326) );
  XNOR U23722 ( .A(n24327), .B(n24328), .Z(n24324) );
  AND U23723 ( .A(n1120), .B(n24329), .Z(n24328) );
  XOR U23724 ( .A(n24330), .B(n24331), .Z(n24322) );
  AND U23725 ( .A(n1124), .B(n24321), .Z(n24331) );
  XNOR U23726 ( .A(n24332), .B(n24319), .Z(n24321) );
  XOR U23727 ( .A(n24333), .B(n24334), .Z(n24319) );
  AND U23728 ( .A(n1147), .B(n24335), .Z(n24334) );
  IV U23729 ( .A(n24330), .Z(n24332) );
  XOR U23730 ( .A(n24336), .B(n24337), .Z(n24330) );
  AND U23731 ( .A(n1131), .B(n24329), .Z(n24337) );
  XNOR U23732 ( .A(n24327), .B(n24336), .Z(n24329) );
  XNOR U23733 ( .A(n24338), .B(n24339), .Z(n24327) );
  AND U23734 ( .A(n1135), .B(n24340), .Z(n24339) );
  XOR U23735 ( .A(p_input[907]), .B(n24338), .Z(n24340) );
  XNOR U23736 ( .A(n24341), .B(n24342), .Z(n24338) );
  AND U23737 ( .A(n1139), .B(n24343), .Z(n24342) );
  XOR U23738 ( .A(n24344), .B(n24345), .Z(n24336) );
  AND U23739 ( .A(n1143), .B(n24335), .Z(n24345) );
  XNOR U23740 ( .A(n24346), .B(n24333), .Z(n24335) );
  XOR U23741 ( .A(n24347), .B(n24348), .Z(n24333) );
  AND U23742 ( .A(n1166), .B(n24349), .Z(n24348) );
  IV U23743 ( .A(n24344), .Z(n24346) );
  XOR U23744 ( .A(n24350), .B(n24351), .Z(n24344) );
  AND U23745 ( .A(n1150), .B(n24343), .Z(n24351) );
  XNOR U23746 ( .A(n24341), .B(n24350), .Z(n24343) );
  XNOR U23747 ( .A(n24352), .B(n24353), .Z(n24341) );
  AND U23748 ( .A(n1154), .B(n24354), .Z(n24353) );
  XOR U23749 ( .A(p_input[923]), .B(n24352), .Z(n24354) );
  XNOR U23750 ( .A(n24355), .B(n24356), .Z(n24352) );
  AND U23751 ( .A(n1158), .B(n24357), .Z(n24356) );
  XOR U23752 ( .A(n24358), .B(n24359), .Z(n24350) );
  AND U23753 ( .A(n1162), .B(n24349), .Z(n24359) );
  XNOR U23754 ( .A(n24360), .B(n24347), .Z(n24349) );
  XOR U23755 ( .A(n24361), .B(n24362), .Z(n24347) );
  AND U23756 ( .A(n1185), .B(n24363), .Z(n24362) );
  IV U23757 ( .A(n24358), .Z(n24360) );
  XOR U23758 ( .A(n24364), .B(n24365), .Z(n24358) );
  AND U23759 ( .A(n1169), .B(n24357), .Z(n24365) );
  XNOR U23760 ( .A(n24355), .B(n24364), .Z(n24357) );
  XNOR U23761 ( .A(n24366), .B(n24367), .Z(n24355) );
  AND U23762 ( .A(n1173), .B(n24368), .Z(n24367) );
  XOR U23763 ( .A(p_input[939]), .B(n24366), .Z(n24368) );
  XNOR U23764 ( .A(n24369), .B(n24370), .Z(n24366) );
  AND U23765 ( .A(n1177), .B(n24371), .Z(n24370) );
  XOR U23766 ( .A(n24372), .B(n24373), .Z(n24364) );
  AND U23767 ( .A(n1181), .B(n24363), .Z(n24373) );
  XNOR U23768 ( .A(n24374), .B(n24361), .Z(n24363) );
  XOR U23769 ( .A(n24375), .B(n24376), .Z(n24361) );
  AND U23770 ( .A(n1204), .B(n24377), .Z(n24376) );
  IV U23771 ( .A(n24372), .Z(n24374) );
  XOR U23772 ( .A(n24378), .B(n24379), .Z(n24372) );
  AND U23773 ( .A(n1188), .B(n24371), .Z(n24379) );
  XNOR U23774 ( .A(n24369), .B(n24378), .Z(n24371) );
  XNOR U23775 ( .A(n24380), .B(n24381), .Z(n24369) );
  AND U23776 ( .A(n1192), .B(n24382), .Z(n24381) );
  XOR U23777 ( .A(p_input[955]), .B(n24380), .Z(n24382) );
  XNOR U23778 ( .A(n24383), .B(n24384), .Z(n24380) );
  AND U23779 ( .A(n1196), .B(n24385), .Z(n24384) );
  XOR U23780 ( .A(n24386), .B(n24387), .Z(n24378) );
  AND U23781 ( .A(n1200), .B(n24377), .Z(n24387) );
  XNOR U23782 ( .A(n24388), .B(n24375), .Z(n24377) );
  XOR U23783 ( .A(n24389), .B(n24390), .Z(n24375) );
  AND U23784 ( .A(n1223), .B(n24391), .Z(n24390) );
  IV U23785 ( .A(n24386), .Z(n24388) );
  XOR U23786 ( .A(n24392), .B(n24393), .Z(n24386) );
  AND U23787 ( .A(n1207), .B(n24385), .Z(n24393) );
  XNOR U23788 ( .A(n24383), .B(n24392), .Z(n24385) );
  XNOR U23789 ( .A(n24394), .B(n24395), .Z(n24383) );
  AND U23790 ( .A(n1211), .B(n24396), .Z(n24395) );
  XOR U23791 ( .A(p_input[971]), .B(n24394), .Z(n24396) );
  XNOR U23792 ( .A(n24397), .B(n24398), .Z(n24394) );
  AND U23793 ( .A(n1215), .B(n24399), .Z(n24398) );
  XOR U23794 ( .A(n24400), .B(n24401), .Z(n24392) );
  AND U23795 ( .A(n1219), .B(n24391), .Z(n24401) );
  XNOR U23796 ( .A(n24402), .B(n24389), .Z(n24391) );
  XOR U23797 ( .A(n24403), .B(n24404), .Z(n24389) );
  AND U23798 ( .A(n1242), .B(n24405), .Z(n24404) );
  IV U23799 ( .A(n24400), .Z(n24402) );
  XOR U23800 ( .A(n24406), .B(n24407), .Z(n24400) );
  AND U23801 ( .A(n1226), .B(n24399), .Z(n24407) );
  XNOR U23802 ( .A(n24397), .B(n24406), .Z(n24399) );
  XNOR U23803 ( .A(n24408), .B(n24409), .Z(n24397) );
  AND U23804 ( .A(n1230), .B(n24410), .Z(n24409) );
  XOR U23805 ( .A(p_input[987]), .B(n24408), .Z(n24410) );
  XNOR U23806 ( .A(n24411), .B(n24412), .Z(n24408) );
  AND U23807 ( .A(n1234), .B(n24413), .Z(n24412) );
  XOR U23808 ( .A(n24414), .B(n24415), .Z(n24406) );
  AND U23809 ( .A(n1238), .B(n24405), .Z(n24415) );
  XNOR U23810 ( .A(n24416), .B(n24403), .Z(n24405) );
  XOR U23811 ( .A(n24417), .B(n24418), .Z(n24403) );
  AND U23812 ( .A(n1261), .B(n24419), .Z(n24418) );
  IV U23813 ( .A(n24414), .Z(n24416) );
  XOR U23814 ( .A(n24420), .B(n24421), .Z(n24414) );
  AND U23815 ( .A(n1245), .B(n24413), .Z(n24421) );
  XNOR U23816 ( .A(n24411), .B(n24420), .Z(n24413) );
  XNOR U23817 ( .A(n24422), .B(n24423), .Z(n24411) );
  AND U23818 ( .A(n1249), .B(n24424), .Z(n24423) );
  XOR U23819 ( .A(p_input[1003]), .B(n24422), .Z(n24424) );
  XNOR U23820 ( .A(n24425), .B(n24426), .Z(n24422) );
  AND U23821 ( .A(n1253), .B(n24427), .Z(n24426) );
  XOR U23822 ( .A(n24428), .B(n24429), .Z(n24420) );
  AND U23823 ( .A(n1257), .B(n24419), .Z(n24429) );
  XNOR U23824 ( .A(n24430), .B(n24417), .Z(n24419) );
  XOR U23825 ( .A(n24431), .B(n24432), .Z(n24417) );
  AND U23826 ( .A(n1280), .B(n24433), .Z(n24432) );
  IV U23827 ( .A(n24428), .Z(n24430) );
  XOR U23828 ( .A(n24434), .B(n24435), .Z(n24428) );
  AND U23829 ( .A(n1264), .B(n24427), .Z(n24435) );
  XNOR U23830 ( .A(n24425), .B(n24434), .Z(n24427) );
  XNOR U23831 ( .A(n24436), .B(n24437), .Z(n24425) );
  AND U23832 ( .A(n1268), .B(n24438), .Z(n24437) );
  XOR U23833 ( .A(p_input[1019]), .B(n24436), .Z(n24438) );
  XNOR U23834 ( .A(n24439), .B(n24440), .Z(n24436) );
  AND U23835 ( .A(n1272), .B(n24441), .Z(n24440) );
  XOR U23836 ( .A(n24442), .B(n24443), .Z(n24434) );
  AND U23837 ( .A(n1276), .B(n24433), .Z(n24443) );
  XNOR U23838 ( .A(n24444), .B(n24431), .Z(n24433) );
  XOR U23839 ( .A(n24445), .B(n24446), .Z(n24431) );
  AND U23840 ( .A(n1299), .B(n24447), .Z(n24446) );
  IV U23841 ( .A(n24442), .Z(n24444) );
  XOR U23842 ( .A(n24448), .B(n24449), .Z(n24442) );
  AND U23843 ( .A(n1283), .B(n24441), .Z(n24449) );
  XNOR U23844 ( .A(n24439), .B(n24448), .Z(n24441) );
  XNOR U23845 ( .A(n24450), .B(n24451), .Z(n24439) );
  AND U23846 ( .A(n1287), .B(n24452), .Z(n24451) );
  XOR U23847 ( .A(p_input[1035]), .B(n24450), .Z(n24452) );
  XNOR U23848 ( .A(n24453), .B(n24454), .Z(n24450) );
  AND U23849 ( .A(n1291), .B(n24455), .Z(n24454) );
  XOR U23850 ( .A(n24456), .B(n24457), .Z(n24448) );
  AND U23851 ( .A(n1295), .B(n24447), .Z(n24457) );
  XNOR U23852 ( .A(n24458), .B(n24445), .Z(n24447) );
  XOR U23853 ( .A(n24459), .B(n24460), .Z(n24445) );
  AND U23854 ( .A(n1318), .B(n24461), .Z(n24460) );
  IV U23855 ( .A(n24456), .Z(n24458) );
  XOR U23856 ( .A(n24462), .B(n24463), .Z(n24456) );
  AND U23857 ( .A(n1302), .B(n24455), .Z(n24463) );
  XNOR U23858 ( .A(n24453), .B(n24462), .Z(n24455) );
  XNOR U23859 ( .A(n24464), .B(n24465), .Z(n24453) );
  AND U23860 ( .A(n1306), .B(n24466), .Z(n24465) );
  XOR U23861 ( .A(p_input[1051]), .B(n24464), .Z(n24466) );
  XNOR U23862 ( .A(n24467), .B(n24468), .Z(n24464) );
  AND U23863 ( .A(n1310), .B(n24469), .Z(n24468) );
  XOR U23864 ( .A(n24470), .B(n24471), .Z(n24462) );
  AND U23865 ( .A(n1314), .B(n24461), .Z(n24471) );
  XNOR U23866 ( .A(n24472), .B(n24459), .Z(n24461) );
  XOR U23867 ( .A(n24473), .B(n24474), .Z(n24459) );
  AND U23868 ( .A(n1337), .B(n24475), .Z(n24474) );
  IV U23869 ( .A(n24470), .Z(n24472) );
  XOR U23870 ( .A(n24476), .B(n24477), .Z(n24470) );
  AND U23871 ( .A(n1321), .B(n24469), .Z(n24477) );
  XNOR U23872 ( .A(n24467), .B(n24476), .Z(n24469) );
  XNOR U23873 ( .A(n24478), .B(n24479), .Z(n24467) );
  AND U23874 ( .A(n1325), .B(n24480), .Z(n24479) );
  XOR U23875 ( .A(p_input[1067]), .B(n24478), .Z(n24480) );
  XNOR U23876 ( .A(n24481), .B(n24482), .Z(n24478) );
  AND U23877 ( .A(n1329), .B(n24483), .Z(n24482) );
  XOR U23878 ( .A(n24484), .B(n24485), .Z(n24476) );
  AND U23879 ( .A(n1333), .B(n24475), .Z(n24485) );
  XNOR U23880 ( .A(n24486), .B(n24473), .Z(n24475) );
  XOR U23881 ( .A(n24487), .B(n24488), .Z(n24473) );
  AND U23882 ( .A(n1356), .B(n24489), .Z(n24488) );
  IV U23883 ( .A(n24484), .Z(n24486) );
  XOR U23884 ( .A(n24490), .B(n24491), .Z(n24484) );
  AND U23885 ( .A(n1340), .B(n24483), .Z(n24491) );
  XNOR U23886 ( .A(n24481), .B(n24490), .Z(n24483) );
  XNOR U23887 ( .A(n24492), .B(n24493), .Z(n24481) );
  AND U23888 ( .A(n1344), .B(n24494), .Z(n24493) );
  XOR U23889 ( .A(p_input[1083]), .B(n24492), .Z(n24494) );
  XNOR U23890 ( .A(n24495), .B(n24496), .Z(n24492) );
  AND U23891 ( .A(n1348), .B(n24497), .Z(n24496) );
  XOR U23892 ( .A(n24498), .B(n24499), .Z(n24490) );
  AND U23893 ( .A(n1352), .B(n24489), .Z(n24499) );
  XNOR U23894 ( .A(n24500), .B(n24487), .Z(n24489) );
  XOR U23895 ( .A(n24501), .B(n24502), .Z(n24487) );
  AND U23896 ( .A(n1375), .B(n24503), .Z(n24502) );
  IV U23897 ( .A(n24498), .Z(n24500) );
  XOR U23898 ( .A(n24504), .B(n24505), .Z(n24498) );
  AND U23899 ( .A(n1359), .B(n24497), .Z(n24505) );
  XNOR U23900 ( .A(n24495), .B(n24504), .Z(n24497) );
  XNOR U23901 ( .A(n24506), .B(n24507), .Z(n24495) );
  AND U23902 ( .A(n1363), .B(n24508), .Z(n24507) );
  XOR U23903 ( .A(p_input[1099]), .B(n24506), .Z(n24508) );
  XNOR U23904 ( .A(n24509), .B(n24510), .Z(n24506) );
  AND U23905 ( .A(n1367), .B(n24511), .Z(n24510) );
  XOR U23906 ( .A(n24512), .B(n24513), .Z(n24504) );
  AND U23907 ( .A(n1371), .B(n24503), .Z(n24513) );
  XNOR U23908 ( .A(n24514), .B(n24501), .Z(n24503) );
  XOR U23909 ( .A(n24515), .B(n24516), .Z(n24501) );
  AND U23910 ( .A(n1394), .B(n24517), .Z(n24516) );
  IV U23911 ( .A(n24512), .Z(n24514) );
  XOR U23912 ( .A(n24518), .B(n24519), .Z(n24512) );
  AND U23913 ( .A(n1378), .B(n24511), .Z(n24519) );
  XNOR U23914 ( .A(n24509), .B(n24518), .Z(n24511) );
  XNOR U23915 ( .A(n24520), .B(n24521), .Z(n24509) );
  AND U23916 ( .A(n1382), .B(n24522), .Z(n24521) );
  XOR U23917 ( .A(p_input[1115]), .B(n24520), .Z(n24522) );
  XNOR U23918 ( .A(n24523), .B(n24524), .Z(n24520) );
  AND U23919 ( .A(n1386), .B(n24525), .Z(n24524) );
  XOR U23920 ( .A(n24526), .B(n24527), .Z(n24518) );
  AND U23921 ( .A(n1390), .B(n24517), .Z(n24527) );
  XNOR U23922 ( .A(n24528), .B(n24515), .Z(n24517) );
  XOR U23923 ( .A(n24529), .B(n24530), .Z(n24515) );
  AND U23924 ( .A(n1413), .B(n24531), .Z(n24530) );
  IV U23925 ( .A(n24526), .Z(n24528) );
  XOR U23926 ( .A(n24532), .B(n24533), .Z(n24526) );
  AND U23927 ( .A(n1397), .B(n24525), .Z(n24533) );
  XNOR U23928 ( .A(n24523), .B(n24532), .Z(n24525) );
  XNOR U23929 ( .A(n24534), .B(n24535), .Z(n24523) );
  AND U23930 ( .A(n1401), .B(n24536), .Z(n24535) );
  XOR U23931 ( .A(p_input[1131]), .B(n24534), .Z(n24536) );
  XNOR U23932 ( .A(n24537), .B(n24538), .Z(n24534) );
  AND U23933 ( .A(n1405), .B(n24539), .Z(n24538) );
  XOR U23934 ( .A(n24540), .B(n24541), .Z(n24532) );
  AND U23935 ( .A(n1409), .B(n24531), .Z(n24541) );
  XNOR U23936 ( .A(n24542), .B(n24529), .Z(n24531) );
  XOR U23937 ( .A(n24543), .B(n24544), .Z(n24529) );
  AND U23938 ( .A(n1432), .B(n24545), .Z(n24544) );
  IV U23939 ( .A(n24540), .Z(n24542) );
  XOR U23940 ( .A(n24546), .B(n24547), .Z(n24540) );
  AND U23941 ( .A(n1416), .B(n24539), .Z(n24547) );
  XNOR U23942 ( .A(n24537), .B(n24546), .Z(n24539) );
  XNOR U23943 ( .A(n24548), .B(n24549), .Z(n24537) );
  AND U23944 ( .A(n1420), .B(n24550), .Z(n24549) );
  XOR U23945 ( .A(p_input[1147]), .B(n24548), .Z(n24550) );
  XNOR U23946 ( .A(n24551), .B(n24552), .Z(n24548) );
  AND U23947 ( .A(n1424), .B(n24553), .Z(n24552) );
  XOR U23948 ( .A(n24554), .B(n24555), .Z(n24546) );
  AND U23949 ( .A(n1428), .B(n24545), .Z(n24555) );
  XNOR U23950 ( .A(n24556), .B(n24543), .Z(n24545) );
  XOR U23951 ( .A(n24557), .B(n24558), .Z(n24543) );
  AND U23952 ( .A(n1451), .B(n24559), .Z(n24558) );
  IV U23953 ( .A(n24554), .Z(n24556) );
  XOR U23954 ( .A(n24560), .B(n24561), .Z(n24554) );
  AND U23955 ( .A(n1435), .B(n24553), .Z(n24561) );
  XNOR U23956 ( .A(n24551), .B(n24560), .Z(n24553) );
  XNOR U23957 ( .A(n24562), .B(n24563), .Z(n24551) );
  AND U23958 ( .A(n1439), .B(n24564), .Z(n24563) );
  XOR U23959 ( .A(p_input[1163]), .B(n24562), .Z(n24564) );
  XNOR U23960 ( .A(n24565), .B(n24566), .Z(n24562) );
  AND U23961 ( .A(n1443), .B(n24567), .Z(n24566) );
  XOR U23962 ( .A(n24568), .B(n24569), .Z(n24560) );
  AND U23963 ( .A(n1447), .B(n24559), .Z(n24569) );
  XNOR U23964 ( .A(n24570), .B(n24557), .Z(n24559) );
  XOR U23965 ( .A(n24571), .B(n24572), .Z(n24557) );
  AND U23966 ( .A(n1470), .B(n24573), .Z(n24572) );
  IV U23967 ( .A(n24568), .Z(n24570) );
  XOR U23968 ( .A(n24574), .B(n24575), .Z(n24568) );
  AND U23969 ( .A(n1454), .B(n24567), .Z(n24575) );
  XNOR U23970 ( .A(n24565), .B(n24574), .Z(n24567) );
  XNOR U23971 ( .A(n24576), .B(n24577), .Z(n24565) );
  AND U23972 ( .A(n1458), .B(n24578), .Z(n24577) );
  XOR U23973 ( .A(p_input[1179]), .B(n24576), .Z(n24578) );
  XNOR U23974 ( .A(n24579), .B(n24580), .Z(n24576) );
  AND U23975 ( .A(n1462), .B(n24581), .Z(n24580) );
  XOR U23976 ( .A(n24582), .B(n24583), .Z(n24574) );
  AND U23977 ( .A(n1466), .B(n24573), .Z(n24583) );
  XNOR U23978 ( .A(n24584), .B(n24571), .Z(n24573) );
  XOR U23979 ( .A(n24585), .B(n24586), .Z(n24571) );
  AND U23980 ( .A(n1489), .B(n24587), .Z(n24586) );
  IV U23981 ( .A(n24582), .Z(n24584) );
  XOR U23982 ( .A(n24588), .B(n24589), .Z(n24582) );
  AND U23983 ( .A(n1473), .B(n24581), .Z(n24589) );
  XNOR U23984 ( .A(n24579), .B(n24588), .Z(n24581) );
  XNOR U23985 ( .A(n24590), .B(n24591), .Z(n24579) );
  AND U23986 ( .A(n1477), .B(n24592), .Z(n24591) );
  XOR U23987 ( .A(p_input[1195]), .B(n24590), .Z(n24592) );
  XNOR U23988 ( .A(n24593), .B(n24594), .Z(n24590) );
  AND U23989 ( .A(n1481), .B(n24595), .Z(n24594) );
  XOR U23990 ( .A(n24596), .B(n24597), .Z(n24588) );
  AND U23991 ( .A(n1485), .B(n24587), .Z(n24597) );
  XNOR U23992 ( .A(n24598), .B(n24585), .Z(n24587) );
  XOR U23993 ( .A(n24599), .B(n24600), .Z(n24585) );
  AND U23994 ( .A(n1508), .B(n24601), .Z(n24600) );
  IV U23995 ( .A(n24596), .Z(n24598) );
  XOR U23996 ( .A(n24602), .B(n24603), .Z(n24596) );
  AND U23997 ( .A(n1492), .B(n24595), .Z(n24603) );
  XNOR U23998 ( .A(n24593), .B(n24602), .Z(n24595) );
  XNOR U23999 ( .A(n24604), .B(n24605), .Z(n24593) );
  AND U24000 ( .A(n1496), .B(n24606), .Z(n24605) );
  XOR U24001 ( .A(p_input[1211]), .B(n24604), .Z(n24606) );
  XNOR U24002 ( .A(n24607), .B(n24608), .Z(n24604) );
  AND U24003 ( .A(n1500), .B(n24609), .Z(n24608) );
  XOR U24004 ( .A(n24610), .B(n24611), .Z(n24602) );
  AND U24005 ( .A(n1504), .B(n24601), .Z(n24611) );
  XNOR U24006 ( .A(n24612), .B(n24599), .Z(n24601) );
  XOR U24007 ( .A(n24613), .B(n24614), .Z(n24599) );
  AND U24008 ( .A(n1527), .B(n24615), .Z(n24614) );
  IV U24009 ( .A(n24610), .Z(n24612) );
  XOR U24010 ( .A(n24616), .B(n24617), .Z(n24610) );
  AND U24011 ( .A(n1511), .B(n24609), .Z(n24617) );
  XNOR U24012 ( .A(n24607), .B(n24616), .Z(n24609) );
  XNOR U24013 ( .A(n24618), .B(n24619), .Z(n24607) );
  AND U24014 ( .A(n1515), .B(n24620), .Z(n24619) );
  XOR U24015 ( .A(p_input[1227]), .B(n24618), .Z(n24620) );
  XNOR U24016 ( .A(n24621), .B(n24622), .Z(n24618) );
  AND U24017 ( .A(n1519), .B(n24623), .Z(n24622) );
  XOR U24018 ( .A(n24624), .B(n24625), .Z(n24616) );
  AND U24019 ( .A(n1523), .B(n24615), .Z(n24625) );
  XNOR U24020 ( .A(n24626), .B(n24613), .Z(n24615) );
  XOR U24021 ( .A(n24627), .B(n24628), .Z(n24613) );
  AND U24022 ( .A(n1546), .B(n24629), .Z(n24628) );
  IV U24023 ( .A(n24624), .Z(n24626) );
  XOR U24024 ( .A(n24630), .B(n24631), .Z(n24624) );
  AND U24025 ( .A(n1530), .B(n24623), .Z(n24631) );
  XNOR U24026 ( .A(n24621), .B(n24630), .Z(n24623) );
  XNOR U24027 ( .A(n24632), .B(n24633), .Z(n24621) );
  AND U24028 ( .A(n1534), .B(n24634), .Z(n24633) );
  XOR U24029 ( .A(p_input[1243]), .B(n24632), .Z(n24634) );
  XNOR U24030 ( .A(n24635), .B(n24636), .Z(n24632) );
  AND U24031 ( .A(n1538), .B(n24637), .Z(n24636) );
  XOR U24032 ( .A(n24638), .B(n24639), .Z(n24630) );
  AND U24033 ( .A(n1542), .B(n24629), .Z(n24639) );
  XNOR U24034 ( .A(n24640), .B(n24627), .Z(n24629) );
  XOR U24035 ( .A(n24641), .B(n24642), .Z(n24627) );
  AND U24036 ( .A(n1565), .B(n24643), .Z(n24642) );
  IV U24037 ( .A(n24638), .Z(n24640) );
  XOR U24038 ( .A(n24644), .B(n24645), .Z(n24638) );
  AND U24039 ( .A(n1549), .B(n24637), .Z(n24645) );
  XNOR U24040 ( .A(n24635), .B(n24644), .Z(n24637) );
  XNOR U24041 ( .A(n24646), .B(n24647), .Z(n24635) );
  AND U24042 ( .A(n1553), .B(n24648), .Z(n24647) );
  XOR U24043 ( .A(p_input[1259]), .B(n24646), .Z(n24648) );
  XNOR U24044 ( .A(n24649), .B(n24650), .Z(n24646) );
  AND U24045 ( .A(n1557), .B(n24651), .Z(n24650) );
  XOR U24046 ( .A(n24652), .B(n24653), .Z(n24644) );
  AND U24047 ( .A(n1561), .B(n24643), .Z(n24653) );
  XNOR U24048 ( .A(n24654), .B(n24641), .Z(n24643) );
  XOR U24049 ( .A(n24655), .B(n24656), .Z(n24641) );
  AND U24050 ( .A(n1584), .B(n24657), .Z(n24656) );
  IV U24051 ( .A(n24652), .Z(n24654) );
  XOR U24052 ( .A(n24658), .B(n24659), .Z(n24652) );
  AND U24053 ( .A(n1568), .B(n24651), .Z(n24659) );
  XNOR U24054 ( .A(n24649), .B(n24658), .Z(n24651) );
  XNOR U24055 ( .A(n24660), .B(n24661), .Z(n24649) );
  AND U24056 ( .A(n1572), .B(n24662), .Z(n24661) );
  XOR U24057 ( .A(p_input[1275]), .B(n24660), .Z(n24662) );
  XNOR U24058 ( .A(n24663), .B(n24664), .Z(n24660) );
  AND U24059 ( .A(n1576), .B(n24665), .Z(n24664) );
  XOR U24060 ( .A(n24666), .B(n24667), .Z(n24658) );
  AND U24061 ( .A(n1580), .B(n24657), .Z(n24667) );
  XNOR U24062 ( .A(n24668), .B(n24655), .Z(n24657) );
  XOR U24063 ( .A(n24669), .B(n24670), .Z(n24655) );
  AND U24064 ( .A(n1603), .B(n24671), .Z(n24670) );
  IV U24065 ( .A(n24666), .Z(n24668) );
  XOR U24066 ( .A(n24672), .B(n24673), .Z(n24666) );
  AND U24067 ( .A(n1587), .B(n24665), .Z(n24673) );
  XNOR U24068 ( .A(n24663), .B(n24672), .Z(n24665) );
  XNOR U24069 ( .A(n24674), .B(n24675), .Z(n24663) );
  AND U24070 ( .A(n1591), .B(n24676), .Z(n24675) );
  XOR U24071 ( .A(p_input[1291]), .B(n24674), .Z(n24676) );
  XNOR U24072 ( .A(n24677), .B(n24678), .Z(n24674) );
  AND U24073 ( .A(n1595), .B(n24679), .Z(n24678) );
  XOR U24074 ( .A(n24680), .B(n24681), .Z(n24672) );
  AND U24075 ( .A(n1599), .B(n24671), .Z(n24681) );
  XNOR U24076 ( .A(n24682), .B(n24669), .Z(n24671) );
  XOR U24077 ( .A(n24683), .B(n24684), .Z(n24669) );
  AND U24078 ( .A(n1622), .B(n24685), .Z(n24684) );
  IV U24079 ( .A(n24680), .Z(n24682) );
  XOR U24080 ( .A(n24686), .B(n24687), .Z(n24680) );
  AND U24081 ( .A(n1606), .B(n24679), .Z(n24687) );
  XNOR U24082 ( .A(n24677), .B(n24686), .Z(n24679) );
  XNOR U24083 ( .A(n24688), .B(n24689), .Z(n24677) );
  AND U24084 ( .A(n1610), .B(n24690), .Z(n24689) );
  XOR U24085 ( .A(p_input[1307]), .B(n24688), .Z(n24690) );
  XNOR U24086 ( .A(n24691), .B(n24692), .Z(n24688) );
  AND U24087 ( .A(n1614), .B(n24693), .Z(n24692) );
  XOR U24088 ( .A(n24694), .B(n24695), .Z(n24686) );
  AND U24089 ( .A(n1618), .B(n24685), .Z(n24695) );
  XNOR U24090 ( .A(n24696), .B(n24683), .Z(n24685) );
  XOR U24091 ( .A(n24697), .B(n24698), .Z(n24683) );
  AND U24092 ( .A(n1641), .B(n24699), .Z(n24698) );
  IV U24093 ( .A(n24694), .Z(n24696) );
  XOR U24094 ( .A(n24700), .B(n24701), .Z(n24694) );
  AND U24095 ( .A(n1625), .B(n24693), .Z(n24701) );
  XNOR U24096 ( .A(n24691), .B(n24700), .Z(n24693) );
  XNOR U24097 ( .A(n24702), .B(n24703), .Z(n24691) );
  AND U24098 ( .A(n1629), .B(n24704), .Z(n24703) );
  XOR U24099 ( .A(p_input[1323]), .B(n24702), .Z(n24704) );
  XNOR U24100 ( .A(n24705), .B(n24706), .Z(n24702) );
  AND U24101 ( .A(n1633), .B(n24707), .Z(n24706) );
  XOR U24102 ( .A(n24708), .B(n24709), .Z(n24700) );
  AND U24103 ( .A(n1637), .B(n24699), .Z(n24709) );
  XNOR U24104 ( .A(n24710), .B(n24697), .Z(n24699) );
  XOR U24105 ( .A(n24711), .B(n24712), .Z(n24697) );
  AND U24106 ( .A(n1660), .B(n24713), .Z(n24712) );
  IV U24107 ( .A(n24708), .Z(n24710) );
  XOR U24108 ( .A(n24714), .B(n24715), .Z(n24708) );
  AND U24109 ( .A(n1644), .B(n24707), .Z(n24715) );
  XNOR U24110 ( .A(n24705), .B(n24714), .Z(n24707) );
  XNOR U24111 ( .A(n24716), .B(n24717), .Z(n24705) );
  AND U24112 ( .A(n1648), .B(n24718), .Z(n24717) );
  XOR U24113 ( .A(p_input[1339]), .B(n24716), .Z(n24718) );
  XNOR U24114 ( .A(n24719), .B(n24720), .Z(n24716) );
  AND U24115 ( .A(n1652), .B(n24721), .Z(n24720) );
  XOR U24116 ( .A(n24722), .B(n24723), .Z(n24714) );
  AND U24117 ( .A(n1656), .B(n24713), .Z(n24723) );
  XNOR U24118 ( .A(n24724), .B(n24711), .Z(n24713) );
  XOR U24119 ( .A(n24725), .B(n24726), .Z(n24711) );
  AND U24120 ( .A(n1679), .B(n24727), .Z(n24726) );
  IV U24121 ( .A(n24722), .Z(n24724) );
  XOR U24122 ( .A(n24728), .B(n24729), .Z(n24722) );
  AND U24123 ( .A(n1663), .B(n24721), .Z(n24729) );
  XNOR U24124 ( .A(n24719), .B(n24728), .Z(n24721) );
  XNOR U24125 ( .A(n24730), .B(n24731), .Z(n24719) );
  AND U24126 ( .A(n1667), .B(n24732), .Z(n24731) );
  XOR U24127 ( .A(p_input[1355]), .B(n24730), .Z(n24732) );
  XNOR U24128 ( .A(n24733), .B(n24734), .Z(n24730) );
  AND U24129 ( .A(n1671), .B(n24735), .Z(n24734) );
  XOR U24130 ( .A(n24736), .B(n24737), .Z(n24728) );
  AND U24131 ( .A(n1675), .B(n24727), .Z(n24737) );
  XNOR U24132 ( .A(n24738), .B(n24725), .Z(n24727) );
  XOR U24133 ( .A(n24739), .B(n24740), .Z(n24725) );
  AND U24134 ( .A(n1698), .B(n24741), .Z(n24740) );
  IV U24135 ( .A(n24736), .Z(n24738) );
  XOR U24136 ( .A(n24742), .B(n24743), .Z(n24736) );
  AND U24137 ( .A(n1682), .B(n24735), .Z(n24743) );
  XNOR U24138 ( .A(n24733), .B(n24742), .Z(n24735) );
  XNOR U24139 ( .A(n24744), .B(n24745), .Z(n24733) );
  AND U24140 ( .A(n1686), .B(n24746), .Z(n24745) );
  XOR U24141 ( .A(p_input[1371]), .B(n24744), .Z(n24746) );
  XNOR U24142 ( .A(n24747), .B(n24748), .Z(n24744) );
  AND U24143 ( .A(n1690), .B(n24749), .Z(n24748) );
  XOR U24144 ( .A(n24750), .B(n24751), .Z(n24742) );
  AND U24145 ( .A(n1694), .B(n24741), .Z(n24751) );
  XNOR U24146 ( .A(n24752), .B(n24739), .Z(n24741) );
  XOR U24147 ( .A(n24753), .B(n24754), .Z(n24739) );
  AND U24148 ( .A(n1717), .B(n24755), .Z(n24754) );
  IV U24149 ( .A(n24750), .Z(n24752) );
  XOR U24150 ( .A(n24756), .B(n24757), .Z(n24750) );
  AND U24151 ( .A(n1701), .B(n24749), .Z(n24757) );
  XNOR U24152 ( .A(n24747), .B(n24756), .Z(n24749) );
  XNOR U24153 ( .A(n24758), .B(n24759), .Z(n24747) );
  AND U24154 ( .A(n1705), .B(n24760), .Z(n24759) );
  XOR U24155 ( .A(p_input[1387]), .B(n24758), .Z(n24760) );
  XNOR U24156 ( .A(n24761), .B(n24762), .Z(n24758) );
  AND U24157 ( .A(n1709), .B(n24763), .Z(n24762) );
  XOR U24158 ( .A(n24764), .B(n24765), .Z(n24756) );
  AND U24159 ( .A(n1713), .B(n24755), .Z(n24765) );
  XNOR U24160 ( .A(n24766), .B(n24753), .Z(n24755) );
  XOR U24161 ( .A(n24767), .B(n24768), .Z(n24753) );
  AND U24162 ( .A(n1736), .B(n24769), .Z(n24768) );
  IV U24163 ( .A(n24764), .Z(n24766) );
  XOR U24164 ( .A(n24770), .B(n24771), .Z(n24764) );
  AND U24165 ( .A(n1720), .B(n24763), .Z(n24771) );
  XNOR U24166 ( .A(n24761), .B(n24770), .Z(n24763) );
  XNOR U24167 ( .A(n24772), .B(n24773), .Z(n24761) );
  AND U24168 ( .A(n1724), .B(n24774), .Z(n24773) );
  XOR U24169 ( .A(p_input[1403]), .B(n24772), .Z(n24774) );
  XNOR U24170 ( .A(n24775), .B(n24776), .Z(n24772) );
  AND U24171 ( .A(n1728), .B(n24777), .Z(n24776) );
  XOR U24172 ( .A(n24778), .B(n24779), .Z(n24770) );
  AND U24173 ( .A(n1732), .B(n24769), .Z(n24779) );
  XNOR U24174 ( .A(n24780), .B(n24767), .Z(n24769) );
  XOR U24175 ( .A(n24781), .B(n24782), .Z(n24767) );
  AND U24176 ( .A(n1755), .B(n24783), .Z(n24782) );
  IV U24177 ( .A(n24778), .Z(n24780) );
  XOR U24178 ( .A(n24784), .B(n24785), .Z(n24778) );
  AND U24179 ( .A(n1739), .B(n24777), .Z(n24785) );
  XNOR U24180 ( .A(n24775), .B(n24784), .Z(n24777) );
  XNOR U24181 ( .A(n24786), .B(n24787), .Z(n24775) );
  AND U24182 ( .A(n1743), .B(n24788), .Z(n24787) );
  XOR U24183 ( .A(p_input[1419]), .B(n24786), .Z(n24788) );
  XNOR U24184 ( .A(n24789), .B(n24790), .Z(n24786) );
  AND U24185 ( .A(n1747), .B(n24791), .Z(n24790) );
  XOR U24186 ( .A(n24792), .B(n24793), .Z(n24784) );
  AND U24187 ( .A(n1751), .B(n24783), .Z(n24793) );
  XNOR U24188 ( .A(n24794), .B(n24781), .Z(n24783) );
  XOR U24189 ( .A(n24795), .B(n24796), .Z(n24781) );
  AND U24190 ( .A(n1774), .B(n24797), .Z(n24796) );
  IV U24191 ( .A(n24792), .Z(n24794) );
  XOR U24192 ( .A(n24798), .B(n24799), .Z(n24792) );
  AND U24193 ( .A(n1758), .B(n24791), .Z(n24799) );
  XNOR U24194 ( .A(n24789), .B(n24798), .Z(n24791) );
  XNOR U24195 ( .A(n24800), .B(n24801), .Z(n24789) );
  AND U24196 ( .A(n1762), .B(n24802), .Z(n24801) );
  XOR U24197 ( .A(p_input[1435]), .B(n24800), .Z(n24802) );
  XNOR U24198 ( .A(n24803), .B(n24804), .Z(n24800) );
  AND U24199 ( .A(n1766), .B(n24805), .Z(n24804) );
  XOR U24200 ( .A(n24806), .B(n24807), .Z(n24798) );
  AND U24201 ( .A(n1770), .B(n24797), .Z(n24807) );
  XNOR U24202 ( .A(n24808), .B(n24795), .Z(n24797) );
  XOR U24203 ( .A(n24809), .B(n24810), .Z(n24795) );
  AND U24204 ( .A(n1793), .B(n24811), .Z(n24810) );
  IV U24205 ( .A(n24806), .Z(n24808) );
  XOR U24206 ( .A(n24812), .B(n24813), .Z(n24806) );
  AND U24207 ( .A(n1777), .B(n24805), .Z(n24813) );
  XNOR U24208 ( .A(n24803), .B(n24812), .Z(n24805) );
  XNOR U24209 ( .A(n24814), .B(n24815), .Z(n24803) );
  AND U24210 ( .A(n1781), .B(n24816), .Z(n24815) );
  XOR U24211 ( .A(p_input[1451]), .B(n24814), .Z(n24816) );
  XNOR U24212 ( .A(n24817), .B(n24818), .Z(n24814) );
  AND U24213 ( .A(n1785), .B(n24819), .Z(n24818) );
  XOR U24214 ( .A(n24820), .B(n24821), .Z(n24812) );
  AND U24215 ( .A(n1789), .B(n24811), .Z(n24821) );
  XNOR U24216 ( .A(n24822), .B(n24809), .Z(n24811) );
  XOR U24217 ( .A(n24823), .B(n24824), .Z(n24809) );
  AND U24218 ( .A(n1812), .B(n24825), .Z(n24824) );
  IV U24219 ( .A(n24820), .Z(n24822) );
  XOR U24220 ( .A(n24826), .B(n24827), .Z(n24820) );
  AND U24221 ( .A(n1796), .B(n24819), .Z(n24827) );
  XNOR U24222 ( .A(n24817), .B(n24826), .Z(n24819) );
  XNOR U24223 ( .A(n24828), .B(n24829), .Z(n24817) );
  AND U24224 ( .A(n1800), .B(n24830), .Z(n24829) );
  XOR U24225 ( .A(p_input[1467]), .B(n24828), .Z(n24830) );
  XNOR U24226 ( .A(n24831), .B(n24832), .Z(n24828) );
  AND U24227 ( .A(n1804), .B(n24833), .Z(n24832) );
  XOR U24228 ( .A(n24834), .B(n24835), .Z(n24826) );
  AND U24229 ( .A(n1808), .B(n24825), .Z(n24835) );
  XNOR U24230 ( .A(n24836), .B(n24823), .Z(n24825) );
  XOR U24231 ( .A(n24837), .B(n24838), .Z(n24823) );
  AND U24232 ( .A(n1831), .B(n24839), .Z(n24838) );
  IV U24233 ( .A(n24834), .Z(n24836) );
  XOR U24234 ( .A(n24840), .B(n24841), .Z(n24834) );
  AND U24235 ( .A(n1815), .B(n24833), .Z(n24841) );
  XNOR U24236 ( .A(n24831), .B(n24840), .Z(n24833) );
  XNOR U24237 ( .A(n24842), .B(n24843), .Z(n24831) );
  AND U24238 ( .A(n1819), .B(n24844), .Z(n24843) );
  XOR U24239 ( .A(p_input[1483]), .B(n24842), .Z(n24844) );
  XNOR U24240 ( .A(n24845), .B(n24846), .Z(n24842) );
  AND U24241 ( .A(n1823), .B(n24847), .Z(n24846) );
  XOR U24242 ( .A(n24848), .B(n24849), .Z(n24840) );
  AND U24243 ( .A(n1827), .B(n24839), .Z(n24849) );
  XNOR U24244 ( .A(n24850), .B(n24837), .Z(n24839) );
  XOR U24245 ( .A(n24851), .B(n24852), .Z(n24837) );
  AND U24246 ( .A(n1850), .B(n24853), .Z(n24852) );
  IV U24247 ( .A(n24848), .Z(n24850) );
  XOR U24248 ( .A(n24854), .B(n24855), .Z(n24848) );
  AND U24249 ( .A(n1834), .B(n24847), .Z(n24855) );
  XNOR U24250 ( .A(n24845), .B(n24854), .Z(n24847) );
  XNOR U24251 ( .A(n24856), .B(n24857), .Z(n24845) );
  AND U24252 ( .A(n1838), .B(n24858), .Z(n24857) );
  XOR U24253 ( .A(p_input[1499]), .B(n24856), .Z(n24858) );
  XNOR U24254 ( .A(n24859), .B(n24860), .Z(n24856) );
  AND U24255 ( .A(n1842), .B(n24861), .Z(n24860) );
  XOR U24256 ( .A(n24862), .B(n24863), .Z(n24854) );
  AND U24257 ( .A(n1846), .B(n24853), .Z(n24863) );
  XNOR U24258 ( .A(n24864), .B(n24851), .Z(n24853) );
  XOR U24259 ( .A(n24865), .B(n24866), .Z(n24851) );
  AND U24260 ( .A(n1869), .B(n24867), .Z(n24866) );
  IV U24261 ( .A(n24862), .Z(n24864) );
  XOR U24262 ( .A(n24868), .B(n24869), .Z(n24862) );
  AND U24263 ( .A(n1853), .B(n24861), .Z(n24869) );
  XNOR U24264 ( .A(n24859), .B(n24868), .Z(n24861) );
  XNOR U24265 ( .A(n24870), .B(n24871), .Z(n24859) );
  AND U24266 ( .A(n1857), .B(n24872), .Z(n24871) );
  XOR U24267 ( .A(p_input[1515]), .B(n24870), .Z(n24872) );
  XNOR U24268 ( .A(n24873), .B(n24874), .Z(n24870) );
  AND U24269 ( .A(n1861), .B(n24875), .Z(n24874) );
  XOR U24270 ( .A(n24876), .B(n24877), .Z(n24868) );
  AND U24271 ( .A(n1865), .B(n24867), .Z(n24877) );
  XNOR U24272 ( .A(n24878), .B(n24865), .Z(n24867) );
  XOR U24273 ( .A(n24879), .B(n24880), .Z(n24865) );
  AND U24274 ( .A(n1888), .B(n24881), .Z(n24880) );
  IV U24275 ( .A(n24876), .Z(n24878) );
  XOR U24276 ( .A(n24882), .B(n24883), .Z(n24876) );
  AND U24277 ( .A(n1872), .B(n24875), .Z(n24883) );
  XNOR U24278 ( .A(n24873), .B(n24882), .Z(n24875) );
  XNOR U24279 ( .A(n24884), .B(n24885), .Z(n24873) );
  AND U24280 ( .A(n1876), .B(n24886), .Z(n24885) );
  XOR U24281 ( .A(p_input[1531]), .B(n24884), .Z(n24886) );
  XNOR U24282 ( .A(n24887), .B(n24888), .Z(n24884) );
  AND U24283 ( .A(n1880), .B(n24889), .Z(n24888) );
  XOR U24284 ( .A(n24890), .B(n24891), .Z(n24882) );
  AND U24285 ( .A(n1884), .B(n24881), .Z(n24891) );
  XNOR U24286 ( .A(n24892), .B(n24879), .Z(n24881) );
  XOR U24287 ( .A(n24893), .B(n24894), .Z(n24879) );
  AND U24288 ( .A(n1907), .B(n24895), .Z(n24894) );
  IV U24289 ( .A(n24890), .Z(n24892) );
  XOR U24290 ( .A(n24896), .B(n24897), .Z(n24890) );
  AND U24291 ( .A(n1891), .B(n24889), .Z(n24897) );
  XNOR U24292 ( .A(n24887), .B(n24896), .Z(n24889) );
  XNOR U24293 ( .A(n24898), .B(n24899), .Z(n24887) );
  AND U24294 ( .A(n1895), .B(n24900), .Z(n24899) );
  XOR U24295 ( .A(p_input[1547]), .B(n24898), .Z(n24900) );
  XNOR U24296 ( .A(n24901), .B(n24902), .Z(n24898) );
  AND U24297 ( .A(n1899), .B(n24903), .Z(n24902) );
  XOR U24298 ( .A(n24904), .B(n24905), .Z(n24896) );
  AND U24299 ( .A(n1903), .B(n24895), .Z(n24905) );
  XNOR U24300 ( .A(n24906), .B(n24893), .Z(n24895) );
  XOR U24301 ( .A(n24907), .B(n24908), .Z(n24893) );
  AND U24302 ( .A(n1926), .B(n24909), .Z(n24908) );
  IV U24303 ( .A(n24904), .Z(n24906) );
  XOR U24304 ( .A(n24910), .B(n24911), .Z(n24904) );
  AND U24305 ( .A(n1910), .B(n24903), .Z(n24911) );
  XNOR U24306 ( .A(n24901), .B(n24910), .Z(n24903) );
  XNOR U24307 ( .A(n24912), .B(n24913), .Z(n24901) );
  AND U24308 ( .A(n1914), .B(n24914), .Z(n24913) );
  XOR U24309 ( .A(p_input[1563]), .B(n24912), .Z(n24914) );
  XNOR U24310 ( .A(n24915), .B(n24916), .Z(n24912) );
  AND U24311 ( .A(n1918), .B(n24917), .Z(n24916) );
  XOR U24312 ( .A(n24918), .B(n24919), .Z(n24910) );
  AND U24313 ( .A(n1922), .B(n24909), .Z(n24919) );
  XNOR U24314 ( .A(n24920), .B(n24907), .Z(n24909) );
  XOR U24315 ( .A(n24921), .B(n24922), .Z(n24907) );
  AND U24316 ( .A(n1945), .B(n24923), .Z(n24922) );
  IV U24317 ( .A(n24918), .Z(n24920) );
  XOR U24318 ( .A(n24924), .B(n24925), .Z(n24918) );
  AND U24319 ( .A(n1929), .B(n24917), .Z(n24925) );
  XNOR U24320 ( .A(n24915), .B(n24924), .Z(n24917) );
  XNOR U24321 ( .A(n24926), .B(n24927), .Z(n24915) );
  AND U24322 ( .A(n1933), .B(n24928), .Z(n24927) );
  XOR U24323 ( .A(p_input[1579]), .B(n24926), .Z(n24928) );
  XNOR U24324 ( .A(n24929), .B(n24930), .Z(n24926) );
  AND U24325 ( .A(n1937), .B(n24931), .Z(n24930) );
  XOR U24326 ( .A(n24932), .B(n24933), .Z(n24924) );
  AND U24327 ( .A(n1941), .B(n24923), .Z(n24933) );
  XNOR U24328 ( .A(n24934), .B(n24921), .Z(n24923) );
  XOR U24329 ( .A(n24935), .B(n24936), .Z(n24921) );
  AND U24330 ( .A(n1964), .B(n24937), .Z(n24936) );
  IV U24331 ( .A(n24932), .Z(n24934) );
  XOR U24332 ( .A(n24938), .B(n24939), .Z(n24932) );
  AND U24333 ( .A(n1948), .B(n24931), .Z(n24939) );
  XNOR U24334 ( .A(n24929), .B(n24938), .Z(n24931) );
  XNOR U24335 ( .A(n24940), .B(n24941), .Z(n24929) );
  AND U24336 ( .A(n1952), .B(n24942), .Z(n24941) );
  XOR U24337 ( .A(p_input[1595]), .B(n24940), .Z(n24942) );
  XNOR U24338 ( .A(n24943), .B(n24944), .Z(n24940) );
  AND U24339 ( .A(n1956), .B(n24945), .Z(n24944) );
  XOR U24340 ( .A(n24946), .B(n24947), .Z(n24938) );
  AND U24341 ( .A(n1960), .B(n24937), .Z(n24947) );
  XNOR U24342 ( .A(n24948), .B(n24935), .Z(n24937) );
  XOR U24343 ( .A(n24949), .B(n24950), .Z(n24935) );
  AND U24344 ( .A(n1983), .B(n24951), .Z(n24950) );
  IV U24345 ( .A(n24946), .Z(n24948) );
  XOR U24346 ( .A(n24952), .B(n24953), .Z(n24946) );
  AND U24347 ( .A(n1967), .B(n24945), .Z(n24953) );
  XNOR U24348 ( .A(n24943), .B(n24952), .Z(n24945) );
  XNOR U24349 ( .A(n24954), .B(n24955), .Z(n24943) );
  AND U24350 ( .A(n1971), .B(n24956), .Z(n24955) );
  XOR U24351 ( .A(p_input[1611]), .B(n24954), .Z(n24956) );
  XNOR U24352 ( .A(n24957), .B(n24958), .Z(n24954) );
  AND U24353 ( .A(n1975), .B(n24959), .Z(n24958) );
  XOR U24354 ( .A(n24960), .B(n24961), .Z(n24952) );
  AND U24355 ( .A(n1979), .B(n24951), .Z(n24961) );
  XNOR U24356 ( .A(n24962), .B(n24949), .Z(n24951) );
  XOR U24357 ( .A(n24963), .B(n24964), .Z(n24949) );
  AND U24358 ( .A(n2002), .B(n24965), .Z(n24964) );
  IV U24359 ( .A(n24960), .Z(n24962) );
  XOR U24360 ( .A(n24966), .B(n24967), .Z(n24960) );
  AND U24361 ( .A(n1986), .B(n24959), .Z(n24967) );
  XNOR U24362 ( .A(n24957), .B(n24966), .Z(n24959) );
  XNOR U24363 ( .A(n24968), .B(n24969), .Z(n24957) );
  AND U24364 ( .A(n1990), .B(n24970), .Z(n24969) );
  XOR U24365 ( .A(p_input[1627]), .B(n24968), .Z(n24970) );
  XNOR U24366 ( .A(n24971), .B(n24972), .Z(n24968) );
  AND U24367 ( .A(n1994), .B(n24973), .Z(n24972) );
  XOR U24368 ( .A(n24974), .B(n24975), .Z(n24966) );
  AND U24369 ( .A(n1998), .B(n24965), .Z(n24975) );
  XNOR U24370 ( .A(n24976), .B(n24963), .Z(n24965) );
  XOR U24371 ( .A(n24977), .B(n24978), .Z(n24963) );
  AND U24372 ( .A(n2021), .B(n24979), .Z(n24978) );
  IV U24373 ( .A(n24974), .Z(n24976) );
  XOR U24374 ( .A(n24980), .B(n24981), .Z(n24974) );
  AND U24375 ( .A(n2005), .B(n24973), .Z(n24981) );
  XNOR U24376 ( .A(n24971), .B(n24980), .Z(n24973) );
  XNOR U24377 ( .A(n24982), .B(n24983), .Z(n24971) );
  AND U24378 ( .A(n2009), .B(n24984), .Z(n24983) );
  XOR U24379 ( .A(p_input[1643]), .B(n24982), .Z(n24984) );
  XNOR U24380 ( .A(n24985), .B(n24986), .Z(n24982) );
  AND U24381 ( .A(n2013), .B(n24987), .Z(n24986) );
  XOR U24382 ( .A(n24988), .B(n24989), .Z(n24980) );
  AND U24383 ( .A(n2017), .B(n24979), .Z(n24989) );
  XNOR U24384 ( .A(n24990), .B(n24977), .Z(n24979) );
  XOR U24385 ( .A(n24991), .B(n24992), .Z(n24977) );
  AND U24386 ( .A(n2040), .B(n24993), .Z(n24992) );
  IV U24387 ( .A(n24988), .Z(n24990) );
  XOR U24388 ( .A(n24994), .B(n24995), .Z(n24988) );
  AND U24389 ( .A(n2024), .B(n24987), .Z(n24995) );
  XNOR U24390 ( .A(n24985), .B(n24994), .Z(n24987) );
  XNOR U24391 ( .A(n24996), .B(n24997), .Z(n24985) );
  AND U24392 ( .A(n2028), .B(n24998), .Z(n24997) );
  XOR U24393 ( .A(p_input[1659]), .B(n24996), .Z(n24998) );
  XNOR U24394 ( .A(n24999), .B(n25000), .Z(n24996) );
  AND U24395 ( .A(n2032), .B(n25001), .Z(n25000) );
  XOR U24396 ( .A(n25002), .B(n25003), .Z(n24994) );
  AND U24397 ( .A(n2036), .B(n24993), .Z(n25003) );
  XNOR U24398 ( .A(n25004), .B(n24991), .Z(n24993) );
  XOR U24399 ( .A(n25005), .B(n25006), .Z(n24991) );
  AND U24400 ( .A(n2059), .B(n25007), .Z(n25006) );
  IV U24401 ( .A(n25002), .Z(n25004) );
  XOR U24402 ( .A(n25008), .B(n25009), .Z(n25002) );
  AND U24403 ( .A(n2043), .B(n25001), .Z(n25009) );
  XNOR U24404 ( .A(n24999), .B(n25008), .Z(n25001) );
  XNOR U24405 ( .A(n25010), .B(n25011), .Z(n24999) );
  AND U24406 ( .A(n2047), .B(n25012), .Z(n25011) );
  XOR U24407 ( .A(p_input[1675]), .B(n25010), .Z(n25012) );
  XNOR U24408 ( .A(n25013), .B(n25014), .Z(n25010) );
  AND U24409 ( .A(n2051), .B(n25015), .Z(n25014) );
  XOR U24410 ( .A(n25016), .B(n25017), .Z(n25008) );
  AND U24411 ( .A(n2055), .B(n25007), .Z(n25017) );
  XNOR U24412 ( .A(n25018), .B(n25005), .Z(n25007) );
  XOR U24413 ( .A(n25019), .B(n25020), .Z(n25005) );
  AND U24414 ( .A(n2078), .B(n25021), .Z(n25020) );
  IV U24415 ( .A(n25016), .Z(n25018) );
  XOR U24416 ( .A(n25022), .B(n25023), .Z(n25016) );
  AND U24417 ( .A(n2062), .B(n25015), .Z(n25023) );
  XNOR U24418 ( .A(n25013), .B(n25022), .Z(n25015) );
  XNOR U24419 ( .A(n25024), .B(n25025), .Z(n25013) );
  AND U24420 ( .A(n2066), .B(n25026), .Z(n25025) );
  XOR U24421 ( .A(p_input[1691]), .B(n25024), .Z(n25026) );
  XNOR U24422 ( .A(n25027), .B(n25028), .Z(n25024) );
  AND U24423 ( .A(n2070), .B(n25029), .Z(n25028) );
  XOR U24424 ( .A(n25030), .B(n25031), .Z(n25022) );
  AND U24425 ( .A(n2074), .B(n25021), .Z(n25031) );
  XNOR U24426 ( .A(n25032), .B(n25019), .Z(n25021) );
  XOR U24427 ( .A(n25033), .B(n25034), .Z(n25019) );
  AND U24428 ( .A(n2097), .B(n25035), .Z(n25034) );
  IV U24429 ( .A(n25030), .Z(n25032) );
  XOR U24430 ( .A(n25036), .B(n25037), .Z(n25030) );
  AND U24431 ( .A(n2081), .B(n25029), .Z(n25037) );
  XNOR U24432 ( .A(n25027), .B(n25036), .Z(n25029) );
  XNOR U24433 ( .A(n25038), .B(n25039), .Z(n25027) );
  AND U24434 ( .A(n2085), .B(n25040), .Z(n25039) );
  XOR U24435 ( .A(p_input[1707]), .B(n25038), .Z(n25040) );
  XNOR U24436 ( .A(n25041), .B(n25042), .Z(n25038) );
  AND U24437 ( .A(n2089), .B(n25043), .Z(n25042) );
  XOR U24438 ( .A(n25044), .B(n25045), .Z(n25036) );
  AND U24439 ( .A(n2093), .B(n25035), .Z(n25045) );
  XNOR U24440 ( .A(n25046), .B(n25033), .Z(n25035) );
  XOR U24441 ( .A(n25047), .B(n25048), .Z(n25033) );
  AND U24442 ( .A(n2116), .B(n25049), .Z(n25048) );
  IV U24443 ( .A(n25044), .Z(n25046) );
  XOR U24444 ( .A(n25050), .B(n25051), .Z(n25044) );
  AND U24445 ( .A(n2100), .B(n25043), .Z(n25051) );
  XNOR U24446 ( .A(n25041), .B(n25050), .Z(n25043) );
  XNOR U24447 ( .A(n25052), .B(n25053), .Z(n25041) );
  AND U24448 ( .A(n2104), .B(n25054), .Z(n25053) );
  XOR U24449 ( .A(p_input[1723]), .B(n25052), .Z(n25054) );
  XNOR U24450 ( .A(n25055), .B(n25056), .Z(n25052) );
  AND U24451 ( .A(n2108), .B(n25057), .Z(n25056) );
  XOR U24452 ( .A(n25058), .B(n25059), .Z(n25050) );
  AND U24453 ( .A(n2112), .B(n25049), .Z(n25059) );
  XNOR U24454 ( .A(n25060), .B(n25047), .Z(n25049) );
  XOR U24455 ( .A(n25061), .B(n25062), .Z(n25047) );
  AND U24456 ( .A(n2135), .B(n25063), .Z(n25062) );
  IV U24457 ( .A(n25058), .Z(n25060) );
  XOR U24458 ( .A(n25064), .B(n25065), .Z(n25058) );
  AND U24459 ( .A(n2119), .B(n25057), .Z(n25065) );
  XNOR U24460 ( .A(n25055), .B(n25064), .Z(n25057) );
  XNOR U24461 ( .A(n25066), .B(n25067), .Z(n25055) );
  AND U24462 ( .A(n2123), .B(n25068), .Z(n25067) );
  XOR U24463 ( .A(p_input[1739]), .B(n25066), .Z(n25068) );
  XNOR U24464 ( .A(n25069), .B(n25070), .Z(n25066) );
  AND U24465 ( .A(n2127), .B(n25071), .Z(n25070) );
  XOR U24466 ( .A(n25072), .B(n25073), .Z(n25064) );
  AND U24467 ( .A(n2131), .B(n25063), .Z(n25073) );
  XNOR U24468 ( .A(n25074), .B(n25061), .Z(n25063) );
  XOR U24469 ( .A(n25075), .B(n25076), .Z(n25061) );
  AND U24470 ( .A(n2154), .B(n25077), .Z(n25076) );
  IV U24471 ( .A(n25072), .Z(n25074) );
  XOR U24472 ( .A(n25078), .B(n25079), .Z(n25072) );
  AND U24473 ( .A(n2138), .B(n25071), .Z(n25079) );
  XNOR U24474 ( .A(n25069), .B(n25078), .Z(n25071) );
  XNOR U24475 ( .A(n25080), .B(n25081), .Z(n25069) );
  AND U24476 ( .A(n2142), .B(n25082), .Z(n25081) );
  XOR U24477 ( .A(p_input[1755]), .B(n25080), .Z(n25082) );
  XNOR U24478 ( .A(n25083), .B(n25084), .Z(n25080) );
  AND U24479 ( .A(n2146), .B(n25085), .Z(n25084) );
  XOR U24480 ( .A(n25086), .B(n25087), .Z(n25078) );
  AND U24481 ( .A(n2150), .B(n25077), .Z(n25087) );
  XNOR U24482 ( .A(n25088), .B(n25075), .Z(n25077) );
  XOR U24483 ( .A(n25089), .B(n25090), .Z(n25075) );
  AND U24484 ( .A(n2173), .B(n25091), .Z(n25090) );
  IV U24485 ( .A(n25086), .Z(n25088) );
  XOR U24486 ( .A(n25092), .B(n25093), .Z(n25086) );
  AND U24487 ( .A(n2157), .B(n25085), .Z(n25093) );
  XNOR U24488 ( .A(n25083), .B(n25092), .Z(n25085) );
  XNOR U24489 ( .A(n25094), .B(n25095), .Z(n25083) );
  AND U24490 ( .A(n2161), .B(n25096), .Z(n25095) );
  XOR U24491 ( .A(p_input[1771]), .B(n25094), .Z(n25096) );
  XNOR U24492 ( .A(n25097), .B(n25098), .Z(n25094) );
  AND U24493 ( .A(n2165), .B(n25099), .Z(n25098) );
  XOR U24494 ( .A(n25100), .B(n25101), .Z(n25092) );
  AND U24495 ( .A(n2169), .B(n25091), .Z(n25101) );
  XNOR U24496 ( .A(n25102), .B(n25089), .Z(n25091) );
  XOR U24497 ( .A(n25103), .B(n25104), .Z(n25089) );
  AND U24498 ( .A(n2192), .B(n25105), .Z(n25104) );
  IV U24499 ( .A(n25100), .Z(n25102) );
  XOR U24500 ( .A(n25106), .B(n25107), .Z(n25100) );
  AND U24501 ( .A(n2176), .B(n25099), .Z(n25107) );
  XNOR U24502 ( .A(n25097), .B(n25106), .Z(n25099) );
  XNOR U24503 ( .A(n25108), .B(n25109), .Z(n25097) );
  AND U24504 ( .A(n2180), .B(n25110), .Z(n25109) );
  XOR U24505 ( .A(p_input[1787]), .B(n25108), .Z(n25110) );
  XNOR U24506 ( .A(n25111), .B(n25112), .Z(n25108) );
  AND U24507 ( .A(n2184), .B(n25113), .Z(n25112) );
  XOR U24508 ( .A(n25114), .B(n25115), .Z(n25106) );
  AND U24509 ( .A(n2188), .B(n25105), .Z(n25115) );
  XNOR U24510 ( .A(n25116), .B(n25103), .Z(n25105) );
  XOR U24511 ( .A(n25117), .B(n25118), .Z(n25103) );
  AND U24512 ( .A(n2211), .B(n25119), .Z(n25118) );
  IV U24513 ( .A(n25114), .Z(n25116) );
  XOR U24514 ( .A(n25120), .B(n25121), .Z(n25114) );
  AND U24515 ( .A(n2195), .B(n25113), .Z(n25121) );
  XNOR U24516 ( .A(n25111), .B(n25120), .Z(n25113) );
  XNOR U24517 ( .A(n25122), .B(n25123), .Z(n25111) );
  AND U24518 ( .A(n2199), .B(n25124), .Z(n25123) );
  XOR U24519 ( .A(p_input[1803]), .B(n25122), .Z(n25124) );
  XNOR U24520 ( .A(n25125), .B(n25126), .Z(n25122) );
  AND U24521 ( .A(n2203), .B(n25127), .Z(n25126) );
  XOR U24522 ( .A(n25128), .B(n25129), .Z(n25120) );
  AND U24523 ( .A(n2207), .B(n25119), .Z(n25129) );
  XNOR U24524 ( .A(n25130), .B(n25117), .Z(n25119) );
  XOR U24525 ( .A(n25131), .B(n25132), .Z(n25117) );
  AND U24526 ( .A(n2230), .B(n25133), .Z(n25132) );
  IV U24527 ( .A(n25128), .Z(n25130) );
  XOR U24528 ( .A(n25134), .B(n25135), .Z(n25128) );
  AND U24529 ( .A(n2214), .B(n25127), .Z(n25135) );
  XNOR U24530 ( .A(n25125), .B(n25134), .Z(n25127) );
  XNOR U24531 ( .A(n25136), .B(n25137), .Z(n25125) );
  AND U24532 ( .A(n2218), .B(n25138), .Z(n25137) );
  XOR U24533 ( .A(p_input[1819]), .B(n25136), .Z(n25138) );
  XNOR U24534 ( .A(n25139), .B(n25140), .Z(n25136) );
  AND U24535 ( .A(n2222), .B(n25141), .Z(n25140) );
  XOR U24536 ( .A(n25142), .B(n25143), .Z(n25134) );
  AND U24537 ( .A(n2226), .B(n25133), .Z(n25143) );
  XNOR U24538 ( .A(n25144), .B(n25131), .Z(n25133) );
  XOR U24539 ( .A(n25145), .B(n25146), .Z(n25131) );
  AND U24540 ( .A(n2249), .B(n25147), .Z(n25146) );
  IV U24541 ( .A(n25142), .Z(n25144) );
  XOR U24542 ( .A(n25148), .B(n25149), .Z(n25142) );
  AND U24543 ( .A(n2233), .B(n25141), .Z(n25149) );
  XNOR U24544 ( .A(n25139), .B(n25148), .Z(n25141) );
  XNOR U24545 ( .A(n25150), .B(n25151), .Z(n25139) );
  AND U24546 ( .A(n2237), .B(n25152), .Z(n25151) );
  XOR U24547 ( .A(p_input[1835]), .B(n25150), .Z(n25152) );
  XNOR U24548 ( .A(n25153), .B(n25154), .Z(n25150) );
  AND U24549 ( .A(n2241), .B(n25155), .Z(n25154) );
  XOR U24550 ( .A(n25156), .B(n25157), .Z(n25148) );
  AND U24551 ( .A(n2245), .B(n25147), .Z(n25157) );
  XNOR U24552 ( .A(n25158), .B(n25145), .Z(n25147) );
  XOR U24553 ( .A(n25159), .B(n25160), .Z(n25145) );
  AND U24554 ( .A(n2268), .B(n25161), .Z(n25160) );
  IV U24555 ( .A(n25156), .Z(n25158) );
  XOR U24556 ( .A(n25162), .B(n25163), .Z(n25156) );
  AND U24557 ( .A(n2252), .B(n25155), .Z(n25163) );
  XNOR U24558 ( .A(n25153), .B(n25162), .Z(n25155) );
  XNOR U24559 ( .A(n25164), .B(n25165), .Z(n25153) );
  AND U24560 ( .A(n2256), .B(n25166), .Z(n25165) );
  XOR U24561 ( .A(p_input[1851]), .B(n25164), .Z(n25166) );
  XNOR U24562 ( .A(n25167), .B(n25168), .Z(n25164) );
  AND U24563 ( .A(n2260), .B(n25169), .Z(n25168) );
  XOR U24564 ( .A(n25170), .B(n25171), .Z(n25162) );
  AND U24565 ( .A(n2264), .B(n25161), .Z(n25171) );
  XNOR U24566 ( .A(n25172), .B(n25159), .Z(n25161) );
  XOR U24567 ( .A(n25173), .B(n25174), .Z(n25159) );
  AND U24568 ( .A(n2287), .B(n25175), .Z(n25174) );
  IV U24569 ( .A(n25170), .Z(n25172) );
  XOR U24570 ( .A(n25176), .B(n25177), .Z(n25170) );
  AND U24571 ( .A(n2271), .B(n25169), .Z(n25177) );
  XNOR U24572 ( .A(n25167), .B(n25176), .Z(n25169) );
  XNOR U24573 ( .A(n25178), .B(n25179), .Z(n25167) );
  AND U24574 ( .A(n2275), .B(n25180), .Z(n25179) );
  XOR U24575 ( .A(p_input[1867]), .B(n25178), .Z(n25180) );
  XNOR U24576 ( .A(n25181), .B(n25182), .Z(n25178) );
  AND U24577 ( .A(n2279), .B(n25183), .Z(n25182) );
  XOR U24578 ( .A(n25184), .B(n25185), .Z(n25176) );
  AND U24579 ( .A(n2283), .B(n25175), .Z(n25185) );
  XNOR U24580 ( .A(n25186), .B(n25173), .Z(n25175) );
  XOR U24581 ( .A(n25187), .B(n25188), .Z(n25173) );
  AND U24582 ( .A(n2306), .B(n25189), .Z(n25188) );
  IV U24583 ( .A(n25184), .Z(n25186) );
  XOR U24584 ( .A(n25190), .B(n25191), .Z(n25184) );
  AND U24585 ( .A(n2290), .B(n25183), .Z(n25191) );
  XNOR U24586 ( .A(n25181), .B(n25190), .Z(n25183) );
  XNOR U24587 ( .A(n25192), .B(n25193), .Z(n25181) );
  AND U24588 ( .A(n2294), .B(n25194), .Z(n25193) );
  XOR U24589 ( .A(p_input[1883]), .B(n25192), .Z(n25194) );
  XNOR U24590 ( .A(n25195), .B(n25196), .Z(n25192) );
  AND U24591 ( .A(n2298), .B(n25197), .Z(n25196) );
  XOR U24592 ( .A(n25198), .B(n25199), .Z(n25190) );
  AND U24593 ( .A(n2302), .B(n25189), .Z(n25199) );
  XNOR U24594 ( .A(n25200), .B(n25187), .Z(n25189) );
  XOR U24595 ( .A(n25201), .B(n25202), .Z(n25187) );
  AND U24596 ( .A(n2325), .B(n25203), .Z(n25202) );
  IV U24597 ( .A(n25198), .Z(n25200) );
  XOR U24598 ( .A(n25204), .B(n25205), .Z(n25198) );
  AND U24599 ( .A(n2309), .B(n25197), .Z(n25205) );
  XNOR U24600 ( .A(n25195), .B(n25204), .Z(n25197) );
  XNOR U24601 ( .A(n25206), .B(n25207), .Z(n25195) );
  AND U24602 ( .A(n2313), .B(n25208), .Z(n25207) );
  XOR U24603 ( .A(p_input[1899]), .B(n25206), .Z(n25208) );
  XNOR U24604 ( .A(n25209), .B(n25210), .Z(n25206) );
  AND U24605 ( .A(n2317), .B(n25211), .Z(n25210) );
  XOR U24606 ( .A(n25212), .B(n25213), .Z(n25204) );
  AND U24607 ( .A(n2321), .B(n25203), .Z(n25213) );
  XNOR U24608 ( .A(n25214), .B(n25201), .Z(n25203) );
  XOR U24609 ( .A(n25215), .B(n25216), .Z(n25201) );
  AND U24610 ( .A(n2344), .B(n25217), .Z(n25216) );
  IV U24611 ( .A(n25212), .Z(n25214) );
  XOR U24612 ( .A(n25218), .B(n25219), .Z(n25212) );
  AND U24613 ( .A(n2328), .B(n25211), .Z(n25219) );
  XNOR U24614 ( .A(n25209), .B(n25218), .Z(n25211) );
  XNOR U24615 ( .A(n25220), .B(n25221), .Z(n25209) );
  AND U24616 ( .A(n2332), .B(n25222), .Z(n25221) );
  XOR U24617 ( .A(p_input[1915]), .B(n25220), .Z(n25222) );
  XNOR U24618 ( .A(n25223), .B(n25224), .Z(n25220) );
  AND U24619 ( .A(n2336), .B(n25225), .Z(n25224) );
  XOR U24620 ( .A(n25226), .B(n25227), .Z(n25218) );
  AND U24621 ( .A(n2340), .B(n25217), .Z(n25227) );
  XNOR U24622 ( .A(n25228), .B(n25215), .Z(n25217) );
  XOR U24623 ( .A(n25229), .B(n25230), .Z(n25215) );
  AND U24624 ( .A(n2363), .B(n25231), .Z(n25230) );
  IV U24625 ( .A(n25226), .Z(n25228) );
  XOR U24626 ( .A(n25232), .B(n25233), .Z(n25226) );
  AND U24627 ( .A(n2347), .B(n25225), .Z(n25233) );
  XNOR U24628 ( .A(n25223), .B(n25232), .Z(n25225) );
  XNOR U24629 ( .A(n25234), .B(n25235), .Z(n25223) );
  AND U24630 ( .A(n2351), .B(n25236), .Z(n25235) );
  XOR U24631 ( .A(p_input[1931]), .B(n25234), .Z(n25236) );
  XNOR U24632 ( .A(n25237), .B(n25238), .Z(n25234) );
  AND U24633 ( .A(n2355), .B(n25239), .Z(n25238) );
  XOR U24634 ( .A(n25240), .B(n25241), .Z(n25232) );
  AND U24635 ( .A(n2359), .B(n25231), .Z(n25241) );
  XNOR U24636 ( .A(n25242), .B(n25229), .Z(n25231) );
  XOR U24637 ( .A(n25243), .B(n25244), .Z(n25229) );
  AND U24638 ( .A(n2382), .B(n25245), .Z(n25244) );
  IV U24639 ( .A(n25240), .Z(n25242) );
  XOR U24640 ( .A(n25246), .B(n25247), .Z(n25240) );
  AND U24641 ( .A(n2366), .B(n25239), .Z(n25247) );
  XNOR U24642 ( .A(n25237), .B(n25246), .Z(n25239) );
  XNOR U24643 ( .A(n25248), .B(n25249), .Z(n25237) );
  AND U24644 ( .A(n2370), .B(n25250), .Z(n25249) );
  XOR U24645 ( .A(p_input[1947]), .B(n25248), .Z(n25250) );
  XNOR U24646 ( .A(n25251), .B(n25252), .Z(n25248) );
  AND U24647 ( .A(n2374), .B(n25253), .Z(n25252) );
  XOR U24648 ( .A(n25254), .B(n25255), .Z(n25246) );
  AND U24649 ( .A(n2378), .B(n25245), .Z(n25255) );
  XNOR U24650 ( .A(n25256), .B(n25243), .Z(n25245) );
  XOR U24651 ( .A(n25257), .B(n25258), .Z(n25243) );
  AND U24652 ( .A(n2401), .B(n25259), .Z(n25258) );
  IV U24653 ( .A(n25254), .Z(n25256) );
  XOR U24654 ( .A(n25260), .B(n25261), .Z(n25254) );
  AND U24655 ( .A(n2385), .B(n25253), .Z(n25261) );
  XNOR U24656 ( .A(n25251), .B(n25260), .Z(n25253) );
  XNOR U24657 ( .A(n25262), .B(n25263), .Z(n25251) );
  AND U24658 ( .A(n2389), .B(n25264), .Z(n25263) );
  XOR U24659 ( .A(p_input[1963]), .B(n25262), .Z(n25264) );
  XNOR U24660 ( .A(n25265), .B(n25266), .Z(n25262) );
  AND U24661 ( .A(n2393), .B(n25267), .Z(n25266) );
  XOR U24662 ( .A(n25268), .B(n25269), .Z(n25260) );
  AND U24663 ( .A(n2397), .B(n25259), .Z(n25269) );
  XNOR U24664 ( .A(n25270), .B(n25257), .Z(n25259) );
  XOR U24665 ( .A(n25271), .B(n25272), .Z(n25257) );
  AND U24666 ( .A(n2420), .B(n25273), .Z(n25272) );
  IV U24667 ( .A(n25268), .Z(n25270) );
  XOR U24668 ( .A(n25274), .B(n25275), .Z(n25268) );
  AND U24669 ( .A(n2404), .B(n25267), .Z(n25275) );
  XNOR U24670 ( .A(n25265), .B(n25274), .Z(n25267) );
  XNOR U24671 ( .A(n25276), .B(n25277), .Z(n25265) );
  AND U24672 ( .A(n2408), .B(n25278), .Z(n25277) );
  XOR U24673 ( .A(p_input[1979]), .B(n25276), .Z(n25278) );
  XNOR U24674 ( .A(n25279), .B(n25280), .Z(n25276) );
  AND U24675 ( .A(n2412), .B(n25281), .Z(n25280) );
  XOR U24676 ( .A(n25282), .B(n25283), .Z(n25274) );
  AND U24677 ( .A(n2416), .B(n25273), .Z(n25283) );
  XNOR U24678 ( .A(n25284), .B(n25271), .Z(n25273) );
  XOR U24679 ( .A(n25285), .B(n25286), .Z(n25271) );
  AND U24680 ( .A(n2438), .B(n25287), .Z(n25286) );
  IV U24681 ( .A(n25282), .Z(n25284) );
  XOR U24682 ( .A(n25288), .B(n25289), .Z(n25282) );
  AND U24683 ( .A(n2423), .B(n25281), .Z(n25289) );
  XNOR U24684 ( .A(n25279), .B(n25288), .Z(n25281) );
  XNOR U24685 ( .A(n25290), .B(n25291), .Z(n25279) );
  AND U24686 ( .A(n2427), .B(n25292), .Z(n25291) );
  XOR U24687 ( .A(p_input[1995]), .B(n25290), .Z(n25292) );
  XOR U24688 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n25293), 
        .Z(n25290) );
  AND U24689 ( .A(n2430), .B(n25294), .Z(n25293) );
  XOR U24690 ( .A(n25295), .B(n25296), .Z(n25288) );
  AND U24691 ( .A(n2434), .B(n25287), .Z(n25296) );
  XNOR U24692 ( .A(n25297), .B(n25285), .Z(n25287) );
  XOR U24693 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n25298), .Z(n25285) );
  AND U24694 ( .A(n2446), .B(n25299), .Z(n25298) );
  IV U24695 ( .A(n25295), .Z(n25297) );
  XOR U24696 ( .A(n25300), .B(n25301), .Z(n25295) );
  AND U24697 ( .A(n2441), .B(n25294), .Z(n25301) );
  XOR U24698 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n25300), 
        .Z(n25294) );
  XOR U24699 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n25302), 
        .Z(n25300) );
  AND U24700 ( .A(n2443), .B(n25299), .Z(n25302) );
  XOR U24701 ( .A(n25303), .B(n25304), .Z(n25299) );
  IV U24702 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n25304)
         );
  IV U24703 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n25303) );
  XOR U24704 ( .A(n59), .B(n25305), .Z(o[10]) );
  AND U24705 ( .A(n62), .B(n25306), .Z(n59) );
  XOR U24706 ( .A(n60), .B(n25305), .Z(n25306) );
  XOR U24707 ( .A(n25307), .B(n25308), .Z(n25305) );
  AND U24708 ( .A(n82), .B(n25309), .Z(n25308) );
  XOR U24709 ( .A(n25310), .B(n23), .Z(n60) );
  AND U24710 ( .A(n65), .B(n25311), .Z(n23) );
  XOR U24711 ( .A(n24), .B(n25310), .Z(n25311) );
  XOR U24712 ( .A(n25312), .B(n25313), .Z(n24) );
  AND U24713 ( .A(n70), .B(n25314), .Z(n25313) );
  XOR U24714 ( .A(p_input[10]), .B(n25312), .Z(n25314) );
  XNOR U24715 ( .A(n25315), .B(n25316), .Z(n25312) );
  AND U24716 ( .A(n74), .B(n25317), .Z(n25316) );
  XOR U24717 ( .A(n25318), .B(n25319), .Z(n25310) );
  AND U24718 ( .A(n78), .B(n25309), .Z(n25319) );
  XNOR U24719 ( .A(n25320), .B(n25307), .Z(n25309) );
  XOR U24720 ( .A(n25321), .B(n25322), .Z(n25307) );
  AND U24721 ( .A(n102), .B(n25323), .Z(n25322) );
  IV U24722 ( .A(n25318), .Z(n25320) );
  XOR U24723 ( .A(n25324), .B(n25325), .Z(n25318) );
  AND U24724 ( .A(n86), .B(n25317), .Z(n25325) );
  XNOR U24725 ( .A(n25315), .B(n25324), .Z(n25317) );
  XNOR U24726 ( .A(n25326), .B(n25327), .Z(n25315) );
  AND U24727 ( .A(n90), .B(n25328), .Z(n25327) );
  XOR U24728 ( .A(p_input[26]), .B(n25326), .Z(n25328) );
  XNOR U24729 ( .A(n25329), .B(n25330), .Z(n25326) );
  AND U24730 ( .A(n94), .B(n25331), .Z(n25330) );
  XOR U24731 ( .A(n25332), .B(n25333), .Z(n25324) );
  AND U24732 ( .A(n98), .B(n25323), .Z(n25333) );
  XNOR U24733 ( .A(n25334), .B(n25321), .Z(n25323) );
  XOR U24734 ( .A(n25335), .B(n25336), .Z(n25321) );
  AND U24735 ( .A(n121), .B(n25337), .Z(n25336) );
  IV U24736 ( .A(n25332), .Z(n25334) );
  XOR U24737 ( .A(n25338), .B(n25339), .Z(n25332) );
  AND U24738 ( .A(n105), .B(n25331), .Z(n25339) );
  XNOR U24739 ( .A(n25329), .B(n25338), .Z(n25331) );
  XNOR U24740 ( .A(n25340), .B(n25341), .Z(n25329) );
  AND U24741 ( .A(n109), .B(n25342), .Z(n25341) );
  XOR U24742 ( .A(p_input[42]), .B(n25340), .Z(n25342) );
  XNOR U24743 ( .A(n25343), .B(n25344), .Z(n25340) );
  AND U24744 ( .A(n113), .B(n25345), .Z(n25344) );
  XOR U24745 ( .A(n25346), .B(n25347), .Z(n25338) );
  AND U24746 ( .A(n117), .B(n25337), .Z(n25347) );
  XNOR U24747 ( .A(n25348), .B(n25335), .Z(n25337) );
  XOR U24748 ( .A(n25349), .B(n25350), .Z(n25335) );
  AND U24749 ( .A(n140), .B(n25351), .Z(n25350) );
  IV U24750 ( .A(n25346), .Z(n25348) );
  XOR U24751 ( .A(n25352), .B(n25353), .Z(n25346) );
  AND U24752 ( .A(n124), .B(n25345), .Z(n25353) );
  XNOR U24753 ( .A(n25343), .B(n25352), .Z(n25345) );
  XNOR U24754 ( .A(n25354), .B(n25355), .Z(n25343) );
  AND U24755 ( .A(n128), .B(n25356), .Z(n25355) );
  XOR U24756 ( .A(p_input[58]), .B(n25354), .Z(n25356) );
  XNOR U24757 ( .A(n25357), .B(n25358), .Z(n25354) );
  AND U24758 ( .A(n132), .B(n25359), .Z(n25358) );
  XOR U24759 ( .A(n25360), .B(n25361), .Z(n25352) );
  AND U24760 ( .A(n136), .B(n25351), .Z(n25361) );
  XNOR U24761 ( .A(n25362), .B(n25349), .Z(n25351) );
  XOR U24762 ( .A(n25363), .B(n25364), .Z(n25349) );
  AND U24763 ( .A(n159), .B(n25365), .Z(n25364) );
  IV U24764 ( .A(n25360), .Z(n25362) );
  XOR U24765 ( .A(n25366), .B(n25367), .Z(n25360) );
  AND U24766 ( .A(n143), .B(n25359), .Z(n25367) );
  XNOR U24767 ( .A(n25357), .B(n25366), .Z(n25359) );
  XNOR U24768 ( .A(n25368), .B(n25369), .Z(n25357) );
  AND U24769 ( .A(n147), .B(n25370), .Z(n25369) );
  XOR U24770 ( .A(p_input[74]), .B(n25368), .Z(n25370) );
  XNOR U24771 ( .A(n25371), .B(n25372), .Z(n25368) );
  AND U24772 ( .A(n151), .B(n25373), .Z(n25372) );
  XOR U24773 ( .A(n25374), .B(n25375), .Z(n25366) );
  AND U24774 ( .A(n155), .B(n25365), .Z(n25375) );
  XNOR U24775 ( .A(n25376), .B(n25363), .Z(n25365) );
  XOR U24776 ( .A(n25377), .B(n25378), .Z(n25363) );
  AND U24777 ( .A(n178), .B(n25379), .Z(n25378) );
  IV U24778 ( .A(n25374), .Z(n25376) );
  XOR U24779 ( .A(n25380), .B(n25381), .Z(n25374) );
  AND U24780 ( .A(n162), .B(n25373), .Z(n25381) );
  XNOR U24781 ( .A(n25371), .B(n25380), .Z(n25373) );
  XNOR U24782 ( .A(n25382), .B(n25383), .Z(n25371) );
  AND U24783 ( .A(n166), .B(n25384), .Z(n25383) );
  XOR U24784 ( .A(p_input[90]), .B(n25382), .Z(n25384) );
  XNOR U24785 ( .A(n25385), .B(n25386), .Z(n25382) );
  AND U24786 ( .A(n170), .B(n25387), .Z(n25386) );
  XOR U24787 ( .A(n25388), .B(n25389), .Z(n25380) );
  AND U24788 ( .A(n174), .B(n25379), .Z(n25389) );
  XNOR U24789 ( .A(n25390), .B(n25377), .Z(n25379) );
  XOR U24790 ( .A(n25391), .B(n25392), .Z(n25377) );
  AND U24791 ( .A(n197), .B(n25393), .Z(n25392) );
  IV U24792 ( .A(n25388), .Z(n25390) );
  XOR U24793 ( .A(n25394), .B(n25395), .Z(n25388) );
  AND U24794 ( .A(n181), .B(n25387), .Z(n25395) );
  XNOR U24795 ( .A(n25385), .B(n25394), .Z(n25387) );
  XNOR U24796 ( .A(n25396), .B(n25397), .Z(n25385) );
  AND U24797 ( .A(n185), .B(n25398), .Z(n25397) );
  XOR U24798 ( .A(p_input[106]), .B(n25396), .Z(n25398) );
  XNOR U24799 ( .A(n25399), .B(n25400), .Z(n25396) );
  AND U24800 ( .A(n189), .B(n25401), .Z(n25400) );
  XOR U24801 ( .A(n25402), .B(n25403), .Z(n25394) );
  AND U24802 ( .A(n193), .B(n25393), .Z(n25403) );
  XNOR U24803 ( .A(n25404), .B(n25391), .Z(n25393) );
  XOR U24804 ( .A(n25405), .B(n25406), .Z(n25391) );
  AND U24805 ( .A(n216), .B(n25407), .Z(n25406) );
  IV U24806 ( .A(n25402), .Z(n25404) );
  XOR U24807 ( .A(n25408), .B(n25409), .Z(n25402) );
  AND U24808 ( .A(n200), .B(n25401), .Z(n25409) );
  XNOR U24809 ( .A(n25399), .B(n25408), .Z(n25401) );
  XNOR U24810 ( .A(n25410), .B(n25411), .Z(n25399) );
  AND U24811 ( .A(n204), .B(n25412), .Z(n25411) );
  XOR U24812 ( .A(p_input[122]), .B(n25410), .Z(n25412) );
  XNOR U24813 ( .A(n25413), .B(n25414), .Z(n25410) );
  AND U24814 ( .A(n208), .B(n25415), .Z(n25414) );
  XOR U24815 ( .A(n25416), .B(n25417), .Z(n25408) );
  AND U24816 ( .A(n212), .B(n25407), .Z(n25417) );
  XNOR U24817 ( .A(n25418), .B(n25405), .Z(n25407) );
  XOR U24818 ( .A(n25419), .B(n25420), .Z(n25405) );
  AND U24819 ( .A(n235), .B(n25421), .Z(n25420) );
  IV U24820 ( .A(n25416), .Z(n25418) );
  XOR U24821 ( .A(n25422), .B(n25423), .Z(n25416) );
  AND U24822 ( .A(n219), .B(n25415), .Z(n25423) );
  XNOR U24823 ( .A(n25413), .B(n25422), .Z(n25415) );
  XNOR U24824 ( .A(n25424), .B(n25425), .Z(n25413) );
  AND U24825 ( .A(n223), .B(n25426), .Z(n25425) );
  XOR U24826 ( .A(p_input[138]), .B(n25424), .Z(n25426) );
  XNOR U24827 ( .A(n25427), .B(n25428), .Z(n25424) );
  AND U24828 ( .A(n227), .B(n25429), .Z(n25428) );
  XOR U24829 ( .A(n25430), .B(n25431), .Z(n25422) );
  AND U24830 ( .A(n231), .B(n25421), .Z(n25431) );
  XNOR U24831 ( .A(n25432), .B(n25419), .Z(n25421) );
  XOR U24832 ( .A(n25433), .B(n25434), .Z(n25419) );
  AND U24833 ( .A(n254), .B(n25435), .Z(n25434) );
  IV U24834 ( .A(n25430), .Z(n25432) );
  XOR U24835 ( .A(n25436), .B(n25437), .Z(n25430) );
  AND U24836 ( .A(n238), .B(n25429), .Z(n25437) );
  XNOR U24837 ( .A(n25427), .B(n25436), .Z(n25429) );
  XNOR U24838 ( .A(n25438), .B(n25439), .Z(n25427) );
  AND U24839 ( .A(n242), .B(n25440), .Z(n25439) );
  XOR U24840 ( .A(p_input[154]), .B(n25438), .Z(n25440) );
  XNOR U24841 ( .A(n25441), .B(n25442), .Z(n25438) );
  AND U24842 ( .A(n246), .B(n25443), .Z(n25442) );
  XOR U24843 ( .A(n25444), .B(n25445), .Z(n25436) );
  AND U24844 ( .A(n250), .B(n25435), .Z(n25445) );
  XNOR U24845 ( .A(n25446), .B(n25433), .Z(n25435) );
  XOR U24846 ( .A(n25447), .B(n25448), .Z(n25433) );
  AND U24847 ( .A(n273), .B(n25449), .Z(n25448) );
  IV U24848 ( .A(n25444), .Z(n25446) );
  XOR U24849 ( .A(n25450), .B(n25451), .Z(n25444) );
  AND U24850 ( .A(n257), .B(n25443), .Z(n25451) );
  XNOR U24851 ( .A(n25441), .B(n25450), .Z(n25443) );
  XNOR U24852 ( .A(n25452), .B(n25453), .Z(n25441) );
  AND U24853 ( .A(n261), .B(n25454), .Z(n25453) );
  XOR U24854 ( .A(p_input[170]), .B(n25452), .Z(n25454) );
  XNOR U24855 ( .A(n25455), .B(n25456), .Z(n25452) );
  AND U24856 ( .A(n265), .B(n25457), .Z(n25456) );
  XOR U24857 ( .A(n25458), .B(n25459), .Z(n25450) );
  AND U24858 ( .A(n269), .B(n25449), .Z(n25459) );
  XNOR U24859 ( .A(n25460), .B(n25447), .Z(n25449) );
  XOR U24860 ( .A(n25461), .B(n25462), .Z(n25447) );
  AND U24861 ( .A(n292), .B(n25463), .Z(n25462) );
  IV U24862 ( .A(n25458), .Z(n25460) );
  XOR U24863 ( .A(n25464), .B(n25465), .Z(n25458) );
  AND U24864 ( .A(n276), .B(n25457), .Z(n25465) );
  XNOR U24865 ( .A(n25455), .B(n25464), .Z(n25457) );
  XNOR U24866 ( .A(n25466), .B(n25467), .Z(n25455) );
  AND U24867 ( .A(n280), .B(n25468), .Z(n25467) );
  XOR U24868 ( .A(p_input[186]), .B(n25466), .Z(n25468) );
  XNOR U24869 ( .A(n25469), .B(n25470), .Z(n25466) );
  AND U24870 ( .A(n284), .B(n25471), .Z(n25470) );
  XOR U24871 ( .A(n25472), .B(n25473), .Z(n25464) );
  AND U24872 ( .A(n288), .B(n25463), .Z(n25473) );
  XNOR U24873 ( .A(n25474), .B(n25461), .Z(n25463) );
  XOR U24874 ( .A(n25475), .B(n25476), .Z(n25461) );
  AND U24875 ( .A(n311), .B(n25477), .Z(n25476) );
  IV U24876 ( .A(n25472), .Z(n25474) );
  XOR U24877 ( .A(n25478), .B(n25479), .Z(n25472) );
  AND U24878 ( .A(n295), .B(n25471), .Z(n25479) );
  XNOR U24879 ( .A(n25469), .B(n25478), .Z(n25471) );
  XNOR U24880 ( .A(n25480), .B(n25481), .Z(n25469) );
  AND U24881 ( .A(n299), .B(n25482), .Z(n25481) );
  XOR U24882 ( .A(p_input[202]), .B(n25480), .Z(n25482) );
  XNOR U24883 ( .A(n25483), .B(n25484), .Z(n25480) );
  AND U24884 ( .A(n303), .B(n25485), .Z(n25484) );
  XOR U24885 ( .A(n25486), .B(n25487), .Z(n25478) );
  AND U24886 ( .A(n307), .B(n25477), .Z(n25487) );
  XNOR U24887 ( .A(n25488), .B(n25475), .Z(n25477) );
  XOR U24888 ( .A(n25489), .B(n25490), .Z(n25475) );
  AND U24889 ( .A(n330), .B(n25491), .Z(n25490) );
  IV U24890 ( .A(n25486), .Z(n25488) );
  XOR U24891 ( .A(n25492), .B(n25493), .Z(n25486) );
  AND U24892 ( .A(n314), .B(n25485), .Z(n25493) );
  XNOR U24893 ( .A(n25483), .B(n25492), .Z(n25485) );
  XNOR U24894 ( .A(n25494), .B(n25495), .Z(n25483) );
  AND U24895 ( .A(n318), .B(n25496), .Z(n25495) );
  XOR U24896 ( .A(p_input[218]), .B(n25494), .Z(n25496) );
  XNOR U24897 ( .A(n25497), .B(n25498), .Z(n25494) );
  AND U24898 ( .A(n322), .B(n25499), .Z(n25498) );
  XOR U24899 ( .A(n25500), .B(n25501), .Z(n25492) );
  AND U24900 ( .A(n326), .B(n25491), .Z(n25501) );
  XNOR U24901 ( .A(n25502), .B(n25489), .Z(n25491) );
  XOR U24902 ( .A(n25503), .B(n25504), .Z(n25489) );
  AND U24903 ( .A(n349), .B(n25505), .Z(n25504) );
  IV U24904 ( .A(n25500), .Z(n25502) );
  XOR U24905 ( .A(n25506), .B(n25507), .Z(n25500) );
  AND U24906 ( .A(n333), .B(n25499), .Z(n25507) );
  XNOR U24907 ( .A(n25497), .B(n25506), .Z(n25499) );
  XNOR U24908 ( .A(n25508), .B(n25509), .Z(n25497) );
  AND U24909 ( .A(n337), .B(n25510), .Z(n25509) );
  XOR U24910 ( .A(p_input[234]), .B(n25508), .Z(n25510) );
  XNOR U24911 ( .A(n25511), .B(n25512), .Z(n25508) );
  AND U24912 ( .A(n341), .B(n25513), .Z(n25512) );
  XOR U24913 ( .A(n25514), .B(n25515), .Z(n25506) );
  AND U24914 ( .A(n345), .B(n25505), .Z(n25515) );
  XNOR U24915 ( .A(n25516), .B(n25503), .Z(n25505) );
  XOR U24916 ( .A(n25517), .B(n25518), .Z(n25503) );
  AND U24917 ( .A(n368), .B(n25519), .Z(n25518) );
  IV U24918 ( .A(n25514), .Z(n25516) );
  XOR U24919 ( .A(n25520), .B(n25521), .Z(n25514) );
  AND U24920 ( .A(n352), .B(n25513), .Z(n25521) );
  XNOR U24921 ( .A(n25511), .B(n25520), .Z(n25513) );
  XNOR U24922 ( .A(n25522), .B(n25523), .Z(n25511) );
  AND U24923 ( .A(n356), .B(n25524), .Z(n25523) );
  XOR U24924 ( .A(p_input[250]), .B(n25522), .Z(n25524) );
  XNOR U24925 ( .A(n25525), .B(n25526), .Z(n25522) );
  AND U24926 ( .A(n360), .B(n25527), .Z(n25526) );
  XOR U24927 ( .A(n25528), .B(n25529), .Z(n25520) );
  AND U24928 ( .A(n364), .B(n25519), .Z(n25529) );
  XNOR U24929 ( .A(n25530), .B(n25517), .Z(n25519) );
  XOR U24930 ( .A(n25531), .B(n25532), .Z(n25517) );
  AND U24931 ( .A(n387), .B(n25533), .Z(n25532) );
  IV U24932 ( .A(n25528), .Z(n25530) );
  XOR U24933 ( .A(n25534), .B(n25535), .Z(n25528) );
  AND U24934 ( .A(n371), .B(n25527), .Z(n25535) );
  XNOR U24935 ( .A(n25525), .B(n25534), .Z(n25527) );
  XNOR U24936 ( .A(n25536), .B(n25537), .Z(n25525) );
  AND U24937 ( .A(n375), .B(n25538), .Z(n25537) );
  XOR U24938 ( .A(p_input[266]), .B(n25536), .Z(n25538) );
  XNOR U24939 ( .A(n25539), .B(n25540), .Z(n25536) );
  AND U24940 ( .A(n379), .B(n25541), .Z(n25540) );
  XOR U24941 ( .A(n25542), .B(n25543), .Z(n25534) );
  AND U24942 ( .A(n383), .B(n25533), .Z(n25543) );
  XNOR U24943 ( .A(n25544), .B(n25531), .Z(n25533) );
  XOR U24944 ( .A(n25545), .B(n25546), .Z(n25531) );
  AND U24945 ( .A(n406), .B(n25547), .Z(n25546) );
  IV U24946 ( .A(n25542), .Z(n25544) );
  XOR U24947 ( .A(n25548), .B(n25549), .Z(n25542) );
  AND U24948 ( .A(n390), .B(n25541), .Z(n25549) );
  XNOR U24949 ( .A(n25539), .B(n25548), .Z(n25541) );
  XNOR U24950 ( .A(n25550), .B(n25551), .Z(n25539) );
  AND U24951 ( .A(n394), .B(n25552), .Z(n25551) );
  XOR U24952 ( .A(p_input[282]), .B(n25550), .Z(n25552) );
  XNOR U24953 ( .A(n25553), .B(n25554), .Z(n25550) );
  AND U24954 ( .A(n398), .B(n25555), .Z(n25554) );
  XOR U24955 ( .A(n25556), .B(n25557), .Z(n25548) );
  AND U24956 ( .A(n402), .B(n25547), .Z(n25557) );
  XNOR U24957 ( .A(n25558), .B(n25545), .Z(n25547) );
  XOR U24958 ( .A(n25559), .B(n25560), .Z(n25545) );
  AND U24959 ( .A(n425), .B(n25561), .Z(n25560) );
  IV U24960 ( .A(n25556), .Z(n25558) );
  XOR U24961 ( .A(n25562), .B(n25563), .Z(n25556) );
  AND U24962 ( .A(n409), .B(n25555), .Z(n25563) );
  XNOR U24963 ( .A(n25553), .B(n25562), .Z(n25555) );
  XNOR U24964 ( .A(n25564), .B(n25565), .Z(n25553) );
  AND U24965 ( .A(n413), .B(n25566), .Z(n25565) );
  XOR U24966 ( .A(p_input[298]), .B(n25564), .Z(n25566) );
  XNOR U24967 ( .A(n25567), .B(n25568), .Z(n25564) );
  AND U24968 ( .A(n417), .B(n25569), .Z(n25568) );
  XOR U24969 ( .A(n25570), .B(n25571), .Z(n25562) );
  AND U24970 ( .A(n421), .B(n25561), .Z(n25571) );
  XNOR U24971 ( .A(n25572), .B(n25559), .Z(n25561) );
  XOR U24972 ( .A(n25573), .B(n25574), .Z(n25559) );
  AND U24973 ( .A(n444), .B(n25575), .Z(n25574) );
  IV U24974 ( .A(n25570), .Z(n25572) );
  XOR U24975 ( .A(n25576), .B(n25577), .Z(n25570) );
  AND U24976 ( .A(n428), .B(n25569), .Z(n25577) );
  XNOR U24977 ( .A(n25567), .B(n25576), .Z(n25569) );
  XNOR U24978 ( .A(n25578), .B(n25579), .Z(n25567) );
  AND U24979 ( .A(n432), .B(n25580), .Z(n25579) );
  XOR U24980 ( .A(p_input[314]), .B(n25578), .Z(n25580) );
  XNOR U24981 ( .A(n25581), .B(n25582), .Z(n25578) );
  AND U24982 ( .A(n436), .B(n25583), .Z(n25582) );
  XOR U24983 ( .A(n25584), .B(n25585), .Z(n25576) );
  AND U24984 ( .A(n440), .B(n25575), .Z(n25585) );
  XNOR U24985 ( .A(n25586), .B(n25573), .Z(n25575) );
  XOR U24986 ( .A(n25587), .B(n25588), .Z(n25573) );
  AND U24987 ( .A(n463), .B(n25589), .Z(n25588) );
  IV U24988 ( .A(n25584), .Z(n25586) );
  XOR U24989 ( .A(n25590), .B(n25591), .Z(n25584) );
  AND U24990 ( .A(n447), .B(n25583), .Z(n25591) );
  XNOR U24991 ( .A(n25581), .B(n25590), .Z(n25583) );
  XNOR U24992 ( .A(n25592), .B(n25593), .Z(n25581) );
  AND U24993 ( .A(n451), .B(n25594), .Z(n25593) );
  XOR U24994 ( .A(p_input[330]), .B(n25592), .Z(n25594) );
  XNOR U24995 ( .A(n25595), .B(n25596), .Z(n25592) );
  AND U24996 ( .A(n455), .B(n25597), .Z(n25596) );
  XOR U24997 ( .A(n25598), .B(n25599), .Z(n25590) );
  AND U24998 ( .A(n459), .B(n25589), .Z(n25599) );
  XNOR U24999 ( .A(n25600), .B(n25587), .Z(n25589) );
  XOR U25000 ( .A(n25601), .B(n25602), .Z(n25587) );
  AND U25001 ( .A(n482), .B(n25603), .Z(n25602) );
  IV U25002 ( .A(n25598), .Z(n25600) );
  XOR U25003 ( .A(n25604), .B(n25605), .Z(n25598) );
  AND U25004 ( .A(n466), .B(n25597), .Z(n25605) );
  XNOR U25005 ( .A(n25595), .B(n25604), .Z(n25597) );
  XNOR U25006 ( .A(n25606), .B(n25607), .Z(n25595) );
  AND U25007 ( .A(n470), .B(n25608), .Z(n25607) );
  XOR U25008 ( .A(p_input[346]), .B(n25606), .Z(n25608) );
  XNOR U25009 ( .A(n25609), .B(n25610), .Z(n25606) );
  AND U25010 ( .A(n474), .B(n25611), .Z(n25610) );
  XOR U25011 ( .A(n25612), .B(n25613), .Z(n25604) );
  AND U25012 ( .A(n478), .B(n25603), .Z(n25613) );
  XNOR U25013 ( .A(n25614), .B(n25601), .Z(n25603) );
  XOR U25014 ( .A(n25615), .B(n25616), .Z(n25601) );
  AND U25015 ( .A(n501), .B(n25617), .Z(n25616) );
  IV U25016 ( .A(n25612), .Z(n25614) );
  XOR U25017 ( .A(n25618), .B(n25619), .Z(n25612) );
  AND U25018 ( .A(n485), .B(n25611), .Z(n25619) );
  XNOR U25019 ( .A(n25609), .B(n25618), .Z(n25611) );
  XNOR U25020 ( .A(n25620), .B(n25621), .Z(n25609) );
  AND U25021 ( .A(n489), .B(n25622), .Z(n25621) );
  XOR U25022 ( .A(p_input[362]), .B(n25620), .Z(n25622) );
  XNOR U25023 ( .A(n25623), .B(n25624), .Z(n25620) );
  AND U25024 ( .A(n493), .B(n25625), .Z(n25624) );
  XOR U25025 ( .A(n25626), .B(n25627), .Z(n25618) );
  AND U25026 ( .A(n497), .B(n25617), .Z(n25627) );
  XNOR U25027 ( .A(n25628), .B(n25615), .Z(n25617) );
  XOR U25028 ( .A(n25629), .B(n25630), .Z(n25615) );
  AND U25029 ( .A(n520), .B(n25631), .Z(n25630) );
  IV U25030 ( .A(n25626), .Z(n25628) );
  XOR U25031 ( .A(n25632), .B(n25633), .Z(n25626) );
  AND U25032 ( .A(n504), .B(n25625), .Z(n25633) );
  XNOR U25033 ( .A(n25623), .B(n25632), .Z(n25625) );
  XNOR U25034 ( .A(n25634), .B(n25635), .Z(n25623) );
  AND U25035 ( .A(n508), .B(n25636), .Z(n25635) );
  XOR U25036 ( .A(p_input[378]), .B(n25634), .Z(n25636) );
  XNOR U25037 ( .A(n25637), .B(n25638), .Z(n25634) );
  AND U25038 ( .A(n512), .B(n25639), .Z(n25638) );
  XOR U25039 ( .A(n25640), .B(n25641), .Z(n25632) );
  AND U25040 ( .A(n516), .B(n25631), .Z(n25641) );
  XNOR U25041 ( .A(n25642), .B(n25629), .Z(n25631) );
  XOR U25042 ( .A(n25643), .B(n25644), .Z(n25629) );
  AND U25043 ( .A(n539), .B(n25645), .Z(n25644) );
  IV U25044 ( .A(n25640), .Z(n25642) );
  XOR U25045 ( .A(n25646), .B(n25647), .Z(n25640) );
  AND U25046 ( .A(n523), .B(n25639), .Z(n25647) );
  XNOR U25047 ( .A(n25637), .B(n25646), .Z(n25639) );
  XNOR U25048 ( .A(n25648), .B(n25649), .Z(n25637) );
  AND U25049 ( .A(n527), .B(n25650), .Z(n25649) );
  XOR U25050 ( .A(p_input[394]), .B(n25648), .Z(n25650) );
  XNOR U25051 ( .A(n25651), .B(n25652), .Z(n25648) );
  AND U25052 ( .A(n531), .B(n25653), .Z(n25652) );
  XOR U25053 ( .A(n25654), .B(n25655), .Z(n25646) );
  AND U25054 ( .A(n535), .B(n25645), .Z(n25655) );
  XNOR U25055 ( .A(n25656), .B(n25643), .Z(n25645) );
  XOR U25056 ( .A(n25657), .B(n25658), .Z(n25643) );
  AND U25057 ( .A(n558), .B(n25659), .Z(n25658) );
  IV U25058 ( .A(n25654), .Z(n25656) );
  XOR U25059 ( .A(n25660), .B(n25661), .Z(n25654) );
  AND U25060 ( .A(n542), .B(n25653), .Z(n25661) );
  XNOR U25061 ( .A(n25651), .B(n25660), .Z(n25653) );
  XNOR U25062 ( .A(n25662), .B(n25663), .Z(n25651) );
  AND U25063 ( .A(n546), .B(n25664), .Z(n25663) );
  XOR U25064 ( .A(p_input[410]), .B(n25662), .Z(n25664) );
  XNOR U25065 ( .A(n25665), .B(n25666), .Z(n25662) );
  AND U25066 ( .A(n550), .B(n25667), .Z(n25666) );
  XOR U25067 ( .A(n25668), .B(n25669), .Z(n25660) );
  AND U25068 ( .A(n554), .B(n25659), .Z(n25669) );
  XNOR U25069 ( .A(n25670), .B(n25657), .Z(n25659) );
  XOR U25070 ( .A(n25671), .B(n25672), .Z(n25657) );
  AND U25071 ( .A(n577), .B(n25673), .Z(n25672) );
  IV U25072 ( .A(n25668), .Z(n25670) );
  XOR U25073 ( .A(n25674), .B(n25675), .Z(n25668) );
  AND U25074 ( .A(n561), .B(n25667), .Z(n25675) );
  XNOR U25075 ( .A(n25665), .B(n25674), .Z(n25667) );
  XNOR U25076 ( .A(n25676), .B(n25677), .Z(n25665) );
  AND U25077 ( .A(n565), .B(n25678), .Z(n25677) );
  XOR U25078 ( .A(p_input[426]), .B(n25676), .Z(n25678) );
  XNOR U25079 ( .A(n25679), .B(n25680), .Z(n25676) );
  AND U25080 ( .A(n569), .B(n25681), .Z(n25680) );
  XOR U25081 ( .A(n25682), .B(n25683), .Z(n25674) );
  AND U25082 ( .A(n573), .B(n25673), .Z(n25683) );
  XNOR U25083 ( .A(n25684), .B(n25671), .Z(n25673) );
  XOR U25084 ( .A(n25685), .B(n25686), .Z(n25671) );
  AND U25085 ( .A(n596), .B(n25687), .Z(n25686) );
  IV U25086 ( .A(n25682), .Z(n25684) );
  XOR U25087 ( .A(n25688), .B(n25689), .Z(n25682) );
  AND U25088 ( .A(n580), .B(n25681), .Z(n25689) );
  XNOR U25089 ( .A(n25679), .B(n25688), .Z(n25681) );
  XNOR U25090 ( .A(n25690), .B(n25691), .Z(n25679) );
  AND U25091 ( .A(n584), .B(n25692), .Z(n25691) );
  XOR U25092 ( .A(p_input[442]), .B(n25690), .Z(n25692) );
  XNOR U25093 ( .A(n25693), .B(n25694), .Z(n25690) );
  AND U25094 ( .A(n588), .B(n25695), .Z(n25694) );
  XOR U25095 ( .A(n25696), .B(n25697), .Z(n25688) );
  AND U25096 ( .A(n592), .B(n25687), .Z(n25697) );
  XNOR U25097 ( .A(n25698), .B(n25685), .Z(n25687) );
  XOR U25098 ( .A(n25699), .B(n25700), .Z(n25685) );
  AND U25099 ( .A(n615), .B(n25701), .Z(n25700) );
  IV U25100 ( .A(n25696), .Z(n25698) );
  XOR U25101 ( .A(n25702), .B(n25703), .Z(n25696) );
  AND U25102 ( .A(n599), .B(n25695), .Z(n25703) );
  XNOR U25103 ( .A(n25693), .B(n25702), .Z(n25695) );
  XNOR U25104 ( .A(n25704), .B(n25705), .Z(n25693) );
  AND U25105 ( .A(n603), .B(n25706), .Z(n25705) );
  XOR U25106 ( .A(p_input[458]), .B(n25704), .Z(n25706) );
  XNOR U25107 ( .A(n25707), .B(n25708), .Z(n25704) );
  AND U25108 ( .A(n607), .B(n25709), .Z(n25708) );
  XOR U25109 ( .A(n25710), .B(n25711), .Z(n25702) );
  AND U25110 ( .A(n611), .B(n25701), .Z(n25711) );
  XNOR U25111 ( .A(n25712), .B(n25699), .Z(n25701) );
  XOR U25112 ( .A(n25713), .B(n25714), .Z(n25699) );
  AND U25113 ( .A(n634), .B(n25715), .Z(n25714) );
  IV U25114 ( .A(n25710), .Z(n25712) );
  XOR U25115 ( .A(n25716), .B(n25717), .Z(n25710) );
  AND U25116 ( .A(n618), .B(n25709), .Z(n25717) );
  XNOR U25117 ( .A(n25707), .B(n25716), .Z(n25709) );
  XNOR U25118 ( .A(n25718), .B(n25719), .Z(n25707) );
  AND U25119 ( .A(n622), .B(n25720), .Z(n25719) );
  XOR U25120 ( .A(p_input[474]), .B(n25718), .Z(n25720) );
  XNOR U25121 ( .A(n25721), .B(n25722), .Z(n25718) );
  AND U25122 ( .A(n626), .B(n25723), .Z(n25722) );
  XOR U25123 ( .A(n25724), .B(n25725), .Z(n25716) );
  AND U25124 ( .A(n630), .B(n25715), .Z(n25725) );
  XNOR U25125 ( .A(n25726), .B(n25713), .Z(n25715) );
  XOR U25126 ( .A(n25727), .B(n25728), .Z(n25713) );
  AND U25127 ( .A(n653), .B(n25729), .Z(n25728) );
  IV U25128 ( .A(n25724), .Z(n25726) );
  XOR U25129 ( .A(n25730), .B(n25731), .Z(n25724) );
  AND U25130 ( .A(n637), .B(n25723), .Z(n25731) );
  XNOR U25131 ( .A(n25721), .B(n25730), .Z(n25723) );
  XNOR U25132 ( .A(n25732), .B(n25733), .Z(n25721) );
  AND U25133 ( .A(n641), .B(n25734), .Z(n25733) );
  XOR U25134 ( .A(p_input[490]), .B(n25732), .Z(n25734) );
  XNOR U25135 ( .A(n25735), .B(n25736), .Z(n25732) );
  AND U25136 ( .A(n645), .B(n25737), .Z(n25736) );
  XOR U25137 ( .A(n25738), .B(n25739), .Z(n25730) );
  AND U25138 ( .A(n649), .B(n25729), .Z(n25739) );
  XNOR U25139 ( .A(n25740), .B(n25727), .Z(n25729) );
  XOR U25140 ( .A(n25741), .B(n25742), .Z(n25727) );
  AND U25141 ( .A(n672), .B(n25743), .Z(n25742) );
  IV U25142 ( .A(n25738), .Z(n25740) );
  XOR U25143 ( .A(n25744), .B(n25745), .Z(n25738) );
  AND U25144 ( .A(n656), .B(n25737), .Z(n25745) );
  XNOR U25145 ( .A(n25735), .B(n25744), .Z(n25737) );
  XNOR U25146 ( .A(n25746), .B(n25747), .Z(n25735) );
  AND U25147 ( .A(n660), .B(n25748), .Z(n25747) );
  XOR U25148 ( .A(p_input[506]), .B(n25746), .Z(n25748) );
  XNOR U25149 ( .A(n25749), .B(n25750), .Z(n25746) );
  AND U25150 ( .A(n664), .B(n25751), .Z(n25750) );
  XOR U25151 ( .A(n25752), .B(n25753), .Z(n25744) );
  AND U25152 ( .A(n668), .B(n25743), .Z(n25753) );
  XNOR U25153 ( .A(n25754), .B(n25741), .Z(n25743) );
  XOR U25154 ( .A(n25755), .B(n25756), .Z(n25741) );
  AND U25155 ( .A(n691), .B(n25757), .Z(n25756) );
  IV U25156 ( .A(n25752), .Z(n25754) );
  XOR U25157 ( .A(n25758), .B(n25759), .Z(n25752) );
  AND U25158 ( .A(n675), .B(n25751), .Z(n25759) );
  XNOR U25159 ( .A(n25749), .B(n25758), .Z(n25751) );
  XNOR U25160 ( .A(n25760), .B(n25761), .Z(n25749) );
  AND U25161 ( .A(n679), .B(n25762), .Z(n25761) );
  XOR U25162 ( .A(p_input[522]), .B(n25760), .Z(n25762) );
  XNOR U25163 ( .A(n25763), .B(n25764), .Z(n25760) );
  AND U25164 ( .A(n683), .B(n25765), .Z(n25764) );
  XOR U25165 ( .A(n25766), .B(n25767), .Z(n25758) );
  AND U25166 ( .A(n687), .B(n25757), .Z(n25767) );
  XNOR U25167 ( .A(n25768), .B(n25755), .Z(n25757) );
  XOR U25168 ( .A(n25769), .B(n25770), .Z(n25755) );
  AND U25169 ( .A(n710), .B(n25771), .Z(n25770) );
  IV U25170 ( .A(n25766), .Z(n25768) );
  XOR U25171 ( .A(n25772), .B(n25773), .Z(n25766) );
  AND U25172 ( .A(n694), .B(n25765), .Z(n25773) );
  XNOR U25173 ( .A(n25763), .B(n25772), .Z(n25765) );
  XNOR U25174 ( .A(n25774), .B(n25775), .Z(n25763) );
  AND U25175 ( .A(n698), .B(n25776), .Z(n25775) );
  XOR U25176 ( .A(p_input[538]), .B(n25774), .Z(n25776) );
  XNOR U25177 ( .A(n25777), .B(n25778), .Z(n25774) );
  AND U25178 ( .A(n702), .B(n25779), .Z(n25778) );
  XOR U25179 ( .A(n25780), .B(n25781), .Z(n25772) );
  AND U25180 ( .A(n706), .B(n25771), .Z(n25781) );
  XNOR U25181 ( .A(n25782), .B(n25769), .Z(n25771) );
  XOR U25182 ( .A(n25783), .B(n25784), .Z(n25769) );
  AND U25183 ( .A(n729), .B(n25785), .Z(n25784) );
  IV U25184 ( .A(n25780), .Z(n25782) );
  XOR U25185 ( .A(n25786), .B(n25787), .Z(n25780) );
  AND U25186 ( .A(n713), .B(n25779), .Z(n25787) );
  XNOR U25187 ( .A(n25777), .B(n25786), .Z(n25779) );
  XNOR U25188 ( .A(n25788), .B(n25789), .Z(n25777) );
  AND U25189 ( .A(n717), .B(n25790), .Z(n25789) );
  XOR U25190 ( .A(p_input[554]), .B(n25788), .Z(n25790) );
  XNOR U25191 ( .A(n25791), .B(n25792), .Z(n25788) );
  AND U25192 ( .A(n721), .B(n25793), .Z(n25792) );
  XOR U25193 ( .A(n25794), .B(n25795), .Z(n25786) );
  AND U25194 ( .A(n725), .B(n25785), .Z(n25795) );
  XNOR U25195 ( .A(n25796), .B(n25783), .Z(n25785) );
  XOR U25196 ( .A(n25797), .B(n25798), .Z(n25783) );
  AND U25197 ( .A(n748), .B(n25799), .Z(n25798) );
  IV U25198 ( .A(n25794), .Z(n25796) );
  XOR U25199 ( .A(n25800), .B(n25801), .Z(n25794) );
  AND U25200 ( .A(n732), .B(n25793), .Z(n25801) );
  XNOR U25201 ( .A(n25791), .B(n25800), .Z(n25793) );
  XNOR U25202 ( .A(n25802), .B(n25803), .Z(n25791) );
  AND U25203 ( .A(n736), .B(n25804), .Z(n25803) );
  XOR U25204 ( .A(p_input[570]), .B(n25802), .Z(n25804) );
  XNOR U25205 ( .A(n25805), .B(n25806), .Z(n25802) );
  AND U25206 ( .A(n740), .B(n25807), .Z(n25806) );
  XOR U25207 ( .A(n25808), .B(n25809), .Z(n25800) );
  AND U25208 ( .A(n744), .B(n25799), .Z(n25809) );
  XNOR U25209 ( .A(n25810), .B(n25797), .Z(n25799) );
  XOR U25210 ( .A(n25811), .B(n25812), .Z(n25797) );
  AND U25211 ( .A(n767), .B(n25813), .Z(n25812) );
  IV U25212 ( .A(n25808), .Z(n25810) );
  XOR U25213 ( .A(n25814), .B(n25815), .Z(n25808) );
  AND U25214 ( .A(n751), .B(n25807), .Z(n25815) );
  XNOR U25215 ( .A(n25805), .B(n25814), .Z(n25807) );
  XNOR U25216 ( .A(n25816), .B(n25817), .Z(n25805) );
  AND U25217 ( .A(n755), .B(n25818), .Z(n25817) );
  XOR U25218 ( .A(p_input[586]), .B(n25816), .Z(n25818) );
  XNOR U25219 ( .A(n25819), .B(n25820), .Z(n25816) );
  AND U25220 ( .A(n759), .B(n25821), .Z(n25820) );
  XOR U25221 ( .A(n25822), .B(n25823), .Z(n25814) );
  AND U25222 ( .A(n763), .B(n25813), .Z(n25823) );
  XNOR U25223 ( .A(n25824), .B(n25811), .Z(n25813) );
  XOR U25224 ( .A(n25825), .B(n25826), .Z(n25811) );
  AND U25225 ( .A(n786), .B(n25827), .Z(n25826) );
  IV U25226 ( .A(n25822), .Z(n25824) );
  XOR U25227 ( .A(n25828), .B(n25829), .Z(n25822) );
  AND U25228 ( .A(n770), .B(n25821), .Z(n25829) );
  XNOR U25229 ( .A(n25819), .B(n25828), .Z(n25821) );
  XNOR U25230 ( .A(n25830), .B(n25831), .Z(n25819) );
  AND U25231 ( .A(n774), .B(n25832), .Z(n25831) );
  XOR U25232 ( .A(p_input[602]), .B(n25830), .Z(n25832) );
  XNOR U25233 ( .A(n25833), .B(n25834), .Z(n25830) );
  AND U25234 ( .A(n778), .B(n25835), .Z(n25834) );
  XOR U25235 ( .A(n25836), .B(n25837), .Z(n25828) );
  AND U25236 ( .A(n782), .B(n25827), .Z(n25837) );
  XNOR U25237 ( .A(n25838), .B(n25825), .Z(n25827) );
  XOR U25238 ( .A(n25839), .B(n25840), .Z(n25825) );
  AND U25239 ( .A(n805), .B(n25841), .Z(n25840) );
  IV U25240 ( .A(n25836), .Z(n25838) );
  XOR U25241 ( .A(n25842), .B(n25843), .Z(n25836) );
  AND U25242 ( .A(n789), .B(n25835), .Z(n25843) );
  XNOR U25243 ( .A(n25833), .B(n25842), .Z(n25835) );
  XNOR U25244 ( .A(n25844), .B(n25845), .Z(n25833) );
  AND U25245 ( .A(n793), .B(n25846), .Z(n25845) );
  XOR U25246 ( .A(p_input[618]), .B(n25844), .Z(n25846) );
  XNOR U25247 ( .A(n25847), .B(n25848), .Z(n25844) );
  AND U25248 ( .A(n797), .B(n25849), .Z(n25848) );
  XOR U25249 ( .A(n25850), .B(n25851), .Z(n25842) );
  AND U25250 ( .A(n801), .B(n25841), .Z(n25851) );
  XNOR U25251 ( .A(n25852), .B(n25839), .Z(n25841) );
  XOR U25252 ( .A(n25853), .B(n25854), .Z(n25839) );
  AND U25253 ( .A(n824), .B(n25855), .Z(n25854) );
  IV U25254 ( .A(n25850), .Z(n25852) );
  XOR U25255 ( .A(n25856), .B(n25857), .Z(n25850) );
  AND U25256 ( .A(n808), .B(n25849), .Z(n25857) );
  XNOR U25257 ( .A(n25847), .B(n25856), .Z(n25849) );
  XNOR U25258 ( .A(n25858), .B(n25859), .Z(n25847) );
  AND U25259 ( .A(n812), .B(n25860), .Z(n25859) );
  XOR U25260 ( .A(p_input[634]), .B(n25858), .Z(n25860) );
  XNOR U25261 ( .A(n25861), .B(n25862), .Z(n25858) );
  AND U25262 ( .A(n816), .B(n25863), .Z(n25862) );
  XOR U25263 ( .A(n25864), .B(n25865), .Z(n25856) );
  AND U25264 ( .A(n820), .B(n25855), .Z(n25865) );
  XNOR U25265 ( .A(n25866), .B(n25853), .Z(n25855) );
  XOR U25266 ( .A(n25867), .B(n25868), .Z(n25853) );
  AND U25267 ( .A(n843), .B(n25869), .Z(n25868) );
  IV U25268 ( .A(n25864), .Z(n25866) );
  XOR U25269 ( .A(n25870), .B(n25871), .Z(n25864) );
  AND U25270 ( .A(n827), .B(n25863), .Z(n25871) );
  XNOR U25271 ( .A(n25861), .B(n25870), .Z(n25863) );
  XNOR U25272 ( .A(n25872), .B(n25873), .Z(n25861) );
  AND U25273 ( .A(n831), .B(n25874), .Z(n25873) );
  XOR U25274 ( .A(p_input[650]), .B(n25872), .Z(n25874) );
  XNOR U25275 ( .A(n25875), .B(n25876), .Z(n25872) );
  AND U25276 ( .A(n835), .B(n25877), .Z(n25876) );
  XOR U25277 ( .A(n25878), .B(n25879), .Z(n25870) );
  AND U25278 ( .A(n839), .B(n25869), .Z(n25879) );
  XNOR U25279 ( .A(n25880), .B(n25867), .Z(n25869) );
  XOR U25280 ( .A(n25881), .B(n25882), .Z(n25867) );
  AND U25281 ( .A(n862), .B(n25883), .Z(n25882) );
  IV U25282 ( .A(n25878), .Z(n25880) );
  XOR U25283 ( .A(n25884), .B(n25885), .Z(n25878) );
  AND U25284 ( .A(n846), .B(n25877), .Z(n25885) );
  XNOR U25285 ( .A(n25875), .B(n25884), .Z(n25877) );
  XNOR U25286 ( .A(n25886), .B(n25887), .Z(n25875) );
  AND U25287 ( .A(n850), .B(n25888), .Z(n25887) );
  XOR U25288 ( .A(p_input[666]), .B(n25886), .Z(n25888) );
  XNOR U25289 ( .A(n25889), .B(n25890), .Z(n25886) );
  AND U25290 ( .A(n854), .B(n25891), .Z(n25890) );
  XOR U25291 ( .A(n25892), .B(n25893), .Z(n25884) );
  AND U25292 ( .A(n858), .B(n25883), .Z(n25893) );
  XNOR U25293 ( .A(n25894), .B(n25881), .Z(n25883) );
  XOR U25294 ( .A(n25895), .B(n25896), .Z(n25881) );
  AND U25295 ( .A(n881), .B(n25897), .Z(n25896) );
  IV U25296 ( .A(n25892), .Z(n25894) );
  XOR U25297 ( .A(n25898), .B(n25899), .Z(n25892) );
  AND U25298 ( .A(n865), .B(n25891), .Z(n25899) );
  XNOR U25299 ( .A(n25889), .B(n25898), .Z(n25891) );
  XNOR U25300 ( .A(n25900), .B(n25901), .Z(n25889) );
  AND U25301 ( .A(n869), .B(n25902), .Z(n25901) );
  XOR U25302 ( .A(p_input[682]), .B(n25900), .Z(n25902) );
  XNOR U25303 ( .A(n25903), .B(n25904), .Z(n25900) );
  AND U25304 ( .A(n873), .B(n25905), .Z(n25904) );
  XOR U25305 ( .A(n25906), .B(n25907), .Z(n25898) );
  AND U25306 ( .A(n877), .B(n25897), .Z(n25907) );
  XNOR U25307 ( .A(n25908), .B(n25895), .Z(n25897) );
  XOR U25308 ( .A(n25909), .B(n25910), .Z(n25895) );
  AND U25309 ( .A(n900), .B(n25911), .Z(n25910) );
  IV U25310 ( .A(n25906), .Z(n25908) );
  XOR U25311 ( .A(n25912), .B(n25913), .Z(n25906) );
  AND U25312 ( .A(n884), .B(n25905), .Z(n25913) );
  XNOR U25313 ( .A(n25903), .B(n25912), .Z(n25905) );
  XNOR U25314 ( .A(n25914), .B(n25915), .Z(n25903) );
  AND U25315 ( .A(n888), .B(n25916), .Z(n25915) );
  XOR U25316 ( .A(p_input[698]), .B(n25914), .Z(n25916) );
  XNOR U25317 ( .A(n25917), .B(n25918), .Z(n25914) );
  AND U25318 ( .A(n892), .B(n25919), .Z(n25918) );
  XOR U25319 ( .A(n25920), .B(n25921), .Z(n25912) );
  AND U25320 ( .A(n896), .B(n25911), .Z(n25921) );
  XNOR U25321 ( .A(n25922), .B(n25909), .Z(n25911) );
  XOR U25322 ( .A(n25923), .B(n25924), .Z(n25909) );
  AND U25323 ( .A(n919), .B(n25925), .Z(n25924) );
  IV U25324 ( .A(n25920), .Z(n25922) );
  XOR U25325 ( .A(n25926), .B(n25927), .Z(n25920) );
  AND U25326 ( .A(n903), .B(n25919), .Z(n25927) );
  XNOR U25327 ( .A(n25917), .B(n25926), .Z(n25919) );
  XNOR U25328 ( .A(n25928), .B(n25929), .Z(n25917) );
  AND U25329 ( .A(n907), .B(n25930), .Z(n25929) );
  XOR U25330 ( .A(p_input[714]), .B(n25928), .Z(n25930) );
  XNOR U25331 ( .A(n25931), .B(n25932), .Z(n25928) );
  AND U25332 ( .A(n911), .B(n25933), .Z(n25932) );
  XOR U25333 ( .A(n25934), .B(n25935), .Z(n25926) );
  AND U25334 ( .A(n915), .B(n25925), .Z(n25935) );
  XNOR U25335 ( .A(n25936), .B(n25923), .Z(n25925) );
  XOR U25336 ( .A(n25937), .B(n25938), .Z(n25923) );
  AND U25337 ( .A(n938), .B(n25939), .Z(n25938) );
  IV U25338 ( .A(n25934), .Z(n25936) );
  XOR U25339 ( .A(n25940), .B(n25941), .Z(n25934) );
  AND U25340 ( .A(n922), .B(n25933), .Z(n25941) );
  XNOR U25341 ( .A(n25931), .B(n25940), .Z(n25933) );
  XNOR U25342 ( .A(n25942), .B(n25943), .Z(n25931) );
  AND U25343 ( .A(n926), .B(n25944), .Z(n25943) );
  XOR U25344 ( .A(p_input[730]), .B(n25942), .Z(n25944) );
  XNOR U25345 ( .A(n25945), .B(n25946), .Z(n25942) );
  AND U25346 ( .A(n930), .B(n25947), .Z(n25946) );
  XOR U25347 ( .A(n25948), .B(n25949), .Z(n25940) );
  AND U25348 ( .A(n934), .B(n25939), .Z(n25949) );
  XNOR U25349 ( .A(n25950), .B(n25937), .Z(n25939) );
  XOR U25350 ( .A(n25951), .B(n25952), .Z(n25937) );
  AND U25351 ( .A(n957), .B(n25953), .Z(n25952) );
  IV U25352 ( .A(n25948), .Z(n25950) );
  XOR U25353 ( .A(n25954), .B(n25955), .Z(n25948) );
  AND U25354 ( .A(n941), .B(n25947), .Z(n25955) );
  XNOR U25355 ( .A(n25945), .B(n25954), .Z(n25947) );
  XNOR U25356 ( .A(n25956), .B(n25957), .Z(n25945) );
  AND U25357 ( .A(n945), .B(n25958), .Z(n25957) );
  XOR U25358 ( .A(p_input[746]), .B(n25956), .Z(n25958) );
  XNOR U25359 ( .A(n25959), .B(n25960), .Z(n25956) );
  AND U25360 ( .A(n949), .B(n25961), .Z(n25960) );
  XOR U25361 ( .A(n25962), .B(n25963), .Z(n25954) );
  AND U25362 ( .A(n953), .B(n25953), .Z(n25963) );
  XNOR U25363 ( .A(n25964), .B(n25951), .Z(n25953) );
  XOR U25364 ( .A(n25965), .B(n25966), .Z(n25951) );
  AND U25365 ( .A(n976), .B(n25967), .Z(n25966) );
  IV U25366 ( .A(n25962), .Z(n25964) );
  XOR U25367 ( .A(n25968), .B(n25969), .Z(n25962) );
  AND U25368 ( .A(n960), .B(n25961), .Z(n25969) );
  XNOR U25369 ( .A(n25959), .B(n25968), .Z(n25961) );
  XNOR U25370 ( .A(n25970), .B(n25971), .Z(n25959) );
  AND U25371 ( .A(n964), .B(n25972), .Z(n25971) );
  XOR U25372 ( .A(p_input[762]), .B(n25970), .Z(n25972) );
  XNOR U25373 ( .A(n25973), .B(n25974), .Z(n25970) );
  AND U25374 ( .A(n968), .B(n25975), .Z(n25974) );
  XOR U25375 ( .A(n25976), .B(n25977), .Z(n25968) );
  AND U25376 ( .A(n972), .B(n25967), .Z(n25977) );
  XNOR U25377 ( .A(n25978), .B(n25965), .Z(n25967) );
  XOR U25378 ( .A(n25979), .B(n25980), .Z(n25965) );
  AND U25379 ( .A(n995), .B(n25981), .Z(n25980) );
  IV U25380 ( .A(n25976), .Z(n25978) );
  XOR U25381 ( .A(n25982), .B(n25983), .Z(n25976) );
  AND U25382 ( .A(n979), .B(n25975), .Z(n25983) );
  XNOR U25383 ( .A(n25973), .B(n25982), .Z(n25975) );
  XNOR U25384 ( .A(n25984), .B(n25985), .Z(n25973) );
  AND U25385 ( .A(n983), .B(n25986), .Z(n25985) );
  XOR U25386 ( .A(p_input[778]), .B(n25984), .Z(n25986) );
  XNOR U25387 ( .A(n25987), .B(n25988), .Z(n25984) );
  AND U25388 ( .A(n987), .B(n25989), .Z(n25988) );
  XOR U25389 ( .A(n25990), .B(n25991), .Z(n25982) );
  AND U25390 ( .A(n991), .B(n25981), .Z(n25991) );
  XNOR U25391 ( .A(n25992), .B(n25979), .Z(n25981) );
  XOR U25392 ( .A(n25993), .B(n25994), .Z(n25979) );
  AND U25393 ( .A(n1014), .B(n25995), .Z(n25994) );
  IV U25394 ( .A(n25990), .Z(n25992) );
  XOR U25395 ( .A(n25996), .B(n25997), .Z(n25990) );
  AND U25396 ( .A(n998), .B(n25989), .Z(n25997) );
  XNOR U25397 ( .A(n25987), .B(n25996), .Z(n25989) );
  XNOR U25398 ( .A(n25998), .B(n25999), .Z(n25987) );
  AND U25399 ( .A(n1002), .B(n26000), .Z(n25999) );
  XOR U25400 ( .A(p_input[794]), .B(n25998), .Z(n26000) );
  XNOR U25401 ( .A(n26001), .B(n26002), .Z(n25998) );
  AND U25402 ( .A(n1006), .B(n26003), .Z(n26002) );
  XOR U25403 ( .A(n26004), .B(n26005), .Z(n25996) );
  AND U25404 ( .A(n1010), .B(n25995), .Z(n26005) );
  XNOR U25405 ( .A(n26006), .B(n25993), .Z(n25995) );
  XOR U25406 ( .A(n26007), .B(n26008), .Z(n25993) );
  AND U25407 ( .A(n1033), .B(n26009), .Z(n26008) );
  IV U25408 ( .A(n26004), .Z(n26006) );
  XOR U25409 ( .A(n26010), .B(n26011), .Z(n26004) );
  AND U25410 ( .A(n1017), .B(n26003), .Z(n26011) );
  XNOR U25411 ( .A(n26001), .B(n26010), .Z(n26003) );
  XNOR U25412 ( .A(n26012), .B(n26013), .Z(n26001) );
  AND U25413 ( .A(n1021), .B(n26014), .Z(n26013) );
  XOR U25414 ( .A(p_input[810]), .B(n26012), .Z(n26014) );
  XNOR U25415 ( .A(n26015), .B(n26016), .Z(n26012) );
  AND U25416 ( .A(n1025), .B(n26017), .Z(n26016) );
  XOR U25417 ( .A(n26018), .B(n26019), .Z(n26010) );
  AND U25418 ( .A(n1029), .B(n26009), .Z(n26019) );
  XNOR U25419 ( .A(n26020), .B(n26007), .Z(n26009) );
  XOR U25420 ( .A(n26021), .B(n26022), .Z(n26007) );
  AND U25421 ( .A(n1052), .B(n26023), .Z(n26022) );
  IV U25422 ( .A(n26018), .Z(n26020) );
  XOR U25423 ( .A(n26024), .B(n26025), .Z(n26018) );
  AND U25424 ( .A(n1036), .B(n26017), .Z(n26025) );
  XNOR U25425 ( .A(n26015), .B(n26024), .Z(n26017) );
  XNOR U25426 ( .A(n26026), .B(n26027), .Z(n26015) );
  AND U25427 ( .A(n1040), .B(n26028), .Z(n26027) );
  XOR U25428 ( .A(p_input[826]), .B(n26026), .Z(n26028) );
  XNOR U25429 ( .A(n26029), .B(n26030), .Z(n26026) );
  AND U25430 ( .A(n1044), .B(n26031), .Z(n26030) );
  XOR U25431 ( .A(n26032), .B(n26033), .Z(n26024) );
  AND U25432 ( .A(n1048), .B(n26023), .Z(n26033) );
  XNOR U25433 ( .A(n26034), .B(n26021), .Z(n26023) );
  XOR U25434 ( .A(n26035), .B(n26036), .Z(n26021) );
  AND U25435 ( .A(n1071), .B(n26037), .Z(n26036) );
  IV U25436 ( .A(n26032), .Z(n26034) );
  XOR U25437 ( .A(n26038), .B(n26039), .Z(n26032) );
  AND U25438 ( .A(n1055), .B(n26031), .Z(n26039) );
  XNOR U25439 ( .A(n26029), .B(n26038), .Z(n26031) );
  XNOR U25440 ( .A(n26040), .B(n26041), .Z(n26029) );
  AND U25441 ( .A(n1059), .B(n26042), .Z(n26041) );
  XOR U25442 ( .A(p_input[842]), .B(n26040), .Z(n26042) );
  XNOR U25443 ( .A(n26043), .B(n26044), .Z(n26040) );
  AND U25444 ( .A(n1063), .B(n26045), .Z(n26044) );
  XOR U25445 ( .A(n26046), .B(n26047), .Z(n26038) );
  AND U25446 ( .A(n1067), .B(n26037), .Z(n26047) );
  XNOR U25447 ( .A(n26048), .B(n26035), .Z(n26037) );
  XOR U25448 ( .A(n26049), .B(n26050), .Z(n26035) );
  AND U25449 ( .A(n1090), .B(n26051), .Z(n26050) );
  IV U25450 ( .A(n26046), .Z(n26048) );
  XOR U25451 ( .A(n26052), .B(n26053), .Z(n26046) );
  AND U25452 ( .A(n1074), .B(n26045), .Z(n26053) );
  XNOR U25453 ( .A(n26043), .B(n26052), .Z(n26045) );
  XNOR U25454 ( .A(n26054), .B(n26055), .Z(n26043) );
  AND U25455 ( .A(n1078), .B(n26056), .Z(n26055) );
  XOR U25456 ( .A(p_input[858]), .B(n26054), .Z(n26056) );
  XNOR U25457 ( .A(n26057), .B(n26058), .Z(n26054) );
  AND U25458 ( .A(n1082), .B(n26059), .Z(n26058) );
  XOR U25459 ( .A(n26060), .B(n26061), .Z(n26052) );
  AND U25460 ( .A(n1086), .B(n26051), .Z(n26061) );
  XNOR U25461 ( .A(n26062), .B(n26049), .Z(n26051) );
  XOR U25462 ( .A(n26063), .B(n26064), .Z(n26049) );
  AND U25463 ( .A(n1109), .B(n26065), .Z(n26064) );
  IV U25464 ( .A(n26060), .Z(n26062) );
  XOR U25465 ( .A(n26066), .B(n26067), .Z(n26060) );
  AND U25466 ( .A(n1093), .B(n26059), .Z(n26067) );
  XNOR U25467 ( .A(n26057), .B(n26066), .Z(n26059) );
  XNOR U25468 ( .A(n26068), .B(n26069), .Z(n26057) );
  AND U25469 ( .A(n1097), .B(n26070), .Z(n26069) );
  XOR U25470 ( .A(p_input[874]), .B(n26068), .Z(n26070) );
  XNOR U25471 ( .A(n26071), .B(n26072), .Z(n26068) );
  AND U25472 ( .A(n1101), .B(n26073), .Z(n26072) );
  XOR U25473 ( .A(n26074), .B(n26075), .Z(n26066) );
  AND U25474 ( .A(n1105), .B(n26065), .Z(n26075) );
  XNOR U25475 ( .A(n26076), .B(n26063), .Z(n26065) );
  XOR U25476 ( .A(n26077), .B(n26078), .Z(n26063) );
  AND U25477 ( .A(n1128), .B(n26079), .Z(n26078) );
  IV U25478 ( .A(n26074), .Z(n26076) );
  XOR U25479 ( .A(n26080), .B(n26081), .Z(n26074) );
  AND U25480 ( .A(n1112), .B(n26073), .Z(n26081) );
  XNOR U25481 ( .A(n26071), .B(n26080), .Z(n26073) );
  XNOR U25482 ( .A(n26082), .B(n26083), .Z(n26071) );
  AND U25483 ( .A(n1116), .B(n26084), .Z(n26083) );
  XOR U25484 ( .A(p_input[890]), .B(n26082), .Z(n26084) );
  XNOR U25485 ( .A(n26085), .B(n26086), .Z(n26082) );
  AND U25486 ( .A(n1120), .B(n26087), .Z(n26086) );
  XOR U25487 ( .A(n26088), .B(n26089), .Z(n26080) );
  AND U25488 ( .A(n1124), .B(n26079), .Z(n26089) );
  XNOR U25489 ( .A(n26090), .B(n26077), .Z(n26079) );
  XOR U25490 ( .A(n26091), .B(n26092), .Z(n26077) );
  AND U25491 ( .A(n1147), .B(n26093), .Z(n26092) );
  IV U25492 ( .A(n26088), .Z(n26090) );
  XOR U25493 ( .A(n26094), .B(n26095), .Z(n26088) );
  AND U25494 ( .A(n1131), .B(n26087), .Z(n26095) );
  XNOR U25495 ( .A(n26085), .B(n26094), .Z(n26087) );
  XNOR U25496 ( .A(n26096), .B(n26097), .Z(n26085) );
  AND U25497 ( .A(n1135), .B(n26098), .Z(n26097) );
  XOR U25498 ( .A(p_input[906]), .B(n26096), .Z(n26098) );
  XNOR U25499 ( .A(n26099), .B(n26100), .Z(n26096) );
  AND U25500 ( .A(n1139), .B(n26101), .Z(n26100) );
  XOR U25501 ( .A(n26102), .B(n26103), .Z(n26094) );
  AND U25502 ( .A(n1143), .B(n26093), .Z(n26103) );
  XNOR U25503 ( .A(n26104), .B(n26091), .Z(n26093) );
  XOR U25504 ( .A(n26105), .B(n26106), .Z(n26091) );
  AND U25505 ( .A(n1166), .B(n26107), .Z(n26106) );
  IV U25506 ( .A(n26102), .Z(n26104) );
  XOR U25507 ( .A(n26108), .B(n26109), .Z(n26102) );
  AND U25508 ( .A(n1150), .B(n26101), .Z(n26109) );
  XNOR U25509 ( .A(n26099), .B(n26108), .Z(n26101) );
  XNOR U25510 ( .A(n26110), .B(n26111), .Z(n26099) );
  AND U25511 ( .A(n1154), .B(n26112), .Z(n26111) );
  XOR U25512 ( .A(p_input[922]), .B(n26110), .Z(n26112) );
  XNOR U25513 ( .A(n26113), .B(n26114), .Z(n26110) );
  AND U25514 ( .A(n1158), .B(n26115), .Z(n26114) );
  XOR U25515 ( .A(n26116), .B(n26117), .Z(n26108) );
  AND U25516 ( .A(n1162), .B(n26107), .Z(n26117) );
  XNOR U25517 ( .A(n26118), .B(n26105), .Z(n26107) );
  XOR U25518 ( .A(n26119), .B(n26120), .Z(n26105) );
  AND U25519 ( .A(n1185), .B(n26121), .Z(n26120) );
  IV U25520 ( .A(n26116), .Z(n26118) );
  XOR U25521 ( .A(n26122), .B(n26123), .Z(n26116) );
  AND U25522 ( .A(n1169), .B(n26115), .Z(n26123) );
  XNOR U25523 ( .A(n26113), .B(n26122), .Z(n26115) );
  XNOR U25524 ( .A(n26124), .B(n26125), .Z(n26113) );
  AND U25525 ( .A(n1173), .B(n26126), .Z(n26125) );
  XOR U25526 ( .A(p_input[938]), .B(n26124), .Z(n26126) );
  XNOR U25527 ( .A(n26127), .B(n26128), .Z(n26124) );
  AND U25528 ( .A(n1177), .B(n26129), .Z(n26128) );
  XOR U25529 ( .A(n26130), .B(n26131), .Z(n26122) );
  AND U25530 ( .A(n1181), .B(n26121), .Z(n26131) );
  XNOR U25531 ( .A(n26132), .B(n26119), .Z(n26121) );
  XOR U25532 ( .A(n26133), .B(n26134), .Z(n26119) );
  AND U25533 ( .A(n1204), .B(n26135), .Z(n26134) );
  IV U25534 ( .A(n26130), .Z(n26132) );
  XOR U25535 ( .A(n26136), .B(n26137), .Z(n26130) );
  AND U25536 ( .A(n1188), .B(n26129), .Z(n26137) );
  XNOR U25537 ( .A(n26127), .B(n26136), .Z(n26129) );
  XNOR U25538 ( .A(n26138), .B(n26139), .Z(n26127) );
  AND U25539 ( .A(n1192), .B(n26140), .Z(n26139) );
  XOR U25540 ( .A(p_input[954]), .B(n26138), .Z(n26140) );
  XNOR U25541 ( .A(n26141), .B(n26142), .Z(n26138) );
  AND U25542 ( .A(n1196), .B(n26143), .Z(n26142) );
  XOR U25543 ( .A(n26144), .B(n26145), .Z(n26136) );
  AND U25544 ( .A(n1200), .B(n26135), .Z(n26145) );
  XNOR U25545 ( .A(n26146), .B(n26133), .Z(n26135) );
  XOR U25546 ( .A(n26147), .B(n26148), .Z(n26133) );
  AND U25547 ( .A(n1223), .B(n26149), .Z(n26148) );
  IV U25548 ( .A(n26144), .Z(n26146) );
  XOR U25549 ( .A(n26150), .B(n26151), .Z(n26144) );
  AND U25550 ( .A(n1207), .B(n26143), .Z(n26151) );
  XNOR U25551 ( .A(n26141), .B(n26150), .Z(n26143) );
  XNOR U25552 ( .A(n26152), .B(n26153), .Z(n26141) );
  AND U25553 ( .A(n1211), .B(n26154), .Z(n26153) );
  XOR U25554 ( .A(p_input[970]), .B(n26152), .Z(n26154) );
  XNOR U25555 ( .A(n26155), .B(n26156), .Z(n26152) );
  AND U25556 ( .A(n1215), .B(n26157), .Z(n26156) );
  XOR U25557 ( .A(n26158), .B(n26159), .Z(n26150) );
  AND U25558 ( .A(n1219), .B(n26149), .Z(n26159) );
  XNOR U25559 ( .A(n26160), .B(n26147), .Z(n26149) );
  XOR U25560 ( .A(n26161), .B(n26162), .Z(n26147) );
  AND U25561 ( .A(n1242), .B(n26163), .Z(n26162) );
  IV U25562 ( .A(n26158), .Z(n26160) );
  XOR U25563 ( .A(n26164), .B(n26165), .Z(n26158) );
  AND U25564 ( .A(n1226), .B(n26157), .Z(n26165) );
  XNOR U25565 ( .A(n26155), .B(n26164), .Z(n26157) );
  XNOR U25566 ( .A(n26166), .B(n26167), .Z(n26155) );
  AND U25567 ( .A(n1230), .B(n26168), .Z(n26167) );
  XOR U25568 ( .A(p_input[986]), .B(n26166), .Z(n26168) );
  XNOR U25569 ( .A(n26169), .B(n26170), .Z(n26166) );
  AND U25570 ( .A(n1234), .B(n26171), .Z(n26170) );
  XOR U25571 ( .A(n26172), .B(n26173), .Z(n26164) );
  AND U25572 ( .A(n1238), .B(n26163), .Z(n26173) );
  XNOR U25573 ( .A(n26174), .B(n26161), .Z(n26163) );
  XOR U25574 ( .A(n26175), .B(n26176), .Z(n26161) );
  AND U25575 ( .A(n1261), .B(n26177), .Z(n26176) );
  IV U25576 ( .A(n26172), .Z(n26174) );
  XOR U25577 ( .A(n26178), .B(n26179), .Z(n26172) );
  AND U25578 ( .A(n1245), .B(n26171), .Z(n26179) );
  XNOR U25579 ( .A(n26169), .B(n26178), .Z(n26171) );
  XNOR U25580 ( .A(n26180), .B(n26181), .Z(n26169) );
  AND U25581 ( .A(n1249), .B(n26182), .Z(n26181) );
  XOR U25582 ( .A(p_input[1002]), .B(n26180), .Z(n26182) );
  XNOR U25583 ( .A(n26183), .B(n26184), .Z(n26180) );
  AND U25584 ( .A(n1253), .B(n26185), .Z(n26184) );
  XOR U25585 ( .A(n26186), .B(n26187), .Z(n26178) );
  AND U25586 ( .A(n1257), .B(n26177), .Z(n26187) );
  XNOR U25587 ( .A(n26188), .B(n26175), .Z(n26177) );
  XOR U25588 ( .A(n26189), .B(n26190), .Z(n26175) );
  AND U25589 ( .A(n1280), .B(n26191), .Z(n26190) );
  IV U25590 ( .A(n26186), .Z(n26188) );
  XOR U25591 ( .A(n26192), .B(n26193), .Z(n26186) );
  AND U25592 ( .A(n1264), .B(n26185), .Z(n26193) );
  XNOR U25593 ( .A(n26183), .B(n26192), .Z(n26185) );
  XNOR U25594 ( .A(n26194), .B(n26195), .Z(n26183) );
  AND U25595 ( .A(n1268), .B(n26196), .Z(n26195) );
  XOR U25596 ( .A(p_input[1018]), .B(n26194), .Z(n26196) );
  XNOR U25597 ( .A(n26197), .B(n26198), .Z(n26194) );
  AND U25598 ( .A(n1272), .B(n26199), .Z(n26198) );
  XOR U25599 ( .A(n26200), .B(n26201), .Z(n26192) );
  AND U25600 ( .A(n1276), .B(n26191), .Z(n26201) );
  XNOR U25601 ( .A(n26202), .B(n26189), .Z(n26191) );
  XOR U25602 ( .A(n26203), .B(n26204), .Z(n26189) );
  AND U25603 ( .A(n1299), .B(n26205), .Z(n26204) );
  IV U25604 ( .A(n26200), .Z(n26202) );
  XOR U25605 ( .A(n26206), .B(n26207), .Z(n26200) );
  AND U25606 ( .A(n1283), .B(n26199), .Z(n26207) );
  XNOR U25607 ( .A(n26197), .B(n26206), .Z(n26199) );
  XNOR U25608 ( .A(n26208), .B(n26209), .Z(n26197) );
  AND U25609 ( .A(n1287), .B(n26210), .Z(n26209) );
  XOR U25610 ( .A(p_input[1034]), .B(n26208), .Z(n26210) );
  XNOR U25611 ( .A(n26211), .B(n26212), .Z(n26208) );
  AND U25612 ( .A(n1291), .B(n26213), .Z(n26212) );
  XOR U25613 ( .A(n26214), .B(n26215), .Z(n26206) );
  AND U25614 ( .A(n1295), .B(n26205), .Z(n26215) );
  XNOR U25615 ( .A(n26216), .B(n26203), .Z(n26205) );
  XOR U25616 ( .A(n26217), .B(n26218), .Z(n26203) );
  AND U25617 ( .A(n1318), .B(n26219), .Z(n26218) );
  IV U25618 ( .A(n26214), .Z(n26216) );
  XOR U25619 ( .A(n26220), .B(n26221), .Z(n26214) );
  AND U25620 ( .A(n1302), .B(n26213), .Z(n26221) );
  XNOR U25621 ( .A(n26211), .B(n26220), .Z(n26213) );
  XNOR U25622 ( .A(n26222), .B(n26223), .Z(n26211) );
  AND U25623 ( .A(n1306), .B(n26224), .Z(n26223) );
  XOR U25624 ( .A(p_input[1050]), .B(n26222), .Z(n26224) );
  XNOR U25625 ( .A(n26225), .B(n26226), .Z(n26222) );
  AND U25626 ( .A(n1310), .B(n26227), .Z(n26226) );
  XOR U25627 ( .A(n26228), .B(n26229), .Z(n26220) );
  AND U25628 ( .A(n1314), .B(n26219), .Z(n26229) );
  XNOR U25629 ( .A(n26230), .B(n26217), .Z(n26219) );
  XOR U25630 ( .A(n26231), .B(n26232), .Z(n26217) );
  AND U25631 ( .A(n1337), .B(n26233), .Z(n26232) );
  IV U25632 ( .A(n26228), .Z(n26230) );
  XOR U25633 ( .A(n26234), .B(n26235), .Z(n26228) );
  AND U25634 ( .A(n1321), .B(n26227), .Z(n26235) );
  XNOR U25635 ( .A(n26225), .B(n26234), .Z(n26227) );
  XNOR U25636 ( .A(n26236), .B(n26237), .Z(n26225) );
  AND U25637 ( .A(n1325), .B(n26238), .Z(n26237) );
  XOR U25638 ( .A(p_input[1066]), .B(n26236), .Z(n26238) );
  XNOR U25639 ( .A(n26239), .B(n26240), .Z(n26236) );
  AND U25640 ( .A(n1329), .B(n26241), .Z(n26240) );
  XOR U25641 ( .A(n26242), .B(n26243), .Z(n26234) );
  AND U25642 ( .A(n1333), .B(n26233), .Z(n26243) );
  XNOR U25643 ( .A(n26244), .B(n26231), .Z(n26233) );
  XOR U25644 ( .A(n26245), .B(n26246), .Z(n26231) );
  AND U25645 ( .A(n1356), .B(n26247), .Z(n26246) );
  IV U25646 ( .A(n26242), .Z(n26244) );
  XOR U25647 ( .A(n26248), .B(n26249), .Z(n26242) );
  AND U25648 ( .A(n1340), .B(n26241), .Z(n26249) );
  XNOR U25649 ( .A(n26239), .B(n26248), .Z(n26241) );
  XNOR U25650 ( .A(n26250), .B(n26251), .Z(n26239) );
  AND U25651 ( .A(n1344), .B(n26252), .Z(n26251) );
  XOR U25652 ( .A(p_input[1082]), .B(n26250), .Z(n26252) );
  XNOR U25653 ( .A(n26253), .B(n26254), .Z(n26250) );
  AND U25654 ( .A(n1348), .B(n26255), .Z(n26254) );
  XOR U25655 ( .A(n26256), .B(n26257), .Z(n26248) );
  AND U25656 ( .A(n1352), .B(n26247), .Z(n26257) );
  XNOR U25657 ( .A(n26258), .B(n26245), .Z(n26247) );
  XOR U25658 ( .A(n26259), .B(n26260), .Z(n26245) );
  AND U25659 ( .A(n1375), .B(n26261), .Z(n26260) );
  IV U25660 ( .A(n26256), .Z(n26258) );
  XOR U25661 ( .A(n26262), .B(n26263), .Z(n26256) );
  AND U25662 ( .A(n1359), .B(n26255), .Z(n26263) );
  XNOR U25663 ( .A(n26253), .B(n26262), .Z(n26255) );
  XNOR U25664 ( .A(n26264), .B(n26265), .Z(n26253) );
  AND U25665 ( .A(n1363), .B(n26266), .Z(n26265) );
  XOR U25666 ( .A(p_input[1098]), .B(n26264), .Z(n26266) );
  XNOR U25667 ( .A(n26267), .B(n26268), .Z(n26264) );
  AND U25668 ( .A(n1367), .B(n26269), .Z(n26268) );
  XOR U25669 ( .A(n26270), .B(n26271), .Z(n26262) );
  AND U25670 ( .A(n1371), .B(n26261), .Z(n26271) );
  XNOR U25671 ( .A(n26272), .B(n26259), .Z(n26261) );
  XOR U25672 ( .A(n26273), .B(n26274), .Z(n26259) );
  AND U25673 ( .A(n1394), .B(n26275), .Z(n26274) );
  IV U25674 ( .A(n26270), .Z(n26272) );
  XOR U25675 ( .A(n26276), .B(n26277), .Z(n26270) );
  AND U25676 ( .A(n1378), .B(n26269), .Z(n26277) );
  XNOR U25677 ( .A(n26267), .B(n26276), .Z(n26269) );
  XNOR U25678 ( .A(n26278), .B(n26279), .Z(n26267) );
  AND U25679 ( .A(n1382), .B(n26280), .Z(n26279) );
  XOR U25680 ( .A(p_input[1114]), .B(n26278), .Z(n26280) );
  XNOR U25681 ( .A(n26281), .B(n26282), .Z(n26278) );
  AND U25682 ( .A(n1386), .B(n26283), .Z(n26282) );
  XOR U25683 ( .A(n26284), .B(n26285), .Z(n26276) );
  AND U25684 ( .A(n1390), .B(n26275), .Z(n26285) );
  XNOR U25685 ( .A(n26286), .B(n26273), .Z(n26275) );
  XOR U25686 ( .A(n26287), .B(n26288), .Z(n26273) );
  AND U25687 ( .A(n1413), .B(n26289), .Z(n26288) );
  IV U25688 ( .A(n26284), .Z(n26286) );
  XOR U25689 ( .A(n26290), .B(n26291), .Z(n26284) );
  AND U25690 ( .A(n1397), .B(n26283), .Z(n26291) );
  XNOR U25691 ( .A(n26281), .B(n26290), .Z(n26283) );
  XNOR U25692 ( .A(n26292), .B(n26293), .Z(n26281) );
  AND U25693 ( .A(n1401), .B(n26294), .Z(n26293) );
  XOR U25694 ( .A(p_input[1130]), .B(n26292), .Z(n26294) );
  XNOR U25695 ( .A(n26295), .B(n26296), .Z(n26292) );
  AND U25696 ( .A(n1405), .B(n26297), .Z(n26296) );
  XOR U25697 ( .A(n26298), .B(n26299), .Z(n26290) );
  AND U25698 ( .A(n1409), .B(n26289), .Z(n26299) );
  XNOR U25699 ( .A(n26300), .B(n26287), .Z(n26289) );
  XOR U25700 ( .A(n26301), .B(n26302), .Z(n26287) );
  AND U25701 ( .A(n1432), .B(n26303), .Z(n26302) );
  IV U25702 ( .A(n26298), .Z(n26300) );
  XOR U25703 ( .A(n26304), .B(n26305), .Z(n26298) );
  AND U25704 ( .A(n1416), .B(n26297), .Z(n26305) );
  XNOR U25705 ( .A(n26295), .B(n26304), .Z(n26297) );
  XNOR U25706 ( .A(n26306), .B(n26307), .Z(n26295) );
  AND U25707 ( .A(n1420), .B(n26308), .Z(n26307) );
  XOR U25708 ( .A(p_input[1146]), .B(n26306), .Z(n26308) );
  XNOR U25709 ( .A(n26309), .B(n26310), .Z(n26306) );
  AND U25710 ( .A(n1424), .B(n26311), .Z(n26310) );
  XOR U25711 ( .A(n26312), .B(n26313), .Z(n26304) );
  AND U25712 ( .A(n1428), .B(n26303), .Z(n26313) );
  XNOR U25713 ( .A(n26314), .B(n26301), .Z(n26303) );
  XOR U25714 ( .A(n26315), .B(n26316), .Z(n26301) );
  AND U25715 ( .A(n1451), .B(n26317), .Z(n26316) );
  IV U25716 ( .A(n26312), .Z(n26314) );
  XOR U25717 ( .A(n26318), .B(n26319), .Z(n26312) );
  AND U25718 ( .A(n1435), .B(n26311), .Z(n26319) );
  XNOR U25719 ( .A(n26309), .B(n26318), .Z(n26311) );
  XNOR U25720 ( .A(n26320), .B(n26321), .Z(n26309) );
  AND U25721 ( .A(n1439), .B(n26322), .Z(n26321) );
  XOR U25722 ( .A(p_input[1162]), .B(n26320), .Z(n26322) );
  XNOR U25723 ( .A(n26323), .B(n26324), .Z(n26320) );
  AND U25724 ( .A(n1443), .B(n26325), .Z(n26324) );
  XOR U25725 ( .A(n26326), .B(n26327), .Z(n26318) );
  AND U25726 ( .A(n1447), .B(n26317), .Z(n26327) );
  XNOR U25727 ( .A(n26328), .B(n26315), .Z(n26317) );
  XOR U25728 ( .A(n26329), .B(n26330), .Z(n26315) );
  AND U25729 ( .A(n1470), .B(n26331), .Z(n26330) );
  IV U25730 ( .A(n26326), .Z(n26328) );
  XOR U25731 ( .A(n26332), .B(n26333), .Z(n26326) );
  AND U25732 ( .A(n1454), .B(n26325), .Z(n26333) );
  XNOR U25733 ( .A(n26323), .B(n26332), .Z(n26325) );
  XNOR U25734 ( .A(n26334), .B(n26335), .Z(n26323) );
  AND U25735 ( .A(n1458), .B(n26336), .Z(n26335) );
  XOR U25736 ( .A(p_input[1178]), .B(n26334), .Z(n26336) );
  XNOR U25737 ( .A(n26337), .B(n26338), .Z(n26334) );
  AND U25738 ( .A(n1462), .B(n26339), .Z(n26338) );
  XOR U25739 ( .A(n26340), .B(n26341), .Z(n26332) );
  AND U25740 ( .A(n1466), .B(n26331), .Z(n26341) );
  XNOR U25741 ( .A(n26342), .B(n26329), .Z(n26331) );
  XOR U25742 ( .A(n26343), .B(n26344), .Z(n26329) );
  AND U25743 ( .A(n1489), .B(n26345), .Z(n26344) );
  IV U25744 ( .A(n26340), .Z(n26342) );
  XOR U25745 ( .A(n26346), .B(n26347), .Z(n26340) );
  AND U25746 ( .A(n1473), .B(n26339), .Z(n26347) );
  XNOR U25747 ( .A(n26337), .B(n26346), .Z(n26339) );
  XNOR U25748 ( .A(n26348), .B(n26349), .Z(n26337) );
  AND U25749 ( .A(n1477), .B(n26350), .Z(n26349) );
  XOR U25750 ( .A(p_input[1194]), .B(n26348), .Z(n26350) );
  XNOR U25751 ( .A(n26351), .B(n26352), .Z(n26348) );
  AND U25752 ( .A(n1481), .B(n26353), .Z(n26352) );
  XOR U25753 ( .A(n26354), .B(n26355), .Z(n26346) );
  AND U25754 ( .A(n1485), .B(n26345), .Z(n26355) );
  XNOR U25755 ( .A(n26356), .B(n26343), .Z(n26345) );
  XOR U25756 ( .A(n26357), .B(n26358), .Z(n26343) );
  AND U25757 ( .A(n1508), .B(n26359), .Z(n26358) );
  IV U25758 ( .A(n26354), .Z(n26356) );
  XOR U25759 ( .A(n26360), .B(n26361), .Z(n26354) );
  AND U25760 ( .A(n1492), .B(n26353), .Z(n26361) );
  XNOR U25761 ( .A(n26351), .B(n26360), .Z(n26353) );
  XNOR U25762 ( .A(n26362), .B(n26363), .Z(n26351) );
  AND U25763 ( .A(n1496), .B(n26364), .Z(n26363) );
  XOR U25764 ( .A(p_input[1210]), .B(n26362), .Z(n26364) );
  XNOR U25765 ( .A(n26365), .B(n26366), .Z(n26362) );
  AND U25766 ( .A(n1500), .B(n26367), .Z(n26366) );
  XOR U25767 ( .A(n26368), .B(n26369), .Z(n26360) );
  AND U25768 ( .A(n1504), .B(n26359), .Z(n26369) );
  XNOR U25769 ( .A(n26370), .B(n26357), .Z(n26359) );
  XOR U25770 ( .A(n26371), .B(n26372), .Z(n26357) );
  AND U25771 ( .A(n1527), .B(n26373), .Z(n26372) );
  IV U25772 ( .A(n26368), .Z(n26370) );
  XOR U25773 ( .A(n26374), .B(n26375), .Z(n26368) );
  AND U25774 ( .A(n1511), .B(n26367), .Z(n26375) );
  XNOR U25775 ( .A(n26365), .B(n26374), .Z(n26367) );
  XNOR U25776 ( .A(n26376), .B(n26377), .Z(n26365) );
  AND U25777 ( .A(n1515), .B(n26378), .Z(n26377) );
  XOR U25778 ( .A(p_input[1226]), .B(n26376), .Z(n26378) );
  XNOR U25779 ( .A(n26379), .B(n26380), .Z(n26376) );
  AND U25780 ( .A(n1519), .B(n26381), .Z(n26380) );
  XOR U25781 ( .A(n26382), .B(n26383), .Z(n26374) );
  AND U25782 ( .A(n1523), .B(n26373), .Z(n26383) );
  XNOR U25783 ( .A(n26384), .B(n26371), .Z(n26373) );
  XOR U25784 ( .A(n26385), .B(n26386), .Z(n26371) );
  AND U25785 ( .A(n1546), .B(n26387), .Z(n26386) );
  IV U25786 ( .A(n26382), .Z(n26384) );
  XOR U25787 ( .A(n26388), .B(n26389), .Z(n26382) );
  AND U25788 ( .A(n1530), .B(n26381), .Z(n26389) );
  XNOR U25789 ( .A(n26379), .B(n26388), .Z(n26381) );
  XNOR U25790 ( .A(n26390), .B(n26391), .Z(n26379) );
  AND U25791 ( .A(n1534), .B(n26392), .Z(n26391) );
  XOR U25792 ( .A(p_input[1242]), .B(n26390), .Z(n26392) );
  XNOR U25793 ( .A(n26393), .B(n26394), .Z(n26390) );
  AND U25794 ( .A(n1538), .B(n26395), .Z(n26394) );
  XOR U25795 ( .A(n26396), .B(n26397), .Z(n26388) );
  AND U25796 ( .A(n1542), .B(n26387), .Z(n26397) );
  XNOR U25797 ( .A(n26398), .B(n26385), .Z(n26387) );
  XOR U25798 ( .A(n26399), .B(n26400), .Z(n26385) );
  AND U25799 ( .A(n1565), .B(n26401), .Z(n26400) );
  IV U25800 ( .A(n26396), .Z(n26398) );
  XOR U25801 ( .A(n26402), .B(n26403), .Z(n26396) );
  AND U25802 ( .A(n1549), .B(n26395), .Z(n26403) );
  XNOR U25803 ( .A(n26393), .B(n26402), .Z(n26395) );
  XNOR U25804 ( .A(n26404), .B(n26405), .Z(n26393) );
  AND U25805 ( .A(n1553), .B(n26406), .Z(n26405) );
  XOR U25806 ( .A(p_input[1258]), .B(n26404), .Z(n26406) );
  XNOR U25807 ( .A(n26407), .B(n26408), .Z(n26404) );
  AND U25808 ( .A(n1557), .B(n26409), .Z(n26408) );
  XOR U25809 ( .A(n26410), .B(n26411), .Z(n26402) );
  AND U25810 ( .A(n1561), .B(n26401), .Z(n26411) );
  XNOR U25811 ( .A(n26412), .B(n26399), .Z(n26401) );
  XOR U25812 ( .A(n26413), .B(n26414), .Z(n26399) );
  AND U25813 ( .A(n1584), .B(n26415), .Z(n26414) );
  IV U25814 ( .A(n26410), .Z(n26412) );
  XOR U25815 ( .A(n26416), .B(n26417), .Z(n26410) );
  AND U25816 ( .A(n1568), .B(n26409), .Z(n26417) );
  XNOR U25817 ( .A(n26407), .B(n26416), .Z(n26409) );
  XNOR U25818 ( .A(n26418), .B(n26419), .Z(n26407) );
  AND U25819 ( .A(n1572), .B(n26420), .Z(n26419) );
  XOR U25820 ( .A(p_input[1274]), .B(n26418), .Z(n26420) );
  XNOR U25821 ( .A(n26421), .B(n26422), .Z(n26418) );
  AND U25822 ( .A(n1576), .B(n26423), .Z(n26422) );
  XOR U25823 ( .A(n26424), .B(n26425), .Z(n26416) );
  AND U25824 ( .A(n1580), .B(n26415), .Z(n26425) );
  XNOR U25825 ( .A(n26426), .B(n26413), .Z(n26415) );
  XOR U25826 ( .A(n26427), .B(n26428), .Z(n26413) );
  AND U25827 ( .A(n1603), .B(n26429), .Z(n26428) );
  IV U25828 ( .A(n26424), .Z(n26426) );
  XOR U25829 ( .A(n26430), .B(n26431), .Z(n26424) );
  AND U25830 ( .A(n1587), .B(n26423), .Z(n26431) );
  XNOR U25831 ( .A(n26421), .B(n26430), .Z(n26423) );
  XNOR U25832 ( .A(n26432), .B(n26433), .Z(n26421) );
  AND U25833 ( .A(n1591), .B(n26434), .Z(n26433) );
  XOR U25834 ( .A(p_input[1290]), .B(n26432), .Z(n26434) );
  XNOR U25835 ( .A(n26435), .B(n26436), .Z(n26432) );
  AND U25836 ( .A(n1595), .B(n26437), .Z(n26436) );
  XOR U25837 ( .A(n26438), .B(n26439), .Z(n26430) );
  AND U25838 ( .A(n1599), .B(n26429), .Z(n26439) );
  XNOR U25839 ( .A(n26440), .B(n26427), .Z(n26429) );
  XOR U25840 ( .A(n26441), .B(n26442), .Z(n26427) );
  AND U25841 ( .A(n1622), .B(n26443), .Z(n26442) );
  IV U25842 ( .A(n26438), .Z(n26440) );
  XOR U25843 ( .A(n26444), .B(n26445), .Z(n26438) );
  AND U25844 ( .A(n1606), .B(n26437), .Z(n26445) );
  XNOR U25845 ( .A(n26435), .B(n26444), .Z(n26437) );
  XNOR U25846 ( .A(n26446), .B(n26447), .Z(n26435) );
  AND U25847 ( .A(n1610), .B(n26448), .Z(n26447) );
  XOR U25848 ( .A(p_input[1306]), .B(n26446), .Z(n26448) );
  XNOR U25849 ( .A(n26449), .B(n26450), .Z(n26446) );
  AND U25850 ( .A(n1614), .B(n26451), .Z(n26450) );
  XOR U25851 ( .A(n26452), .B(n26453), .Z(n26444) );
  AND U25852 ( .A(n1618), .B(n26443), .Z(n26453) );
  XNOR U25853 ( .A(n26454), .B(n26441), .Z(n26443) );
  XOR U25854 ( .A(n26455), .B(n26456), .Z(n26441) );
  AND U25855 ( .A(n1641), .B(n26457), .Z(n26456) );
  IV U25856 ( .A(n26452), .Z(n26454) );
  XOR U25857 ( .A(n26458), .B(n26459), .Z(n26452) );
  AND U25858 ( .A(n1625), .B(n26451), .Z(n26459) );
  XNOR U25859 ( .A(n26449), .B(n26458), .Z(n26451) );
  XNOR U25860 ( .A(n26460), .B(n26461), .Z(n26449) );
  AND U25861 ( .A(n1629), .B(n26462), .Z(n26461) );
  XOR U25862 ( .A(p_input[1322]), .B(n26460), .Z(n26462) );
  XNOR U25863 ( .A(n26463), .B(n26464), .Z(n26460) );
  AND U25864 ( .A(n1633), .B(n26465), .Z(n26464) );
  XOR U25865 ( .A(n26466), .B(n26467), .Z(n26458) );
  AND U25866 ( .A(n1637), .B(n26457), .Z(n26467) );
  XNOR U25867 ( .A(n26468), .B(n26455), .Z(n26457) );
  XOR U25868 ( .A(n26469), .B(n26470), .Z(n26455) );
  AND U25869 ( .A(n1660), .B(n26471), .Z(n26470) );
  IV U25870 ( .A(n26466), .Z(n26468) );
  XOR U25871 ( .A(n26472), .B(n26473), .Z(n26466) );
  AND U25872 ( .A(n1644), .B(n26465), .Z(n26473) );
  XNOR U25873 ( .A(n26463), .B(n26472), .Z(n26465) );
  XNOR U25874 ( .A(n26474), .B(n26475), .Z(n26463) );
  AND U25875 ( .A(n1648), .B(n26476), .Z(n26475) );
  XOR U25876 ( .A(p_input[1338]), .B(n26474), .Z(n26476) );
  XNOR U25877 ( .A(n26477), .B(n26478), .Z(n26474) );
  AND U25878 ( .A(n1652), .B(n26479), .Z(n26478) );
  XOR U25879 ( .A(n26480), .B(n26481), .Z(n26472) );
  AND U25880 ( .A(n1656), .B(n26471), .Z(n26481) );
  XNOR U25881 ( .A(n26482), .B(n26469), .Z(n26471) );
  XOR U25882 ( .A(n26483), .B(n26484), .Z(n26469) );
  AND U25883 ( .A(n1679), .B(n26485), .Z(n26484) );
  IV U25884 ( .A(n26480), .Z(n26482) );
  XOR U25885 ( .A(n26486), .B(n26487), .Z(n26480) );
  AND U25886 ( .A(n1663), .B(n26479), .Z(n26487) );
  XNOR U25887 ( .A(n26477), .B(n26486), .Z(n26479) );
  XNOR U25888 ( .A(n26488), .B(n26489), .Z(n26477) );
  AND U25889 ( .A(n1667), .B(n26490), .Z(n26489) );
  XOR U25890 ( .A(p_input[1354]), .B(n26488), .Z(n26490) );
  XNOR U25891 ( .A(n26491), .B(n26492), .Z(n26488) );
  AND U25892 ( .A(n1671), .B(n26493), .Z(n26492) );
  XOR U25893 ( .A(n26494), .B(n26495), .Z(n26486) );
  AND U25894 ( .A(n1675), .B(n26485), .Z(n26495) );
  XNOR U25895 ( .A(n26496), .B(n26483), .Z(n26485) );
  XOR U25896 ( .A(n26497), .B(n26498), .Z(n26483) );
  AND U25897 ( .A(n1698), .B(n26499), .Z(n26498) );
  IV U25898 ( .A(n26494), .Z(n26496) );
  XOR U25899 ( .A(n26500), .B(n26501), .Z(n26494) );
  AND U25900 ( .A(n1682), .B(n26493), .Z(n26501) );
  XNOR U25901 ( .A(n26491), .B(n26500), .Z(n26493) );
  XNOR U25902 ( .A(n26502), .B(n26503), .Z(n26491) );
  AND U25903 ( .A(n1686), .B(n26504), .Z(n26503) );
  XOR U25904 ( .A(p_input[1370]), .B(n26502), .Z(n26504) );
  XNOR U25905 ( .A(n26505), .B(n26506), .Z(n26502) );
  AND U25906 ( .A(n1690), .B(n26507), .Z(n26506) );
  XOR U25907 ( .A(n26508), .B(n26509), .Z(n26500) );
  AND U25908 ( .A(n1694), .B(n26499), .Z(n26509) );
  XNOR U25909 ( .A(n26510), .B(n26497), .Z(n26499) );
  XOR U25910 ( .A(n26511), .B(n26512), .Z(n26497) );
  AND U25911 ( .A(n1717), .B(n26513), .Z(n26512) );
  IV U25912 ( .A(n26508), .Z(n26510) );
  XOR U25913 ( .A(n26514), .B(n26515), .Z(n26508) );
  AND U25914 ( .A(n1701), .B(n26507), .Z(n26515) );
  XNOR U25915 ( .A(n26505), .B(n26514), .Z(n26507) );
  XNOR U25916 ( .A(n26516), .B(n26517), .Z(n26505) );
  AND U25917 ( .A(n1705), .B(n26518), .Z(n26517) );
  XOR U25918 ( .A(p_input[1386]), .B(n26516), .Z(n26518) );
  XNOR U25919 ( .A(n26519), .B(n26520), .Z(n26516) );
  AND U25920 ( .A(n1709), .B(n26521), .Z(n26520) );
  XOR U25921 ( .A(n26522), .B(n26523), .Z(n26514) );
  AND U25922 ( .A(n1713), .B(n26513), .Z(n26523) );
  XNOR U25923 ( .A(n26524), .B(n26511), .Z(n26513) );
  XOR U25924 ( .A(n26525), .B(n26526), .Z(n26511) );
  AND U25925 ( .A(n1736), .B(n26527), .Z(n26526) );
  IV U25926 ( .A(n26522), .Z(n26524) );
  XOR U25927 ( .A(n26528), .B(n26529), .Z(n26522) );
  AND U25928 ( .A(n1720), .B(n26521), .Z(n26529) );
  XNOR U25929 ( .A(n26519), .B(n26528), .Z(n26521) );
  XNOR U25930 ( .A(n26530), .B(n26531), .Z(n26519) );
  AND U25931 ( .A(n1724), .B(n26532), .Z(n26531) );
  XOR U25932 ( .A(p_input[1402]), .B(n26530), .Z(n26532) );
  XNOR U25933 ( .A(n26533), .B(n26534), .Z(n26530) );
  AND U25934 ( .A(n1728), .B(n26535), .Z(n26534) );
  XOR U25935 ( .A(n26536), .B(n26537), .Z(n26528) );
  AND U25936 ( .A(n1732), .B(n26527), .Z(n26537) );
  XNOR U25937 ( .A(n26538), .B(n26525), .Z(n26527) );
  XOR U25938 ( .A(n26539), .B(n26540), .Z(n26525) );
  AND U25939 ( .A(n1755), .B(n26541), .Z(n26540) );
  IV U25940 ( .A(n26536), .Z(n26538) );
  XOR U25941 ( .A(n26542), .B(n26543), .Z(n26536) );
  AND U25942 ( .A(n1739), .B(n26535), .Z(n26543) );
  XNOR U25943 ( .A(n26533), .B(n26542), .Z(n26535) );
  XNOR U25944 ( .A(n26544), .B(n26545), .Z(n26533) );
  AND U25945 ( .A(n1743), .B(n26546), .Z(n26545) );
  XOR U25946 ( .A(p_input[1418]), .B(n26544), .Z(n26546) );
  XNOR U25947 ( .A(n26547), .B(n26548), .Z(n26544) );
  AND U25948 ( .A(n1747), .B(n26549), .Z(n26548) );
  XOR U25949 ( .A(n26550), .B(n26551), .Z(n26542) );
  AND U25950 ( .A(n1751), .B(n26541), .Z(n26551) );
  XNOR U25951 ( .A(n26552), .B(n26539), .Z(n26541) );
  XOR U25952 ( .A(n26553), .B(n26554), .Z(n26539) );
  AND U25953 ( .A(n1774), .B(n26555), .Z(n26554) );
  IV U25954 ( .A(n26550), .Z(n26552) );
  XOR U25955 ( .A(n26556), .B(n26557), .Z(n26550) );
  AND U25956 ( .A(n1758), .B(n26549), .Z(n26557) );
  XNOR U25957 ( .A(n26547), .B(n26556), .Z(n26549) );
  XNOR U25958 ( .A(n26558), .B(n26559), .Z(n26547) );
  AND U25959 ( .A(n1762), .B(n26560), .Z(n26559) );
  XOR U25960 ( .A(p_input[1434]), .B(n26558), .Z(n26560) );
  XNOR U25961 ( .A(n26561), .B(n26562), .Z(n26558) );
  AND U25962 ( .A(n1766), .B(n26563), .Z(n26562) );
  XOR U25963 ( .A(n26564), .B(n26565), .Z(n26556) );
  AND U25964 ( .A(n1770), .B(n26555), .Z(n26565) );
  XNOR U25965 ( .A(n26566), .B(n26553), .Z(n26555) );
  XOR U25966 ( .A(n26567), .B(n26568), .Z(n26553) );
  AND U25967 ( .A(n1793), .B(n26569), .Z(n26568) );
  IV U25968 ( .A(n26564), .Z(n26566) );
  XOR U25969 ( .A(n26570), .B(n26571), .Z(n26564) );
  AND U25970 ( .A(n1777), .B(n26563), .Z(n26571) );
  XNOR U25971 ( .A(n26561), .B(n26570), .Z(n26563) );
  XNOR U25972 ( .A(n26572), .B(n26573), .Z(n26561) );
  AND U25973 ( .A(n1781), .B(n26574), .Z(n26573) );
  XOR U25974 ( .A(p_input[1450]), .B(n26572), .Z(n26574) );
  XNOR U25975 ( .A(n26575), .B(n26576), .Z(n26572) );
  AND U25976 ( .A(n1785), .B(n26577), .Z(n26576) );
  XOR U25977 ( .A(n26578), .B(n26579), .Z(n26570) );
  AND U25978 ( .A(n1789), .B(n26569), .Z(n26579) );
  XNOR U25979 ( .A(n26580), .B(n26567), .Z(n26569) );
  XOR U25980 ( .A(n26581), .B(n26582), .Z(n26567) );
  AND U25981 ( .A(n1812), .B(n26583), .Z(n26582) );
  IV U25982 ( .A(n26578), .Z(n26580) );
  XOR U25983 ( .A(n26584), .B(n26585), .Z(n26578) );
  AND U25984 ( .A(n1796), .B(n26577), .Z(n26585) );
  XNOR U25985 ( .A(n26575), .B(n26584), .Z(n26577) );
  XNOR U25986 ( .A(n26586), .B(n26587), .Z(n26575) );
  AND U25987 ( .A(n1800), .B(n26588), .Z(n26587) );
  XOR U25988 ( .A(p_input[1466]), .B(n26586), .Z(n26588) );
  XNOR U25989 ( .A(n26589), .B(n26590), .Z(n26586) );
  AND U25990 ( .A(n1804), .B(n26591), .Z(n26590) );
  XOR U25991 ( .A(n26592), .B(n26593), .Z(n26584) );
  AND U25992 ( .A(n1808), .B(n26583), .Z(n26593) );
  XNOR U25993 ( .A(n26594), .B(n26581), .Z(n26583) );
  XOR U25994 ( .A(n26595), .B(n26596), .Z(n26581) );
  AND U25995 ( .A(n1831), .B(n26597), .Z(n26596) );
  IV U25996 ( .A(n26592), .Z(n26594) );
  XOR U25997 ( .A(n26598), .B(n26599), .Z(n26592) );
  AND U25998 ( .A(n1815), .B(n26591), .Z(n26599) );
  XNOR U25999 ( .A(n26589), .B(n26598), .Z(n26591) );
  XNOR U26000 ( .A(n26600), .B(n26601), .Z(n26589) );
  AND U26001 ( .A(n1819), .B(n26602), .Z(n26601) );
  XOR U26002 ( .A(p_input[1482]), .B(n26600), .Z(n26602) );
  XNOR U26003 ( .A(n26603), .B(n26604), .Z(n26600) );
  AND U26004 ( .A(n1823), .B(n26605), .Z(n26604) );
  XOR U26005 ( .A(n26606), .B(n26607), .Z(n26598) );
  AND U26006 ( .A(n1827), .B(n26597), .Z(n26607) );
  XNOR U26007 ( .A(n26608), .B(n26595), .Z(n26597) );
  XOR U26008 ( .A(n26609), .B(n26610), .Z(n26595) );
  AND U26009 ( .A(n1850), .B(n26611), .Z(n26610) );
  IV U26010 ( .A(n26606), .Z(n26608) );
  XOR U26011 ( .A(n26612), .B(n26613), .Z(n26606) );
  AND U26012 ( .A(n1834), .B(n26605), .Z(n26613) );
  XNOR U26013 ( .A(n26603), .B(n26612), .Z(n26605) );
  XNOR U26014 ( .A(n26614), .B(n26615), .Z(n26603) );
  AND U26015 ( .A(n1838), .B(n26616), .Z(n26615) );
  XOR U26016 ( .A(p_input[1498]), .B(n26614), .Z(n26616) );
  XNOR U26017 ( .A(n26617), .B(n26618), .Z(n26614) );
  AND U26018 ( .A(n1842), .B(n26619), .Z(n26618) );
  XOR U26019 ( .A(n26620), .B(n26621), .Z(n26612) );
  AND U26020 ( .A(n1846), .B(n26611), .Z(n26621) );
  XNOR U26021 ( .A(n26622), .B(n26609), .Z(n26611) );
  XOR U26022 ( .A(n26623), .B(n26624), .Z(n26609) );
  AND U26023 ( .A(n1869), .B(n26625), .Z(n26624) );
  IV U26024 ( .A(n26620), .Z(n26622) );
  XOR U26025 ( .A(n26626), .B(n26627), .Z(n26620) );
  AND U26026 ( .A(n1853), .B(n26619), .Z(n26627) );
  XNOR U26027 ( .A(n26617), .B(n26626), .Z(n26619) );
  XNOR U26028 ( .A(n26628), .B(n26629), .Z(n26617) );
  AND U26029 ( .A(n1857), .B(n26630), .Z(n26629) );
  XOR U26030 ( .A(p_input[1514]), .B(n26628), .Z(n26630) );
  XNOR U26031 ( .A(n26631), .B(n26632), .Z(n26628) );
  AND U26032 ( .A(n1861), .B(n26633), .Z(n26632) );
  XOR U26033 ( .A(n26634), .B(n26635), .Z(n26626) );
  AND U26034 ( .A(n1865), .B(n26625), .Z(n26635) );
  XNOR U26035 ( .A(n26636), .B(n26623), .Z(n26625) );
  XOR U26036 ( .A(n26637), .B(n26638), .Z(n26623) );
  AND U26037 ( .A(n1888), .B(n26639), .Z(n26638) );
  IV U26038 ( .A(n26634), .Z(n26636) );
  XOR U26039 ( .A(n26640), .B(n26641), .Z(n26634) );
  AND U26040 ( .A(n1872), .B(n26633), .Z(n26641) );
  XNOR U26041 ( .A(n26631), .B(n26640), .Z(n26633) );
  XNOR U26042 ( .A(n26642), .B(n26643), .Z(n26631) );
  AND U26043 ( .A(n1876), .B(n26644), .Z(n26643) );
  XOR U26044 ( .A(p_input[1530]), .B(n26642), .Z(n26644) );
  XNOR U26045 ( .A(n26645), .B(n26646), .Z(n26642) );
  AND U26046 ( .A(n1880), .B(n26647), .Z(n26646) );
  XOR U26047 ( .A(n26648), .B(n26649), .Z(n26640) );
  AND U26048 ( .A(n1884), .B(n26639), .Z(n26649) );
  XNOR U26049 ( .A(n26650), .B(n26637), .Z(n26639) );
  XOR U26050 ( .A(n26651), .B(n26652), .Z(n26637) );
  AND U26051 ( .A(n1907), .B(n26653), .Z(n26652) );
  IV U26052 ( .A(n26648), .Z(n26650) );
  XOR U26053 ( .A(n26654), .B(n26655), .Z(n26648) );
  AND U26054 ( .A(n1891), .B(n26647), .Z(n26655) );
  XNOR U26055 ( .A(n26645), .B(n26654), .Z(n26647) );
  XNOR U26056 ( .A(n26656), .B(n26657), .Z(n26645) );
  AND U26057 ( .A(n1895), .B(n26658), .Z(n26657) );
  XOR U26058 ( .A(p_input[1546]), .B(n26656), .Z(n26658) );
  XNOR U26059 ( .A(n26659), .B(n26660), .Z(n26656) );
  AND U26060 ( .A(n1899), .B(n26661), .Z(n26660) );
  XOR U26061 ( .A(n26662), .B(n26663), .Z(n26654) );
  AND U26062 ( .A(n1903), .B(n26653), .Z(n26663) );
  XNOR U26063 ( .A(n26664), .B(n26651), .Z(n26653) );
  XOR U26064 ( .A(n26665), .B(n26666), .Z(n26651) );
  AND U26065 ( .A(n1926), .B(n26667), .Z(n26666) );
  IV U26066 ( .A(n26662), .Z(n26664) );
  XOR U26067 ( .A(n26668), .B(n26669), .Z(n26662) );
  AND U26068 ( .A(n1910), .B(n26661), .Z(n26669) );
  XNOR U26069 ( .A(n26659), .B(n26668), .Z(n26661) );
  XNOR U26070 ( .A(n26670), .B(n26671), .Z(n26659) );
  AND U26071 ( .A(n1914), .B(n26672), .Z(n26671) );
  XOR U26072 ( .A(p_input[1562]), .B(n26670), .Z(n26672) );
  XNOR U26073 ( .A(n26673), .B(n26674), .Z(n26670) );
  AND U26074 ( .A(n1918), .B(n26675), .Z(n26674) );
  XOR U26075 ( .A(n26676), .B(n26677), .Z(n26668) );
  AND U26076 ( .A(n1922), .B(n26667), .Z(n26677) );
  XNOR U26077 ( .A(n26678), .B(n26665), .Z(n26667) );
  XOR U26078 ( .A(n26679), .B(n26680), .Z(n26665) );
  AND U26079 ( .A(n1945), .B(n26681), .Z(n26680) );
  IV U26080 ( .A(n26676), .Z(n26678) );
  XOR U26081 ( .A(n26682), .B(n26683), .Z(n26676) );
  AND U26082 ( .A(n1929), .B(n26675), .Z(n26683) );
  XNOR U26083 ( .A(n26673), .B(n26682), .Z(n26675) );
  XNOR U26084 ( .A(n26684), .B(n26685), .Z(n26673) );
  AND U26085 ( .A(n1933), .B(n26686), .Z(n26685) );
  XOR U26086 ( .A(p_input[1578]), .B(n26684), .Z(n26686) );
  XNOR U26087 ( .A(n26687), .B(n26688), .Z(n26684) );
  AND U26088 ( .A(n1937), .B(n26689), .Z(n26688) );
  XOR U26089 ( .A(n26690), .B(n26691), .Z(n26682) );
  AND U26090 ( .A(n1941), .B(n26681), .Z(n26691) );
  XNOR U26091 ( .A(n26692), .B(n26679), .Z(n26681) );
  XOR U26092 ( .A(n26693), .B(n26694), .Z(n26679) );
  AND U26093 ( .A(n1964), .B(n26695), .Z(n26694) );
  IV U26094 ( .A(n26690), .Z(n26692) );
  XOR U26095 ( .A(n26696), .B(n26697), .Z(n26690) );
  AND U26096 ( .A(n1948), .B(n26689), .Z(n26697) );
  XNOR U26097 ( .A(n26687), .B(n26696), .Z(n26689) );
  XNOR U26098 ( .A(n26698), .B(n26699), .Z(n26687) );
  AND U26099 ( .A(n1952), .B(n26700), .Z(n26699) );
  XOR U26100 ( .A(p_input[1594]), .B(n26698), .Z(n26700) );
  XNOR U26101 ( .A(n26701), .B(n26702), .Z(n26698) );
  AND U26102 ( .A(n1956), .B(n26703), .Z(n26702) );
  XOR U26103 ( .A(n26704), .B(n26705), .Z(n26696) );
  AND U26104 ( .A(n1960), .B(n26695), .Z(n26705) );
  XNOR U26105 ( .A(n26706), .B(n26693), .Z(n26695) );
  XOR U26106 ( .A(n26707), .B(n26708), .Z(n26693) );
  AND U26107 ( .A(n1983), .B(n26709), .Z(n26708) );
  IV U26108 ( .A(n26704), .Z(n26706) );
  XOR U26109 ( .A(n26710), .B(n26711), .Z(n26704) );
  AND U26110 ( .A(n1967), .B(n26703), .Z(n26711) );
  XNOR U26111 ( .A(n26701), .B(n26710), .Z(n26703) );
  XNOR U26112 ( .A(n26712), .B(n26713), .Z(n26701) );
  AND U26113 ( .A(n1971), .B(n26714), .Z(n26713) );
  XOR U26114 ( .A(p_input[1610]), .B(n26712), .Z(n26714) );
  XNOR U26115 ( .A(n26715), .B(n26716), .Z(n26712) );
  AND U26116 ( .A(n1975), .B(n26717), .Z(n26716) );
  XOR U26117 ( .A(n26718), .B(n26719), .Z(n26710) );
  AND U26118 ( .A(n1979), .B(n26709), .Z(n26719) );
  XNOR U26119 ( .A(n26720), .B(n26707), .Z(n26709) );
  XOR U26120 ( .A(n26721), .B(n26722), .Z(n26707) );
  AND U26121 ( .A(n2002), .B(n26723), .Z(n26722) );
  IV U26122 ( .A(n26718), .Z(n26720) );
  XOR U26123 ( .A(n26724), .B(n26725), .Z(n26718) );
  AND U26124 ( .A(n1986), .B(n26717), .Z(n26725) );
  XNOR U26125 ( .A(n26715), .B(n26724), .Z(n26717) );
  XNOR U26126 ( .A(n26726), .B(n26727), .Z(n26715) );
  AND U26127 ( .A(n1990), .B(n26728), .Z(n26727) );
  XOR U26128 ( .A(p_input[1626]), .B(n26726), .Z(n26728) );
  XNOR U26129 ( .A(n26729), .B(n26730), .Z(n26726) );
  AND U26130 ( .A(n1994), .B(n26731), .Z(n26730) );
  XOR U26131 ( .A(n26732), .B(n26733), .Z(n26724) );
  AND U26132 ( .A(n1998), .B(n26723), .Z(n26733) );
  XNOR U26133 ( .A(n26734), .B(n26721), .Z(n26723) );
  XOR U26134 ( .A(n26735), .B(n26736), .Z(n26721) );
  AND U26135 ( .A(n2021), .B(n26737), .Z(n26736) );
  IV U26136 ( .A(n26732), .Z(n26734) );
  XOR U26137 ( .A(n26738), .B(n26739), .Z(n26732) );
  AND U26138 ( .A(n2005), .B(n26731), .Z(n26739) );
  XNOR U26139 ( .A(n26729), .B(n26738), .Z(n26731) );
  XNOR U26140 ( .A(n26740), .B(n26741), .Z(n26729) );
  AND U26141 ( .A(n2009), .B(n26742), .Z(n26741) );
  XOR U26142 ( .A(p_input[1642]), .B(n26740), .Z(n26742) );
  XNOR U26143 ( .A(n26743), .B(n26744), .Z(n26740) );
  AND U26144 ( .A(n2013), .B(n26745), .Z(n26744) );
  XOR U26145 ( .A(n26746), .B(n26747), .Z(n26738) );
  AND U26146 ( .A(n2017), .B(n26737), .Z(n26747) );
  XNOR U26147 ( .A(n26748), .B(n26735), .Z(n26737) );
  XOR U26148 ( .A(n26749), .B(n26750), .Z(n26735) );
  AND U26149 ( .A(n2040), .B(n26751), .Z(n26750) );
  IV U26150 ( .A(n26746), .Z(n26748) );
  XOR U26151 ( .A(n26752), .B(n26753), .Z(n26746) );
  AND U26152 ( .A(n2024), .B(n26745), .Z(n26753) );
  XNOR U26153 ( .A(n26743), .B(n26752), .Z(n26745) );
  XNOR U26154 ( .A(n26754), .B(n26755), .Z(n26743) );
  AND U26155 ( .A(n2028), .B(n26756), .Z(n26755) );
  XOR U26156 ( .A(p_input[1658]), .B(n26754), .Z(n26756) );
  XNOR U26157 ( .A(n26757), .B(n26758), .Z(n26754) );
  AND U26158 ( .A(n2032), .B(n26759), .Z(n26758) );
  XOR U26159 ( .A(n26760), .B(n26761), .Z(n26752) );
  AND U26160 ( .A(n2036), .B(n26751), .Z(n26761) );
  XNOR U26161 ( .A(n26762), .B(n26749), .Z(n26751) );
  XOR U26162 ( .A(n26763), .B(n26764), .Z(n26749) );
  AND U26163 ( .A(n2059), .B(n26765), .Z(n26764) );
  IV U26164 ( .A(n26760), .Z(n26762) );
  XOR U26165 ( .A(n26766), .B(n26767), .Z(n26760) );
  AND U26166 ( .A(n2043), .B(n26759), .Z(n26767) );
  XNOR U26167 ( .A(n26757), .B(n26766), .Z(n26759) );
  XNOR U26168 ( .A(n26768), .B(n26769), .Z(n26757) );
  AND U26169 ( .A(n2047), .B(n26770), .Z(n26769) );
  XOR U26170 ( .A(p_input[1674]), .B(n26768), .Z(n26770) );
  XNOR U26171 ( .A(n26771), .B(n26772), .Z(n26768) );
  AND U26172 ( .A(n2051), .B(n26773), .Z(n26772) );
  XOR U26173 ( .A(n26774), .B(n26775), .Z(n26766) );
  AND U26174 ( .A(n2055), .B(n26765), .Z(n26775) );
  XNOR U26175 ( .A(n26776), .B(n26763), .Z(n26765) );
  XOR U26176 ( .A(n26777), .B(n26778), .Z(n26763) );
  AND U26177 ( .A(n2078), .B(n26779), .Z(n26778) );
  IV U26178 ( .A(n26774), .Z(n26776) );
  XOR U26179 ( .A(n26780), .B(n26781), .Z(n26774) );
  AND U26180 ( .A(n2062), .B(n26773), .Z(n26781) );
  XNOR U26181 ( .A(n26771), .B(n26780), .Z(n26773) );
  XNOR U26182 ( .A(n26782), .B(n26783), .Z(n26771) );
  AND U26183 ( .A(n2066), .B(n26784), .Z(n26783) );
  XOR U26184 ( .A(p_input[1690]), .B(n26782), .Z(n26784) );
  XNOR U26185 ( .A(n26785), .B(n26786), .Z(n26782) );
  AND U26186 ( .A(n2070), .B(n26787), .Z(n26786) );
  XOR U26187 ( .A(n26788), .B(n26789), .Z(n26780) );
  AND U26188 ( .A(n2074), .B(n26779), .Z(n26789) );
  XNOR U26189 ( .A(n26790), .B(n26777), .Z(n26779) );
  XOR U26190 ( .A(n26791), .B(n26792), .Z(n26777) );
  AND U26191 ( .A(n2097), .B(n26793), .Z(n26792) );
  IV U26192 ( .A(n26788), .Z(n26790) );
  XOR U26193 ( .A(n26794), .B(n26795), .Z(n26788) );
  AND U26194 ( .A(n2081), .B(n26787), .Z(n26795) );
  XNOR U26195 ( .A(n26785), .B(n26794), .Z(n26787) );
  XNOR U26196 ( .A(n26796), .B(n26797), .Z(n26785) );
  AND U26197 ( .A(n2085), .B(n26798), .Z(n26797) );
  XOR U26198 ( .A(p_input[1706]), .B(n26796), .Z(n26798) );
  XNOR U26199 ( .A(n26799), .B(n26800), .Z(n26796) );
  AND U26200 ( .A(n2089), .B(n26801), .Z(n26800) );
  XOR U26201 ( .A(n26802), .B(n26803), .Z(n26794) );
  AND U26202 ( .A(n2093), .B(n26793), .Z(n26803) );
  XNOR U26203 ( .A(n26804), .B(n26791), .Z(n26793) );
  XOR U26204 ( .A(n26805), .B(n26806), .Z(n26791) );
  AND U26205 ( .A(n2116), .B(n26807), .Z(n26806) );
  IV U26206 ( .A(n26802), .Z(n26804) );
  XOR U26207 ( .A(n26808), .B(n26809), .Z(n26802) );
  AND U26208 ( .A(n2100), .B(n26801), .Z(n26809) );
  XNOR U26209 ( .A(n26799), .B(n26808), .Z(n26801) );
  XNOR U26210 ( .A(n26810), .B(n26811), .Z(n26799) );
  AND U26211 ( .A(n2104), .B(n26812), .Z(n26811) );
  XOR U26212 ( .A(p_input[1722]), .B(n26810), .Z(n26812) );
  XNOR U26213 ( .A(n26813), .B(n26814), .Z(n26810) );
  AND U26214 ( .A(n2108), .B(n26815), .Z(n26814) );
  XOR U26215 ( .A(n26816), .B(n26817), .Z(n26808) );
  AND U26216 ( .A(n2112), .B(n26807), .Z(n26817) );
  XNOR U26217 ( .A(n26818), .B(n26805), .Z(n26807) );
  XOR U26218 ( .A(n26819), .B(n26820), .Z(n26805) );
  AND U26219 ( .A(n2135), .B(n26821), .Z(n26820) );
  IV U26220 ( .A(n26816), .Z(n26818) );
  XOR U26221 ( .A(n26822), .B(n26823), .Z(n26816) );
  AND U26222 ( .A(n2119), .B(n26815), .Z(n26823) );
  XNOR U26223 ( .A(n26813), .B(n26822), .Z(n26815) );
  XNOR U26224 ( .A(n26824), .B(n26825), .Z(n26813) );
  AND U26225 ( .A(n2123), .B(n26826), .Z(n26825) );
  XOR U26226 ( .A(p_input[1738]), .B(n26824), .Z(n26826) );
  XNOR U26227 ( .A(n26827), .B(n26828), .Z(n26824) );
  AND U26228 ( .A(n2127), .B(n26829), .Z(n26828) );
  XOR U26229 ( .A(n26830), .B(n26831), .Z(n26822) );
  AND U26230 ( .A(n2131), .B(n26821), .Z(n26831) );
  XNOR U26231 ( .A(n26832), .B(n26819), .Z(n26821) );
  XOR U26232 ( .A(n26833), .B(n26834), .Z(n26819) );
  AND U26233 ( .A(n2154), .B(n26835), .Z(n26834) );
  IV U26234 ( .A(n26830), .Z(n26832) );
  XOR U26235 ( .A(n26836), .B(n26837), .Z(n26830) );
  AND U26236 ( .A(n2138), .B(n26829), .Z(n26837) );
  XNOR U26237 ( .A(n26827), .B(n26836), .Z(n26829) );
  XNOR U26238 ( .A(n26838), .B(n26839), .Z(n26827) );
  AND U26239 ( .A(n2142), .B(n26840), .Z(n26839) );
  XOR U26240 ( .A(p_input[1754]), .B(n26838), .Z(n26840) );
  XNOR U26241 ( .A(n26841), .B(n26842), .Z(n26838) );
  AND U26242 ( .A(n2146), .B(n26843), .Z(n26842) );
  XOR U26243 ( .A(n26844), .B(n26845), .Z(n26836) );
  AND U26244 ( .A(n2150), .B(n26835), .Z(n26845) );
  XNOR U26245 ( .A(n26846), .B(n26833), .Z(n26835) );
  XOR U26246 ( .A(n26847), .B(n26848), .Z(n26833) );
  AND U26247 ( .A(n2173), .B(n26849), .Z(n26848) );
  IV U26248 ( .A(n26844), .Z(n26846) );
  XOR U26249 ( .A(n26850), .B(n26851), .Z(n26844) );
  AND U26250 ( .A(n2157), .B(n26843), .Z(n26851) );
  XNOR U26251 ( .A(n26841), .B(n26850), .Z(n26843) );
  XNOR U26252 ( .A(n26852), .B(n26853), .Z(n26841) );
  AND U26253 ( .A(n2161), .B(n26854), .Z(n26853) );
  XOR U26254 ( .A(p_input[1770]), .B(n26852), .Z(n26854) );
  XNOR U26255 ( .A(n26855), .B(n26856), .Z(n26852) );
  AND U26256 ( .A(n2165), .B(n26857), .Z(n26856) );
  XOR U26257 ( .A(n26858), .B(n26859), .Z(n26850) );
  AND U26258 ( .A(n2169), .B(n26849), .Z(n26859) );
  XNOR U26259 ( .A(n26860), .B(n26847), .Z(n26849) );
  XOR U26260 ( .A(n26861), .B(n26862), .Z(n26847) );
  AND U26261 ( .A(n2192), .B(n26863), .Z(n26862) );
  IV U26262 ( .A(n26858), .Z(n26860) );
  XOR U26263 ( .A(n26864), .B(n26865), .Z(n26858) );
  AND U26264 ( .A(n2176), .B(n26857), .Z(n26865) );
  XNOR U26265 ( .A(n26855), .B(n26864), .Z(n26857) );
  XNOR U26266 ( .A(n26866), .B(n26867), .Z(n26855) );
  AND U26267 ( .A(n2180), .B(n26868), .Z(n26867) );
  XOR U26268 ( .A(p_input[1786]), .B(n26866), .Z(n26868) );
  XNOR U26269 ( .A(n26869), .B(n26870), .Z(n26866) );
  AND U26270 ( .A(n2184), .B(n26871), .Z(n26870) );
  XOR U26271 ( .A(n26872), .B(n26873), .Z(n26864) );
  AND U26272 ( .A(n2188), .B(n26863), .Z(n26873) );
  XNOR U26273 ( .A(n26874), .B(n26861), .Z(n26863) );
  XOR U26274 ( .A(n26875), .B(n26876), .Z(n26861) );
  AND U26275 ( .A(n2211), .B(n26877), .Z(n26876) );
  IV U26276 ( .A(n26872), .Z(n26874) );
  XOR U26277 ( .A(n26878), .B(n26879), .Z(n26872) );
  AND U26278 ( .A(n2195), .B(n26871), .Z(n26879) );
  XNOR U26279 ( .A(n26869), .B(n26878), .Z(n26871) );
  XNOR U26280 ( .A(n26880), .B(n26881), .Z(n26869) );
  AND U26281 ( .A(n2199), .B(n26882), .Z(n26881) );
  XOR U26282 ( .A(p_input[1802]), .B(n26880), .Z(n26882) );
  XNOR U26283 ( .A(n26883), .B(n26884), .Z(n26880) );
  AND U26284 ( .A(n2203), .B(n26885), .Z(n26884) );
  XOR U26285 ( .A(n26886), .B(n26887), .Z(n26878) );
  AND U26286 ( .A(n2207), .B(n26877), .Z(n26887) );
  XNOR U26287 ( .A(n26888), .B(n26875), .Z(n26877) );
  XOR U26288 ( .A(n26889), .B(n26890), .Z(n26875) );
  AND U26289 ( .A(n2230), .B(n26891), .Z(n26890) );
  IV U26290 ( .A(n26886), .Z(n26888) );
  XOR U26291 ( .A(n26892), .B(n26893), .Z(n26886) );
  AND U26292 ( .A(n2214), .B(n26885), .Z(n26893) );
  XNOR U26293 ( .A(n26883), .B(n26892), .Z(n26885) );
  XNOR U26294 ( .A(n26894), .B(n26895), .Z(n26883) );
  AND U26295 ( .A(n2218), .B(n26896), .Z(n26895) );
  XOR U26296 ( .A(p_input[1818]), .B(n26894), .Z(n26896) );
  XNOR U26297 ( .A(n26897), .B(n26898), .Z(n26894) );
  AND U26298 ( .A(n2222), .B(n26899), .Z(n26898) );
  XOR U26299 ( .A(n26900), .B(n26901), .Z(n26892) );
  AND U26300 ( .A(n2226), .B(n26891), .Z(n26901) );
  XNOR U26301 ( .A(n26902), .B(n26889), .Z(n26891) );
  XOR U26302 ( .A(n26903), .B(n26904), .Z(n26889) );
  AND U26303 ( .A(n2249), .B(n26905), .Z(n26904) );
  IV U26304 ( .A(n26900), .Z(n26902) );
  XOR U26305 ( .A(n26906), .B(n26907), .Z(n26900) );
  AND U26306 ( .A(n2233), .B(n26899), .Z(n26907) );
  XNOR U26307 ( .A(n26897), .B(n26906), .Z(n26899) );
  XNOR U26308 ( .A(n26908), .B(n26909), .Z(n26897) );
  AND U26309 ( .A(n2237), .B(n26910), .Z(n26909) );
  XOR U26310 ( .A(p_input[1834]), .B(n26908), .Z(n26910) );
  XNOR U26311 ( .A(n26911), .B(n26912), .Z(n26908) );
  AND U26312 ( .A(n2241), .B(n26913), .Z(n26912) );
  XOR U26313 ( .A(n26914), .B(n26915), .Z(n26906) );
  AND U26314 ( .A(n2245), .B(n26905), .Z(n26915) );
  XNOR U26315 ( .A(n26916), .B(n26903), .Z(n26905) );
  XOR U26316 ( .A(n26917), .B(n26918), .Z(n26903) );
  AND U26317 ( .A(n2268), .B(n26919), .Z(n26918) );
  IV U26318 ( .A(n26914), .Z(n26916) );
  XOR U26319 ( .A(n26920), .B(n26921), .Z(n26914) );
  AND U26320 ( .A(n2252), .B(n26913), .Z(n26921) );
  XNOR U26321 ( .A(n26911), .B(n26920), .Z(n26913) );
  XNOR U26322 ( .A(n26922), .B(n26923), .Z(n26911) );
  AND U26323 ( .A(n2256), .B(n26924), .Z(n26923) );
  XOR U26324 ( .A(p_input[1850]), .B(n26922), .Z(n26924) );
  XNOR U26325 ( .A(n26925), .B(n26926), .Z(n26922) );
  AND U26326 ( .A(n2260), .B(n26927), .Z(n26926) );
  XOR U26327 ( .A(n26928), .B(n26929), .Z(n26920) );
  AND U26328 ( .A(n2264), .B(n26919), .Z(n26929) );
  XNOR U26329 ( .A(n26930), .B(n26917), .Z(n26919) );
  XOR U26330 ( .A(n26931), .B(n26932), .Z(n26917) );
  AND U26331 ( .A(n2287), .B(n26933), .Z(n26932) );
  IV U26332 ( .A(n26928), .Z(n26930) );
  XOR U26333 ( .A(n26934), .B(n26935), .Z(n26928) );
  AND U26334 ( .A(n2271), .B(n26927), .Z(n26935) );
  XNOR U26335 ( .A(n26925), .B(n26934), .Z(n26927) );
  XNOR U26336 ( .A(n26936), .B(n26937), .Z(n26925) );
  AND U26337 ( .A(n2275), .B(n26938), .Z(n26937) );
  XOR U26338 ( .A(p_input[1866]), .B(n26936), .Z(n26938) );
  XNOR U26339 ( .A(n26939), .B(n26940), .Z(n26936) );
  AND U26340 ( .A(n2279), .B(n26941), .Z(n26940) );
  XOR U26341 ( .A(n26942), .B(n26943), .Z(n26934) );
  AND U26342 ( .A(n2283), .B(n26933), .Z(n26943) );
  XNOR U26343 ( .A(n26944), .B(n26931), .Z(n26933) );
  XOR U26344 ( .A(n26945), .B(n26946), .Z(n26931) );
  AND U26345 ( .A(n2306), .B(n26947), .Z(n26946) );
  IV U26346 ( .A(n26942), .Z(n26944) );
  XOR U26347 ( .A(n26948), .B(n26949), .Z(n26942) );
  AND U26348 ( .A(n2290), .B(n26941), .Z(n26949) );
  XNOR U26349 ( .A(n26939), .B(n26948), .Z(n26941) );
  XNOR U26350 ( .A(n26950), .B(n26951), .Z(n26939) );
  AND U26351 ( .A(n2294), .B(n26952), .Z(n26951) );
  XOR U26352 ( .A(p_input[1882]), .B(n26950), .Z(n26952) );
  XNOR U26353 ( .A(n26953), .B(n26954), .Z(n26950) );
  AND U26354 ( .A(n2298), .B(n26955), .Z(n26954) );
  XOR U26355 ( .A(n26956), .B(n26957), .Z(n26948) );
  AND U26356 ( .A(n2302), .B(n26947), .Z(n26957) );
  XNOR U26357 ( .A(n26958), .B(n26945), .Z(n26947) );
  XOR U26358 ( .A(n26959), .B(n26960), .Z(n26945) );
  AND U26359 ( .A(n2325), .B(n26961), .Z(n26960) );
  IV U26360 ( .A(n26956), .Z(n26958) );
  XOR U26361 ( .A(n26962), .B(n26963), .Z(n26956) );
  AND U26362 ( .A(n2309), .B(n26955), .Z(n26963) );
  XNOR U26363 ( .A(n26953), .B(n26962), .Z(n26955) );
  XNOR U26364 ( .A(n26964), .B(n26965), .Z(n26953) );
  AND U26365 ( .A(n2313), .B(n26966), .Z(n26965) );
  XOR U26366 ( .A(p_input[1898]), .B(n26964), .Z(n26966) );
  XNOR U26367 ( .A(n26967), .B(n26968), .Z(n26964) );
  AND U26368 ( .A(n2317), .B(n26969), .Z(n26968) );
  XOR U26369 ( .A(n26970), .B(n26971), .Z(n26962) );
  AND U26370 ( .A(n2321), .B(n26961), .Z(n26971) );
  XNOR U26371 ( .A(n26972), .B(n26959), .Z(n26961) );
  XOR U26372 ( .A(n26973), .B(n26974), .Z(n26959) );
  AND U26373 ( .A(n2344), .B(n26975), .Z(n26974) );
  IV U26374 ( .A(n26970), .Z(n26972) );
  XOR U26375 ( .A(n26976), .B(n26977), .Z(n26970) );
  AND U26376 ( .A(n2328), .B(n26969), .Z(n26977) );
  XNOR U26377 ( .A(n26967), .B(n26976), .Z(n26969) );
  XNOR U26378 ( .A(n26978), .B(n26979), .Z(n26967) );
  AND U26379 ( .A(n2332), .B(n26980), .Z(n26979) );
  XOR U26380 ( .A(p_input[1914]), .B(n26978), .Z(n26980) );
  XNOR U26381 ( .A(n26981), .B(n26982), .Z(n26978) );
  AND U26382 ( .A(n2336), .B(n26983), .Z(n26982) );
  XOR U26383 ( .A(n26984), .B(n26985), .Z(n26976) );
  AND U26384 ( .A(n2340), .B(n26975), .Z(n26985) );
  XNOR U26385 ( .A(n26986), .B(n26973), .Z(n26975) );
  XOR U26386 ( .A(n26987), .B(n26988), .Z(n26973) );
  AND U26387 ( .A(n2363), .B(n26989), .Z(n26988) );
  IV U26388 ( .A(n26984), .Z(n26986) );
  XOR U26389 ( .A(n26990), .B(n26991), .Z(n26984) );
  AND U26390 ( .A(n2347), .B(n26983), .Z(n26991) );
  XNOR U26391 ( .A(n26981), .B(n26990), .Z(n26983) );
  XNOR U26392 ( .A(n26992), .B(n26993), .Z(n26981) );
  AND U26393 ( .A(n2351), .B(n26994), .Z(n26993) );
  XOR U26394 ( .A(p_input[1930]), .B(n26992), .Z(n26994) );
  XNOR U26395 ( .A(n26995), .B(n26996), .Z(n26992) );
  AND U26396 ( .A(n2355), .B(n26997), .Z(n26996) );
  XOR U26397 ( .A(n26998), .B(n26999), .Z(n26990) );
  AND U26398 ( .A(n2359), .B(n26989), .Z(n26999) );
  XNOR U26399 ( .A(n27000), .B(n26987), .Z(n26989) );
  XOR U26400 ( .A(n27001), .B(n27002), .Z(n26987) );
  AND U26401 ( .A(n2382), .B(n27003), .Z(n27002) );
  IV U26402 ( .A(n26998), .Z(n27000) );
  XOR U26403 ( .A(n27004), .B(n27005), .Z(n26998) );
  AND U26404 ( .A(n2366), .B(n26997), .Z(n27005) );
  XNOR U26405 ( .A(n26995), .B(n27004), .Z(n26997) );
  XNOR U26406 ( .A(n27006), .B(n27007), .Z(n26995) );
  AND U26407 ( .A(n2370), .B(n27008), .Z(n27007) );
  XOR U26408 ( .A(p_input[1946]), .B(n27006), .Z(n27008) );
  XNOR U26409 ( .A(n27009), .B(n27010), .Z(n27006) );
  AND U26410 ( .A(n2374), .B(n27011), .Z(n27010) );
  XOR U26411 ( .A(n27012), .B(n27013), .Z(n27004) );
  AND U26412 ( .A(n2378), .B(n27003), .Z(n27013) );
  XNOR U26413 ( .A(n27014), .B(n27001), .Z(n27003) );
  XOR U26414 ( .A(n27015), .B(n27016), .Z(n27001) );
  AND U26415 ( .A(n2401), .B(n27017), .Z(n27016) );
  IV U26416 ( .A(n27012), .Z(n27014) );
  XOR U26417 ( .A(n27018), .B(n27019), .Z(n27012) );
  AND U26418 ( .A(n2385), .B(n27011), .Z(n27019) );
  XNOR U26419 ( .A(n27009), .B(n27018), .Z(n27011) );
  XNOR U26420 ( .A(n27020), .B(n27021), .Z(n27009) );
  AND U26421 ( .A(n2389), .B(n27022), .Z(n27021) );
  XOR U26422 ( .A(p_input[1962]), .B(n27020), .Z(n27022) );
  XNOR U26423 ( .A(n27023), .B(n27024), .Z(n27020) );
  AND U26424 ( .A(n2393), .B(n27025), .Z(n27024) );
  XOR U26425 ( .A(n27026), .B(n27027), .Z(n27018) );
  AND U26426 ( .A(n2397), .B(n27017), .Z(n27027) );
  XNOR U26427 ( .A(n27028), .B(n27015), .Z(n27017) );
  XOR U26428 ( .A(n27029), .B(n27030), .Z(n27015) );
  AND U26429 ( .A(n2420), .B(n27031), .Z(n27030) );
  IV U26430 ( .A(n27026), .Z(n27028) );
  XOR U26431 ( .A(n27032), .B(n27033), .Z(n27026) );
  AND U26432 ( .A(n2404), .B(n27025), .Z(n27033) );
  XNOR U26433 ( .A(n27023), .B(n27032), .Z(n27025) );
  XNOR U26434 ( .A(n27034), .B(n27035), .Z(n27023) );
  AND U26435 ( .A(n2408), .B(n27036), .Z(n27035) );
  XOR U26436 ( .A(p_input[1978]), .B(n27034), .Z(n27036) );
  XNOR U26437 ( .A(n27037), .B(n27038), .Z(n27034) );
  AND U26438 ( .A(n2412), .B(n27039), .Z(n27038) );
  XOR U26439 ( .A(n27040), .B(n27041), .Z(n27032) );
  AND U26440 ( .A(n2416), .B(n27031), .Z(n27041) );
  XNOR U26441 ( .A(n27042), .B(n27029), .Z(n27031) );
  XOR U26442 ( .A(n27043), .B(n27044), .Z(n27029) );
  AND U26443 ( .A(n2438), .B(n27045), .Z(n27044) );
  IV U26444 ( .A(n27040), .Z(n27042) );
  XOR U26445 ( .A(n27046), .B(n27047), .Z(n27040) );
  AND U26446 ( .A(n2423), .B(n27039), .Z(n27047) );
  XNOR U26447 ( .A(n27037), .B(n27046), .Z(n27039) );
  XNOR U26448 ( .A(n27048), .B(n27049), .Z(n27037) );
  AND U26449 ( .A(n2427), .B(n27050), .Z(n27049) );
  XOR U26450 ( .A(p_input[1994]), .B(n27048), .Z(n27050) );
  XOR U26451 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n27051), 
        .Z(n27048) );
  AND U26452 ( .A(n2430), .B(n27052), .Z(n27051) );
  XOR U26453 ( .A(n27053), .B(n27054), .Z(n27046) );
  AND U26454 ( .A(n2434), .B(n27045), .Z(n27054) );
  XNOR U26455 ( .A(n27055), .B(n27043), .Z(n27045) );
  XOR U26456 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n27056), .Z(n27043) );
  AND U26457 ( .A(n2446), .B(n27057), .Z(n27056) );
  IV U26458 ( .A(n27053), .Z(n27055) );
  XOR U26459 ( .A(n27058), .B(n27059), .Z(n27053) );
  AND U26460 ( .A(n2441), .B(n27052), .Z(n27059) );
  XOR U26461 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n27058), 
        .Z(n27052) );
  XOR U26462 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n27060), 
        .Z(n27058) );
  AND U26463 ( .A(n2443), .B(n27057), .Z(n27060) );
  XOR U26464 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n27057) );
  XOR U26465 ( .A(n16517), .B(n27061), .Z(o[0]) );
  AND U26466 ( .A(n62), .B(n27062), .Z(n16517) );
  XOR U26467 ( .A(n16518), .B(n27061), .Z(n27062) );
  XOR U26468 ( .A(n27063), .B(n27064), .Z(n27061) );
  AND U26469 ( .A(n82), .B(n27065), .Z(n27064) );
  XOR U26470 ( .A(n27066), .B(n45), .Z(n16518) );
  AND U26471 ( .A(n65), .B(n27067), .Z(n45) );
  XOR U26472 ( .A(n46), .B(n27066), .Z(n27067) );
  XOR U26473 ( .A(n27068), .B(n27069), .Z(n46) );
  AND U26474 ( .A(n70), .B(n27070), .Z(n27069) );
  XOR U26475 ( .A(p_input[0]), .B(n27068), .Z(n27070) );
  XNOR U26476 ( .A(n27071), .B(n27072), .Z(n27068) );
  AND U26477 ( .A(n74), .B(n27073), .Z(n27072) );
  XOR U26478 ( .A(n27074), .B(n27075), .Z(n27066) );
  AND U26479 ( .A(n78), .B(n27065), .Z(n27075) );
  XNOR U26480 ( .A(n27076), .B(n27063), .Z(n27065) );
  XOR U26481 ( .A(n27077), .B(n27078), .Z(n27063) );
  AND U26482 ( .A(n102), .B(n27079), .Z(n27078) );
  IV U26483 ( .A(n27074), .Z(n27076) );
  XOR U26484 ( .A(n27080), .B(n27081), .Z(n27074) );
  AND U26485 ( .A(n86), .B(n27073), .Z(n27081) );
  XNOR U26486 ( .A(n27071), .B(n27080), .Z(n27073) );
  XNOR U26487 ( .A(n27082), .B(n27083), .Z(n27071) );
  AND U26488 ( .A(n90), .B(n27084), .Z(n27083) );
  XOR U26489 ( .A(p_input[16]), .B(n27082), .Z(n27084) );
  XNOR U26490 ( .A(n27085), .B(n27086), .Z(n27082) );
  AND U26491 ( .A(n94), .B(n27087), .Z(n27086) );
  XOR U26492 ( .A(n27088), .B(n27089), .Z(n27080) );
  AND U26493 ( .A(n98), .B(n27079), .Z(n27089) );
  XNOR U26494 ( .A(n27090), .B(n27077), .Z(n27079) );
  XOR U26495 ( .A(n27091), .B(n27092), .Z(n27077) );
  AND U26496 ( .A(n121), .B(n27093), .Z(n27092) );
  IV U26497 ( .A(n27088), .Z(n27090) );
  XOR U26498 ( .A(n27094), .B(n27095), .Z(n27088) );
  AND U26499 ( .A(n105), .B(n27087), .Z(n27095) );
  XNOR U26500 ( .A(n27085), .B(n27094), .Z(n27087) );
  XNOR U26501 ( .A(n27096), .B(n27097), .Z(n27085) );
  AND U26502 ( .A(n109), .B(n27098), .Z(n27097) );
  XOR U26503 ( .A(p_input[32]), .B(n27096), .Z(n27098) );
  XNOR U26504 ( .A(n27099), .B(n27100), .Z(n27096) );
  AND U26505 ( .A(n113), .B(n27101), .Z(n27100) );
  XOR U26506 ( .A(n27102), .B(n27103), .Z(n27094) );
  AND U26507 ( .A(n117), .B(n27093), .Z(n27103) );
  XNOR U26508 ( .A(n27104), .B(n27091), .Z(n27093) );
  XOR U26509 ( .A(n27105), .B(n27106), .Z(n27091) );
  AND U26510 ( .A(n140), .B(n27107), .Z(n27106) );
  IV U26511 ( .A(n27102), .Z(n27104) );
  XOR U26512 ( .A(n27108), .B(n27109), .Z(n27102) );
  AND U26513 ( .A(n124), .B(n27101), .Z(n27109) );
  XNOR U26514 ( .A(n27099), .B(n27108), .Z(n27101) );
  XNOR U26515 ( .A(n27110), .B(n27111), .Z(n27099) );
  AND U26516 ( .A(n128), .B(n27112), .Z(n27111) );
  XOR U26517 ( .A(p_input[48]), .B(n27110), .Z(n27112) );
  XNOR U26518 ( .A(n27113), .B(n27114), .Z(n27110) );
  AND U26519 ( .A(n132), .B(n27115), .Z(n27114) );
  XOR U26520 ( .A(n27116), .B(n27117), .Z(n27108) );
  AND U26521 ( .A(n136), .B(n27107), .Z(n27117) );
  XNOR U26522 ( .A(n27118), .B(n27105), .Z(n27107) );
  XOR U26523 ( .A(n27119), .B(n27120), .Z(n27105) );
  AND U26524 ( .A(n159), .B(n27121), .Z(n27120) );
  IV U26525 ( .A(n27116), .Z(n27118) );
  XOR U26526 ( .A(n27122), .B(n27123), .Z(n27116) );
  AND U26527 ( .A(n143), .B(n27115), .Z(n27123) );
  XNOR U26528 ( .A(n27113), .B(n27122), .Z(n27115) );
  XNOR U26529 ( .A(n27124), .B(n27125), .Z(n27113) );
  AND U26530 ( .A(n147), .B(n27126), .Z(n27125) );
  XOR U26531 ( .A(p_input[64]), .B(n27124), .Z(n27126) );
  XNOR U26532 ( .A(n27127), .B(n27128), .Z(n27124) );
  AND U26533 ( .A(n151), .B(n27129), .Z(n27128) );
  XOR U26534 ( .A(n27130), .B(n27131), .Z(n27122) );
  AND U26535 ( .A(n155), .B(n27121), .Z(n27131) );
  XNOR U26536 ( .A(n27132), .B(n27119), .Z(n27121) );
  XOR U26537 ( .A(n27133), .B(n27134), .Z(n27119) );
  AND U26538 ( .A(n178), .B(n27135), .Z(n27134) );
  IV U26539 ( .A(n27130), .Z(n27132) );
  XOR U26540 ( .A(n27136), .B(n27137), .Z(n27130) );
  AND U26541 ( .A(n162), .B(n27129), .Z(n27137) );
  XNOR U26542 ( .A(n27127), .B(n27136), .Z(n27129) );
  XNOR U26543 ( .A(n27138), .B(n27139), .Z(n27127) );
  AND U26544 ( .A(n166), .B(n27140), .Z(n27139) );
  XOR U26545 ( .A(p_input[80]), .B(n27138), .Z(n27140) );
  XNOR U26546 ( .A(n27141), .B(n27142), .Z(n27138) );
  AND U26547 ( .A(n170), .B(n27143), .Z(n27142) );
  XOR U26548 ( .A(n27144), .B(n27145), .Z(n27136) );
  AND U26549 ( .A(n174), .B(n27135), .Z(n27145) );
  XNOR U26550 ( .A(n27146), .B(n27133), .Z(n27135) );
  XOR U26551 ( .A(n27147), .B(n27148), .Z(n27133) );
  AND U26552 ( .A(n197), .B(n27149), .Z(n27148) );
  IV U26553 ( .A(n27144), .Z(n27146) );
  XOR U26554 ( .A(n27150), .B(n27151), .Z(n27144) );
  AND U26555 ( .A(n181), .B(n27143), .Z(n27151) );
  XNOR U26556 ( .A(n27141), .B(n27150), .Z(n27143) );
  XNOR U26557 ( .A(n27152), .B(n27153), .Z(n27141) );
  AND U26558 ( .A(n185), .B(n27154), .Z(n27153) );
  XOR U26559 ( .A(p_input[96]), .B(n27152), .Z(n27154) );
  XNOR U26560 ( .A(n27155), .B(n27156), .Z(n27152) );
  AND U26561 ( .A(n189), .B(n27157), .Z(n27156) );
  XOR U26562 ( .A(n27158), .B(n27159), .Z(n27150) );
  AND U26563 ( .A(n193), .B(n27149), .Z(n27159) );
  XNOR U26564 ( .A(n27160), .B(n27147), .Z(n27149) );
  XOR U26565 ( .A(n27161), .B(n27162), .Z(n27147) );
  AND U26566 ( .A(n216), .B(n27163), .Z(n27162) );
  IV U26567 ( .A(n27158), .Z(n27160) );
  XOR U26568 ( .A(n27164), .B(n27165), .Z(n27158) );
  AND U26569 ( .A(n200), .B(n27157), .Z(n27165) );
  XNOR U26570 ( .A(n27155), .B(n27164), .Z(n27157) );
  XNOR U26571 ( .A(n27166), .B(n27167), .Z(n27155) );
  AND U26572 ( .A(n204), .B(n27168), .Z(n27167) );
  XOR U26573 ( .A(p_input[112]), .B(n27166), .Z(n27168) );
  XNOR U26574 ( .A(n27169), .B(n27170), .Z(n27166) );
  AND U26575 ( .A(n208), .B(n27171), .Z(n27170) );
  XOR U26576 ( .A(n27172), .B(n27173), .Z(n27164) );
  AND U26577 ( .A(n212), .B(n27163), .Z(n27173) );
  XNOR U26578 ( .A(n27174), .B(n27161), .Z(n27163) );
  XOR U26579 ( .A(n27175), .B(n27176), .Z(n27161) );
  AND U26580 ( .A(n235), .B(n27177), .Z(n27176) );
  IV U26581 ( .A(n27172), .Z(n27174) );
  XOR U26582 ( .A(n27178), .B(n27179), .Z(n27172) );
  AND U26583 ( .A(n219), .B(n27171), .Z(n27179) );
  XNOR U26584 ( .A(n27169), .B(n27178), .Z(n27171) );
  XNOR U26585 ( .A(n27180), .B(n27181), .Z(n27169) );
  AND U26586 ( .A(n223), .B(n27182), .Z(n27181) );
  XOR U26587 ( .A(p_input[128]), .B(n27180), .Z(n27182) );
  XNOR U26588 ( .A(n27183), .B(n27184), .Z(n27180) );
  AND U26589 ( .A(n227), .B(n27185), .Z(n27184) );
  XOR U26590 ( .A(n27186), .B(n27187), .Z(n27178) );
  AND U26591 ( .A(n231), .B(n27177), .Z(n27187) );
  XNOR U26592 ( .A(n27188), .B(n27175), .Z(n27177) );
  XOR U26593 ( .A(n27189), .B(n27190), .Z(n27175) );
  AND U26594 ( .A(n254), .B(n27191), .Z(n27190) );
  IV U26595 ( .A(n27186), .Z(n27188) );
  XOR U26596 ( .A(n27192), .B(n27193), .Z(n27186) );
  AND U26597 ( .A(n238), .B(n27185), .Z(n27193) );
  XNOR U26598 ( .A(n27183), .B(n27192), .Z(n27185) );
  XNOR U26599 ( .A(n27194), .B(n27195), .Z(n27183) );
  AND U26600 ( .A(n242), .B(n27196), .Z(n27195) );
  XOR U26601 ( .A(p_input[144]), .B(n27194), .Z(n27196) );
  XNOR U26602 ( .A(n27197), .B(n27198), .Z(n27194) );
  AND U26603 ( .A(n246), .B(n27199), .Z(n27198) );
  XOR U26604 ( .A(n27200), .B(n27201), .Z(n27192) );
  AND U26605 ( .A(n250), .B(n27191), .Z(n27201) );
  XNOR U26606 ( .A(n27202), .B(n27189), .Z(n27191) );
  XOR U26607 ( .A(n27203), .B(n27204), .Z(n27189) );
  AND U26608 ( .A(n273), .B(n27205), .Z(n27204) );
  IV U26609 ( .A(n27200), .Z(n27202) );
  XOR U26610 ( .A(n27206), .B(n27207), .Z(n27200) );
  AND U26611 ( .A(n257), .B(n27199), .Z(n27207) );
  XNOR U26612 ( .A(n27197), .B(n27206), .Z(n27199) );
  XNOR U26613 ( .A(n27208), .B(n27209), .Z(n27197) );
  AND U26614 ( .A(n261), .B(n27210), .Z(n27209) );
  XOR U26615 ( .A(p_input[160]), .B(n27208), .Z(n27210) );
  XNOR U26616 ( .A(n27211), .B(n27212), .Z(n27208) );
  AND U26617 ( .A(n265), .B(n27213), .Z(n27212) );
  XOR U26618 ( .A(n27214), .B(n27215), .Z(n27206) );
  AND U26619 ( .A(n269), .B(n27205), .Z(n27215) );
  XNOR U26620 ( .A(n27216), .B(n27203), .Z(n27205) );
  XOR U26621 ( .A(n27217), .B(n27218), .Z(n27203) );
  AND U26622 ( .A(n292), .B(n27219), .Z(n27218) );
  IV U26623 ( .A(n27214), .Z(n27216) );
  XOR U26624 ( .A(n27220), .B(n27221), .Z(n27214) );
  AND U26625 ( .A(n276), .B(n27213), .Z(n27221) );
  XNOR U26626 ( .A(n27211), .B(n27220), .Z(n27213) );
  XNOR U26627 ( .A(n27222), .B(n27223), .Z(n27211) );
  AND U26628 ( .A(n280), .B(n27224), .Z(n27223) );
  XOR U26629 ( .A(p_input[176]), .B(n27222), .Z(n27224) );
  XNOR U26630 ( .A(n27225), .B(n27226), .Z(n27222) );
  AND U26631 ( .A(n284), .B(n27227), .Z(n27226) );
  XOR U26632 ( .A(n27228), .B(n27229), .Z(n27220) );
  AND U26633 ( .A(n288), .B(n27219), .Z(n27229) );
  XNOR U26634 ( .A(n27230), .B(n27217), .Z(n27219) );
  XOR U26635 ( .A(n27231), .B(n27232), .Z(n27217) );
  AND U26636 ( .A(n311), .B(n27233), .Z(n27232) );
  IV U26637 ( .A(n27228), .Z(n27230) );
  XOR U26638 ( .A(n27234), .B(n27235), .Z(n27228) );
  AND U26639 ( .A(n295), .B(n27227), .Z(n27235) );
  XNOR U26640 ( .A(n27225), .B(n27234), .Z(n27227) );
  XNOR U26641 ( .A(n27236), .B(n27237), .Z(n27225) );
  AND U26642 ( .A(n299), .B(n27238), .Z(n27237) );
  XOR U26643 ( .A(p_input[192]), .B(n27236), .Z(n27238) );
  XNOR U26644 ( .A(n27239), .B(n27240), .Z(n27236) );
  AND U26645 ( .A(n303), .B(n27241), .Z(n27240) );
  XOR U26646 ( .A(n27242), .B(n27243), .Z(n27234) );
  AND U26647 ( .A(n307), .B(n27233), .Z(n27243) );
  XNOR U26648 ( .A(n27244), .B(n27231), .Z(n27233) );
  XOR U26649 ( .A(n27245), .B(n27246), .Z(n27231) );
  AND U26650 ( .A(n330), .B(n27247), .Z(n27246) );
  IV U26651 ( .A(n27242), .Z(n27244) );
  XOR U26652 ( .A(n27248), .B(n27249), .Z(n27242) );
  AND U26653 ( .A(n314), .B(n27241), .Z(n27249) );
  XNOR U26654 ( .A(n27239), .B(n27248), .Z(n27241) );
  XNOR U26655 ( .A(n27250), .B(n27251), .Z(n27239) );
  AND U26656 ( .A(n318), .B(n27252), .Z(n27251) );
  XOR U26657 ( .A(p_input[208]), .B(n27250), .Z(n27252) );
  XNOR U26658 ( .A(n27253), .B(n27254), .Z(n27250) );
  AND U26659 ( .A(n322), .B(n27255), .Z(n27254) );
  XOR U26660 ( .A(n27256), .B(n27257), .Z(n27248) );
  AND U26661 ( .A(n326), .B(n27247), .Z(n27257) );
  XNOR U26662 ( .A(n27258), .B(n27245), .Z(n27247) );
  XOR U26663 ( .A(n27259), .B(n27260), .Z(n27245) );
  AND U26664 ( .A(n349), .B(n27261), .Z(n27260) );
  IV U26665 ( .A(n27256), .Z(n27258) );
  XOR U26666 ( .A(n27262), .B(n27263), .Z(n27256) );
  AND U26667 ( .A(n333), .B(n27255), .Z(n27263) );
  XNOR U26668 ( .A(n27253), .B(n27262), .Z(n27255) );
  XNOR U26669 ( .A(n27264), .B(n27265), .Z(n27253) );
  AND U26670 ( .A(n337), .B(n27266), .Z(n27265) );
  XOR U26671 ( .A(p_input[224]), .B(n27264), .Z(n27266) );
  XNOR U26672 ( .A(n27267), .B(n27268), .Z(n27264) );
  AND U26673 ( .A(n341), .B(n27269), .Z(n27268) );
  XOR U26674 ( .A(n27270), .B(n27271), .Z(n27262) );
  AND U26675 ( .A(n345), .B(n27261), .Z(n27271) );
  XNOR U26676 ( .A(n27272), .B(n27259), .Z(n27261) );
  XOR U26677 ( .A(n27273), .B(n27274), .Z(n27259) );
  AND U26678 ( .A(n368), .B(n27275), .Z(n27274) );
  IV U26679 ( .A(n27270), .Z(n27272) );
  XOR U26680 ( .A(n27276), .B(n27277), .Z(n27270) );
  AND U26681 ( .A(n352), .B(n27269), .Z(n27277) );
  XNOR U26682 ( .A(n27267), .B(n27276), .Z(n27269) );
  XNOR U26683 ( .A(n27278), .B(n27279), .Z(n27267) );
  AND U26684 ( .A(n356), .B(n27280), .Z(n27279) );
  XOR U26685 ( .A(p_input[240]), .B(n27278), .Z(n27280) );
  XNOR U26686 ( .A(n27281), .B(n27282), .Z(n27278) );
  AND U26687 ( .A(n360), .B(n27283), .Z(n27282) );
  XOR U26688 ( .A(n27284), .B(n27285), .Z(n27276) );
  AND U26689 ( .A(n364), .B(n27275), .Z(n27285) );
  XNOR U26690 ( .A(n27286), .B(n27273), .Z(n27275) );
  XOR U26691 ( .A(n27287), .B(n27288), .Z(n27273) );
  AND U26692 ( .A(n387), .B(n27289), .Z(n27288) );
  IV U26693 ( .A(n27284), .Z(n27286) );
  XOR U26694 ( .A(n27290), .B(n27291), .Z(n27284) );
  AND U26695 ( .A(n371), .B(n27283), .Z(n27291) );
  XNOR U26696 ( .A(n27281), .B(n27290), .Z(n27283) );
  XNOR U26697 ( .A(n27292), .B(n27293), .Z(n27281) );
  AND U26698 ( .A(n375), .B(n27294), .Z(n27293) );
  XOR U26699 ( .A(p_input[256]), .B(n27292), .Z(n27294) );
  XNOR U26700 ( .A(n27295), .B(n27296), .Z(n27292) );
  AND U26701 ( .A(n379), .B(n27297), .Z(n27296) );
  XOR U26702 ( .A(n27298), .B(n27299), .Z(n27290) );
  AND U26703 ( .A(n383), .B(n27289), .Z(n27299) );
  XNOR U26704 ( .A(n27300), .B(n27287), .Z(n27289) );
  XOR U26705 ( .A(n27301), .B(n27302), .Z(n27287) );
  AND U26706 ( .A(n406), .B(n27303), .Z(n27302) );
  IV U26707 ( .A(n27298), .Z(n27300) );
  XOR U26708 ( .A(n27304), .B(n27305), .Z(n27298) );
  AND U26709 ( .A(n390), .B(n27297), .Z(n27305) );
  XNOR U26710 ( .A(n27295), .B(n27304), .Z(n27297) );
  XNOR U26711 ( .A(n27306), .B(n27307), .Z(n27295) );
  AND U26712 ( .A(n394), .B(n27308), .Z(n27307) );
  XOR U26713 ( .A(p_input[272]), .B(n27306), .Z(n27308) );
  XNOR U26714 ( .A(n27309), .B(n27310), .Z(n27306) );
  AND U26715 ( .A(n398), .B(n27311), .Z(n27310) );
  XOR U26716 ( .A(n27312), .B(n27313), .Z(n27304) );
  AND U26717 ( .A(n402), .B(n27303), .Z(n27313) );
  XNOR U26718 ( .A(n27314), .B(n27301), .Z(n27303) );
  XOR U26719 ( .A(n27315), .B(n27316), .Z(n27301) );
  AND U26720 ( .A(n425), .B(n27317), .Z(n27316) );
  IV U26721 ( .A(n27312), .Z(n27314) );
  XOR U26722 ( .A(n27318), .B(n27319), .Z(n27312) );
  AND U26723 ( .A(n409), .B(n27311), .Z(n27319) );
  XNOR U26724 ( .A(n27309), .B(n27318), .Z(n27311) );
  XNOR U26725 ( .A(n27320), .B(n27321), .Z(n27309) );
  AND U26726 ( .A(n413), .B(n27322), .Z(n27321) );
  XOR U26727 ( .A(p_input[288]), .B(n27320), .Z(n27322) );
  XNOR U26728 ( .A(n27323), .B(n27324), .Z(n27320) );
  AND U26729 ( .A(n417), .B(n27325), .Z(n27324) );
  XOR U26730 ( .A(n27326), .B(n27327), .Z(n27318) );
  AND U26731 ( .A(n421), .B(n27317), .Z(n27327) );
  XNOR U26732 ( .A(n27328), .B(n27315), .Z(n27317) );
  XOR U26733 ( .A(n27329), .B(n27330), .Z(n27315) );
  AND U26734 ( .A(n444), .B(n27331), .Z(n27330) );
  IV U26735 ( .A(n27326), .Z(n27328) );
  XOR U26736 ( .A(n27332), .B(n27333), .Z(n27326) );
  AND U26737 ( .A(n428), .B(n27325), .Z(n27333) );
  XNOR U26738 ( .A(n27323), .B(n27332), .Z(n27325) );
  XNOR U26739 ( .A(n27334), .B(n27335), .Z(n27323) );
  AND U26740 ( .A(n432), .B(n27336), .Z(n27335) );
  XOR U26741 ( .A(p_input[304]), .B(n27334), .Z(n27336) );
  XNOR U26742 ( .A(n27337), .B(n27338), .Z(n27334) );
  AND U26743 ( .A(n436), .B(n27339), .Z(n27338) );
  XOR U26744 ( .A(n27340), .B(n27341), .Z(n27332) );
  AND U26745 ( .A(n440), .B(n27331), .Z(n27341) );
  XNOR U26746 ( .A(n27342), .B(n27329), .Z(n27331) );
  XOR U26747 ( .A(n27343), .B(n27344), .Z(n27329) );
  AND U26748 ( .A(n463), .B(n27345), .Z(n27344) );
  IV U26749 ( .A(n27340), .Z(n27342) );
  XOR U26750 ( .A(n27346), .B(n27347), .Z(n27340) );
  AND U26751 ( .A(n447), .B(n27339), .Z(n27347) );
  XNOR U26752 ( .A(n27337), .B(n27346), .Z(n27339) );
  XNOR U26753 ( .A(n27348), .B(n27349), .Z(n27337) );
  AND U26754 ( .A(n451), .B(n27350), .Z(n27349) );
  XOR U26755 ( .A(p_input[320]), .B(n27348), .Z(n27350) );
  XNOR U26756 ( .A(n27351), .B(n27352), .Z(n27348) );
  AND U26757 ( .A(n455), .B(n27353), .Z(n27352) );
  XOR U26758 ( .A(n27354), .B(n27355), .Z(n27346) );
  AND U26759 ( .A(n459), .B(n27345), .Z(n27355) );
  XNOR U26760 ( .A(n27356), .B(n27343), .Z(n27345) );
  XOR U26761 ( .A(n27357), .B(n27358), .Z(n27343) );
  AND U26762 ( .A(n482), .B(n27359), .Z(n27358) );
  IV U26763 ( .A(n27354), .Z(n27356) );
  XOR U26764 ( .A(n27360), .B(n27361), .Z(n27354) );
  AND U26765 ( .A(n466), .B(n27353), .Z(n27361) );
  XNOR U26766 ( .A(n27351), .B(n27360), .Z(n27353) );
  XNOR U26767 ( .A(n27362), .B(n27363), .Z(n27351) );
  AND U26768 ( .A(n470), .B(n27364), .Z(n27363) );
  XOR U26769 ( .A(p_input[336]), .B(n27362), .Z(n27364) );
  XNOR U26770 ( .A(n27365), .B(n27366), .Z(n27362) );
  AND U26771 ( .A(n474), .B(n27367), .Z(n27366) );
  XOR U26772 ( .A(n27368), .B(n27369), .Z(n27360) );
  AND U26773 ( .A(n478), .B(n27359), .Z(n27369) );
  XNOR U26774 ( .A(n27370), .B(n27357), .Z(n27359) );
  XOR U26775 ( .A(n27371), .B(n27372), .Z(n27357) );
  AND U26776 ( .A(n501), .B(n27373), .Z(n27372) );
  IV U26777 ( .A(n27368), .Z(n27370) );
  XOR U26778 ( .A(n27374), .B(n27375), .Z(n27368) );
  AND U26779 ( .A(n485), .B(n27367), .Z(n27375) );
  XNOR U26780 ( .A(n27365), .B(n27374), .Z(n27367) );
  XNOR U26781 ( .A(n27376), .B(n27377), .Z(n27365) );
  AND U26782 ( .A(n489), .B(n27378), .Z(n27377) );
  XOR U26783 ( .A(p_input[352]), .B(n27376), .Z(n27378) );
  XNOR U26784 ( .A(n27379), .B(n27380), .Z(n27376) );
  AND U26785 ( .A(n493), .B(n27381), .Z(n27380) );
  XOR U26786 ( .A(n27382), .B(n27383), .Z(n27374) );
  AND U26787 ( .A(n497), .B(n27373), .Z(n27383) );
  XNOR U26788 ( .A(n27384), .B(n27371), .Z(n27373) );
  XOR U26789 ( .A(n27385), .B(n27386), .Z(n27371) );
  AND U26790 ( .A(n520), .B(n27387), .Z(n27386) );
  IV U26791 ( .A(n27382), .Z(n27384) );
  XOR U26792 ( .A(n27388), .B(n27389), .Z(n27382) );
  AND U26793 ( .A(n504), .B(n27381), .Z(n27389) );
  XNOR U26794 ( .A(n27379), .B(n27388), .Z(n27381) );
  XNOR U26795 ( .A(n27390), .B(n27391), .Z(n27379) );
  AND U26796 ( .A(n508), .B(n27392), .Z(n27391) );
  XOR U26797 ( .A(p_input[368]), .B(n27390), .Z(n27392) );
  XNOR U26798 ( .A(n27393), .B(n27394), .Z(n27390) );
  AND U26799 ( .A(n512), .B(n27395), .Z(n27394) );
  XOR U26800 ( .A(n27396), .B(n27397), .Z(n27388) );
  AND U26801 ( .A(n516), .B(n27387), .Z(n27397) );
  XNOR U26802 ( .A(n27398), .B(n27385), .Z(n27387) );
  XOR U26803 ( .A(n27399), .B(n27400), .Z(n27385) );
  AND U26804 ( .A(n539), .B(n27401), .Z(n27400) );
  IV U26805 ( .A(n27396), .Z(n27398) );
  XOR U26806 ( .A(n27402), .B(n27403), .Z(n27396) );
  AND U26807 ( .A(n523), .B(n27395), .Z(n27403) );
  XNOR U26808 ( .A(n27393), .B(n27402), .Z(n27395) );
  XNOR U26809 ( .A(n27404), .B(n27405), .Z(n27393) );
  AND U26810 ( .A(n527), .B(n27406), .Z(n27405) );
  XOR U26811 ( .A(p_input[384]), .B(n27404), .Z(n27406) );
  XNOR U26812 ( .A(n27407), .B(n27408), .Z(n27404) );
  AND U26813 ( .A(n531), .B(n27409), .Z(n27408) );
  XOR U26814 ( .A(n27410), .B(n27411), .Z(n27402) );
  AND U26815 ( .A(n535), .B(n27401), .Z(n27411) );
  XNOR U26816 ( .A(n27412), .B(n27399), .Z(n27401) );
  XOR U26817 ( .A(n27413), .B(n27414), .Z(n27399) );
  AND U26818 ( .A(n558), .B(n27415), .Z(n27414) );
  IV U26819 ( .A(n27410), .Z(n27412) );
  XOR U26820 ( .A(n27416), .B(n27417), .Z(n27410) );
  AND U26821 ( .A(n542), .B(n27409), .Z(n27417) );
  XNOR U26822 ( .A(n27407), .B(n27416), .Z(n27409) );
  XNOR U26823 ( .A(n27418), .B(n27419), .Z(n27407) );
  AND U26824 ( .A(n546), .B(n27420), .Z(n27419) );
  XOR U26825 ( .A(p_input[400]), .B(n27418), .Z(n27420) );
  XNOR U26826 ( .A(n27421), .B(n27422), .Z(n27418) );
  AND U26827 ( .A(n550), .B(n27423), .Z(n27422) );
  XOR U26828 ( .A(n27424), .B(n27425), .Z(n27416) );
  AND U26829 ( .A(n554), .B(n27415), .Z(n27425) );
  XNOR U26830 ( .A(n27426), .B(n27413), .Z(n27415) );
  XOR U26831 ( .A(n27427), .B(n27428), .Z(n27413) );
  AND U26832 ( .A(n577), .B(n27429), .Z(n27428) );
  IV U26833 ( .A(n27424), .Z(n27426) );
  XOR U26834 ( .A(n27430), .B(n27431), .Z(n27424) );
  AND U26835 ( .A(n561), .B(n27423), .Z(n27431) );
  XNOR U26836 ( .A(n27421), .B(n27430), .Z(n27423) );
  XNOR U26837 ( .A(n27432), .B(n27433), .Z(n27421) );
  AND U26838 ( .A(n565), .B(n27434), .Z(n27433) );
  XOR U26839 ( .A(p_input[416]), .B(n27432), .Z(n27434) );
  XNOR U26840 ( .A(n27435), .B(n27436), .Z(n27432) );
  AND U26841 ( .A(n569), .B(n27437), .Z(n27436) );
  XOR U26842 ( .A(n27438), .B(n27439), .Z(n27430) );
  AND U26843 ( .A(n573), .B(n27429), .Z(n27439) );
  XNOR U26844 ( .A(n27440), .B(n27427), .Z(n27429) );
  XOR U26845 ( .A(n27441), .B(n27442), .Z(n27427) );
  AND U26846 ( .A(n596), .B(n27443), .Z(n27442) );
  IV U26847 ( .A(n27438), .Z(n27440) );
  XOR U26848 ( .A(n27444), .B(n27445), .Z(n27438) );
  AND U26849 ( .A(n580), .B(n27437), .Z(n27445) );
  XNOR U26850 ( .A(n27435), .B(n27444), .Z(n27437) );
  XNOR U26851 ( .A(n27446), .B(n27447), .Z(n27435) );
  AND U26852 ( .A(n584), .B(n27448), .Z(n27447) );
  XOR U26853 ( .A(p_input[432]), .B(n27446), .Z(n27448) );
  XNOR U26854 ( .A(n27449), .B(n27450), .Z(n27446) );
  AND U26855 ( .A(n588), .B(n27451), .Z(n27450) );
  XOR U26856 ( .A(n27452), .B(n27453), .Z(n27444) );
  AND U26857 ( .A(n592), .B(n27443), .Z(n27453) );
  XNOR U26858 ( .A(n27454), .B(n27441), .Z(n27443) );
  XOR U26859 ( .A(n27455), .B(n27456), .Z(n27441) );
  AND U26860 ( .A(n615), .B(n27457), .Z(n27456) );
  IV U26861 ( .A(n27452), .Z(n27454) );
  XOR U26862 ( .A(n27458), .B(n27459), .Z(n27452) );
  AND U26863 ( .A(n599), .B(n27451), .Z(n27459) );
  XNOR U26864 ( .A(n27449), .B(n27458), .Z(n27451) );
  XNOR U26865 ( .A(n27460), .B(n27461), .Z(n27449) );
  AND U26866 ( .A(n603), .B(n27462), .Z(n27461) );
  XOR U26867 ( .A(p_input[448]), .B(n27460), .Z(n27462) );
  XNOR U26868 ( .A(n27463), .B(n27464), .Z(n27460) );
  AND U26869 ( .A(n607), .B(n27465), .Z(n27464) );
  XOR U26870 ( .A(n27466), .B(n27467), .Z(n27458) );
  AND U26871 ( .A(n611), .B(n27457), .Z(n27467) );
  XNOR U26872 ( .A(n27468), .B(n27455), .Z(n27457) );
  XOR U26873 ( .A(n27469), .B(n27470), .Z(n27455) );
  AND U26874 ( .A(n634), .B(n27471), .Z(n27470) );
  IV U26875 ( .A(n27466), .Z(n27468) );
  XOR U26876 ( .A(n27472), .B(n27473), .Z(n27466) );
  AND U26877 ( .A(n618), .B(n27465), .Z(n27473) );
  XNOR U26878 ( .A(n27463), .B(n27472), .Z(n27465) );
  XNOR U26879 ( .A(n27474), .B(n27475), .Z(n27463) );
  AND U26880 ( .A(n622), .B(n27476), .Z(n27475) );
  XOR U26881 ( .A(p_input[464]), .B(n27474), .Z(n27476) );
  XNOR U26882 ( .A(n27477), .B(n27478), .Z(n27474) );
  AND U26883 ( .A(n626), .B(n27479), .Z(n27478) );
  XOR U26884 ( .A(n27480), .B(n27481), .Z(n27472) );
  AND U26885 ( .A(n630), .B(n27471), .Z(n27481) );
  XNOR U26886 ( .A(n27482), .B(n27469), .Z(n27471) );
  XOR U26887 ( .A(n27483), .B(n27484), .Z(n27469) );
  AND U26888 ( .A(n653), .B(n27485), .Z(n27484) );
  IV U26889 ( .A(n27480), .Z(n27482) );
  XOR U26890 ( .A(n27486), .B(n27487), .Z(n27480) );
  AND U26891 ( .A(n637), .B(n27479), .Z(n27487) );
  XNOR U26892 ( .A(n27477), .B(n27486), .Z(n27479) );
  XNOR U26893 ( .A(n27488), .B(n27489), .Z(n27477) );
  AND U26894 ( .A(n641), .B(n27490), .Z(n27489) );
  XOR U26895 ( .A(p_input[480]), .B(n27488), .Z(n27490) );
  XNOR U26896 ( .A(n27491), .B(n27492), .Z(n27488) );
  AND U26897 ( .A(n645), .B(n27493), .Z(n27492) );
  XOR U26898 ( .A(n27494), .B(n27495), .Z(n27486) );
  AND U26899 ( .A(n649), .B(n27485), .Z(n27495) );
  XNOR U26900 ( .A(n27496), .B(n27483), .Z(n27485) );
  XOR U26901 ( .A(n27497), .B(n27498), .Z(n27483) );
  AND U26902 ( .A(n672), .B(n27499), .Z(n27498) );
  IV U26903 ( .A(n27494), .Z(n27496) );
  XOR U26904 ( .A(n27500), .B(n27501), .Z(n27494) );
  AND U26905 ( .A(n656), .B(n27493), .Z(n27501) );
  XNOR U26906 ( .A(n27491), .B(n27500), .Z(n27493) );
  XNOR U26907 ( .A(n27502), .B(n27503), .Z(n27491) );
  AND U26908 ( .A(n660), .B(n27504), .Z(n27503) );
  XOR U26909 ( .A(p_input[496]), .B(n27502), .Z(n27504) );
  XNOR U26910 ( .A(n27505), .B(n27506), .Z(n27502) );
  AND U26911 ( .A(n664), .B(n27507), .Z(n27506) );
  XOR U26912 ( .A(n27508), .B(n27509), .Z(n27500) );
  AND U26913 ( .A(n668), .B(n27499), .Z(n27509) );
  XNOR U26914 ( .A(n27510), .B(n27497), .Z(n27499) );
  XOR U26915 ( .A(n27511), .B(n27512), .Z(n27497) );
  AND U26916 ( .A(n691), .B(n27513), .Z(n27512) );
  IV U26917 ( .A(n27508), .Z(n27510) );
  XOR U26918 ( .A(n27514), .B(n27515), .Z(n27508) );
  AND U26919 ( .A(n675), .B(n27507), .Z(n27515) );
  XNOR U26920 ( .A(n27505), .B(n27514), .Z(n27507) );
  XNOR U26921 ( .A(n27516), .B(n27517), .Z(n27505) );
  AND U26922 ( .A(n679), .B(n27518), .Z(n27517) );
  XOR U26923 ( .A(p_input[512]), .B(n27516), .Z(n27518) );
  XNOR U26924 ( .A(n27519), .B(n27520), .Z(n27516) );
  AND U26925 ( .A(n683), .B(n27521), .Z(n27520) );
  XOR U26926 ( .A(n27522), .B(n27523), .Z(n27514) );
  AND U26927 ( .A(n687), .B(n27513), .Z(n27523) );
  XNOR U26928 ( .A(n27524), .B(n27511), .Z(n27513) );
  XOR U26929 ( .A(n27525), .B(n27526), .Z(n27511) );
  AND U26930 ( .A(n710), .B(n27527), .Z(n27526) );
  IV U26931 ( .A(n27522), .Z(n27524) );
  XOR U26932 ( .A(n27528), .B(n27529), .Z(n27522) );
  AND U26933 ( .A(n694), .B(n27521), .Z(n27529) );
  XNOR U26934 ( .A(n27519), .B(n27528), .Z(n27521) );
  XNOR U26935 ( .A(n27530), .B(n27531), .Z(n27519) );
  AND U26936 ( .A(n698), .B(n27532), .Z(n27531) );
  XOR U26937 ( .A(p_input[528]), .B(n27530), .Z(n27532) );
  XNOR U26938 ( .A(n27533), .B(n27534), .Z(n27530) );
  AND U26939 ( .A(n702), .B(n27535), .Z(n27534) );
  XOR U26940 ( .A(n27536), .B(n27537), .Z(n27528) );
  AND U26941 ( .A(n706), .B(n27527), .Z(n27537) );
  XNOR U26942 ( .A(n27538), .B(n27525), .Z(n27527) );
  XOR U26943 ( .A(n27539), .B(n27540), .Z(n27525) );
  AND U26944 ( .A(n729), .B(n27541), .Z(n27540) );
  IV U26945 ( .A(n27536), .Z(n27538) );
  XOR U26946 ( .A(n27542), .B(n27543), .Z(n27536) );
  AND U26947 ( .A(n713), .B(n27535), .Z(n27543) );
  XNOR U26948 ( .A(n27533), .B(n27542), .Z(n27535) );
  XNOR U26949 ( .A(n27544), .B(n27545), .Z(n27533) );
  AND U26950 ( .A(n717), .B(n27546), .Z(n27545) );
  XOR U26951 ( .A(p_input[544]), .B(n27544), .Z(n27546) );
  XNOR U26952 ( .A(n27547), .B(n27548), .Z(n27544) );
  AND U26953 ( .A(n721), .B(n27549), .Z(n27548) );
  XOR U26954 ( .A(n27550), .B(n27551), .Z(n27542) );
  AND U26955 ( .A(n725), .B(n27541), .Z(n27551) );
  XNOR U26956 ( .A(n27552), .B(n27539), .Z(n27541) );
  XOR U26957 ( .A(n27553), .B(n27554), .Z(n27539) );
  AND U26958 ( .A(n748), .B(n27555), .Z(n27554) );
  IV U26959 ( .A(n27550), .Z(n27552) );
  XOR U26960 ( .A(n27556), .B(n27557), .Z(n27550) );
  AND U26961 ( .A(n732), .B(n27549), .Z(n27557) );
  XNOR U26962 ( .A(n27547), .B(n27556), .Z(n27549) );
  XNOR U26963 ( .A(n27558), .B(n27559), .Z(n27547) );
  AND U26964 ( .A(n736), .B(n27560), .Z(n27559) );
  XOR U26965 ( .A(p_input[560]), .B(n27558), .Z(n27560) );
  XNOR U26966 ( .A(n27561), .B(n27562), .Z(n27558) );
  AND U26967 ( .A(n740), .B(n27563), .Z(n27562) );
  XOR U26968 ( .A(n27564), .B(n27565), .Z(n27556) );
  AND U26969 ( .A(n744), .B(n27555), .Z(n27565) );
  XNOR U26970 ( .A(n27566), .B(n27553), .Z(n27555) );
  XOR U26971 ( .A(n27567), .B(n27568), .Z(n27553) );
  AND U26972 ( .A(n767), .B(n27569), .Z(n27568) );
  IV U26973 ( .A(n27564), .Z(n27566) );
  XOR U26974 ( .A(n27570), .B(n27571), .Z(n27564) );
  AND U26975 ( .A(n751), .B(n27563), .Z(n27571) );
  XNOR U26976 ( .A(n27561), .B(n27570), .Z(n27563) );
  XNOR U26977 ( .A(n27572), .B(n27573), .Z(n27561) );
  AND U26978 ( .A(n755), .B(n27574), .Z(n27573) );
  XOR U26979 ( .A(p_input[576]), .B(n27572), .Z(n27574) );
  XNOR U26980 ( .A(n27575), .B(n27576), .Z(n27572) );
  AND U26981 ( .A(n759), .B(n27577), .Z(n27576) );
  XOR U26982 ( .A(n27578), .B(n27579), .Z(n27570) );
  AND U26983 ( .A(n763), .B(n27569), .Z(n27579) );
  XNOR U26984 ( .A(n27580), .B(n27567), .Z(n27569) );
  XOR U26985 ( .A(n27581), .B(n27582), .Z(n27567) );
  AND U26986 ( .A(n786), .B(n27583), .Z(n27582) );
  IV U26987 ( .A(n27578), .Z(n27580) );
  XOR U26988 ( .A(n27584), .B(n27585), .Z(n27578) );
  AND U26989 ( .A(n770), .B(n27577), .Z(n27585) );
  XNOR U26990 ( .A(n27575), .B(n27584), .Z(n27577) );
  XNOR U26991 ( .A(n27586), .B(n27587), .Z(n27575) );
  AND U26992 ( .A(n774), .B(n27588), .Z(n27587) );
  XOR U26993 ( .A(p_input[592]), .B(n27586), .Z(n27588) );
  XNOR U26994 ( .A(n27589), .B(n27590), .Z(n27586) );
  AND U26995 ( .A(n778), .B(n27591), .Z(n27590) );
  XOR U26996 ( .A(n27592), .B(n27593), .Z(n27584) );
  AND U26997 ( .A(n782), .B(n27583), .Z(n27593) );
  XNOR U26998 ( .A(n27594), .B(n27581), .Z(n27583) );
  XOR U26999 ( .A(n27595), .B(n27596), .Z(n27581) );
  AND U27000 ( .A(n805), .B(n27597), .Z(n27596) );
  IV U27001 ( .A(n27592), .Z(n27594) );
  XOR U27002 ( .A(n27598), .B(n27599), .Z(n27592) );
  AND U27003 ( .A(n789), .B(n27591), .Z(n27599) );
  XNOR U27004 ( .A(n27589), .B(n27598), .Z(n27591) );
  XNOR U27005 ( .A(n27600), .B(n27601), .Z(n27589) );
  AND U27006 ( .A(n793), .B(n27602), .Z(n27601) );
  XOR U27007 ( .A(p_input[608]), .B(n27600), .Z(n27602) );
  XNOR U27008 ( .A(n27603), .B(n27604), .Z(n27600) );
  AND U27009 ( .A(n797), .B(n27605), .Z(n27604) );
  XOR U27010 ( .A(n27606), .B(n27607), .Z(n27598) );
  AND U27011 ( .A(n801), .B(n27597), .Z(n27607) );
  XNOR U27012 ( .A(n27608), .B(n27595), .Z(n27597) );
  XOR U27013 ( .A(n27609), .B(n27610), .Z(n27595) );
  AND U27014 ( .A(n824), .B(n27611), .Z(n27610) );
  IV U27015 ( .A(n27606), .Z(n27608) );
  XOR U27016 ( .A(n27612), .B(n27613), .Z(n27606) );
  AND U27017 ( .A(n808), .B(n27605), .Z(n27613) );
  XNOR U27018 ( .A(n27603), .B(n27612), .Z(n27605) );
  XNOR U27019 ( .A(n27614), .B(n27615), .Z(n27603) );
  AND U27020 ( .A(n812), .B(n27616), .Z(n27615) );
  XOR U27021 ( .A(p_input[624]), .B(n27614), .Z(n27616) );
  XNOR U27022 ( .A(n27617), .B(n27618), .Z(n27614) );
  AND U27023 ( .A(n816), .B(n27619), .Z(n27618) );
  XOR U27024 ( .A(n27620), .B(n27621), .Z(n27612) );
  AND U27025 ( .A(n820), .B(n27611), .Z(n27621) );
  XNOR U27026 ( .A(n27622), .B(n27609), .Z(n27611) );
  XOR U27027 ( .A(n27623), .B(n27624), .Z(n27609) );
  AND U27028 ( .A(n843), .B(n27625), .Z(n27624) );
  IV U27029 ( .A(n27620), .Z(n27622) );
  XOR U27030 ( .A(n27626), .B(n27627), .Z(n27620) );
  AND U27031 ( .A(n827), .B(n27619), .Z(n27627) );
  XNOR U27032 ( .A(n27617), .B(n27626), .Z(n27619) );
  XNOR U27033 ( .A(n27628), .B(n27629), .Z(n27617) );
  AND U27034 ( .A(n831), .B(n27630), .Z(n27629) );
  XOR U27035 ( .A(p_input[640]), .B(n27628), .Z(n27630) );
  XNOR U27036 ( .A(n27631), .B(n27632), .Z(n27628) );
  AND U27037 ( .A(n835), .B(n27633), .Z(n27632) );
  XOR U27038 ( .A(n27634), .B(n27635), .Z(n27626) );
  AND U27039 ( .A(n839), .B(n27625), .Z(n27635) );
  XNOR U27040 ( .A(n27636), .B(n27623), .Z(n27625) );
  XOR U27041 ( .A(n27637), .B(n27638), .Z(n27623) );
  AND U27042 ( .A(n862), .B(n27639), .Z(n27638) );
  IV U27043 ( .A(n27634), .Z(n27636) );
  XOR U27044 ( .A(n27640), .B(n27641), .Z(n27634) );
  AND U27045 ( .A(n846), .B(n27633), .Z(n27641) );
  XNOR U27046 ( .A(n27631), .B(n27640), .Z(n27633) );
  XNOR U27047 ( .A(n27642), .B(n27643), .Z(n27631) );
  AND U27048 ( .A(n850), .B(n27644), .Z(n27643) );
  XOR U27049 ( .A(p_input[656]), .B(n27642), .Z(n27644) );
  XNOR U27050 ( .A(n27645), .B(n27646), .Z(n27642) );
  AND U27051 ( .A(n854), .B(n27647), .Z(n27646) );
  XOR U27052 ( .A(n27648), .B(n27649), .Z(n27640) );
  AND U27053 ( .A(n858), .B(n27639), .Z(n27649) );
  XNOR U27054 ( .A(n27650), .B(n27637), .Z(n27639) );
  XOR U27055 ( .A(n27651), .B(n27652), .Z(n27637) );
  AND U27056 ( .A(n881), .B(n27653), .Z(n27652) );
  IV U27057 ( .A(n27648), .Z(n27650) );
  XOR U27058 ( .A(n27654), .B(n27655), .Z(n27648) );
  AND U27059 ( .A(n865), .B(n27647), .Z(n27655) );
  XNOR U27060 ( .A(n27645), .B(n27654), .Z(n27647) );
  XNOR U27061 ( .A(n27656), .B(n27657), .Z(n27645) );
  AND U27062 ( .A(n869), .B(n27658), .Z(n27657) );
  XOR U27063 ( .A(p_input[672]), .B(n27656), .Z(n27658) );
  XNOR U27064 ( .A(n27659), .B(n27660), .Z(n27656) );
  AND U27065 ( .A(n873), .B(n27661), .Z(n27660) );
  XOR U27066 ( .A(n27662), .B(n27663), .Z(n27654) );
  AND U27067 ( .A(n877), .B(n27653), .Z(n27663) );
  XNOR U27068 ( .A(n27664), .B(n27651), .Z(n27653) );
  XOR U27069 ( .A(n27665), .B(n27666), .Z(n27651) );
  AND U27070 ( .A(n900), .B(n27667), .Z(n27666) );
  IV U27071 ( .A(n27662), .Z(n27664) );
  XOR U27072 ( .A(n27668), .B(n27669), .Z(n27662) );
  AND U27073 ( .A(n884), .B(n27661), .Z(n27669) );
  XNOR U27074 ( .A(n27659), .B(n27668), .Z(n27661) );
  XNOR U27075 ( .A(n27670), .B(n27671), .Z(n27659) );
  AND U27076 ( .A(n888), .B(n27672), .Z(n27671) );
  XOR U27077 ( .A(p_input[688]), .B(n27670), .Z(n27672) );
  XNOR U27078 ( .A(n27673), .B(n27674), .Z(n27670) );
  AND U27079 ( .A(n892), .B(n27675), .Z(n27674) );
  XOR U27080 ( .A(n27676), .B(n27677), .Z(n27668) );
  AND U27081 ( .A(n896), .B(n27667), .Z(n27677) );
  XNOR U27082 ( .A(n27678), .B(n27665), .Z(n27667) );
  XOR U27083 ( .A(n27679), .B(n27680), .Z(n27665) );
  AND U27084 ( .A(n919), .B(n27681), .Z(n27680) );
  IV U27085 ( .A(n27676), .Z(n27678) );
  XOR U27086 ( .A(n27682), .B(n27683), .Z(n27676) );
  AND U27087 ( .A(n903), .B(n27675), .Z(n27683) );
  XNOR U27088 ( .A(n27673), .B(n27682), .Z(n27675) );
  XNOR U27089 ( .A(n27684), .B(n27685), .Z(n27673) );
  AND U27090 ( .A(n907), .B(n27686), .Z(n27685) );
  XOR U27091 ( .A(p_input[704]), .B(n27684), .Z(n27686) );
  XNOR U27092 ( .A(n27687), .B(n27688), .Z(n27684) );
  AND U27093 ( .A(n911), .B(n27689), .Z(n27688) );
  XOR U27094 ( .A(n27690), .B(n27691), .Z(n27682) );
  AND U27095 ( .A(n915), .B(n27681), .Z(n27691) );
  XNOR U27096 ( .A(n27692), .B(n27679), .Z(n27681) );
  XOR U27097 ( .A(n27693), .B(n27694), .Z(n27679) );
  AND U27098 ( .A(n938), .B(n27695), .Z(n27694) );
  IV U27099 ( .A(n27690), .Z(n27692) );
  XOR U27100 ( .A(n27696), .B(n27697), .Z(n27690) );
  AND U27101 ( .A(n922), .B(n27689), .Z(n27697) );
  XNOR U27102 ( .A(n27687), .B(n27696), .Z(n27689) );
  XNOR U27103 ( .A(n27698), .B(n27699), .Z(n27687) );
  AND U27104 ( .A(n926), .B(n27700), .Z(n27699) );
  XOR U27105 ( .A(p_input[720]), .B(n27698), .Z(n27700) );
  XNOR U27106 ( .A(n27701), .B(n27702), .Z(n27698) );
  AND U27107 ( .A(n930), .B(n27703), .Z(n27702) );
  XOR U27108 ( .A(n27704), .B(n27705), .Z(n27696) );
  AND U27109 ( .A(n934), .B(n27695), .Z(n27705) );
  XNOR U27110 ( .A(n27706), .B(n27693), .Z(n27695) );
  XOR U27111 ( .A(n27707), .B(n27708), .Z(n27693) );
  AND U27112 ( .A(n957), .B(n27709), .Z(n27708) );
  IV U27113 ( .A(n27704), .Z(n27706) );
  XOR U27114 ( .A(n27710), .B(n27711), .Z(n27704) );
  AND U27115 ( .A(n941), .B(n27703), .Z(n27711) );
  XNOR U27116 ( .A(n27701), .B(n27710), .Z(n27703) );
  XNOR U27117 ( .A(n27712), .B(n27713), .Z(n27701) );
  AND U27118 ( .A(n945), .B(n27714), .Z(n27713) );
  XOR U27119 ( .A(p_input[736]), .B(n27712), .Z(n27714) );
  XNOR U27120 ( .A(n27715), .B(n27716), .Z(n27712) );
  AND U27121 ( .A(n949), .B(n27717), .Z(n27716) );
  XOR U27122 ( .A(n27718), .B(n27719), .Z(n27710) );
  AND U27123 ( .A(n953), .B(n27709), .Z(n27719) );
  XNOR U27124 ( .A(n27720), .B(n27707), .Z(n27709) );
  XOR U27125 ( .A(n27721), .B(n27722), .Z(n27707) );
  AND U27126 ( .A(n976), .B(n27723), .Z(n27722) );
  IV U27127 ( .A(n27718), .Z(n27720) );
  XOR U27128 ( .A(n27724), .B(n27725), .Z(n27718) );
  AND U27129 ( .A(n960), .B(n27717), .Z(n27725) );
  XNOR U27130 ( .A(n27715), .B(n27724), .Z(n27717) );
  XNOR U27131 ( .A(n27726), .B(n27727), .Z(n27715) );
  AND U27132 ( .A(n964), .B(n27728), .Z(n27727) );
  XOR U27133 ( .A(p_input[752]), .B(n27726), .Z(n27728) );
  XNOR U27134 ( .A(n27729), .B(n27730), .Z(n27726) );
  AND U27135 ( .A(n968), .B(n27731), .Z(n27730) );
  XOR U27136 ( .A(n27732), .B(n27733), .Z(n27724) );
  AND U27137 ( .A(n972), .B(n27723), .Z(n27733) );
  XNOR U27138 ( .A(n27734), .B(n27721), .Z(n27723) );
  XOR U27139 ( .A(n27735), .B(n27736), .Z(n27721) );
  AND U27140 ( .A(n995), .B(n27737), .Z(n27736) );
  IV U27141 ( .A(n27732), .Z(n27734) );
  XOR U27142 ( .A(n27738), .B(n27739), .Z(n27732) );
  AND U27143 ( .A(n979), .B(n27731), .Z(n27739) );
  XNOR U27144 ( .A(n27729), .B(n27738), .Z(n27731) );
  XNOR U27145 ( .A(n27740), .B(n27741), .Z(n27729) );
  AND U27146 ( .A(n983), .B(n27742), .Z(n27741) );
  XOR U27147 ( .A(p_input[768]), .B(n27740), .Z(n27742) );
  XNOR U27148 ( .A(n27743), .B(n27744), .Z(n27740) );
  AND U27149 ( .A(n987), .B(n27745), .Z(n27744) );
  XOR U27150 ( .A(n27746), .B(n27747), .Z(n27738) );
  AND U27151 ( .A(n991), .B(n27737), .Z(n27747) );
  XNOR U27152 ( .A(n27748), .B(n27735), .Z(n27737) );
  XOR U27153 ( .A(n27749), .B(n27750), .Z(n27735) );
  AND U27154 ( .A(n1014), .B(n27751), .Z(n27750) );
  IV U27155 ( .A(n27746), .Z(n27748) );
  XOR U27156 ( .A(n27752), .B(n27753), .Z(n27746) );
  AND U27157 ( .A(n998), .B(n27745), .Z(n27753) );
  XNOR U27158 ( .A(n27743), .B(n27752), .Z(n27745) );
  XNOR U27159 ( .A(n27754), .B(n27755), .Z(n27743) );
  AND U27160 ( .A(n1002), .B(n27756), .Z(n27755) );
  XOR U27161 ( .A(p_input[784]), .B(n27754), .Z(n27756) );
  XNOR U27162 ( .A(n27757), .B(n27758), .Z(n27754) );
  AND U27163 ( .A(n1006), .B(n27759), .Z(n27758) );
  XOR U27164 ( .A(n27760), .B(n27761), .Z(n27752) );
  AND U27165 ( .A(n1010), .B(n27751), .Z(n27761) );
  XNOR U27166 ( .A(n27762), .B(n27749), .Z(n27751) );
  XOR U27167 ( .A(n27763), .B(n27764), .Z(n27749) );
  AND U27168 ( .A(n1033), .B(n27765), .Z(n27764) );
  IV U27169 ( .A(n27760), .Z(n27762) );
  XOR U27170 ( .A(n27766), .B(n27767), .Z(n27760) );
  AND U27171 ( .A(n1017), .B(n27759), .Z(n27767) );
  XNOR U27172 ( .A(n27757), .B(n27766), .Z(n27759) );
  XNOR U27173 ( .A(n27768), .B(n27769), .Z(n27757) );
  AND U27174 ( .A(n1021), .B(n27770), .Z(n27769) );
  XOR U27175 ( .A(p_input[800]), .B(n27768), .Z(n27770) );
  XNOR U27176 ( .A(n27771), .B(n27772), .Z(n27768) );
  AND U27177 ( .A(n1025), .B(n27773), .Z(n27772) );
  XOR U27178 ( .A(n27774), .B(n27775), .Z(n27766) );
  AND U27179 ( .A(n1029), .B(n27765), .Z(n27775) );
  XNOR U27180 ( .A(n27776), .B(n27763), .Z(n27765) );
  XOR U27181 ( .A(n27777), .B(n27778), .Z(n27763) );
  AND U27182 ( .A(n1052), .B(n27779), .Z(n27778) );
  IV U27183 ( .A(n27774), .Z(n27776) );
  XOR U27184 ( .A(n27780), .B(n27781), .Z(n27774) );
  AND U27185 ( .A(n1036), .B(n27773), .Z(n27781) );
  XNOR U27186 ( .A(n27771), .B(n27780), .Z(n27773) );
  XNOR U27187 ( .A(n27782), .B(n27783), .Z(n27771) );
  AND U27188 ( .A(n1040), .B(n27784), .Z(n27783) );
  XOR U27189 ( .A(p_input[816]), .B(n27782), .Z(n27784) );
  XNOR U27190 ( .A(n27785), .B(n27786), .Z(n27782) );
  AND U27191 ( .A(n1044), .B(n27787), .Z(n27786) );
  XOR U27192 ( .A(n27788), .B(n27789), .Z(n27780) );
  AND U27193 ( .A(n1048), .B(n27779), .Z(n27789) );
  XNOR U27194 ( .A(n27790), .B(n27777), .Z(n27779) );
  XOR U27195 ( .A(n27791), .B(n27792), .Z(n27777) );
  AND U27196 ( .A(n1071), .B(n27793), .Z(n27792) );
  IV U27197 ( .A(n27788), .Z(n27790) );
  XOR U27198 ( .A(n27794), .B(n27795), .Z(n27788) );
  AND U27199 ( .A(n1055), .B(n27787), .Z(n27795) );
  XNOR U27200 ( .A(n27785), .B(n27794), .Z(n27787) );
  XNOR U27201 ( .A(n27796), .B(n27797), .Z(n27785) );
  AND U27202 ( .A(n1059), .B(n27798), .Z(n27797) );
  XOR U27203 ( .A(p_input[832]), .B(n27796), .Z(n27798) );
  XNOR U27204 ( .A(n27799), .B(n27800), .Z(n27796) );
  AND U27205 ( .A(n1063), .B(n27801), .Z(n27800) );
  XOR U27206 ( .A(n27802), .B(n27803), .Z(n27794) );
  AND U27207 ( .A(n1067), .B(n27793), .Z(n27803) );
  XNOR U27208 ( .A(n27804), .B(n27791), .Z(n27793) );
  XOR U27209 ( .A(n27805), .B(n27806), .Z(n27791) );
  AND U27210 ( .A(n1090), .B(n27807), .Z(n27806) );
  IV U27211 ( .A(n27802), .Z(n27804) );
  XOR U27212 ( .A(n27808), .B(n27809), .Z(n27802) );
  AND U27213 ( .A(n1074), .B(n27801), .Z(n27809) );
  XNOR U27214 ( .A(n27799), .B(n27808), .Z(n27801) );
  XNOR U27215 ( .A(n27810), .B(n27811), .Z(n27799) );
  AND U27216 ( .A(n1078), .B(n27812), .Z(n27811) );
  XOR U27217 ( .A(p_input[848]), .B(n27810), .Z(n27812) );
  XNOR U27218 ( .A(n27813), .B(n27814), .Z(n27810) );
  AND U27219 ( .A(n1082), .B(n27815), .Z(n27814) );
  XOR U27220 ( .A(n27816), .B(n27817), .Z(n27808) );
  AND U27221 ( .A(n1086), .B(n27807), .Z(n27817) );
  XNOR U27222 ( .A(n27818), .B(n27805), .Z(n27807) );
  XOR U27223 ( .A(n27819), .B(n27820), .Z(n27805) );
  AND U27224 ( .A(n1109), .B(n27821), .Z(n27820) );
  IV U27225 ( .A(n27816), .Z(n27818) );
  XOR U27226 ( .A(n27822), .B(n27823), .Z(n27816) );
  AND U27227 ( .A(n1093), .B(n27815), .Z(n27823) );
  XNOR U27228 ( .A(n27813), .B(n27822), .Z(n27815) );
  XNOR U27229 ( .A(n27824), .B(n27825), .Z(n27813) );
  AND U27230 ( .A(n1097), .B(n27826), .Z(n27825) );
  XOR U27231 ( .A(p_input[864]), .B(n27824), .Z(n27826) );
  XNOR U27232 ( .A(n27827), .B(n27828), .Z(n27824) );
  AND U27233 ( .A(n1101), .B(n27829), .Z(n27828) );
  XOR U27234 ( .A(n27830), .B(n27831), .Z(n27822) );
  AND U27235 ( .A(n1105), .B(n27821), .Z(n27831) );
  XNOR U27236 ( .A(n27832), .B(n27819), .Z(n27821) );
  XOR U27237 ( .A(n27833), .B(n27834), .Z(n27819) );
  AND U27238 ( .A(n1128), .B(n27835), .Z(n27834) );
  IV U27239 ( .A(n27830), .Z(n27832) );
  XOR U27240 ( .A(n27836), .B(n27837), .Z(n27830) );
  AND U27241 ( .A(n1112), .B(n27829), .Z(n27837) );
  XNOR U27242 ( .A(n27827), .B(n27836), .Z(n27829) );
  XNOR U27243 ( .A(n27838), .B(n27839), .Z(n27827) );
  AND U27244 ( .A(n1116), .B(n27840), .Z(n27839) );
  XOR U27245 ( .A(p_input[880]), .B(n27838), .Z(n27840) );
  XNOR U27246 ( .A(n27841), .B(n27842), .Z(n27838) );
  AND U27247 ( .A(n1120), .B(n27843), .Z(n27842) );
  XOR U27248 ( .A(n27844), .B(n27845), .Z(n27836) );
  AND U27249 ( .A(n1124), .B(n27835), .Z(n27845) );
  XNOR U27250 ( .A(n27846), .B(n27833), .Z(n27835) );
  XOR U27251 ( .A(n27847), .B(n27848), .Z(n27833) );
  AND U27252 ( .A(n1147), .B(n27849), .Z(n27848) );
  IV U27253 ( .A(n27844), .Z(n27846) );
  XOR U27254 ( .A(n27850), .B(n27851), .Z(n27844) );
  AND U27255 ( .A(n1131), .B(n27843), .Z(n27851) );
  XNOR U27256 ( .A(n27841), .B(n27850), .Z(n27843) );
  XNOR U27257 ( .A(n27852), .B(n27853), .Z(n27841) );
  AND U27258 ( .A(n1135), .B(n27854), .Z(n27853) );
  XOR U27259 ( .A(p_input[896]), .B(n27852), .Z(n27854) );
  XNOR U27260 ( .A(n27855), .B(n27856), .Z(n27852) );
  AND U27261 ( .A(n1139), .B(n27857), .Z(n27856) );
  XOR U27262 ( .A(n27858), .B(n27859), .Z(n27850) );
  AND U27263 ( .A(n1143), .B(n27849), .Z(n27859) );
  XNOR U27264 ( .A(n27860), .B(n27847), .Z(n27849) );
  XOR U27265 ( .A(n27861), .B(n27862), .Z(n27847) );
  AND U27266 ( .A(n1166), .B(n27863), .Z(n27862) );
  IV U27267 ( .A(n27858), .Z(n27860) );
  XOR U27268 ( .A(n27864), .B(n27865), .Z(n27858) );
  AND U27269 ( .A(n1150), .B(n27857), .Z(n27865) );
  XNOR U27270 ( .A(n27855), .B(n27864), .Z(n27857) );
  XNOR U27271 ( .A(n27866), .B(n27867), .Z(n27855) );
  AND U27272 ( .A(n1154), .B(n27868), .Z(n27867) );
  XOR U27273 ( .A(p_input[912]), .B(n27866), .Z(n27868) );
  XNOR U27274 ( .A(n27869), .B(n27870), .Z(n27866) );
  AND U27275 ( .A(n1158), .B(n27871), .Z(n27870) );
  XOR U27276 ( .A(n27872), .B(n27873), .Z(n27864) );
  AND U27277 ( .A(n1162), .B(n27863), .Z(n27873) );
  XNOR U27278 ( .A(n27874), .B(n27861), .Z(n27863) );
  XOR U27279 ( .A(n27875), .B(n27876), .Z(n27861) );
  AND U27280 ( .A(n1185), .B(n27877), .Z(n27876) );
  IV U27281 ( .A(n27872), .Z(n27874) );
  XOR U27282 ( .A(n27878), .B(n27879), .Z(n27872) );
  AND U27283 ( .A(n1169), .B(n27871), .Z(n27879) );
  XNOR U27284 ( .A(n27869), .B(n27878), .Z(n27871) );
  XNOR U27285 ( .A(n27880), .B(n27881), .Z(n27869) );
  AND U27286 ( .A(n1173), .B(n27882), .Z(n27881) );
  XOR U27287 ( .A(p_input[928]), .B(n27880), .Z(n27882) );
  XNOR U27288 ( .A(n27883), .B(n27884), .Z(n27880) );
  AND U27289 ( .A(n1177), .B(n27885), .Z(n27884) );
  XOR U27290 ( .A(n27886), .B(n27887), .Z(n27878) );
  AND U27291 ( .A(n1181), .B(n27877), .Z(n27887) );
  XNOR U27292 ( .A(n27888), .B(n27875), .Z(n27877) );
  XOR U27293 ( .A(n27889), .B(n27890), .Z(n27875) );
  AND U27294 ( .A(n1204), .B(n27891), .Z(n27890) );
  IV U27295 ( .A(n27886), .Z(n27888) );
  XOR U27296 ( .A(n27892), .B(n27893), .Z(n27886) );
  AND U27297 ( .A(n1188), .B(n27885), .Z(n27893) );
  XNOR U27298 ( .A(n27883), .B(n27892), .Z(n27885) );
  XNOR U27299 ( .A(n27894), .B(n27895), .Z(n27883) );
  AND U27300 ( .A(n1192), .B(n27896), .Z(n27895) );
  XOR U27301 ( .A(p_input[944]), .B(n27894), .Z(n27896) );
  XNOR U27302 ( .A(n27897), .B(n27898), .Z(n27894) );
  AND U27303 ( .A(n1196), .B(n27899), .Z(n27898) );
  XOR U27304 ( .A(n27900), .B(n27901), .Z(n27892) );
  AND U27305 ( .A(n1200), .B(n27891), .Z(n27901) );
  XNOR U27306 ( .A(n27902), .B(n27889), .Z(n27891) );
  XOR U27307 ( .A(n27903), .B(n27904), .Z(n27889) );
  AND U27308 ( .A(n1223), .B(n27905), .Z(n27904) );
  IV U27309 ( .A(n27900), .Z(n27902) );
  XOR U27310 ( .A(n27906), .B(n27907), .Z(n27900) );
  AND U27311 ( .A(n1207), .B(n27899), .Z(n27907) );
  XNOR U27312 ( .A(n27897), .B(n27906), .Z(n27899) );
  XNOR U27313 ( .A(n27908), .B(n27909), .Z(n27897) );
  AND U27314 ( .A(n1211), .B(n27910), .Z(n27909) );
  XOR U27315 ( .A(p_input[960]), .B(n27908), .Z(n27910) );
  XNOR U27316 ( .A(n27911), .B(n27912), .Z(n27908) );
  AND U27317 ( .A(n1215), .B(n27913), .Z(n27912) );
  XOR U27318 ( .A(n27914), .B(n27915), .Z(n27906) );
  AND U27319 ( .A(n1219), .B(n27905), .Z(n27915) );
  XNOR U27320 ( .A(n27916), .B(n27903), .Z(n27905) );
  XOR U27321 ( .A(n27917), .B(n27918), .Z(n27903) );
  AND U27322 ( .A(n1242), .B(n27919), .Z(n27918) );
  IV U27323 ( .A(n27914), .Z(n27916) );
  XOR U27324 ( .A(n27920), .B(n27921), .Z(n27914) );
  AND U27325 ( .A(n1226), .B(n27913), .Z(n27921) );
  XNOR U27326 ( .A(n27911), .B(n27920), .Z(n27913) );
  XNOR U27327 ( .A(n27922), .B(n27923), .Z(n27911) );
  AND U27328 ( .A(n1230), .B(n27924), .Z(n27923) );
  XOR U27329 ( .A(p_input[976]), .B(n27922), .Z(n27924) );
  XNOR U27330 ( .A(n27925), .B(n27926), .Z(n27922) );
  AND U27331 ( .A(n1234), .B(n27927), .Z(n27926) );
  XOR U27332 ( .A(n27928), .B(n27929), .Z(n27920) );
  AND U27333 ( .A(n1238), .B(n27919), .Z(n27929) );
  XNOR U27334 ( .A(n27930), .B(n27917), .Z(n27919) );
  XOR U27335 ( .A(n27931), .B(n27932), .Z(n27917) );
  AND U27336 ( .A(n1261), .B(n27933), .Z(n27932) );
  IV U27337 ( .A(n27928), .Z(n27930) );
  XOR U27338 ( .A(n27934), .B(n27935), .Z(n27928) );
  AND U27339 ( .A(n1245), .B(n27927), .Z(n27935) );
  XNOR U27340 ( .A(n27925), .B(n27934), .Z(n27927) );
  XNOR U27341 ( .A(n27936), .B(n27937), .Z(n27925) );
  AND U27342 ( .A(n1249), .B(n27938), .Z(n27937) );
  XOR U27343 ( .A(p_input[992]), .B(n27936), .Z(n27938) );
  XNOR U27344 ( .A(n27939), .B(n27940), .Z(n27936) );
  AND U27345 ( .A(n1253), .B(n27941), .Z(n27940) );
  XOR U27346 ( .A(n27942), .B(n27943), .Z(n27934) );
  AND U27347 ( .A(n1257), .B(n27933), .Z(n27943) );
  XNOR U27348 ( .A(n27944), .B(n27931), .Z(n27933) );
  XOR U27349 ( .A(n27945), .B(n27946), .Z(n27931) );
  AND U27350 ( .A(n1280), .B(n27947), .Z(n27946) );
  IV U27351 ( .A(n27942), .Z(n27944) );
  XOR U27352 ( .A(n27948), .B(n27949), .Z(n27942) );
  AND U27353 ( .A(n1264), .B(n27941), .Z(n27949) );
  XNOR U27354 ( .A(n27939), .B(n27948), .Z(n27941) );
  XNOR U27355 ( .A(n27950), .B(n27951), .Z(n27939) );
  AND U27356 ( .A(n1268), .B(n27952), .Z(n27951) );
  XOR U27357 ( .A(p_input[1008]), .B(n27950), .Z(n27952) );
  XNOR U27358 ( .A(n27953), .B(n27954), .Z(n27950) );
  AND U27359 ( .A(n1272), .B(n27955), .Z(n27954) );
  XOR U27360 ( .A(n27956), .B(n27957), .Z(n27948) );
  AND U27361 ( .A(n1276), .B(n27947), .Z(n27957) );
  XNOR U27362 ( .A(n27958), .B(n27945), .Z(n27947) );
  XOR U27363 ( .A(n27959), .B(n27960), .Z(n27945) );
  AND U27364 ( .A(n1299), .B(n27961), .Z(n27960) );
  IV U27365 ( .A(n27956), .Z(n27958) );
  XOR U27366 ( .A(n27962), .B(n27963), .Z(n27956) );
  AND U27367 ( .A(n1283), .B(n27955), .Z(n27963) );
  XNOR U27368 ( .A(n27953), .B(n27962), .Z(n27955) );
  XNOR U27369 ( .A(n27964), .B(n27965), .Z(n27953) );
  AND U27370 ( .A(n1287), .B(n27966), .Z(n27965) );
  XOR U27371 ( .A(p_input[1024]), .B(n27964), .Z(n27966) );
  XNOR U27372 ( .A(n27967), .B(n27968), .Z(n27964) );
  AND U27373 ( .A(n1291), .B(n27969), .Z(n27968) );
  XOR U27374 ( .A(n27970), .B(n27971), .Z(n27962) );
  AND U27375 ( .A(n1295), .B(n27961), .Z(n27971) );
  XNOR U27376 ( .A(n27972), .B(n27959), .Z(n27961) );
  XOR U27377 ( .A(n27973), .B(n27974), .Z(n27959) );
  AND U27378 ( .A(n1318), .B(n27975), .Z(n27974) );
  IV U27379 ( .A(n27970), .Z(n27972) );
  XOR U27380 ( .A(n27976), .B(n27977), .Z(n27970) );
  AND U27381 ( .A(n1302), .B(n27969), .Z(n27977) );
  XNOR U27382 ( .A(n27967), .B(n27976), .Z(n27969) );
  XNOR U27383 ( .A(n27978), .B(n27979), .Z(n27967) );
  AND U27384 ( .A(n1306), .B(n27980), .Z(n27979) );
  XOR U27385 ( .A(p_input[1040]), .B(n27978), .Z(n27980) );
  XNOR U27386 ( .A(n27981), .B(n27982), .Z(n27978) );
  AND U27387 ( .A(n1310), .B(n27983), .Z(n27982) );
  XOR U27388 ( .A(n27984), .B(n27985), .Z(n27976) );
  AND U27389 ( .A(n1314), .B(n27975), .Z(n27985) );
  XNOR U27390 ( .A(n27986), .B(n27973), .Z(n27975) );
  XOR U27391 ( .A(n27987), .B(n27988), .Z(n27973) );
  AND U27392 ( .A(n1337), .B(n27989), .Z(n27988) );
  IV U27393 ( .A(n27984), .Z(n27986) );
  XOR U27394 ( .A(n27990), .B(n27991), .Z(n27984) );
  AND U27395 ( .A(n1321), .B(n27983), .Z(n27991) );
  XNOR U27396 ( .A(n27981), .B(n27990), .Z(n27983) );
  XNOR U27397 ( .A(n27992), .B(n27993), .Z(n27981) );
  AND U27398 ( .A(n1325), .B(n27994), .Z(n27993) );
  XOR U27399 ( .A(p_input[1056]), .B(n27992), .Z(n27994) );
  XNOR U27400 ( .A(n27995), .B(n27996), .Z(n27992) );
  AND U27401 ( .A(n1329), .B(n27997), .Z(n27996) );
  XOR U27402 ( .A(n27998), .B(n27999), .Z(n27990) );
  AND U27403 ( .A(n1333), .B(n27989), .Z(n27999) );
  XNOR U27404 ( .A(n28000), .B(n27987), .Z(n27989) );
  XOR U27405 ( .A(n28001), .B(n28002), .Z(n27987) );
  AND U27406 ( .A(n1356), .B(n28003), .Z(n28002) );
  IV U27407 ( .A(n27998), .Z(n28000) );
  XOR U27408 ( .A(n28004), .B(n28005), .Z(n27998) );
  AND U27409 ( .A(n1340), .B(n27997), .Z(n28005) );
  XNOR U27410 ( .A(n27995), .B(n28004), .Z(n27997) );
  XNOR U27411 ( .A(n28006), .B(n28007), .Z(n27995) );
  AND U27412 ( .A(n1344), .B(n28008), .Z(n28007) );
  XOR U27413 ( .A(p_input[1072]), .B(n28006), .Z(n28008) );
  XNOR U27414 ( .A(n28009), .B(n28010), .Z(n28006) );
  AND U27415 ( .A(n1348), .B(n28011), .Z(n28010) );
  XOR U27416 ( .A(n28012), .B(n28013), .Z(n28004) );
  AND U27417 ( .A(n1352), .B(n28003), .Z(n28013) );
  XNOR U27418 ( .A(n28014), .B(n28001), .Z(n28003) );
  XOR U27419 ( .A(n28015), .B(n28016), .Z(n28001) );
  AND U27420 ( .A(n1375), .B(n28017), .Z(n28016) );
  IV U27421 ( .A(n28012), .Z(n28014) );
  XOR U27422 ( .A(n28018), .B(n28019), .Z(n28012) );
  AND U27423 ( .A(n1359), .B(n28011), .Z(n28019) );
  XNOR U27424 ( .A(n28009), .B(n28018), .Z(n28011) );
  XNOR U27425 ( .A(n28020), .B(n28021), .Z(n28009) );
  AND U27426 ( .A(n1363), .B(n28022), .Z(n28021) );
  XOR U27427 ( .A(p_input[1088]), .B(n28020), .Z(n28022) );
  XNOR U27428 ( .A(n28023), .B(n28024), .Z(n28020) );
  AND U27429 ( .A(n1367), .B(n28025), .Z(n28024) );
  XOR U27430 ( .A(n28026), .B(n28027), .Z(n28018) );
  AND U27431 ( .A(n1371), .B(n28017), .Z(n28027) );
  XNOR U27432 ( .A(n28028), .B(n28015), .Z(n28017) );
  XOR U27433 ( .A(n28029), .B(n28030), .Z(n28015) );
  AND U27434 ( .A(n1394), .B(n28031), .Z(n28030) );
  IV U27435 ( .A(n28026), .Z(n28028) );
  XOR U27436 ( .A(n28032), .B(n28033), .Z(n28026) );
  AND U27437 ( .A(n1378), .B(n28025), .Z(n28033) );
  XNOR U27438 ( .A(n28023), .B(n28032), .Z(n28025) );
  XNOR U27439 ( .A(n28034), .B(n28035), .Z(n28023) );
  AND U27440 ( .A(n1382), .B(n28036), .Z(n28035) );
  XOR U27441 ( .A(p_input[1104]), .B(n28034), .Z(n28036) );
  XNOR U27442 ( .A(n28037), .B(n28038), .Z(n28034) );
  AND U27443 ( .A(n1386), .B(n28039), .Z(n28038) );
  XOR U27444 ( .A(n28040), .B(n28041), .Z(n28032) );
  AND U27445 ( .A(n1390), .B(n28031), .Z(n28041) );
  XNOR U27446 ( .A(n28042), .B(n28029), .Z(n28031) );
  XOR U27447 ( .A(n28043), .B(n28044), .Z(n28029) );
  AND U27448 ( .A(n1413), .B(n28045), .Z(n28044) );
  IV U27449 ( .A(n28040), .Z(n28042) );
  XOR U27450 ( .A(n28046), .B(n28047), .Z(n28040) );
  AND U27451 ( .A(n1397), .B(n28039), .Z(n28047) );
  XNOR U27452 ( .A(n28037), .B(n28046), .Z(n28039) );
  XNOR U27453 ( .A(n28048), .B(n28049), .Z(n28037) );
  AND U27454 ( .A(n1401), .B(n28050), .Z(n28049) );
  XOR U27455 ( .A(p_input[1120]), .B(n28048), .Z(n28050) );
  XNOR U27456 ( .A(n28051), .B(n28052), .Z(n28048) );
  AND U27457 ( .A(n1405), .B(n28053), .Z(n28052) );
  XOR U27458 ( .A(n28054), .B(n28055), .Z(n28046) );
  AND U27459 ( .A(n1409), .B(n28045), .Z(n28055) );
  XNOR U27460 ( .A(n28056), .B(n28043), .Z(n28045) );
  XOR U27461 ( .A(n28057), .B(n28058), .Z(n28043) );
  AND U27462 ( .A(n1432), .B(n28059), .Z(n28058) );
  IV U27463 ( .A(n28054), .Z(n28056) );
  XOR U27464 ( .A(n28060), .B(n28061), .Z(n28054) );
  AND U27465 ( .A(n1416), .B(n28053), .Z(n28061) );
  XNOR U27466 ( .A(n28051), .B(n28060), .Z(n28053) );
  XNOR U27467 ( .A(n28062), .B(n28063), .Z(n28051) );
  AND U27468 ( .A(n1420), .B(n28064), .Z(n28063) );
  XOR U27469 ( .A(p_input[1136]), .B(n28062), .Z(n28064) );
  XNOR U27470 ( .A(n28065), .B(n28066), .Z(n28062) );
  AND U27471 ( .A(n1424), .B(n28067), .Z(n28066) );
  XOR U27472 ( .A(n28068), .B(n28069), .Z(n28060) );
  AND U27473 ( .A(n1428), .B(n28059), .Z(n28069) );
  XNOR U27474 ( .A(n28070), .B(n28057), .Z(n28059) );
  XOR U27475 ( .A(n28071), .B(n28072), .Z(n28057) );
  AND U27476 ( .A(n1451), .B(n28073), .Z(n28072) );
  IV U27477 ( .A(n28068), .Z(n28070) );
  XOR U27478 ( .A(n28074), .B(n28075), .Z(n28068) );
  AND U27479 ( .A(n1435), .B(n28067), .Z(n28075) );
  XNOR U27480 ( .A(n28065), .B(n28074), .Z(n28067) );
  XNOR U27481 ( .A(n28076), .B(n28077), .Z(n28065) );
  AND U27482 ( .A(n1439), .B(n28078), .Z(n28077) );
  XOR U27483 ( .A(p_input[1152]), .B(n28076), .Z(n28078) );
  XNOR U27484 ( .A(n28079), .B(n28080), .Z(n28076) );
  AND U27485 ( .A(n1443), .B(n28081), .Z(n28080) );
  XOR U27486 ( .A(n28082), .B(n28083), .Z(n28074) );
  AND U27487 ( .A(n1447), .B(n28073), .Z(n28083) );
  XNOR U27488 ( .A(n28084), .B(n28071), .Z(n28073) );
  XOR U27489 ( .A(n28085), .B(n28086), .Z(n28071) );
  AND U27490 ( .A(n1470), .B(n28087), .Z(n28086) );
  IV U27491 ( .A(n28082), .Z(n28084) );
  XOR U27492 ( .A(n28088), .B(n28089), .Z(n28082) );
  AND U27493 ( .A(n1454), .B(n28081), .Z(n28089) );
  XNOR U27494 ( .A(n28079), .B(n28088), .Z(n28081) );
  XNOR U27495 ( .A(n28090), .B(n28091), .Z(n28079) );
  AND U27496 ( .A(n1458), .B(n28092), .Z(n28091) );
  XOR U27497 ( .A(p_input[1168]), .B(n28090), .Z(n28092) );
  XNOR U27498 ( .A(n28093), .B(n28094), .Z(n28090) );
  AND U27499 ( .A(n1462), .B(n28095), .Z(n28094) );
  XOR U27500 ( .A(n28096), .B(n28097), .Z(n28088) );
  AND U27501 ( .A(n1466), .B(n28087), .Z(n28097) );
  XNOR U27502 ( .A(n28098), .B(n28085), .Z(n28087) );
  XOR U27503 ( .A(n28099), .B(n28100), .Z(n28085) );
  AND U27504 ( .A(n1489), .B(n28101), .Z(n28100) );
  IV U27505 ( .A(n28096), .Z(n28098) );
  XOR U27506 ( .A(n28102), .B(n28103), .Z(n28096) );
  AND U27507 ( .A(n1473), .B(n28095), .Z(n28103) );
  XNOR U27508 ( .A(n28093), .B(n28102), .Z(n28095) );
  XNOR U27509 ( .A(n28104), .B(n28105), .Z(n28093) );
  AND U27510 ( .A(n1477), .B(n28106), .Z(n28105) );
  XOR U27511 ( .A(p_input[1184]), .B(n28104), .Z(n28106) );
  XNOR U27512 ( .A(n28107), .B(n28108), .Z(n28104) );
  AND U27513 ( .A(n1481), .B(n28109), .Z(n28108) );
  XOR U27514 ( .A(n28110), .B(n28111), .Z(n28102) );
  AND U27515 ( .A(n1485), .B(n28101), .Z(n28111) );
  XNOR U27516 ( .A(n28112), .B(n28099), .Z(n28101) );
  XOR U27517 ( .A(n28113), .B(n28114), .Z(n28099) );
  AND U27518 ( .A(n1508), .B(n28115), .Z(n28114) );
  IV U27519 ( .A(n28110), .Z(n28112) );
  XOR U27520 ( .A(n28116), .B(n28117), .Z(n28110) );
  AND U27521 ( .A(n1492), .B(n28109), .Z(n28117) );
  XNOR U27522 ( .A(n28107), .B(n28116), .Z(n28109) );
  XNOR U27523 ( .A(n28118), .B(n28119), .Z(n28107) );
  AND U27524 ( .A(n1496), .B(n28120), .Z(n28119) );
  XOR U27525 ( .A(p_input[1200]), .B(n28118), .Z(n28120) );
  XNOR U27526 ( .A(n28121), .B(n28122), .Z(n28118) );
  AND U27527 ( .A(n1500), .B(n28123), .Z(n28122) );
  XOR U27528 ( .A(n28124), .B(n28125), .Z(n28116) );
  AND U27529 ( .A(n1504), .B(n28115), .Z(n28125) );
  XNOR U27530 ( .A(n28126), .B(n28113), .Z(n28115) );
  XOR U27531 ( .A(n28127), .B(n28128), .Z(n28113) );
  AND U27532 ( .A(n1527), .B(n28129), .Z(n28128) );
  IV U27533 ( .A(n28124), .Z(n28126) );
  XOR U27534 ( .A(n28130), .B(n28131), .Z(n28124) );
  AND U27535 ( .A(n1511), .B(n28123), .Z(n28131) );
  XNOR U27536 ( .A(n28121), .B(n28130), .Z(n28123) );
  XNOR U27537 ( .A(n28132), .B(n28133), .Z(n28121) );
  AND U27538 ( .A(n1515), .B(n28134), .Z(n28133) );
  XOR U27539 ( .A(p_input[1216]), .B(n28132), .Z(n28134) );
  XNOR U27540 ( .A(n28135), .B(n28136), .Z(n28132) );
  AND U27541 ( .A(n1519), .B(n28137), .Z(n28136) );
  XOR U27542 ( .A(n28138), .B(n28139), .Z(n28130) );
  AND U27543 ( .A(n1523), .B(n28129), .Z(n28139) );
  XNOR U27544 ( .A(n28140), .B(n28127), .Z(n28129) );
  XOR U27545 ( .A(n28141), .B(n28142), .Z(n28127) );
  AND U27546 ( .A(n1546), .B(n28143), .Z(n28142) );
  IV U27547 ( .A(n28138), .Z(n28140) );
  XOR U27548 ( .A(n28144), .B(n28145), .Z(n28138) );
  AND U27549 ( .A(n1530), .B(n28137), .Z(n28145) );
  XNOR U27550 ( .A(n28135), .B(n28144), .Z(n28137) );
  XNOR U27551 ( .A(n28146), .B(n28147), .Z(n28135) );
  AND U27552 ( .A(n1534), .B(n28148), .Z(n28147) );
  XOR U27553 ( .A(p_input[1232]), .B(n28146), .Z(n28148) );
  XNOR U27554 ( .A(n28149), .B(n28150), .Z(n28146) );
  AND U27555 ( .A(n1538), .B(n28151), .Z(n28150) );
  XOR U27556 ( .A(n28152), .B(n28153), .Z(n28144) );
  AND U27557 ( .A(n1542), .B(n28143), .Z(n28153) );
  XNOR U27558 ( .A(n28154), .B(n28141), .Z(n28143) );
  XOR U27559 ( .A(n28155), .B(n28156), .Z(n28141) );
  AND U27560 ( .A(n1565), .B(n28157), .Z(n28156) );
  IV U27561 ( .A(n28152), .Z(n28154) );
  XOR U27562 ( .A(n28158), .B(n28159), .Z(n28152) );
  AND U27563 ( .A(n1549), .B(n28151), .Z(n28159) );
  XNOR U27564 ( .A(n28149), .B(n28158), .Z(n28151) );
  XNOR U27565 ( .A(n28160), .B(n28161), .Z(n28149) );
  AND U27566 ( .A(n1553), .B(n28162), .Z(n28161) );
  XOR U27567 ( .A(p_input[1248]), .B(n28160), .Z(n28162) );
  XNOR U27568 ( .A(n28163), .B(n28164), .Z(n28160) );
  AND U27569 ( .A(n1557), .B(n28165), .Z(n28164) );
  XOR U27570 ( .A(n28166), .B(n28167), .Z(n28158) );
  AND U27571 ( .A(n1561), .B(n28157), .Z(n28167) );
  XNOR U27572 ( .A(n28168), .B(n28155), .Z(n28157) );
  XOR U27573 ( .A(n28169), .B(n28170), .Z(n28155) );
  AND U27574 ( .A(n1584), .B(n28171), .Z(n28170) );
  IV U27575 ( .A(n28166), .Z(n28168) );
  XOR U27576 ( .A(n28172), .B(n28173), .Z(n28166) );
  AND U27577 ( .A(n1568), .B(n28165), .Z(n28173) );
  XNOR U27578 ( .A(n28163), .B(n28172), .Z(n28165) );
  XNOR U27579 ( .A(n28174), .B(n28175), .Z(n28163) );
  AND U27580 ( .A(n1572), .B(n28176), .Z(n28175) );
  XOR U27581 ( .A(p_input[1264]), .B(n28174), .Z(n28176) );
  XNOR U27582 ( .A(n28177), .B(n28178), .Z(n28174) );
  AND U27583 ( .A(n1576), .B(n28179), .Z(n28178) );
  XOR U27584 ( .A(n28180), .B(n28181), .Z(n28172) );
  AND U27585 ( .A(n1580), .B(n28171), .Z(n28181) );
  XNOR U27586 ( .A(n28182), .B(n28169), .Z(n28171) );
  XOR U27587 ( .A(n28183), .B(n28184), .Z(n28169) );
  AND U27588 ( .A(n1603), .B(n28185), .Z(n28184) );
  IV U27589 ( .A(n28180), .Z(n28182) );
  XOR U27590 ( .A(n28186), .B(n28187), .Z(n28180) );
  AND U27591 ( .A(n1587), .B(n28179), .Z(n28187) );
  XNOR U27592 ( .A(n28177), .B(n28186), .Z(n28179) );
  XNOR U27593 ( .A(n28188), .B(n28189), .Z(n28177) );
  AND U27594 ( .A(n1591), .B(n28190), .Z(n28189) );
  XOR U27595 ( .A(p_input[1280]), .B(n28188), .Z(n28190) );
  XNOR U27596 ( .A(n28191), .B(n28192), .Z(n28188) );
  AND U27597 ( .A(n1595), .B(n28193), .Z(n28192) );
  XOR U27598 ( .A(n28194), .B(n28195), .Z(n28186) );
  AND U27599 ( .A(n1599), .B(n28185), .Z(n28195) );
  XNOR U27600 ( .A(n28196), .B(n28183), .Z(n28185) );
  XOR U27601 ( .A(n28197), .B(n28198), .Z(n28183) );
  AND U27602 ( .A(n1622), .B(n28199), .Z(n28198) );
  IV U27603 ( .A(n28194), .Z(n28196) );
  XOR U27604 ( .A(n28200), .B(n28201), .Z(n28194) );
  AND U27605 ( .A(n1606), .B(n28193), .Z(n28201) );
  XNOR U27606 ( .A(n28191), .B(n28200), .Z(n28193) );
  XNOR U27607 ( .A(n28202), .B(n28203), .Z(n28191) );
  AND U27608 ( .A(n1610), .B(n28204), .Z(n28203) );
  XOR U27609 ( .A(p_input[1296]), .B(n28202), .Z(n28204) );
  XNOR U27610 ( .A(n28205), .B(n28206), .Z(n28202) );
  AND U27611 ( .A(n1614), .B(n28207), .Z(n28206) );
  XOR U27612 ( .A(n28208), .B(n28209), .Z(n28200) );
  AND U27613 ( .A(n1618), .B(n28199), .Z(n28209) );
  XNOR U27614 ( .A(n28210), .B(n28197), .Z(n28199) );
  XOR U27615 ( .A(n28211), .B(n28212), .Z(n28197) );
  AND U27616 ( .A(n1641), .B(n28213), .Z(n28212) );
  IV U27617 ( .A(n28208), .Z(n28210) );
  XOR U27618 ( .A(n28214), .B(n28215), .Z(n28208) );
  AND U27619 ( .A(n1625), .B(n28207), .Z(n28215) );
  XNOR U27620 ( .A(n28205), .B(n28214), .Z(n28207) );
  XNOR U27621 ( .A(n28216), .B(n28217), .Z(n28205) );
  AND U27622 ( .A(n1629), .B(n28218), .Z(n28217) );
  XOR U27623 ( .A(p_input[1312]), .B(n28216), .Z(n28218) );
  XNOR U27624 ( .A(n28219), .B(n28220), .Z(n28216) );
  AND U27625 ( .A(n1633), .B(n28221), .Z(n28220) );
  XOR U27626 ( .A(n28222), .B(n28223), .Z(n28214) );
  AND U27627 ( .A(n1637), .B(n28213), .Z(n28223) );
  XNOR U27628 ( .A(n28224), .B(n28211), .Z(n28213) );
  XOR U27629 ( .A(n28225), .B(n28226), .Z(n28211) );
  AND U27630 ( .A(n1660), .B(n28227), .Z(n28226) );
  IV U27631 ( .A(n28222), .Z(n28224) );
  XOR U27632 ( .A(n28228), .B(n28229), .Z(n28222) );
  AND U27633 ( .A(n1644), .B(n28221), .Z(n28229) );
  XNOR U27634 ( .A(n28219), .B(n28228), .Z(n28221) );
  XNOR U27635 ( .A(n28230), .B(n28231), .Z(n28219) );
  AND U27636 ( .A(n1648), .B(n28232), .Z(n28231) );
  XOR U27637 ( .A(p_input[1328]), .B(n28230), .Z(n28232) );
  XNOR U27638 ( .A(n28233), .B(n28234), .Z(n28230) );
  AND U27639 ( .A(n1652), .B(n28235), .Z(n28234) );
  XOR U27640 ( .A(n28236), .B(n28237), .Z(n28228) );
  AND U27641 ( .A(n1656), .B(n28227), .Z(n28237) );
  XNOR U27642 ( .A(n28238), .B(n28225), .Z(n28227) );
  XOR U27643 ( .A(n28239), .B(n28240), .Z(n28225) );
  AND U27644 ( .A(n1679), .B(n28241), .Z(n28240) );
  IV U27645 ( .A(n28236), .Z(n28238) );
  XOR U27646 ( .A(n28242), .B(n28243), .Z(n28236) );
  AND U27647 ( .A(n1663), .B(n28235), .Z(n28243) );
  XNOR U27648 ( .A(n28233), .B(n28242), .Z(n28235) );
  XNOR U27649 ( .A(n28244), .B(n28245), .Z(n28233) );
  AND U27650 ( .A(n1667), .B(n28246), .Z(n28245) );
  XOR U27651 ( .A(p_input[1344]), .B(n28244), .Z(n28246) );
  XNOR U27652 ( .A(n28247), .B(n28248), .Z(n28244) );
  AND U27653 ( .A(n1671), .B(n28249), .Z(n28248) );
  XOR U27654 ( .A(n28250), .B(n28251), .Z(n28242) );
  AND U27655 ( .A(n1675), .B(n28241), .Z(n28251) );
  XNOR U27656 ( .A(n28252), .B(n28239), .Z(n28241) );
  XOR U27657 ( .A(n28253), .B(n28254), .Z(n28239) );
  AND U27658 ( .A(n1698), .B(n28255), .Z(n28254) );
  IV U27659 ( .A(n28250), .Z(n28252) );
  XOR U27660 ( .A(n28256), .B(n28257), .Z(n28250) );
  AND U27661 ( .A(n1682), .B(n28249), .Z(n28257) );
  XNOR U27662 ( .A(n28247), .B(n28256), .Z(n28249) );
  XNOR U27663 ( .A(n28258), .B(n28259), .Z(n28247) );
  AND U27664 ( .A(n1686), .B(n28260), .Z(n28259) );
  XOR U27665 ( .A(p_input[1360]), .B(n28258), .Z(n28260) );
  XNOR U27666 ( .A(n28261), .B(n28262), .Z(n28258) );
  AND U27667 ( .A(n1690), .B(n28263), .Z(n28262) );
  XOR U27668 ( .A(n28264), .B(n28265), .Z(n28256) );
  AND U27669 ( .A(n1694), .B(n28255), .Z(n28265) );
  XNOR U27670 ( .A(n28266), .B(n28253), .Z(n28255) );
  XOR U27671 ( .A(n28267), .B(n28268), .Z(n28253) );
  AND U27672 ( .A(n1717), .B(n28269), .Z(n28268) );
  IV U27673 ( .A(n28264), .Z(n28266) );
  XOR U27674 ( .A(n28270), .B(n28271), .Z(n28264) );
  AND U27675 ( .A(n1701), .B(n28263), .Z(n28271) );
  XNOR U27676 ( .A(n28261), .B(n28270), .Z(n28263) );
  XNOR U27677 ( .A(n28272), .B(n28273), .Z(n28261) );
  AND U27678 ( .A(n1705), .B(n28274), .Z(n28273) );
  XOR U27679 ( .A(p_input[1376]), .B(n28272), .Z(n28274) );
  XNOR U27680 ( .A(n28275), .B(n28276), .Z(n28272) );
  AND U27681 ( .A(n1709), .B(n28277), .Z(n28276) );
  XOR U27682 ( .A(n28278), .B(n28279), .Z(n28270) );
  AND U27683 ( .A(n1713), .B(n28269), .Z(n28279) );
  XNOR U27684 ( .A(n28280), .B(n28267), .Z(n28269) );
  XOR U27685 ( .A(n28281), .B(n28282), .Z(n28267) );
  AND U27686 ( .A(n1736), .B(n28283), .Z(n28282) );
  IV U27687 ( .A(n28278), .Z(n28280) );
  XOR U27688 ( .A(n28284), .B(n28285), .Z(n28278) );
  AND U27689 ( .A(n1720), .B(n28277), .Z(n28285) );
  XNOR U27690 ( .A(n28275), .B(n28284), .Z(n28277) );
  XNOR U27691 ( .A(n28286), .B(n28287), .Z(n28275) );
  AND U27692 ( .A(n1724), .B(n28288), .Z(n28287) );
  XOR U27693 ( .A(p_input[1392]), .B(n28286), .Z(n28288) );
  XNOR U27694 ( .A(n28289), .B(n28290), .Z(n28286) );
  AND U27695 ( .A(n1728), .B(n28291), .Z(n28290) );
  XOR U27696 ( .A(n28292), .B(n28293), .Z(n28284) );
  AND U27697 ( .A(n1732), .B(n28283), .Z(n28293) );
  XNOR U27698 ( .A(n28294), .B(n28281), .Z(n28283) );
  XOR U27699 ( .A(n28295), .B(n28296), .Z(n28281) );
  AND U27700 ( .A(n1755), .B(n28297), .Z(n28296) );
  IV U27701 ( .A(n28292), .Z(n28294) );
  XOR U27702 ( .A(n28298), .B(n28299), .Z(n28292) );
  AND U27703 ( .A(n1739), .B(n28291), .Z(n28299) );
  XNOR U27704 ( .A(n28289), .B(n28298), .Z(n28291) );
  XNOR U27705 ( .A(n28300), .B(n28301), .Z(n28289) );
  AND U27706 ( .A(n1743), .B(n28302), .Z(n28301) );
  XOR U27707 ( .A(p_input[1408]), .B(n28300), .Z(n28302) );
  XNOR U27708 ( .A(n28303), .B(n28304), .Z(n28300) );
  AND U27709 ( .A(n1747), .B(n28305), .Z(n28304) );
  XOR U27710 ( .A(n28306), .B(n28307), .Z(n28298) );
  AND U27711 ( .A(n1751), .B(n28297), .Z(n28307) );
  XNOR U27712 ( .A(n28308), .B(n28295), .Z(n28297) );
  XOR U27713 ( .A(n28309), .B(n28310), .Z(n28295) );
  AND U27714 ( .A(n1774), .B(n28311), .Z(n28310) );
  IV U27715 ( .A(n28306), .Z(n28308) );
  XOR U27716 ( .A(n28312), .B(n28313), .Z(n28306) );
  AND U27717 ( .A(n1758), .B(n28305), .Z(n28313) );
  XNOR U27718 ( .A(n28303), .B(n28312), .Z(n28305) );
  XNOR U27719 ( .A(n28314), .B(n28315), .Z(n28303) );
  AND U27720 ( .A(n1762), .B(n28316), .Z(n28315) );
  XOR U27721 ( .A(p_input[1424]), .B(n28314), .Z(n28316) );
  XNOR U27722 ( .A(n28317), .B(n28318), .Z(n28314) );
  AND U27723 ( .A(n1766), .B(n28319), .Z(n28318) );
  XOR U27724 ( .A(n28320), .B(n28321), .Z(n28312) );
  AND U27725 ( .A(n1770), .B(n28311), .Z(n28321) );
  XNOR U27726 ( .A(n28322), .B(n28309), .Z(n28311) );
  XOR U27727 ( .A(n28323), .B(n28324), .Z(n28309) );
  AND U27728 ( .A(n1793), .B(n28325), .Z(n28324) );
  IV U27729 ( .A(n28320), .Z(n28322) );
  XOR U27730 ( .A(n28326), .B(n28327), .Z(n28320) );
  AND U27731 ( .A(n1777), .B(n28319), .Z(n28327) );
  XNOR U27732 ( .A(n28317), .B(n28326), .Z(n28319) );
  XNOR U27733 ( .A(n28328), .B(n28329), .Z(n28317) );
  AND U27734 ( .A(n1781), .B(n28330), .Z(n28329) );
  XOR U27735 ( .A(p_input[1440]), .B(n28328), .Z(n28330) );
  XNOR U27736 ( .A(n28331), .B(n28332), .Z(n28328) );
  AND U27737 ( .A(n1785), .B(n28333), .Z(n28332) );
  XOR U27738 ( .A(n28334), .B(n28335), .Z(n28326) );
  AND U27739 ( .A(n1789), .B(n28325), .Z(n28335) );
  XNOR U27740 ( .A(n28336), .B(n28323), .Z(n28325) );
  XOR U27741 ( .A(n28337), .B(n28338), .Z(n28323) );
  AND U27742 ( .A(n1812), .B(n28339), .Z(n28338) );
  IV U27743 ( .A(n28334), .Z(n28336) );
  XOR U27744 ( .A(n28340), .B(n28341), .Z(n28334) );
  AND U27745 ( .A(n1796), .B(n28333), .Z(n28341) );
  XNOR U27746 ( .A(n28331), .B(n28340), .Z(n28333) );
  XNOR U27747 ( .A(n28342), .B(n28343), .Z(n28331) );
  AND U27748 ( .A(n1800), .B(n28344), .Z(n28343) );
  XOR U27749 ( .A(p_input[1456]), .B(n28342), .Z(n28344) );
  XNOR U27750 ( .A(n28345), .B(n28346), .Z(n28342) );
  AND U27751 ( .A(n1804), .B(n28347), .Z(n28346) );
  XOR U27752 ( .A(n28348), .B(n28349), .Z(n28340) );
  AND U27753 ( .A(n1808), .B(n28339), .Z(n28349) );
  XNOR U27754 ( .A(n28350), .B(n28337), .Z(n28339) );
  XOR U27755 ( .A(n28351), .B(n28352), .Z(n28337) );
  AND U27756 ( .A(n1831), .B(n28353), .Z(n28352) );
  IV U27757 ( .A(n28348), .Z(n28350) );
  XOR U27758 ( .A(n28354), .B(n28355), .Z(n28348) );
  AND U27759 ( .A(n1815), .B(n28347), .Z(n28355) );
  XNOR U27760 ( .A(n28345), .B(n28354), .Z(n28347) );
  XNOR U27761 ( .A(n28356), .B(n28357), .Z(n28345) );
  AND U27762 ( .A(n1819), .B(n28358), .Z(n28357) );
  XOR U27763 ( .A(p_input[1472]), .B(n28356), .Z(n28358) );
  XNOR U27764 ( .A(n28359), .B(n28360), .Z(n28356) );
  AND U27765 ( .A(n1823), .B(n28361), .Z(n28360) );
  XOR U27766 ( .A(n28362), .B(n28363), .Z(n28354) );
  AND U27767 ( .A(n1827), .B(n28353), .Z(n28363) );
  XNOR U27768 ( .A(n28364), .B(n28351), .Z(n28353) );
  XOR U27769 ( .A(n28365), .B(n28366), .Z(n28351) );
  AND U27770 ( .A(n1850), .B(n28367), .Z(n28366) );
  IV U27771 ( .A(n28362), .Z(n28364) );
  XOR U27772 ( .A(n28368), .B(n28369), .Z(n28362) );
  AND U27773 ( .A(n1834), .B(n28361), .Z(n28369) );
  XNOR U27774 ( .A(n28359), .B(n28368), .Z(n28361) );
  XNOR U27775 ( .A(n28370), .B(n28371), .Z(n28359) );
  AND U27776 ( .A(n1838), .B(n28372), .Z(n28371) );
  XOR U27777 ( .A(p_input[1488]), .B(n28370), .Z(n28372) );
  XNOR U27778 ( .A(n28373), .B(n28374), .Z(n28370) );
  AND U27779 ( .A(n1842), .B(n28375), .Z(n28374) );
  XOR U27780 ( .A(n28376), .B(n28377), .Z(n28368) );
  AND U27781 ( .A(n1846), .B(n28367), .Z(n28377) );
  XNOR U27782 ( .A(n28378), .B(n28365), .Z(n28367) );
  XOR U27783 ( .A(n28379), .B(n28380), .Z(n28365) );
  AND U27784 ( .A(n1869), .B(n28381), .Z(n28380) );
  IV U27785 ( .A(n28376), .Z(n28378) );
  XOR U27786 ( .A(n28382), .B(n28383), .Z(n28376) );
  AND U27787 ( .A(n1853), .B(n28375), .Z(n28383) );
  XNOR U27788 ( .A(n28373), .B(n28382), .Z(n28375) );
  XNOR U27789 ( .A(n28384), .B(n28385), .Z(n28373) );
  AND U27790 ( .A(n1857), .B(n28386), .Z(n28385) );
  XOR U27791 ( .A(p_input[1504]), .B(n28384), .Z(n28386) );
  XNOR U27792 ( .A(n28387), .B(n28388), .Z(n28384) );
  AND U27793 ( .A(n1861), .B(n28389), .Z(n28388) );
  XOR U27794 ( .A(n28390), .B(n28391), .Z(n28382) );
  AND U27795 ( .A(n1865), .B(n28381), .Z(n28391) );
  XNOR U27796 ( .A(n28392), .B(n28379), .Z(n28381) );
  XOR U27797 ( .A(n28393), .B(n28394), .Z(n28379) );
  AND U27798 ( .A(n1888), .B(n28395), .Z(n28394) );
  IV U27799 ( .A(n28390), .Z(n28392) );
  XOR U27800 ( .A(n28396), .B(n28397), .Z(n28390) );
  AND U27801 ( .A(n1872), .B(n28389), .Z(n28397) );
  XNOR U27802 ( .A(n28387), .B(n28396), .Z(n28389) );
  XNOR U27803 ( .A(n28398), .B(n28399), .Z(n28387) );
  AND U27804 ( .A(n1876), .B(n28400), .Z(n28399) );
  XOR U27805 ( .A(p_input[1520]), .B(n28398), .Z(n28400) );
  XNOR U27806 ( .A(n28401), .B(n28402), .Z(n28398) );
  AND U27807 ( .A(n1880), .B(n28403), .Z(n28402) );
  XOR U27808 ( .A(n28404), .B(n28405), .Z(n28396) );
  AND U27809 ( .A(n1884), .B(n28395), .Z(n28405) );
  XNOR U27810 ( .A(n28406), .B(n28393), .Z(n28395) );
  XOR U27811 ( .A(n28407), .B(n28408), .Z(n28393) );
  AND U27812 ( .A(n1907), .B(n28409), .Z(n28408) );
  IV U27813 ( .A(n28404), .Z(n28406) );
  XOR U27814 ( .A(n28410), .B(n28411), .Z(n28404) );
  AND U27815 ( .A(n1891), .B(n28403), .Z(n28411) );
  XNOR U27816 ( .A(n28401), .B(n28410), .Z(n28403) );
  XNOR U27817 ( .A(n28412), .B(n28413), .Z(n28401) );
  AND U27818 ( .A(n1895), .B(n28414), .Z(n28413) );
  XOR U27819 ( .A(p_input[1536]), .B(n28412), .Z(n28414) );
  XNOR U27820 ( .A(n28415), .B(n28416), .Z(n28412) );
  AND U27821 ( .A(n1899), .B(n28417), .Z(n28416) );
  XOR U27822 ( .A(n28418), .B(n28419), .Z(n28410) );
  AND U27823 ( .A(n1903), .B(n28409), .Z(n28419) );
  XNOR U27824 ( .A(n28420), .B(n28407), .Z(n28409) );
  XOR U27825 ( .A(n28421), .B(n28422), .Z(n28407) );
  AND U27826 ( .A(n1926), .B(n28423), .Z(n28422) );
  IV U27827 ( .A(n28418), .Z(n28420) );
  XOR U27828 ( .A(n28424), .B(n28425), .Z(n28418) );
  AND U27829 ( .A(n1910), .B(n28417), .Z(n28425) );
  XNOR U27830 ( .A(n28415), .B(n28424), .Z(n28417) );
  XNOR U27831 ( .A(n28426), .B(n28427), .Z(n28415) );
  AND U27832 ( .A(n1914), .B(n28428), .Z(n28427) );
  XOR U27833 ( .A(p_input[1552]), .B(n28426), .Z(n28428) );
  XNOR U27834 ( .A(n28429), .B(n28430), .Z(n28426) );
  AND U27835 ( .A(n1918), .B(n28431), .Z(n28430) );
  XOR U27836 ( .A(n28432), .B(n28433), .Z(n28424) );
  AND U27837 ( .A(n1922), .B(n28423), .Z(n28433) );
  XNOR U27838 ( .A(n28434), .B(n28421), .Z(n28423) );
  XOR U27839 ( .A(n28435), .B(n28436), .Z(n28421) );
  AND U27840 ( .A(n1945), .B(n28437), .Z(n28436) );
  IV U27841 ( .A(n28432), .Z(n28434) );
  XOR U27842 ( .A(n28438), .B(n28439), .Z(n28432) );
  AND U27843 ( .A(n1929), .B(n28431), .Z(n28439) );
  XNOR U27844 ( .A(n28429), .B(n28438), .Z(n28431) );
  XNOR U27845 ( .A(n28440), .B(n28441), .Z(n28429) );
  AND U27846 ( .A(n1933), .B(n28442), .Z(n28441) );
  XOR U27847 ( .A(p_input[1568]), .B(n28440), .Z(n28442) );
  XNOR U27848 ( .A(n28443), .B(n28444), .Z(n28440) );
  AND U27849 ( .A(n1937), .B(n28445), .Z(n28444) );
  XOR U27850 ( .A(n28446), .B(n28447), .Z(n28438) );
  AND U27851 ( .A(n1941), .B(n28437), .Z(n28447) );
  XNOR U27852 ( .A(n28448), .B(n28435), .Z(n28437) );
  XOR U27853 ( .A(n28449), .B(n28450), .Z(n28435) );
  AND U27854 ( .A(n1964), .B(n28451), .Z(n28450) );
  IV U27855 ( .A(n28446), .Z(n28448) );
  XOR U27856 ( .A(n28452), .B(n28453), .Z(n28446) );
  AND U27857 ( .A(n1948), .B(n28445), .Z(n28453) );
  XNOR U27858 ( .A(n28443), .B(n28452), .Z(n28445) );
  XNOR U27859 ( .A(n28454), .B(n28455), .Z(n28443) );
  AND U27860 ( .A(n1952), .B(n28456), .Z(n28455) );
  XOR U27861 ( .A(p_input[1584]), .B(n28454), .Z(n28456) );
  XNOR U27862 ( .A(n28457), .B(n28458), .Z(n28454) );
  AND U27863 ( .A(n1956), .B(n28459), .Z(n28458) );
  XOR U27864 ( .A(n28460), .B(n28461), .Z(n28452) );
  AND U27865 ( .A(n1960), .B(n28451), .Z(n28461) );
  XNOR U27866 ( .A(n28462), .B(n28449), .Z(n28451) );
  XOR U27867 ( .A(n28463), .B(n28464), .Z(n28449) );
  AND U27868 ( .A(n1983), .B(n28465), .Z(n28464) );
  IV U27869 ( .A(n28460), .Z(n28462) );
  XOR U27870 ( .A(n28466), .B(n28467), .Z(n28460) );
  AND U27871 ( .A(n1967), .B(n28459), .Z(n28467) );
  XNOR U27872 ( .A(n28457), .B(n28466), .Z(n28459) );
  XNOR U27873 ( .A(n28468), .B(n28469), .Z(n28457) );
  AND U27874 ( .A(n1971), .B(n28470), .Z(n28469) );
  XOR U27875 ( .A(p_input[1600]), .B(n28468), .Z(n28470) );
  XNOR U27876 ( .A(n28471), .B(n28472), .Z(n28468) );
  AND U27877 ( .A(n1975), .B(n28473), .Z(n28472) );
  XOR U27878 ( .A(n28474), .B(n28475), .Z(n28466) );
  AND U27879 ( .A(n1979), .B(n28465), .Z(n28475) );
  XNOR U27880 ( .A(n28476), .B(n28463), .Z(n28465) );
  XOR U27881 ( .A(n28477), .B(n28478), .Z(n28463) );
  AND U27882 ( .A(n2002), .B(n28479), .Z(n28478) );
  IV U27883 ( .A(n28474), .Z(n28476) );
  XOR U27884 ( .A(n28480), .B(n28481), .Z(n28474) );
  AND U27885 ( .A(n1986), .B(n28473), .Z(n28481) );
  XNOR U27886 ( .A(n28471), .B(n28480), .Z(n28473) );
  XNOR U27887 ( .A(n28482), .B(n28483), .Z(n28471) );
  AND U27888 ( .A(n1990), .B(n28484), .Z(n28483) );
  XOR U27889 ( .A(p_input[1616]), .B(n28482), .Z(n28484) );
  XNOR U27890 ( .A(n28485), .B(n28486), .Z(n28482) );
  AND U27891 ( .A(n1994), .B(n28487), .Z(n28486) );
  XOR U27892 ( .A(n28488), .B(n28489), .Z(n28480) );
  AND U27893 ( .A(n1998), .B(n28479), .Z(n28489) );
  XNOR U27894 ( .A(n28490), .B(n28477), .Z(n28479) );
  XOR U27895 ( .A(n28491), .B(n28492), .Z(n28477) );
  AND U27896 ( .A(n2021), .B(n28493), .Z(n28492) );
  IV U27897 ( .A(n28488), .Z(n28490) );
  XOR U27898 ( .A(n28494), .B(n28495), .Z(n28488) );
  AND U27899 ( .A(n2005), .B(n28487), .Z(n28495) );
  XNOR U27900 ( .A(n28485), .B(n28494), .Z(n28487) );
  XNOR U27901 ( .A(n28496), .B(n28497), .Z(n28485) );
  AND U27902 ( .A(n2009), .B(n28498), .Z(n28497) );
  XOR U27903 ( .A(p_input[1632]), .B(n28496), .Z(n28498) );
  XNOR U27904 ( .A(n28499), .B(n28500), .Z(n28496) );
  AND U27905 ( .A(n2013), .B(n28501), .Z(n28500) );
  XOR U27906 ( .A(n28502), .B(n28503), .Z(n28494) );
  AND U27907 ( .A(n2017), .B(n28493), .Z(n28503) );
  XNOR U27908 ( .A(n28504), .B(n28491), .Z(n28493) );
  XOR U27909 ( .A(n28505), .B(n28506), .Z(n28491) );
  AND U27910 ( .A(n2040), .B(n28507), .Z(n28506) );
  IV U27911 ( .A(n28502), .Z(n28504) );
  XOR U27912 ( .A(n28508), .B(n28509), .Z(n28502) );
  AND U27913 ( .A(n2024), .B(n28501), .Z(n28509) );
  XNOR U27914 ( .A(n28499), .B(n28508), .Z(n28501) );
  XNOR U27915 ( .A(n28510), .B(n28511), .Z(n28499) );
  AND U27916 ( .A(n2028), .B(n28512), .Z(n28511) );
  XOR U27917 ( .A(p_input[1648]), .B(n28510), .Z(n28512) );
  XNOR U27918 ( .A(n28513), .B(n28514), .Z(n28510) );
  AND U27919 ( .A(n2032), .B(n28515), .Z(n28514) );
  XOR U27920 ( .A(n28516), .B(n28517), .Z(n28508) );
  AND U27921 ( .A(n2036), .B(n28507), .Z(n28517) );
  XNOR U27922 ( .A(n28518), .B(n28505), .Z(n28507) );
  XOR U27923 ( .A(n28519), .B(n28520), .Z(n28505) );
  AND U27924 ( .A(n2059), .B(n28521), .Z(n28520) );
  IV U27925 ( .A(n28516), .Z(n28518) );
  XOR U27926 ( .A(n28522), .B(n28523), .Z(n28516) );
  AND U27927 ( .A(n2043), .B(n28515), .Z(n28523) );
  XNOR U27928 ( .A(n28513), .B(n28522), .Z(n28515) );
  XNOR U27929 ( .A(n28524), .B(n28525), .Z(n28513) );
  AND U27930 ( .A(n2047), .B(n28526), .Z(n28525) );
  XOR U27931 ( .A(p_input[1664]), .B(n28524), .Z(n28526) );
  XNOR U27932 ( .A(n28527), .B(n28528), .Z(n28524) );
  AND U27933 ( .A(n2051), .B(n28529), .Z(n28528) );
  XOR U27934 ( .A(n28530), .B(n28531), .Z(n28522) );
  AND U27935 ( .A(n2055), .B(n28521), .Z(n28531) );
  XNOR U27936 ( .A(n28532), .B(n28519), .Z(n28521) );
  XOR U27937 ( .A(n28533), .B(n28534), .Z(n28519) );
  AND U27938 ( .A(n2078), .B(n28535), .Z(n28534) );
  IV U27939 ( .A(n28530), .Z(n28532) );
  XOR U27940 ( .A(n28536), .B(n28537), .Z(n28530) );
  AND U27941 ( .A(n2062), .B(n28529), .Z(n28537) );
  XNOR U27942 ( .A(n28527), .B(n28536), .Z(n28529) );
  XNOR U27943 ( .A(n28538), .B(n28539), .Z(n28527) );
  AND U27944 ( .A(n2066), .B(n28540), .Z(n28539) );
  XOR U27945 ( .A(p_input[1680]), .B(n28538), .Z(n28540) );
  XNOR U27946 ( .A(n28541), .B(n28542), .Z(n28538) );
  AND U27947 ( .A(n2070), .B(n28543), .Z(n28542) );
  XOR U27948 ( .A(n28544), .B(n28545), .Z(n28536) );
  AND U27949 ( .A(n2074), .B(n28535), .Z(n28545) );
  XNOR U27950 ( .A(n28546), .B(n28533), .Z(n28535) );
  XOR U27951 ( .A(n28547), .B(n28548), .Z(n28533) );
  AND U27952 ( .A(n2097), .B(n28549), .Z(n28548) );
  IV U27953 ( .A(n28544), .Z(n28546) );
  XOR U27954 ( .A(n28550), .B(n28551), .Z(n28544) );
  AND U27955 ( .A(n2081), .B(n28543), .Z(n28551) );
  XNOR U27956 ( .A(n28541), .B(n28550), .Z(n28543) );
  XNOR U27957 ( .A(n28552), .B(n28553), .Z(n28541) );
  AND U27958 ( .A(n2085), .B(n28554), .Z(n28553) );
  XOR U27959 ( .A(p_input[1696]), .B(n28552), .Z(n28554) );
  XNOR U27960 ( .A(n28555), .B(n28556), .Z(n28552) );
  AND U27961 ( .A(n2089), .B(n28557), .Z(n28556) );
  XOR U27962 ( .A(n28558), .B(n28559), .Z(n28550) );
  AND U27963 ( .A(n2093), .B(n28549), .Z(n28559) );
  XNOR U27964 ( .A(n28560), .B(n28547), .Z(n28549) );
  XOR U27965 ( .A(n28561), .B(n28562), .Z(n28547) );
  AND U27966 ( .A(n2116), .B(n28563), .Z(n28562) );
  IV U27967 ( .A(n28558), .Z(n28560) );
  XOR U27968 ( .A(n28564), .B(n28565), .Z(n28558) );
  AND U27969 ( .A(n2100), .B(n28557), .Z(n28565) );
  XNOR U27970 ( .A(n28555), .B(n28564), .Z(n28557) );
  XNOR U27971 ( .A(n28566), .B(n28567), .Z(n28555) );
  AND U27972 ( .A(n2104), .B(n28568), .Z(n28567) );
  XOR U27973 ( .A(p_input[1712]), .B(n28566), .Z(n28568) );
  XNOR U27974 ( .A(n28569), .B(n28570), .Z(n28566) );
  AND U27975 ( .A(n2108), .B(n28571), .Z(n28570) );
  XOR U27976 ( .A(n28572), .B(n28573), .Z(n28564) );
  AND U27977 ( .A(n2112), .B(n28563), .Z(n28573) );
  XNOR U27978 ( .A(n28574), .B(n28561), .Z(n28563) );
  XOR U27979 ( .A(n28575), .B(n28576), .Z(n28561) );
  AND U27980 ( .A(n2135), .B(n28577), .Z(n28576) );
  IV U27981 ( .A(n28572), .Z(n28574) );
  XOR U27982 ( .A(n28578), .B(n28579), .Z(n28572) );
  AND U27983 ( .A(n2119), .B(n28571), .Z(n28579) );
  XNOR U27984 ( .A(n28569), .B(n28578), .Z(n28571) );
  XNOR U27985 ( .A(n28580), .B(n28581), .Z(n28569) );
  AND U27986 ( .A(n2123), .B(n28582), .Z(n28581) );
  XOR U27987 ( .A(p_input[1728]), .B(n28580), .Z(n28582) );
  XNOR U27988 ( .A(n28583), .B(n28584), .Z(n28580) );
  AND U27989 ( .A(n2127), .B(n28585), .Z(n28584) );
  XOR U27990 ( .A(n28586), .B(n28587), .Z(n28578) );
  AND U27991 ( .A(n2131), .B(n28577), .Z(n28587) );
  XNOR U27992 ( .A(n28588), .B(n28575), .Z(n28577) );
  XOR U27993 ( .A(n28589), .B(n28590), .Z(n28575) );
  AND U27994 ( .A(n2154), .B(n28591), .Z(n28590) );
  IV U27995 ( .A(n28586), .Z(n28588) );
  XOR U27996 ( .A(n28592), .B(n28593), .Z(n28586) );
  AND U27997 ( .A(n2138), .B(n28585), .Z(n28593) );
  XNOR U27998 ( .A(n28583), .B(n28592), .Z(n28585) );
  XNOR U27999 ( .A(n28594), .B(n28595), .Z(n28583) );
  AND U28000 ( .A(n2142), .B(n28596), .Z(n28595) );
  XOR U28001 ( .A(p_input[1744]), .B(n28594), .Z(n28596) );
  XNOR U28002 ( .A(n28597), .B(n28598), .Z(n28594) );
  AND U28003 ( .A(n2146), .B(n28599), .Z(n28598) );
  XOR U28004 ( .A(n28600), .B(n28601), .Z(n28592) );
  AND U28005 ( .A(n2150), .B(n28591), .Z(n28601) );
  XNOR U28006 ( .A(n28602), .B(n28589), .Z(n28591) );
  XOR U28007 ( .A(n28603), .B(n28604), .Z(n28589) );
  AND U28008 ( .A(n2173), .B(n28605), .Z(n28604) );
  IV U28009 ( .A(n28600), .Z(n28602) );
  XOR U28010 ( .A(n28606), .B(n28607), .Z(n28600) );
  AND U28011 ( .A(n2157), .B(n28599), .Z(n28607) );
  XNOR U28012 ( .A(n28597), .B(n28606), .Z(n28599) );
  XNOR U28013 ( .A(n28608), .B(n28609), .Z(n28597) );
  AND U28014 ( .A(n2161), .B(n28610), .Z(n28609) );
  XOR U28015 ( .A(p_input[1760]), .B(n28608), .Z(n28610) );
  XNOR U28016 ( .A(n28611), .B(n28612), .Z(n28608) );
  AND U28017 ( .A(n2165), .B(n28613), .Z(n28612) );
  XOR U28018 ( .A(n28614), .B(n28615), .Z(n28606) );
  AND U28019 ( .A(n2169), .B(n28605), .Z(n28615) );
  XNOR U28020 ( .A(n28616), .B(n28603), .Z(n28605) );
  XOR U28021 ( .A(n28617), .B(n28618), .Z(n28603) );
  AND U28022 ( .A(n2192), .B(n28619), .Z(n28618) );
  IV U28023 ( .A(n28614), .Z(n28616) );
  XOR U28024 ( .A(n28620), .B(n28621), .Z(n28614) );
  AND U28025 ( .A(n2176), .B(n28613), .Z(n28621) );
  XNOR U28026 ( .A(n28611), .B(n28620), .Z(n28613) );
  XNOR U28027 ( .A(n28622), .B(n28623), .Z(n28611) );
  AND U28028 ( .A(n2180), .B(n28624), .Z(n28623) );
  XOR U28029 ( .A(p_input[1776]), .B(n28622), .Z(n28624) );
  XNOR U28030 ( .A(n28625), .B(n28626), .Z(n28622) );
  AND U28031 ( .A(n2184), .B(n28627), .Z(n28626) );
  XOR U28032 ( .A(n28628), .B(n28629), .Z(n28620) );
  AND U28033 ( .A(n2188), .B(n28619), .Z(n28629) );
  XNOR U28034 ( .A(n28630), .B(n28617), .Z(n28619) );
  XOR U28035 ( .A(n28631), .B(n28632), .Z(n28617) );
  AND U28036 ( .A(n2211), .B(n28633), .Z(n28632) );
  IV U28037 ( .A(n28628), .Z(n28630) );
  XOR U28038 ( .A(n28634), .B(n28635), .Z(n28628) );
  AND U28039 ( .A(n2195), .B(n28627), .Z(n28635) );
  XNOR U28040 ( .A(n28625), .B(n28634), .Z(n28627) );
  XNOR U28041 ( .A(n28636), .B(n28637), .Z(n28625) );
  AND U28042 ( .A(n2199), .B(n28638), .Z(n28637) );
  XOR U28043 ( .A(p_input[1792]), .B(n28636), .Z(n28638) );
  XNOR U28044 ( .A(n28639), .B(n28640), .Z(n28636) );
  AND U28045 ( .A(n2203), .B(n28641), .Z(n28640) );
  XOR U28046 ( .A(n28642), .B(n28643), .Z(n28634) );
  AND U28047 ( .A(n2207), .B(n28633), .Z(n28643) );
  XNOR U28048 ( .A(n28644), .B(n28631), .Z(n28633) );
  XOR U28049 ( .A(n28645), .B(n28646), .Z(n28631) );
  AND U28050 ( .A(n2230), .B(n28647), .Z(n28646) );
  IV U28051 ( .A(n28642), .Z(n28644) );
  XOR U28052 ( .A(n28648), .B(n28649), .Z(n28642) );
  AND U28053 ( .A(n2214), .B(n28641), .Z(n28649) );
  XNOR U28054 ( .A(n28639), .B(n28648), .Z(n28641) );
  XNOR U28055 ( .A(n28650), .B(n28651), .Z(n28639) );
  AND U28056 ( .A(n2218), .B(n28652), .Z(n28651) );
  XOR U28057 ( .A(p_input[1808]), .B(n28650), .Z(n28652) );
  XNOR U28058 ( .A(n28653), .B(n28654), .Z(n28650) );
  AND U28059 ( .A(n2222), .B(n28655), .Z(n28654) );
  XOR U28060 ( .A(n28656), .B(n28657), .Z(n28648) );
  AND U28061 ( .A(n2226), .B(n28647), .Z(n28657) );
  XNOR U28062 ( .A(n28658), .B(n28645), .Z(n28647) );
  XOR U28063 ( .A(n28659), .B(n28660), .Z(n28645) );
  AND U28064 ( .A(n2249), .B(n28661), .Z(n28660) );
  IV U28065 ( .A(n28656), .Z(n28658) );
  XOR U28066 ( .A(n28662), .B(n28663), .Z(n28656) );
  AND U28067 ( .A(n2233), .B(n28655), .Z(n28663) );
  XNOR U28068 ( .A(n28653), .B(n28662), .Z(n28655) );
  XNOR U28069 ( .A(n28664), .B(n28665), .Z(n28653) );
  AND U28070 ( .A(n2237), .B(n28666), .Z(n28665) );
  XOR U28071 ( .A(p_input[1824]), .B(n28664), .Z(n28666) );
  XNOR U28072 ( .A(n28667), .B(n28668), .Z(n28664) );
  AND U28073 ( .A(n2241), .B(n28669), .Z(n28668) );
  XOR U28074 ( .A(n28670), .B(n28671), .Z(n28662) );
  AND U28075 ( .A(n2245), .B(n28661), .Z(n28671) );
  XNOR U28076 ( .A(n28672), .B(n28659), .Z(n28661) );
  XOR U28077 ( .A(n28673), .B(n28674), .Z(n28659) );
  AND U28078 ( .A(n2268), .B(n28675), .Z(n28674) );
  IV U28079 ( .A(n28670), .Z(n28672) );
  XOR U28080 ( .A(n28676), .B(n28677), .Z(n28670) );
  AND U28081 ( .A(n2252), .B(n28669), .Z(n28677) );
  XNOR U28082 ( .A(n28667), .B(n28676), .Z(n28669) );
  XNOR U28083 ( .A(n28678), .B(n28679), .Z(n28667) );
  AND U28084 ( .A(n2256), .B(n28680), .Z(n28679) );
  XOR U28085 ( .A(p_input[1840]), .B(n28678), .Z(n28680) );
  XNOR U28086 ( .A(n28681), .B(n28682), .Z(n28678) );
  AND U28087 ( .A(n2260), .B(n28683), .Z(n28682) );
  XOR U28088 ( .A(n28684), .B(n28685), .Z(n28676) );
  AND U28089 ( .A(n2264), .B(n28675), .Z(n28685) );
  XNOR U28090 ( .A(n28686), .B(n28673), .Z(n28675) );
  XOR U28091 ( .A(n28687), .B(n28688), .Z(n28673) );
  AND U28092 ( .A(n2287), .B(n28689), .Z(n28688) );
  IV U28093 ( .A(n28684), .Z(n28686) );
  XOR U28094 ( .A(n28690), .B(n28691), .Z(n28684) );
  AND U28095 ( .A(n2271), .B(n28683), .Z(n28691) );
  XNOR U28096 ( .A(n28681), .B(n28690), .Z(n28683) );
  XNOR U28097 ( .A(n28692), .B(n28693), .Z(n28681) );
  AND U28098 ( .A(n2275), .B(n28694), .Z(n28693) );
  XOR U28099 ( .A(p_input[1856]), .B(n28692), .Z(n28694) );
  XNOR U28100 ( .A(n28695), .B(n28696), .Z(n28692) );
  AND U28101 ( .A(n2279), .B(n28697), .Z(n28696) );
  XOR U28102 ( .A(n28698), .B(n28699), .Z(n28690) );
  AND U28103 ( .A(n2283), .B(n28689), .Z(n28699) );
  XNOR U28104 ( .A(n28700), .B(n28687), .Z(n28689) );
  XOR U28105 ( .A(n28701), .B(n28702), .Z(n28687) );
  AND U28106 ( .A(n2306), .B(n28703), .Z(n28702) );
  IV U28107 ( .A(n28698), .Z(n28700) );
  XOR U28108 ( .A(n28704), .B(n28705), .Z(n28698) );
  AND U28109 ( .A(n2290), .B(n28697), .Z(n28705) );
  XNOR U28110 ( .A(n28695), .B(n28704), .Z(n28697) );
  XNOR U28111 ( .A(n28706), .B(n28707), .Z(n28695) );
  AND U28112 ( .A(n2294), .B(n28708), .Z(n28707) );
  XOR U28113 ( .A(p_input[1872]), .B(n28706), .Z(n28708) );
  XNOR U28114 ( .A(n28709), .B(n28710), .Z(n28706) );
  AND U28115 ( .A(n2298), .B(n28711), .Z(n28710) );
  XOR U28116 ( .A(n28712), .B(n28713), .Z(n28704) );
  AND U28117 ( .A(n2302), .B(n28703), .Z(n28713) );
  XNOR U28118 ( .A(n28714), .B(n28701), .Z(n28703) );
  XOR U28119 ( .A(n28715), .B(n28716), .Z(n28701) );
  AND U28120 ( .A(n2325), .B(n28717), .Z(n28716) );
  IV U28121 ( .A(n28712), .Z(n28714) );
  XOR U28122 ( .A(n28718), .B(n28719), .Z(n28712) );
  AND U28123 ( .A(n2309), .B(n28711), .Z(n28719) );
  XNOR U28124 ( .A(n28709), .B(n28718), .Z(n28711) );
  XNOR U28125 ( .A(n28720), .B(n28721), .Z(n28709) );
  AND U28126 ( .A(n2313), .B(n28722), .Z(n28721) );
  XOR U28127 ( .A(p_input[1888]), .B(n28720), .Z(n28722) );
  XNOR U28128 ( .A(n28723), .B(n28724), .Z(n28720) );
  AND U28129 ( .A(n2317), .B(n28725), .Z(n28724) );
  XOR U28130 ( .A(n28726), .B(n28727), .Z(n28718) );
  AND U28131 ( .A(n2321), .B(n28717), .Z(n28727) );
  XNOR U28132 ( .A(n28728), .B(n28715), .Z(n28717) );
  XOR U28133 ( .A(n28729), .B(n28730), .Z(n28715) );
  AND U28134 ( .A(n2344), .B(n28731), .Z(n28730) );
  IV U28135 ( .A(n28726), .Z(n28728) );
  XOR U28136 ( .A(n28732), .B(n28733), .Z(n28726) );
  AND U28137 ( .A(n2328), .B(n28725), .Z(n28733) );
  XNOR U28138 ( .A(n28723), .B(n28732), .Z(n28725) );
  XNOR U28139 ( .A(n28734), .B(n28735), .Z(n28723) );
  AND U28140 ( .A(n2332), .B(n28736), .Z(n28735) );
  XOR U28141 ( .A(p_input[1904]), .B(n28734), .Z(n28736) );
  XNOR U28142 ( .A(n28737), .B(n28738), .Z(n28734) );
  AND U28143 ( .A(n2336), .B(n28739), .Z(n28738) );
  XOR U28144 ( .A(n28740), .B(n28741), .Z(n28732) );
  AND U28145 ( .A(n2340), .B(n28731), .Z(n28741) );
  XNOR U28146 ( .A(n28742), .B(n28729), .Z(n28731) );
  XOR U28147 ( .A(n28743), .B(n28744), .Z(n28729) );
  AND U28148 ( .A(n2363), .B(n28745), .Z(n28744) );
  IV U28149 ( .A(n28740), .Z(n28742) );
  XOR U28150 ( .A(n28746), .B(n28747), .Z(n28740) );
  AND U28151 ( .A(n2347), .B(n28739), .Z(n28747) );
  XNOR U28152 ( .A(n28737), .B(n28746), .Z(n28739) );
  XNOR U28153 ( .A(n28748), .B(n28749), .Z(n28737) );
  AND U28154 ( .A(n2351), .B(n28750), .Z(n28749) );
  XOR U28155 ( .A(p_input[1920]), .B(n28748), .Z(n28750) );
  XNOR U28156 ( .A(n28751), .B(n28752), .Z(n28748) );
  AND U28157 ( .A(n2355), .B(n28753), .Z(n28752) );
  XOR U28158 ( .A(n28754), .B(n28755), .Z(n28746) );
  AND U28159 ( .A(n2359), .B(n28745), .Z(n28755) );
  XNOR U28160 ( .A(n28756), .B(n28743), .Z(n28745) );
  XOR U28161 ( .A(n28757), .B(n28758), .Z(n28743) );
  AND U28162 ( .A(n2382), .B(n28759), .Z(n28758) );
  IV U28163 ( .A(n28754), .Z(n28756) );
  XOR U28164 ( .A(n28760), .B(n28761), .Z(n28754) );
  AND U28165 ( .A(n2366), .B(n28753), .Z(n28761) );
  XNOR U28166 ( .A(n28751), .B(n28760), .Z(n28753) );
  XNOR U28167 ( .A(n28762), .B(n28763), .Z(n28751) );
  AND U28168 ( .A(n2370), .B(n28764), .Z(n28763) );
  XOR U28169 ( .A(p_input[1936]), .B(n28762), .Z(n28764) );
  XNOR U28170 ( .A(n28765), .B(n28766), .Z(n28762) );
  AND U28171 ( .A(n2374), .B(n28767), .Z(n28766) );
  XOR U28172 ( .A(n28768), .B(n28769), .Z(n28760) );
  AND U28173 ( .A(n2378), .B(n28759), .Z(n28769) );
  XNOR U28174 ( .A(n28770), .B(n28757), .Z(n28759) );
  XOR U28175 ( .A(n28771), .B(n28772), .Z(n28757) );
  AND U28176 ( .A(n2401), .B(n28773), .Z(n28772) );
  IV U28177 ( .A(n28768), .Z(n28770) );
  XOR U28178 ( .A(n28774), .B(n28775), .Z(n28768) );
  AND U28179 ( .A(n2385), .B(n28767), .Z(n28775) );
  XNOR U28180 ( .A(n28765), .B(n28774), .Z(n28767) );
  XNOR U28181 ( .A(n28776), .B(n28777), .Z(n28765) );
  AND U28182 ( .A(n2389), .B(n28778), .Z(n28777) );
  XOR U28183 ( .A(p_input[1952]), .B(n28776), .Z(n28778) );
  XNOR U28184 ( .A(n28779), .B(n28780), .Z(n28776) );
  AND U28185 ( .A(n2393), .B(n28781), .Z(n28780) );
  XOR U28186 ( .A(n28782), .B(n28783), .Z(n28774) );
  AND U28187 ( .A(n2397), .B(n28773), .Z(n28783) );
  XNOR U28188 ( .A(n28784), .B(n28771), .Z(n28773) );
  XOR U28189 ( .A(n28785), .B(n28786), .Z(n28771) );
  AND U28190 ( .A(n2420), .B(n28787), .Z(n28786) );
  IV U28191 ( .A(n28782), .Z(n28784) );
  XOR U28192 ( .A(n28788), .B(n28789), .Z(n28782) );
  AND U28193 ( .A(n2404), .B(n28781), .Z(n28789) );
  XNOR U28194 ( .A(n28779), .B(n28788), .Z(n28781) );
  XNOR U28195 ( .A(n28790), .B(n28791), .Z(n28779) );
  AND U28196 ( .A(n2408), .B(n28792), .Z(n28791) );
  XOR U28197 ( .A(p_input[1968]), .B(n28790), .Z(n28792) );
  XNOR U28198 ( .A(n28793), .B(n28794), .Z(n28790) );
  AND U28199 ( .A(n2412), .B(n28795), .Z(n28794) );
  XOR U28200 ( .A(n28796), .B(n28797), .Z(n28788) );
  AND U28201 ( .A(n2416), .B(n28787), .Z(n28797) );
  XNOR U28202 ( .A(n28798), .B(n28785), .Z(n28787) );
  XOR U28203 ( .A(n28799), .B(n28800), .Z(n28785) );
  AND U28204 ( .A(n2438), .B(n28801), .Z(n28800) );
  IV U28205 ( .A(n28796), .Z(n28798) );
  XOR U28206 ( .A(n28802), .B(n28803), .Z(n28796) );
  AND U28207 ( .A(n2423), .B(n28795), .Z(n28803) );
  XNOR U28208 ( .A(n28793), .B(n28802), .Z(n28795) );
  XNOR U28209 ( .A(n28804), .B(n28805), .Z(n28793) );
  AND U28210 ( .A(n2427), .B(n28806), .Z(n28805) );
  XOR U28211 ( .A(p_input[1984]), .B(n28804), .Z(n28806) );
  XOR U28212 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n28807), 
        .Z(n28804) );
  AND U28213 ( .A(n2430), .B(n28808), .Z(n28807) );
  XOR U28214 ( .A(n28809), .B(n28810), .Z(n28802) );
  AND U28215 ( .A(n2434), .B(n28801), .Z(n28810) );
  XNOR U28216 ( .A(n28811), .B(n28799), .Z(n28801) );
  XOR U28217 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n28812), .Z(n28799) );
  AND U28218 ( .A(n2446), .B(n28813), .Z(n28812) );
  IV U28219 ( .A(n28809), .Z(n28811) );
  XOR U28220 ( .A(n28814), .B(n28815), .Z(n28809) );
  AND U28221 ( .A(n2441), .B(n28808), .Z(n28815) );
  XOR U28222 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n28814), 
        .Z(n28808) );
  XOR U28223 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n28816), 
        .Z(n28814) );
  AND U28224 ( .A(n2443), .B(n28813), .Z(n28816) );
  XOR U28225 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n28813) );
  XNOR U28226 ( .A(n28817), .B(n28818), .Z(n62) );
  AND U28227 ( .A(n28819), .B(n28820), .Z(n28818) );
  XNOR U28228 ( .A(n28817), .B(n28821), .Z(n28820) );
  XOR U28229 ( .A(n28822), .B(n28823), .Z(n28821) );
  AND U28230 ( .A(n65), .B(n28824), .Z(n28823) );
  XNOR U28231 ( .A(n28822), .B(n28825), .Z(n28824) );
  IV U28232 ( .A(n28826), .Z(n28822) );
  XNOR U28233 ( .A(n28817), .B(n28827), .Z(n28819) );
  XOR U28234 ( .A(n28828), .B(n28829), .Z(n28827) );
  AND U28235 ( .A(n82), .B(n28830), .Z(n28829) );
  XOR U28236 ( .A(n28831), .B(n28832), .Z(n28817) );
  AND U28237 ( .A(n28833), .B(n28834), .Z(n28832) );
  XOR U28238 ( .A(n28835), .B(n28831), .Z(n28834) );
  XNOR U28239 ( .A(n28836), .B(n28837), .Z(n28835) );
  AND U28240 ( .A(n65), .B(n28838), .Z(n28837) );
  XNOR U28241 ( .A(n28839), .B(n28836), .Z(n28838) );
  XNOR U28242 ( .A(n28831), .B(n28840), .Z(n28833) );
  XOR U28243 ( .A(n28841), .B(n28842), .Z(n28840) );
  AND U28244 ( .A(n82), .B(n28843), .Z(n28842) );
  XOR U28245 ( .A(n28844), .B(n28845), .Z(n28831) );
  AND U28246 ( .A(n28846), .B(n28847), .Z(n28845) );
  XOR U28247 ( .A(n28848), .B(n28844), .Z(n28847) );
  XNOR U28248 ( .A(n28849), .B(n28850), .Z(n28848) );
  AND U28249 ( .A(n65), .B(n28851), .Z(n28850) );
  XNOR U28250 ( .A(n28852), .B(n28849), .Z(n28851) );
  XNOR U28251 ( .A(n28844), .B(n28853), .Z(n28846) );
  XOR U28252 ( .A(n28854), .B(n28855), .Z(n28853) );
  AND U28253 ( .A(n82), .B(n28856), .Z(n28855) );
  XOR U28254 ( .A(n28857), .B(n28858), .Z(n28844) );
  AND U28255 ( .A(n28859), .B(n28860), .Z(n28858) );
  XOR U28256 ( .A(n28857), .B(n28861), .Z(n28860) );
  XOR U28257 ( .A(n28862), .B(n28863), .Z(n28861) );
  AND U28258 ( .A(n65), .B(n28864), .Z(n28863) );
  XOR U28259 ( .A(n28865), .B(n28862), .Z(n28864) );
  XNOR U28260 ( .A(n28866), .B(n28857), .Z(n28859) );
  XNOR U28261 ( .A(n28867), .B(n28868), .Z(n28866) );
  AND U28262 ( .A(n82), .B(n28869), .Z(n28868) );
  AND U28263 ( .A(n28870), .B(n28871), .Z(n28857) );
  XNOR U28264 ( .A(n28872), .B(n28873), .Z(n28871) );
  AND U28265 ( .A(n65), .B(n28874), .Z(n28873) );
  XNOR U28266 ( .A(n28875), .B(n28872), .Z(n28874) );
  XNOR U28267 ( .A(n28876), .B(n28877), .Z(n65) );
  AND U28268 ( .A(n28878), .B(n28879), .Z(n28877) );
  XOR U28269 ( .A(n28825), .B(n28876), .Z(n28879) );
  XOR U28270 ( .A(n28880), .B(n28881), .Z(n28825) );
  AND U28271 ( .A(n70), .B(n28882), .Z(n28881) );
  XOR U28272 ( .A(n28883), .B(n28880), .Z(n28882) );
  XNOR U28273 ( .A(n28826), .B(n28876), .Z(n28878) );
  XOR U28274 ( .A(n28884), .B(n28885), .Z(n28826) );
  AND U28275 ( .A(n78), .B(n28830), .Z(n28885) );
  XOR U28276 ( .A(n28828), .B(n28884), .Z(n28830) );
  XOR U28277 ( .A(n28886), .B(n28887), .Z(n28876) );
  AND U28278 ( .A(n28888), .B(n28889), .Z(n28887) );
  XOR U28279 ( .A(n28839), .B(n28886), .Z(n28889) );
  XOR U28280 ( .A(n28890), .B(n28891), .Z(n28839) );
  AND U28281 ( .A(n70), .B(n28892), .Z(n28891) );
  XOR U28282 ( .A(n28893), .B(n28890), .Z(n28892) );
  XOR U28283 ( .A(n28886), .B(n28836), .Z(n28888) );
  XOR U28284 ( .A(n28894), .B(n28895), .Z(n28836) );
  AND U28285 ( .A(n78), .B(n28843), .Z(n28895) );
  XOR U28286 ( .A(n28894), .B(n28896), .Z(n28843) );
  XOR U28287 ( .A(n28897), .B(n28898), .Z(n28886) );
  AND U28288 ( .A(n28899), .B(n28900), .Z(n28898) );
  XOR U28289 ( .A(n28852), .B(n28897), .Z(n28900) );
  XOR U28290 ( .A(n28901), .B(n28902), .Z(n28852) );
  AND U28291 ( .A(n70), .B(n28903), .Z(n28902) );
  XNOR U28292 ( .A(n28904), .B(n28901), .Z(n28903) );
  XOR U28293 ( .A(n28897), .B(n28849), .Z(n28899) );
  XOR U28294 ( .A(n28905), .B(n28906), .Z(n28849) );
  AND U28295 ( .A(n78), .B(n28856), .Z(n28906) );
  XOR U28296 ( .A(n28905), .B(n28907), .Z(n28856) );
  XOR U28297 ( .A(n28908), .B(n28909), .Z(n28897) );
  AND U28298 ( .A(n28910), .B(n28911), .Z(n28909) );
  XOR U28299 ( .A(n28908), .B(n28865), .Z(n28911) );
  XOR U28300 ( .A(n28912), .B(n28913), .Z(n28865) );
  AND U28301 ( .A(n70), .B(n28914), .Z(n28913) );
  XOR U28302 ( .A(n28915), .B(n28912), .Z(n28914) );
  XNOR U28303 ( .A(n28862), .B(n28908), .Z(n28910) );
  XNOR U28304 ( .A(n28916), .B(n28917), .Z(n28862) );
  AND U28305 ( .A(n78), .B(n28869), .Z(n28917) );
  XOR U28306 ( .A(n28916), .B(n28867), .Z(n28869) );
  AND U28307 ( .A(n28872), .B(n28875), .Z(n28908) );
  XOR U28308 ( .A(n28918), .B(n28919), .Z(n28875) );
  AND U28309 ( .A(n70), .B(n28920), .Z(n28919) );
  XNOR U28310 ( .A(n28921), .B(n28922), .Z(n28920) );
  XNOR U28311 ( .A(n28923), .B(n28924), .Z(n70) );
  AND U28312 ( .A(n28925), .B(n28926), .Z(n28924) );
  XOR U28313 ( .A(n28883), .B(n28923), .Z(n28926) );
  AND U28314 ( .A(n28927), .B(n28928), .Z(n28883) );
  XNOR U28315 ( .A(n28880), .B(n28923), .Z(n28925) );
  XNOR U28316 ( .A(n28929), .B(n28930), .Z(n28880) );
  AND U28317 ( .A(n74), .B(n28931), .Z(n28930) );
  XNOR U28318 ( .A(n28932), .B(n28933), .Z(n28931) );
  XOR U28319 ( .A(n28934), .B(n28935), .Z(n28923) );
  AND U28320 ( .A(n28936), .B(n28937), .Z(n28935) );
  XNOR U28321 ( .A(n28934), .B(n28927), .Z(n28937) );
  IV U28322 ( .A(n28893), .Z(n28927) );
  XOR U28323 ( .A(n28938), .B(n28939), .Z(n28893) );
  XOR U28324 ( .A(n28940), .B(n28928), .Z(n28939) );
  AND U28325 ( .A(n28904), .B(n28941), .Z(n28928) );
  AND U28326 ( .A(n28942), .B(n28943), .Z(n28940) );
  XOR U28327 ( .A(n28944), .B(n28938), .Z(n28942) );
  XNOR U28328 ( .A(n28890), .B(n28934), .Z(n28936) );
  XNOR U28329 ( .A(n28945), .B(n28946), .Z(n28890) );
  AND U28330 ( .A(n74), .B(n28947), .Z(n28946) );
  XNOR U28331 ( .A(n28948), .B(n28949), .Z(n28947) );
  XOR U28332 ( .A(n28950), .B(n28951), .Z(n28934) );
  AND U28333 ( .A(n28952), .B(n28953), .Z(n28951) );
  XNOR U28334 ( .A(n28950), .B(n28904), .Z(n28953) );
  XOR U28335 ( .A(n28954), .B(n28943), .Z(n28904) );
  XNOR U28336 ( .A(n28955), .B(n28938), .Z(n28943) );
  XOR U28337 ( .A(n28956), .B(n28957), .Z(n28938) );
  AND U28338 ( .A(n28958), .B(n28959), .Z(n28957) );
  XOR U28339 ( .A(n28960), .B(n28956), .Z(n28958) );
  XNOR U28340 ( .A(n28961), .B(n28962), .Z(n28955) );
  AND U28341 ( .A(n28963), .B(n28964), .Z(n28962) );
  XOR U28342 ( .A(n28961), .B(n28965), .Z(n28963) );
  XNOR U28343 ( .A(n28944), .B(n28941), .Z(n28954) );
  AND U28344 ( .A(n28966), .B(n28967), .Z(n28941) );
  XOR U28345 ( .A(n28968), .B(n28969), .Z(n28944) );
  AND U28346 ( .A(n28970), .B(n28971), .Z(n28969) );
  XOR U28347 ( .A(n28968), .B(n28972), .Z(n28970) );
  XNOR U28348 ( .A(n28901), .B(n28950), .Z(n28952) );
  XNOR U28349 ( .A(n28973), .B(n28974), .Z(n28901) );
  AND U28350 ( .A(n74), .B(n28975), .Z(n28974) );
  XNOR U28351 ( .A(n28976), .B(n28977), .Z(n28975) );
  XOR U28352 ( .A(n28978), .B(n28979), .Z(n28950) );
  AND U28353 ( .A(n28980), .B(n28981), .Z(n28979) );
  XNOR U28354 ( .A(n28978), .B(n28966), .Z(n28981) );
  IV U28355 ( .A(n28915), .Z(n28966) );
  XNOR U28356 ( .A(n28982), .B(n28959), .Z(n28915) );
  XNOR U28357 ( .A(n28983), .B(n28965), .Z(n28959) );
  XNOR U28358 ( .A(n28984), .B(n28985), .Z(n28965) );
  NOR U28359 ( .A(n28986), .B(n28987), .Z(n28985) );
  XOR U28360 ( .A(n28984), .B(n28988), .Z(n28986) );
  XNOR U28361 ( .A(n28964), .B(n28956), .Z(n28983) );
  XOR U28362 ( .A(n28989), .B(n28990), .Z(n28956) );
  AND U28363 ( .A(n28991), .B(n28992), .Z(n28990) );
  XNOR U28364 ( .A(n28989), .B(n28993), .Z(n28991) );
  XNOR U28365 ( .A(n28994), .B(n28961), .Z(n28964) );
  XOR U28366 ( .A(n28995), .B(n28996), .Z(n28961) );
  AND U28367 ( .A(n28997), .B(n28998), .Z(n28996) );
  XOR U28368 ( .A(n28995), .B(n28999), .Z(n28997) );
  XNOR U28369 ( .A(n29000), .B(n29001), .Z(n28994) );
  NOR U28370 ( .A(n29002), .B(n29003), .Z(n29001) );
  XNOR U28371 ( .A(n29000), .B(n29004), .Z(n29002) );
  XNOR U28372 ( .A(n28960), .B(n28967), .Z(n28982) );
  NOR U28373 ( .A(n28921), .B(n29005), .Z(n28967) );
  XOR U28374 ( .A(n28972), .B(n28971), .Z(n28960) );
  XNOR U28375 ( .A(n29006), .B(n28968), .Z(n28971) );
  XOR U28376 ( .A(n29007), .B(n29008), .Z(n28968) );
  AND U28377 ( .A(n29009), .B(n29010), .Z(n29008) );
  XOR U28378 ( .A(n29007), .B(n29011), .Z(n29009) );
  XNOR U28379 ( .A(n29012), .B(n29013), .Z(n29006) );
  NOR U28380 ( .A(n29014), .B(n29015), .Z(n29013) );
  XNOR U28381 ( .A(n29012), .B(n29016), .Z(n29014) );
  XOR U28382 ( .A(n29017), .B(n29018), .Z(n28972) );
  NOR U28383 ( .A(n29019), .B(n29020), .Z(n29018) );
  XNOR U28384 ( .A(n29017), .B(n29021), .Z(n29019) );
  XNOR U28385 ( .A(n28912), .B(n28978), .Z(n28980) );
  XNOR U28386 ( .A(n29022), .B(n29023), .Z(n28912) );
  AND U28387 ( .A(n74), .B(n29024), .Z(n29023) );
  XNOR U28388 ( .A(n29025), .B(n29026), .Z(n29024) );
  AND U28389 ( .A(n28922), .B(n28921), .Z(n28978) );
  XOR U28390 ( .A(n29027), .B(n29005), .Z(n28921) );
  XNOR U28391 ( .A(p_input[0]), .B(p_input[2048]), .Z(n29005) );
  XOR U28392 ( .A(n28993), .B(n28992), .Z(n29027) );
  XNOR U28393 ( .A(n29028), .B(n28999), .Z(n28992) );
  XNOR U28394 ( .A(n28988), .B(n28987), .Z(n28999) );
  XNOR U28395 ( .A(n29029), .B(n28984), .Z(n28987) );
  XNOR U28396 ( .A(p_input[10]), .B(p_input[2058]), .Z(n28984) );
  XOR U28397 ( .A(p_input[11]), .B(n29030), .Z(n29029) );
  XOR U28398 ( .A(p_input[12]), .B(p_input[2060]), .Z(n28988) );
  XOR U28399 ( .A(n28998), .B(n29031), .Z(n29028) );
  IV U28400 ( .A(n28989), .Z(n29031) );
  XOR U28401 ( .A(p_input[1]), .B(p_input[2049]), .Z(n28989) );
  XNOR U28402 ( .A(n29032), .B(n29004), .Z(n28998) );
  XNOR U28403 ( .A(p_input[15]), .B(n29033), .Z(n29004) );
  XOR U28404 ( .A(n28995), .B(n29003), .Z(n29032) );
  XOR U28405 ( .A(n29034), .B(n29000), .Z(n29003) );
  XOR U28406 ( .A(p_input[13]), .B(p_input[2061]), .Z(n29000) );
  XOR U28407 ( .A(p_input[14]), .B(n29035), .Z(n29034) );
  XNOR U28408 ( .A(n29036), .B(p_input[9]), .Z(n28995) );
  XNOR U28409 ( .A(n29011), .B(n29010), .Z(n28993) );
  XNOR U28410 ( .A(n29037), .B(n29016), .Z(n29010) );
  XOR U28411 ( .A(p_input[2056]), .B(p_input[8]), .Z(n29016) );
  XOR U28412 ( .A(n29007), .B(n29015), .Z(n29037) );
  XOR U28413 ( .A(n29038), .B(n29012), .Z(n29015) );
  XOR U28414 ( .A(p_input[2054]), .B(p_input[6]), .Z(n29012) );
  XNOR U28415 ( .A(p_input[2055]), .B(p_input[7]), .Z(n29038) );
  XNOR U28416 ( .A(n29039), .B(p_input[2]), .Z(n29007) );
  XNOR U28417 ( .A(n29021), .B(n29020), .Z(n29011) );
  XOR U28418 ( .A(n29040), .B(n29017), .Z(n29020) );
  XOR U28419 ( .A(p_input[2051]), .B(p_input[3]), .Z(n29017) );
  XNOR U28420 ( .A(p_input[2052]), .B(p_input[4]), .Z(n29040) );
  XOR U28421 ( .A(p_input[2053]), .B(p_input[5]), .Z(n29021) );
  IV U28422 ( .A(n28918), .Z(n28922) );
  XOR U28423 ( .A(n29041), .B(n29042), .Z(n28918) );
  AND U28424 ( .A(n74), .B(n29043), .Z(n29042) );
  XNOR U28425 ( .A(n29044), .B(n29045), .Z(n74) );
  AND U28426 ( .A(n29046), .B(n29047), .Z(n29045) );
  XOR U28427 ( .A(n28933), .B(n29044), .Z(n29047) );
  XNOR U28428 ( .A(n29048), .B(n29044), .Z(n29046) );
  XOR U28429 ( .A(n29049), .B(n29050), .Z(n29044) );
  AND U28430 ( .A(n29051), .B(n29052), .Z(n29050) );
  XOR U28431 ( .A(n28948), .B(n29049), .Z(n29052) );
  XOR U28432 ( .A(n29049), .B(n28949), .Z(n29051) );
  XOR U28433 ( .A(n29053), .B(n29054), .Z(n29049) );
  AND U28434 ( .A(n29055), .B(n29056), .Z(n29054) );
  XOR U28435 ( .A(n28976), .B(n29053), .Z(n29056) );
  XOR U28436 ( .A(n29053), .B(n28977), .Z(n29055) );
  XOR U28437 ( .A(n29057), .B(n29058), .Z(n29053) );
  AND U28438 ( .A(n29059), .B(n29060), .Z(n29058) );
  XOR U28439 ( .A(n29057), .B(n29025), .Z(n29060) );
  XNOR U28440 ( .A(n29061), .B(n29062), .Z(n28872) );
  AND U28441 ( .A(n78), .B(n29063), .Z(n29062) );
  XNOR U28442 ( .A(n29064), .B(n29065), .Z(n78) );
  AND U28443 ( .A(n29066), .B(n29067), .Z(n29065) );
  XOR U28444 ( .A(n29064), .B(n28884), .Z(n29067) );
  XNOR U28445 ( .A(n29064), .B(n28828), .Z(n29066) );
  XOR U28446 ( .A(n29068), .B(n29069), .Z(n29064) );
  AND U28447 ( .A(n29070), .B(n29071), .Z(n29069) );
  XNOR U28448 ( .A(n28894), .B(n29068), .Z(n29071) );
  XOR U28449 ( .A(n29068), .B(n28896), .Z(n29070) );
  XOR U28450 ( .A(n29072), .B(n29073), .Z(n29068) );
  AND U28451 ( .A(n29074), .B(n29075), .Z(n29073) );
  XOR U28452 ( .A(n29072), .B(n28907), .Z(n29074) );
  IV U28453 ( .A(n28854), .Z(n28907) );
  XOR U28454 ( .A(n29076), .B(n29077), .Z(n28870) );
  AND U28455 ( .A(n82), .B(n29063), .Z(n29077) );
  XNOR U28456 ( .A(n29061), .B(n29076), .Z(n29063) );
  XNOR U28457 ( .A(n29078), .B(n29079), .Z(n82) );
  AND U28458 ( .A(n29080), .B(n29081), .Z(n29079) );
  XNOR U28459 ( .A(n29082), .B(n29078), .Z(n29081) );
  IV U28460 ( .A(n28884), .Z(n29082) );
  XOR U28461 ( .A(n29048), .B(n29083), .Z(n28884) );
  AND U28462 ( .A(n86), .B(n29084), .Z(n29083) );
  XOR U28463 ( .A(n28932), .B(n28929), .Z(n29084) );
  IV U28464 ( .A(n29048), .Z(n28932) );
  XNOR U28465 ( .A(n28828), .B(n29078), .Z(n29080) );
  XOR U28466 ( .A(n29085), .B(n29086), .Z(n28828) );
  AND U28467 ( .A(n102), .B(n29087), .Z(n29086) );
  XOR U28468 ( .A(n29088), .B(n29089), .Z(n29078) );
  AND U28469 ( .A(n29090), .B(n29091), .Z(n29089) );
  XNOR U28470 ( .A(n29088), .B(n28894), .Z(n29091) );
  XOR U28471 ( .A(n28949), .B(n29092), .Z(n28894) );
  AND U28472 ( .A(n86), .B(n29093), .Z(n29092) );
  XOR U28473 ( .A(n28945), .B(n28949), .Z(n29093) );
  XNOR U28474 ( .A(n28841), .B(n29088), .Z(n29090) );
  IV U28475 ( .A(n28896), .Z(n28841) );
  XOR U28476 ( .A(n29094), .B(n29095), .Z(n28896) );
  AND U28477 ( .A(n102), .B(n29096), .Z(n29095) );
  XOR U28478 ( .A(n29072), .B(n29097), .Z(n29088) );
  AND U28479 ( .A(n29098), .B(n29075), .Z(n29097) );
  XNOR U28480 ( .A(n28905), .B(n29072), .Z(n29075) );
  XOR U28481 ( .A(n28977), .B(n29099), .Z(n28905) );
  AND U28482 ( .A(n86), .B(n29100), .Z(n29099) );
  XOR U28483 ( .A(n28973), .B(n28977), .Z(n29100) );
  XNOR U28484 ( .A(n28854), .B(n29072), .Z(n29098) );
  XNOR U28485 ( .A(n29101), .B(n29102), .Z(n28854) );
  AND U28486 ( .A(n102), .B(n29103), .Z(n29102) );
  XOR U28487 ( .A(n29104), .B(n29105), .Z(n29072) );
  AND U28488 ( .A(n29106), .B(n29107), .Z(n29105) );
  XNOR U28489 ( .A(n29104), .B(n28916), .Z(n29107) );
  XOR U28490 ( .A(n29026), .B(n29108), .Z(n28916) );
  AND U28491 ( .A(n86), .B(n29109), .Z(n29108) );
  XOR U28492 ( .A(n29022), .B(n29026), .Z(n29109) );
  XNOR U28493 ( .A(n29110), .B(n29104), .Z(n29106) );
  IV U28494 ( .A(n28867), .Z(n29110) );
  XOR U28495 ( .A(n29111), .B(n29112), .Z(n28867) );
  AND U28496 ( .A(n102), .B(n29113), .Z(n29112) );
  AND U28497 ( .A(n29076), .B(n29061), .Z(n29104) );
  XNOR U28498 ( .A(n29114), .B(n29115), .Z(n29061) );
  AND U28499 ( .A(n86), .B(n29043), .Z(n29115) );
  XNOR U28500 ( .A(n29041), .B(n29114), .Z(n29043) );
  XNOR U28501 ( .A(n29116), .B(n29117), .Z(n86) );
  AND U28502 ( .A(n29118), .B(n29119), .Z(n29117) );
  XNOR U28503 ( .A(n29116), .B(n28929), .Z(n29119) );
  IV U28504 ( .A(n28933), .Z(n28929) );
  XOR U28505 ( .A(n29120), .B(n29121), .Z(n28933) );
  AND U28506 ( .A(n90), .B(n29122), .Z(n29121) );
  XOR U28507 ( .A(n29123), .B(n29120), .Z(n29122) );
  XNOR U28508 ( .A(n29116), .B(n29048), .Z(n29118) );
  XOR U28509 ( .A(n29124), .B(n29125), .Z(n29048) );
  AND U28510 ( .A(n98), .B(n29087), .Z(n29125) );
  XOR U28511 ( .A(n29085), .B(n29124), .Z(n29087) );
  XOR U28512 ( .A(n29126), .B(n29127), .Z(n29116) );
  AND U28513 ( .A(n29128), .B(n29129), .Z(n29127) );
  XNOR U28514 ( .A(n29126), .B(n28945), .Z(n29129) );
  IV U28515 ( .A(n28948), .Z(n28945) );
  XOR U28516 ( .A(n29130), .B(n29131), .Z(n28948) );
  AND U28517 ( .A(n90), .B(n29132), .Z(n29131) );
  XOR U28518 ( .A(n29133), .B(n29130), .Z(n29132) );
  XOR U28519 ( .A(n28949), .B(n29126), .Z(n29128) );
  XOR U28520 ( .A(n29134), .B(n29135), .Z(n28949) );
  AND U28521 ( .A(n98), .B(n29096), .Z(n29135) );
  XOR U28522 ( .A(n29134), .B(n29094), .Z(n29096) );
  XOR U28523 ( .A(n29136), .B(n29137), .Z(n29126) );
  AND U28524 ( .A(n29138), .B(n29139), .Z(n29137) );
  XNOR U28525 ( .A(n29136), .B(n28973), .Z(n29139) );
  IV U28526 ( .A(n28976), .Z(n28973) );
  XOR U28527 ( .A(n29140), .B(n29141), .Z(n28976) );
  AND U28528 ( .A(n90), .B(n29142), .Z(n29141) );
  XNOR U28529 ( .A(n29143), .B(n29140), .Z(n29142) );
  XOR U28530 ( .A(n28977), .B(n29136), .Z(n29138) );
  XOR U28531 ( .A(n29144), .B(n29145), .Z(n28977) );
  AND U28532 ( .A(n98), .B(n29103), .Z(n29145) );
  XOR U28533 ( .A(n29144), .B(n29101), .Z(n29103) );
  XOR U28534 ( .A(n29057), .B(n29146), .Z(n29136) );
  AND U28535 ( .A(n29059), .B(n29147), .Z(n29146) );
  XNOR U28536 ( .A(n29057), .B(n29022), .Z(n29147) );
  IV U28537 ( .A(n29025), .Z(n29022) );
  XOR U28538 ( .A(n29148), .B(n29149), .Z(n29025) );
  AND U28539 ( .A(n90), .B(n29150), .Z(n29149) );
  XOR U28540 ( .A(n29151), .B(n29148), .Z(n29150) );
  XOR U28541 ( .A(n29026), .B(n29057), .Z(n29059) );
  XOR U28542 ( .A(n29152), .B(n29153), .Z(n29026) );
  AND U28543 ( .A(n98), .B(n29113), .Z(n29153) );
  XOR U28544 ( .A(n29152), .B(n29111), .Z(n29113) );
  AND U28545 ( .A(n29114), .B(n29041), .Z(n29057) );
  XNOR U28546 ( .A(n29154), .B(n29155), .Z(n29041) );
  AND U28547 ( .A(n90), .B(n29156), .Z(n29155) );
  XNOR U28548 ( .A(n29157), .B(n29154), .Z(n29156) );
  XNOR U28549 ( .A(n29158), .B(n29159), .Z(n90) );
  AND U28550 ( .A(n29160), .B(n29161), .Z(n29159) );
  XOR U28551 ( .A(n29123), .B(n29158), .Z(n29161) );
  AND U28552 ( .A(n29162), .B(n29163), .Z(n29123) );
  XNOR U28553 ( .A(n29120), .B(n29158), .Z(n29160) );
  XNOR U28554 ( .A(n29164), .B(n29165), .Z(n29120) );
  AND U28555 ( .A(n94), .B(n29166), .Z(n29165) );
  XNOR U28556 ( .A(n29167), .B(n29168), .Z(n29166) );
  XOR U28557 ( .A(n29169), .B(n29170), .Z(n29158) );
  AND U28558 ( .A(n29171), .B(n29172), .Z(n29170) );
  XNOR U28559 ( .A(n29169), .B(n29162), .Z(n29172) );
  IV U28560 ( .A(n29133), .Z(n29162) );
  XOR U28561 ( .A(n29173), .B(n29174), .Z(n29133) );
  XOR U28562 ( .A(n29175), .B(n29163), .Z(n29174) );
  AND U28563 ( .A(n29143), .B(n29176), .Z(n29163) );
  AND U28564 ( .A(n29177), .B(n29178), .Z(n29175) );
  XOR U28565 ( .A(n29179), .B(n29173), .Z(n29177) );
  XNOR U28566 ( .A(n29130), .B(n29169), .Z(n29171) );
  XNOR U28567 ( .A(n29180), .B(n29181), .Z(n29130) );
  AND U28568 ( .A(n94), .B(n29182), .Z(n29181) );
  XNOR U28569 ( .A(n29183), .B(n29184), .Z(n29182) );
  XOR U28570 ( .A(n29185), .B(n29186), .Z(n29169) );
  AND U28571 ( .A(n29187), .B(n29188), .Z(n29186) );
  XNOR U28572 ( .A(n29185), .B(n29143), .Z(n29188) );
  XOR U28573 ( .A(n29189), .B(n29178), .Z(n29143) );
  XNOR U28574 ( .A(n29190), .B(n29173), .Z(n29178) );
  XOR U28575 ( .A(n29191), .B(n29192), .Z(n29173) );
  AND U28576 ( .A(n29193), .B(n29194), .Z(n29192) );
  XOR U28577 ( .A(n29195), .B(n29191), .Z(n29193) );
  XNOR U28578 ( .A(n29196), .B(n29197), .Z(n29190) );
  AND U28579 ( .A(n29198), .B(n29199), .Z(n29197) );
  XOR U28580 ( .A(n29196), .B(n29200), .Z(n29198) );
  XNOR U28581 ( .A(n29179), .B(n29176), .Z(n29189) );
  AND U28582 ( .A(n29201), .B(n29202), .Z(n29176) );
  XOR U28583 ( .A(n29203), .B(n29204), .Z(n29179) );
  AND U28584 ( .A(n29205), .B(n29206), .Z(n29204) );
  XOR U28585 ( .A(n29203), .B(n29207), .Z(n29205) );
  XNOR U28586 ( .A(n29140), .B(n29185), .Z(n29187) );
  XNOR U28587 ( .A(n29208), .B(n29209), .Z(n29140) );
  AND U28588 ( .A(n94), .B(n29210), .Z(n29209) );
  XNOR U28589 ( .A(n29211), .B(n29212), .Z(n29210) );
  XOR U28590 ( .A(n29213), .B(n29214), .Z(n29185) );
  AND U28591 ( .A(n29215), .B(n29216), .Z(n29214) );
  XNOR U28592 ( .A(n29213), .B(n29201), .Z(n29216) );
  IV U28593 ( .A(n29151), .Z(n29201) );
  XNOR U28594 ( .A(n29217), .B(n29194), .Z(n29151) );
  XNOR U28595 ( .A(n29218), .B(n29200), .Z(n29194) );
  XOR U28596 ( .A(n29219), .B(n29220), .Z(n29200) );
  NOR U28597 ( .A(n29221), .B(n29222), .Z(n29220) );
  XNOR U28598 ( .A(n29219), .B(n29223), .Z(n29221) );
  XNOR U28599 ( .A(n29199), .B(n29191), .Z(n29218) );
  XOR U28600 ( .A(n29224), .B(n29225), .Z(n29191) );
  AND U28601 ( .A(n29226), .B(n29227), .Z(n29225) );
  XNOR U28602 ( .A(n29224), .B(n29228), .Z(n29226) );
  XNOR U28603 ( .A(n29229), .B(n29196), .Z(n29199) );
  XOR U28604 ( .A(n29230), .B(n29231), .Z(n29196) );
  AND U28605 ( .A(n29232), .B(n29233), .Z(n29231) );
  XOR U28606 ( .A(n29230), .B(n29234), .Z(n29232) );
  XNOR U28607 ( .A(n29235), .B(n29236), .Z(n29229) );
  NOR U28608 ( .A(n29237), .B(n29238), .Z(n29236) );
  XOR U28609 ( .A(n29235), .B(n29239), .Z(n29237) );
  XNOR U28610 ( .A(n29195), .B(n29202), .Z(n29217) );
  NOR U28611 ( .A(n29157), .B(n29240), .Z(n29202) );
  XOR U28612 ( .A(n29207), .B(n29206), .Z(n29195) );
  XNOR U28613 ( .A(n29241), .B(n29203), .Z(n29206) );
  XOR U28614 ( .A(n29242), .B(n29243), .Z(n29203) );
  AND U28615 ( .A(n29244), .B(n29245), .Z(n29243) );
  XNOR U28616 ( .A(n29246), .B(n29247), .Z(n29244) );
  IV U28617 ( .A(n29242), .Z(n29246) );
  XNOR U28618 ( .A(n29248), .B(n29249), .Z(n29241) );
  NOR U28619 ( .A(n29250), .B(n29251), .Z(n29249) );
  XNOR U28620 ( .A(n29248), .B(n29252), .Z(n29250) );
  XOR U28621 ( .A(n29253), .B(n29254), .Z(n29207) );
  NOR U28622 ( .A(n29255), .B(n29256), .Z(n29254) );
  XNOR U28623 ( .A(n29253), .B(n29257), .Z(n29255) );
  XNOR U28624 ( .A(n29148), .B(n29213), .Z(n29215) );
  XNOR U28625 ( .A(n29258), .B(n29259), .Z(n29148) );
  AND U28626 ( .A(n94), .B(n29260), .Z(n29259) );
  XNOR U28627 ( .A(n29261), .B(n29262), .Z(n29260) );
  AND U28628 ( .A(n29154), .B(n29157), .Z(n29213) );
  XOR U28629 ( .A(n29263), .B(n29240), .Z(n29157) );
  XNOR U28630 ( .A(p_input[16]), .B(p_input[2048]), .Z(n29240) );
  XOR U28631 ( .A(n29228), .B(n29227), .Z(n29263) );
  XNOR U28632 ( .A(n29264), .B(n29234), .Z(n29227) );
  XNOR U28633 ( .A(n29223), .B(n29222), .Z(n29234) );
  XOR U28634 ( .A(n29265), .B(n29219), .Z(n29222) );
  XNOR U28635 ( .A(n29266), .B(p_input[26]), .Z(n29219) );
  XNOR U28636 ( .A(p_input[2059]), .B(p_input[27]), .Z(n29265) );
  XOR U28637 ( .A(p_input[2060]), .B(p_input[28]), .Z(n29223) );
  XOR U28638 ( .A(n29233), .B(n29267), .Z(n29264) );
  IV U28639 ( .A(n29224), .Z(n29267) );
  XOR U28640 ( .A(p_input[17]), .B(p_input[2049]), .Z(n29224) );
  XOR U28641 ( .A(n29268), .B(n29239), .Z(n29233) );
  XNOR U28642 ( .A(p_input[2063]), .B(p_input[31]), .Z(n29239) );
  XOR U28643 ( .A(n29230), .B(n29238), .Z(n29268) );
  XOR U28644 ( .A(n29269), .B(n29235), .Z(n29238) );
  XOR U28645 ( .A(p_input[2061]), .B(p_input[29]), .Z(n29235) );
  XNOR U28646 ( .A(p_input[2062]), .B(p_input[30]), .Z(n29269) );
  XNOR U28647 ( .A(n29036), .B(p_input[25]), .Z(n29230) );
  XNOR U28648 ( .A(n29247), .B(n29245), .Z(n29228) );
  XNOR U28649 ( .A(n29270), .B(n29252), .Z(n29245) );
  XOR U28650 ( .A(p_input[2056]), .B(p_input[24]), .Z(n29252) );
  XOR U28651 ( .A(n29242), .B(n29251), .Z(n29270) );
  XOR U28652 ( .A(n29271), .B(n29248), .Z(n29251) );
  XOR U28653 ( .A(p_input[2054]), .B(p_input[22]), .Z(n29248) );
  XNOR U28654 ( .A(p_input[2055]), .B(p_input[23]), .Z(n29271) );
  XOR U28655 ( .A(p_input[18]), .B(p_input[2050]), .Z(n29242) );
  XNOR U28656 ( .A(n29257), .B(n29256), .Z(n29247) );
  XOR U28657 ( .A(n29272), .B(n29253), .Z(n29256) );
  XOR U28658 ( .A(p_input[19]), .B(p_input[2051]), .Z(n29253) );
  XNOR U28659 ( .A(p_input[2052]), .B(p_input[20]), .Z(n29272) );
  XOR U28660 ( .A(p_input[2053]), .B(p_input[21]), .Z(n29257) );
  XNOR U28661 ( .A(n29273), .B(n29274), .Z(n29154) );
  AND U28662 ( .A(n94), .B(n29275), .Z(n29274) );
  XNOR U28663 ( .A(n29276), .B(n29277), .Z(n94) );
  AND U28664 ( .A(n29278), .B(n29279), .Z(n29277) );
  XOR U28665 ( .A(n29168), .B(n29276), .Z(n29279) );
  XNOR U28666 ( .A(n29280), .B(n29276), .Z(n29278) );
  XOR U28667 ( .A(n29281), .B(n29282), .Z(n29276) );
  AND U28668 ( .A(n29283), .B(n29284), .Z(n29282) );
  XOR U28669 ( .A(n29183), .B(n29281), .Z(n29284) );
  XOR U28670 ( .A(n29281), .B(n29184), .Z(n29283) );
  XOR U28671 ( .A(n29285), .B(n29286), .Z(n29281) );
  AND U28672 ( .A(n29287), .B(n29288), .Z(n29286) );
  XOR U28673 ( .A(n29211), .B(n29285), .Z(n29288) );
  XOR U28674 ( .A(n29285), .B(n29212), .Z(n29287) );
  XOR U28675 ( .A(n29289), .B(n29290), .Z(n29285) );
  AND U28676 ( .A(n29291), .B(n29292), .Z(n29290) );
  XOR U28677 ( .A(n29289), .B(n29261), .Z(n29292) );
  XNOR U28678 ( .A(n29293), .B(n29294), .Z(n29114) );
  AND U28679 ( .A(n98), .B(n29295), .Z(n29294) );
  XNOR U28680 ( .A(n29296), .B(n29297), .Z(n98) );
  AND U28681 ( .A(n29298), .B(n29299), .Z(n29297) );
  XOR U28682 ( .A(n29296), .B(n29124), .Z(n29299) );
  XNOR U28683 ( .A(n29296), .B(n29085), .Z(n29298) );
  XOR U28684 ( .A(n29300), .B(n29301), .Z(n29296) );
  AND U28685 ( .A(n29302), .B(n29303), .Z(n29301) );
  XOR U28686 ( .A(n29300), .B(n29094), .Z(n29302) );
  XOR U28687 ( .A(n29304), .B(n29305), .Z(n29076) );
  AND U28688 ( .A(n102), .B(n29295), .Z(n29305) );
  XNOR U28689 ( .A(n29293), .B(n29304), .Z(n29295) );
  XNOR U28690 ( .A(n29306), .B(n29307), .Z(n102) );
  AND U28691 ( .A(n29308), .B(n29309), .Z(n29307) );
  XNOR U28692 ( .A(n29310), .B(n29306), .Z(n29309) );
  IV U28693 ( .A(n29124), .Z(n29310) );
  XOR U28694 ( .A(n29280), .B(n29311), .Z(n29124) );
  AND U28695 ( .A(n105), .B(n29312), .Z(n29311) );
  XOR U28696 ( .A(n29167), .B(n29164), .Z(n29312) );
  IV U28697 ( .A(n29280), .Z(n29167) );
  XNOR U28698 ( .A(n29085), .B(n29306), .Z(n29308) );
  XOR U28699 ( .A(n29313), .B(n29314), .Z(n29085) );
  AND U28700 ( .A(n121), .B(n29315), .Z(n29314) );
  XOR U28701 ( .A(n29300), .B(n29316), .Z(n29306) );
  AND U28702 ( .A(n29317), .B(n29303), .Z(n29316) );
  XNOR U28703 ( .A(n29134), .B(n29300), .Z(n29303) );
  XOR U28704 ( .A(n29184), .B(n29318), .Z(n29134) );
  AND U28705 ( .A(n105), .B(n29319), .Z(n29318) );
  XOR U28706 ( .A(n29180), .B(n29184), .Z(n29319) );
  XNOR U28707 ( .A(n29320), .B(n29300), .Z(n29317) );
  IV U28708 ( .A(n29094), .Z(n29320) );
  XOR U28709 ( .A(n29321), .B(n29322), .Z(n29094) );
  AND U28710 ( .A(n121), .B(n29323), .Z(n29322) );
  XOR U28711 ( .A(n29324), .B(n29325), .Z(n29300) );
  AND U28712 ( .A(n29326), .B(n29327), .Z(n29325) );
  XNOR U28713 ( .A(n29144), .B(n29324), .Z(n29327) );
  XOR U28714 ( .A(n29212), .B(n29328), .Z(n29144) );
  AND U28715 ( .A(n105), .B(n29329), .Z(n29328) );
  XOR U28716 ( .A(n29208), .B(n29212), .Z(n29329) );
  XOR U28717 ( .A(n29324), .B(n29101), .Z(n29326) );
  XOR U28718 ( .A(n29330), .B(n29331), .Z(n29101) );
  AND U28719 ( .A(n121), .B(n29332), .Z(n29331) );
  XOR U28720 ( .A(n29333), .B(n29334), .Z(n29324) );
  AND U28721 ( .A(n29335), .B(n29336), .Z(n29334) );
  XNOR U28722 ( .A(n29333), .B(n29152), .Z(n29336) );
  XOR U28723 ( .A(n29262), .B(n29337), .Z(n29152) );
  AND U28724 ( .A(n105), .B(n29338), .Z(n29337) );
  XOR U28725 ( .A(n29258), .B(n29262), .Z(n29338) );
  XNOR U28726 ( .A(n29339), .B(n29333), .Z(n29335) );
  IV U28727 ( .A(n29111), .Z(n29339) );
  XOR U28728 ( .A(n29340), .B(n29341), .Z(n29111) );
  AND U28729 ( .A(n121), .B(n29342), .Z(n29341) );
  AND U28730 ( .A(n29304), .B(n29293), .Z(n29333) );
  XNOR U28731 ( .A(n29343), .B(n29344), .Z(n29293) );
  AND U28732 ( .A(n105), .B(n29275), .Z(n29344) );
  XNOR U28733 ( .A(n29273), .B(n29343), .Z(n29275) );
  XNOR U28734 ( .A(n29345), .B(n29346), .Z(n105) );
  AND U28735 ( .A(n29347), .B(n29348), .Z(n29346) );
  XNOR U28736 ( .A(n29345), .B(n29164), .Z(n29348) );
  IV U28737 ( .A(n29168), .Z(n29164) );
  XOR U28738 ( .A(n29349), .B(n29350), .Z(n29168) );
  AND U28739 ( .A(n109), .B(n29351), .Z(n29350) );
  XOR U28740 ( .A(n29352), .B(n29349), .Z(n29351) );
  XNOR U28741 ( .A(n29345), .B(n29280), .Z(n29347) );
  XOR U28742 ( .A(n29353), .B(n29354), .Z(n29280) );
  AND U28743 ( .A(n117), .B(n29315), .Z(n29354) );
  XOR U28744 ( .A(n29313), .B(n29353), .Z(n29315) );
  XOR U28745 ( .A(n29355), .B(n29356), .Z(n29345) );
  AND U28746 ( .A(n29357), .B(n29358), .Z(n29356) );
  XNOR U28747 ( .A(n29355), .B(n29180), .Z(n29358) );
  IV U28748 ( .A(n29183), .Z(n29180) );
  XOR U28749 ( .A(n29359), .B(n29360), .Z(n29183) );
  AND U28750 ( .A(n109), .B(n29361), .Z(n29360) );
  XOR U28751 ( .A(n29362), .B(n29359), .Z(n29361) );
  XOR U28752 ( .A(n29184), .B(n29355), .Z(n29357) );
  XOR U28753 ( .A(n29363), .B(n29364), .Z(n29184) );
  AND U28754 ( .A(n117), .B(n29323), .Z(n29364) );
  XOR U28755 ( .A(n29363), .B(n29321), .Z(n29323) );
  XOR U28756 ( .A(n29365), .B(n29366), .Z(n29355) );
  AND U28757 ( .A(n29367), .B(n29368), .Z(n29366) );
  XNOR U28758 ( .A(n29365), .B(n29208), .Z(n29368) );
  IV U28759 ( .A(n29211), .Z(n29208) );
  XOR U28760 ( .A(n29369), .B(n29370), .Z(n29211) );
  AND U28761 ( .A(n109), .B(n29371), .Z(n29370) );
  XNOR U28762 ( .A(n29372), .B(n29369), .Z(n29371) );
  XOR U28763 ( .A(n29212), .B(n29365), .Z(n29367) );
  XOR U28764 ( .A(n29373), .B(n29374), .Z(n29212) );
  AND U28765 ( .A(n117), .B(n29332), .Z(n29374) );
  XOR U28766 ( .A(n29373), .B(n29330), .Z(n29332) );
  XOR U28767 ( .A(n29289), .B(n29375), .Z(n29365) );
  AND U28768 ( .A(n29291), .B(n29376), .Z(n29375) );
  XNOR U28769 ( .A(n29289), .B(n29258), .Z(n29376) );
  IV U28770 ( .A(n29261), .Z(n29258) );
  XOR U28771 ( .A(n29377), .B(n29378), .Z(n29261) );
  AND U28772 ( .A(n109), .B(n29379), .Z(n29378) );
  XOR U28773 ( .A(n29380), .B(n29377), .Z(n29379) );
  XOR U28774 ( .A(n29262), .B(n29289), .Z(n29291) );
  XOR U28775 ( .A(n29381), .B(n29382), .Z(n29262) );
  AND U28776 ( .A(n117), .B(n29342), .Z(n29382) );
  XOR U28777 ( .A(n29381), .B(n29340), .Z(n29342) );
  AND U28778 ( .A(n29343), .B(n29273), .Z(n29289) );
  XNOR U28779 ( .A(n29383), .B(n29384), .Z(n29273) );
  AND U28780 ( .A(n109), .B(n29385), .Z(n29384) );
  XNOR U28781 ( .A(n29386), .B(n29383), .Z(n29385) );
  XNOR U28782 ( .A(n29387), .B(n29388), .Z(n109) );
  AND U28783 ( .A(n29389), .B(n29390), .Z(n29388) );
  XOR U28784 ( .A(n29352), .B(n29387), .Z(n29390) );
  AND U28785 ( .A(n29391), .B(n29392), .Z(n29352) );
  XNOR U28786 ( .A(n29349), .B(n29387), .Z(n29389) );
  XNOR U28787 ( .A(n29393), .B(n29394), .Z(n29349) );
  AND U28788 ( .A(n113), .B(n29395), .Z(n29394) );
  XNOR U28789 ( .A(n29396), .B(n29397), .Z(n29395) );
  XOR U28790 ( .A(n29398), .B(n29399), .Z(n29387) );
  AND U28791 ( .A(n29400), .B(n29401), .Z(n29399) );
  XNOR U28792 ( .A(n29398), .B(n29391), .Z(n29401) );
  IV U28793 ( .A(n29362), .Z(n29391) );
  XOR U28794 ( .A(n29402), .B(n29403), .Z(n29362) );
  XOR U28795 ( .A(n29404), .B(n29392), .Z(n29403) );
  AND U28796 ( .A(n29372), .B(n29405), .Z(n29392) );
  AND U28797 ( .A(n29406), .B(n29407), .Z(n29404) );
  XOR U28798 ( .A(n29408), .B(n29402), .Z(n29406) );
  XNOR U28799 ( .A(n29359), .B(n29398), .Z(n29400) );
  XNOR U28800 ( .A(n29409), .B(n29410), .Z(n29359) );
  AND U28801 ( .A(n113), .B(n29411), .Z(n29410) );
  XNOR U28802 ( .A(n29412), .B(n29413), .Z(n29411) );
  XOR U28803 ( .A(n29414), .B(n29415), .Z(n29398) );
  AND U28804 ( .A(n29416), .B(n29417), .Z(n29415) );
  XNOR U28805 ( .A(n29414), .B(n29372), .Z(n29417) );
  XOR U28806 ( .A(n29418), .B(n29407), .Z(n29372) );
  XNOR U28807 ( .A(n29419), .B(n29402), .Z(n29407) );
  XOR U28808 ( .A(n29420), .B(n29421), .Z(n29402) );
  AND U28809 ( .A(n29422), .B(n29423), .Z(n29421) );
  XOR U28810 ( .A(n29424), .B(n29420), .Z(n29422) );
  XNOR U28811 ( .A(n29425), .B(n29426), .Z(n29419) );
  AND U28812 ( .A(n29427), .B(n29428), .Z(n29426) );
  XOR U28813 ( .A(n29425), .B(n29429), .Z(n29427) );
  XNOR U28814 ( .A(n29408), .B(n29405), .Z(n29418) );
  AND U28815 ( .A(n29430), .B(n29431), .Z(n29405) );
  XOR U28816 ( .A(n29432), .B(n29433), .Z(n29408) );
  AND U28817 ( .A(n29434), .B(n29435), .Z(n29433) );
  XOR U28818 ( .A(n29432), .B(n29436), .Z(n29434) );
  XNOR U28819 ( .A(n29369), .B(n29414), .Z(n29416) );
  XNOR U28820 ( .A(n29437), .B(n29438), .Z(n29369) );
  AND U28821 ( .A(n113), .B(n29439), .Z(n29438) );
  XNOR U28822 ( .A(n29440), .B(n29441), .Z(n29439) );
  XOR U28823 ( .A(n29442), .B(n29443), .Z(n29414) );
  AND U28824 ( .A(n29444), .B(n29445), .Z(n29443) );
  XNOR U28825 ( .A(n29442), .B(n29430), .Z(n29445) );
  IV U28826 ( .A(n29380), .Z(n29430) );
  XNOR U28827 ( .A(n29446), .B(n29423), .Z(n29380) );
  XNOR U28828 ( .A(n29447), .B(n29429), .Z(n29423) );
  XOR U28829 ( .A(n29448), .B(n29449), .Z(n29429) );
  NOR U28830 ( .A(n29450), .B(n29451), .Z(n29449) );
  XNOR U28831 ( .A(n29448), .B(n29452), .Z(n29450) );
  XNOR U28832 ( .A(n29428), .B(n29420), .Z(n29447) );
  XOR U28833 ( .A(n29453), .B(n29454), .Z(n29420) );
  AND U28834 ( .A(n29455), .B(n29456), .Z(n29454) );
  XNOR U28835 ( .A(n29453), .B(n29457), .Z(n29455) );
  XNOR U28836 ( .A(n29458), .B(n29425), .Z(n29428) );
  XOR U28837 ( .A(n29459), .B(n29460), .Z(n29425) );
  AND U28838 ( .A(n29461), .B(n29462), .Z(n29460) );
  XOR U28839 ( .A(n29459), .B(n29463), .Z(n29461) );
  XNOR U28840 ( .A(n29464), .B(n29465), .Z(n29458) );
  NOR U28841 ( .A(n29466), .B(n29467), .Z(n29465) );
  XOR U28842 ( .A(n29464), .B(n29468), .Z(n29466) );
  XNOR U28843 ( .A(n29424), .B(n29431), .Z(n29446) );
  NOR U28844 ( .A(n29386), .B(n29469), .Z(n29431) );
  XOR U28845 ( .A(n29436), .B(n29435), .Z(n29424) );
  XNOR U28846 ( .A(n29470), .B(n29432), .Z(n29435) );
  XOR U28847 ( .A(n29471), .B(n29472), .Z(n29432) );
  AND U28848 ( .A(n29473), .B(n29474), .Z(n29472) );
  XOR U28849 ( .A(n29471), .B(n29475), .Z(n29473) );
  XNOR U28850 ( .A(n29476), .B(n29477), .Z(n29470) );
  NOR U28851 ( .A(n29478), .B(n29479), .Z(n29477) );
  XNOR U28852 ( .A(n29476), .B(n29480), .Z(n29478) );
  XOR U28853 ( .A(n29481), .B(n29482), .Z(n29436) );
  NOR U28854 ( .A(n29483), .B(n29484), .Z(n29482) );
  XNOR U28855 ( .A(n29481), .B(n29485), .Z(n29483) );
  XNOR U28856 ( .A(n29377), .B(n29442), .Z(n29444) );
  XNOR U28857 ( .A(n29486), .B(n29487), .Z(n29377) );
  AND U28858 ( .A(n113), .B(n29488), .Z(n29487) );
  XNOR U28859 ( .A(n29489), .B(n29490), .Z(n29488) );
  AND U28860 ( .A(n29383), .B(n29386), .Z(n29442) );
  XOR U28861 ( .A(n29491), .B(n29469), .Z(n29386) );
  XNOR U28862 ( .A(p_input[2048]), .B(p_input[32]), .Z(n29469) );
  XOR U28863 ( .A(n29457), .B(n29456), .Z(n29491) );
  XNOR U28864 ( .A(n29492), .B(n29463), .Z(n29456) );
  XNOR U28865 ( .A(n29452), .B(n29451), .Z(n29463) );
  XOR U28866 ( .A(n29493), .B(n29448), .Z(n29451) );
  XNOR U28867 ( .A(n29266), .B(p_input[42]), .Z(n29448) );
  XNOR U28868 ( .A(p_input[2059]), .B(p_input[43]), .Z(n29493) );
  XOR U28869 ( .A(p_input[2060]), .B(p_input[44]), .Z(n29452) );
  XNOR U28870 ( .A(n29462), .B(n29453), .Z(n29492) );
  XNOR U28871 ( .A(n29494), .B(p_input[33]), .Z(n29453) );
  XOR U28872 ( .A(n29495), .B(n29468), .Z(n29462) );
  XNOR U28873 ( .A(p_input[2063]), .B(p_input[47]), .Z(n29468) );
  XOR U28874 ( .A(n29459), .B(n29467), .Z(n29495) );
  XOR U28875 ( .A(n29496), .B(n29464), .Z(n29467) );
  XOR U28876 ( .A(p_input[2061]), .B(p_input[45]), .Z(n29464) );
  XNOR U28877 ( .A(p_input[2062]), .B(p_input[46]), .Z(n29496) );
  XNOR U28878 ( .A(n29036), .B(p_input[41]), .Z(n29459) );
  XNOR U28879 ( .A(n29475), .B(n29474), .Z(n29457) );
  XNOR U28880 ( .A(n29497), .B(n29480), .Z(n29474) );
  XOR U28881 ( .A(p_input[2056]), .B(p_input[40]), .Z(n29480) );
  XOR U28882 ( .A(n29471), .B(n29479), .Z(n29497) );
  XOR U28883 ( .A(n29498), .B(n29476), .Z(n29479) );
  XOR U28884 ( .A(p_input[2054]), .B(p_input[38]), .Z(n29476) );
  XNOR U28885 ( .A(p_input[2055]), .B(p_input[39]), .Z(n29498) );
  XNOR U28886 ( .A(n29039), .B(p_input[34]), .Z(n29471) );
  XNOR U28887 ( .A(n29485), .B(n29484), .Z(n29475) );
  XOR U28888 ( .A(n29499), .B(n29481), .Z(n29484) );
  XOR U28889 ( .A(p_input[2051]), .B(p_input[35]), .Z(n29481) );
  XNOR U28890 ( .A(p_input[2052]), .B(p_input[36]), .Z(n29499) );
  XOR U28891 ( .A(p_input[2053]), .B(p_input[37]), .Z(n29485) );
  XNOR U28892 ( .A(n29500), .B(n29501), .Z(n29383) );
  AND U28893 ( .A(n113), .B(n29502), .Z(n29501) );
  XNOR U28894 ( .A(n29503), .B(n29504), .Z(n113) );
  AND U28895 ( .A(n29505), .B(n29506), .Z(n29504) );
  XOR U28896 ( .A(n29397), .B(n29503), .Z(n29506) );
  XNOR U28897 ( .A(n29507), .B(n29503), .Z(n29505) );
  XOR U28898 ( .A(n29508), .B(n29509), .Z(n29503) );
  AND U28899 ( .A(n29510), .B(n29511), .Z(n29509) );
  XOR U28900 ( .A(n29412), .B(n29508), .Z(n29511) );
  XOR U28901 ( .A(n29508), .B(n29413), .Z(n29510) );
  XOR U28902 ( .A(n29512), .B(n29513), .Z(n29508) );
  AND U28903 ( .A(n29514), .B(n29515), .Z(n29513) );
  XOR U28904 ( .A(n29440), .B(n29512), .Z(n29515) );
  XOR U28905 ( .A(n29512), .B(n29441), .Z(n29514) );
  XOR U28906 ( .A(n29516), .B(n29517), .Z(n29512) );
  AND U28907 ( .A(n29518), .B(n29519), .Z(n29517) );
  XOR U28908 ( .A(n29516), .B(n29489), .Z(n29519) );
  XNOR U28909 ( .A(n29520), .B(n29521), .Z(n29343) );
  AND U28910 ( .A(n117), .B(n29522), .Z(n29521) );
  XNOR U28911 ( .A(n29523), .B(n29524), .Z(n117) );
  AND U28912 ( .A(n29525), .B(n29526), .Z(n29524) );
  XOR U28913 ( .A(n29523), .B(n29353), .Z(n29526) );
  XNOR U28914 ( .A(n29523), .B(n29313), .Z(n29525) );
  XOR U28915 ( .A(n29527), .B(n29528), .Z(n29523) );
  AND U28916 ( .A(n29529), .B(n29530), .Z(n29528) );
  XOR U28917 ( .A(n29527), .B(n29321), .Z(n29529) );
  XOR U28918 ( .A(n29531), .B(n29532), .Z(n29304) );
  AND U28919 ( .A(n121), .B(n29522), .Z(n29532) );
  XNOR U28920 ( .A(n29520), .B(n29531), .Z(n29522) );
  XNOR U28921 ( .A(n29533), .B(n29534), .Z(n121) );
  AND U28922 ( .A(n29535), .B(n29536), .Z(n29534) );
  XNOR U28923 ( .A(n29537), .B(n29533), .Z(n29536) );
  IV U28924 ( .A(n29353), .Z(n29537) );
  XOR U28925 ( .A(n29507), .B(n29538), .Z(n29353) );
  AND U28926 ( .A(n124), .B(n29539), .Z(n29538) );
  XOR U28927 ( .A(n29396), .B(n29393), .Z(n29539) );
  IV U28928 ( .A(n29507), .Z(n29396) );
  XNOR U28929 ( .A(n29313), .B(n29533), .Z(n29535) );
  XOR U28930 ( .A(n29540), .B(n29541), .Z(n29313) );
  AND U28931 ( .A(n140), .B(n29542), .Z(n29541) );
  XOR U28932 ( .A(n29527), .B(n29543), .Z(n29533) );
  AND U28933 ( .A(n29544), .B(n29530), .Z(n29543) );
  XNOR U28934 ( .A(n29363), .B(n29527), .Z(n29530) );
  XOR U28935 ( .A(n29413), .B(n29545), .Z(n29363) );
  AND U28936 ( .A(n124), .B(n29546), .Z(n29545) );
  XOR U28937 ( .A(n29409), .B(n29413), .Z(n29546) );
  XNOR U28938 ( .A(n29547), .B(n29527), .Z(n29544) );
  IV U28939 ( .A(n29321), .Z(n29547) );
  XOR U28940 ( .A(n29548), .B(n29549), .Z(n29321) );
  AND U28941 ( .A(n140), .B(n29550), .Z(n29549) );
  XOR U28942 ( .A(n29551), .B(n29552), .Z(n29527) );
  AND U28943 ( .A(n29553), .B(n29554), .Z(n29552) );
  XNOR U28944 ( .A(n29373), .B(n29551), .Z(n29554) );
  XOR U28945 ( .A(n29441), .B(n29555), .Z(n29373) );
  AND U28946 ( .A(n124), .B(n29556), .Z(n29555) );
  XOR U28947 ( .A(n29437), .B(n29441), .Z(n29556) );
  XOR U28948 ( .A(n29551), .B(n29330), .Z(n29553) );
  XOR U28949 ( .A(n29557), .B(n29558), .Z(n29330) );
  AND U28950 ( .A(n140), .B(n29559), .Z(n29558) );
  XOR U28951 ( .A(n29560), .B(n29561), .Z(n29551) );
  AND U28952 ( .A(n29562), .B(n29563), .Z(n29561) );
  XNOR U28953 ( .A(n29560), .B(n29381), .Z(n29563) );
  XOR U28954 ( .A(n29490), .B(n29564), .Z(n29381) );
  AND U28955 ( .A(n124), .B(n29565), .Z(n29564) );
  XOR U28956 ( .A(n29486), .B(n29490), .Z(n29565) );
  XNOR U28957 ( .A(n29566), .B(n29560), .Z(n29562) );
  IV U28958 ( .A(n29340), .Z(n29566) );
  XOR U28959 ( .A(n29567), .B(n29568), .Z(n29340) );
  AND U28960 ( .A(n140), .B(n29569), .Z(n29568) );
  AND U28961 ( .A(n29531), .B(n29520), .Z(n29560) );
  XNOR U28962 ( .A(n29570), .B(n29571), .Z(n29520) );
  AND U28963 ( .A(n124), .B(n29502), .Z(n29571) );
  XNOR U28964 ( .A(n29500), .B(n29570), .Z(n29502) );
  XNOR U28965 ( .A(n29572), .B(n29573), .Z(n124) );
  AND U28966 ( .A(n29574), .B(n29575), .Z(n29573) );
  XNOR U28967 ( .A(n29572), .B(n29393), .Z(n29575) );
  IV U28968 ( .A(n29397), .Z(n29393) );
  XOR U28969 ( .A(n29576), .B(n29577), .Z(n29397) );
  AND U28970 ( .A(n128), .B(n29578), .Z(n29577) );
  XOR U28971 ( .A(n29579), .B(n29576), .Z(n29578) );
  XNOR U28972 ( .A(n29572), .B(n29507), .Z(n29574) );
  XOR U28973 ( .A(n29580), .B(n29581), .Z(n29507) );
  AND U28974 ( .A(n136), .B(n29542), .Z(n29581) );
  XOR U28975 ( .A(n29540), .B(n29580), .Z(n29542) );
  XOR U28976 ( .A(n29582), .B(n29583), .Z(n29572) );
  AND U28977 ( .A(n29584), .B(n29585), .Z(n29583) );
  XNOR U28978 ( .A(n29582), .B(n29409), .Z(n29585) );
  IV U28979 ( .A(n29412), .Z(n29409) );
  XOR U28980 ( .A(n29586), .B(n29587), .Z(n29412) );
  AND U28981 ( .A(n128), .B(n29588), .Z(n29587) );
  XOR U28982 ( .A(n29589), .B(n29586), .Z(n29588) );
  XOR U28983 ( .A(n29413), .B(n29582), .Z(n29584) );
  XOR U28984 ( .A(n29590), .B(n29591), .Z(n29413) );
  AND U28985 ( .A(n136), .B(n29550), .Z(n29591) );
  XOR U28986 ( .A(n29590), .B(n29548), .Z(n29550) );
  XOR U28987 ( .A(n29592), .B(n29593), .Z(n29582) );
  AND U28988 ( .A(n29594), .B(n29595), .Z(n29593) );
  XNOR U28989 ( .A(n29592), .B(n29437), .Z(n29595) );
  IV U28990 ( .A(n29440), .Z(n29437) );
  XOR U28991 ( .A(n29596), .B(n29597), .Z(n29440) );
  AND U28992 ( .A(n128), .B(n29598), .Z(n29597) );
  XNOR U28993 ( .A(n29599), .B(n29596), .Z(n29598) );
  XOR U28994 ( .A(n29441), .B(n29592), .Z(n29594) );
  XOR U28995 ( .A(n29600), .B(n29601), .Z(n29441) );
  AND U28996 ( .A(n136), .B(n29559), .Z(n29601) );
  XOR U28997 ( .A(n29600), .B(n29557), .Z(n29559) );
  XOR U28998 ( .A(n29516), .B(n29602), .Z(n29592) );
  AND U28999 ( .A(n29518), .B(n29603), .Z(n29602) );
  XNOR U29000 ( .A(n29516), .B(n29486), .Z(n29603) );
  IV U29001 ( .A(n29489), .Z(n29486) );
  XOR U29002 ( .A(n29604), .B(n29605), .Z(n29489) );
  AND U29003 ( .A(n128), .B(n29606), .Z(n29605) );
  XOR U29004 ( .A(n29607), .B(n29604), .Z(n29606) );
  XOR U29005 ( .A(n29490), .B(n29516), .Z(n29518) );
  XOR U29006 ( .A(n29608), .B(n29609), .Z(n29490) );
  AND U29007 ( .A(n136), .B(n29569), .Z(n29609) );
  XOR U29008 ( .A(n29608), .B(n29567), .Z(n29569) );
  AND U29009 ( .A(n29570), .B(n29500), .Z(n29516) );
  XNOR U29010 ( .A(n29610), .B(n29611), .Z(n29500) );
  AND U29011 ( .A(n128), .B(n29612), .Z(n29611) );
  XNOR U29012 ( .A(n29613), .B(n29610), .Z(n29612) );
  XNOR U29013 ( .A(n29614), .B(n29615), .Z(n128) );
  AND U29014 ( .A(n29616), .B(n29617), .Z(n29615) );
  XOR U29015 ( .A(n29579), .B(n29614), .Z(n29617) );
  AND U29016 ( .A(n29618), .B(n29619), .Z(n29579) );
  XNOR U29017 ( .A(n29576), .B(n29614), .Z(n29616) );
  XNOR U29018 ( .A(n29620), .B(n29621), .Z(n29576) );
  AND U29019 ( .A(n132), .B(n29622), .Z(n29621) );
  XNOR U29020 ( .A(n29623), .B(n29624), .Z(n29622) );
  XOR U29021 ( .A(n29625), .B(n29626), .Z(n29614) );
  AND U29022 ( .A(n29627), .B(n29628), .Z(n29626) );
  XNOR U29023 ( .A(n29625), .B(n29618), .Z(n29628) );
  IV U29024 ( .A(n29589), .Z(n29618) );
  XOR U29025 ( .A(n29629), .B(n29630), .Z(n29589) );
  XOR U29026 ( .A(n29631), .B(n29619), .Z(n29630) );
  AND U29027 ( .A(n29599), .B(n29632), .Z(n29619) );
  AND U29028 ( .A(n29633), .B(n29634), .Z(n29631) );
  XOR U29029 ( .A(n29635), .B(n29629), .Z(n29633) );
  XNOR U29030 ( .A(n29586), .B(n29625), .Z(n29627) );
  XNOR U29031 ( .A(n29636), .B(n29637), .Z(n29586) );
  AND U29032 ( .A(n132), .B(n29638), .Z(n29637) );
  XNOR U29033 ( .A(n29639), .B(n29640), .Z(n29638) );
  XOR U29034 ( .A(n29641), .B(n29642), .Z(n29625) );
  AND U29035 ( .A(n29643), .B(n29644), .Z(n29642) );
  XNOR U29036 ( .A(n29641), .B(n29599), .Z(n29644) );
  XOR U29037 ( .A(n29645), .B(n29634), .Z(n29599) );
  XNOR U29038 ( .A(n29646), .B(n29629), .Z(n29634) );
  XOR U29039 ( .A(n29647), .B(n29648), .Z(n29629) );
  AND U29040 ( .A(n29649), .B(n29650), .Z(n29648) );
  XOR U29041 ( .A(n29651), .B(n29647), .Z(n29649) );
  XNOR U29042 ( .A(n29652), .B(n29653), .Z(n29646) );
  AND U29043 ( .A(n29654), .B(n29655), .Z(n29653) );
  XOR U29044 ( .A(n29652), .B(n29656), .Z(n29654) );
  XNOR U29045 ( .A(n29635), .B(n29632), .Z(n29645) );
  AND U29046 ( .A(n29657), .B(n29658), .Z(n29632) );
  XOR U29047 ( .A(n29659), .B(n29660), .Z(n29635) );
  AND U29048 ( .A(n29661), .B(n29662), .Z(n29660) );
  XOR U29049 ( .A(n29659), .B(n29663), .Z(n29661) );
  XNOR U29050 ( .A(n29596), .B(n29641), .Z(n29643) );
  XNOR U29051 ( .A(n29664), .B(n29665), .Z(n29596) );
  AND U29052 ( .A(n132), .B(n29666), .Z(n29665) );
  XNOR U29053 ( .A(n29667), .B(n29668), .Z(n29666) );
  XOR U29054 ( .A(n29669), .B(n29670), .Z(n29641) );
  AND U29055 ( .A(n29671), .B(n29672), .Z(n29670) );
  XNOR U29056 ( .A(n29669), .B(n29657), .Z(n29672) );
  IV U29057 ( .A(n29607), .Z(n29657) );
  XNOR U29058 ( .A(n29673), .B(n29650), .Z(n29607) );
  XNOR U29059 ( .A(n29674), .B(n29656), .Z(n29650) );
  XOR U29060 ( .A(n29675), .B(n29676), .Z(n29656) );
  NOR U29061 ( .A(n29677), .B(n29678), .Z(n29676) );
  XNOR U29062 ( .A(n29675), .B(n29679), .Z(n29677) );
  XNOR U29063 ( .A(n29655), .B(n29647), .Z(n29674) );
  XOR U29064 ( .A(n29680), .B(n29681), .Z(n29647) );
  AND U29065 ( .A(n29682), .B(n29683), .Z(n29681) );
  XNOR U29066 ( .A(n29680), .B(n29684), .Z(n29682) );
  XNOR U29067 ( .A(n29685), .B(n29652), .Z(n29655) );
  XOR U29068 ( .A(n29686), .B(n29687), .Z(n29652) );
  AND U29069 ( .A(n29688), .B(n29689), .Z(n29687) );
  XOR U29070 ( .A(n29686), .B(n29690), .Z(n29688) );
  XNOR U29071 ( .A(n29691), .B(n29692), .Z(n29685) );
  NOR U29072 ( .A(n29693), .B(n29694), .Z(n29692) );
  XOR U29073 ( .A(n29691), .B(n29695), .Z(n29693) );
  XNOR U29074 ( .A(n29651), .B(n29658), .Z(n29673) );
  NOR U29075 ( .A(n29613), .B(n29696), .Z(n29658) );
  XOR U29076 ( .A(n29663), .B(n29662), .Z(n29651) );
  XNOR U29077 ( .A(n29697), .B(n29659), .Z(n29662) );
  XOR U29078 ( .A(n29698), .B(n29699), .Z(n29659) );
  AND U29079 ( .A(n29700), .B(n29701), .Z(n29699) );
  XOR U29080 ( .A(n29698), .B(n29702), .Z(n29700) );
  XNOR U29081 ( .A(n29703), .B(n29704), .Z(n29697) );
  NOR U29082 ( .A(n29705), .B(n29706), .Z(n29704) );
  XNOR U29083 ( .A(n29703), .B(n29707), .Z(n29705) );
  XOR U29084 ( .A(n29708), .B(n29709), .Z(n29663) );
  NOR U29085 ( .A(n29710), .B(n29711), .Z(n29709) );
  XNOR U29086 ( .A(n29708), .B(n29712), .Z(n29710) );
  XNOR U29087 ( .A(n29604), .B(n29669), .Z(n29671) );
  XNOR U29088 ( .A(n29713), .B(n29714), .Z(n29604) );
  AND U29089 ( .A(n132), .B(n29715), .Z(n29714) );
  XNOR U29090 ( .A(n29716), .B(n29717), .Z(n29715) );
  AND U29091 ( .A(n29610), .B(n29613), .Z(n29669) );
  XOR U29092 ( .A(n29718), .B(n29696), .Z(n29613) );
  XNOR U29093 ( .A(p_input[2048]), .B(p_input[48]), .Z(n29696) );
  XOR U29094 ( .A(n29684), .B(n29683), .Z(n29718) );
  XNOR U29095 ( .A(n29719), .B(n29690), .Z(n29683) );
  XNOR U29096 ( .A(n29679), .B(n29678), .Z(n29690) );
  XOR U29097 ( .A(n29720), .B(n29675), .Z(n29678) );
  XNOR U29098 ( .A(n29266), .B(p_input[58]), .Z(n29675) );
  XNOR U29099 ( .A(p_input[2059]), .B(p_input[59]), .Z(n29720) );
  XOR U29100 ( .A(p_input[2060]), .B(p_input[60]), .Z(n29679) );
  XNOR U29101 ( .A(n29689), .B(n29680), .Z(n29719) );
  XNOR U29102 ( .A(n29494), .B(p_input[49]), .Z(n29680) );
  XOR U29103 ( .A(n29721), .B(n29695), .Z(n29689) );
  XNOR U29104 ( .A(p_input[2063]), .B(p_input[63]), .Z(n29695) );
  XOR U29105 ( .A(n29686), .B(n29694), .Z(n29721) );
  XOR U29106 ( .A(n29722), .B(n29691), .Z(n29694) );
  XOR U29107 ( .A(p_input[2061]), .B(p_input[61]), .Z(n29691) );
  XNOR U29108 ( .A(p_input[2062]), .B(p_input[62]), .Z(n29722) );
  XNOR U29109 ( .A(n29036), .B(p_input[57]), .Z(n29686) );
  XNOR U29110 ( .A(n29702), .B(n29701), .Z(n29684) );
  XNOR U29111 ( .A(n29723), .B(n29707), .Z(n29701) );
  XOR U29112 ( .A(p_input[2056]), .B(p_input[56]), .Z(n29707) );
  XOR U29113 ( .A(n29698), .B(n29706), .Z(n29723) );
  XOR U29114 ( .A(n29724), .B(n29703), .Z(n29706) );
  XOR U29115 ( .A(p_input[2054]), .B(p_input[54]), .Z(n29703) );
  XNOR U29116 ( .A(p_input[2055]), .B(p_input[55]), .Z(n29724) );
  XNOR U29117 ( .A(n29039), .B(p_input[50]), .Z(n29698) );
  XNOR U29118 ( .A(n29712), .B(n29711), .Z(n29702) );
  XOR U29119 ( .A(n29725), .B(n29708), .Z(n29711) );
  XOR U29120 ( .A(p_input[2051]), .B(p_input[51]), .Z(n29708) );
  XNOR U29121 ( .A(p_input[2052]), .B(p_input[52]), .Z(n29725) );
  XOR U29122 ( .A(p_input[2053]), .B(p_input[53]), .Z(n29712) );
  XNOR U29123 ( .A(n29726), .B(n29727), .Z(n29610) );
  AND U29124 ( .A(n132), .B(n29728), .Z(n29727) );
  XNOR U29125 ( .A(n29729), .B(n29730), .Z(n132) );
  AND U29126 ( .A(n29731), .B(n29732), .Z(n29730) );
  XOR U29127 ( .A(n29624), .B(n29729), .Z(n29732) );
  XNOR U29128 ( .A(n29733), .B(n29729), .Z(n29731) );
  XOR U29129 ( .A(n29734), .B(n29735), .Z(n29729) );
  AND U29130 ( .A(n29736), .B(n29737), .Z(n29735) );
  XOR U29131 ( .A(n29639), .B(n29734), .Z(n29737) );
  XOR U29132 ( .A(n29734), .B(n29640), .Z(n29736) );
  XOR U29133 ( .A(n29738), .B(n29739), .Z(n29734) );
  AND U29134 ( .A(n29740), .B(n29741), .Z(n29739) );
  XOR U29135 ( .A(n29667), .B(n29738), .Z(n29741) );
  XOR U29136 ( .A(n29738), .B(n29668), .Z(n29740) );
  XOR U29137 ( .A(n29742), .B(n29743), .Z(n29738) );
  AND U29138 ( .A(n29744), .B(n29745), .Z(n29743) );
  XOR U29139 ( .A(n29742), .B(n29716), .Z(n29745) );
  XNOR U29140 ( .A(n29746), .B(n29747), .Z(n29570) );
  AND U29141 ( .A(n136), .B(n29748), .Z(n29747) );
  XNOR U29142 ( .A(n29749), .B(n29750), .Z(n136) );
  AND U29143 ( .A(n29751), .B(n29752), .Z(n29750) );
  XOR U29144 ( .A(n29749), .B(n29580), .Z(n29752) );
  XNOR U29145 ( .A(n29749), .B(n29540), .Z(n29751) );
  XOR U29146 ( .A(n29753), .B(n29754), .Z(n29749) );
  AND U29147 ( .A(n29755), .B(n29756), .Z(n29754) );
  XOR U29148 ( .A(n29753), .B(n29548), .Z(n29755) );
  XOR U29149 ( .A(n29757), .B(n29758), .Z(n29531) );
  AND U29150 ( .A(n140), .B(n29748), .Z(n29758) );
  XNOR U29151 ( .A(n29746), .B(n29757), .Z(n29748) );
  XNOR U29152 ( .A(n29759), .B(n29760), .Z(n140) );
  AND U29153 ( .A(n29761), .B(n29762), .Z(n29760) );
  XNOR U29154 ( .A(n29763), .B(n29759), .Z(n29762) );
  IV U29155 ( .A(n29580), .Z(n29763) );
  XOR U29156 ( .A(n29733), .B(n29764), .Z(n29580) );
  AND U29157 ( .A(n143), .B(n29765), .Z(n29764) );
  XOR U29158 ( .A(n29623), .B(n29620), .Z(n29765) );
  IV U29159 ( .A(n29733), .Z(n29623) );
  XNOR U29160 ( .A(n29540), .B(n29759), .Z(n29761) );
  XOR U29161 ( .A(n29766), .B(n29767), .Z(n29540) );
  AND U29162 ( .A(n159), .B(n29768), .Z(n29767) );
  XOR U29163 ( .A(n29753), .B(n29769), .Z(n29759) );
  AND U29164 ( .A(n29770), .B(n29756), .Z(n29769) );
  XNOR U29165 ( .A(n29590), .B(n29753), .Z(n29756) );
  XOR U29166 ( .A(n29640), .B(n29771), .Z(n29590) );
  AND U29167 ( .A(n143), .B(n29772), .Z(n29771) );
  XOR U29168 ( .A(n29636), .B(n29640), .Z(n29772) );
  XNOR U29169 ( .A(n29773), .B(n29753), .Z(n29770) );
  IV U29170 ( .A(n29548), .Z(n29773) );
  XOR U29171 ( .A(n29774), .B(n29775), .Z(n29548) );
  AND U29172 ( .A(n159), .B(n29776), .Z(n29775) );
  XOR U29173 ( .A(n29777), .B(n29778), .Z(n29753) );
  AND U29174 ( .A(n29779), .B(n29780), .Z(n29778) );
  XNOR U29175 ( .A(n29600), .B(n29777), .Z(n29780) );
  XOR U29176 ( .A(n29668), .B(n29781), .Z(n29600) );
  AND U29177 ( .A(n143), .B(n29782), .Z(n29781) );
  XOR U29178 ( .A(n29664), .B(n29668), .Z(n29782) );
  XOR U29179 ( .A(n29777), .B(n29557), .Z(n29779) );
  XOR U29180 ( .A(n29783), .B(n29784), .Z(n29557) );
  AND U29181 ( .A(n159), .B(n29785), .Z(n29784) );
  XOR U29182 ( .A(n29786), .B(n29787), .Z(n29777) );
  AND U29183 ( .A(n29788), .B(n29789), .Z(n29787) );
  XNOR U29184 ( .A(n29786), .B(n29608), .Z(n29789) );
  XOR U29185 ( .A(n29717), .B(n29790), .Z(n29608) );
  AND U29186 ( .A(n143), .B(n29791), .Z(n29790) );
  XOR U29187 ( .A(n29713), .B(n29717), .Z(n29791) );
  XNOR U29188 ( .A(n29792), .B(n29786), .Z(n29788) );
  IV U29189 ( .A(n29567), .Z(n29792) );
  XOR U29190 ( .A(n29793), .B(n29794), .Z(n29567) );
  AND U29191 ( .A(n159), .B(n29795), .Z(n29794) );
  AND U29192 ( .A(n29757), .B(n29746), .Z(n29786) );
  XNOR U29193 ( .A(n29796), .B(n29797), .Z(n29746) );
  AND U29194 ( .A(n143), .B(n29728), .Z(n29797) );
  XNOR U29195 ( .A(n29726), .B(n29796), .Z(n29728) );
  XNOR U29196 ( .A(n29798), .B(n29799), .Z(n143) );
  AND U29197 ( .A(n29800), .B(n29801), .Z(n29799) );
  XNOR U29198 ( .A(n29798), .B(n29620), .Z(n29801) );
  IV U29199 ( .A(n29624), .Z(n29620) );
  XOR U29200 ( .A(n29802), .B(n29803), .Z(n29624) );
  AND U29201 ( .A(n147), .B(n29804), .Z(n29803) );
  XOR U29202 ( .A(n29805), .B(n29802), .Z(n29804) );
  XNOR U29203 ( .A(n29798), .B(n29733), .Z(n29800) );
  XOR U29204 ( .A(n29806), .B(n29807), .Z(n29733) );
  AND U29205 ( .A(n155), .B(n29768), .Z(n29807) );
  XOR U29206 ( .A(n29766), .B(n29806), .Z(n29768) );
  XOR U29207 ( .A(n29808), .B(n29809), .Z(n29798) );
  AND U29208 ( .A(n29810), .B(n29811), .Z(n29809) );
  XNOR U29209 ( .A(n29808), .B(n29636), .Z(n29811) );
  IV U29210 ( .A(n29639), .Z(n29636) );
  XOR U29211 ( .A(n29812), .B(n29813), .Z(n29639) );
  AND U29212 ( .A(n147), .B(n29814), .Z(n29813) );
  XOR U29213 ( .A(n29815), .B(n29812), .Z(n29814) );
  XOR U29214 ( .A(n29640), .B(n29808), .Z(n29810) );
  XOR U29215 ( .A(n29816), .B(n29817), .Z(n29640) );
  AND U29216 ( .A(n155), .B(n29776), .Z(n29817) );
  XOR U29217 ( .A(n29816), .B(n29774), .Z(n29776) );
  XOR U29218 ( .A(n29818), .B(n29819), .Z(n29808) );
  AND U29219 ( .A(n29820), .B(n29821), .Z(n29819) );
  XNOR U29220 ( .A(n29818), .B(n29664), .Z(n29821) );
  IV U29221 ( .A(n29667), .Z(n29664) );
  XOR U29222 ( .A(n29822), .B(n29823), .Z(n29667) );
  AND U29223 ( .A(n147), .B(n29824), .Z(n29823) );
  XNOR U29224 ( .A(n29825), .B(n29822), .Z(n29824) );
  XOR U29225 ( .A(n29668), .B(n29818), .Z(n29820) );
  XOR U29226 ( .A(n29826), .B(n29827), .Z(n29668) );
  AND U29227 ( .A(n155), .B(n29785), .Z(n29827) );
  XOR U29228 ( .A(n29826), .B(n29783), .Z(n29785) );
  XOR U29229 ( .A(n29742), .B(n29828), .Z(n29818) );
  AND U29230 ( .A(n29744), .B(n29829), .Z(n29828) );
  XNOR U29231 ( .A(n29742), .B(n29713), .Z(n29829) );
  IV U29232 ( .A(n29716), .Z(n29713) );
  XOR U29233 ( .A(n29830), .B(n29831), .Z(n29716) );
  AND U29234 ( .A(n147), .B(n29832), .Z(n29831) );
  XOR U29235 ( .A(n29833), .B(n29830), .Z(n29832) );
  XOR U29236 ( .A(n29717), .B(n29742), .Z(n29744) );
  XOR U29237 ( .A(n29834), .B(n29835), .Z(n29717) );
  AND U29238 ( .A(n155), .B(n29795), .Z(n29835) );
  XOR U29239 ( .A(n29834), .B(n29793), .Z(n29795) );
  AND U29240 ( .A(n29796), .B(n29726), .Z(n29742) );
  XNOR U29241 ( .A(n29836), .B(n29837), .Z(n29726) );
  AND U29242 ( .A(n147), .B(n29838), .Z(n29837) );
  XNOR U29243 ( .A(n29839), .B(n29836), .Z(n29838) );
  XNOR U29244 ( .A(n29840), .B(n29841), .Z(n147) );
  AND U29245 ( .A(n29842), .B(n29843), .Z(n29841) );
  XOR U29246 ( .A(n29805), .B(n29840), .Z(n29843) );
  AND U29247 ( .A(n29844), .B(n29845), .Z(n29805) );
  XNOR U29248 ( .A(n29802), .B(n29840), .Z(n29842) );
  XNOR U29249 ( .A(n29846), .B(n29847), .Z(n29802) );
  AND U29250 ( .A(n151), .B(n29848), .Z(n29847) );
  XNOR U29251 ( .A(n29849), .B(n29850), .Z(n29848) );
  XOR U29252 ( .A(n29851), .B(n29852), .Z(n29840) );
  AND U29253 ( .A(n29853), .B(n29854), .Z(n29852) );
  XNOR U29254 ( .A(n29851), .B(n29844), .Z(n29854) );
  IV U29255 ( .A(n29815), .Z(n29844) );
  XOR U29256 ( .A(n29855), .B(n29856), .Z(n29815) );
  XOR U29257 ( .A(n29857), .B(n29845), .Z(n29856) );
  AND U29258 ( .A(n29825), .B(n29858), .Z(n29845) );
  AND U29259 ( .A(n29859), .B(n29860), .Z(n29857) );
  XOR U29260 ( .A(n29861), .B(n29855), .Z(n29859) );
  XNOR U29261 ( .A(n29812), .B(n29851), .Z(n29853) );
  XNOR U29262 ( .A(n29862), .B(n29863), .Z(n29812) );
  AND U29263 ( .A(n151), .B(n29864), .Z(n29863) );
  XNOR U29264 ( .A(n29865), .B(n29866), .Z(n29864) );
  XOR U29265 ( .A(n29867), .B(n29868), .Z(n29851) );
  AND U29266 ( .A(n29869), .B(n29870), .Z(n29868) );
  XNOR U29267 ( .A(n29867), .B(n29825), .Z(n29870) );
  XOR U29268 ( .A(n29871), .B(n29860), .Z(n29825) );
  XNOR U29269 ( .A(n29872), .B(n29855), .Z(n29860) );
  XOR U29270 ( .A(n29873), .B(n29874), .Z(n29855) );
  AND U29271 ( .A(n29875), .B(n29876), .Z(n29874) );
  XOR U29272 ( .A(n29877), .B(n29873), .Z(n29875) );
  XNOR U29273 ( .A(n29878), .B(n29879), .Z(n29872) );
  AND U29274 ( .A(n29880), .B(n29881), .Z(n29879) );
  XOR U29275 ( .A(n29878), .B(n29882), .Z(n29880) );
  XNOR U29276 ( .A(n29861), .B(n29858), .Z(n29871) );
  AND U29277 ( .A(n29883), .B(n29884), .Z(n29858) );
  XOR U29278 ( .A(n29885), .B(n29886), .Z(n29861) );
  AND U29279 ( .A(n29887), .B(n29888), .Z(n29886) );
  XOR U29280 ( .A(n29885), .B(n29889), .Z(n29887) );
  XNOR U29281 ( .A(n29822), .B(n29867), .Z(n29869) );
  XNOR U29282 ( .A(n29890), .B(n29891), .Z(n29822) );
  AND U29283 ( .A(n151), .B(n29892), .Z(n29891) );
  XNOR U29284 ( .A(n29893), .B(n29894), .Z(n29892) );
  XOR U29285 ( .A(n29895), .B(n29896), .Z(n29867) );
  AND U29286 ( .A(n29897), .B(n29898), .Z(n29896) );
  XNOR U29287 ( .A(n29895), .B(n29883), .Z(n29898) );
  IV U29288 ( .A(n29833), .Z(n29883) );
  XNOR U29289 ( .A(n29899), .B(n29876), .Z(n29833) );
  XNOR U29290 ( .A(n29900), .B(n29882), .Z(n29876) );
  XOR U29291 ( .A(n29901), .B(n29902), .Z(n29882) );
  NOR U29292 ( .A(n29903), .B(n29904), .Z(n29902) );
  XNOR U29293 ( .A(n29901), .B(n29905), .Z(n29903) );
  XNOR U29294 ( .A(n29881), .B(n29873), .Z(n29900) );
  XOR U29295 ( .A(n29906), .B(n29907), .Z(n29873) );
  AND U29296 ( .A(n29908), .B(n29909), .Z(n29907) );
  XNOR U29297 ( .A(n29906), .B(n29910), .Z(n29908) );
  XNOR U29298 ( .A(n29911), .B(n29878), .Z(n29881) );
  XOR U29299 ( .A(n29912), .B(n29913), .Z(n29878) );
  AND U29300 ( .A(n29914), .B(n29915), .Z(n29913) );
  XOR U29301 ( .A(n29912), .B(n29916), .Z(n29914) );
  XNOR U29302 ( .A(n29917), .B(n29918), .Z(n29911) );
  NOR U29303 ( .A(n29919), .B(n29920), .Z(n29918) );
  XOR U29304 ( .A(n29917), .B(n29921), .Z(n29919) );
  XNOR U29305 ( .A(n29877), .B(n29884), .Z(n29899) );
  NOR U29306 ( .A(n29839), .B(n29922), .Z(n29884) );
  XOR U29307 ( .A(n29889), .B(n29888), .Z(n29877) );
  XNOR U29308 ( .A(n29923), .B(n29885), .Z(n29888) );
  XOR U29309 ( .A(n29924), .B(n29925), .Z(n29885) );
  AND U29310 ( .A(n29926), .B(n29927), .Z(n29925) );
  XOR U29311 ( .A(n29924), .B(n29928), .Z(n29926) );
  XNOR U29312 ( .A(n29929), .B(n29930), .Z(n29923) );
  NOR U29313 ( .A(n29931), .B(n29932), .Z(n29930) );
  XNOR U29314 ( .A(n29929), .B(n29933), .Z(n29931) );
  XOR U29315 ( .A(n29934), .B(n29935), .Z(n29889) );
  NOR U29316 ( .A(n29936), .B(n29937), .Z(n29935) );
  XNOR U29317 ( .A(n29934), .B(n29938), .Z(n29936) );
  XNOR U29318 ( .A(n29830), .B(n29895), .Z(n29897) );
  XNOR U29319 ( .A(n29939), .B(n29940), .Z(n29830) );
  AND U29320 ( .A(n151), .B(n29941), .Z(n29940) );
  XNOR U29321 ( .A(n29942), .B(n29943), .Z(n29941) );
  AND U29322 ( .A(n29836), .B(n29839), .Z(n29895) );
  XOR U29323 ( .A(n29944), .B(n29922), .Z(n29839) );
  XNOR U29324 ( .A(p_input[2048]), .B(p_input[64]), .Z(n29922) );
  XOR U29325 ( .A(n29910), .B(n29909), .Z(n29944) );
  XNOR U29326 ( .A(n29945), .B(n29916), .Z(n29909) );
  XNOR U29327 ( .A(n29905), .B(n29904), .Z(n29916) );
  XOR U29328 ( .A(n29946), .B(n29901), .Z(n29904) );
  XNOR U29329 ( .A(n29266), .B(p_input[74]), .Z(n29901) );
  XNOR U29330 ( .A(p_input[2059]), .B(p_input[75]), .Z(n29946) );
  XOR U29331 ( .A(p_input[2060]), .B(p_input[76]), .Z(n29905) );
  XNOR U29332 ( .A(n29915), .B(n29906), .Z(n29945) );
  XNOR U29333 ( .A(n29494), .B(p_input[65]), .Z(n29906) );
  XOR U29334 ( .A(n29947), .B(n29921), .Z(n29915) );
  XNOR U29335 ( .A(p_input[2063]), .B(p_input[79]), .Z(n29921) );
  XOR U29336 ( .A(n29912), .B(n29920), .Z(n29947) );
  XOR U29337 ( .A(n29948), .B(n29917), .Z(n29920) );
  XOR U29338 ( .A(p_input[2061]), .B(p_input[77]), .Z(n29917) );
  XNOR U29339 ( .A(p_input[2062]), .B(p_input[78]), .Z(n29948) );
  XNOR U29340 ( .A(n29036), .B(p_input[73]), .Z(n29912) );
  XNOR U29341 ( .A(n29928), .B(n29927), .Z(n29910) );
  XNOR U29342 ( .A(n29949), .B(n29933), .Z(n29927) );
  XOR U29343 ( .A(p_input[2056]), .B(p_input[72]), .Z(n29933) );
  XOR U29344 ( .A(n29924), .B(n29932), .Z(n29949) );
  XOR U29345 ( .A(n29950), .B(n29929), .Z(n29932) );
  XOR U29346 ( .A(p_input[2054]), .B(p_input[70]), .Z(n29929) );
  XNOR U29347 ( .A(p_input[2055]), .B(p_input[71]), .Z(n29950) );
  XNOR U29348 ( .A(n29039), .B(p_input[66]), .Z(n29924) );
  XNOR U29349 ( .A(n29938), .B(n29937), .Z(n29928) );
  XOR U29350 ( .A(n29951), .B(n29934), .Z(n29937) );
  XOR U29351 ( .A(p_input[2051]), .B(p_input[67]), .Z(n29934) );
  XNOR U29352 ( .A(p_input[2052]), .B(p_input[68]), .Z(n29951) );
  XOR U29353 ( .A(p_input[2053]), .B(p_input[69]), .Z(n29938) );
  XNOR U29354 ( .A(n29952), .B(n29953), .Z(n29836) );
  AND U29355 ( .A(n151), .B(n29954), .Z(n29953) );
  XNOR U29356 ( .A(n29955), .B(n29956), .Z(n151) );
  AND U29357 ( .A(n29957), .B(n29958), .Z(n29956) );
  XOR U29358 ( .A(n29850), .B(n29955), .Z(n29958) );
  XNOR U29359 ( .A(n29959), .B(n29955), .Z(n29957) );
  XOR U29360 ( .A(n29960), .B(n29961), .Z(n29955) );
  AND U29361 ( .A(n29962), .B(n29963), .Z(n29961) );
  XOR U29362 ( .A(n29865), .B(n29960), .Z(n29963) );
  XOR U29363 ( .A(n29960), .B(n29866), .Z(n29962) );
  XOR U29364 ( .A(n29964), .B(n29965), .Z(n29960) );
  AND U29365 ( .A(n29966), .B(n29967), .Z(n29965) );
  XOR U29366 ( .A(n29893), .B(n29964), .Z(n29967) );
  XOR U29367 ( .A(n29964), .B(n29894), .Z(n29966) );
  XOR U29368 ( .A(n29968), .B(n29969), .Z(n29964) );
  AND U29369 ( .A(n29970), .B(n29971), .Z(n29969) );
  XOR U29370 ( .A(n29968), .B(n29942), .Z(n29971) );
  XNOR U29371 ( .A(n29972), .B(n29973), .Z(n29796) );
  AND U29372 ( .A(n155), .B(n29974), .Z(n29973) );
  XNOR U29373 ( .A(n29975), .B(n29976), .Z(n155) );
  AND U29374 ( .A(n29977), .B(n29978), .Z(n29976) );
  XOR U29375 ( .A(n29975), .B(n29806), .Z(n29978) );
  XNOR U29376 ( .A(n29975), .B(n29766), .Z(n29977) );
  XOR U29377 ( .A(n29979), .B(n29980), .Z(n29975) );
  AND U29378 ( .A(n29981), .B(n29982), .Z(n29980) );
  XOR U29379 ( .A(n29979), .B(n29774), .Z(n29981) );
  XOR U29380 ( .A(n29983), .B(n29984), .Z(n29757) );
  AND U29381 ( .A(n159), .B(n29974), .Z(n29984) );
  XNOR U29382 ( .A(n29972), .B(n29983), .Z(n29974) );
  XNOR U29383 ( .A(n29985), .B(n29986), .Z(n159) );
  AND U29384 ( .A(n29987), .B(n29988), .Z(n29986) );
  XNOR U29385 ( .A(n29989), .B(n29985), .Z(n29988) );
  IV U29386 ( .A(n29806), .Z(n29989) );
  XOR U29387 ( .A(n29959), .B(n29990), .Z(n29806) );
  AND U29388 ( .A(n162), .B(n29991), .Z(n29990) );
  XOR U29389 ( .A(n29849), .B(n29846), .Z(n29991) );
  IV U29390 ( .A(n29959), .Z(n29849) );
  XNOR U29391 ( .A(n29766), .B(n29985), .Z(n29987) );
  XOR U29392 ( .A(n29992), .B(n29993), .Z(n29766) );
  AND U29393 ( .A(n178), .B(n29994), .Z(n29993) );
  XOR U29394 ( .A(n29979), .B(n29995), .Z(n29985) );
  AND U29395 ( .A(n29996), .B(n29982), .Z(n29995) );
  XNOR U29396 ( .A(n29816), .B(n29979), .Z(n29982) );
  XOR U29397 ( .A(n29866), .B(n29997), .Z(n29816) );
  AND U29398 ( .A(n162), .B(n29998), .Z(n29997) );
  XOR U29399 ( .A(n29862), .B(n29866), .Z(n29998) );
  XNOR U29400 ( .A(n29999), .B(n29979), .Z(n29996) );
  IV U29401 ( .A(n29774), .Z(n29999) );
  XOR U29402 ( .A(n30000), .B(n30001), .Z(n29774) );
  AND U29403 ( .A(n178), .B(n30002), .Z(n30001) );
  XOR U29404 ( .A(n30003), .B(n30004), .Z(n29979) );
  AND U29405 ( .A(n30005), .B(n30006), .Z(n30004) );
  XNOR U29406 ( .A(n29826), .B(n30003), .Z(n30006) );
  XOR U29407 ( .A(n29894), .B(n30007), .Z(n29826) );
  AND U29408 ( .A(n162), .B(n30008), .Z(n30007) );
  XOR U29409 ( .A(n29890), .B(n29894), .Z(n30008) );
  XOR U29410 ( .A(n30003), .B(n29783), .Z(n30005) );
  XOR U29411 ( .A(n30009), .B(n30010), .Z(n29783) );
  AND U29412 ( .A(n178), .B(n30011), .Z(n30010) );
  XOR U29413 ( .A(n30012), .B(n30013), .Z(n30003) );
  AND U29414 ( .A(n30014), .B(n30015), .Z(n30013) );
  XNOR U29415 ( .A(n30012), .B(n29834), .Z(n30015) );
  XOR U29416 ( .A(n29943), .B(n30016), .Z(n29834) );
  AND U29417 ( .A(n162), .B(n30017), .Z(n30016) );
  XOR U29418 ( .A(n29939), .B(n29943), .Z(n30017) );
  XNOR U29419 ( .A(n30018), .B(n30012), .Z(n30014) );
  IV U29420 ( .A(n29793), .Z(n30018) );
  XOR U29421 ( .A(n30019), .B(n30020), .Z(n29793) );
  AND U29422 ( .A(n178), .B(n30021), .Z(n30020) );
  AND U29423 ( .A(n29983), .B(n29972), .Z(n30012) );
  XNOR U29424 ( .A(n30022), .B(n30023), .Z(n29972) );
  AND U29425 ( .A(n162), .B(n29954), .Z(n30023) );
  XNOR U29426 ( .A(n29952), .B(n30022), .Z(n29954) );
  XNOR U29427 ( .A(n30024), .B(n30025), .Z(n162) );
  AND U29428 ( .A(n30026), .B(n30027), .Z(n30025) );
  XNOR U29429 ( .A(n30024), .B(n29846), .Z(n30027) );
  IV U29430 ( .A(n29850), .Z(n29846) );
  XOR U29431 ( .A(n30028), .B(n30029), .Z(n29850) );
  AND U29432 ( .A(n166), .B(n30030), .Z(n30029) );
  XOR U29433 ( .A(n30031), .B(n30028), .Z(n30030) );
  XNOR U29434 ( .A(n30024), .B(n29959), .Z(n30026) );
  XOR U29435 ( .A(n30032), .B(n30033), .Z(n29959) );
  AND U29436 ( .A(n174), .B(n29994), .Z(n30033) );
  XOR U29437 ( .A(n29992), .B(n30032), .Z(n29994) );
  XOR U29438 ( .A(n30034), .B(n30035), .Z(n30024) );
  AND U29439 ( .A(n30036), .B(n30037), .Z(n30035) );
  XNOR U29440 ( .A(n30034), .B(n29862), .Z(n30037) );
  IV U29441 ( .A(n29865), .Z(n29862) );
  XOR U29442 ( .A(n30038), .B(n30039), .Z(n29865) );
  AND U29443 ( .A(n166), .B(n30040), .Z(n30039) );
  XOR U29444 ( .A(n30041), .B(n30038), .Z(n30040) );
  XOR U29445 ( .A(n29866), .B(n30034), .Z(n30036) );
  XOR U29446 ( .A(n30042), .B(n30043), .Z(n29866) );
  AND U29447 ( .A(n174), .B(n30002), .Z(n30043) );
  XOR U29448 ( .A(n30042), .B(n30000), .Z(n30002) );
  XOR U29449 ( .A(n30044), .B(n30045), .Z(n30034) );
  AND U29450 ( .A(n30046), .B(n30047), .Z(n30045) );
  XNOR U29451 ( .A(n30044), .B(n29890), .Z(n30047) );
  IV U29452 ( .A(n29893), .Z(n29890) );
  XOR U29453 ( .A(n30048), .B(n30049), .Z(n29893) );
  AND U29454 ( .A(n166), .B(n30050), .Z(n30049) );
  XNOR U29455 ( .A(n30051), .B(n30048), .Z(n30050) );
  XOR U29456 ( .A(n29894), .B(n30044), .Z(n30046) );
  XOR U29457 ( .A(n30052), .B(n30053), .Z(n29894) );
  AND U29458 ( .A(n174), .B(n30011), .Z(n30053) );
  XOR U29459 ( .A(n30052), .B(n30009), .Z(n30011) );
  XOR U29460 ( .A(n29968), .B(n30054), .Z(n30044) );
  AND U29461 ( .A(n29970), .B(n30055), .Z(n30054) );
  XNOR U29462 ( .A(n29968), .B(n29939), .Z(n30055) );
  IV U29463 ( .A(n29942), .Z(n29939) );
  XOR U29464 ( .A(n30056), .B(n30057), .Z(n29942) );
  AND U29465 ( .A(n166), .B(n30058), .Z(n30057) );
  XOR U29466 ( .A(n30059), .B(n30056), .Z(n30058) );
  XOR U29467 ( .A(n29943), .B(n29968), .Z(n29970) );
  XOR U29468 ( .A(n30060), .B(n30061), .Z(n29943) );
  AND U29469 ( .A(n174), .B(n30021), .Z(n30061) );
  XOR U29470 ( .A(n30060), .B(n30019), .Z(n30021) );
  AND U29471 ( .A(n30022), .B(n29952), .Z(n29968) );
  XNOR U29472 ( .A(n30062), .B(n30063), .Z(n29952) );
  AND U29473 ( .A(n166), .B(n30064), .Z(n30063) );
  XNOR U29474 ( .A(n30065), .B(n30062), .Z(n30064) );
  XNOR U29475 ( .A(n30066), .B(n30067), .Z(n166) );
  AND U29476 ( .A(n30068), .B(n30069), .Z(n30067) );
  XOR U29477 ( .A(n30031), .B(n30066), .Z(n30069) );
  AND U29478 ( .A(n30070), .B(n30071), .Z(n30031) );
  XNOR U29479 ( .A(n30028), .B(n30066), .Z(n30068) );
  XNOR U29480 ( .A(n30072), .B(n30073), .Z(n30028) );
  AND U29481 ( .A(n170), .B(n30074), .Z(n30073) );
  XNOR U29482 ( .A(n30075), .B(n30076), .Z(n30074) );
  XOR U29483 ( .A(n30077), .B(n30078), .Z(n30066) );
  AND U29484 ( .A(n30079), .B(n30080), .Z(n30078) );
  XNOR U29485 ( .A(n30077), .B(n30070), .Z(n30080) );
  IV U29486 ( .A(n30041), .Z(n30070) );
  XOR U29487 ( .A(n30081), .B(n30082), .Z(n30041) );
  XOR U29488 ( .A(n30083), .B(n30071), .Z(n30082) );
  AND U29489 ( .A(n30051), .B(n30084), .Z(n30071) );
  AND U29490 ( .A(n30085), .B(n30086), .Z(n30083) );
  XOR U29491 ( .A(n30087), .B(n30081), .Z(n30085) );
  XNOR U29492 ( .A(n30038), .B(n30077), .Z(n30079) );
  XNOR U29493 ( .A(n30088), .B(n30089), .Z(n30038) );
  AND U29494 ( .A(n170), .B(n30090), .Z(n30089) );
  XNOR U29495 ( .A(n30091), .B(n30092), .Z(n30090) );
  XOR U29496 ( .A(n30093), .B(n30094), .Z(n30077) );
  AND U29497 ( .A(n30095), .B(n30096), .Z(n30094) );
  XNOR U29498 ( .A(n30093), .B(n30051), .Z(n30096) );
  XOR U29499 ( .A(n30097), .B(n30086), .Z(n30051) );
  XNOR U29500 ( .A(n30098), .B(n30081), .Z(n30086) );
  XOR U29501 ( .A(n30099), .B(n30100), .Z(n30081) );
  AND U29502 ( .A(n30101), .B(n30102), .Z(n30100) );
  XOR U29503 ( .A(n30103), .B(n30099), .Z(n30101) );
  XNOR U29504 ( .A(n30104), .B(n30105), .Z(n30098) );
  AND U29505 ( .A(n30106), .B(n30107), .Z(n30105) );
  XOR U29506 ( .A(n30104), .B(n30108), .Z(n30106) );
  XNOR U29507 ( .A(n30087), .B(n30084), .Z(n30097) );
  AND U29508 ( .A(n30109), .B(n30110), .Z(n30084) );
  XOR U29509 ( .A(n30111), .B(n30112), .Z(n30087) );
  AND U29510 ( .A(n30113), .B(n30114), .Z(n30112) );
  XOR U29511 ( .A(n30111), .B(n30115), .Z(n30113) );
  XNOR U29512 ( .A(n30048), .B(n30093), .Z(n30095) );
  XNOR U29513 ( .A(n30116), .B(n30117), .Z(n30048) );
  AND U29514 ( .A(n170), .B(n30118), .Z(n30117) );
  XNOR U29515 ( .A(n30119), .B(n30120), .Z(n30118) );
  XOR U29516 ( .A(n30121), .B(n30122), .Z(n30093) );
  AND U29517 ( .A(n30123), .B(n30124), .Z(n30122) );
  XNOR U29518 ( .A(n30121), .B(n30109), .Z(n30124) );
  IV U29519 ( .A(n30059), .Z(n30109) );
  XNOR U29520 ( .A(n30125), .B(n30102), .Z(n30059) );
  XNOR U29521 ( .A(n30126), .B(n30108), .Z(n30102) );
  XOR U29522 ( .A(n30127), .B(n30128), .Z(n30108) );
  NOR U29523 ( .A(n30129), .B(n30130), .Z(n30128) );
  XNOR U29524 ( .A(n30127), .B(n30131), .Z(n30129) );
  XNOR U29525 ( .A(n30107), .B(n30099), .Z(n30126) );
  XOR U29526 ( .A(n30132), .B(n30133), .Z(n30099) );
  AND U29527 ( .A(n30134), .B(n30135), .Z(n30133) );
  XNOR U29528 ( .A(n30132), .B(n30136), .Z(n30134) );
  XNOR U29529 ( .A(n30137), .B(n30104), .Z(n30107) );
  XOR U29530 ( .A(n30138), .B(n30139), .Z(n30104) );
  AND U29531 ( .A(n30140), .B(n30141), .Z(n30139) );
  XOR U29532 ( .A(n30138), .B(n30142), .Z(n30140) );
  XNOR U29533 ( .A(n30143), .B(n30144), .Z(n30137) );
  NOR U29534 ( .A(n30145), .B(n30146), .Z(n30144) );
  XOR U29535 ( .A(n30143), .B(n30147), .Z(n30145) );
  XNOR U29536 ( .A(n30103), .B(n30110), .Z(n30125) );
  NOR U29537 ( .A(n30065), .B(n30148), .Z(n30110) );
  XOR U29538 ( .A(n30115), .B(n30114), .Z(n30103) );
  XNOR U29539 ( .A(n30149), .B(n30111), .Z(n30114) );
  XOR U29540 ( .A(n30150), .B(n30151), .Z(n30111) );
  AND U29541 ( .A(n30152), .B(n30153), .Z(n30151) );
  XOR U29542 ( .A(n30150), .B(n30154), .Z(n30152) );
  XNOR U29543 ( .A(n30155), .B(n30156), .Z(n30149) );
  NOR U29544 ( .A(n30157), .B(n30158), .Z(n30156) );
  XNOR U29545 ( .A(n30155), .B(n30159), .Z(n30157) );
  XOR U29546 ( .A(n30160), .B(n30161), .Z(n30115) );
  NOR U29547 ( .A(n30162), .B(n30163), .Z(n30161) );
  XNOR U29548 ( .A(n30160), .B(n30164), .Z(n30162) );
  XNOR U29549 ( .A(n30056), .B(n30121), .Z(n30123) );
  XNOR U29550 ( .A(n30165), .B(n30166), .Z(n30056) );
  AND U29551 ( .A(n170), .B(n30167), .Z(n30166) );
  XNOR U29552 ( .A(n30168), .B(n30169), .Z(n30167) );
  AND U29553 ( .A(n30062), .B(n30065), .Z(n30121) );
  XOR U29554 ( .A(n30170), .B(n30148), .Z(n30065) );
  XNOR U29555 ( .A(p_input[2048]), .B(p_input[80]), .Z(n30148) );
  XOR U29556 ( .A(n30136), .B(n30135), .Z(n30170) );
  XNOR U29557 ( .A(n30171), .B(n30142), .Z(n30135) );
  XNOR U29558 ( .A(n30131), .B(n30130), .Z(n30142) );
  XOR U29559 ( .A(n30172), .B(n30127), .Z(n30130) );
  XNOR U29560 ( .A(n29266), .B(p_input[90]), .Z(n30127) );
  XNOR U29561 ( .A(p_input[2059]), .B(p_input[91]), .Z(n30172) );
  XOR U29562 ( .A(p_input[2060]), .B(p_input[92]), .Z(n30131) );
  XNOR U29563 ( .A(n30141), .B(n30132), .Z(n30171) );
  XNOR U29564 ( .A(n29494), .B(p_input[81]), .Z(n30132) );
  XOR U29565 ( .A(n30173), .B(n30147), .Z(n30141) );
  XNOR U29566 ( .A(p_input[2063]), .B(p_input[95]), .Z(n30147) );
  XOR U29567 ( .A(n30138), .B(n30146), .Z(n30173) );
  XOR U29568 ( .A(n30174), .B(n30143), .Z(n30146) );
  XOR U29569 ( .A(p_input[2061]), .B(p_input[93]), .Z(n30143) );
  XNOR U29570 ( .A(p_input[2062]), .B(p_input[94]), .Z(n30174) );
  XNOR U29571 ( .A(n29036), .B(p_input[89]), .Z(n30138) );
  XNOR U29572 ( .A(n30154), .B(n30153), .Z(n30136) );
  XNOR U29573 ( .A(n30175), .B(n30159), .Z(n30153) );
  XOR U29574 ( .A(p_input[2056]), .B(p_input[88]), .Z(n30159) );
  XOR U29575 ( .A(n30150), .B(n30158), .Z(n30175) );
  XOR U29576 ( .A(n30176), .B(n30155), .Z(n30158) );
  XOR U29577 ( .A(p_input[2054]), .B(p_input[86]), .Z(n30155) );
  XNOR U29578 ( .A(p_input[2055]), .B(p_input[87]), .Z(n30176) );
  XNOR U29579 ( .A(n29039), .B(p_input[82]), .Z(n30150) );
  XNOR U29580 ( .A(n30164), .B(n30163), .Z(n30154) );
  XOR U29581 ( .A(n30177), .B(n30160), .Z(n30163) );
  XOR U29582 ( .A(p_input[2051]), .B(p_input[83]), .Z(n30160) );
  XNOR U29583 ( .A(p_input[2052]), .B(p_input[84]), .Z(n30177) );
  XOR U29584 ( .A(p_input[2053]), .B(p_input[85]), .Z(n30164) );
  XNOR U29585 ( .A(n30178), .B(n30179), .Z(n30062) );
  AND U29586 ( .A(n170), .B(n30180), .Z(n30179) );
  XNOR U29587 ( .A(n30181), .B(n30182), .Z(n170) );
  AND U29588 ( .A(n30183), .B(n30184), .Z(n30182) );
  XOR U29589 ( .A(n30076), .B(n30181), .Z(n30184) );
  XNOR U29590 ( .A(n30185), .B(n30181), .Z(n30183) );
  XOR U29591 ( .A(n30186), .B(n30187), .Z(n30181) );
  AND U29592 ( .A(n30188), .B(n30189), .Z(n30187) );
  XOR U29593 ( .A(n30091), .B(n30186), .Z(n30189) );
  XOR U29594 ( .A(n30186), .B(n30092), .Z(n30188) );
  XOR U29595 ( .A(n30190), .B(n30191), .Z(n30186) );
  AND U29596 ( .A(n30192), .B(n30193), .Z(n30191) );
  XOR U29597 ( .A(n30119), .B(n30190), .Z(n30193) );
  XOR U29598 ( .A(n30190), .B(n30120), .Z(n30192) );
  XOR U29599 ( .A(n30194), .B(n30195), .Z(n30190) );
  AND U29600 ( .A(n30196), .B(n30197), .Z(n30195) );
  XOR U29601 ( .A(n30194), .B(n30168), .Z(n30197) );
  XNOR U29602 ( .A(n30198), .B(n30199), .Z(n30022) );
  AND U29603 ( .A(n174), .B(n30200), .Z(n30199) );
  XNOR U29604 ( .A(n30201), .B(n30202), .Z(n174) );
  AND U29605 ( .A(n30203), .B(n30204), .Z(n30202) );
  XOR U29606 ( .A(n30201), .B(n30032), .Z(n30204) );
  XNOR U29607 ( .A(n30201), .B(n29992), .Z(n30203) );
  XOR U29608 ( .A(n30205), .B(n30206), .Z(n30201) );
  AND U29609 ( .A(n30207), .B(n30208), .Z(n30206) );
  XOR U29610 ( .A(n30205), .B(n30000), .Z(n30207) );
  XOR U29611 ( .A(n30209), .B(n30210), .Z(n29983) );
  AND U29612 ( .A(n178), .B(n30200), .Z(n30210) );
  XNOR U29613 ( .A(n30198), .B(n30209), .Z(n30200) );
  XNOR U29614 ( .A(n30211), .B(n30212), .Z(n178) );
  AND U29615 ( .A(n30213), .B(n30214), .Z(n30212) );
  XNOR U29616 ( .A(n30215), .B(n30211), .Z(n30214) );
  IV U29617 ( .A(n30032), .Z(n30215) );
  XOR U29618 ( .A(n30185), .B(n30216), .Z(n30032) );
  AND U29619 ( .A(n181), .B(n30217), .Z(n30216) );
  XOR U29620 ( .A(n30075), .B(n30072), .Z(n30217) );
  IV U29621 ( .A(n30185), .Z(n30075) );
  XNOR U29622 ( .A(n29992), .B(n30211), .Z(n30213) );
  XOR U29623 ( .A(n30218), .B(n30219), .Z(n29992) );
  AND U29624 ( .A(n197), .B(n30220), .Z(n30219) );
  XOR U29625 ( .A(n30205), .B(n30221), .Z(n30211) );
  AND U29626 ( .A(n30222), .B(n30208), .Z(n30221) );
  XNOR U29627 ( .A(n30042), .B(n30205), .Z(n30208) );
  XOR U29628 ( .A(n30092), .B(n30223), .Z(n30042) );
  AND U29629 ( .A(n181), .B(n30224), .Z(n30223) );
  XOR U29630 ( .A(n30088), .B(n30092), .Z(n30224) );
  XNOR U29631 ( .A(n30225), .B(n30205), .Z(n30222) );
  IV U29632 ( .A(n30000), .Z(n30225) );
  XOR U29633 ( .A(n30226), .B(n30227), .Z(n30000) );
  AND U29634 ( .A(n197), .B(n30228), .Z(n30227) );
  XOR U29635 ( .A(n30229), .B(n30230), .Z(n30205) );
  AND U29636 ( .A(n30231), .B(n30232), .Z(n30230) );
  XNOR U29637 ( .A(n30052), .B(n30229), .Z(n30232) );
  XOR U29638 ( .A(n30120), .B(n30233), .Z(n30052) );
  AND U29639 ( .A(n181), .B(n30234), .Z(n30233) );
  XOR U29640 ( .A(n30116), .B(n30120), .Z(n30234) );
  XOR U29641 ( .A(n30229), .B(n30009), .Z(n30231) );
  XOR U29642 ( .A(n30235), .B(n30236), .Z(n30009) );
  AND U29643 ( .A(n197), .B(n30237), .Z(n30236) );
  XOR U29644 ( .A(n30238), .B(n30239), .Z(n30229) );
  AND U29645 ( .A(n30240), .B(n30241), .Z(n30239) );
  XNOR U29646 ( .A(n30238), .B(n30060), .Z(n30241) );
  XOR U29647 ( .A(n30169), .B(n30242), .Z(n30060) );
  AND U29648 ( .A(n181), .B(n30243), .Z(n30242) );
  XOR U29649 ( .A(n30165), .B(n30169), .Z(n30243) );
  XNOR U29650 ( .A(n30244), .B(n30238), .Z(n30240) );
  IV U29651 ( .A(n30019), .Z(n30244) );
  XOR U29652 ( .A(n30245), .B(n30246), .Z(n30019) );
  AND U29653 ( .A(n197), .B(n30247), .Z(n30246) );
  AND U29654 ( .A(n30209), .B(n30198), .Z(n30238) );
  XNOR U29655 ( .A(n30248), .B(n30249), .Z(n30198) );
  AND U29656 ( .A(n181), .B(n30180), .Z(n30249) );
  XNOR U29657 ( .A(n30178), .B(n30248), .Z(n30180) );
  XNOR U29658 ( .A(n30250), .B(n30251), .Z(n181) );
  AND U29659 ( .A(n30252), .B(n30253), .Z(n30251) );
  XNOR U29660 ( .A(n30250), .B(n30072), .Z(n30253) );
  IV U29661 ( .A(n30076), .Z(n30072) );
  XOR U29662 ( .A(n30254), .B(n30255), .Z(n30076) );
  AND U29663 ( .A(n185), .B(n30256), .Z(n30255) );
  XOR U29664 ( .A(n30257), .B(n30254), .Z(n30256) );
  XNOR U29665 ( .A(n30250), .B(n30185), .Z(n30252) );
  XOR U29666 ( .A(n30258), .B(n30259), .Z(n30185) );
  AND U29667 ( .A(n193), .B(n30220), .Z(n30259) );
  XOR U29668 ( .A(n30218), .B(n30258), .Z(n30220) );
  XOR U29669 ( .A(n30260), .B(n30261), .Z(n30250) );
  AND U29670 ( .A(n30262), .B(n30263), .Z(n30261) );
  XNOR U29671 ( .A(n30260), .B(n30088), .Z(n30263) );
  IV U29672 ( .A(n30091), .Z(n30088) );
  XOR U29673 ( .A(n30264), .B(n30265), .Z(n30091) );
  AND U29674 ( .A(n185), .B(n30266), .Z(n30265) );
  XOR U29675 ( .A(n30267), .B(n30264), .Z(n30266) );
  XOR U29676 ( .A(n30092), .B(n30260), .Z(n30262) );
  XOR U29677 ( .A(n30268), .B(n30269), .Z(n30092) );
  AND U29678 ( .A(n193), .B(n30228), .Z(n30269) );
  XOR U29679 ( .A(n30268), .B(n30226), .Z(n30228) );
  XOR U29680 ( .A(n30270), .B(n30271), .Z(n30260) );
  AND U29681 ( .A(n30272), .B(n30273), .Z(n30271) );
  XNOR U29682 ( .A(n30270), .B(n30116), .Z(n30273) );
  IV U29683 ( .A(n30119), .Z(n30116) );
  XOR U29684 ( .A(n30274), .B(n30275), .Z(n30119) );
  AND U29685 ( .A(n185), .B(n30276), .Z(n30275) );
  XNOR U29686 ( .A(n30277), .B(n30274), .Z(n30276) );
  XOR U29687 ( .A(n30120), .B(n30270), .Z(n30272) );
  XOR U29688 ( .A(n30278), .B(n30279), .Z(n30120) );
  AND U29689 ( .A(n193), .B(n30237), .Z(n30279) );
  XOR U29690 ( .A(n30278), .B(n30235), .Z(n30237) );
  XOR U29691 ( .A(n30194), .B(n30280), .Z(n30270) );
  AND U29692 ( .A(n30196), .B(n30281), .Z(n30280) );
  XNOR U29693 ( .A(n30194), .B(n30165), .Z(n30281) );
  IV U29694 ( .A(n30168), .Z(n30165) );
  XOR U29695 ( .A(n30282), .B(n30283), .Z(n30168) );
  AND U29696 ( .A(n185), .B(n30284), .Z(n30283) );
  XOR U29697 ( .A(n30285), .B(n30282), .Z(n30284) );
  XOR U29698 ( .A(n30169), .B(n30194), .Z(n30196) );
  XOR U29699 ( .A(n30286), .B(n30287), .Z(n30169) );
  AND U29700 ( .A(n193), .B(n30247), .Z(n30287) );
  XOR U29701 ( .A(n30286), .B(n30245), .Z(n30247) );
  AND U29702 ( .A(n30248), .B(n30178), .Z(n30194) );
  XNOR U29703 ( .A(n30288), .B(n30289), .Z(n30178) );
  AND U29704 ( .A(n185), .B(n30290), .Z(n30289) );
  XNOR U29705 ( .A(n30291), .B(n30288), .Z(n30290) );
  XNOR U29706 ( .A(n30292), .B(n30293), .Z(n185) );
  AND U29707 ( .A(n30294), .B(n30295), .Z(n30293) );
  XOR U29708 ( .A(n30257), .B(n30292), .Z(n30295) );
  AND U29709 ( .A(n30296), .B(n30297), .Z(n30257) );
  XNOR U29710 ( .A(n30254), .B(n30292), .Z(n30294) );
  XNOR U29711 ( .A(n30298), .B(n30299), .Z(n30254) );
  AND U29712 ( .A(n189), .B(n30300), .Z(n30299) );
  XNOR U29713 ( .A(n30301), .B(n30302), .Z(n30300) );
  XOR U29714 ( .A(n30303), .B(n30304), .Z(n30292) );
  AND U29715 ( .A(n30305), .B(n30306), .Z(n30304) );
  XNOR U29716 ( .A(n30303), .B(n30296), .Z(n30306) );
  IV U29717 ( .A(n30267), .Z(n30296) );
  XOR U29718 ( .A(n30307), .B(n30308), .Z(n30267) );
  XOR U29719 ( .A(n30309), .B(n30297), .Z(n30308) );
  AND U29720 ( .A(n30277), .B(n30310), .Z(n30297) );
  AND U29721 ( .A(n30311), .B(n30312), .Z(n30309) );
  XOR U29722 ( .A(n30313), .B(n30307), .Z(n30311) );
  XNOR U29723 ( .A(n30264), .B(n30303), .Z(n30305) );
  XNOR U29724 ( .A(n30314), .B(n30315), .Z(n30264) );
  AND U29725 ( .A(n189), .B(n30316), .Z(n30315) );
  XNOR U29726 ( .A(n30317), .B(n30318), .Z(n30316) );
  XOR U29727 ( .A(n30319), .B(n30320), .Z(n30303) );
  AND U29728 ( .A(n30321), .B(n30322), .Z(n30320) );
  XNOR U29729 ( .A(n30319), .B(n30277), .Z(n30322) );
  XOR U29730 ( .A(n30323), .B(n30312), .Z(n30277) );
  XNOR U29731 ( .A(n30324), .B(n30307), .Z(n30312) );
  XOR U29732 ( .A(n30325), .B(n30326), .Z(n30307) );
  AND U29733 ( .A(n30327), .B(n30328), .Z(n30326) );
  XOR U29734 ( .A(n30329), .B(n30325), .Z(n30327) );
  XNOR U29735 ( .A(n30330), .B(n30331), .Z(n30324) );
  AND U29736 ( .A(n30332), .B(n30333), .Z(n30331) );
  XOR U29737 ( .A(n30330), .B(n30334), .Z(n30332) );
  XNOR U29738 ( .A(n30313), .B(n30310), .Z(n30323) );
  AND U29739 ( .A(n30335), .B(n30336), .Z(n30310) );
  XOR U29740 ( .A(n30337), .B(n30338), .Z(n30313) );
  AND U29741 ( .A(n30339), .B(n30340), .Z(n30338) );
  XOR U29742 ( .A(n30337), .B(n30341), .Z(n30339) );
  XNOR U29743 ( .A(n30274), .B(n30319), .Z(n30321) );
  XNOR U29744 ( .A(n30342), .B(n30343), .Z(n30274) );
  AND U29745 ( .A(n189), .B(n30344), .Z(n30343) );
  XNOR U29746 ( .A(n30345), .B(n30346), .Z(n30344) );
  XOR U29747 ( .A(n30347), .B(n30348), .Z(n30319) );
  AND U29748 ( .A(n30349), .B(n30350), .Z(n30348) );
  XNOR U29749 ( .A(n30347), .B(n30335), .Z(n30350) );
  IV U29750 ( .A(n30285), .Z(n30335) );
  XNOR U29751 ( .A(n30351), .B(n30328), .Z(n30285) );
  XNOR U29752 ( .A(n30352), .B(n30334), .Z(n30328) );
  XNOR U29753 ( .A(n30353), .B(n30354), .Z(n30334) );
  NOR U29754 ( .A(n30355), .B(n30356), .Z(n30354) );
  XOR U29755 ( .A(n30353), .B(n30357), .Z(n30355) );
  XNOR U29756 ( .A(n30333), .B(n30325), .Z(n30352) );
  XOR U29757 ( .A(n30358), .B(n30359), .Z(n30325) );
  AND U29758 ( .A(n30360), .B(n30361), .Z(n30359) );
  XOR U29759 ( .A(n30358), .B(n30362), .Z(n30360) );
  XNOR U29760 ( .A(n30363), .B(n30330), .Z(n30333) );
  XOR U29761 ( .A(n30364), .B(n30365), .Z(n30330) );
  AND U29762 ( .A(n30366), .B(n30367), .Z(n30365) );
  XNOR U29763 ( .A(n30368), .B(n30369), .Z(n30366) );
  IV U29764 ( .A(n30364), .Z(n30368) );
  XNOR U29765 ( .A(n30370), .B(n30371), .Z(n30363) );
  NOR U29766 ( .A(n30372), .B(n30373), .Z(n30371) );
  XNOR U29767 ( .A(n30370), .B(n30374), .Z(n30372) );
  XNOR U29768 ( .A(n30329), .B(n30336), .Z(n30351) );
  NOR U29769 ( .A(n30291), .B(n30375), .Z(n30336) );
  XOR U29770 ( .A(n30341), .B(n30340), .Z(n30329) );
  XNOR U29771 ( .A(n30376), .B(n30337), .Z(n30340) );
  XOR U29772 ( .A(n30377), .B(n30378), .Z(n30337) );
  AND U29773 ( .A(n30379), .B(n30380), .Z(n30378) );
  XOR U29774 ( .A(n30377), .B(n30381), .Z(n30379) );
  XNOR U29775 ( .A(n30382), .B(n30383), .Z(n30376) );
  NOR U29776 ( .A(n30384), .B(n30385), .Z(n30383) );
  XNOR U29777 ( .A(n30382), .B(n30386), .Z(n30384) );
  XOR U29778 ( .A(n30387), .B(n30388), .Z(n30341) );
  NOR U29779 ( .A(n30389), .B(n30390), .Z(n30388) );
  XNOR U29780 ( .A(n30387), .B(n30391), .Z(n30389) );
  XNOR U29781 ( .A(n30282), .B(n30347), .Z(n30349) );
  XNOR U29782 ( .A(n30392), .B(n30393), .Z(n30282) );
  AND U29783 ( .A(n189), .B(n30394), .Z(n30393) );
  XNOR U29784 ( .A(n30395), .B(n30396), .Z(n30394) );
  AND U29785 ( .A(n30288), .B(n30291), .Z(n30347) );
  XOR U29786 ( .A(n30397), .B(n30375), .Z(n30291) );
  XNOR U29787 ( .A(p_input[2048]), .B(p_input[96]), .Z(n30375) );
  XNOR U29788 ( .A(n30362), .B(n30361), .Z(n30397) );
  XNOR U29789 ( .A(n30398), .B(n30369), .Z(n30361) );
  XNOR U29790 ( .A(n30357), .B(n30356), .Z(n30369) );
  XNOR U29791 ( .A(n30399), .B(n30353), .Z(n30356) );
  XNOR U29792 ( .A(p_input[106]), .B(p_input[2058]), .Z(n30353) );
  XOR U29793 ( .A(p_input[107]), .B(n29030), .Z(n30399) );
  XOR U29794 ( .A(p_input[108]), .B(p_input[2060]), .Z(n30357) );
  XNOR U29795 ( .A(n30367), .B(n30358), .Z(n30398) );
  XNOR U29796 ( .A(n29494), .B(p_input[97]), .Z(n30358) );
  XNOR U29797 ( .A(n30400), .B(n30374), .Z(n30367) );
  XNOR U29798 ( .A(p_input[111]), .B(n29033), .Z(n30374) );
  XOR U29799 ( .A(n30364), .B(n30373), .Z(n30400) );
  XOR U29800 ( .A(n30401), .B(n30370), .Z(n30373) );
  XOR U29801 ( .A(p_input[109]), .B(p_input[2061]), .Z(n30370) );
  XOR U29802 ( .A(p_input[110]), .B(n29035), .Z(n30401) );
  XOR U29803 ( .A(p_input[105]), .B(p_input[2057]), .Z(n30364) );
  XOR U29804 ( .A(n30381), .B(n30380), .Z(n30362) );
  XNOR U29805 ( .A(n30402), .B(n30386), .Z(n30380) );
  XOR U29806 ( .A(p_input[104]), .B(p_input[2056]), .Z(n30386) );
  XOR U29807 ( .A(n30377), .B(n30385), .Z(n30402) );
  XOR U29808 ( .A(n30403), .B(n30382), .Z(n30385) );
  XOR U29809 ( .A(p_input[102]), .B(p_input[2054]), .Z(n30382) );
  XOR U29810 ( .A(p_input[103]), .B(n30404), .Z(n30403) );
  XNOR U29811 ( .A(n29039), .B(p_input[98]), .Z(n30377) );
  XNOR U29812 ( .A(n30391), .B(n30390), .Z(n30381) );
  XOR U29813 ( .A(n30405), .B(n30387), .Z(n30390) );
  XOR U29814 ( .A(p_input[2051]), .B(p_input[99]), .Z(n30387) );
  XOR U29815 ( .A(p_input[100]), .B(n30406), .Z(n30405) );
  XOR U29816 ( .A(p_input[101]), .B(p_input[2053]), .Z(n30391) );
  XNOR U29817 ( .A(n30407), .B(n30408), .Z(n30288) );
  AND U29818 ( .A(n189), .B(n30409), .Z(n30408) );
  XNOR U29819 ( .A(n30410), .B(n30411), .Z(n189) );
  AND U29820 ( .A(n30412), .B(n30413), .Z(n30411) );
  XOR U29821 ( .A(n30302), .B(n30410), .Z(n30413) );
  XNOR U29822 ( .A(n30414), .B(n30410), .Z(n30412) );
  XOR U29823 ( .A(n30415), .B(n30416), .Z(n30410) );
  AND U29824 ( .A(n30417), .B(n30418), .Z(n30416) );
  XOR U29825 ( .A(n30317), .B(n30415), .Z(n30418) );
  XOR U29826 ( .A(n30415), .B(n30318), .Z(n30417) );
  XOR U29827 ( .A(n30419), .B(n30420), .Z(n30415) );
  AND U29828 ( .A(n30421), .B(n30422), .Z(n30420) );
  XOR U29829 ( .A(n30345), .B(n30419), .Z(n30422) );
  XOR U29830 ( .A(n30419), .B(n30346), .Z(n30421) );
  XOR U29831 ( .A(n30423), .B(n30424), .Z(n30419) );
  AND U29832 ( .A(n30425), .B(n30426), .Z(n30424) );
  XOR U29833 ( .A(n30423), .B(n30395), .Z(n30426) );
  XNOR U29834 ( .A(n30427), .B(n30428), .Z(n30248) );
  AND U29835 ( .A(n193), .B(n30429), .Z(n30428) );
  XNOR U29836 ( .A(n30430), .B(n30431), .Z(n193) );
  AND U29837 ( .A(n30432), .B(n30433), .Z(n30431) );
  XOR U29838 ( .A(n30430), .B(n30258), .Z(n30433) );
  XNOR U29839 ( .A(n30430), .B(n30218), .Z(n30432) );
  XOR U29840 ( .A(n30434), .B(n30435), .Z(n30430) );
  AND U29841 ( .A(n30436), .B(n30437), .Z(n30435) );
  XOR U29842 ( .A(n30434), .B(n30226), .Z(n30436) );
  XOR U29843 ( .A(n30438), .B(n30439), .Z(n30209) );
  AND U29844 ( .A(n197), .B(n30429), .Z(n30439) );
  XNOR U29845 ( .A(n30427), .B(n30438), .Z(n30429) );
  XNOR U29846 ( .A(n30440), .B(n30441), .Z(n197) );
  AND U29847 ( .A(n30442), .B(n30443), .Z(n30441) );
  XNOR U29848 ( .A(n30444), .B(n30440), .Z(n30443) );
  IV U29849 ( .A(n30258), .Z(n30444) );
  XOR U29850 ( .A(n30414), .B(n30445), .Z(n30258) );
  AND U29851 ( .A(n200), .B(n30446), .Z(n30445) );
  XOR U29852 ( .A(n30301), .B(n30298), .Z(n30446) );
  IV U29853 ( .A(n30414), .Z(n30301) );
  XNOR U29854 ( .A(n30218), .B(n30440), .Z(n30442) );
  XOR U29855 ( .A(n30447), .B(n30448), .Z(n30218) );
  AND U29856 ( .A(n216), .B(n30449), .Z(n30448) );
  XOR U29857 ( .A(n30434), .B(n30450), .Z(n30440) );
  AND U29858 ( .A(n30451), .B(n30437), .Z(n30450) );
  XNOR U29859 ( .A(n30268), .B(n30434), .Z(n30437) );
  XOR U29860 ( .A(n30318), .B(n30452), .Z(n30268) );
  AND U29861 ( .A(n200), .B(n30453), .Z(n30452) );
  XOR U29862 ( .A(n30314), .B(n30318), .Z(n30453) );
  XNOR U29863 ( .A(n30454), .B(n30434), .Z(n30451) );
  IV U29864 ( .A(n30226), .Z(n30454) );
  XOR U29865 ( .A(n30455), .B(n30456), .Z(n30226) );
  AND U29866 ( .A(n216), .B(n30457), .Z(n30456) );
  XOR U29867 ( .A(n30458), .B(n30459), .Z(n30434) );
  AND U29868 ( .A(n30460), .B(n30461), .Z(n30459) );
  XNOR U29869 ( .A(n30278), .B(n30458), .Z(n30461) );
  XOR U29870 ( .A(n30346), .B(n30462), .Z(n30278) );
  AND U29871 ( .A(n200), .B(n30463), .Z(n30462) );
  XOR U29872 ( .A(n30342), .B(n30346), .Z(n30463) );
  XOR U29873 ( .A(n30458), .B(n30235), .Z(n30460) );
  XOR U29874 ( .A(n30464), .B(n30465), .Z(n30235) );
  AND U29875 ( .A(n216), .B(n30466), .Z(n30465) );
  XOR U29876 ( .A(n30467), .B(n30468), .Z(n30458) );
  AND U29877 ( .A(n30469), .B(n30470), .Z(n30468) );
  XNOR U29878 ( .A(n30467), .B(n30286), .Z(n30470) );
  XOR U29879 ( .A(n30396), .B(n30471), .Z(n30286) );
  AND U29880 ( .A(n200), .B(n30472), .Z(n30471) );
  XOR U29881 ( .A(n30392), .B(n30396), .Z(n30472) );
  XNOR U29882 ( .A(n30473), .B(n30467), .Z(n30469) );
  IV U29883 ( .A(n30245), .Z(n30473) );
  XOR U29884 ( .A(n30474), .B(n30475), .Z(n30245) );
  AND U29885 ( .A(n216), .B(n30476), .Z(n30475) );
  AND U29886 ( .A(n30438), .B(n30427), .Z(n30467) );
  XNOR U29887 ( .A(n30477), .B(n30478), .Z(n30427) );
  AND U29888 ( .A(n200), .B(n30409), .Z(n30478) );
  XNOR U29889 ( .A(n30407), .B(n30477), .Z(n30409) );
  XNOR U29890 ( .A(n30479), .B(n30480), .Z(n200) );
  AND U29891 ( .A(n30481), .B(n30482), .Z(n30480) );
  XNOR U29892 ( .A(n30479), .B(n30298), .Z(n30482) );
  IV U29893 ( .A(n30302), .Z(n30298) );
  XOR U29894 ( .A(n30483), .B(n30484), .Z(n30302) );
  AND U29895 ( .A(n204), .B(n30485), .Z(n30484) );
  XOR U29896 ( .A(n30486), .B(n30483), .Z(n30485) );
  XNOR U29897 ( .A(n30479), .B(n30414), .Z(n30481) );
  XOR U29898 ( .A(n30487), .B(n30488), .Z(n30414) );
  AND U29899 ( .A(n212), .B(n30449), .Z(n30488) );
  XOR U29900 ( .A(n30447), .B(n30487), .Z(n30449) );
  XOR U29901 ( .A(n30489), .B(n30490), .Z(n30479) );
  AND U29902 ( .A(n30491), .B(n30492), .Z(n30490) );
  XNOR U29903 ( .A(n30489), .B(n30314), .Z(n30492) );
  IV U29904 ( .A(n30317), .Z(n30314) );
  XOR U29905 ( .A(n30493), .B(n30494), .Z(n30317) );
  AND U29906 ( .A(n204), .B(n30495), .Z(n30494) );
  XOR U29907 ( .A(n30496), .B(n30493), .Z(n30495) );
  XOR U29908 ( .A(n30318), .B(n30489), .Z(n30491) );
  XOR U29909 ( .A(n30497), .B(n30498), .Z(n30318) );
  AND U29910 ( .A(n212), .B(n30457), .Z(n30498) );
  XOR U29911 ( .A(n30497), .B(n30455), .Z(n30457) );
  XOR U29912 ( .A(n30499), .B(n30500), .Z(n30489) );
  AND U29913 ( .A(n30501), .B(n30502), .Z(n30500) );
  XNOR U29914 ( .A(n30499), .B(n30342), .Z(n30502) );
  IV U29915 ( .A(n30345), .Z(n30342) );
  XOR U29916 ( .A(n30503), .B(n30504), .Z(n30345) );
  AND U29917 ( .A(n204), .B(n30505), .Z(n30504) );
  XNOR U29918 ( .A(n30506), .B(n30503), .Z(n30505) );
  XOR U29919 ( .A(n30346), .B(n30499), .Z(n30501) );
  XOR U29920 ( .A(n30507), .B(n30508), .Z(n30346) );
  AND U29921 ( .A(n212), .B(n30466), .Z(n30508) );
  XOR U29922 ( .A(n30507), .B(n30464), .Z(n30466) );
  XOR U29923 ( .A(n30423), .B(n30509), .Z(n30499) );
  AND U29924 ( .A(n30425), .B(n30510), .Z(n30509) );
  XNOR U29925 ( .A(n30423), .B(n30392), .Z(n30510) );
  IV U29926 ( .A(n30395), .Z(n30392) );
  XOR U29927 ( .A(n30511), .B(n30512), .Z(n30395) );
  AND U29928 ( .A(n204), .B(n30513), .Z(n30512) );
  XOR U29929 ( .A(n30514), .B(n30511), .Z(n30513) );
  XOR U29930 ( .A(n30396), .B(n30423), .Z(n30425) );
  XOR U29931 ( .A(n30515), .B(n30516), .Z(n30396) );
  AND U29932 ( .A(n212), .B(n30476), .Z(n30516) );
  XOR U29933 ( .A(n30515), .B(n30474), .Z(n30476) );
  AND U29934 ( .A(n30477), .B(n30407), .Z(n30423) );
  XNOR U29935 ( .A(n30517), .B(n30518), .Z(n30407) );
  AND U29936 ( .A(n204), .B(n30519), .Z(n30518) );
  XNOR U29937 ( .A(n30520), .B(n30517), .Z(n30519) );
  XNOR U29938 ( .A(n30521), .B(n30522), .Z(n204) );
  AND U29939 ( .A(n30523), .B(n30524), .Z(n30522) );
  XOR U29940 ( .A(n30486), .B(n30521), .Z(n30524) );
  AND U29941 ( .A(n30525), .B(n30526), .Z(n30486) );
  XNOR U29942 ( .A(n30483), .B(n30521), .Z(n30523) );
  XNOR U29943 ( .A(n30527), .B(n30528), .Z(n30483) );
  AND U29944 ( .A(n208), .B(n30529), .Z(n30528) );
  XNOR U29945 ( .A(n30530), .B(n30531), .Z(n30529) );
  XOR U29946 ( .A(n30532), .B(n30533), .Z(n30521) );
  AND U29947 ( .A(n30534), .B(n30535), .Z(n30533) );
  XNOR U29948 ( .A(n30532), .B(n30525), .Z(n30535) );
  IV U29949 ( .A(n30496), .Z(n30525) );
  XOR U29950 ( .A(n30536), .B(n30537), .Z(n30496) );
  XOR U29951 ( .A(n30538), .B(n30526), .Z(n30537) );
  AND U29952 ( .A(n30506), .B(n30539), .Z(n30526) );
  AND U29953 ( .A(n30540), .B(n30541), .Z(n30538) );
  XOR U29954 ( .A(n30542), .B(n30536), .Z(n30540) );
  XNOR U29955 ( .A(n30493), .B(n30532), .Z(n30534) );
  XNOR U29956 ( .A(n30543), .B(n30544), .Z(n30493) );
  AND U29957 ( .A(n208), .B(n30545), .Z(n30544) );
  XNOR U29958 ( .A(n30546), .B(n30547), .Z(n30545) );
  XOR U29959 ( .A(n30548), .B(n30549), .Z(n30532) );
  AND U29960 ( .A(n30550), .B(n30551), .Z(n30549) );
  XNOR U29961 ( .A(n30548), .B(n30506), .Z(n30551) );
  XOR U29962 ( .A(n30552), .B(n30541), .Z(n30506) );
  XNOR U29963 ( .A(n30553), .B(n30536), .Z(n30541) );
  XOR U29964 ( .A(n30554), .B(n30555), .Z(n30536) );
  AND U29965 ( .A(n30556), .B(n30557), .Z(n30555) );
  XOR U29966 ( .A(n30558), .B(n30554), .Z(n30556) );
  XNOR U29967 ( .A(n30559), .B(n30560), .Z(n30553) );
  AND U29968 ( .A(n30561), .B(n30562), .Z(n30560) );
  XOR U29969 ( .A(n30559), .B(n30563), .Z(n30561) );
  XNOR U29970 ( .A(n30542), .B(n30539), .Z(n30552) );
  AND U29971 ( .A(n30564), .B(n30565), .Z(n30539) );
  XOR U29972 ( .A(n30566), .B(n30567), .Z(n30542) );
  AND U29973 ( .A(n30568), .B(n30569), .Z(n30567) );
  XOR U29974 ( .A(n30566), .B(n30570), .Z(n30568) );
  XNOR U29975 ( .A(n30503), .B(n30548), .Z(n30550) );
  XNOR U29976 ( .A(n30571), .B(n30572), .Z(n30503) );
  AND U29977 ( .A(n208), .B(n30573), .Z(n30572) );
  XNOR U29978 ( .A(n30574), .B(n30575), .Z(n30573) );
  XOR U29979 ( .A(n30576), .B(n30577), .Z(n30548) );
  AND U29980 ( .A(n30578), .B(n30579), .Z(n30577) );
  XNOR U29981 ( .A(n30576), .B(n30564), .Z(n30579) );
  IV U29982 ( .A(n30514), .Z(n30564) );
  XNOR U29983 ( .A(n30580), .B(n30557), .Z(n30514) );
  XNOR U29984 ( .A(n30581), .B(n30563), .Z(n30557) );
  XNOR U29985 ( .A(n30582), .B(n30583), .Z(n30563) );
  NOR U29986 ( .A(n30584), .B(n30585), .Z(n30583) );
  XOR U29987 ( .A(n30582), .B(n30586), .Z(n30584) );
  XNOR U29988 ( .A(n30562), .B(n30554), .Z(n30581) );
  XOR U29989 ( .A(n30587), .B(n30588), .Z(n30554) );
  AND U29990 ( .A(n30589), .B(n30590), .Z(n30588) );
  XOR U29991 ( .A(n30587), .B(n30591), .Z(n30589) );
  XNOR U29992 ( .A(n30592), .B(n30559), .Z(n30562) );
  XOR U29993 ( .A(n30593), .B(n30594), .Z(n30559) );
  AND U29994 ( .A(n30595), .B(n30596), .Z(n30594) );
  XNOR U29995 ( .A(n30597), .B(n30598), .Z(n30595) );
  IV U29996 ( .A(n30593), .Z(n30597) );
  XNOR U29997 ( .A(n30599), .B(n30600), .Z(n30592) );
  NOR U29998 ( .A(n30601), .B(n30602), .Z(n30600) );
  XNOR U29999 ( .A(n30599), .B(n30603), .Z(n30601) );
  XNOR U30000 ( .A(n30558), .B(n30565), .Z(n30580) );
  NOR U30001 ( .A(n30520), .B(n30604), .Z(n30565) );
  XOR U30002 ( .A(n30570), .B(n30569), .Z(n30558) );
  XNOR U30003 ( .A(n30605), .B(n30566), .Z(n30569) );
  XOR U30004 ( .A(n30606), .B(n30607), .Z(n30566) );
  AND U30005 ( .A(n30608), .B(n30609), .Z(n30607) );
  XNOR U30006 ( .A(n30610), .B(n30611), .Z(n30608) );
  IV U30007 ( .A(n30606), .Z(n30610) );
  XNOR U30008 ( .A(n30612), .B(n30613), .Z(n30605) );
  NOR U30009 ( .A(n30614), .B(n30615), .Z(n30613) );
  XNOR U30010 ( .A(n30612), .B(n30616), .Z(n30614) );
  XOR U30011 ( .A(n30617), .B(n30618), .Z(n30570) );
  NOR U30012 ( .A(n30619), .B(n30620), .Z(n30618) );
  XNOR U30013 ( .A(n30617), .B(n30621), .Z(n30619) );
  XNOR U30014 ( .A(n30511), .B(n30576), .Z(n30578) );
  XNOR U30015 ( .A(n30622), .B(n30623), .Z(n30511) );
  AND U30016 ( .A(n208), .B(n30624), .Z(n30623) );
  XNOR U30017 ( .A(n30625), .B(n30626), .Z(n30624) );
  AND U30018 ( .A(n30517), .B(n30520), .Z(n30576) );
  XOR U30019 ( .A(n30627), .B(n30604), .Z(n30520) );
  XNOR U30020 ( .A(p_input[112]), .B(p_input[2048]), .Z(n30604) );
  XNOR U30021 ( .A(n30591), .B(n30590), .Z(n30627) );
  XNOR U30022 ( .A(n30628), .B(n30598), .Z(n30590) );
  XNOR U30023 ( .A(n30586), .B(n30585), .Z(n30598) );
  XNOR U30024 ( .A(n30629), .B(n30582), .Z(n30585) );
  XNOR U30025 ( .A(p_input[122]), .B(p_input[2058]), .Z(n30582) );
  XOR U30026 ( .A(p_input[123]), .B(n29030), .Z(n30629) );
  XOR U30027 ( .A(p_input[124]), .B(p_input[2060]), .Z(n30586) );
  XOR U30028 ( .A(n30596), .B(n30630), .Z(n30628) );
  IV U30029 ( .A(n30587), .Z(n30630) );
  XOR U30030 ( .A(p_input[113]), .B(p_input[2049]), .Z(n30587) );
  XNOR U30031 ( .A(n30631), .B(n30603), .Z(n30596) );
  XNOR U30032 ( .A(p_input[127]), .B(n29033), .Z(n30603) );
  XOR U30033 ( .A(n30593), .B(n30602), .Z(n30631) );
  XOR U30034 ( .A(n30632), .B(n30599), .Z(n30602) );
  XOR U30035 ( .A(p_input[125]), .B(p_input[2061]), .Z(n30599) );
  XOR U30036 ( .A(p_input[126]), .B(n29035), .Z(n30632) );
  XOR U30037 ( .A(p_input[121]), .B(p_input[2057]), .Z(n30593) );
  XOR U30038 ( .A(n30611), .B(n30609), .Z(n30591) );
  XNOR U30039 ( .A(n30633), .B(n30616), .Z(n30609) );
  XOR U30040 ( .A(p_input[120]), .B(p_input[2056]), .Z(n30616) );
  XOR U30041 ( .A(n30606), .B(n30615), .Z(n30633) );
  XOR U30042 ( .A(n30634), .B(n30612), .Z(n30615) );
  XOR U30043 ( .A(p_input[118]), .B(p_input[2054]), .Z(n30612) );
  XOR U30044 ( .A(p_input[119]), .B(n30404), .Z(n30634) );
  XOR U30045 ( .A(p_input[114]), .B(p_input[2050]), .Z(n30606) );
  XNOR U30046 ( .A(n30621), .B(n30620), .Z(n30611) );
  XOR U30047 ( .A(n30635), .B(n30617), .Z(n30620) );
  XOR U30048 ( .A(p_input[115]), .B(p_input[2051]), .Z(n30617) );
  XOR U30049 ( .A(p_input[116]), .B(n30406), .Z(n30635) );
  XOR U30050 ( .A(p_input[117]), .B(p_input[2053]), .Z(n30621) );
  XNOR U30051 ( .A(n30636), .B(n30637), .Z(n30517) );
  AND U30052 ( .A(n208), .B(n30638), .Z(n30637) );
  XNOR U30053 ( .A(n30639), .B(n30640), .Z(n208) );
  AND U30054 ( .A(n30641), .B(n30642), .Z(n30640) );
  XOR U30055 ( .A(n30531), .B(n30639), .Z(n30642) );
  XNOR U30056 ( .A(n30643), .B(n30639), .Z(n30641) );
  XOR U30057 ( .A(n30644), .B(n30645), .Z(n30639) );
  AND U30058 ( .A(n30646), .B(n30647), .Z(n30645) );
  XOR U30059 ( .A(n30546), .B(n30644), .Z(n30647) );
  XOR U30060 ( .A(n30644), .B(n30547), .Z(n30646) );
  XOR U30061 ( .A(n30648), .B(n30649), .Z(n30644) );
  AND U30062 ( .A(n30650), .B(n30651), .Z(n30649) );
  XOR U30063 ( .A(n30574), .B(n30648), .Z(n30651) );
  XOR U30064 ( .A(n30648), .B(n30575), .Z(n30650) );
  XOR U30065 ( .A(n30652), .B(n30653), .Z(n30648) );
  AND U30066 ( .A(n30654), .B(n30655), .Z(n30653) );
  XOR U30067 ( .A(n30652), .B(n30625), .Z(n30655) );
  XNOR U30068 ( .A(n30656), .B(n30657), .Z(n30477) );
  AND U30069 ( .A(n212), .B(n30658), .Z(n30657) );
  XNOR U30070 ( .A(n30659), .B(n30660), .Z(n212) );
  AND U30071 ( .A(n30661), .B(n30662), .Z(n30660) );
  XOR U30072 ( .A(n30659), .B(n30487), .Z(n30662) );
  XNOR U30073 ( .A(n30659), .B(n30447), .Z(n30661) );
  XOR U30074 ( .A(n30663), .B(n30664), .Z(n30659) );
  AND U30075 ( .A(n30665), .B(n30666), .Z(n30664) );
  XOR U30076 ( .A(n30663), .B(n30455), .Z(n30665) );
  XOR U30077 ( .A(n30667), .B(n30668), .Z(n30438) );
  AND U30078 ( .A(n216), .B(n30658), .Z(n30668) );
  XNOR U30079 ( .A(n30656), .B(n30667), .Z(n30658) );
  XNOR U30080 ( .A(n30669), .B(n30670), .Z(n216) );
  AND U30081 ( .A(n30671), .B(n30672), .Z(n30670) );
  XNOR U30082 ( .A(n30673), .B(n30669), .Z(n30672) );
  IV U30083 ( .A(n30487), .Z(n30673) );
  XOR U30084 ( .A(n30643), .B(n30674), .Z(n30487) );
  AND U30085 ( .A(n219), .B(n30675), .Z(n30674) );
  XOR U30086 ( .A(n30530), .B(n30527), .Z(n30675) );
  IV U30087 ( .A(n30643), .Z(n30530) );
  XNOR U30088 ( .A(n30447), .B(n30669), .Z(n30671) );
  XOR U30089 ( .A(n30676), .B(n30677), .Z(n30447) );
  AND U30090 ( .A(n235), .B(n30678), .Z(n30677) );
  XOR U30091 ( .A(n30663), .B(n30679), .Z(n30669) );
  AND U30092 ( .A(n30680), .B(n30666), .Z(n30679) );
  XNOR U30093 ( .A(n30497), .B(n30663), .Z(n30666) );
  XOR U30094 ( .A(n30547), .B(n30681), .Z(n30497) );
  AND U30095 ( .A(n219), .B(n30682), .Z(n30681) );
  XOR U30096 ( .A(n30543), .B(n30547), .Z(n30682) );
  XNOR U30097 ( .A(n30683), .B(n30663), .Z(n30680) );
  IV U30098 ( .A(n30455), .Z(n30683) );
  XOR U30099 ( .A(n30684), .B(n30685), .Z(n30455) );
  AND U30100 ( .A(n235), .B(n30686), .Z(n30685) );
  XOR U30101 ( .A(n30687), .B(n30688), .Z(n30663) );
  AND U30102 ( .A(n30689), .B(n30690), .Z(n30688) );
  XNOR U30103 ( .A(n30507), .B(n30687), .Z(n30690) );
  XOR U30104 ( .A(n30575), .B(n30691), .Z(n30507) );
  AND U30105 ( .A(n219), .B(n30692), .Z(n30691) );
  XOR U30106 ( .A(n30571), .B(n30575), .Z(n30692) );
  XOR U30107 ( .A(n30687), .B(n30464), .Z(n30689) );
  XOR U30108 ( .A(n30693), .B(n30694), .Z(n30464) );
  AND U30109 ( .A(n235), .B(n30695), .Z(n30694) );
  XOR U30110 ( .A(n30696), .B(n30697), .Z(n30687) );
  AND U30111 ( .A(n30698), .B(n30699), .Z(n30697) );
  XNOR U30112 ( .A(n30696), .B(n30515), .Z(n30699) );
  XOR U30113 ( .A(n30626), .B(n30700), .Z(n30515) );
  AND U30114 ( .A(n219), .B(n30701), .Z(n30700) );
  XOR U30115 ( .A(n30622), .B(n30626), .Z(n30701) );
  XNOR U30116 ( .A(n30702), .B(n30696), .Z(n30698) );
  IV U30117 ( .A(n30474), .Z(n30702) );
  XOR U30118 ( .A(n30703), .B(n30704), .Z(n30474) );
  AND U30119 ( .A(n235), .B(n30705), .Z(n30704) );
  AND U30120 ( .A(n30667), .B(n30656), .Z(n30696) );
  XNOR U30121 ( .A(n30706), .B(n30707), .Z(n30656) );
  AND U30122 ( .A(n219), .B(n30638), .Z(n30707) );
  XNOR U30123 ( .A(n30636), .B(n30706), .Z(n30638) );
  XNOR U30124 ( .A(n30708), .B(n30709), .Z(n219) );
  AND U30125 ( .A(n30710), .B(n30711), .Z(n30709) );
  XNOR U30126 ( .A(n30708), .B(n30527), .Z(n30711) );
  IV U30127 ( .A(n30531), .Z(n30527) );
  XOR U30128 ( .A(n30712), .B(n30713), .Z(n30531) );
  AND U30129 ( .A(n223), .B(n30714), .Z(n30713) );
  XOR U30130 ( .A(n30715), .B(n30712), .Z(n30714) );
  XNOR U30131 ( .A(n30708), .B(n30643), .Z(n30710) );
  XOR U30132 ( .A(n30716), .B(n30717), .Z(n30643) );
  AND U30133 ( .A(n231), .B(n30678), .Z(n30717) );
  XOR U30134 ( .A(n30676), .B(n30716), .Z(n30678) );
  XOR U30135 ( .A(n30718), .B(n30719), .Z(n30708) );
  AND U30136 ( .A(n30720), .B(n30721), .Z(n30719) );
  XNOR U30137 ( .A(n30718), .B(n30543), .Z(n30721) );
  IV U30138 ( .A(n30546), .Z(n30543) );
  XOR U30139 ( .A(n30722), .B(n30723), .Z(n30546) );
  AND U30140 ( .A(n223), .B(n30724), .Z(n30723) );
  XOR U30141 ( .A(n30725), .B(n30722), .Z(n30724) );
  XOR U30142 ( .A(n30547), .B(n30718), .Z(n30720) );
  XOR U30143 ( .A(n30726), .B(n30727), .Z(n30547) );
  AND U30144 ( .A(n231), .B(n30686), .Z(n30727) );
  XOR U30145 ( .A(n30726), .B(n30684), .Z(n30686) );
  XOR U30146 ( .A(n30728), .B(n30729), .Z(n30718) );
  AND U30147 ( .A(n30730), .B(n30731), .Z(n30729) );
  XNOR U30148 ( .A(n30728), .B(n30571), .Z(n30731) );
  IV U30149 ( .A(n30574), .Z(n30571) );
  XOR U30150 ( .A(n30732), .B(n30733), .Z(n30574) );
  AND U30151 ( .A(n223), .B(n30734), .Z(n30733) );
  XNOR U30152 ( .A(n30735), .B(n30732), .Z(n30734) );
  XOR U30153 ( .A(n30575), .B(n30728), .Z(n30730) );
  XOR U30154 ( .A(n30736), .B(n30737), .Z(n30575) );
  AND U30155 ( .A(n231), .B(n30695), .Z(n30737) );
  XOR U30156 ( .A(n30736), .B(n30693), .Z(n30695) );
  XOR U30157 ( .A(n30652), .B(n30738), .Z(n30728) );
  AND U30158 ( .A(n30654), .B(n30739), .Z(n30738) );
  XNOR U30159 ( .A(n30652), .B(n30622), .Z(n30739) );
  IV U30160 ( .A(n30625), .Z(n30622) );
  XOR U30161 ( .A(n30740), .B(n30741), .Z(n30625) );
  AND U30162 ( .A(n223), .B(n30742), .Z(n30741) );
  XOR U30163 ( .A(n30743), .B(n30740), .Z(n30742) );
  XOR U30164 ( .A(n30626), .B(n30652), .Z(n30654) );
  XOR U30165 ( .A(n30744), .B(n30745), .Z(n30626) );
  AND U30166 ( .A(n231), .B(n30705), .Z(n30745) );
  XOR U30167 ( .A(n30744), .B(n30703), .Z(n30705) );
  AND U30168 ( .A(n30706), .B(n30636), .Z(n30652) );
  XNOR U30169 ( .A(n30746), .B(n30747), .Z(n30636) );
  AND U30170 ( .A(n223), .B(n30748), .Z(n30747) );
  XNOR U30171 ( .A(n30749), .B(n30746), .Z(n30748) );
  XNOR U30172 ( .A(n30750), .B(n30751), .Z(n223) );
  AND U30173 ( .A(n30752), .B(n30753), .Z(n30751) );
  XOR U30174 ( .A(n30715), .B(n30750), .Z(n30753) );
  AND U30175 ( .A(n30754), .B(n30755), .Z(n30715) );
  XNOR U30176 ( .A(n30712), .B(n30750), .Z(n30752) );
  XNOR U30177 ( .A(n30756), .B(n30757), .Z(n30712) );
  AND U30178 ( .A(n227), .B(n30758), .Z(n30757) );
  XNOR U30179 ( .A(n30759), .B(n30760), .Z(n30758) );
  XOR U30180 ( .A(n30761), .B(n30762), .Z(n30750) );
  AND U30181 ( .A(n30763), .B(n30764), .Z(n30762) );
  XNOR U30182 ( .A(n30761), .B(n30754), .Z(n30764) );
  IV U30183 ( .A(n30725), .Z(n30754) );
  XOR U30184 ( .A(n30765), .B(n30766), .Z(n30725) );
  XOR U30185 ( .A(n30767), .B(n30755), .Z(n30766) );
  AND U30186 ( .A(n30735), .B(n30768), .Z(n30755) );
  AND U30187 ( .A(n30769), .B(n30770), .Z(n30767) );
  XOR U30188 ( .A(n30771), .B(n30765), .Z(n30769) );
  XNOR U30189 ( .A(n30722), .B(n30761), .Z(n30763) );
  XNOR U30190 ( .A(n30772), .B(n30773), .Z(n30722) );
  AND U30191 ( .A(n227), .B(n30774), .Z(n30773) );
  XNOR U30192 ( .A(n30775), .B(n30776), .Z(n30774) );
  XOR U30193 ( .A(n30777), .B(n30778), .Z(n30761) );
  AND U30194 ( .A(n30779), .B(n30780), .Z(n30778) );
  XNOR U30195 ( .A(n30777), .B(n30735), .Z(n30780) );
  XOR U30196 ( .A(n30781), .B(n30770), .Z(n30735) );
  XNOR U30197 ( .A(n30782), .B(n30765), .Z(n30770) );
  XOR U30198 ( .A(n30783), .B(n30784), .Z(n30765) );
  AND U30199 ( .A(n30785), .B(n30786), .Z(n30784) );
  XOR U30200 ( .A(n30787), .B(n30783), .Z(n30785) );
  XNOR U30201 ( .A(n30788), .B(n30789), .Z(n30782) );
  AND U30202 ( .A(n30790), .B(n30791), .Z(n30789) );
  XOR U30203 ( .A(n30788), .B(n30792), .Z(n30790) );
  XNOR U30204 ( .A(n30771), .B(n30768), .Z(n30781) );
  AND U30205 ( .A(n30793), .B(n30794), .Z(n30768) );
  XOR U30206 ( .A(n30795), .B(n30796), .Z(n30771) );
  AND U30207 ( .A(n30797), .B(n30798), .Z(n30796) );
  XOR U30208 ( .A(n30795), .B(n30799), .Z(n30797) );
  XNOR U30209 ( .A(n30732), .B(n30777), .Z(n30779) );
  XNOR U30210 ( .A(n30800), .B(n30801), .Z(n30732) );
  AND U30211 ( .A(n227), .B(n30802), .Z(n30801) );
  XNOR U30212 ( .A(n30803), .B(n30804), .Z(n30802) );
  XOR U30213 ( .A(n30805), .B(n30806), .Z(n30777) );
  AND U30214 ( .A(n30807), .B(n30808), .Z(n30806) );
  XNOR U30215 ( .A(n30805), .B(n30793), .Z(n30808) );
  IV U30216 ( .A(n30743), .Z(n30793) );
  XNOR U30217 ( .A(n30809), .B(n30786), .Z(n30743) );
  XNOR U30218 ( .A(n30810), .B(n30792), .Z(n30786) );
  XNOR U30219 ( .A(n30811), .B(n30812), .Z(n30792) );
  NOR U30220 ( .A(n30813), .B(n30814), .Z(n30812) );
  XOR U30221 ( .A(n30811), .B(n30815), .Z(n30813) );
  XNOR U30222 ( .A(n30791), .B(n30783), .Z(n30810) );
  XOR U30223 ( .A(n30816), .B(n30817), .Z(n30783) );
  AND U30224 ( .A(n30818), .B(n30819), .Z(n30817) );
  XOR U30225 ( .A(n30816), .B(n30820), .Z(n30818) );
  XNOR U30226 ( .A(n30821), .B(n30788), .Z(n30791) );
  XOR U30227 ( .A(n30822), .B(n30823), .Z(n30788) );
  AND U30228 ( .A(n30824), .B(n30825), .Z(n30823) );
  XNOR U30229 ( .A(n30826), .B(n30827), .Z(n30824) );
  IV U30230 ( .A(n30822), .Z(n30826) );
  XNOR U30231 ( .A(n30828), .B(n30829), .Z(n30821) );
  NOR U30232 ( .A(n30830), .B(n30831), .Z(n30829) );
  XNOR U30233 ( .A(n30828), .B(n30832), .Z(n30830) );
  XNOR U30234 ( .A(n30787), .B(n30794), .Z(n30809) );
  NOR U30235 ( .A(n30749), .B(n30833), .Z(n30794) );
  XOR U30236 ( .A(n30799), .B(n30798), .Z(n30787) );
  XNOR U30237 ( .A(n30834), .B(n30795), .Z(n30798) );
  XOR U30238 ( .A(n30835), .B(n30836), .Z(n30795) );
  AND U30239 ( .A(n30837), .B(n30838), .Z(n30836) );
  XNOR U30240 ( .A(n30839), .B(n30840), .Z(n30837) );
  IV U30241 ( .A(n30835), .Z(n30839) );
  XNOR U30242 ( .A(n30841), .B(n30842), .Z(n30834) );
  NOR U30243 ( .A(n30843), .B(n30844), .Z(n30842) );
  XNOR U30244 ( .A(n30841), .B(n30845), .Z(n30843) );
  XOR U30245 ( .A(n30846), .B(n30847), .Z(n30799) );
  NOR U30246 ( .A(n30848), .B(n30849), .Z(n30847) );
  XNOR U30247 ( .A(n30846), .B(n30850), .Z(n30848) );
  XNOR U30248 ( .A(n30740), .B(n30805), .Z(n30807) );
  XNOR U30249 ( .A(n30851), .B(n30852), .Z(n30740) );
  AND U30250 ( .A(n227), .B(n30853), .Z(n30852) );
  XNOR U30251 ( .A(n30854), .B(n30855), .Z(n30853) );
  AND U30252 ( .A(n30746), .B(n30749), .Z(n30805) );
  XOR U30253 ( .A(n30856), .B(n30833), .Z(n30749) );
  XNOR U30254 ( .A(p_input[128]), .B(p_input[2048]), .Z(n30833) );
  XNOR U30255 ( .A(n30820), .B(n30819), .Z(n30856) );
  XNOR U30256 ( .A(n30857), .B(n30827), .Z(n30819) );
  XNOR U30257 ( .A(n30815), .B(n30814), .Z(n30827) );
  XNOR U30258 ( .A(n30858), .B(n30811), .Z(n30814) );
  XNOR U30259 ( .A(p_input[138]), .B(p_input[2058]), .Z(n30811) );
  XOR U30260 ( .A(p_input[139]), .B(n29030), .Z(n30858) );
  XOR U30261 ( .A(p_input[140]), .B(p_input[2060]), .Z(n30815) );
  XOR U30262 ( .A(n30825), .B(n30859), .Z(n30857) );
  IV U30263 ( .A(n30816), .Z(n30859) );
  XOR U30264 ( .A(p_input[129]), .B(p_input[2049]), .Z(n30816) );
  XNOR U30265 ( .A(n30860), .B(n30832), .Z(n30825) );
  XNOR U30266 ( .A(p_input[143]), .B(n29033), .Z(n30832) );
  XOR U30267 ( .A(n30822), .B(n30831), .Z(n30860) );
  XOR U30268 ( .A(n30861), .B(n30828), .Z(n30831) );
  XOR U30269 ( .A(p_input[141]), .B(p_input[2061]), .Z(n30828) );
  XOR U30270 ( .A(p_input[142]), .B(n29035), .Z(n30861) );
  XOR U30271 ( .A(p_input[137]), .B(p_input[2057]), .Z(n30822) );
  XOR U30272 ( .A(n30840), .B(n30838), .Z(n30820) );
  XNOR U30273 ( .A(n30862), .B(n30845), .Z(n30838) );
  XOR U30274 ( .A(p_input[136]), .B(p_input[2056]), .Z(n30845) );
  XOR U30275 ( .A(n30835), .B(n30844), .Z(n30862) );
  XOR U30276 ( .A(n30863), .B(n30841), .Z(n30844) );
  XOR U30277 ( .A(p_input[134]), .B(p_input[2054]), .Z(n30841) );
  XOR U30278 ( .A(p_input[135]), .B(n30404), .Z(n30863) );
  XOR U30279 ( .A(p_input[130]), .B(p_input[2050]), .Z(n30835) );
  XNOR U30280 ( .A(n30850), .B(n30849), .Z(n30840) );
  XOR U30281 ( .A(n30864), .B(n30846), .Z(n30849) );
  XOR U30282 ( .A(p_input[131]), .B(p_input[2051]), .Z(n30846) );
  XOR U30283 ( .A(p_input[132]), .B(n30406), .Z(n30864) );
  XOR U30284 ( .A(p_input[133]), .B(p_input[2053]), .Z(n30850) );
  XNOR U30285 ( .A(n30865), .B(n30866), .Z(n30746) );
  AND U30286 ( .A(n227), .B(n30867), .Z(n30866) );
  XNOR U30287 ( .A(n30868), .B(n30869), .Z(n227) );
  AND U30288 ( .A(n30870), .B(n30871), .Z(n30869) );
  XOR U30289 ( .A(n30760), .B(n30868), .Z(n30871) );
  XNOR U30290 ( .A(n30872), .B(n30868), .Z(n30870) );
  XOR U30291 ( .A(n30873), .B(n30874), .Z(n30868) );
  AND U30292 ( .A(n30875), .B(n30876), .Z(n30874) );
  XOR U30293 ( .A(n30775), .B(n30873), .Z(n30876) );
  XOR U30294 ( .A(n30873), .B(n30776), .Z(n30875) );
  XOR U30295 ( .A(n30877), .B(n30878), .Z(n30873) );
  AND U30296 ( .A(n30879), .B(n30880), .Z(n30878) );
  XOR U30297 ( .A(n30803), .B(n30877), .Z(n30880) );
  XOR U30298 ( .A(n30877), .B(n30804), .Z(n30879) );
  XOR U30299 ( .A(n30881), .B(n30882), .Z(n30877) );
  AND U30300 ( .A(n30883), .B(n30884), .Z(n30882) );
  XOR U30301 ( .A(n30881), .B(n30854), .Z(n30884) );
  XNOR U30302 ( .A(n30885), .B(n30886), .Z(n30706) );
  AND U30303 ( .A(n231), .B(n30887), .Z(n30886) );
  XNOR U30304 ( .A(n30888), .B(n30889), .Z(n231) );
  AND U30305 ( .A(n30890), .B(n30891), .Z(n30889) );
  XOR U30306 ( .A(n30888), .B(n30716), .Z(n30891) );
  XNOR U30307 ( .A(n30888), .B(n30676), .Z(n30890) );
  XOR U30308 ( .A(n30892), .B(n30893), .Z(n30888) );
  AND U30309 ( .A(n30894), .B(n30895), .Z(n30893) );
  XOR U30310 ( .A(n30892), .B(n30684), .Z(n30894) );
  XOR U30311 ( .A(n30896), .B(n30897), .Z(n30667) );
  AND U30312 ( .A(n235), .B(n30887), .Z(n30897) );
  XNOR U30313 ( .A(n30885), .B(n30896), .Z(n30887) );
  XNOR U30314 ( .A(n30898), .B(n30899), .Z(n235) );
  AND U30315 ( .A(n30900), .B(n30901), .Z(n30899) );
  XNOR U30316 ( .A(n30902), .B(n30898), .Z(n30901) );
  IV U30317 ( .A(n30716), .Z(n30902) );
  XOR U30318 ( .A(n30872), .B(n30903), .Z(n30716) );
  AND U30319 ( .A(n238), .B(n30904), .Z(n30903) );
  XOR U30320 ( .A(n30759), .B(n30756), .Z(n30904) );
  IV U30321 ( .A(n30872), .Z(n30759) );
  XNOR U30322 ( .A(n30676), .B(n30898), .Z(n30900) );
  XOR U30323 ( .A(n30905), .B(n30906), .Z(n30676) );
  AND U30324 ( .A(n254), .B(n30907), .Z(n30906) );
  XOR U30325 ( .A(n30892), .B(n30908), .Z(n30898) );
  AND U30326 ( .A(n30909), .B(n30895), .Z(n30908) );
  XNOR U30327 ( .A(n30726), .B(n30892), .Z(n30895) );
  XOR U30328 ( .A(n30776), .B(n30910), .Z(n30726) );
  AND U30329 ( .A(n238), .B(n30911), .Z(n30910) );
  XOR U30330 ( .A(n30772), .B(n30776), .Z(n30911) );
  XNOR U30331 ( .A(n30912), .B(n30892), .Z(n30909) );
  IV U30332 ( .A(n30684), .Z(n30912) );
  XOR U30333 ( .A(n30913), .B(n30914), .Z(n30684) );
  AND U30334 ( .A(n254), .B(n30915), .Z(n30914) );
  XOR U30335 ( .A(n30916), .B(n30917), .Z(n30892) );
  AND U30336 ( .A(n30918), .B(n30919), .Z(n30917) );
  XNOR U30337 ( .A(n30736), .B(n30916), .Z(n30919) );
  XOR U30338 ( .A(n30804), .B(n30920), .Z(n30736) );
  AND U30339 ( .A(n238), .B(n30921), .Z(n30920) );
  XOR U30340 ( .A(n30800), .B(n30804), .Z(n30921) );
  XOR U30341 ( .A(n30916), .B(n30693), .Z(n30918) );
  XOR U30342 ( .A(n30922), .B(n30923), .Z(n30693) );
  AND U30343 ( .A(n254), .B(n30924), .Z(n30923) );
  XOR U30344 ( .A(n30925), .B(n30926), .Z(n30916) );
  AND U30345 ( .A(n30927), .B(n30928), .Z(n30926) );
  XNOR U30346 ( .A(n30925), .B(n30744), .Z(n30928) );
  XOR U30347 ( .A(n30855), .B(n30929), .Z(n30744) );
  AND U30348 ( .A(n238), .B(n30930), .Z(n30929) );
  XOR U30349 ( .A(n30851), .B(n30855), .Z(n30930) );
  XNOR U30350 ( .A(n30931), .B(n30925), .Z(n30927) );
  IV U30351 ( .A(n30703), .Z(n30931) );
  XOR U30352 ( .A(n30932), .B(n30933), .Z(n30703) );
  AND U30353 ( .A(n254), .B(n30934), .Z(n30933) );
  AND U30354 ( .A(n30896), .B(n30885), .Z(n30925) );
  XNOR U30355 ( .A(n30935), .B(n30936), .Z(n30885) );
  AND U30356 ( .A(n238), .B(n30867), .Z(n30936) );
  XNOR U30357 ( .A(n30865), .B(n30935), .Z(n30867) );
  XNOR U30358 ( .A(n30937), .B(n30938), .Z(n238) );
  AND U30359 ( .A(n30939), .B(n30940), .Z(n30938) );
  XNOR U30360 ( .A(n30937), .B(n30756), .Z(n30940) );
  IV U30361 ( .A(n30760), .Z(n30756) );
  XOR U30362 ( .A(n30941), .B(n30942), .Z(n30760) );
  AND U30363 ( .A(n242), .B(n30943), .Z(n30942) );
  XOR U30364 ( .A(n30944), .B(n30941), .Z(n30943) );
  XNOR U30365 ( .A(n30937), .B(n30872), .Z(n30939) );
  XOR U30366 ( .A(n30945), .B(n30946), .Z(n30872) );
  AND U30367 ( .A(n250), .B(n30907), .Z(n30946) );
  XOR U30368 ( .A(n30905), .B(n30945), .Z(n30907) );
  XOR U30369 ( .A(n30947), .B(n30948), .Z(n30937) );
  AND U30370 ( .A(n30949), .B(n30950), .Z(n30948) );
  XNOR U30371 ( .A(n30947), .B(n30772), .Z(n30950) );
  IV U30372 ( .A(n30775), .Z(n30772) );
  XOR U30373 ( .A(n30951), .B(n30952), .Z(n30775) );
  AND U30374 ( .A(n242), .B(n30953), .Z(n30952) );
  XOR U30375 ( .A(n30954), .B(n30951), .Z(n30953) );
  XOR U30376 ( .A(n30776), .B(n30947), .Z(n30949) );
  XOR U30377 ( .A(n30955), .B(n30956), .Z(n30776) );
  AND U30378 ( .A(n250), .B(n30915), .Z(n30956) );
  XOR U30379 ( .A(n30955), .B(n30913), .Z(n30915) );
  XOR U30380 ( .A(n30957), .B(n30958), .Z(n30947) );
  AND U30381 ( .A(n30959), .B(n30960), .Z(n30958) );
  XNOR U30382 ( .A(n30957), .B(n30800), .Z(n30960) );
  IV U30383 ( .A(n30803), .Z(n30800) );
  XOR U30384 ( .A(n30961), .B(n30962), .Z(n30803) );
  AND U30385 ( .A(n242), .B(n30963), .Z(n30962) );
  XNOR U30386 ( .A(n30964), .B(n30961), .Z(n30963) );
  XOR U30387 ( .A(n30804), .B(n30957), .Z(n30959) );
  XOR U30388 ( .A(n30965), .B(n30966), .Z(n30804) );
  AND U30389 ( .A(n250), .B(n30924), .Z(n30966) );
  XOR U30390 ( .A(n30965), .B(n30922), .Z(n30924) );
  XOR U30391 ( .A(n30881), .B(n30967), .Z(n30957) );
  AND U30392 ( .A(n30883), .B(n30968), .Z(n30967) );
  XNOR U30393 ( .A(n30881), .B(n30851), .Z(n30968) );
  IV U30394 ( .A(n30854), .Z(n30851) );
  XOR U30395 ( .A(n30969), .B(n30970), .Z(n30854) );
  AND U30396 ( .A(n242), .B(n30971), .Z(n30970) );
  XOR U30397 ( .A(n30972), .B(n30969), .Z(n30971) );
  XOR U30398 ( .A(n30855), .B(n30881), .Z(n30883) );
  XOR U30399 ( .A(n30973), .B(n30974), .Z(n30855) );
  AND U30400 ( .A(n250), .B(n30934), .Z(n30974) );
  XOR U30401 ( .A(n30973), .B(n30932), .Z(n30934) );
  AND U30402 ( .A(n30935), .B(n30865), .Z(n30881) );
  XNOR U30403 ( .A(n30975), .B(n30976), .Z(n30865) );
  AND U30404 ( .A(n242), .B(n30977), .Z(n30976) );
  XNOR U30405 ( .A(n30978), .B(n30975), .Z(n30977) );
  XNOR U30406 ( .A(n30979), .B(n30980), .Z(n242) );
  AND U30407 ( .A(n30981), .B(n30982), .Z(n30980) );
  XOR U30408 ( .A(n30944), .B(n30979), .Z(n30982) );
  AND U30409 ( .A(n30983), .B(n30984), .Z(n30944) );
  XNOR U30410 ( .A(n30941), .B(n30979), .Z(n30981) );
  XNOR U30411 ( .A(n30985), .B(n30986), .Z(n30941) );
  AND U30412 ( .A(n246), .B(n30987), .Z(n30986) );
  XNOR U30413 ( .A(n30988), .B(n30989), .Z(n30987) );
  XOR U30414 ( .A(n30990), .B(n30991), .Z(n30979) );
  AND U30415 ( .A(n30992), .B(n30993), .Z(n30991) );
  XNOR U30416 ( .A(n30990), .B(n30983), .Z(n30993) );
  IV U30417 ( .A(n30954), .Z(n30983) );
  XOR U30418 ( .A(n30994), .B(n30995), .Z(n30954) );
  XOR U30419 ( .A(n30996), .B(n30984), .Z(n30995) );
  AND U30420 ( .A(n30964), .B(n30997), .Z(n30984) );
  AND U30421 ( .A(n30998), .B(n30999), .Z(n30996) );
  XOR U30422 ( .A(n31000), .B(n30994), .Z(n30998) );
  XNOR U30423 ( .A(n30951), .B(n30990), .Z(n30992) );
  XNOR U30424 ( .A(n31001), .B(n31002), .Z(n30951) );
  AND U30425 ( .A(n246), .B(n31003), .Z(n31002) );
  XNOR U30426 ( .A(n31004), .B(n31005), .Z(n31003) );
  XOR U30427 ( .A(n31006), .B(n31007), .Z(n30990) );
  AND U30428 ( .A(n31008), .B(n31009), .Z(n31007) );
  XNOR U30429 ( .A(n31006), .B(n30964), .Z(n31009) );
  XOR U30430 ( .A(n31010), .B(n30999), .Z(n30964) );
  XNOR U30431 ( .A(n31011), .B(n30994), .Z(n30999) );
  XOR U30432 ( .A(n31012), .B(n31013), .Z(n30994) );
  AND U30433 ( .A(n31014), .B(n31015), .Z(n31013) );
  XOR U30434 ( .A(n31016), .B(n31012), .Z(n31014) );
  XNOR U30435 ( .A(n31017), .B(n31018), .Z(n31011) );
  AND U30436 ( .A(n31019), .B(n31020), .Z(n31018) );
  XOR U30437 ( .A(n31017), .B(n31021), .Z(n31019) );
  XNOR U30438 ( .A(n31000), .B(n30997), .Z(n31010) );
  AND U30439 ( .A(n31022), .B(n31023), .Z(n30997) );
  XOR U30440 ( .A(n31024), .B(n31025), .Z(n31000) );
  AND U30441 ( .A(n31026), .B(n31027), .Z(n31025) );
  XOR U30442 ( .A(n31024), .B(n31028), .Z(n31026) );
  XNOR U30443 ( .A(n30961), .B(n31006), .Z(n31008) );
  XNOR U30444 ( .A(n31029), .B(n31030), .Z(n30961) );
  AND U30445 ( .A(n246), .B(n31031), .Z(n31030) );
  XNOR U30446 ( .A(n31032), .B(n31033), .Z(n31031) );
  XOR U30447 ( .A(n31034), .B(n31035), .Z(n31006) );
  AND U30448 ( .A(n31036), .B(n31037), .Z(n31035) );
  XNOR U30449 ( .A(n31034), .B(n31022), .Z(n31037) );
  IV U30450 ( .A(n30972), .Z(n31022) );
  XNOR U30451 ( .A(n31038), .B(n31015), .Z(n30972) );
  XNOR U30452 ( .A(n31039), .B(n31021), .Z(n31015) );
  XNOR U30453 ( .A(n31040), .B(n31041), .Z(n31021) );
  NOR U30454 ( .A(n31042), .B(n31043), .Z(n31041) );
  XOR U30455 ( .A(n31040), .B(n31044), .Z(n31042) );
  XNOR U30456 ( .A(n31020), .B(n31012), .Z(n31039) );
  XOR U30457 ( .A(n31045), .B(n31046), .Z(n31012) );
  AND U30458 ( .A(n31047), .B(n31048), .Z(n31046) );
  XOR U30459 ( .A(n31045), .B(n31049), .Z(n31047) );
  XNOR U30460 ( .A(n31050), .B(n31017), .Z(n31020) );
  XOR U30461 ( .A(n31051), .B(n31052), .Z(n31017) );
  AND U30462 ( .A(n31053), .B(n31054), .Z(n31052) );
  XNOR U30463 ( .A(n31055), .B(n31056), .Z(n31053) );
  IV U30464 ( .A(n31051), .Z(n31055) );
  XNOR U30465 ( .A(n31057), .B(n31058), .Z(n31050) );
  NOR U30466 ( .A(n31059), .B(n31060), .Z(n31058) );
  XNOR U30467 ( .A(n31057), .B(n31061), .Z(n31059) );
  XNOR U30468 ( .A(n31016), .B(n31023), .Z(n31038) );
  NOR U30469 ( .A(n30978), .B(n31062), .Z(n31023) );
  XOR U30470 ( .A(n31028), .B(n31027), .Z(n31016) );
  XNOR U30471 ( .A(n31063), .B(n31024), .Z(n31027) );
  XOR U30472 ( .A(n31064), .B(n31065), .Z(n31024) );
  AND U30473 ( .A(n31066), .B(n31067), .Z(n31065) );
  XNOR U30474 ( .A(n31068), .B(n31069), .Z(n31066) );
  IV U30475 ( .A(n31064), .Z(n31068) );
  XNOR U30476 ( .A(n31070), .B(n31071), .Z(n31063) );
  NOR U30477 ( .A(n31072), .B(n31073), .Z(n31071) );
  XNOR U30478 ( .A(n31070), .B(n31074), .Z(n31072) );
  XOR U30479 ( .A(n31075), .B(n31076), .Z(n31028) );
  NOR U30480 ( .A(n31077), .B(n31078), .Z(n31076) );
  XNOR U30481 ( .A(n31075), .B(n31079), .Z(n31077) );
  XNOR U30482 ( .A(n30969), .B(n31034), .Z(n31036) );
  XNOR U30483 ( .A(n31080), .B(n31081), .Z(n30969) );
  AND U30484 ( .A(n246), .B(n31082), .Z(n31081) );
  XNOR U30485 ( .A(n31083), .B(n31084), .Z(n31082) );
  AND U30486 ( .A(n30975), .B(n30978), .Z(n31034) );
  XOR U30487 ( .A(n31085), .B(n31062), .Z(n30978) );
  XNOR U30488 ( .A(p_input[144]), .B(p_input[2048]), .Z(n31062) );
  XNOR U30489 ( .A(n31049), .B(n31048), .Z(n31085) );
  XNOR U30490 ( .A(n31086), .B(n31056), .Z(n31048) );
  XNOR U30491 ( .A(n31044), .B(n31043), .Z(n31056) );
  XNOR U30492 ( .A(n31087), .B(n31040), .Z(n31043) );
  XNOR U30493 ( .A(p_input[154]), .B(p_input[2058]), .Z(n31040) );
  XOR U30494 ( .A(p_input[155]), .B(n29030), .Z(n31087) );
  XOR U30495 ( .A(p_input[156]), .B(p_input[2060]), .Z(n31044) );
  XOR U30496 ( .A(n31054), .B(n31088), .Z(n31086) );
  IV U30497 ( .A(n31045), .Z(n31088) );
  XOR U30498 ( .A(p_input[145]), .B(p_input[2049]), .Z(n31045) );
  XNOR U30499 ( .A(n31089), .B(n31061), .Z(n31054) );
  XNOR U30500 ( .A(p_input[159]), .B(n29033), .Z(n31061) );
  XOR U30501 ( .A(n31051), .B(n31060), .Z(n31089) );
  XOR U30502 ( .A(n31090), .B(n31057), .Z(n31060) );
  XOR U30503 ( .A(p_input[157]), .B(p_input[2061]), .Z(n31057) );
  XOR U30504 ( .A(p_input[158]), .B(n29035), .Z(n31090) );
  XOR U30505 ( .A(p_input[153]), .B(p_input[2057]), .Z(n31051) );
  XOR U30506 ( .A(n31069), .B(n31067), .Z(n31049) );
  XNOR U30507 ( .A(n31091), .B(n31074), .Z(n31067) );
  XOR U30508 ( .A(p_input[152]), .B(p_input[2056]), .Z(n31074) );
  XOR U30509 ( .A(n31064), .B(n31073), .Z(n31091) );
  XOR U30510 ( .A(n31092), .B(n31070), .Z(n31073) );
  XOR U30511 ( .A(p_input[150]), .B(p_input[2054]), .Z(n31070) );
  XOR U30512 ( .A(p_input[151]), .B(n30404), .Z(n31092) );
  XOR U30513 ( .A(p_input[146]), .B(p_input[2050]), .Z(n31064) );
  XNOR U30514 ( .A(n31079), .B(n31078), .Z(n31069) );
  XOR U30515 ( .A(n31093), .B(n31075), .Z(n31078) );
  XOR U30516 ( .A(p_input[147]), .B(p_input[2051]), .Z(n31075) );
  XOR U30517 ( .A(p_input[148]), .B(n30406), .Z(n31093) );
  XOR U30518 ( .A(p_input[149]), .B(p_input[2053]), .Z(n31079) );
  XNOR U30519 ( .A(n31094), .B(n31095), .Z(n30975) );
  AND U30520 ( .A(n246), .B(n31096), .Z(n31095) );
  XNOR U30521 ( .A(n31097), .B(n31098), .Z(n246) );
  AND U30522 ( .A(n31099), .B(n31100), .Z(n31098) );
  XOR U30523 ( .A(n30989), .B(n31097), .Z(n31100) );
  XNOR U30524 ( .A(n31101), .B(n31097), .Z(n31099) );
  XOR U30525 ( .A(n31102), .B(n31103), .Z(n31097) );
  AND U30526 ( .A(n31104), .B(n31105), .Z(n31103) );
  XOR U30527 ( .A(n31004), .B(n31102), .Z(n31105) );
  XOR U30528 ( .A(n31102), .B(n31005), .Z(n31104) );
  XOR U30529 ( .A(n31106), .B(n31107), .Z(n31102) );
  AND U30530 ( .A(n31108), .B(n31109), .Z(n31107) );
  XOR U30531 ( .A(n31032), .B(n31106), .Z(n31109) );
  XOR U30532 ( .A(n31106), .B(n31033), .Z(n31108) );
  XOR U30533 ( .A(n31110), .B(n31111), .Z(n31106) );
  AND U30534 ( .A(n31112), .B(n31113), .Z(n31111) );
  XOR U30535 ( .A(n31110), .B(n31083), .Z(n31113) );
  XNOR U30536 ( .A(n31114), .B(n31115), .Z(n30935) );
  AND U30537 ( .A(n250), .B(n31116), .Z(n31115) );
  XNOR U30538 ( .A(n31117), .B(n31118), .Z(n250) );
  AND U30539 ( .A(n31119), .B(n31120), .Z(n31118) );
  XOR U30540 ( .A(n31117), .B(n30945), .Z(n31120) );
  XNOR U30541 ( .A(n31117), .B(n30905), .Z(n31119) );
  XOR U30542 ( .A(n31121), .B(n31122), .Z(n31117) );
  AND U30543 ( .A(n31123), .B(n31124), .Z(n31122) );
  XOR U30544 ( .A(n31121), .B(n30913), .Z(n31123) );
  XOR U30545 ( .A(n31125), .B(n31126), .Z(n30896) );
  AND U30546 ( .A(n254), .B(n31116), .Z(n31126) );
  XNOR U30547 ( .A(n31114), .B(n31125), .Z(n31116) );
  XNOR U30548 ( .A(n31127), .B(n31128), .Z(n254) );
  AND U30549 ( .A(n31129), .B(n31130), .Z(n31128) );
  XNOR U30550 ( .A(n31131), .B(n31127), .Z(n31130) );
  IV U30551 ( .A(n30945), .Z(n31131) );
  XOR U30552 ( .A(n31101), .B(n31132), .Z(n30945) );
  AND U30553 ( .A(n257), .B(n31133), .Z(n31132) );
  XOR U30554 ( .A(n30988), .B(n30985), .Z(n31133) );
  IV U30555 ( .A(n31101), .Z(n30988) );
  XNOR U30556 ( .A(n30905), .B(n31127), .Z(n31129) );
  XOR U30557 ( .A(n31134), .B(n31135), .Z(n30905) );
  AND U30558 ( .A(n273), .B(n31136), .Z(n31135) );
  XOR U30559 ( .A(n31121), .B(n31137), .Z(n31127) );
  AND U30560 ( .A(n31138), .B(n31124), .Z(n31137) );
  XNOR U30561 ( .A(n30955), .B(n31121), .Z(n31124) );
  XOR U30562 ( .A(n31005), .B(n31139), .Z(n30955) );
  AND U30563 ( .A(n257), .B(n31140), .Z(n31139) );
  XOR U30564 ( .A(n31001), .B(n31005), .Z(n31140) );
  XNOR U30565 ( .A(n31141), .B(n31121), .Z(n31138) );
  IV U30566 ( .A(n30913), .Z(n31141) );
  XOR U30567 ( .A(n31142), .B(n31143), .Z(n30913) );
  AND U30568 ( .A(n273), .B(n31144), .Z(n31143) );
  XOR U30569 ( .A(n31145), .B(n31146), .Z(n31121) );
  AND U30570 ( .A(n31147), .B(n31148), .Z(n31146) );
  XNOR U30571 ( .A(n30965), .B(n31145), .Z(n31148) );
  XOR U30572 ( .A(n31033), .B(n31149), .Z(n30965) );
  AND U30573 ( .A(n257), .B(n31150), .Z(n31149) );
  XOR U30574 ( .A(n31029), .B(n31033), .Z(n31150) );
  XOR U30575 ( .A(n31145), .B(n30922), .Z(n31147) );
  XOR U30576 ( .A(n31151), .B(n31152), .Z(n30922) );
  AND U30577 ( .A(n273), .B(n31153), .Z(n31152) );
  XOR U30578 ( .A(n31154), .B(n31155), .Z(n31145) );
  AND U30579 ( .A(n31156), .B(n31157), .Z(n31155) );
  XNOR U30580 ( .A(n31154), .B(n30973), .Z(n31157) );
  XOR U30581 ( .A(n31084), .B(n31158), .Z(n30973) );
  AND U30582 ( .A(n257), .B(n31159), .Z(n31158) );
  XOR U30583 ( .A(n31080), .B(n31084), .Z(n31159) );
  XNOR U30584 ( .A(n31160), .B(n31154), .Z(n31156) );
  IV U30585 ( .A(n30932), .Z(n31160) );
  XOR U30586 ( .A(n31161), .B(n31162), .Z(n30932) );
  AND U30587 ( .A(n273), .B(n31163), .Z(n31162) );
  AND U30588 ( .A(n31125), .B(n31114), .Z(n31154) );
  XNOR U30589 ( .A(n31164), .B(n31165), .Z(n31114) );
  AND U30590 ( .A(n257), .B(n31096), .Z(n31165) );
  XNOR U30591 ( .A(n31094), .B(n31164), .Z(n31096) );
  XNOR U30592 ( .A(n31166), .B(n31167), .Z(n257) );
  AND U30593 ( .A(n31168), .B(n31169), .Z(n31167) );
  XNOR U30594 ( .A(n31166), .B(n30985), .Z(n31169) );
  IV U30595 ( .A(n30989), .Z(n30985) );
  XOR U30596 ( .A(n31170), .B(n31171), .Z(n30989) );
  AND U30597 ( .A(n261), .B(n31172), .Z(n31171) );
  XOR U30598 ( .A(n31173), .B(n31170), .Z(n31172) );
  XNOR U30599 ( .A(n31166), .B(n31101), .Z(n31168) );
  XOR U30600 ( .A(n31174), .B(n31175), .Z(n31101) );
  AND U30601 ( .A(n269), .B(n31136), .Z(n31175) );
  XOR U30602 ( .A(n31134), .B(n31174), .Z(n31136) );
  XOR U30603 ( .A(n31176), .B(n31177), .Z(n31166) );
  AND U30604 ( .A(n31178), .B(n31179), .Z(n31177) );
  XNOR U30605 ( .A(n31176), .B(n31001), .Z(n31179) );
  IV U30606 ( .A(n31004), .Z(n31001) );
  XOR U30607 ( .A(n31180), .B(n31181), .Z(n31004) );
  AND U30608 ( .A(n261), .B(n31182), .Z(n31181) );
  XOR U30609 ( .A(n31183), .B(n31180), .Z(n31182) );
  XOR U30610 ( .A(n31005), .B(n31176), .Z(n31178) );
  XOR U30611 ( .A(n31184), .B(n31185), .Z(n31005) );
  AND U30612 ( .A(n269), .B(n31144), .Z(n31185) );
  XOR U30613 ( .A(n31184), .B(n31142), .Z(n31144) );
  XOR U30614 ( .A(n31186), .B(n31187), .Z(n31176) );
  AND U30615 ( .A(n31188), .B(n31189), .Z(n31187) );
  XNOR U30616 ( .A(n31186), .B(n31029), .Z(n31189) );
  IV U30617 ( .A(n31032), .Z(n31029) );
  XOR U30618 ( .A(n31190), .B(n31191), .Z(n31032) );
  AND U30619 ( .A(n261), .B(n31192), .Z(n31191) );
  XNOR U30620 ( .A(n31193), .B(n31190), .Z(n31192) );
  XOR U30621 ( .A(n31033), .B(n31186), .Z(n31188) );
  XOR U30622 ( .A(n31194), .B(n31195), .Z(n31033) );
  AND U30623 ( .A(n269), .B(n31153), .Z(n31195) );
  XOR U30624 ( .A(n31194), .B(n31151), .Z(n31153) );
  XOR U30625 ( .A(n31110), .B(n31196), .Z(n31186) );
  AND U30626 ( .A(n31112), .B(n31197), .Z(n31196) );
  XNOR U30627 ( .A(n31110), .B(n31080), .Z(n31197) );
  IV U30628 ( .A(n31083), .Z(n31080) );
  XOR U30629 ( .A(n31198), .B(n31199), .Z(n31083) );
  AND U30630 ( .A(n261), .B(n31200), .Z(n31199) );
  XOR U30631 ( .A(n31201), .B(n31198), .Z(n31200) );
  XOR U30632 ( .A(n31084), .B(n31110), .Z(n31112) );
  XOR U30633 ( .A(n31202), .B(n31203), .Z(n31084) );
  AND U30634 ( .A(n269), .B(n31163), .Z(n31203) );
  XOR U30635 ( .A(n31202), .B(n31161), .Z(n31163) );
  AND U30636 ( .A(n31164), .B(n31094), .Z(n31110) );
  XNOR U30637 ( .A(n31204), .B(n31205), .Z(n31094) );
  AND U30638 ( .A(n261), .B(n31206), .Z(n31205) );
  XNOR U30639 ( .A(n31207), .B(n31204), .Z(n31206) );
  XNOR U30640 ( .A(n31208), .B(n31209), .Z(n261) );
  AND U30641 ( .A(n31210), .B(n31211), .Z(n31209) );
  XOR U30642 ( .A(n31173), .B(n31208), .Z(n31211) );
  AND U30643 ( .A(n31212), .B(n31213), .Z(n31173) );
  XNOR U30644 ( .A(n31170), .B(n31208), .Z(n31210) );
  XNOR U30645 ( .A(n31214), .B(n31215), .Z(n31170) );
  AND U30646 ( .A(n265), .B(n31216), .Z(n31215) );
  XNOR U30647 ( .A(n31217), .B(n31218), .Z(n31216) );
  XOR U30648 ( .A(n31219), .B(n31220), .Z(n31208) );
  AND U30649 ( .A(n31221), .B(n31222), .Z(n31220) );
  XNOR U30650 ( .A(n31219), .B(n31212), .Z(n31222) );
  IV U30651 ( .A(n31183), .Z(n31212) );
  XOR U30652 ( .A(n31223), .B(n31224), .Z(n31183) );
  XOR U30653 ( .A(n31225), .B(n31213), .Z(n31224) );
  AND U30654 ( .A(n31193), .B(n31226), .Z(n31213) );
  AND U30655 ( .A(n31227), .B(n31228), .Z(n31225) );
  XOR U30656 ( .A(n31229), .B(n31223), .Z(n31227) );
  XNOR U30657 ( .A(n31180), .B(n31219), .Z(n31221) );
  XNOR U30658 ( .A(n31230), .B(n31231), .Z(n31180) );
  AND U30659 ( .A(n265), .B(n31232), .Z(n31231) );
  XNOR U30660 ( .A(n31233), .B(n31234), .Z(n31232) );
  XOR U30661 ( .A(n31235), .B(n31236), .Z(n31219) );
  AND U30662 ( .A(n31237), .B(n31238), .Z(n31236) );
  XNOR U30663 ( .A(n31235), .B(n31193), .Z(n31238) );
  XOR U30664 ( .A(n31239), .B(n31228), .Z(n31193) );
  XNOR U30665 ( .A(n31240), .B(n31223), .Z(n31228) );
  XOR U30666 ( .A(n31241), .B(n31242), .Z(n31223) );
  AND U30667 ( .A(n31243), .B(n31244), .Z(n31242) );
  XOR U30668 ( .A(n31245), .B(n31241), .Z(n31243) );
  XNOR U30669 ( .A(n31246), .B(n31247), .Z(n31240) );
  AND U30670 ( .A(n31248), .B(n31249), .Z(n31247) );
  XOR U30671 ( .A(n31246), .B(n31250), .Z(n31248) );
  XNOR U30672 ( .A(n31229), .B(n31226), .Z(n31239) );
  AND U30673 ( .A(n31251), .B(n31252), .Z(n31226) );
  XOR U30674 ( .A(n31253), .B(n31254), .Z(n31229) );
  AND U30675 ( .A(n31255), .B(n31256), .Z(n31254) );
  XOR U30676 ( .A(n31253), .B(n31257), .Z(n31255) );
  XNOR U30677 ( .A(n31190), .B(n31235), .Z(n31237) );
  XNOR U30678 ( .A(n31258), .B(n31259), .Z(n31190) );
  AND U30679 ( .A(n265), .B(n31260), .Z(n31259) );
  XNOR U30680 ( .A(n31261), .B(n31262), .Z(n31260) );
  XOR U30681 ( .A(n31263), .B(n31264), .Z(n31235) );
  AND U30682 ( .A(n31265), .B(n31266), .Z(n31264) );
  XNOR U30683 ( .A(n31263), .B(n31251), .Z(n31266) );
  IV U30684 ( .A(n31201), .Z(n31251) );
  XNOR U30685 ( .A(n31267), .B(n31244), .Z(n31201) );
  XNOR U30686 ( .A(n31268), .B(n31250), .Z(n31244) );
  XNOR U30687 ( .A(n31269), .B(n31270), .Z(n31250) );
  NOR U30688 ( .A(n31271), .B(n31272), .Z(n31270) );
  XOR U30689 ( .A(n31269), .B(n31273), .Z(n31271) );
  XNOR U30690 ( .A(n31249), .B(n31241), .Z(n31268) );
  XOR U30691 ( .A(n31274), .B(n31275), .Z(n31241) );
  AND U30692 ( .A(n31276), .B(n31277), .Z(n31275) );
  XOR U30693 ( .A(n31274), .B(n31278), .Z(n31276) );
  XNOR U30694 ( .A(n31279), .B(n31246), .Z(n31249) );
  XOR U30695 ( .A(n31280), .B(n31281), .Z(n31246) );
  AND U30696 ( .A(n31282), .B(n31283), .Z(n31281) );
  XNOR U30697 ( .A(n31284), .B(n31285), .Z(n31282) );
  IV U30698 ( .A(n31280), .Z(n31284) );
  XNOR U30699 ( .A(n31286), .B(n31287), .Z(n31279) );
  NOR U30700 ( .A(n31288), .B(n31289), .Z(n31287) );
  XNOR U30701 ( .A(n31286), .B(n31290), .Z(n31288) );
  XNOR U30702 ( .A(n31245), .B(n31252), .Z(n31267) );
  NOR U30703 ( .A(n31207), .B(n31291), .Z(n31252) );
  XOR U30704 ( .A(n31257), .B(n31256), .Z(n31245) );
  XNOR U30705 ( .A(n31292), .B(n31253), .Z(n31256) );
  XOR U30706 ( .A(n31293), .B(n31294), .Z(n31253) );
  AND U30707 ( .A(n31295), .B(n31296), .Z(n31294) );
  XNOR U30708 ( .A(n31297), .B(n31298), .Z(n31295) );
  IV U30709 ( .A(n31293), .Z(n31297) );
  XNOR U30710 ( .A(n31299), .B(n31300), .Z(n31292) );
  NOR U30711 ( .A(n31301), .B(n31302), .Z(n31300) );
  XNOR U30712 ( .A(n31299), .B(n31303), .Z(n31301) );
  XOR U30713 ( .A(n31304), .B(n31305), .Z(n31257) );
  NOR U30714 ( .A(n31306), .B(n31307), .Z(n31305) );
  XNOR U30715 ( .A(n31304), .B(n31308), .Z(n31306) );
  XNOR U30716 ( .A(n31198), .B(n31263), .Z(n31265) );
  XNOR U30717 ( .A(n31309), .B(n31310), .Z(n31198) );
  AND U30718 ( .A(n265), .B(n31311), .Z(n31310) );
  XNOR U30719 ( .A(n31312), .B(n31313), .Z(n31311) );
  AND U30720 ( .A(n31204), .B(n31207), .Z(n31263) );
  XOR U30721 ( .A(n31314), .B(n31291), .Z(n31207) );
  XNOR U30722 ( .A(p_input[160]), .B(p_input[2048]), .Z(n31291) );
  XNOR U30723 ( .A(n31278), .B(n31277), .Z(n31314) );
  XNOR U30724 ( .A(n31315), .B(n31285), .Z(n31277) );
  XNOR U30725 ( .A(n31273), .B(n31272), .Z(n31285) );
  XNOR U30726 ( .A(n31316), .B(n31269), .Z(n31272) );
  XNOR U30727 ( .A(p_input[170]), .B(p_input[2058]), .Z(n31269) );
  XOR U30728 ( .A(p_input[171]), .B(n29030), .Z(n31316) );
  XOR U30729 ( .A(p_input[172]), .B(p_input[2060]), .Z(n31273) );
  XOR U30730 ( .A(n31283), .B(n31317), .Z(n31315) );
  IV U30731 ( .A(n31274), .Z(n31317) );
  XOR U30732 ( .A(p_input[161]), .B(p_input[2049]), .Z(n31274) );
  XNOR U30733 ( .A(n31318), .B(n31290), .Z(n31283) );
  XNOR U30734 ( .A(p_input[175]), .B(n29033), .Z(n31290) );
  XOR U30735 ( .A(n31280), .B(n31289), .Z(n31318) );
  XOR U30736 ( .A(n31319), .B(n31286), .Z(n31289) );
  XOR U30737 ( .A(p_input[173]), .B(p_input[2061]), .Z(n31286) );
  XOR U30738 ( .A(p_input[174]), .B(n29035), .Z(n31319) );
  XOR U30739 ( .A(p_input[169]), .B(p_input[2057]), .Z(n31280) );
  XOR U30740 ( .A(n31298), .B(n31296), .Z(n31278) );
  XNOR U30741 ( .A(n31320), .B(n31303), .Z(n31296) );
  XOR U30742 ( .A(p_input[168]), .B(p_input[2056]), .Z(n31303) );
  XOR U30743 ( .A(n31293), .B(n31302), .Z(n31320) );
  XOR U30744 ( .A(n31321), .B(n31299), .Z(n31302) );
  XOR U30745 ( .A(p_input[166]), .B(p_input[2054]), .Z(n31299) );
  XOR U30746 ( .A(p_input[167]), .B(n30404), .Z(n31321) );
  XOR U30747 ( .A(p_input[162]), .B(p_input[2050]), .Z(n31293) );
  XNOR U30748 ( .A(n31308), .B(n31307), .Z(n31298) );
  XOR U30749 ( .A(n31322), .B(n31304), .Z(n31307) );
  XOR U30750 ( .A(p_input[163]), .B(p_input[2051]), .Z(n31304) );
  XOR U30751 ( .A(p_input[164]), .B(n30406), .Z(n31322) );
  XOR U30752 ( .A(p_input[165]), .B(p_input[2053]), .Z(n31308) );
  XNOR U30753 ( .A(n31323), .B(n31324), .Z(n31204) );
  AND U30754 ( .A(n265), .B(n31325), .Z(n31324) );
  XNOR U30755 ( .A(n31326), .B(n31327), .Z(n265) );
  AND U30756 ( .A(n31328), .B(n31329), .Z(n31327) );
  XOR U30757 ( .A(n31218), .B(n31326), .Z(n31329) );
  XNOR U30758 ( .A(n31330), .B(n31326), .Z(n31328) );
  XOR U30759 ( .A(n31331), .B(n31332), .Z(n31326) );
  AND U30760 ( .A(n31333), .B(n31334), .Z(n31332) );
  XOR U30761 ( .A(n31233), .B(n31331), .Z(n31334) );
  XOR U30762 ( .A(n31331), .B(n31234), .Z(n31333) );
  XOR U30763 ( .A(n31335), .B(n31336), .Z(n31331) );
  AND U30764 ( .A(n31337), .B(n31338), .Z(n31336) );
  XOR U30765 ( .A(n31261), .B(n31335), .Z(n31338) );
  XOR U30766 ( .A(n31335), .B(n31262), .Z(n31337) );
  XOR U30767 ( .A(n31339), .B(n31340), .Z(n31335) );
  AND U30768 ( .A(n31341), .B(n31342), .Z(n31340) );
  XOR U30769 ( .A(n31339), .B(n31312), .Z(n31342) );
  XNOR U30770 ( .A(n31343), .B(n31344), .Z(n31164) );
  AND U30771 ( .A(n269), .B(n31345), .Z(n31344) );
  XNOR U30772 ( .A(n31346), .B(n31347), .Z(n269) );
  AND U30773 ( .A(n31348), .B(n31349), .Z(n31347) );
  XOR U30774 ( .A(n31346), .B(n31174), .Z(n31349) );
  XNOR U30775 ( .A(n31346), .B(n31134), .Z(n31348) );
  XOR U30776 ( .A(n31350), .B(n31351), .Z(n31346) );
  AND U30777 ( .A(n31352), .B(n31353), .Z(n31351) );
  XOR U30778 ( .A(n31350), .B(n31142), .Z(n31352) );
  XOR U30779 ( .A(n31354), .B(n31355), .Z(n31125) );
  AND U30780 ( .A(n273), .B(n31345), .Z(n31355) );
  XNOR U30781 ( .A(n31343), .B(n31354), .Z(n31345) );
  XNOR U30782 ( .A(n31356), .B(n31357), .Z(n273) );
  AND U30783 ( .A(n31358), .B(n31359), .Z(n31357) );
  XNOR U30784 ( .A(n31360), .B(n31356), .Z(n31359) );
  IV U30785 ( .A(n31174), .Z(n31360) );
  XOR U30786 ( .A(n31330), .B(n31361), .Z(n31174) );
  AND U30787 ( .A(n276), .B(n31362), .Z(n31361) );
  XOR U30788 ( .A(n31217), .B(n31214), .Z(n31362) );
  IV U30789 ( .A(n31330), .Z(n31217) );
  XNOR U30790 ( .A(n31134), .B(n31356), .Z(n31358) );
  XOR U30791 ( .A(n31363), .B(n31364), .Z(n31134) );
  AND U30792 ( .A(n292), .B(n31365), .Z(n31364) );
  XOR U30793 ( .A(n31350), .B(n31366), .Z(n31356) );
  AND U30794 ( .A(n31367), .B(n31353), .Z(n31366) );
  XNOR U30795 ( .A(n31184), .B(n31350), .Z(n31353) );
  XOR U30796 ( .A(n31234), .B(n31368), .Z(n31184) );
  AND U30797 ( .A(n276), .B(n31369), .Z(n31368) );
  XOR U30798 ( .A(n31230), .B(n31234), .Z(n31369) );
  XNOR U30799 ( .A(n31370), .B(n31350), .Z(n31367) );
  IV U30800 ( .A(n31142), .Z(n31370) );
  XOR U30801 ( .A(n31371), .B(n31372), .Z(n31142) );
  AND U30802 ( .A(n292), .B(n31373), .Z(n31372) );
  XOR U30803 ( .A(n31374), .B(n31375), .Z(n31350) );
  AND U30804 ( .A(n31376), .B(n31377), .Z(n31375) );
  XNOR U30805 ( .A(n31194), .B(n31374), .Z(n31377) );
  XOR U30806 ( .A(n31262), .B(n31378), .Z(n31194) );
  AND U30807 ( .A(n276), .B(n31379), .Z(n31378) );
  XOR U30808 ( .A(n31258), .B(n31262), .Z(n31379) );
  XOR U30809 ( .A(n31374), .B(n31151), .Z(n31376) );
  XOR U30810 ( .A(n31380), .B(n31381), .Z(n31151) );
  AND U30811 ( .A(n292), .B(n31382), .Z(n31381) );
  XOR U30812 ( .A(n31383), .B(n31384), .Z(n31374) );
  AND U30813 ( .A(n31385), .B(n31386), .Z(n31384) );
  XNOR U30814 ( .A(n31383), .B(n31202), .Z(n31386) );
  XOR U30815 ( .A(n31313), .B(n31387), .Z(n31202) );
  AND U30816 ( .A(n276), .B(n31388), .Z(n31387) );
  XOR U30817 ( .A(n31309), .B(n31313), .Z(n31388) );
  XNOR U30818 ( .A(n31389), .B(n31383), .Z(n31385) );
  IV U30819 ( .A(n31161), .Z(n31389) );
  XOR U30820 ( .A(n31390), .B(n31391), .Z(n31161) );
  AND U30821 ( .A(n292), .B(n31392), .Z(n31391) );
  AND U30822 ( .A(n31354), .B(n31343), .Z(n31383) );
  XNOR U30823 ( .A(n31393), .B(n31394), .Z(n31343) );
  AND U30824 ( .A(n276), .B(n31325), .Z(n31394) );
  XNOR U30825 ( .A(n31323), .B(n31393), .Z(n31325) );
  XNOR U30826 ( .A(n31395), .B(n31396), .Z(n276) );
  AND U30827 ( .A(n31397), .B(n31398), .Z(n31396) );
  XNOR U30828 ( .A(n31395), .B(n31214), .Z(n31398) );
  IV U30829 ( .A(n31218), .Z(n31214) );
  XOR U30830 ( .A(n31399), .B(n31400), .Z(n31218) );
  AND U30831 ( .A(n280), .B(n31401), .Z(n31400) );
  XOR U30832 ( .A(n31402), .B(n31399), .Z(n31401) );
  XNOR U30833 ( .A(n31395), .B(n31330), .Z(n31397) );
  XOR U30834 ( .A(n31403), .B(n31404), .Z(n31330) );
  AND U30835 ( .A(n288), .B(n31365), .Z(n31404) );
  XOR U30836 ( .A(n31363), .B(n31403), .Z(n31365) );
  XOR U30837 ( .A(n31405), .B(n31406), .Z(n31395) );
  AND U30838 ( .A(n31407), .B(n31408), .Z(n31406) );
  XNOR U30839 ( .A(n31405), .B(n31230), .Z(n31408) );
  IV U30840 ( .A(n31233), .Z(n31230) );
  XOR U30841 ( .A(n31409), .B(n31410), .Z(n31233) );
  AND U30842 ( .A(n280), .B(n31411), .Z(n31410) );
  XOR U30843 ( .A(n31412), .B(n31409), .Z(n31411) );
  XOR U30844 ( .A(n31234), .B(n31405), .Z(n31407) );
  XOR U30845 ( .A(n31413), .B(n31414), .Z(n31234) );
  AND U30846 ( .A(n288), .B(n31373), .Z(n31414) );
  XOR U30847 ( .A(n31413), .B(n31371), .Z(n31373) );
  XOR U30848 ( .A(n31415), .B(n31416), .Z(n31405) );
  AND U30849 ( .A(n31417), .B(n31418), .Z(n31416) );
  XNOR U30850 ( .A(n31415), .B(n31258), .Z(n31418) );
  IV U30851 ( .A(n31261), .Z(n31258) );
  XOR U30852 ( .A(n31419), .B(n31420), .Z(n31261) );
  AND U30853 ( .A(n280), .B(n31421), .Z(n31420) );
  XNOR U30854 ( .A(n31422), .B(n31419), .Z(n31421) );
  XOR U30855 ( .A(n31262), .B(n31415), .Z(n31417) );
  XOR U30856 ( .A(n31423), .B(n31424), .Z(n31262) );
  AND U30857 ( .A(n288), .B(n31382), .Z(n31424) );
  XOR U30858 ( .A(n31423), .B(n31380), .Z(n31382) );
  XOR U30859 ( .A(n31339), .B(n31425), .Z(n31415) );
  AND U30860 ( .A(n31341), .B(n31426), .Z(n31425) );
  XNOR U30861 ( .A(n31339), .B(n31309), .Z(n31426) );
  IV U30862 ( .A(n31312), .Z(n31309) );
  XOR U30863 ( .A(n31427), .B(n31428), .Z(n31312) );
  AND U30864 ( .A(n280), .B(n31429), .Z(n31428) );
  XOR U30865 ( .A(n31430), .B(n31427), .Z(n31429) );
  XOR U30866 ( .A(n31313), .B(n31339), .Z(n31341) );
  XOR U30867 ( .A(n31431), .B(n31432), .Z(n31313) );
  AND U30868 ( .A(n288), .B(n31392), .Z(n31432) );
  XOR U30869 ( .A(n31431), .B(n31390), .Z(n31392) );
  AND U30870 ( .A(n31393), .B(n31323), .Z(n31339) );
  XNOR U30871 ( .A(n31433), .B(n31434), .Z(n31323) );
  AND U30872 ( .A(n280), .B(n31435), .Z(n31434) );
  XNOR U30873 ( .A(n31436), .B(n31433), .Z(n31435) );
  XNOR U30874 ( .A(n31437), .B(n31438), .Z(n280) );
  AND U30875 ( .A(n31439), .B(n31440), .Z(n31438) );
  XOR U30876 ( .A(n31402), .B(n31437), .Z(n31440) );
  AND U30877 ( .A(n31441), .B(n31442), .Z(n31402) );
  XNOR U30878 ( .A(n31399), .B(n31437), .Z(n31439) );
  XNOR U30879 ( .A(n31443), .B(n31444), .Z(n31399) );
  AND U30880 ( .A(n284), .B(n31445), .Z(n31444) );
  XNOR U30881 ( .A(n31446), .B(n31447), .Z(n31445) );
  XOR U30882 ( .A(n31448), .B(n31449), .Z(n31437) );
  AND U30883 ( .A(n31450), .B(n31451), .Z(n31449) );
  XNOR U30884 ( .A(n31448), .B(n31441), .Z(n31451) );
  IV U30885 ( .A(n31412), .Z(n31441) );
  XOR U30886 ( .A(n31452), .B(n31453), .Z(n31412) );
  XOR U30887 ( .A(n31454), .B(n31442), .Z(n31453) );
  AND U30888 ( .A(n31422), .B(n31455), .Z(n31442) );
  AND U30889 ( .A(n31456), .B(n31457), .Z(n31454) );
  XOR U30890 ( .A(n31458), .B(n31452), .Z(n31456) );
  XNOR U30891 ( .A(n31409), .B(n31448), .Z(n31450) );
  XNOR U30892 ( .A(n31459), .B(n31460), .Z(n31409) );
  AND U30893 ( .A(n284), .B(n31461), .Z(n31460) );
  XNOR U30894 ( .A(n31462), .B(n31463), .Z(n31461) );
  XOR U30895 ( .A(n31464), .B(n31465), .Z(n31448) );
  AND U30896 ( .A(n31466), .B(n31467), .Z(n31465) );
  XNOR U30897 ( .A(n31464), .B(n31422), .Z(n31467) );
  XOR U30898 ( .A(n31468), .B(n31457), .Z(n31422) );
  XNOR U30899 ( .A(n31469), .B(n31452), .Z(n31457) );
  XOR U30900 ( .A(n31470), .B(n31471), .Z(n31452) );
  AND U30901 ( .A(n31472), .B(n31473), .Z(n31471) );
  XOR U30902 ( .A(n31474), .B(n31470), .Z(n31472) );
  XNOR U30903 ( .A(n31475), .B(n31476), .Z(n31469) );
  AND U30904 ( .A(n31477), .B(n31478), .Z(n31476) );
  XOR U30905 ( .A(n31475), .B(n31479), .Z(n31477) );
  XNOR U30906 ( .A(n31458), .B(n31455), .Z(n31468) );
  AND U30907 ( .A(n31480), .B(n31481), .Z(n31455) );
  XOR U30908 ( .A(n31482), .B(n31483), .Z(n31458) );
  AND U30909 ( .A(n31484), .B(n31485), .Z(n31483) );
  XOR U30910 ( .A(n31482), .B(n31486), .Z(n31484) );
  XNOR U30911 ( .A(n31419), .B(n31464), .Z(n31466) );
  XNOR U30912 ( .A(n31487), .B(n31488), .Z(n31419) );
  AND U30913 ( .A(n284), .B(n31489), .Z(n31488) );
  XNOR U30914 ( .A(n31490), .B(n31491), .Z(n31489) );
  XOR U30915 ( .A(n31492), .B(n31493), .Z(n31464) );
  AND U30916 ( .A(n31494), .B(n31495), .Z(n31493) );
  XNOR U30917 ( .A(n31492), .B(n31480), .Z(n31495) );
  IV U30918 ( .A(n31430), .Z(n31480) );
  XNOR U30919 ( .A(n31496), .B(n31473), .Z(n31430) );
  XNOR U30920 ( .A(n31497), .B(n31479), .Z(n31473) );
  XNOR U30921 ( .A(n31498), .B(n31499), .Z(n31479) );
  NOR U30922 ( .A(n31500), .B(n31501), .Z(n31499) );
  XOR U30923 ( .A(n31498), .B(n31502), .Z(n31500) );
  XNOR U30924 ( .A(n31478), .B(n31470), .Z(n31497) );
  XOR U30925 ( .A(n31503), .B(n31504), .Z(n31470) );
  AND U30926 ( .A(n31505), .B(n31506), .Z(n31504) );
  XOR U30927 ( .A(n31503), .B(n31507), .Z(n31505) );
  XNOR U30928 ( .A(n31508), .B(n31475), .Z(n31478) );
  XOR U30929 ( .A(n31509), .B(n31510), .Z(n31475) );
  AND U30930 ( .A(n31511), .B(n31512), .Z(n31510) );
  XNOR U30931 ( .A(n31513), .B(n31514), .Z(n31511) );
  IV U30932 ( .A(n31509), .Z(n31513) );
  XNOR U30933 ( .A(n31515), .B(n31516), .Z(n31508) );
  NOR U30934 ( .A(n31517), .B(n31518), .Z(n31516) );
  XNOR U30935 ( .A(n31515), .B(n31519), .Z(n31517) );
  XNOR U30936 ( .A(n31474), .B(n31481), .Z(n31496) );
  NOR U30937 ( .A(n31436), .B(n31520), .Z(n31481) );
  XOR U30938 ( .A(n31486), .B(n31485), .Z(n31474) );
  XNOR U30939 ( .A(n31521), .B(n31482), .Z(n31485) );
  XOR U30940 ( .A(n31522), .B(n31523), .Z(n31482) );
  AND U30941 ( .A(n31524), .B(n31525), .Z(n31523) );
  XNOR U30942 ( .A(n31526), .B(n31527), .Z(n31524) );
  IV U30943 ( .A(n31522), .Z(n31526) );
  XNOR U30944 ( .A(n31528), .B(n31529), .Z(n31521) );
  NOR U30945 ( .A(n31530), .B(n31531), .Z(n31529) );
  XNOR U30946 ( .A(n31528), .B(n31532), .Z(n31530) );
  XOR U30947 ( .A(n31533), .B(n31534), .Z(n31486) );
  NOR U30948 ( .A(n31535), .B(n31536), .Z(n31534) );
  XNOR U30949 ( .A(n31533), .B(n31537), .Z(n31535) );
  XNOR U30950 ( .A(n31427), .B(n31492), .Z(n31494) );
  XNOR U30951 ( .A(n31538), .B(n31539), .Z(n31427) );
  AND U30952 ( .A(n284), .B(n31540), .Z(n31539) );
  XNOR U30953 ( .A(n31541), .B(n31542), .Z(n31540) );
  AND U30954 ( .A(n31433), .B(n31436), .Z(n31492) );
  XOR U30955 ( .A(n31543), .B(n31520), .Z(n31436) );
  XNOR U30956 ( .A(p_input[176]), .B(p_input[2048]), .Z(n31520) );
  XNOR U30957 ( .A(n31507), .B(n31506), .Z(n31543) );
  XNOR U30958 ( .A(n31544), .B(n31514), .Z(n31506) );
  XNOR U30959 ( .A(n31502), .B(n31501), .Z(n31514) );
  XNOR U30960 ( .A(n31545), .B(n31498), .Z(n31501) );
  XNOR U30961 ( .A(p_input[186]), .B(p_input[2058]), .Z(n31498) );
  XOR U30962 ( .A(p_input[187]), .B(n29030), .Z(n31545) );
  XOR U30963 ( .A(p_input[188]), .B(p_input[2060]), .Z(n31502) );
  XOR U30964 ( .A(n31512), .B(n31546), .Z(n31544) );
  IV U30965 ( .A(n31503), .Z(n31546) );
  XOR U30966 ( .A(p_input[177]), .B(p_input[2049]), .Z(n31503) );
  XNOR U30967 ( .A(n31547), .B(n31519), .Z(n31512) );
  XNOR U30968 ( .A(p_input[191]), .B(n29033), .Z(n31519) );
  XOR U30969 ( .A(n31509), .B(n31518), .Z(n31547) );
  XOR U30970 ( .A(n31548), .B(n31515), .Z(n31518) );
  XOR U30971 ( .A(p_input[189]), .B(p_input[2061]), .Z(n31515) );
  XOR U30972 ( .A(p_input[190]), .B(n29035), .Z(n31548) );
  XOR U30973 ( .A(p_input[185]), .B(p_input[2057]), .Z(n31509) );
  XOR U30974 ( .A(n31527), .B(n31525), .Z(n31507) );
  XNOR U30975 ( .A(n31549), .B(n31532), .Z(n31525) );
  XOR U30976 ( .A(p_input[184]), .B(p_input[2056]), .Z(n31532) );
  XOR U30977 ( .A(n31522), .B(n31531), .Z(n31549) );
  XOR U30978 ( .A(n31550), .B(n31528), .Z(n31531) );
  XOR U30979 ( .A(p_input[182]), .B(p_input[2054]), .Z(n31528) );
  XOR U30980 ( .A(p_input[183]), .B(n30404), .Z(n31550) );
  XOR U30981 ( .A(p_input[178]), .B(p_input[2050]), .Z(n31522) );
  XNOR U30982 ( .A(n31537), .B(n31536), .Z(n31527) );
  XOR U30983 ( .A(n31551), .B(n31533), .Z(n31536) );
  XOR U30984 ( .A(p_input[179]), .B(p_input[2051]), .Z(n31533) );
  XOR U30985 ( .A(p_input[180]), .B(n30406), .Z(n31551) );
  XOR U30986 ( .A(p_input[181]), .B(p_input[2053]), .Z(n31537) );
  XNOR U30987 ( .A(n31552), .B(n31553), .Z(n31433) );
  AND U30988 ( .A(n284), .B(n31554), .Z(n31553) );
  XNOR U30989 ( .A(n31555), .B(n31556), .Z(n284) );
  AND U30990 ( .A(n31557), .B(n31558), .Z(n31556) );
  XOR U30991 ( .A(n31447), .B(n31555), .Z(n31558) );
  XNOR U30992 ( .A(n31559), .B(n31555), .Z(n31557) );
  XOR U30993 ( .A(n31560), .B(n31561), .Z(n31555) );
  AND U30994 ( .A(n31562), .B(n31563), .Z(n31561) );
  XOR U30995 ( .A(n31462), .B(n31560), .Z(n31563) );
  XOR U30996 ( .A(n31560), .B(n31463), .Z(n31562) );
  XOR U30997 ( .A(n31564), .B(n31565), .Z(n31560) );
  AND U30998 ( .A(n31566), .B(n31567), .Z(n31565) );
  XOR U30999 ( .A(n31490), .B(n31564), .Z(n31567) );
  XOR U31000 ( .A(n31564), .B(n31491), .Z(n31566) );
  XOR U31001 ( .A(n31568), .B(n31569), .Z(n31564) );
  AND U31002 ( .A(n31570), .B(n31571), .Z(n31569) );
  XOR U31003 ( .A(n31568), .B(n31541), .Z(n31571) );
  XNOR U31004 ( .A(n31572), .B(n31573), .Z(n31393) );
  AND U31005 ( .A(n288), .B(n31574), .Z(n31573) );
  XNOR U31006 ( .A(n31575), .B(n31576), .Z(n288) );
  AND U31007 ( .A(n31577), .B(n31578), .Z(n31576) );
  XOR U31008 ( .A(n31575), .B(n31403), .Z(n31578) );
  XNOR U31009 ( .A(n31575), .B(n31363), .Z(n31577) );
  XOR U31010 ( .A(n31579), .B(n31580), .Z(n31575) );
  AND U31011 ( .A(n31581), .B(n31582), .Z(n31580) );
  XOR U31012 ( .A(n31579), .B(n31371), .Z(n31581) );
  XOR U31013 ( .A(n31583), .B(n31584), .Z(n31354) );
  AND U31014 ( .A(n292), .B(n31574), .Z(n31584) );
  XNOR U31015 ( .A(n31572), .B(n31583), .Z(n31574) );
  XNOR U31016 ( .A(n31585), .B(n31586), .Z(n292) );
  AND U31017 ( .A(n31587), .B(n31588), .Z(n31586) );
  XNOR U31018 ( .A(n31589), .B(n31585), .Z(n31588) );
  IV U31019 ( .A(n31403), .Z(n31589) );
  XOR U31020 ( .A(n31559), .B(n31590), .Z(n31403) );
  AND U31021 ( .A(n295), .B(n31591), .Z(n31590) );
  XOR U31022 ( .A(n31446), .B(n31443), .Z(n31591) );
  IV U31023 ( .A(n31559), .Z(n31446) );
  XNOR U31024 ( .A(n31363), .B(n31585), .Z(n31587) );
  XOR U31025 ( .A(n31592), .B(n31593), .Z(n31363) );
  AND U31026 ( .A(n311), .B(n31594), .Z(n31593) );
  XOR U31027 ( .A(n31579), .B(n31595), .Z(n31585) );
  AND U31028 ( .A(n31596), .B(n31582), .Z(n31595) );
  XNOR U31029 ( .A(n31413), .B(n31579), .Z(n31582) );
  XOR U31030 ( .A(n31463), .B(n31597), .Z(n31413) );
  AND U31031 ( .A(n295), .B(n31598), .Z(n31597) );
  XOR U31032 ( .A(n31459), .B(n31463), .Z(n31598) );
  XNOR U31033 ( .A(n31599), .B(n31579), .Z(n31596) );
  IV U31034 ( .A(n31371), .Z(n31599) );
  XOR U31035 ( .A(n31600), .B(n31601), .Z(n31371) );
  AND U31036 ( .A(n311), .B(n31602), .Z(n31601) );
  XOR U31037 ( .A(n31603), .B(n31604), .Z(n31579) );
  AND U31038 ( .A(n31605), .B(n31606), .Z(n31604) );
  XNOR U31039 ( .A(n31423), .B(n31603), .Z(n31606) );
  XOR U31040 ( .A(n31491), .B(n31607), .Z(n31423) );
  AND U31041 ( .A(n295), .B(n31608), .Z(n31607) );
  XOR U31042 ( .A(n31487), .B(n31491), .Z(n31608) );
  XOR U31043 ( .A(n31603), .B(n31380), .Z(n31605) );
  XOR U31044 ( .A(n31609), .B(n31610), .Z(n31380) );
  AND U31045 ( .A(n311), .B(n31611), .Z(n31610) );
  XOR U31046 ( .A(n31612), .B(n31613), .Z(n31603) );
  AND U31047 ( .A(n31614), .B(n31615), .Z(n31613) );
  XNOR U31048 ( .A(n31612), .B(n31431), .Z(n31615) );
  XOR U31049 ( .A(n31542), .B(n31616), .Z(n31431) );
  AND U31050 ( .A(n295), .B(n31617), .Z(n31616) );
  XOR U31051 ( .A(n31538), .B(n31542), .Z(n31617) );
  XNOR U31052 ( .A(n31618), .B(n31612), .Z(n31614) );
  IV U31053 ( .A(n31390), .Z(n31618) );
  XOR U31054 ( .A(n31619), .B(n31620), .Z(n31390) );
  AND U31055 ( .A(n311), .B(n31621), .Z(n31620) );
  AND U31056 ( .A(n31583), .B(n31572), .Z(n31612) );
  XNOR U31057 ( .A(n31622), .B(n31623), .Z(n31572) );
  AND U31058 ( .A(n295), .B(n31554), .Z(n31623) );
  XNOR U31059 ( .A(n31552), .B(n31622), .Z(n31554) );
  XNOR U31060 ( .A(n31624), .B(n31625), .Z(n295) );
  AND U31061 ( .A(n31626), .B(n31627), .Z(n31625) );
  XNOR U31062 ( .A(n31624), .B(n31443), .Z(n31627) );
  IV U31063 ( .A(n31447), .Z(n31443) );
  XOR U31064 ( .A(n31628), .B(n31629), .Z(n31447) );
  AND U31065 ( .A(n299), .B(n31630), .Z(n31629) );
  XOR U31066 ( .A(n31631), .B(n31628), .Z(n31630) );
  XNOR U31067 ( .A(n31624), .B(n31559), .Z(n31626) );
  XOR U31068 ( .A(n31632), .B(n31633), .Z(n31559) );
  AND U31069 ( .A(n307), .B(n31594), .Z(n31633) );
  XOR U31070 ( .A(n31592), .B(n31632), .Z(n31594) );
  XOR U31071 ( .A(n31634), .B(n31635), .Z(n31624) );
  AND U31072 ( .A(n31636), .B(n31637), .Z(n31635) );
  XNOR U31073 ( .A(n31634), .B(n31459), .Z(n31637) );
  IV U31074 ( .A(n31462), .Z(n31459) );
  XOR U31075 ( .A(n31638), .B(n31639), .Z(n31462) );
  AND U31076 ( .A(n299), .B(n31640), .Z(n31639) );
  XOR U31077 ( .A(n31641), .B(n31638), .Z(n31640) );
  XOR U31078 ( .A(n31463), .B(n31634), .Z(n31636) );
  XOR U31079 ( .A(n31642), .B(n31643), .Z(n31463) );
  AND U31080 ( .A(n307), .B(n31602), .Z(n31643) );
  XOR U31081 ( .A(n31642), .B(n31600), .Z(n31602) );
  XOR U31082 ( .A(n31644), .B(n31645), .Z(n31634) );
  AND U31083 ( .A(n31646), .B(n31647), .Z(n31645) );
  XNOR U31084 ( .A(n31644), .B(n31487), .Z(n31647) );
  IV U31085 ( .A(n31490), .Z(n31487) );
  XOR U31086 ( .A(n31648), .B(n31649), .Z(n31490) );
  AND U31087 ( .A(n299), .B(n31650), .Z(n31649) );
  XNOR U31088 ( .A(n31651), .B(n31648), .Z(n31650) );
  XOR U31089 ( .A(n31491), .B(n31644), .Z(n31646) );
  XOR U31090 ( .A(n31652), .B(n31653), .Z(n31491) );
  AND U31091 ( .A(n307), .B(n31611), .Z(n31653) );
  XOR U31092 ( .A(n31652), .B(n31609), .Z(n31611) );
  XOR U31093 ( .A(n31568), .B(n31654), .Z(n31644) );
  AND U31094 ( .A(n31570), .B(n31655), .Z(n31654) );
  XNOR U31095 ( .A(n31568), .B(n31538), .Z(n31655) );
  IV U31096 ( .A(n31541), .Z(n31538) );
  XOR U31097 ( .A(n31656), .B(n31657), .Z(n31541) );
  AND U31098 ( .A(n299), .B(n31658), .Z(n31657) );
  XOR U31099 ( .A(n31659), .B(n31656), .Z(n31658) );
  XOR U31100 ( .A(n31542), .B(n31568), .Z(n31570) );
  XOR U31101 ( .A(n31660), .B(n31661), .Z(n31542) );
  AND U31102 ( .A(n307), .B(n31621), .Z(n31661) );
  XOR U31103 ( .A(n31660), .B(n31619), .Z(n31621) );
  AND U31104 ( .A(n31622), .B(n31552), .Z(n31568) );
  XNOR U31105 ( .A(n31662), .B(n31663), .Z(n31552) );
  AND U31106 ( .A(n299), .B(n31664), .Z(n31663) );
  XNOR U31107 ( .A(n31665), .B(n31662), .Z(n31664) );
  XNOR U31108 ( .A(n31666), .B(n31667), .Z(n299) );
  AND U31109 ( .A(n31668), .B(n31669), .Z(n31667) );
  XOR U31110 ( .A(n31631), .B(n31666), .Z(n31669) );
  AND U31111 ( .A(n31670), .B(n31671), .Z(n31631) );
  XNOR U31112 ( .A(n31628), .B(n31666), .Z(n31668) );
  XNOR U31113 ( .A(n31672), .B(n31673), .Z(n31628) );
  AND U31114 ( .A(n303), .B(n31674), .Z(n31673) );
  XNOR U31115 ( .A(n31675), .B(n31676), .Z(n31674) );
  XOR U31116 ( .A(n31677), .B(n31678), .Z(n31666) );
  AND U31117 ( .A(n31679), .B(n31680), .Z(n31678) );
  XNOR U31118 ( .A(n31677), .B(n31670), .Z(n31680) );
  IV U31119 ( .A(n31641), .Z(n31670) );
  XOR U31120 ( .A(n31681), .B(n31682), .Z(n31641) );
  XOR U31121 ( .A(n31683), .B(n31671), .Z(n31682) );
  AND U31122 ( .A(n31651), .B(n31684), .Z(n31671) );
  AND U31123 ( .A(n31685), .B(n31686), .Z(n31683) );
  XOR U31124 ( .A(n31687), .B(n31681), .Z(n31685) );
  XNOR U31125 ( .A(n31638), .B(n31677), .Z(n31679) );
  XNOR U31126 ( .A(n31688), .B(n31689), .Z(n31638) );
  AND U31127 ( .A(n303), .B(n31690), .Z(n31689) );
  XNOR U31128 ( .A(n31691), .B(n31692), .Z(n31690) );
  XOR U31129 ( .A(n31693), .B(n31694), .Z(n31677) );
  AND U31130 ( .A(n31695), .B(n31696), .Z(n31694) );
  XNOR U31131 ( .A(n31693), .B(n31651), .Z(n31696) );
  XOR U31132 ( .A(n31697), .B(n31686), .Z(n31651) );
  XNOR U31133 ( .A(n31698), .B(n31681), .Z(n31686) );
  XOR U31134 ( .A(n31699), .B(n31700), .Z(n31681) );
  AND U31135 ( .A(n31701), .B(n31702), .Z(n31700) );
  XOR U31136 ( .A(n31703), .B(n31699), .Z(n31701) );
  XNOR U31137 ( .A(n31704), .B(n31705), .Z(n31698) );
  AND U31138 ( .A(n31706), .B(n31707), .Z(n31705) );
  XOR U31139 ( .A(n31704), .B(n31708), .Z(n31706) );
  XNOR U31140 ( .A(n31687), .B(n31684), .Z(n31697) );
  AND U31141 ( .A(n31709), .B(n31710), .Z(n31684) );
  XOR U31142 ( .A(n31711), .B(n31712), .Z(n31687) );
  AND U31143 ( .A(n31713), .B(n31714), .Z(n31712) );
  XOR U31144 ( .A(n31711), .B(n31715), .Z(n31713) );
  XNOR U31145 ( .A(n31648), .B(n31693), .Z(n31695) );
  XNOR U31146 ( .A(n31716), .B(n31717), .Z(n31648) );
  AND U31147 ( .A(n303), .B(n31718), .Z(n31717) );
  XNOR U31148 ( .A(n31719), .B(n31720), .Z(n31718) );
  XOR U31149 ( .A(n31721), .B(n31722), .Z(n31693) );
  AND U31150 ( .A(n31723), .B(n31724), .Z(n31722) );
  XNOR U31151 ( .A(n31721), .B(n31709), .Z(n31724) );
  IV U31152 ( .A(n31659), .Z(n31709) );
  XNOR U31153 ( .A(n31725), .B(n31702), .Z(n31659) );
  XNOR U31154 ( .A(n31726), .B(n31708), .Z(n31702) );
  XNOR U31155 ( .A(n31727), .B(n31728), .Z(n31708) );
  NOR U31156 ( .A(n31729), .B(n31730), .Z(n31728) );
  XOR U31157 ( .A(n31727), .B(n31731), .Z(n31729) );
  XNOR U31158 ( .A(n31707), .B(n31699), .Z(n31726) );
  XOR U31159 ( .A(n31732), .B(n31733), .Z(n31699) );
  AND U31160 ( .A(n31734), .B(n31735), .Z(n31733) );
  XOR U31161 ( .A(n31732), .B(n31736), .Z(n31734) );
  XNOR U31162 ( .A(n31737), .B(n31704), .Z(n31707) );
  XOR U31163 ( .A(n31738), .B(n31739), .Z(n31704) );
  AND U31164 ( .A(n31740), .B(n31741), .Z(n31739) );
  XNOR U31165 ( .A(n31742), .B(n31743), .Z(n31740) );
  IV U31166 ( .A(n31738), .Z(n31742) );
  XNOR U31167 ( .A(n31744), .B(n31745), .Z(n31737) );
  NOR U31168 ( .A(n31746), .B(n31747), .Z(n31745) );
  XOR U31169 ( .A(n31744), .B(n31748), .Z(n31746) );
  XNOR U31170 ( .A(n31703), .B(n31710), .Z(n31725) );
  NOR U31171 ( .A(n31665), .B(n31749), .Z(n31710) );
  XOR U31172 ( .A(n31715), .B(n31714), .Z(n31703) );
  XNOR U31173 ( .A(n31750), .B(n31711), .Z(n31714) );
  XOR U31174 ( .A(n31751), .B(n31752), .Z(n31711) );
  AND U31175 ( .A(n31753), .B(n31754), .Z(n31752) );
  XNOR U31176 ( .A(n31755), .B(n31756), .Z(n31753) );
  IV U31177 ( .A(n31751), .Z(n31755) );
  XNOR U31178 ( .A(n31757), .B(n31758), .Z(n31750) );
  NOR U31179 ( .A(n31759), .B(n31760), .Z(n31758) );
  XNOR U31180 ( .A(n31757), .B(n31761), .Z(n31759) );
  XOR U31181 ( .A(n31762), .B(n31763), .Z(n31715) );
  NOR U31182 ( .A(n31764), .B(n31765), .Z(n31763) );
  XNOR U31183 ( .A(n31762), .B(n31766), .Z(n31764) );
  XNOR U31184 ( .A(n31656), .B(n31721), .Z(n31723) );
  XNOR U31185 ( .A(n31767), .B(n31768), .Z(n31656) );
  AND U31186 ( .A(n303), .B(n31769), .Z(n31768) );
  XNOR U31187 ( .A(n31770), .B(n31771), .Z(n31769) );
  AND U31188 ( .A(n31662), .B(n31665), .Z(n31721) );
  XOR U31189 ( .A(n31772), .B(n31749), .Z(n31665) );
  XNOR U31190 ( .A(p_input[192]), .B(p_input[2048]), .Z(n31749) );
  XNOR U31191 ( .A(n31736), .B(n31735), .Z(n31772) );
  XNOR U31192 ( .A(n31773), .B(n31743), .Z(n31735) );
  XNOR U31193 ( .A(n31731), .B(n31730), .Z(n31743) );
  XNOR U31194 ( .A(n31774), .B(n31727), .Z(n31730) );
  XNOR U31195 ( .A(p_input[202]), .B(p_input[2058]), .Z(n31727) );
  XOR U31196 ( .A(p_input[203]), .B(n29030), .Z(n31774) );
  XOR U31197 ( .A(p_input[204]), .B(p_input[2060]), .Z(n31731) );
  XOR U31198 ( .A(n31741), .B(n31775), .Z(n31773) );
  IV U31199 ( .A(n31732), .Z(n31775) );
  XOR U31200 ( .A(p_input[193]), .B(p_input[2049]), .Z(n31732) );
  XOR U31201 ( .A(n31776), .B(n31748), .Z(n31741) );
  XNOR U31202 ( .A(p_input[2063]), .B(p_input[207]), .Z(n31748) );
  XOR U31203 ( .A(n31738), .B(n31747), .Z(n31776) );
  XOR U31204 ( .A(n31777), .B(n31744), .Z(n31747) );
  XOR U31205 ( .A(p_input[205]), .B(p_input[2061]), .Z(n31744) );
  XNOR U31206 ( .A(p_input[2062]), .B(p_input[206]), .Z(n31777) );
  XOR U31207 ( .A(p_input[201]), .B(p_input[2057]), .Z(n31738) );
  XOR U31208 ( .A(n31756), .B(n31754), .Z(n31736) );
  XNOR U31209 ( .A(n31778), .B(n31761), .Z(n31754) );
  XOR U31210 ( .A(p_input[200]), .B(p_input[2056]), .Z(n31761) );
  XOR U31211 ( .A(n31751), .B(n31760), .Z(n31778) );
  XOR U31212 ( .A(n31779), .B(n31757), .Z(n31760) );
  XOR U31213 ( .A(p_input[198]), .B(p_input[2054]), .Z(n31757) );
  XOR U31214 ( .A(p_input[199]), .B(n30404), .Z(n31779) );
  XOR U31215 ( .A(p_input[194]), .B(p_input[2050]), .Z(n31751) );
  XNOR U31216 ( .A(n31766), .B(n31765), .Z(n31756) );
  XOR U31217 ( .A(n31780), .B(n31762), .Z(n31765) );
  XOR U31218 ( .A(p_input[195]), .B(p_input[2051]), .Z(n31762) );
  XOR U31219 ( .A(p_input[196]), .B(n30406), .Z(n31780) );
  XOR U31220 ( .A(p_input[197]), .B(p_input[2053]), .Z(n31766) );
  XNOR U31221 ( .A(n31781), .B(n31782), .Z(n31662) );
  AND U31222 ( .A(n303), .B(n31783), .Z(n31782) );
  XNOR U31223 ( .A(n31784), .B(n31785), .Z(n303) );
  AND U31224 ( .A(n31786), .B(n31787), .Z(n31785) );
  XOR U31225 ( .A(n31676), .B(n31784), .Z(n31787) );
  XNOR U31226 ( .A(n31788), .B(n31784), .Z(n31786) );
  XOR U31227 ( .A(n31789), .B(n31790), .Z(n31784) );
  AND U31228 ( .A(n31791), .B(n31792), .Z(n31790) );
  XOR U31229 ( .A(n31691), .B(n31789), .Z(n31792) );
  XOR U31230 ( .A(n31789), .B(n31692), .Z(n31791) );
  XOR U31231 ( .A(n31793), .B(n31794), .Z(n31789) );
  AND U31232 ( .A(n31795), .B(n31796), .Z(n31794) );
  XOR U31233 ( .A(n31719), .B(n31793), .Z(n31796) );
  XOR U31234 ( .A(n31793), .B(n31720), .Z(n31795) );
  XOR U31235 ( .A(n31797), .B(n31798), .Z(n31793) );
  AND U31236 ( .A(n31799), .B(n31800), .Z(n31798) );
  XOR U31237 ( .A(n31797), .B(n31770), .Z(n31800) );
  XNOR U31238 ( .A(n31801), .B(n31802), .Z(n31622) );
  AND U31239 ( .A(n307), .B(n31803), .Z(n31802) );
  XNOR U31240 ( .A(n31804), .B(n31805), .Z(n307) );
  AND U31241 ( .A(n31806), .B(n31807), .Z(n31805) );
  XOR U31242 ( .A(n31804), .B(n31632), .Z(n31807) );
  XNOR U31243 ( .A(n31804), .B(n31592), .Z(n31806) );
  XOR U31244 ( .A(n31808), .B(n31809), .Z(n31804) );
  AND U31245 ( .A(n31810), .B(n31811), .Z(n31809) );
  XOR U31246 ( .A(n31808), .B(n31600), .Z(n31810) );
  XOR U31247 ( .A(n31812), .B(n31813), .Z(n31583) );
  AND U31248 ( .A(n311), .B(n31803), .Z(n31813) );
  XNOR U31249 ( .A(n31801), .B(n31812), .Z(n31803) );
  XNOR U31250 ( .A(n31814), .B(n31815), .Z(n311) );
  AND U31251 ( .A(n31816), .B(n31817), .Z(n31815) );
  XNOR U31252 ( .A(n31818), .B(n31814), .Z(n31817) );
  IV U31253 ( .A(n31632), .Z(n31818) );
  XOR U31254 ( .A(n31788), .B(n31819), .Z(n31632) );
  AND U31255 ( .A(n314), .B(n31820), .Z(n31819) );
  XOR U31256 ( .A(n31675), .B(n31672), .Z(n31820) );
  IV U31257 ( .A(n31788), .Z(n31675) );
  XNOR U31258 ( .A(n31592), .B(n31814), .Z(n31816) );
  XOR U31259 ( .A(n31821), .B(n31822), .Z(n31592) );
  AND U31260 ( .A(n330), .B(n31823), .Z(n31822) );
  XOR U31261 ( .A(n31808), .B(n31824), .Z(n31814) );
  AND U31262 ( .A(n31825), .B(n31811), .Z(n31824) );
  XNOR U31263 ( .A(n31642), .B(n31808), .Z(n31811) );
  XOR U31264 ( .A(n31692), .B(n31826), .Z(n31642) );
  AND U31265 ( .A(n314), .B(n31827), .Z(n31826) );
  XOR U31266 ( .A(n31688), .B(n31692), .Z(n31827) );
  XNOR U31267 ( .A(n31828), .B(n31808), .Z(n31825) );
  IV U31268 ( .A(n31600), .Z(n31828) );
  XOR U31269 ( .A(n31829), .B(n31830), .Z(n31600) );
  AND U31270 ( .A(n330), .B(n31831), .Z(n31830) );
  XOR U31271 ( .A(n31832), .B(n31833), .Z(n31808) );
  AND U31272 ( .A(n31834), .B(n31835), .Z(n31833) );
  XNOR U31273 ( .A(n31652), .B(n31832), .Z(n31835) );
  XOR U31274 ( .A(n31720), .B(n31836), .Z(n31652) );
  AND U31275 ( .A(n314), .B(n31837), .Z(n31836) );
  XOR U31276 ( .A(n31716), .B(n31720), .Z(n31837) );
  XOR U31277 ( .A(n31832), .B(n31609), .Z(n31834) );
  XOR U31278 ( .A(n31838), .B(n31839), .Z(n31609) );
  AND U31279 ( .A(n330), .B(n31840), .Z(n31839) );
  XOR U31280 ( .A(n31841), .B(n31842), .Z(n31832) );
  AND U31281 ( .A(n31843), .B(n31844), .Z(n31842) );
  XNOR U31282 ( .A(n31841), .B(n31660), .Z(n31844) );
  XOR U31283 ( .A(n31771), .B(n31845), .Z(n31660) );
  AND U31284 ( .A(n314), .B(n31846), .Z(n31845) );
  XOR U31285 ( .A(n31767), .B(n31771), .Z(n31846) );
  XNOR U31286 ( .A(n31847), .B(n31841), .Z(n31843) );
  IV U31287 ( .A(n31619), .Z(n31847) );
  XOR U31288 ( .A(n31848), .B(n31849), .Z(n31619) );
  AND U31289 ( .A(n330), .B(n31850), .Z(n31849) );
  AND U31290 ( .A(n31812), .B(n31801), .Z(n31841) );
  XNOR U31291 ( .A(n31851), .B(n31852), .Z(n31801) );
  AND U31292 ( .A(n314), .B(n31783), .Z(n31852) );
  XNOR U31293 ( .A(n31781), .B(n31851), .Z(n31783) );
  XNOR U31294 ( .A(n31853), .B(n31854), .Z(n314) );
  AND U31295 ( .A(n31855), .B(n31856), .Z(n31854) );
  XNOR U31296 ( .A(n31853), .B(n31672), .Z(n31856) );
  IV U31297 ( .A(n31676), .Z(n31672) );
  XOR U31298 ( .A(n31857), .B(n31858), .Z(n31676) );
  AND U31299 ( .A(n318), .B(n31859), .Z(n31858) );
  XOR U31300 ( .A(n31860), .B(n31857), .Z(n31859) );
  XNOR U31301 ( .A(n31853), .B(n31788), .Z(n31855) );
  XOR U31302 ( .A(n31861), .B(n31862), .Z(n31788) );
  AND U31303 ( .A(n326), .B(n31823), .Z(n31862) );
  XOR U31304 ( .A(n31821), .B(n31861), .Z(n31823) );
  XOR U31305 ( .A(n31863), .B(n31864), .Z(n31853) );
  AND U31306 ( .A(n31865), .B(n31866), .Z(n31864) );
  XNOR U31307 ( .A(n31863), .B(n31688), .Z(n31866) );
  IV U31308 ( .A(n31691), .Z(n31688) );
  XOR U31309 ( .A(n31867), .B(n31868), .Z(n31691) );
  AND U31310 ( .A(n318), .B(n31869), .Z(n31868) );
  XOR U31311 ( .A(n31870), .B(n31867), .Z(n31869) );
  XOR U31312 ( .A(n31692), .B(n31863), .Z(n31865) );
  XOR U31313 ( .A(n31871), .B(n31872), .Z(n31692) );
  AND U31314 ( .A(n326), .B(n31831), .Z(n31872) );
  XOR U31315 ( .A(n31871), .B(n31829), .Z(n31831) );
  XOR U31316 ( .A(n31873), .B(n31874), .Z(n31863) );
  AND U31317 ( .A(n31875), .B(n31876), .Z(n31874) );
  XNOR U31318 ( .A(n31873), .B(n31716), .Z(n31876) );
  IV U31319 ( .A(n31719), .Z(n31716) );
  XOR U31320 ( .A(n31877), .B(n31878), .Z(n31719) );
  AND U31321 ( .A(n318), .B(n31879), .Z(n31878) );
  XNOR U31322 ( .A(n31880), .B(n31877), .Z(n31879) );
  XOR U31323 ( .A(n31720), .B(n31873), .Z(n31875) );
  XOR U31324 ( .A(n31881), .B(n31882), .Z(n31720) );
  AND U31325 ( .A(n326), .B(n31840), .Z(n31882) );
  XOR U31326 ( .A(n31881), .B(n31838), .Z(n31840) );
  XOR U31327 ( .A(n31797), .B(n31883), .Z(n31873) );
  AND U31328 ( .A(n31799), .B(n31884), .Z(n31883) );
  XNOR U31329 ( .A(n31797), .B(n31767), .Z(n31884) );
  IV U31330 ( .A(n31770), .Z(n31767) );
  XOR U31331 ( .A(n31885), .B(n31886), .Z(n31770) );
  AND U31332 ( .A(n318), .B(n31887), .Z(n31886) );
  XOR U31333 ( .A(n31888), .B(n31885), .Z(n31887) );
  XOR U31334 ( .A(n31771), .B(n31797), .Z(n31799) );
  XOR U31335 ( .A(n31889), .B(n31890), .Z(n31771) );
  AND U31336 ( .A(n326), .B(n31850), .Z(n31890) );
  XOR U31337 ( .A(n31889), .B(n31848), .Z(n31850) );
  AND U31338 ( .A(n31851), .B(n31781), .Z(n31797) );
  XNOR U31339 ( .A(n31891), .B(n31892), .Z(n31781) );
  AND U31340 ( .A(n318), .B(n31893), .Z(n31892) );
  XNOR U31341 ( .A(n31894), .B(n31891), .Z(n31893) );
  XNOR U31342 ( .A(n31895), .B(n31896), .Z(n318) );
  AND U31343 ( .A(n31897), .B(n31898), .Z(n31896) );
  XOR U31344 ( .A(n31860), .B(n31895), .Z(n31898) );
  AND U31345 ( .A(n31899), .B(n31900), .Z(n31860) );
  XNOR U31346 ( .A(n31857), .B(n31895), .Z(n31897) );
  XNOR U31347 ( .A(n31901), .B(n31902), .Z(n31857) );
  AND U31348 ( .A(n322), .B(n31903), .Z(n31902) );
  XNOR U31349 ( .A(n31904), .B(n31905), .Z(n31903) );
  XOR U31350 ( .A(n31906), .B(n31907), .Z(n31895) );
  AND U31351 ( .A(n31908), .B(n31909), .Z(n31907) );
  XNOR U31352 ( .A(n31906), .B(n31899), .Z(n31909) );
  IV U31353 ( .A(n31870), .Z(n31899) );
  XOR U31354 ( .A(n31910), .B(n31911), .Z(n31870) );
  XOR U31355 ( .A(n31912), .B(n31900), .Z(n31911) );
  AND U31356 ( .A(n31880), .B(n31913), .Z(n31900) );
  AND U31357 ( .A(n31914), .B(n31915), .Z(n31912) );
  XOR U31358 ( .A(n31916), .B(n31910), .Z(n31914) );
  XNOR U31359 ( .A(n31867), .B(n31906), .Z(n31908) );
  XNOR U31360 ( .A(n31917), .B(n31918), .Z(n31867) );
  AND U31361 ( .A(n322), .B(n31919), .Z(n31918) );
  XNOR U31362 ( .A(n31920), .B(n31921), .Z(n31919) );
  XOR U31363 ( .A(n31922), .B(n31923), .Z(n31906) );
  AND U31364 ( .A(n31924), .B(n31925), .Z(n31923) );
  XNOR U31365 ( .A(n31922), .B(n31880), .Z(n31925) );
  XOR U31366 ( .A(n31926), .B(n31915), .Z(n31880) );
  XNOR U31367 ( .A(n31927), .B(n31910), .Z(n31915) );
  XOR U31368 ( .A(n31928), .B(n31929), .Z(n31910) );
  AND U31369 ( .A(n31930), .B(n31931), .Z(n31929) );
  XOR U31370 ( .A(n31932), .B(n31928), .Z(n31930) );
  XNOR U31371 ( .A(n31933), .B(n31934), .Z(n31927) );
  AND U31372 ( .A(n31935), .B(n31936), .Z(n31934) );
  XOR U31373 ( .A(n31933), .B(n31937), .Z(n31935) );
  XNOR U31374 ( .A(n31916), .B(n31913), .Z(n31926) );
  AND U31375 ( .A(n31938), .B(n31939), .Z(n31913) );
  XOR U31376 ( .A(n31940), .B(n31941), .Z(n31916) );
  AND U31377 ( .A(n31942), .B(n31943), .Z(n31941) );
  XOR U31378 ( .A(n31940), .B(n31944), .Z(n31942) );
  XNOR U31379 ( .A(n31877), .B(n31922), .Z(n31924) );
  XNOR U31380 ( .A(n31945), .B(n31946), .Z(n31877) );
  AND U31381 ( .A(n322), .B(n31947), .Z(n31946) );
  XNOR U31382 ( .A(n31948), .B(n31949), .Z(n31947) );
  XOR U31383 ( .A(n31950), .B(n31951), .Z(n31922) );
  AND U31384 ( .A(n31952), .B(n31953), .Z(n31951) );
  XNOR U31385 ( .A(n31950), .B(n31938), .Z(n31953) );
  IV U31386 ( .A(n31888), .Z(n31938) );
  XNOR U31387 ( .A(n31954), .B(n31931), .Z(n31888) );
  XNOR U31388 ( .A(n31955), .B(n31937), .Z(n31931) );
  XOR U31389 ( .A(n31956), .B(n31957), .Z(n31937) );
  NOR U31390 ( .A(n31958), .B(n31959), .Z(n31957) );
  XNOR U31391 ( .A(n31956), .B(n31960), .Z(n31958) );
  XNOR U31392 ( .A(n31936), .B(n31928), .Z(n31955) );
  XOR U31393 ( .A(n31961), .B(n31962), .Z(n31928) );
  AND U31394 ( .A(n31963), .B(n31964), .Z(n31962) );
  XNOR U31395 ( .A(n31961), .B(n31965), .Z(n31963) );
  XNOR U31396 ( .A(n31966), .B(n31933), .Z(n31936) );
  XOR U31397 ( .A(n31967), .B(n31968), .Z(n31933) );
  AND U31398 ( .A(n31969), .B(n31970), .Z(n31968) );
  XOR U31399 ( .A(n31967), .B(n31971), .Z(n31969) );
  XNOR U31400 ( .A(n31972), .B(n31973), .Z(n31966) );
  NOR U31401 ( .A(n31974), .B(n31975), .Z(n31973) );
  XOR U31402 ( .A(n31972), .B(n31976), .Z(n31974) );
  XNOR U31403 ( .A(n31932), .B(n31939), .Z(n31954) );
  NOR U31404 ( .A(n31894), .B(n31977), .Z(n31939) );
  XOR U31405 ( .A(n31944), .B(n31943), .Z(n31932) );
  XNOR U31406 ( .A(n31978), .B(n31940), .Z(n31943) );
  XOR U31407 ( .A(n31979), .B(n31980), .Z(n31940) );
  AND U31408 ( .A(n31981), .B(n31982), .Z(n31980) );
  XOR U31409 ( .A(n31979), .B(n31983), .Z(n31981) );
  XNOR U31410 ( .A(n31984), .B(n31985), .Z(n31978) );
  NOR U31411 ( .A(n31986), .B(n31987), .Z(n31985) );
  XNOR U31412 ( .A(n31984), .B(n31988), .Z(n31986) );
  XOR U31413 ( .A(n31989), .B(n31990), .Z(n31944) );
  NOR U31414 ( .A(n31991), .B(n31992), .Z(n31990) );
  XNOR U31415 ( .A(n31989), .B(n31993), .Z(n31991) );
  XNOR U31416 ( .A(n31885), .B(n31950), .Z(n31952) );
  XNOR U31417 ( .A(n31994), .B(n31995), .Z(n31885) );
  AND U31418 ( .A(n322), .B(n31996), .Z(n31995) );
  XNOR U31419 ( .A(n31997), .B(n31998), .Z(n31996) );
  AND U31420 ( .A(n31891), .B(n31894), .Z(n31950) );
  XOR U31421 ( .A(n31999), .B(n31977), .Z(n31894) );
  XNOR U31422 ( .A(p_input[2048]), .B(p_input[208]), .Z(n31977) );
  XOR U31423 ( .A(n31965), .B(n31964), .Z(n31999) );
  XNOR U31424 ( .A(n32000), .B(n31971), .Z(n31964) );
  XNOR U31425 ( .A(n31960), .B(n31959), .Z(n31971) );
  XOR U31426 ( .A(n32001), .B(n31956), .Z(n31959) );
  XNOR U31427 ( .A(n29266), .B(p_input[218]), .Z(n31956) );
  XNOR U31428 ( .A(p_input[2059]), .B(p_input[219]), .Z(n32001) );
  XOR U31429 ( .A(p_input[2060]), .B(p_input[220]), .Z(n31960) );
  XNOR U31430 ( .A(n31970), .B(n31961), .Z(n32000) );
  XNOR U31431 ( .A(n29494), .B(p_input[209]), .Z(n31961) );
  XOR U31432 ( .A(n32002), .B(n31976), .Z(n31970) );
  XNOR U31433 ( .A(p_input[2063]), .B(p_input[223]), .Z(n31976) );
  XOR U31434 ( .A(n31967), .B(n31975), .Z(n32002) );
  XOR U31435 ( .A(n32003), .B(n31972), .Z(n31975) );
  XOR U31436 ( .A(p_input[2061]), .B(p_input[221]), .Z(n31972) );
  XNOR U31437 ( .A(p_input[2062]), .B(p_input[222]), .Z(n32003) );
  XNOR U31438 ( .A(n29036), .B(p_input[217]), .Z(n31967) );
  XNOR U31439 ( .A(n31983), .B(n31982), .Z(n31965) );
  XNOR U31440 ( .A(n32004), .B(n31988), .Z(n31982) );
  XOR U31441 ( .A(p_input[2056]), .B(p_input[216]), .Z(n31988) );
  XOR U31442 ( .A(n31979), .B(n31987), .Z(n32004) );
  XOR U31443 ( .A(n32005), .B(n31984), .Z(n31987) );
  XOR U31444 ( .A(p_input[2054]), .B(p_input[214]), .Z(n31984) );
  XNOR U31445 ( .A(p_input[2055]), .B(p_input[215]), .Z(n32005) );
  XNOR U31446 ( .A(n29039), .B(p_input[210]), .Z(n31979) );
  XNOR U31447 ( .A(n31993), .B(n31992), .Z(n31983) );
  XOR U31448 ( .A(n32006), .B(n31989), .Z(n31992) );
  XOR U31449 ( .A(p_input[2051]), .B(p_input[211]), .Z(n31989) );
  XNOR U31450 ( .A(p_input[2052]), .B(p_input[212]), .Z(n32006) );
  XOR U31451 ( .A(p_input[2053]), .B(p_input[213]), .Z(n31993) );
  XNOR U31452 ( .A(n32007), .B(n32008), .Z(n31891) );
  AND U31453 ( .A(n322), .B(n32009), .Z(n32008) );
  XNOR U31454 ( .A(n32010), .B(n32011), .Z(n322) );
  AND U31455 ( .A(n32012), .B(n32013), .Z(n32011) );
  XOR U31456 ( .A(n31905), .B(n32010), .Z(n32013) );
  XNOR U31457 ( .A(n32014), .B(n32010), .Z(n32012) );
  XOR U31458 ( .A(n32015), .B(n32016), .Z(n32010) );
  AND U31459 ( .A(n32017), .B(n32018), .Z(n32016) );
  XOR U31460 ( .A(n31920), .B(n32015), .Z(n32018) );
  XOR U31461 ( .A(n32015), .B(n31921), .Z(n32017) );
  XOR U31462 ( .A(n32019), .B(n32020), .Z(n32015) );
  AND U31463 ( .A(n32021), .B(n32022), .Z(n32020) );
  XOR U31464 ( .A(n31948), .B(n32019), .Z(n32022) );
  XOR U31465 ( .A(n32019), .B(n31949), .Z(n32021) );
  XOR U31466 ( .A(n32023), .B(n32024), .Z(n32019) );
  AND U31467 ( .A(n32025), .B(n32026), .Z(n32024) );
  XOR U31468 ( .A(n32023), .B(n31997), .Z(n32026) );
  XNOR U31469 ( .A(n32027), .B(n32028), .Z(n31851) );
  AND U31470 ( .A(n326), .B(n32029), .Z(n32028) );
  XNOR U31471 ( .A(n32030), .B(n32031), .Z(n326) );
  AND U31472 ( .A(n32032), .B(n32033), .Z(n32031) );
  XOR U31473 ( .A(n32030), .B(n31861), .Z(n32033) );
  XNOR U31474 ( .A(n32030), .B(n31821), .Z(n32032) );
  XOR U31475 ( .A(n32034), .B(n32035), .Z(n32030) );
  AND U31476 ( .A(n32036), .B(n32037), .Z(n32035) );
  XOR U31477 ( .A(n32034), .B(n31829), .Z(n32036) );
  XOR U31478 ( .A(n32038), .B(n32039), .Z(n31812) );
  AND U31479 ( .A(n330), .B(n32029), .Z(n32039) );
  XNOR U31480 ( .A(n32027), .B(n32038), .Z(n32029) );
  XNOR U31481 ( .A(n32040), .B(n32041), .Z(n330) );
  AND U31482 ( .A(n32042), .B(n32043), .Z(n32041) );
  XNOR U31483 ( .A(n32044), .B(n32040), .Z(n32043) );
  IV U31484 ( .A(n31861), .Z(n32044) );
  XOR U31485 ( .A(n32014), .B(n32045), .Z(n31861) );
  AND U31486 ( .A(n333), .B(n32046), .Z(n32045) );
  XOR U31487 ( .A(n31904), .B(n31901), .Z(n32046) );
  IV U31488 ( .A(n32014), .Z(n31904) );
  XNOR U31489 ( .A(n31821), .B(n32040), .Z(n32042) );
  XOR U31490 ( .A(n32047), .B(n32048), .Z(n31821) );
  AND U31491 ( .A(n349), .B(n32049), .Z(n32048) );
  XOR U31492 ( .A(n32034), .B(n32050), .Z(n32040) );
  AND U31493 ( .A(n32051), .B(n32037), .Z(n32050) );
  XNOR U31494 ( .A(n31871), .B(n32034), .Z(n32037) );
  XOR U31495 ( .A(n31921), .B(n32052), .Z(n31871) );
  AND U31496 ( .A(n333), .B(n32053), .Z(n32052) );
  XOR U31497 ( .A(n31917), .B(n31921), .Z(n32053) );
  XNOR U31498 ( .A(n32054), .B(n32034), .Z(n32051) );
  IV U31499 ( .A(n31829), .Z(n32054) );
  XOR U31500 ( .A(n32055), .B(n32056), .Z(n31829) );
  AND U31501 ( .A(n349), .B(n32057), .Z(n32056) );
  XOR U31502 ( .A(n32058), .B(n32059), .Z(n32034) );
  AND U31503 ( .A(n32060), .B(n32061), .Z(n32059) );
  XNOR U31504 ( .A(n31881), .B(n32058), .Z(n32061) );
  XOR U31505 ( .A(n31949), .B(n32062), .Z(n31881) );
  AND U31506 ( .A(n333), .B(n32063), .Z(n32062) );
  XOR U31507 ( .A(n31945), .B(n31949), .Z(n32063) );
  XOR U31508 ( .A(n32058), .B(n31838), .Z(n32060) );
  XOR U31509 ( .A(n32064), .B(n32065), .Z(n31838) );
  AND U31510 ( .A(n349), .B(n32066), .Z(n32065) );
  XOR U31511 ( .A(n32067), .B(n32068), .Z(n32058) );
  AND U31512 ( .A(n32069), .B(n32070), .Z(n32068) );
  XNOR U31513 ( .A(n32067), .B(n31889), .Z(n32070) );
  XOR U31514 ( .A(n31998), .B(n32071), .Z(n31889) );
  AND U31515 ( .A(n333), .B(n32072), .Z(n32071) );
  XOR U31516 ( .A(n31994), .B(n31998), .Z(n32072) );
  XNOR U31517 ( .A(n32073), .B(n32067), .Z(n32069) );
  IV U31518 ( .A(n31848), .Z(n32073) );
  XOR U31519 ( .A(n32074), .B(n32075), .Z(n31848) );
  AND U31520 ( .A(n349), .B(n32076), .Z(n32075) );
  AND U31521 ( .A(n32038), .B(n32027), .Z(n32067) );
  XNOR U31522 ( .A(n32077), .B(n32078), .Z(n32027) );
  AND U31523 ( .A(n333), .B(n32009), .Z(n32078) );
  XNOR U31524 ( .A(n32007), .B(n32077), .Z(n32009) );
  XNOR U31525 ( .A(n32079), .B(n32080), .Z(n333) );
  AND U31526 ( .A(n32081), .B(n32082), .Z(n32080) );
  XNOR U31527 ( .A(n32079), .B(n31901), .Z(n32082) );
  IV U31528 ( .A(n31905), .Z(n31901) );
  XOR U31529 ( .A(n32083), .B(n32084), .Z(n31905) );
  AND U31530 ( .A(n337), .B(n32085), .Z(n32084) );
  XOR U31531 ( .A(n32086), .B(n32083), .Z(n32085) );
  XNOR U31532 ( .A(n32079), .B(n32014), .Z(n32081) );
  XOR U31533 ( .A(n32087), .B(n32088), .Z(n32014) );
  AND U31534 ( .A(n345), .B(n32049), .Z(n32088) );
  XOR U31535 ( .A(n32047), .B(n32087), .Z(n32049) );
  XOR U31536 ( .A(n32089), .B(n32090), .Z(n32079) );
  AND U31537 ( .A(n32091), .B(n32092), .Z(n32090) );
  XNOR U31538 ( .A(n32089), .B(n31917), .Z(n32092) );
  IV U31539 ( .A(n31920), .Z(n31917) );
  XOR U31540 ( .A(n32093), .B(n32094), .Z(n31920) );
  AND U31541 ( .A(n337), .B(n32095), .Z(n32094) );
  XOR U31542 ( .A(n32096), .B(n32093), .Z(n32095) );
  XOR U31543 ( .A(n31921), .B(n32089), .Z(n32091) );
  XOR U31544 ( .A(n32097), .B(n32098), .Z(n31921) );
  AND U31545 ( .A(n345), .B(n32057), .Z(n32098) );
  XOR U31546 ( .A(n32097), .B(n32055), .Z(n32057) );
  XOR U31547 ( .A(n32099), .B(n32100), .Z(n32089) );
  AND U31548 ( .A(n32101), .B(n32102), .Z(n32100) );
  XNOR U31549 ( .A(n32099), .B(n31945), .Z(n32102) );
  IV U31550 ( .A(n31948), .Z(n31945) );
  XOR U31551 ( .A(n32103), .B(n32104), .Z(n31948) );
  AND U31552 ( .A(n337), .B(n32105), .Z(n32104) );
  XNOR U31553 ( .A(n32106), .B(n32103), .Z(n32105) );
  XOR U31554 ( .A(n31949), .B(n32099), .Z(n32101) );
  XOR U31555 ( .A(n32107), .B(n32108), .Z(n31949) );
  AND U31556 ( .A(n345), .B(n32066), .Z(n32108) );
  XOR U31557 ( .A(n32107), .B(n32064), .Z(n32066) );
  XOR U31558 ( .A(n32023), .B(n32109), .Z(n32099) );
  AND U31559 ( .A(n32025), .B(n32110), .Z(n32109) );
  XNOR U31560 ( .A(n32023), .B(n31994), .Z(n32110) );
  IV U31561 ( .A(n31997), .Z(n31994) );
  XOR U31562 ( .A(n32111), .B(n32112), .Z(n31997) );
  AND U31563 ( .A(n337), .B(n32113), .Z(n32112) );
  XOR U31564 ( .A(n32114), .B(n32111), .Z(n32113) );
  XOR U31565 ( .A(n31998), .B(n32023), .Z(n32025) );
  XOR U31566 ( .A(n32115), .B(n32116), .Z(n31998) );
  AND U31567 ( .A(n345), .B(n32076), .Z(n32116) );
  XOR U31568 ( .A(n32115), .B(n32074), .Z(n32076) );
  AND U31569 ( .A(n32077), .B(n32007), .Z(n32023) );
  XNOR U31570 ( .A(n32117), .B(n32118), .Z(n32007) );
  AND U31571 ( .A(n337), .B(n32119), .Z(n32118) );
  XNOR U31572 ( .A(n32120), .B(n32117), .Z(n32119) );
  XNOR U31573 ( .A(n32121), .B(n32122), .Z(n337) );
  AND U31574 ( .A(n32123), .B(n32124), .Z(n32122) );
  XOR U31575 ( .A(n32086), .B(n32121), .Z(n32124) );
  AND U31576 ( .A(n32125), .B(n32126), .Z(n32086) );
  XNOR U31577 ( .A(n32083), .B(n32121), .Z(n32123) );
  XNOR U31578 ( .A(n32127), .B(n32128), .Z(n32083) );
  AND U31579 ( .A(n341), .B(n32129), .Z(n32128) );
  XNOR U31580 ( .A(n32130), .B(n32131), .Z(n32129) );
  XOR U31581 ( .A(n32132), .B(n32133), .Z(n32121) );
  AND U31582 ( .A(n32134), .B(n32135), .Z(n32133) );
  XNOR U31583 ( .A(n32132), .B(n32125), .Z(n32135) );
  IV U31584 ( .A(n32096), .Z(n32125) );
  XOR U31585 ( .A(n32136), .B(n32137), .Z(n32096) );
  XOR U31586 ( .A(n32138), .B(n32126), .Z(n32137) );
  AND U31587 ( .A(n32106), .B(n32139), .Z(n32126) );
  AND U31588 ( .A(n32140), .B(n32141), .Z(n32138) );
  XOR U31589 ( .A(n32142), .B(n32136), .Z(n32140) );
  XNOR U31590 ( .A(n32093), .B(n32132), .Z(n32134) );
  XNOR U31591 ( .A(n32143), .B(n32144), .Z(n32093) );
  AND U31592 ( .A(n341), .B(n32145), .Z(n32144) );
  XNOR U31593 ( .A(n32146), .B(n32147), .Z(n32145) );
  XOR U31594 ( .A(n32148), .B(n32149), .Z(n32132) );
  AND U31595 ( .A(n32150), .B(n32151), .Z(n32149) );
  XNOR U31596 ( .A(n32148), .B(n32106), .Z(n32151) );
  XOR U31597 ( .A(n32152), .B(n32141), .Z(n32106) );
  XNOR U31598 ( .A(n32153), .B(n32136), .Z(n32141) );
  XOR U31599 ( .A(n32154), .B(n32155), .Z(n32136) );
  AND U31600 ( .A(n32156), .B(n32157), .Z(n32155) );
  XOR U31601 ( .A(n32158), .B(n32154), .Z(n32156) );
  XNOR U31602 ( .A(n32159), .B(n32160), .Z(n32153) );
  AND U31603 ( .A(n32161), .B(n32162), .Z(n32160) );
  XOR U31604 ( .A(n32159), .B(n32163), .Z(n32161) );
  XNOR U31605 ( .A(n32142), .B(n32139), .Z(n32152) );
  AND U31606 ( .A(n32164), .B(n32165), .Z(n32139) );
  XOR U31607 ( .A(n32166), .B(n32167), .Z(n32142) );
  AND U31608 ( .A(n32168), .B(n32169), .Z(n32167) );
  XOR U31609 ( .A(n32166), .B(n32170), .Z(n32168) );
  XNOR U31610 ( .A(n32103), .B(n32148), .Z(n32150) );
  XNOR U31611 ( .A(n32171), .B(n32172), .Z(n32103) );
  AND U31612 ( .A(n341), .B(n32173), .Z(n32172) );
  XNOR U31613 ( .A(n32174), .B(n32175), .Z(n32173) );
  XOR U31614 ( .A(n32176), .B(n32177), .Z(n32148) );
  AND U31615 ( .A(n32178), .B(n32179), .Z(n32177) );
  XNOR U31616 ( .A(n32176), .B(n32164), .Z(n32179) );
  IV U31617 ( .A(n32114), .Z(n32164) );
  XNOR U31618 ( .A(n32180), .B(n32157), .Z(n32114) );
  XNOR U31619 ( .A(n32181), .B(n32163), .Z(n32157) );
  XOR U31620 ( .A(n32182), .B(n32183), .Z(n32163) );
  NOR U31621 ( .A(n32184), .B(n32185), .Z(n32183) );
  XNOR U31622 ( .A(n32182), .B(n32186), .Z(n32184) );
  XNOR U31623 ( .A(n32162), .B(n32154), .Z(n32181) );
  XOR U31624 ( .A(n32187), .B(n32188), .Z(n32154) );
  AND U31625 ( .A(n32189), .B(n32190), .Z(n32188) );
  XNOR U31626 ( .A(n32187), .B(n32191), .Z(n32189) );
  XNOR U31627 ( .A(n32192), .B(n32159), .Z(n32162) );
  XOR U31628 ( .A(n32193), .B(n32194), .Z(n32159) );
  AND U31629 ( .A(n32195), .B(n32196), .Z(n32194) );
  XOR U31630 ( .A(n32193), .B(n32197), .Z(n32195) );
  XNOR U31631 ( .A(n32198), .B(n32199), .Z(n32192) );
  NOR U31632 ( .A(n32200), .B(n32201), .Z(n32199) );
  XOR U31633 ( .A(n32198), .B(n32202), .Z(n32200) );
  XNOR U31634 ( .A(n32158), .B(n32165), .Z(n32180) );
  NOR U31635 ( .A(n32120), .B(n32203), .Z(n32165) );
  XOR U31636 ( .A(n32170), .B(n32169), .Z(n32158) );
  XNOR U31637 ( .A(n32204), .B(n32166), .Z(n32169) );
  XOR U31638 ( .A(n32205), .B(n32206), .Z(n32166) );
  AND U31639 ( .A(n32207), .B(n32208), .Z(n32206) );
  XOR U31640 ( .A(n32205), .B(n32209), .Z(n32207) );
  XNOR U31641 ( .A(n32210), .B(n32211), .Z(n32204) );
  NOR U31642 ( .A(n32212), .B(n32213), .Z(n32211) );
  XNOR U31643 ( .A(n32210), .B(n32214), .Z(n32212) );
  XOR U31644 ( .A(n32215), .B(n32216), .Z(n32170) );
  NOR U31645 ( .A(n32217), .B(n32218), .Z(n32216) );
  XNOR U31646 ( .A(n32215), .B(n32219), .Z(n32217) );
  XNOR U31647 ( .A(n32111), .B(n32176), .Z(n32178) );
  XNOR U31648 ( .A(n32220), .B(n32221), .Z(n32111) );
  AND U31649 ( .A(n341), .B(n32222), .Z(n32221) );
  XNOR U31650 ( .A(n32223), .B(n32224), .Z(n32222) );
  AND U31651 ( .A(n32117), .B(n32120), .Z(n32176) );
  XOR U31652 ( .A(n32225), .B(n32203), .Z(n32120) );
  XNOR U31653 ( .A(p_input[2048]), .B(p_input[224]), .Z(n32203) );
  XOR U31654 ( .A(n32191), .B(n32190), .Z(n32225) );
  XNOR U31655 ( .A(n32226), .B(n32197), .Z(n32190) );
  XNOR U31656 ( .A(n32186), .B(n32185), .Z(n32197) );
  XOR U31657 ( .A(n32227), .B(n32182), .Z(n32185) );
  XNOR U31658 ( .A(n29266), .B(p_input[234]), .Z(n32182) );
  XNOR U31659 ( .A(p_input[2059]), .B(p_input[235]), .Z(n32227) );
  XOR U31660 ( .A(p_input[2060]), .B(p_input[236]), .Z(n32186) );
  XNOR U31661 ( .A(n32196), .B(n32187), .Z(n32226) );
  XNOR U31662 ( .A(n29494), .B(p_input[225]), .Z(n32187) );
  XOR U31663 ( .A(n32228), .B(n32202), .Z(n32196) );
  XNOR U31664 ( .A(p_input[2063]), .B(p_input[239]), .Z(n32202) );
  XOR U31665 ( .A(n32193), .B(n32201), .Z(n32228) );
  XOR U31666 ( .A(n32229), .B(n32198), .Z(n32201) );
  XOR U31667 ( .A(p_input[2061]), .B(p_input[237]), .Z(n32198) );
  XNOR U31668 ( .A(p_input[2062]), .B(p_input[238]), .Z(n32229) );
  XNOR U31669 ( .A(n29036), .B(p_input[233]), .Z(n32193) );
  XNOR U31670 ( .A(n32209), .B(n32208), .Z(n32191) );
  XNOR U31671 ( .A(n32230), .B(n32214), .Z(n32208) );
  XOR U31672 ( .A(p_input[2056]), .B(p_input[232]), .Z(n32214) );
  XOR U31673 ( .A(n32205), .B(n32213), .Z(n32230) );
  XOR U31674 ( .A(n32231), .B(n32210), .Z(n32213) );
  XOR U31675 ( .A(p_input[2054]), .B(p_input[230]), .Z(n32210) );
  XNOR U31676 ( .A(p_input[2055]), .B(p_input[231]), .Z(n32231) );
  XNOR U31677 ( .A(n29039), .B(p_input[226]), .Z(n32205) );
  XNOR U31678 ( .A(n32219), .B(n32218), .Z(n32209) );
  XOR U31679 ( .A(n32232), .B(n32215), .Z(n32218) );
  XOR U31680 ( .A(p_input[2051]), .B(p_input[227]), .Z(n32215) );
  XNOR U31681 ( .A(p_input[2052]), .B(p_input[228]), .Z(n32232) );
  XOR U31682 ( .A(p_input[2053]), .B(p_input[229]), .Z(n32219) );
  XNOR U31683 ( .A(n32233), .B(n32234), .Z(n32117) );
  AND U31684 ( .A(n341), .B(n32235), .Z(n32234) );
  XNOR U31685 ( .A(n32236), .B(n32237), .Z(n341) );
  AND U31686 ( .A(n32238), .B(n32239), .Z(n32237) );
  XOR U31687 ( .A(n32131), .B(n32236), .Z(n32239) );
  XNOR U31688 ( .A(n32240), .B(n32236), .Z(n32238) );
  XOR U31689 ( .A(n32241), .B(n32242), .Z(n32236) );
  AND U31690 ( .A(n32243), .B(n32244), .Z(n32242) );
  XOR U31691 ( .A(n32146), .B(n32241), .Z(n32244) );
  XOR U31692 ( .A(n32241), .B(n32147), .Z(n32243) );
  XOR U31693 ( .A(n32245), .B(n32246), .Z(n32241) );
  AND U31694 ( .A(n32247), .B(n32248), .Z(n32246) );
  XOR U31695 ( .A(n32174), .B(n32245), .Z(n32248) );
  XOR U31696 ( .A(n32245), .B(n32175), .Z(n32247) );
  XOR U31697 ( .A(n32249), .B(n32250), .Z(n32245) );
  AND U31698 ( .A(n32251), .B(n32252), .Z(n32250) );
  XOR U31699 ( .A(n32249), .B(n32223), .Z(n32252) );
  XNOR U31700 ( .A(n32253), .B(n32254), .Z(n32077) );
  AND U31701 ( .A(n345), .B(n32255), .Z(n32254) );
  XNOR U31702 ( .A(n32256), .B(n32257), .Z(n345) );
  AND U31703 ( .A(n32258), .B(n32259), .Z(n32257) );
  XOR U31704 ( .A(n32256), .B(n32087), .Z(n32259) );
  XNOR U31705 ( .A(n32256), .B(n32047), .Z(n32258) );
  XOR U31706 ( .A(n32260), .B(n32261), .Z(n32256) );
  AND U31707 ( .A(n32262), .B(n32263), .Z(n32261) );
  XOR U31708 ( .A(n32260), .B(n32055), .Z(n32262) );
  XOR U31709 ( .A(n32264), .B(n32265), .Z(n32038) );
  AND U31710 ( .A(n349), .B(n32255), .Z(n32265) );
  XNOR U31711 ( .A(n32253), .B(n32264), .Z(n32255) );
  XNOR U31712 ( .A(n32266), .B(n32267), .Z(n349) );
  AND U31713 ( .A(n32268), .B(n32269), .Z(n32267) );
  XNOR U31714 ( .A(n32270), .B(n32266), .Z(n32269) );
  IV U31715 ( .A(n32087), .Z(n32270) );
  XOR U31716 ( .A(n32240), .B(n32271), .Z(n32087) );
  AND U31717 ( .A(n352), .B(n32272), .Z(n32271) );
  XOR U31718 ( .A(n32130), .B(n32127), .Z(n32272) );
  IV U31719 ( .A(n32240), .Z(n32130) );
  XNOR U31720 ( .A(n32047), .B(n32266), .Z(n32268) );
  XOR U31721 ( .A(n32273), .B(n32274), .Z(n32047) );
  AND U31722 ( .A(n368), .B(n32275), .Z(n32274) );
  XOR U31723 ( .A(n32260), .B(n32276), .Z(n32266) );
  AND U31724 ( .A(n32277), .B(n32263), .Z(n32276) );
  XNOR U31725 ( .A(n32097), .B(n32260), .Z(n32263) );
  XOR U31726 ( .A(n32147), .B(n32278), .Z(n32097) );
  AND U31727 ( .A(n352), .B(n32279), .Z(n32278) );
  XOR U31728 ( .A(n32143), .B(n32147), .Z(n32279) );
  XNOR U31729 ( .A(n32280), .B(n32260), .Z(n32277) );
  IV U31730 ( .A(n32055), .Z(n32280) );
  XOR U31731 ( .A(n32281), .B(n32282), .Z(n32055) );
  AND U31732 ( .A(n368), .B(n32283), .Z(n32282) );
  XOR U31733 ( .A(n32284), .B(n32285), .Z(n32260) );
  AND U31734 ( .A(n32286), .B(n32287), .Z(n32285) );
  XNOR U31735 ( .A(n32107), .B(n32284), .Z(n32287) );
  XOR U31736 ( .A(n32175), .B(n32288), .Z(n32107) );
  AND U31737 ( .A(n352), .B(n32289), .Z(n32288) );
  XOR U31738 ( .A(n32171), .B(n32175), .Z(n32289) );
  XOR U31739 ( .A(n32284), .B(n32064), .Z(n32286) );
  XOR U31740 ( .A(n32290), .B(n32291), .Z(n32064) );
  AND U31741 ( .A(n368), .B(n32292), .Z(n32291) );
  XOR U31742 ( .A(n32293), .B(n32294), .Z(n32284) );
  AND U31743 ( .A(n32295), .B(n32296), .Z(n32294) );
  XNOR U31744 ( .A(n32293), .B(n32115), .Z(n32296) );
  XOR U31745 ( .A(n32224), .B(n32297), .Z(n32115) );
  AND U31746 ( .A(n352), .B(n32298), .Z(n32297) );
  XOR U31747 ( .A(n32220), .B(n32224), .Z(n32298) );
  XNOR U31748 ( .A(n32299), .B(n32293), .Z(n32295) );
  IV U31749 ( .A(n32074), .Z(n32299) );
  XOR U31750 ( .A(n32300), .B(n32301), .Z(n32074) );
  AND U31751 ( .A(n368), .B(n32302), .Z(n32301) );
  AND U31752 ( .A(n32264), .B(n32253), .Z(n32293) );
  XNOR U31753 ( .A(n32303), .B(n32304), .Z(n32253) );
  AND U31754 ( .A(n352), .B(n32235), .Z(n32304) );
  XNOR U31755 ( .A(n32233), .B(n32303), .Z(n32235) );
  XNOR U31756 ( .A(n32305), .B(n32306), .Z(n352) );
  AND U31757 ( .A(n32307), .B(n32308), .Z(n32306) );
  XNOR U31758 ( .A(n32305), .B(n32127), .Z(n32308) );
  IV U31759 ( .A(n32131), .Z(n32127) );
  XOR U31760 ( .A(n32309), .B(n32310), .Z(n32131) );
  AND U31761 ( .A(n356), .B(n32311), .Z(n32310) );
  XOR U31762 ( .A(n32312), .B(n32309), .Z(n32311) );
  XNOR U31763 ( .A(n32305), .B(n32240), .Z(n32307) );
  XOR U31764 ( .A(n32313), .B(n32314), .Z(n32240) );
  AND U31765 ( .A(n364), .B(n32275), .Z(n32314) );
  XOR U31766 ( .A(n32273), .B(n32313), .Z(n32275) );
  XOR U31767 ( .A(n32315), .B(n32316), .Z(n32305) );
  AND U31768 ( .A(n32317), .B(n32318), .Z(n32316) );
  XNOR U31769 ( .A(n32315), .B(n32143), .Z(n32318) );
  IV U31770 ( .A(n32146), .Z(n32143) );
  XOR U31771 ( .A(n32319), .B(n32320), .Z(n32146) );
  AND U31772 ( .A(n356), .B(n32321), .Z(n32320) );
  XOR U31773 ( .A(n32322), .B(n32319), .Z(n32321) );
  XOR U31774 ( .A(n32147), .B(n32315), .Z(n32317) );
  XOR U31775 ( .A(n32323), .B(n32324), .Z(n32147) );
  AND U31776 ( .A(n364), .B(n32283), .Z(n32324) );
  XOR U31777 ( .A(n32323), .B(n32281), .Z(n32283) );
  XOR U31778 ( .A(n32325), .B(n32326), .Z(n32315) );
  AND U31779 ( .A(n32327), .B(n32328), .Z(n32326) );
  XNOR U31780 ( .A(n32325), .B(n32171), .Z(n32328) );
  IV U31781 ( .A(n32174), .Z(n32171) );
  XOR U31782 ( .A(n32329), .B(n32330), .Z(n32174) );
  AND U31783 ( .A(n356), .B(n32331), .Z(n32330) );
  XNOR U31784 ( .A(n32332), .B(n32329), .Z(n32331) );
  XOR U31785 ( .A(n32175), .B(n32325), .Z(n32327) );
  XOR U31786 ( .A(n32333), .B(n32334), .Z(n32175) );
  AND U31787 ( .A(n364), .B(n32292), .Z(n32334) );
  XOR U31788 ( .A(n32333), .B(n32290), .Z(n32292) );
  XOR U31789 ( .A(n32249), .B(n32335), .Z(n32325) );
  AND U31790 ( .A(n32251), .B(n32336), .Z(n32335) );
  XNOR U31791 ( .A(n32249), .B(n32220), .Z(n32336) );
  IV U31792 ( .A(n32223), .Z(n32220) );
  XOR U31793 ( .A(n32337), .B(n32338), .Z(n32223) );
  AND U31794 ( .A(n356), .B(n32339), .Z(n32338) );
  XOR U31795 ( .A(n32340), .B(n32337), .Z(n32339) );
  XOR U31796 ( .A(n32224), .B(n32249), .Z(n32251) );
  XOR U31797 ( .A(n32341), .B(n32342), .Z(n32224) );
  AND U31798 ( .A(n364), .B(n32302), .Z(n32342) );
  XOR U31799 ( .A(n32341), .B(n32300), .Z(n32302) );
  AND U31800 ( .A(n32303), .B(n32233), .Z(n32249) );
  XNOR U31801 ( .A(n32343), .B(n32344), .Z(n32233) );
  AND U31802 ( .A(n356), .B(n32345), .Z(n32344) );
  XNOR U31803 ( .A(n32346), .B(n32343), .Z(n32345) );
  XNOR U31804 ( .A(n32347), .B(n32348), .Z(n356) );
  AND U31805 ( .A(n32349), .B(n32350), .Z(n32348) );
  XOR U31806 ( .A(n32312), .B(n32347), .Z(n32350) );
  AND U31807 ( .A(n32351), .B(n32352), .Z(n32312) );
  XNOR U31808 ( .A(n32309), .B(n32347), .Z(n32349) );
  XNOR U31809 ( .A(n32353), .B(n32354), .Z(n32309) );
  AND U31810 ( .A(n360), .B(n32355), .Z(n32354) );
  XNOR U31811 ( .A(n32356), .B(n32357), .Z(n32355) );
  XOR U31812 ( .A(n32358), .B(n32359), .Z(n32347) );
  AND U31813 ( .A(n32360), .B(n32361), .Z(n32359) );
  XNOR U31814 ( .A(n32358), .B(n32351), .Z(n32361) );
  IV U31815 ( .A(n32322), .Z(n32351) );
  XOR U31816 ( .A(n32362), .B(n32363), .Z(n32322) );
  XOR U31817 ( .A(n32364), .B(n32352), .Z(n32363) );
  AND U31818 ( .A(n32332), .B(n32365), .Z(n32352) );
  AND U31819 ( .A(n32366), .B(n32367), .Z(n32364) );
  XOR U31820 ( .A(n32368), .B(n32362), .Z(n32366) );
  XNOR U31821 ( .A(n32319), .B(n32358), .Z(n32360) );
  XNOR U31822 ( .A(n32369), .B(n32370), .Z(n32319) );
  AND U31823 ( .A(n360), .B(n32371), .Z(n32370) );
  XNOR U31824 ( .A(n32372), .B(n32373), .Z(n32371) );
  XOR U31825 ( .A(n32374), .B(n32375), .Z(n32358) );
  AND U31826 ( .A(n32376), .B(n32377), .Z(n32375) );
  XNOR U31827 ( .A(n32374), .B(n32332), .Z(n32377) );
  XOR U31828 ( .A(n32378), .B(n32367), .Z(n32332) );
  XNOR U31829 ( .A(n32379), .B(n32362), .Z(n32367) );
  XOR U31830 ( .A(n32380), .B(n32381), .Z(n32362) );
  AND U31831 ( .A(n32382), .B(n32383), .Z(n32381) );
  XOR U31832 ( .A(n32384), .B(n32380), .Z(n32382) );
  XNOR U31833 ( .A(n32385), .B(n32386), .Z(n32379) );
  AND U31834 ( .A(n32387), .B(n32388), .Z(n32386) );
  XOR U31835 ( .A(n32385), .B(n32389), .Z(n32387) );
  XNOR U31836 ( .A(n32368), .B(n32365), .Z(n32378) );
  AND U31837 ( .A(n32390), .B(n32391), .Z(n32365) );
  XOR U31838 ( .A(n32392), .B(n32393), .Z(n32368) );
  AND U31839 ( .A(n32394), .B(n32395), .Z(n32393) );
  XOR U31840 ( .A(n32392), .B(n32396), .Z(n32394) );
  XNOR U31841 ( .A(n32329), .B(n32374), .Z(n32376) );
  XNOR U31842 ( .A(n32397), .B(n32398), .Z(n32329) );
  AND U31843 ( .A(n360), .B(n32399), .Z(n32398) );
  XNOR U31844 ( .A(n32400), .B(n32401), .Z(n32399) );
  XOR U31845 ( .A(n32402), .B(n32403), .Z(n32374) );
  AND U31846 ( .A(n32404), .B(n32405), .Z(n32403) );
  XNOR U31847 ( .A(n32402), .B(n32390), .Z(n32405) );
  IV U31848 ( .A(n32340), .Z(n32390) );
  XNOR U31849 ( .A(n32406), .B(n32383), .Z(n32340) );
  XNOR U31850 ( .A(n32407), .B(n32389), .Z(n32383) );
  XOR U31851 ( .A(n32408), .B(n32409), .Z(n32389) );
  NOR U31852 ( .A(n32410), .B(n32411), .Z(n32409) );
  XNOR U31853 ( .A(n32408), .B(n32412), .Z(n32410) );
  XNOR U31854 ( .A(n32388), .B(n32380), .Z(n32407) );
  XOR U31855 ( .A(n32413), .B(n32414), .Z(n32380) );
  AND U31856 ( .A(n32415), .B(n32416), .Z(n32414) );
  XNOR U31857 ( .A(n32413), .B(n32417), .Z(n32415) );
  XNOR U31858 ( .A(n32418), .B(n32385), .Z(n32388) );
  XOR U31859 ( .A(n32419), .B(n32420), .Z(n32385) );
  AND U31860 ( .A(n32421), .B(n32422), .Z(n32420) );
  XOR U31861 ( .A(n32419), .B(n32423), .Z(n32421) );
  XNOR U31862 ( .A(n32424), .B(n32425), .Z(n32418) );
  NOR U31863 ( .A(n32426), .B(n32427), .Z(n32425) );
  XOR U31864 ( .A(n32424), .B(n32428), .Z(n32426) );
  XNOR U31865 ( .A(n32384), .B(n32391), .Z(n32406) );
  NOR U31866 ( .A(n32346), .B(n32429), .Z(n32391) );
  XOR U31867 ( .A(n32396), .B(n32395), .Z(n32384) );
  XNOR U31868 ( .A(n32430), .B(n32392), .Z(n32395) );
  XOR U31869 ( .A(n32431), .B(n32432), .Z(n32392) );
  AND U31870 ( .A(n32433), .B(n32434), .Z(n32432) );
  XOR U31871 ( .A(n32431), .B(n32435), .Z(n32433) );
  XNOR U31872 ( .A(n32436), .B(n32437), .Z(n32430) );
  NOR U31873 ( .A(n32438), .B(n32439), .Z(n32437) );
  XNOR U31874 ( .A(n32436), .B(n32440), .Z(n32438) );
  XOR U31875 ( .A(n32441), .B(n32442), .Z(n32396) );
  NOR U31876 ( .A(n32443), .B(n32444), .Z(n32442) );
  XNOR U31877 ( .A(n32441), .B(n32445), .Z(n32443) );
  XNOR U31878 ( .A(n32337), .B(n32402), .Z(n32404) );
  XNOR U31879 ( .A(n32446), .B(n32447), .Z(n32337) );
  AND U31880 ( .A(n360), .B(n32448), .Z(n32447) );
  XNOR U31881 ( .A(n32449), .B(n32450), .Z(n32448) );
  AND U31882 ( .A(n32343), .B(n32346), .Z(n32402) );
  XOR U31883 ( .A(n32451), .B(n32429), .Z(n32346) );
  XNOR U31884 ( .A(p_input[2048]), .B(p_input[240]), .Z(n32429) );
  XOR U31885 ( .A(n32417), .B(n32416), .Z(n32451) );
  XNOR U31886 ( .A(n32452), .B(n32423), .Z(n32416) );
  XNOR U31887 ( .A(n32412), .B(n32411), .Z(n32423) );
  XOR U31888 ( .A(n32453), .B(n32408), .Z(n32411) );
  XNOR U31889 ( .A(n29266), .B(p_input[250]), .Z(n32408) );
  XNOR U31890 ( .A(p_input[2059]), .B(p_input[251]), .Z(n32453) );
  XOR U31891 ( .A(p_input[2060]), .B(p_input[252]), .Z(n32412) );
  XNOR U31892 ( .A(n32422), .B(n32413), .Z(n32452) );
  XNOR U31893 ( .A(n29494), .B(p_input[241]), .Z(n32413) );
  XOR U31894 ( .A(n32454), .B(n32428), .Z(n32422) );
  XNOR U31895 ( .A(p_input[2063]), .B(p_input[255]), .Z(n32428) );
  XOR U31896 ( .A(n32419), .B(n32427), .Z(n32454) );
  XOR U31897 ( .A(n32455), .B(n32424), .Z(n32427) );
  XOR U31898 ( .A(p_input[2061]), .B(p_input[253]), .Z(n32424) );
  XNOR U31899 ( .A(p_input[2062]), .B(p_input[254]), .Z(n32455) );
  XNOR U31900 ( .A(n29036), .B(p_input[249]), .Z(n32419) );
  XNOR U31901 ( .A(n32435), .B(n32434), .Z(n32417) );
  XNOR U31902 ( .A(n32456), .B(n32440), .Z(n32434) );
  XOR U31903 ( .A(p_input[2056]), .B(p_input[248]), .Z(n32440) );
  XOR U31904 ( .A(n32431), .B(n32439), .Z(n32456) );
  XOR U31905 ( .A(n32457), .B(n32436), .Z(n32439) );
  XOR U31906 ( .A(p_input[2054]), .B(p_input[246]), .Z(n32436) );
  XNOR U31907 ( .A(p_input[2055]), .B(p_input[247]), .Z(n32457) );
  XNOR U31908 ( .A(n29039), .B(p_input[242]), .Z(n32431) );
  XNOR U31909 ( .A(n32445), .B(n32444), .Z(n32435) );
  XOR U31910 ( .A(n32458), .B(n32441), .Z(n32444) );
  XOR U31911 ( .A(p_input[2051]), .B(p_input[243]), .Z(n32441) );
  XNOR U31912 ( .A(p_input[2052]), .B(p_input[244]), .Z(n32458) );
  XOR U31913 ( .A(p_input[2053]), .B(p_input[245]), .Z(n32445) );
  XNOR U31914 ( .A(n32459), .B(n32460), .Z(n32343) );
  AND U31915 ( .A(n360), .B(n32461), .Z(n32460) );
  XNOR U31916 ( .A(n32462), .B(n32463), .Z(n360) );
  AND U31917 ( .A(n32464), .B(n32465), .Z(n32463) );
  XOR U31918 ( .A(n32357), .B(n32462), .Z(n32465) );
  XNOR U31919 ( .A(n32466), .B(n32462), .Z(n32464) );
  XOR U31920 ( .A(n32467), .B(n32468), .Z(n32462) );
  AND U31921 ( .A(n32469), .B(n32470), .Z(n32468) );
  XOR U31922 ( .A(n32372), .B(n32467), .Z(n32470) );
  XOR U31923 ( .A(n32467), .B(n32373), .Z(n32469) );
  XOR U31924 ( .A(n32471), .B(n32472), .Z(n32467) );
  AND U31925 ( .A(n32473), .B(n32474), .Z(n32472) );
  XOR U31926 ( .A(n32400), .B(n32471), .Z(n32474) );
  XOR U31927 ( .A(n32471), .B(n32401), .Z(n32473) );
  XOR U31928 ( .A(n32475), .B(n32476), .Z(n32471) );
  AND U31929 ( .A(n32477), .B(n32478), .Z(n32476) );
  XOR U31930 ( .A(n32475), .B(n32449), .Z(n32478) );
  XNOR U31931 ( .A(n32479), .B(n32480), .Z(n32303) );
  AND U31932 ( .A(n364), .B(n32481), .Z(n32480) );
  XNOR U31933 ( .A(n32482), .B(n32483), .Z(n364) );
  AND U31934 ( .A(n32484), .B(n32485), .Z(n32483) );
  XOR U31935 ( .A(n32482), .B(n32313), .Z(n32485) );
  XNOR U31936 ( .A(n32482), .B(n32273), .Z(n32484) );
  XOR U31937 ( .A(n32486), .B(n32487), .Z(n32482) );
  AND U31938 ( .A(n32488), .B(n32489), .Z(n32487) );
  XOR U31939 ( .A(n32486), .B(n32281), .Z(n32488) );
  XOR U31940 ( .A(n32490), .B(n32491), .Z(n32264) );
  AND U31941 ( .A(n368), .B(n32481), .Z(n32491) );
  XNOR U31942 ( .A(n32479), .B(n32490), .Z(n32481) );
  XNOR U31943 ( .A(n32492), .B(n32493), .Z(n368) );
  AND U31944 ( .A(n32494), .B(n32495), .Z(n32493) );
  XNOR U31945 ( .A(n32496), .B(n32492), .Z(n32495) );
  IV U31946 ( .A(n32313), .Z(n32496) );
  XOR U31947 ( .A(n32466), .B(n32497), .Z(n32313) );
  AND U31948 ( .A(n371), .B(n32498), .Z(n32497) );
  XOR U31949 ( .A(n32356), .B(n32353), .Z(n32498) );
  IV U31950 ( .A(n32466), .Z(n32356) );
  XNOR U31951 ( .A(n32273), .B(n32492), .Z(n32494) );
  XOR U31952 ( .A(n32499), .B(n32500), .Z(n32273) );
  AND U31953 ( .A(n387), .B(n32501), .Z(n32500) );
  XOR U31954 ( .A(n32486), .B(n32502), .Z(n32492) );
  AND U31955 ( .A(n32503), .B(n32489), .Z(n32502) );
  XNOR U31956 ( .A(n32323), .B(n32486), .Z(n32489) );
  XOR U31957 ( .A(n32373), .B(n32504), .Z(n32323) );
  AND U31958 ( .A(n371), .B(n32505), .Z(n32504) );
  XOR U31959 ( .A(n32369), .B(n32373), .Z(n32505) );
  XNOR U31960 ( .A(n32506), .B(n32486), .Z(n32503) );
  IV U31961 ( .A(n32281), .Z(n32506) );
  XOR U31962 ( .A(n32507), .B(n32508), .Z(n32281) );
  AND U31963 ( .A(n387), .B(n32509), .Z(n32508) );
  XOR U31964 ( .A(n32510), .B(n32511), .Z(n32486) );
  AND U31965 ( .A(n32512), .B(n32513), .Z(n32511) );
  XNOR U31966 ( .A(n32333), .B(n32510), .Z(n32513) );
  XOR U31967 ( .A(n32401), .B(n32514), .Z(n32333) );
  AND U31968 ( .A(n371), .B(n32515), .Z(n32514) );
  XOR U31969 ( .A(n32397), .B(n32401), .Z(n32515) );
  XOR U31970 ( .A(n32510), .B(n32290), .Z(n32512) );
  XOR U31971 ( .A(n32516), .B(n32517), .Z(n32290) );
  AND U31972 ( .A(n387), .B(n32518), .Z(n32517) );
  XOR U31973 ( .A(n32519), .B(n32520), .Z(n32510) );
  AND U31974 ( .A(n32521), .B(n32522), .Z(n32520) );
  XNOR U31975 ( .A(n32519), .B(n32341), .Z(n32522) );
  XOR U31976 ( .A(n32450), .B(n32523), .Z(n32341) );
  AND U31977 ( .A(n371), .B(n32524), .Z(n32523) );
  XOR U31978 ( .A(n32446), .B(n32450), .Z(n32524) );
  XNOR U31979 ( .A(n32525), .B(n32519), .Z(n32521) );
  IV U31980 ( .A(n32300), .Z(n32525) );
  XOR U31981 ( .A(n32526), .B(n32527), .Z(n32300) );
  AND U31982 ( .A(n387), .B(n32528), .Z(n32527) );
  AND U31983 ( .A(n32490), .B(n32479), .Z(n32519) );
  XNOR U31984 ( .A(n32529), .B(n32530), .Z(n32479) );
  AND U31985 ( .A(n371), .B(n32461), .Z(n32530) );
  XNOR U31986 ( .A(n32459), .B(n32529), .Z(n32461) );
  XNOR U31987 ( .A(n32531), .B(n32532), .Z(n371) );
  AND U31988 ( .A(n32533), .B(n32534), .Z(n32532) );
  XNOR U31989 ( .A(n32531), .B(n32353), .Z(n32534) );
  IV U31990 ( .A(n32357), .Z(n32353) );
  XOR U31991 ( .A(n32535), .B(n32536), .Z(n32357) );
  AND U31992 ( .A(n375), .B(n32537), .Z(n32536) );
  XOR U31993 ( .A(n32538), .B(n32535), .Z(n32537) );
  XNOR U31994 ( .A(n32531), .B(n32466), .Z(n32533) );
  XOR U31995 ( .A(n32539), .B(n32540), .Z(n32466) );
  AND U31996 ( .A(n383), .B(n32501), .Z(n32540) );
  XOR U31997 ( .A(n32499), .B(n32539), .Z(n32501) );
  XOR U31998 ( .A(n32541), .B(n32542), .Z(n32531) );
  AND U31999 ( .A(n32543), .B(n32544), .Z(n32542) );
  XNOR U32000 ( .A(n32541), .B(n32369), .Z(n32544) );
  IV U32001 ( .A(n32372), .Z(n32369) );
  XOR U32002 ( .A(n32545), .B(n32546), .Z(n32372) );
  AND U32003 ( .A(n375), .B(n32547), .Z(n32546) );
  XOR U32004 ( .A(n32548), .B(n32545), .Z(n32547) );
  XOR U32005 ( .A(n32373), .B(n32541), .Z(n32543) );
  XOR U32006 ( .A(n32549), .B(n32550), .Z(n32373) );
  AND U32007 ( .A(n383), .B(n32509), .Z(n32550) );
  XOR U32008 ( .A(n32549), .B(n32507), .Z(n32509) );
  XOR U32009 ( .A(n32551), .B(n32552), .Z(n32541) );
  AND U32010 ( .A(n32553), .B(n32554), .Z(n32552) );
  XNOR U32011 ( .A(n32551), .B(n32397), .Z(n32554) );
  IV U32012 ( .A(n32400), .Z(n32397) );
  XOR U32013 ( .A(n32555), .B(n32556), .Z(n32400) );
  AND U32014 ( .A(n375), .B(n32557), .Z(n32556) );
  XNOR U32015 ( .A(n32558), .B(n32555), .Z(n32557) );
  XOR U32016 ( .A(n32401), .B(n32551), .Z(n32553) );
  XOR U32017 ( .A(n32559), .B(n32560), .Z(n32401) );
  AND U32018 ( .A(n383), .B(n32518), .Z(n32560) );
  XOR U32019 ( .A(n32559), .B(n32516), .Z(n32518) );
  XOR U32020 ( .A(n32475), .B(n32561), .Z(n32551) );
  AND U32021 ( .A(n32477), .B(n32562), .Z(n32561) );
  XNOR U32022 ( .A(n32475), .B(n32446), .Z(n32562) );
  IV U32023 ( .A(n32449), .Z(n32446) );
  XOR U32024 ( .A(n32563), .B(n32564), .Z(n32449) );
  AND U32025 ( .A(n375), .B(n32565), .Z(n32564) );
  XOR U32026 ( .A(n32566), .B(n32563), .Z(n32565) );
  XOR U32027 ( .A(n32450), .B(n32475), .Z(n32477) );
  XOR U32028 ( .A(n32567), .B(n32568), .Z(n32450) );
  AND U32029 ( .A(n383), .B(n32528), .Z(n32568) );
  XOR U32030 ( .A(n32567), .B(n32526), .Z(n32528) );
  AND U32031 ( .A(n32529), .B(n32459), .Z(n32475) );
  XNOR U32032 ( .A(n32569), .B(n32570), .Z(n32459) );
  AND U32033 ( .A(n375), .B(n32571), .Z(n32570) );
  XNOR U32034 ( .A(n32572), .B(n32569), .Z(n32571) );
  XNOR U32035 ( .A(n32573), .B(n32574), .Z(n375) );
  AND U32036 ( .A(n32575), .B(n32576), .Z(n32574) );
  XOR U32037 ( .A(n32538), .B(n32573), .Z(n32576) );
  AND U32038 ( .A(n32577), .B(n32578), .Z(n32538) );
  XNOR U32039 ( .A(n32535), .B(n32573), .Z(n32575) );
  XNOR U32040 ( .A(n32579), .B(n32580), .Z(n32535) );
  AND U32041 ( .A(n379), .B(n32581), .Z(n32580) );
  XNOR U32042 ( .A(n32582), .B(n32583), .Z(n32581) );
  XOR U32043 ( .A(n32584), .B(n32585), .Z(n32573) );
  AND U32044 ( .A(n32586), .B(n32587), .Z(n32585) );
  XNOR U32045 ( .A(n32584), .B(n32577), .Z(n32587) );
  IV U32046 ( .A(n32548), .Z(n32577) );
  XOR U32047 ( .A(n32588), .B(n32589), .Z(n32548) );
  XOR U32048 ( .A(n32590), .B(n32578), .Z(n32589) );
  AND U32049 ( .A(n32558), .B(n32591), .Z(n32578) );
  AND U32050 ( .A(n32592), .B(n32593), .Z(n32590) );
  XOR U32051 ( .A(n32594), .B(n32588), .Z(n32592) );
  XNOR U32052 ( .A(n32545), .B(n32584), .Z(n32586) );
  XNOR U32053 ( .A(n32595), .B(n32596), .Z(n32545) );
  AND U32054 ( .A(n379), .B(n32597), .Z(n32596) );
  XNOR U32055 ( .A(n32598), .B(n32599), .Z(n32597) );
  XOR U32056 ( .A(n32600), .B(n32601), .Z(n32584) );
  AND U32057 ( .A(n32602), .B(n32603), .Z(n32601) );
  XNOR U32058 ( .A(n32600), .B(n32558), .Z(n32603) );
  XOR U32059 ( .A(n32604), .B(n32593), .Z(n32558) );
  XNOR U32060 ( .A(n32605), .B(n32588), .Z(n32593) );
  XOR U32061 ( .A(n32606), .B(n32607), .Z(n32588) );
  AND U32062 ( .A(n32608), .B(n32609), .Z(n32607) );
  XOR U32063 ( .A(n32610), .B(n32606), .Z(n32608) );
  XNOR U32064 ( .A(n32611), .B(n32612), .Z(n32605) );
  AND U32065 ( .A(n32613), .B(n32614), .Z(n32612) );
  XOR U32066 ( .A(n32611), .B(n32615), .Z(n32613) );
  XNOR U32067 ( .A(n32594), .B(n32591), .Z(n32604) );
  AND U32068 ( .A(n32616), .B(n32617), .Z(n32591) );
  XOR U32069 ( .A(n32618), .B(n32619), .Z(n32594) );
  AND U32070 ( .A(n32620), .B(n32621), .Z(n32619) );
  XOR U32071 ( .A(n32618), .B(n32622), .Z(n32620) );
  XNOR U32072 ( .A(n32555), .B(n32600), .Z(n32602) );
  XNOR U32073 ( .A(n32623), .B(n32624), .Z(n32555) );
  AND U32074 ( .A(n379), .B(n32625), .Z(n32624) );
  XNOR U32075 ( .A(n32626), .B(n32627), .Z(n32625) );
  XOR U32076 ( .A(n32628), .B(n32629), .Z(n32600) );
  AND U32077 ( .A(n32630), .B(n32631), .Z(n32629) );
  XNOR U32078 ( .A(n32628), .B(n32616), .Z(n32631) );
  IV U32079 ( .A(n32566), .Z(n32616) );
  XNOR U32080 ( .A(n32632), .B(n32609), .Z(n32566) );
  XNOR U32081 ( .A(n32633), .B(n32615), .Z(n32609) );
  XOR U32082 ( .A(n32634), .B(n32635), .Z(n32615) );
  NOR U32083 ( .A(n32636), .B(n32637), .Z(n32635) );
  XNOR U32084 ( .A(n32634), .B(n32638), .Z(n32636) );
  XNOR U32085 ( .A(n32614), .B(n32606), .Z(n32633) );
  XOR U32086 ( .A(n32639), .B(n32640), .Z(n32606) );
  AND U32087 ( .A(n32641), .B(n32642), .Z(n32640) );
  XNOR U32088 ( .A(n32639), .B(n32643), .Z(n32641) );
  XNOR U32089 ( .A(n32644), .B(n32611), .Z(n32614) );
  XOR U32090 ( .A(n32645), .B(n32646), .Z(n32611) );
  AND U32091 ( .A(n32647), .B(n32648), .Z(n32646) );
  XOR U32092 ( .A(n32645), .B(n32649), .Z(n32647) );
  XNOR U32093 ( .A(n32650), .B(n32651), .Z(n32644) );
  NOR U32094 ( .A(n32652), .B(n32653), .Z(n32651) );
  XOR U32095 ( .A(n32650), .B(n32654), .Z(n32652) );
  XNOR U32096 ( .A(n32610), .B(n32617), .Z(n32632) );
  NOR U32097 ( .A(n32572), .B(n32655), .Z(n32617) );
  XOR U32098 ( .A(n32622), .B(n32621), .Z(n32610) );
  XNOR U32099 ( .A(n32656), .B(n32618), .Z(n32621) );
  XOR U32100 ( .A(n32657), .B(n32658), .Z(n32618) );
  AND U32101 ( .A(n32659), .B(n32660), .Z(n32658) );
  XOR U32102 ( .A(n32657), .B(n32661), .Z(n32659) );
  XNOR U32103 ( .A(n32662), .B(n32663), .Z(n32656) );
  NOR U32104 ( .A(n32664), .B(n32665), .Z(n32663) );
  XNOR U32105 ( .A(n32662), .B(n32666), .Z(n32664) );
  XOR U32106 ( .A(n32667), .B(n32668), .Z(n32622) );
  NOR U32107 ( .A(n32669), .B(n32670), .Z(n32668) );
  XNOR U32108 ( .A(n32667), .B(n32671), .Z(n32669) );
  XNOR U32109 ( .A(n32563), .B(n32628), .Z(n32630) );
  XNOR U32110 ( .A(n32672), .B(n32673), .Z(n32563) );
  AND U32111 ( .A(n379), .B(n32674), .Z(n32673) );
  XNOR U32112 ( .A(n32675), .B(n32676), .Z(n32674) );
  AND U32113 ( .A(n32569), .B(n32572), .Z(n32628) );
  XOR U32114 ( .A(n32677), .B(n32655), .Z(n32572) );
  XNOR U32115 ( .A(p_input[2048]), .B(p_input[256]), .Z(n32655) );
  XOR U32116 ( .A(n32643), .B(n32642), .Z(n32677) );
  XNOR U32117 ( .A(n32678), .B(n32649), .Z(n32642) );
  XNOR U32118 ( .A(n32638), .B(n32637), .Z(n32649) );
  XOR U32119 ( .A(n32679), .B(n32634), .Z(n32637) );
  XNOR U32120 ( .A(n29266), .B(p_input[266]), .Z(n32634) );
  XNOR U32121 ( .A(p_input[2059]), .B(p_input[267]), .Z(n32679) );
  XOR U32122 ( .A(p_input[2060]), .B(p_input[268]), .Z(n32638) );
  XNOR U32123 ( .A(n32648), .B(n32639), .Z(n32678) );
  XNOR U32124 ( .A(n29494), .B(p_input[257]), .Z(n32639) );
  XOR U32125 ( .A(n32680), .B(n32654), .Z(n32648) );
  XNOR U32126 ( .A(p_input[2063]), .B(p_input[271]), .Z(n32654) );
  XOR U32127 ( .A(n32645), .B(n32653), .Z(n32680) );
  XOR U32128 ( .A(n32681), .B(n32650), .Z(n32653) );
  XOR U32129 ( .A(p_input[2061]), .B(p_input[269]), .Z(n32650) );
  XNOR U32130 ( .A(p_input[2062]), .B(p_input[270]), .Z(n32681) );
  XNOR U32131 ( .A(n29036), .B(p_input[265]), .Z(n32645) );
  XNOR U32132 ( .A(n32661), .B(n32660), .Z(n32643) );
  XNOR U32133 ( .A(n32682), .B(n32666), .Z(n32660) );
  XOR U32134 ( .A(p_input[2056]), .B(p_input[264]), .Z(n32666) );
  XOR U32135 ( .A(n32657), .B(n32665), .Z(n32682) );
  XOR U32136 ( .A(n32683), .B(n32662), .Z(n32665) );
  XOR U32137 ( .A(p_input[2054]), .B(p_input[262]), .Z(n32662) );
  XNOR U32138 ( .A(p_input[2055]), .B(p_input[263]), .Z(n32683) );
  XNOR U32139 ( .A(n29039), .B(p_input[258]), .Z(n32657) );
  XNOR U32140 ( .A(n32671), .B(n32670), .Z(n32661) );
  XOR U32141 ( .A(n32684), .B(n32667), .Z(n32670) );
  XOR U32142 ( .A(p_input[2051]), .B(p_input[259]), .Z(n32667) );
  XNOR U32143 ( .A(p_input[2052]), .B(p_input[260]), .Z(n32684) );
  XOR U32144 ( .A(p_input[2053]), .B(p_input[261]), .Z(n32671) );
  XNOR U32145 ( .A(n32685), .B(n32686), .Z(n32569) );
  AND U32146 ( .A(n379), .B(n32687), .Z(n32686) );
  XNOR U32147 ( .A(n32688), .B(n32689), .Z(n379) );
  AND U32148 ( .A(n32690), .B(n32691), .Z(n32689) );
  XOR U32149 ( .A(n32583), .B(n32688), .Z(n32691) );
  XNOR U32150 ( .A(n32692), .B(n32688), .Z(n32690) );
  XOR U32151 ( .A(n32693), .B(n32694), .Z(n32688) );
  AND U32152 ( .A(n32695), .B(n32696), .Z(n32694) );
  XOR U32153 ( .A(n32598), .B(n32693), .Z(n32696) );
  XOR U32154 ( .A(n32693), .B(n32599), .Z(n32695) );
  XOR U32155 ( .A(n32697), .B(n32698), .Z(n32693) );
  AND U32156 ( .A(n32699), .B(n32700), .Z(n32698) );
  XOR U32157 ( .A(n32626), .B(n32697), .Z(n32700) );
  XOR U32158 ( .A(n32697), .B(n32627), .Z(n32699) );
  XOR U32159 ( .A(n32701), .B(n32702), .Z(n32697) );
  AND U32160 ( .A(n32703), .B(n32704), .Z(n32702) );
  XOR U32161 ( .A(n32701), .B(n32675), .Z(n32704) );
  XNOR U32162 ( .A(n32705), .B(n32706), .Z(n32529) );
  AND U32163 ( .A(n383), .B(n32707), .Z(n32706) );
  XNOR U32164 ( .A(n32708), .B(n32709), .Z(n383) );
  AND U32165 ( .A(n32710), .B(n32711), .Z(n32709) );
  XOR U32166 ( .A(n32708), .B(n32539), .Z(n32711) );
  XNOR U32167 ( .A(n32708), .B(n32499), .Z(n32710) );
  XOR U32168 ( .A(n32712), .B(n32713), .Z(n32708) );
  AND U32169 ( .A(n32714), .B(n32715), .Z(n32713) );
  XOR U32170 ( .A(n32712), .B(n32507), .Z(n32714) );
  XOR U32171 ( .A(n32716), .B(n32717), .Z(n32490) );
  AND U32172 ( .A(n387), .B(n32707), .Z(n32717) );
  XNOR U32173 ( .A(n32705), .B(n32716), .Z(n32707) );
  XNOR U32174 ( .A(n32718), .B(n32719), .Z(n387) );
  AND U32175 ( .A(n32720), .B(n32721), .Z(n32719) );
  XNOR U32176 ( .A(n32722), .B(n32718), .Z(n32721) );
  IV U32177 ( .A(n32539), .Z(n32722) );
  XOR U32178 ( .A(n32692), .B(n32723), .Z(n32539) );
  AND U32179 ( .A(n390), .B(n32724), .Z(n32723) );
  XOR U32180 ( .A(n32582), .B(n32579), .Z(n32724) );
  IV U32181 ( .A(n32692), .Z(n32582) );
  XNOR U32182 ( .A(n32499), .B(n32718), .Z(n32720) );
  XOR U32183 ( .A(n32725), .B(n32726), .Z(n32499) );
  AND U32184 ( .A(n406), .B(n32727), .Z(n32726) );
  XOR U32185 ( .A(n32712), .B(n32728), .Z(n32718) );
  AND U32186 ( .A(n32729), .B(n32715), .Z(n32728) );
  XNOR U32187 ( .A(n32549), .B(n32712), .Z(n32715) );
  XOR U32188 ( .A(n32599), .B(n32730), .Z(n32549) );
  AND U32189 ( .A(n390), .B(n32731), .Z(n32730) );
  XOR U32190 ( .A(n32595), .B(n32599), .Z(n32731) );
  XNOR U32191 ( .A(n32732), .B(n32712), .Z(n32729) );
  IV U32192 ( .A(n32507), .Z(n32732) );
  XOR U32193 ( .A(n32733), .B(n32734), .Z(n32507) );
  AND U32194 ( .A(n406), .B(n32735), .Z(n32734) );
  XOR U32195 ( .A(n32736), .B(n32737), .Z(n32712) );
  AND U32196 ( .A(n32738), .B(n32739), .Z(n32737) );
  XNOR U32197 ( .A(n32559), .B(n32736), .Z(n32739) );
  XOR U32198 ( .A(n32627), .B(n32740), .Z(n32559) );
  AND U32199 ( .A(n390), .B(n32741), .Z(n32740) );
  XOR U32200 ( .A(n32623), .B(n32627), .Z(n32741) );
  XOR U32201 ( .A(n32736), .B(n32516), .Z(n32738) );
  XOR U32202 ( .A(n32742), .B(n32743), .Z(n32516) );
  AND U32203 ( .A(n406), .B(n32744), .Z(n32743) );
  XOR U32204 ( .A(n32745), .B(n32746), .Z(n32736) );
  AND U32205 ( .A(n32747), .B(n32748), .Z(n32746) );
  XNOR U32206 ( .A(n32745), .B(n32567), .Z(n32748) );
  XOR U32207 ( .A(n32676), .B(n32749), .Z(n32567) );
  AND U32208 ( .A(n390), .B(n32750), .Z(n32749) );
  XOR U32209 ( .A(n32672), .B(n32676), .Z(n32750) );
  XNOR U32210 ( .A(n32751), .B(n32745), .Z(n32747) );
  IV U32211 ( .A(n32526), .Z(n32751) );
  XOR U32212 ( .A(n32752), .B(n32753), .Z(n32526) );
  AND U32213 ( .A(n406), .B(n32754), .Z(n32753) );
  AND U32214 ( .A(n32716), .B(n32705), .Z(n32745) );
  XNOR U32215 ( .A(n32755), .B(n32756), .Z(n32705) );
  AND U32216 ( .A(n390), .B(n32687), .Z(n32756) );
  XNOR U32217 ( .A(n32685), .B(n32755), .Z(n32687) );
  XNOR U32218 ( .A(n32757), .B(n32758), .Z(n390) );
  AND U32219 ( .A(n32759), .B(n32760), .Z(n32758) );
  XNOR U32220 ( .A(n32757), .B(n32579), .Z(n32760) );
  IV U32221 ( .A(n32583), .Z(n32579) );
  XOR U32222 ( .A(n32761), .B(n32762), .Z(n32583) );
  AND U32223 ( .A(n394), .B(n32763), .Z(n32762) );
  XOR U32224 ( .A(n32764), .B(n32761), .Z(n32763) );
  XNOR U32225 ( .A(n32757), .B(n32692), .Z(n32759) );
  XOR U32226 ( .A(n32765), .B(n32766), .Z(n32692) );
  AND U32227 ( .A(n402), .B(n32727), .Z(n32766) );
  XOR U32228 ( .A(n32725), .B(n32765), .Z(n32727) );
  XOR U32229 ( .A(n32767), .B(n32768), .Z(n32757) );
  AND U32230 ( .A(n32769), .B(n32770), .Z(n32768) );
  XNOR U32231 ( .A(n32767), .B(n32595), .Z(n32770) );
  IV U32232 ( .A(n32598), .Z(n32595) );
  XOR U32233 ( .A(n32771), .B(n32772), .Z(n32598) );
  AND U32234 ( .A(n394), .B(n32773), .Z(n32772) );
  XOR U32235 ( .A(n32774), .B(n32771), .Z(n32773) );
  XOR U32236 ( .A(n32599), .B(n32767), .Z(n32769) );
  XOR U32237 ( .A(n32775), .B(n32776), .Z(n32599) );
  AND U32238 ( .A(n402), .B(n32735), .Z(n32776) );
  XOR U32239 ( .A(n32775), .B(n32733), .Z(n32735) );
  XOR U32240 ( .A(n32777), .B(n32778), .Z(n32767) );
  AND U32241 ( .A(n32779), .B(n32780), .Z(n32778) );
  XNOR U32242 ( .A(n32777), .B(n32623), .Z(n32780) );
  IV U32243 ( .A(n32626), .Z(n32623) );
  XOR U32244 ( .A(n32781), .B(n32782), .Z(n32626) );
  AND U32245 ( .A(n394), .B(n32783), .Z(n32782) );
  XNOR U32246 ( .A(n32784), .B(n32781), .Z(n32783) );
  XOR U32247 ( .A(n32627), .B(n32777), .Z(n32779) );
  XOR U32248 ( .A(n32785), .B(n32786), .Z(n32627) );
  AND U32249 ( .A(n402), .B(n32744), .Z(n32786) );
  XOR U32250 ( .A(n32785), .B(n32742), .Z(n32744) );
  XOR U32251 ( .A(n32701), .B(n32787), .Z(n32777) );
  AND U32252 ( .A(n32703), .B(n32788), .Z(n32787) );
  XNOR U32253 ( .A(n32701), .B(n32672), .Z(n32788) );
  IV U32254 ( .A(n32675), .Z(n32672) );
  XOR U32255 ( .A(n32789), .B(n32790), .Z(n32675) );
  AND U32256 ( .A(n394), .B(n32791), .Z(n32790) );
  XOR U32257 ( .A(n32792), .B(n32789), .Z(n32791) );
  XOR U32258 ( .A(n32676), .B(n32701), .Z(n32703) );
  XOR U32259 ( .A(n32793), .B(n32794), .Z(n32676) );
  AND U32260 ( .A(n402), .B(n32754), .Z(n32794) );
  XOR U32261 ( .A(n32793), .B(n32752), .Z(n32754) );
  AND U32262 ( .A(n32755), .B(n32685), .Z(n32701) );
  XNOR U32263 ( .A(n32795), .B(n32796), .Z(n32685) );
  AND U32264 ( .A(n394), .B(n32797), .Z(n32796) );
  XNOR U32265 ( .A(n32798), .B(n32795), .Z(n32797) );
  XNOR U32266 ( .A(n32799), .B(n32800), .Z(n394) );
  AND U32267 ( .A(n32801), .B(n32802), .Z(n32800) );
  XOR U32268 ( .A(n32764), .B(n32799), .Z(n32802) );
  AND U32269 ( .A(n32803), .B(n32804), .Z(n32764) );
  XNOR U32270 ( .A(n32761), .B(n32799), .Z(n32801) );
  XNOR U32271 ( .A(n32805), .B(n32806), .Z(n32761) );
  AND U32272 ( .A(n398), .B(n32807), .Z(n32806) );
  XNOR U32273 ( .A(n32808), .B(n32809), .Z(n32807) );
  XOR U32274 ( .A(n32810), .B(n32811), .Z(n32799) );
  AND U32275 ( .A(n32812), .B(n32813), .Z(n32811) );
  XNOR U32276 ( .A(n32810), .B(n32803), .Z(n32813) );
  IV U32277 ( .A(n32774), .Z(n32803) );
  XOR U32278 ( .A(n32814), .B(n32815), .Z(n32774) );
  XOR U32279 ( .A(n32816), .B(n32804), .Z(n32815) );
  AND U32280 ( .A(n32784), .B(n32817), .Z(n32804) );
  AND U32281 ( .A(n32818), .B(n32819), .Z(n32816) );
  XOR U32282 ( .A(n32820), .B(n32814), .Z(n32818) );
  XNOR U32283 ( .A(n32771), .B(n32810), .Z(n32812) );
  XNOR U32284 ( .A(n32821), .B(n32822), .Z(n32771) );
  AND U32285 ( .A(n398), .B(n32823), .Z(n32822) );
  XNOR U32286 ( .A(n32824), .B(n32825), .Z(n32823) );
  XOR U32287 ( .A(n32826), .B(n32827), .Z(n32810) );
  AND U32288 ( .A(n32828), .B(n32829), .Z(n32827) );
  XNOR U32289 ( .A(n32826), .B(n32784), .Z(n32829) );
  XOR U32290 ( .A(n32830), .B(n32819), .Z(n32784) );
  XNOR U32291 ( .A(n32831), .B(n32814), .Z(n32819) );
  XOR U32292 ( .A(n32832), .B(n32833), .Z(n32814) );
  AND U32293 ( .A(n32834), .B(n32835), .Z(n32833) );
  XOR U32294 ( .A(n32836), .B(n32832), .Z(n32834) );
  XNOR U32295 ( .A(n32837), .B(n32838), .Z(n32831) );
  AND U32296 ( .A(n32839), .B(n32840), .Z(n32838) );
  XOR U32297 ( .A(n32837), .B(n32841), .Z(n32839) );
  XNOR U32298 ( .A(n32820), .B(n32817), .Z(n32830) );
  AND U32299 ( .A(n32842), .B(n32843), .Z(n32817) );
  XOR U32300 ( .A(n32844), .B(n32845), .Z(n32820) );
  AND U32301 ( .A(n32846), .B(n32847), .Z(n32845) );
  XOR U32302 ( .A(n32844), .B(n32848), .Z(n32846) );
  XNOR U32303 ( .A(n32781), .B(n32826), .Z(n32828) );
  XNOR U32304 ( .A(n32849), .B(n32850), .Z(n32781) );
  AND U32305 ( .A(n398), .B(n32851), .Z(n32850) );
  XNOR U32306 ( .A(n32852), .B(n32853), .Z(n32851) );
  XOR U32307 ( .A(n32854), .B(n32855), .Z(n32826) );
  AND U32308 ( .A(n32856), .B(n32857), .Z(n32855) );
  XNOR U32309 ( .A(n32854), .B(n32842), .Z(n32857) );
  IV U32310 ( .A(n32792), .Z(n32842) );
  XNOR U32311 ( .A(n32858), .B(n32835), .Z(n32792) );
  XNOR U32312 ( .A(n32859), .B(n32841), .Z(n32835) );
  XOR U32313 ( .A(n32860), .B(n32861), .Z(n32841) );
  NOR U32314 ( .A(n32862), .B(n32863), .Z(n32861) );
  XNOR U32315 ( .A(n32860), .B(n32864), .Z(n32862) );
  XNOR U32316 ( .A(n32840), .B(n32832), .Z(n32859) );
  XOR U32317 ( .A(n32865), .B(n32866), .Z(n32832) );
  AND U32318 ( .A(n32867), .B(n32868), .Z(n32866) );
  XNOR U32319 ( .A(n32865), .B(n32869), .Z(n32867) );
  XNOR U32320 ( .A(n32870), .B(n32837), .Z(n32840) );
  XOR U32321 ( .A(n32871), .B(n32872), .Z(n32837) );
  AND U32322 ( .A(n32873), .B(n32874), .Z(n32872) );
  XOR U32323 ( .A(n32871), .B(n32875), .Z(n32873) );
  XNOR U32324 ( .A(n32876), .B(n32877), .Z(n32870) );
  NOR U32325 ( .A(n32878), .B(n32879), .Z(n32877) );
  XOR U32326 ( .A(n32876), .B(n32880), .Z(n32878) );
  XNOR U32327 ( .A(n32836), .B(n32843), .Z(n32858) );
  NOR U32328 ( .A(n32798), .B(n32881), .Z(n32843) );
  XOR U32329 ( .A(n32848), .B(n32847), .Z(n32836) );
  XNOR U32330 ( .A(n32882), .B(n32844), .Z(n32847) );
  XOR U32331 ( .A(n32883), .B(n32884), .Z(n32844) );
  AND U32332 ( .A(n32885), .B(n32886), .Z(n32884) );
  XOR U32333 ( .A(n32883), .B(n32887), .Z(n32885) );
  XNOR U32334 ( .A(n32888), .B(n32889), .Z(n32882) );
  NOR U32335 ( .A(n32890), .B(n32891), .Z(n32889) );
  XNOR U32336 ( .A(n32888), .B(n32892), .Z(n32890) );
  XOR U32337 ( .A(n32893), .B(n32894), .Z(n32848) );
  NOR U32338 ( .A(n32895), .B(n32896), .Z(n32894) );
  XNOR U32339 ( .A(n32893), .B(n32897), .Z(n32895) );
  XNOR U32340 ( .A(n32789), .B(n32854), .Z(n32856) );
  XNOR U32341 ( .A(n32898), .B(n32899), .Z(n32789) );
  AND U32342 ( .A(n398), .B(n32900), .Z(n32899) );
  XNOR U32343 ( .A(n32901), .B(n32902), .Z(n32900) );
  AND U32344 ( .A(n32795), .B(n32798), .Z(n32854) );
  XOR U32345 ( .A(n32903), .B(n32881), .Z(n32798) );
  XNOR U32346 ( .A(p_input[2048]), .B(p_input[272]), .Z(n32881) );
  XOR U32347 ( .A(n32869), .B(n32868), .Z(n32903) );
  XNOR U32348 ( .A(n32904), .B(n32875), .Z(n32868) );
  XNOR U32349 ( .A(n32864), .B(n32863), .Z(n32875) );
  XOR U32350 ( .A(n32905), .B(n32860), .Z(n32863) );
  XNOR U32351 ( .A(n29266), .B(p_input[282]), .Z(n32860) );
  XNOR U32352 ( .A(p_input[2059]), .B(p_input[283]), .Z(n32905) );
  XOR U32353 ( .A(p_input[2060]), .B(p_input[284]), .Z(n32864) );
  XNOR U32354 ( .A(n32874), .B(n32865), .Z(n32904) );
  XNOR U32355 ( .A(n29494), .B(p_input[273]), .Z(n32865) );
  XOR U32356 ( .A(n32906), .B(n32880), .Z(n32874) );
  XNOR U32357 ( .A(p_input[2063]), .B(p_input[287]), .Z(n32880) );
  XOR U32358 ( .A(n32871), .B(n32879), .Z(n32906) );
  XOR U32359 ( .A(n32907), .B(n32876), .Z(n32879) );
  XOR U32360 ( .A(p_input[2061]), .B(p_input[285]), .Z(n32876) );
  XNOR U32361 ( .A(p_input[2062]), .B(p_input[286]), .Z(n32907) );
  XNOR U32362 ( .A(n29036), .B(p_input[281]), .Z(n32871) );
  XNOR U32363 ( .A(n32887), .B(n32886), .Z(n32869) );
  XNOR U32364 ( .A(n32908), .B(n32892), .Z(n32886) );
  XOR U32365 ( .A(p_input[2056]), .B(p_input[280]), .Z(n32892) );
  XOR U32366 ( .A(n32883), .B(n32891), .Z(n32908) );
  XOR U32367 ( .A(n32909), .B(n32888), .Z(n32891) );
  XOR U32368 ( .A(p_input[2054]), .B(p_input[278]), .Z(n32888) );
  XNOR U32369 ( .A(p_input[2055]), .B(p_input[279]), .Z(n32909) );
  XNOR U32370 ( .A(n29039), .B(p_input[274]), .Z(n32883) );
  XNOR U32371 ( .A(n32897), .B(n32896), .Z(n32887) );
  XOR U32372 ( .A(n32910), .B(n32893), .Z(n32896) );
  XOR U32373 ( .A(p_input[2051]), .B(p_input[275]), .Z(n32893) );
  XNOR U32374 ( .A(p_input[2052]), .B(p_input[276]), .Z(n32910) );
  XOR U32375 ( .A(p_input[2053]), .B(p_input[277]), .Z(n32897) );
  XNOR U32376 ( .A(n32911), .B(n32912), .Z(n32795) );
  AND U32377 ( .A(n398), .B(n32913), .Z(n32912) );
  XNOR U32378 ( .A(n32914), .B(n32915), .Z(n398) );
  AND U32379 ( .A(n32916), .B(n32917), .Z(n32915) );
  XOR U32380 ( .A(n32809), .B(n32914), .Z(n32917) );
  XNOR U32381 ( .A(n32918), .B(n32914), .Z(n32916) );
  XOR U32382 ( .A(n32919), .B(n32920), .Z(n32914) );
  AND U32383 ( .A(n32921), .B(n32922), .Z(n32920) );
  XOR U32384 ( .A(n32824), .B(n32919), .Z(n32922) );
  XOR U32385 ( .A(n32919), .B(n32825), .Z(n32921) );
  XOR U32386 ( .A(n32923), .B(n32924), .Z(n32919) );
  AND U32387 ( .A(n32925), .B(n32926), .Z(n32924) );
  XOR U32388 ( .A(n32852), .B(n32923), .Z(n32926) );
  XOR U32389 ( .A(n32923), .B(n32853), .Z(n32925) );
  XOR U32390 ( .A(n32927), .B(n32928), .Z(n32923) );
  AND U32391 ( .A(n32929), .B(n32930), .Z(n32928) );
  XOR U32392 ( .A(n32927), .B(n32901), .Z(n32930) );
  XNOR U32393 ( .A(n32931), .B(n32932), .Z(n32755) );
  AND U32394 ( .A(n402), .B(n32933), .Z(n32932) );
  XNOR U32395 ( .A(n32934), .B(n32935), .Z(n402) );
  AND U32396 ( .A(n32936), .B(n32937), .Z(n32935) );
  XOR U32397 ( .A(n32934), .B(n32765), .Z(n32937) );
  XNOR U32398 ( .A(n32934), .B(n32725), .Z(n32936) );
  XOR U32399 ( .A(n32938), .B(n32939), .Z(n32934) );
  AND U32400 ( .A(n32940), .B(n32941), .Z(n32939) );
  XOR U32401 ( .A(n32938), .B(n32733), .Z(n32940) );
  XOR U32402 ( .A(n32942), .B(n32943), .Z(n32716) );
  AND U32403 ( .A(n406), .B(n32933), .Z(n32943) );
  XNOR U32404 ( .A(n32931), .B(n32942), .Z(n32933) );
  XNOR U32405 ( .A(n32944), .B(n32945), .Z(n406) );
  AND U32406 ( .A(n32946), .B(n32947), .Z(n32945) );
  XNOR U32407 ( .A(n32948), .B(n32944), .Z(n32947) );
  IV U32408 ( .A(n32765), .Z(n32948) );
  XOR U32409 ( .A(n32918), .B(n32949), .Z(n32765) );
  AND U32410 ( .A(n409), .B(n32950), .Z(n32949) );
  XOR U32411 ( .A(n32808), .B(n32805), .Z(n32950) );
  IV U32412 ( .A(n32918), .Z(n32808) );
  XNOR U32413 ( .A(n32725), .B(n32944), .Z(n32946) );
  XOR U32414 ( .A(n32951), .B(n32952), .Z(n32725) );
  AND U32415 ( .A(n425), .B(n32953), .Z(n32952) );
  XOR U32416 ( .A(n32938), .B(n32954), .Z(n32944) );
  AND U32417 ( .A(n32955), .B(n32941), .Z(n32954) );
  XNOR U32418 ( .A(n32775), .B(n32938), .Z(n32941) );
  XOR U32419 ( .A(n32825), .B(n32956), .Z(n32775) );
  AND U32420 ( .A(n409), .B(n32957), .Z(n32956) );
  XOR U32421 ( .A(n32821), .B(n32825), .Z(n32957) );
  XNOR U32422 ( .A(n32958), .B(n32938), .Z(n32955) );
  IV U32423 ( .A(n32733), .Z(n32958) );
  XOR U32424 ( .A(n32959), .B(n32960), .Z(n32733) );
  AND U32425 ( .A(n425), .B(n32961), .Z(n32960) );
  XOR U32426 ( .A(n32962), .B(n32963), .Z(n32938) );
  AND U32427 ( .A(n32964), .B(n32965), .Z(n32963) );
  XNOR U32428 ( .A(n32785), .B(n32962), .Z(n32965) );
  XOR U32429 ( .A(n32853), .B(n32966), .Z(n32785) );
  AND U32430 ( .A(n409), .B(n32967), .Z(n32966) );
  XOR U32431 ( .A(n32849), .B(n32853), .Z(n32967) );
  XOR U32432 ( .A(n32962), .B(n32742), .Z(n32964) );
  XOR U32433 ( .A(n32968), .B(n32969), .Z(n32742) );
  AND U32434 ( .A(n425), .B(n32970), .Z(n32969) );
  XOR U32435 ( .A(n32971), .B(n32972), .Z(n32962) );
  AND U32436 ( .A(n32973), .B(n32974), .Z(n32972) );
  XNOR U32437 ( .A(n32971), .B(n32793), .Z(n32974) );
  XOR U32438 ( .A(n32902), .B(n32975), .Z(n32793) );
  AND U32439 ( .A(n409), .B(n32976), .Z(n32975) );
  XOR U32440 ( .A(n32898), .B(n32902), .Z(n32976) );
  XNOR U32441 ( .A(n32977), .B(n32971), .Z(n32973) );
  IV U32442 ( .A(n32752), .Z(n32977) );
  XOR U32443 ( .A(n32978), .B(n32979), .Z(n32752) );
  AND U32444 ( .A(n425), .B(n32980), .Z(n32979) );
  AND U32445 ( .A(n32942), .B(n32931), .Z(n32971) );
  XNOR U32446 ( .A(n32981), .B(n32982), .Z(n32931) );
  AND U32447 ( .A(n409), .B(n32913), .Z(n32982) );
  XNOR U32448 ( .A(n32911), .B(n32981), .Z(n32913) );
  XNOR U32449 ( .A(n32983), .B(n32984), .Z(n409) );
  AND U32450 ( .A(n32985), .B(n32986), .Z(n32984) );
  XNOR U32451 ( .A(n32983), .B(n32805), .Z(n32986) );
  IV U32452 ( .A(n32809), .Z(n32805) );
  XOR U32453 ( .A(n32987), .B(n32988), .Z(n32809) );
  AND U32454 ( .A(n413), .B(n32989), .Z(n32988) );
  XOR U32455 ( .A(n32990), .B(n32987), .Z(n32989) );
  XNOR U32456 ( .A(n32983), .B(n32918), .Z(n32985) );
  XOR U32457 ( .A(n32991), .B(n32992), .Z(n32918) );
  AND U32458 ( .A(n421), .B(n32953), .Z(n32992) );
  XOR U32459 ( .A(n32951), .B(n32991), .Z(n32953) );
  XOR U32460 ( .A(n32993), .B(n32994), .Z(n32983) );
  AND U32461 ( .A(n32995), .B(n32996), .Z(n32994) );
  XNOR U32462 ( .A(n32993), .B(n32821), .Z(n32996) );
  IV U32463 ( .A(n32824), .Z(n32821) );
  XOR U32464 ( .A(n32997), .B(n32998), .Z(n32824) );
  AND U32465 ( .A(n413), .B(n32999), .Z(n32998) );
  XOR U32466 ( .A(n33000), .B(n32997), .Z(n32999) );
  XOR U32467 ( .A(n32825), .B(n32993), .Z(n32995) );
  XOR U32468 ( .A(n33001), .B(n33002), .Z(n32825) );
  AND U32469 ( .A(n421), .B(n32961), .Z(n33002) );
  XOR U32470 ( .A(n33001), .B(n32959), .Z(n32961) );
  XOR U32471 ( .A(n33003), .B(n33004), .Z(n32993) );
  AND U32472 ( .A(n33005), .B(n33006), .Z(n33004) );
  XNOR U32473 ( .A(n33003), .B(n32849), .Z(n33006) );
  IV U32474 ( .A(n32852), .Z(n32849) );
  XOR U32475 ( .A(n33007), .B(n33008), .Z(n32852) );
  AND U32476 ( .A(n413), .B(n33009), .Z(n33008) );
  XNOR U32477 ( .A(n33010), .B(n33007), .Z(n33009) );
  XOR U32478 ( .A(n32853), .B(n33003), .Z(n33005) );
  XOR U32479 ( .A(n33011), .B(n33012), .Z(n32853) );
  AND U32480 ( .A(n421), .B(n32970), .Z(n33012) );
  XOR U32481 ( .A(n33011), .B(n32968), .Z(n32970) );
  XOR U32482 ( .A(n32927), .B(n33013), .Z(n33003) );
  AND U32483 ( .A(n32929), .B(n33014), .Z(n33013) );
  XNOR U32484 ( .A(n32927), .B(n32898), .Z(n33014) );
  IV U32485 ( .A(n32901), .Z(n32898) );
  XOR U32486 ( .A(n33015), .B(n33016), .Z(n32901) );
  AND U32487 ( .A(n413), .B(n33017), .Z(n33016) );
  XOR U32488 ( .A(n33018), .B(n33015), .Z(n33017) );
  XOR U32489 ( .A(n32902), .B(n32927), .Z(n32929) );
  XOR U32490 ( .A(n33019), .B(n33020), .Z(n32902) );
  AND U32491 ( .A(n421), .B(n32980), .Z(n33020) );
  XOR U32492 ( .A(n33019), .B(n32978), .Z(n32980) );
  AND U32493 ( .A(n32981), .B(n32911), .Z(n32927) );
  XNOR U32494 ( .A(n33021), .B(n33022), .Z(n32911) );
  AND U32495 ( .A(n413), .B(n33023), .Z(n33022) );
  XNOR U32496 ( .A(n33024), .B(n33021), .Z(n33023) );
  XNOR U32497 ( .A(n33025), .B(n33026), .Z(n413) );
  AND U32498 ( .A(n33027), .B(n33028), .Z(n33026) );
  XOR U32499 ( .A(n32990), .B(n33025), .Z(n33028) );
  AND U32500 ( .A(n33029), .B(n33030), .Z(n32990) );
  XNOR U32501 ( .A(n32987), .B(n33025), .Z(n33027) );
  XNOR U32502 ( .A(n33031), .B(n33032), .Z(n32987) );
  AND U32503 ( .A(n417), .B(n33033), .Z(n33032) );
  XNOR U32504 ( .A(n33034), .B(n33035), .Z(n33033) );
  XOR U32505 ( .A(n33036), .B(n33037), .Z(n33025) );
  AND U32506 ( .A(n33038), .B(n33039), .Z(n33037) );
  XNOR U32507 ( .A(n33036), .B(n33029), .Z(n33039) );
  IV U32508 ( .A(n33000), .Z(n33029) );
  XOR U32509 ( .A(n33040), .B(n33041), .Z(n33000) );
  XOR U32510 ( .A(n33042), .B(n33030), .Z(n33041) );
  AND U32511 ( .A(n33010), .B(n33043), .Z(n33030) );
  AND U32512 ( .A(n33044), .B(n33045), .Z(n33042) );
  XOR U32513 ( .A(n33046), .B(n33040), .Z(n33044) );
  XNOR U32514 ( .A(n32997), .B(n33036), .Z(n33038) );
  XNOR U32515 ( .A(n33047), .B(n33048), .Z(n32997) );
  AND U32516 ( .A(n417), .B(n33049), .Z(n33048) );
  XNOR U32517 ( .A(n33050), .B(n33051), .Z(n33049) );
  XOR U32518 ( .A(n33052), .B(n33053), .Z(n33036) );
  AND U32519 ( .A(n33054), .B(n33055), .Z(n33053) );
  XNOR U32520 ( .A(n33052), .B(n33010), .Z(n33055) );
  XOR U32521 ( .A(n33056), .B(n33045), .Z(n33010) );
  XNOR U32522 ( .A(n33057), .B(n33040), .Z(n33045) );
  XOR U32523 ( .A(n33058), .B(n33059), .Z(n33040) );
  AND U32524 ( .A(n33060), .B(n33061), .Z(n33059) );
  XOR U32525 ( .A(n33062), .B(n33058), .Z(n33060) );
  XNOR U32526 ( .A(n33063), .B(n33064), .Z(n33057) );
  AND U32527 ( .A(n33065), .B(n33066), .Z(n33064) );
  XOR U32528 ( .A(n33063), .B(n33067), .Z(n33065) );
  XNOR U32529 ( .A(n33046), .B(n33043), .Z(n33056) );
  AND U32530 ( .A(n33068), .B(n33069), .Z(n33043) );
  XOR U32531 ( .A(n33070), .B(n33071), .Z(n33046) );
  AND U32532 ( .A(n33072), .B(n33073), .Z(n33071) );
  XOR U32533 ( .A(n33070), .B(n33074), .Z(n33072) );
  XNOR U32534 ( .A(n33007), .B(n33052), .Z(n33054) );
  XNOR U32535 ( .A(n33075), .B(n33076), .Z(n33007) );
  AND U32536 ( .A(n417), .B(n33077), .Z(n33076) );
  XNOR U32537 ( .A(n33078), .B(n33079), .Z(n33077) );
  XOR U32538 ( .A(n33080), .B(n33081), .Z(n33052) );
  AND U32539 ( .A(n33082), .B(n33083), .Z(n33081) );
  XNOR U32540 ( .A(n33080), .B(n33068), .Z(n33083) );
  IV U32541 ( .A(n33018), .Z(n33068) );
  XNOR U32542 ( .A(n33084), .B(n33061), .Z(n33018) );
  XNOR U32543 ( .A(n33085), .B(n33067), .Z(n33061) );
  XOR U32544 ( .A(n33086), .B(n33087), .Z(n33067) );
  NOR U32545 ( .A(n33088), .B(n33089), .Z(n33087) );
  XNOR U32546 ( .A(n33086), .B(n33090), .Z(n33088) );
  XNOR U32547 ( .A(n33066), .B(n33058), .Z(n33085) );
  XOR U32548 ( .A(n33091), .B(n33092), .Z(n33058) );
  AND U32549 ( .A(n33093), .B(n33094), .Z(n33092) );
  XNOR U32550 ( .A(n33091), .B(n33095), .Z(n33093) );
  XNOR U32551 ( .A(n33096), .B(n33063), .Z(n33066) );
  XOR U32552 ( .A(n33097), .B(n33098), .Z(n33063) );
  AND U32553 ( .A(n33099), .B(n33100), .Z(n33098) );
  XOR U32554 ( .A(n33097), .B(n33101), .Z(n33099) );
  XNOR U32555 ( .A(n33102), .B(n33103), .Z(n33096) );
  NOR U32556 ( .A(n33104), .B(n33105), .Z(n33103) );
  XOR U32557 ( .A(n33102), .B(n33106), .Z(n33104) );
  XNOR U32558 ( .A(n33062), .B(n33069), .Z(n33084) );
  NOR U32559 ( .A(n33024), .B(n33107), .Z(n33069) );
  XOR U32560 ( .A(n33074), .B(n33073), .Z(n33062) );
  XNOR U32561 ( .A(n33108), .B(n33070), .Z(n33073) );
  XOR U32562 ( .A(n33109), .B(n33110), .Z(n33070) );
  AND U32563 ( .A(n33111), .B(n33112), .Z(n33110) );
  XOR U32564 ( .A(n33109), .B(n33113), .Z(n33111) );
  XNOR U32565 ( .A(n33114), .B(n33115), .Z(n33108) );
  NOR U32566 ( .A(n33116), .B(n33117), .Z(n33115) );
  XNOR U32567 ( .A(n33114), .B(n33118), .Z(n33116) );
  XOR U32568 ( .A(n33119), .B(n33120), .Z(n33074) );
  NOR U32569 ( .A(n33121), .B(n33122), .Z(n33120) );
  XNOR U32570 ( .A(n33119), .B(n33123), .Z(n33121) );
  XNOR U32571 ( .A(n33015), .B(n33080), .Z(n33082) );
  XNOR U32572 ( .A(n33124), .B(n33125), .Z(n33015) );
  AND U32573 ( .A(n417), .B(n33126), .Z(n33125) );
  XNOR U32574 ( .A(n33127), .B(n33128), .Z(n33126) );
  AND U32575 ( .A(n33021), .B(n33024), .Z(n33080) );
  XOR U32576 ( .A(n33129), .B(n33107), .Z(n33024) );
  XNOR U32577 ( .A(p_input[2048]), .B(p_input[288]), .Z(n33107) );
  XOR U32578 ( .A(n33095), .B(n33094), .Z(n33129) );
  XNOR U32579 ( .A(n33130), .B(n33101), .Z(n33094) );
  XNOR U32580 ( .A(n33090), .B(n33089), .Z(n33101) );
  XOR U32581 ( .A(n33131), .B(n33086), .Z(n33089) );
  XNOR U32582 ( .A(n29266), .B(p_input[298]), .Z(n33086) );
  XNOR U32583 ( .A(p_input[2059]), .B(p_input[299]), .Z(n33131) );
  XOR U32584 ( .A(p_input[2060]), .B(p_input[300]), .Z(n33090) );
  XNOR U32585 ( .A(n33100), .B(n33091), .Z(n33130) );
  XNOR U32586 ( .A(n29494), .B(p_input[289]), .Z(n33091) );
  XOR U32587 ( .A(n33132), .B(n33106), .Z(n33100) );
  XNOR U32588 ( .A(p_input[2063]), .B(p_input[303]), .Z(n33106) );
  XOR U32589 ( .A(n33097), .B(n33105), .Z(n33132) );
  XOR U32590 ( .A(n33133), .B(n33102), .Z(n33105) );
  XOR U32591 ( .A(p_input[2061]), .B(p_input[301]), .Z(n33102) );
  XNOR U32592 ( .A(p_input[2062]), .B(p_input[302]), .Z(n33133) );
  XNOR U32593 ( .A(n29036), .B(p_input[297]), .Z(n33097) );
  XNOR U32594 ( .A(n33113), .B(n33112), .Z(n33095) );
  XNOR U32595 ( .A(n33134), .B(n33118), .Z(n33112) );
  XOR U32596 ( .A(p_input[2056]), .B(p_input[296]), .Z(n33118) );
  XOR U32597 ( .A(n33109), .B(n33117), .Z(n33134) );
  XOR U32598 ( .A(n33135), .B(n33114), .Z(n33117) );
  XOR U32599 ( .A(p_input[2054]), .B(p_input[294]), .Z(n33114) );
  XNOR U32600 ( .A(p_input[2055]), .B(p_input[295]), .Z(n33135) );
  XNOR U32601 ( .A(n29039), .B(p_input[290]), .Z(n33109) );
  XNOR U32602 ( .A(n33123), .B(n33122), .Z(n33113) );
  XOR U32603 ( .A(n33136), .B(n33119), .Z(n33122) );
  XOR U32604 ( .A(p_input[2051]), .B(p_input[291]), .Z(n33119) );
  XNOR U32605 ( .A(p_input[2052]), .B(p_input[292]), .Z(n33136) );
  XOR U32606 ( .A(p_input[2053]), .B(p_input[293]), .Z(n33123) );
  XNOR U32607 ( .A(n33137), .B(n33138), .Z(n33021) );
  AND U32608 ( .A(n417), .B(n33139), .Z(n33138) );
  XNOR U32609 ( .A(n33140), .B(n33141), .Z(n417) );
  AND U32610 ( .A(n33142), .B(n33143), .Z(n33141) );
  XOR U32611 ( .A(n33035), .B(n33140), .Z(n33143) );
  XNOR U32612 ( .A(n33144), .B(n33140), .Z(n33142) );
  XOR U32613 ( .A(n33145), .B(n33146), .Z(n33140) );
  AND U32614 ( .A(n33147), .B(n33148), .Z(n33146) );
  XOR U32615 ( .A(n33050), .B(n33145), .Z(n33148) );
  XOR U32616 ( .A(n33145), .B(n33051), .Z(n33147) );
  XOR U32617 ( .A(n33149), .B(n33150), .Z(n33145) );
  AND U32618 ( .A(n33151), .B(n33152), .Z(n33150) );
  XOR U32619 ( .A(n33078), .B(n33149), .Z(n33152) );
  XOR U32620 ( .A(n33149), .B(n33079), .Z(n33151) );
  XOR U32621 ( .A(n33153), .B(n33154), .Z(n33149) );
  AND U32622 ( .A(n33155), .B(n33156), .Z(n33154) );
  XOR U32623 ( .A(n33153), .B(n33127), .Z(n33156) );
  XNOR U32624 ( .A(n33157), .B(n33158), .Z(n32981) );
  AND U32625 ( .A(n421), .B(n33159), .Z(n33158) );
  XNOR U32626 ( .A(n33160), .B(n33161), .Z(n421) );
  AND U32627 ( .A(n33162), .B(n33163), .Z(n33161) );
  XOR U32628 ( .A(n33160), .B(n32991), .Z(n33163) );
  XNOR U32629 ( .A(n33160), .B(n32951), .Z(n33162) );
  XOR U32630 ( .A(n33164), .B(n33165), .Z(n33160) );
  AND U32631 ( .A(n33166), .B(n33167), .Z(n33165) );
  XOR U32632 ( .A(n33164), .B(n32959), .Z(n33166) );
  XOR U32633 ( .A(n33168), .B(n33169), .Z(n32942) );
  AND U32634 ( .A(n425), .B(n33159), .Z(n33169) );
  XNOR U32635 ( .A(n33157), .B(n33168), .Z(n33159) );
  XNOR U32636 ( .A(n33170), .B(n33171), .Z(n425) );
  AND U32637 ( .A(n33172), .B(n33173), .Z(n33171) );
  XNOR U32638 ( .A(n33174), .B(n33170), .Z(n33173) );
  IV U32639 ( .A(n32991), .Z(n33174) );
  XOR U32640 ( .A(n33144), .B(n33175), .Z(n32991) );
  AND U32641 ( .A(n428), .B(n33176), .Z(n33175) );
  XOR U32642 ( .A(n33034), .B(n33031), .Z(n33176) );
  IV U32643 ( .A(n33144), .Z(n33034) );
  XNOR U32644 ( .A(n32951), .B(n33170), .Z(n33172) );
  XOR U32645 ( .A(n33177), .B(n33178), .Z(n32951) );
  AND U32646 ( .A(n444), .B(n33179), .Z(n33178) );
  XOR U32647 ( .A(n33164), .B(n33180), .Z(n33170) );
  AND U32648 ( .A(n33181), .B(n33167), .Z(n33180) );
  XNOR U32649 ( .A(n33001), .B(n33164), .Z(n33167) );
  XOR U32650 ( .A(n33051), .B(n33182), .Z(n33001) );
  AND U32651 ( .A(n428), .B(n33183), .Z(n33182) );
  XOR U32652 ( .A(n33047), .B(n33051), .Z(n33183) );
  XNOR U32653 ( .A(n33184), .B(n33164), .Z(n33181) );
  IV U32654 ( .A(n32959), .Z(n33184) );
  XOR U32655 ( .A(n33185), .B(n33186), .Z(n32959) );
  AND U32656 ( .A(n444), .B(n33187), .Z(n33186) );
  XOR U32657 ( .A(n33188), .B(n33189), .Z(n33164) );
  AND U32658 ( .A(n33190), .B(n33191), .Z(n33189) );
  XNOR U32659 ( .A(n33011), .B(n33188), .Z(n33191) );
  XOR U32660 ( .A(n33079), .B(n33192), .Z(n33011) );
  AND U32661 ( .A(n428), .B(n33193), .Z(n33192) );
  XOR U32662 ( .A(n33075), .B(n33079), .Z(n33193) );
  XOR U32663 ( .A(n33188), .B(n32968), .Z(n33190) );
  XOR U32664 ( .A(n33194), .B(n33195), .Z(n32968) );
  AND U32665 ( .A(n444), .B(n33196), .Z(n33195) );
  XOR U32666 ( .A(n33197), .B(n33198), .Z(n33188) );
  AND U32667 ( .A(n33199), .B(n33200), .Z(n33198) );
  XNOR U32668 ( .A(n33197), .B(n33019), .Z(n33200) );
  XOR U32669 ( .A(n33128), .B(n33201), .Z(n33019) );
  AND U32670 ( .A(n428), .B(n33202), .Z(n33201) );
  XOR U32671 ( .A(n33124), .B(n33128), .Z(n33202) );
  XNOR U32672 ( .A(n33203), .B(n33197), .Z(n33199) );
  IV U32673 ( .A(n32978), .Z(n33203) );
  XOR U32674 ( .A(n33204), .B(n33205), .Z(n32978) );
  AND U32675 ( .A(n444), .B(n33206), .Z(n33205) );
  AND U32676 ( .A(n33168), .B(n33157), .Z(n33197) );
  XNOR U32677 ( .A(n33207), .B(n33208), .Z(n33157) );
  AND U32678 ( .A(n428), .B(n33139), .Z(n33208) );
  XNOR U32679 ( .A(n33137), .B(n33207), .Z(n33139) );
  XNOR U32680 ( .A(n33209), .B(n33210), .Z(n428) );
  AND U32681 ( .A(n33211), .B(n33212), .Z(n33210) );
  XNOR U32682 ( .A(n33209), .B(n33031), .Z(n33212) );
  IV U32683 ( .A(n33035), .Z(n33031) );
  XOR U32684 ( .A(n33213), .B(n33214), .Z(n33035) );
  AND U32685 ( .A(n432), .B(n33215), .Z(n33214) );
  XOR U32686 ( .A(n33216), .B(n33213), .Z(n33215) );
  XNOR U32687 ( .A(n33209), .B(n33144), .Z(n33211) );
  XOR U32688 ( .A(n33217), .B(n33218), .Z(n33144) );
  AND U32689 ( .A(n440), .B(n33179), .Z(n33218) );
  XOR U32690 ( .A(n33177), .B(n33217), .Z(n33179) );
  XOR U32691 ( .A(n33219), .B(n33220), .Z(n33209) );
  AND U32692 ( .A(n33221), .B(n33222), .Z(n33220) );
  XNOR U32693 ( .A(n33219), .B(n33047), .Z(n33222) );
  IV U32694 ( .A(n33050), .Z(n33047) );
  XOR U32695 ( .A(n33223), .B(n33224), .Z(n33050) );
  AND U32696 ( .A(n432), .B(n33225), .Z(n33224) );
  XOR U32697 ( .A(n33226), .B(n33223), .Z(n33225) );
  XOR U32698 ( .A(n33051), .B(n33219), .Z(n33221) );
  XOR U32699 ( .A(n33227), .B(n33228), .Z(n33051) );
  AND U32700 ( .A(n440), .B(n33187), .Z(n33228) );
  XOR U32701 ( .A(n33227), .B(n33185), .Z(n33187) );
  XOR U32702 ( .A(n33229), .B(n33230), .Z(n33219) );
  AND U32703 ( .A(n33231), .B(n33232), .Z(n33230) );
  XNOR U32704 ( .A(n33229), .B(n33075), .Z(n33232) );
  IV U32705 ( .A(n33078), .Z(n33075) );
  XOR U32706 ( .A(n33233), .B(n33234), .Z(n33078) );
  AND U32707 ( .A(n432), .B(n33235), .Z(n33234) );
  XNOR U32708 ( .A(n33236), .B(n33233), .Z(n33235) );
  XOR U32709 ( .A(n33079), .B(n33229), .Z(n33231) );
  XOR U32710 ( .A(n33237), .B(n33238), .Z(n33079) );
  AND U32711 ( .A(n440), .B(n33196), .Z(n33238) );
  XOR U32712 ( .A(n33237), .B(n33194), .Z(n33196) );
  XOR U32713 ( .A(n33153), .B(n33239), .Z(n33229) );
  AND U32714 ( .A(n33155), .B(n33240), .Z(n33239) );
  XNOR U32715 ( .A(n33153), .B(n33124), .Z(n33240) );
  IV U32716 ( .A(n33127), .Z(n33124) );
  XOR U32717 ( .A(n33241), .B(n33242), .Z(n33127) );
  AND U32718 ( .A(n432), .B(n33243), .Z(n33242) );
  XOR U32719 ( .A(n33244), .B(n33241), .Z(n33243) );
  XOR U32720 ( .A(n33128), .B(n33153), .Z(n33155) );
  XOR U32721 ( .A(n33245), .B(n33246), .Z(n33128) );
  AND U32722 ( .A(n440), .B(n33206), .Z(n33246) );
  XOR U32723 ( .A(n33245), .B(n33204), .Z(n33206) );
  AND U32724 ( .A(n33207), .B(n33137), .Z(n33153) );
  XNOR U32725 ( .A(n33247), .B(n33248), .Z(n33137) );
  AND U32726 ( .A(n432), .B(n33249), .Z(n33248) );
  XNOR U32727 ( .A(n33250), .B(n33247), .Z(n33249) );
  XNOR U32728 ( .A(n33251), .B(n33252), .Z(n432) );
  AND U32729 ( .A(n33253), .B(n33254), .Z(n33252) );
  XOR U32730 ( .A(n33216), .B(n33251), .Z(n33254) );
  AND U32731 ( .A(n33255), .B(n33256), .Z(n33216) );
  XNOR U32732 ( .A(n33213), .B(n33251), .Z(n33253) );
  XNOR U32733 ( .A(n33257), .B(n33258), .Z(n33213) );
  AND U32734 ( .A(n436), .B(n33259), .Z(n33258) );
  XNOR U32735 ( .A(n33260), .B(n33261), .Z(n33259) );
  XOR U32736 ( .A(n33262), .B(n33263), .Z(n33251) );
  AND U32737 ( .A(n33264), .B(n33265), .Z(n33263) );
  XNOR U32738 ( .A(n33262), .B(n33255), .Z(n33265) );
  IV U32739 ( .A(n33226), .Z(n33255) );
  XOR U32740 ( .A(n33266), .B(n33267), .Z(n33226) );
  XOR U32741 ( .A(n33268), .B(n33256), .Z(n33267) );
  AND U32742 ( .A(n33236), .B(n33269), .Z(n33256) );
  AND U32743 ( .A(n33270), .B(n33271), .Z(n33268) );
  XOR U32744 ( .A(n33272), .B(n33266), .Z(n33270) );
  XNOR U32745 ( .A(n33223), .B(n33262), .Z(n33264) );
  XNOR U32746 ( .A(n33273), .B(n33274), .Z(n33223) );
  AND U32747 ( .A(n436), .B(n33275), .Z(n33274) );
  XNOR U32748 ( .A(n33276), .B(n33277), .Z(n33275) );
  XOR U32749 ( .A(n33278), .B(n33279), .Z(n33262) );
  AND U32750 ( .A(n33280), .B(n33281), .Z(n33279) );
  XNOR U32751 ( .A(n33278), .B(n33236), .Z(n33281) );
  XOR U32752 ( .A(n33282), .B(n33271), .Z(n33236) );
  XNOR U32753 ( .A(n33283), .B(n33266), .Z(n33271) );
  XOR U32754 ( .A(n33284), .B(n33285), .Z(n33266) );
  AND U32755 ( .A(n33286), .B(n33287), .Z(n33285) );
  XOR U32756 ( .A(n33288), .B(n33284), .Z(n33286) );
  XNOR U32757 ( .A(n33289), .B(n33290), .Z(n33283) );
  AND U32758 ( .A(n33291), .B(n33292), .Z(n33290) );
  XOR U32759 ( .A(n33289), .B(n33293), .Z(n33291) );
  XNOR U32760 ( .A(n33272), .B(n33269), .Z(n33282) );
  AND U32761 ( .A(n33294), .B(n33295), .Z(n33269) );
  XOR U32762 ( .A(n33296), .B(n33297), .Z(n33272) );
  AND U32763 ( .A(n33298), .B(n33299), .Z(n33297) );
  XOR U32764 ( .A(n33296), .B(n33300), .Z(n33298) );
  XNOR U32765 ( .A(n33233), .B(n33278), .Z(n33280) );
  XNOR U32766 ( .A(n33301), .B(n33302), .Z(n33233) );
  AND U32767 ( .A(n436), .B(n33303), .Z(n33302) );
  XNOR U32768 ( .A(n33304), .B(n33305), .Z(n33303) );
  XOR U32769 ( .A(n33306), .B(n33307), .Z(n33278) );
  AND U32770 ( .A(n33308), .B(n33309), .Z(n33307) );
  XNOR U32771 ( .A(n33306), .B(n33294), .Z(n33309) );
  IV U32772 ( .A(n33244), .Z(n33294) );
  XNOR U32773 ( .A(n33310), .B(n33287), .Z(n33244) );
  XNOR U32774 ( .A(n33311), .B(n33293), .Z(n33287) );
  XOR U32775 ( .A(n33312), .B(n33313), .Z(n33293) );
  NOR U32776 ( .A(n33314), .B(n33315), .Z(n33313) );
  XNOR U32777 ( .A(n33312), .B(n33316), .Z(n33314) );
  XNOR U32778 ( .A(n33292), .B(n33284), .Z(n33311) );
  XOR U32779 ( .A(n33317), .B(n33318), .Z(n33284) );
  AND U32780 ( .A(n33319), .B(n33320), .Z(n33318) );
  XNOR U32781 ( .A(n33317), .B(n33321), .Z(n33319) );
  XNOR U32782 ( .A(n33322), .B(n33289), .Z(n33292) );
  XOR U32783 ( .A(n33323), .B(n33324), .Z(n33289) );
  AND U32784 ( .A(n33325), .B(n33326), .Z(n33324) );
  XOR U32785 ( .A(n33323), .B(n33327), .Z(n33325) );
  XNOR U32786 ( .A(n33328), .B(n33329), .Z(n33322) );
  NOR U32787 ( .A(n33330), .B(n33331), .Z(n33329) );
  XOR U32788 ( .A(n33328), .B(n33332), .Z(n33330) );
  XNOR U32789 ( .A(n33288), .B(n33295), .Z(n33310) );
  NOR U32790 ( .A(n33250), .B(n33333), .Z(n33295) );
  XOR U32791 ( .A(n33300), .B(n33299), .Z(n33288) );
  XNOR U32792 ( .A(n33334), .B(n33296), .Z(n33299) );
  XOR U32793 ( .A(n33335), .B(n33336), .Z(n33296) );
  AND U32794 ( .A(n33337), .B(n33338), .Z(n33336) );
  XOR U32795 ( .A(n33335), .B(n33339), .Z(n33337) );
  XNOR U32796 ( .A(n33340), .B(n33341), .Z(n33334) );
  NOR U32797 ( .A(n33342), .B(n33343), .Z(n33341) );
  XNOR U32798 ( .A(n33340), .B(n33344), .Z(n33342) );
  XOR U32799 ( .A(n33345), .B(n33346), .Z(n33300) );
  NOR U32800 ( .A(n33347), .B(n33348), .Z(n33346) );
  XNOR U32801 ( .A(n33345), .B(n33349), .Z(n33347) );
  XNOR U32802 ( .A(n33241), .B(n33306), .Z(n33308) );
  XNOR U32803 ( .A(n33350), .B(n33351), .Z(n33241) );
  AND U32804 ( .A(n436), .B(n33352), .Z(n33351) );
  XNOR U32805 ( .A(n33353), .B(n33354), .Z(n33352) );
  AND U32806 ( .A(n33247), .B(n33250), .Z(n33306) );
  XOR U32807 ( .A(n33355), .B(n33333), .Z(n33250) );
  XNOR U32808 ( .A(p_input[2048]), .B(p_input[304]), .Z(n33333) );
  XOR U32809 ( .A(n33321), .B(n33320), .Z(n33355) );
  XNOR U32810 ( .A(n33356), .B(n33327), .Z(n33320) );
  XNOR U32811 ( .A(n33316), .B(n33315), .Z(n33327) );
  XOR U32812 ( .A(n33357), .B(n33312), .Z(n33315) );
  XNOR U32813 ( .A(n29266), .B(p_input[314]), .Z(n33312) );
  XNOR U32814 ( .A(p_input[2059]), .B(p_input[315]), .Z(n33357) );
  XOR U32815 ( .A(p_input[2060]), .B(p_input[316]), .Z(n33316) );
  XNOR U32816 ( .A(n33326), .B(n33317), .Z(n33356) );
  XNOR U32817 ( .A(n29494), .B(p_input[305]), .Z(n33317) );
  XOR U32818 ( .A(n33358), .B(n33332), .Z(n33326) );
  XNOR U32819 ( .A(p_input[2063]), .B(p_input[319]), .Z(n33332) );
  XOR U32820 ( .A(n33323), .B(n33331), .Z(n33358) );
  XOR U32821 ( .A(n33359), .B(n33328), .Z(n33331) );
  XOR U32822 ( .A(p_input[2061]), .B(p_input[317]), .Z(n33328) );
  XNOR U32823 ( .A(p_input[2062]), .B(p_input[318]), .Z(n33359) );
  XNOR U32824 ( .A(n29036), .B(p_input[313]), .Z(n33323) );
  XNOR U32825 ( .A(n33339), .B(n33338), .Z(n33321) );
  XNOR U32826 ( .A(n33360), .B(n33344), .Z(n33338) );
  XOR U32827 ( .A(p_input[2056]), .B(p_input[312]), .Z(n33344) );
  XOR U32828 ( .A(n33335), .B(n33343), .Z(n33360) );
  XOR U32829 ( .A(n33361), .B(n33340), .Z(n33343) );
  XOR U32830 ( .A(p_input[2054]), .B(p_input[310]), .Z(n33340) );
  XNOR U32831 ( .A(p_input[2055]), .B(p_input[311]), .Z(n33361) );
  XNOR U32832 ( .A(n29039), .B(p_input[306]), .Z(n33335) );
  XNOR U32833 ( .A(n33349), .B(n33348), .Z(n33339) );
  XOR U32834 ( .A(n33362), .B(n33345), .Z(n33348) );
  XOR U32835 ( .A(p_input[2051]), .B(p_input[307]), .Z(n33345) );
  XNOR U32836 ( .A(p_input[2052]), .B(p_input[308]), .Z(n33362) );
  XOR U32837 ( .A(p_input[2053]), .B(p_input[309]), .Z(n33349) );
  XNOR U32838 ( .A(n33363), .B(n33364), .Z(n33247) );
  AND U32839 ( .A(n436), .B(n33365), .Z(n33364) );
  XNOR U32840 ( .A(n33366), .B(n33367), .Z(n436) );
  AND U32841 ( .A(n33368), .B(n33369), .Z(n33367) );
  XOR U32842 ( .A(n33261), .B(n33366), .Z(n33369) );
  XNOR U32843 ( .A(n33370), .B(n33366), .Z(n33368) );
  XOR U32844 ( .A(n33371), .B(n33372), .Z(n33366) );
  AND U32845 ( .A(n33373), .B(n33374), .Z(n33372) );
  XOR U32846 ( .A(n33276), .B(n33371), .Z(n33374) );
  XOR U32847 ( .A(n33371), .B(n33277), .Z(n33373) );
  XOR U32848 ( .A(n33375), .B(n33376), .Z(n33371) );
  AND U32849 ( .A(n33377), .B(n33378), .Z(n33376) );
  XOR U32850 ( .A(n33304), .B(n33375), .Z(n33378) );
  XOR U32851 ( .A(n33375), .B(n33305), .Z(n33377) );
  XOR U32852 ( .A(n33379), .B(n33380), .Z(n33375) );
  AND U32853 ( .A(n33381), .B(n33382), .Z(n33380) );
  XOR U32854 ( .A(n33379), .B(n33353), .Z(n33382) );
  XNOR U32855 ( .A(n33383), .B(n33384), .Z(n33207) );
  AND U32856 ( .A(n440), .B(n33385), .Z(n33384) );
  XNOR U32857 ( .A(n33386), .B(n33387), .Z(n440) );
  AND U32858 ( .A(n33388), .B(n33389), .Z(n33387) );
  XOR U32859 ( .A(n33386), .B(n33217), .Z(n33389) );
  XNOR U32860 ( .A(n33386), .B(n33177), .Z(n33388) );
  XOR U32861 ( .A(n33390), .B(n33391), .Z(n33386) );
  AND U32862 ( .A(n33392), .B(n33393), .Z(n33391) );
  XOR U32863 ( .A(n33390), .B(n33185), .Z(n33392) );
  XOR U32864 ( .A(n33394), .B(n33395), .Z(n33168) );
  AND U32865 ( .A(n444), .B(n33385), .Z(n33395) );
  XNOR U32866 ( .A(n33383), .B(n33394), .Z(n33385) );
  XNOR U32867 ( .A(n33396), .B(n33397), .Z(n444) );
  AND U32868 ( .A(n33398), .B(n33399), .Z(n33397) );
  XNOR U32869 ( .A(n33400), .B(n33396), .Z(n33399) );
  IV U32870 ( .A(n33217), .Z(n33400) );
  XOR U32871 ( .A(n33370), .B(n33401), .Z(n33217) );
  AND U32872 ( .A(n447), .B(n33402), .Z(n33401) );
  XOR U32873 ( .A(n33260), .B(n33257), .Z(n33402) );
  IV U32874 ( .A(n33370), .Z(n33260) );
  XNOR U32875 ( .A(n33177), .B(n33396), .Z(n33398) );
  XOR U32876 ( .A(n33403), .B(n33404), .Z(n33177) );
  AND U32877 ( .A(n463), .B(n33405), .Z(n33404) );
  XOR U32878 ( .A(n33390), .B(n33406), .Z(n33396) );
  AND U32879 ( .A(n33407), .B(n33393), .Z(n33406) );
  XNOR U32880 ( .A(n33227), .B(n33390), .Z(n33393) );
  XOR U32881 ( .A(n33277), .B(n33408), .Z(n33227) );
  AND U32882 ( .A(n447), .B(n33409), .Z(n33408) );
  XOR U32883 ( .A(n33273), .B(n33277), .Z(n33409) );
  XNOR U32884 ( .A(n33410), .B(n33390), .Z(n33407) );
  IV U32885 ( .A(n33185), .Z(n33410) );
  XOR U32886 ( .A(n33411), .B(n33412), .Z(n33185) );
  AND U32887 ( .A(n463), .B(n33413), .Z(n33412) );
  XOR U32888 ( .A(n33414), .B(n33415), .Z(n33390) );
  AND U32889 ( .A(n33416), .B(n33417), .Z(n33415) );
  XNOR U32890 ( .A(n33237), .B(n33414), .Z(n33417) );
  XOR U32891 ( .A(n33305), .B(n33418), .Z(n33237) );
  AND U32892 ( .A(n447), .B(n33419), .Z(n33418) );
  XOR U32893 ( .A(n33301), .B(n33305), .Z(n33419) );
  XOR U32894 ( .A(n33414), .B(n33194), .Z(n33416) );
  XOR U32895 ( .A(n33420), .B(n33421), .Z(n33194) );
  AND U32896 ( .A(n463), .B(n33422), .Z(n33421) );
  XOR U32897 ( .A(n33423), .B(n33424), .Z(n33414) );
  AND U32898 ( .A(n33425), .B(n33426), .Z(n33424) );
  XNOR U32899 ( .A(n33423), .B(n33245), .Z(n33426) );
  XOR U32900 ( .A(n33354), .B(n33427), .Z(n33245) );
  AND U32901 ( .A(n447), .B(n33428), .Z(n33427) );
  XOR U32902 ( .A(n33350), .B(n33354), .Z(n33428) );
  XNOR U32903 ( .A(n33429), .B(n33423), .Z(n33425) );
  IV U32904 ( .A(n33204), .Z(n33429) );
  XOR U32905 ( .A(n33430), .B(n33431), .Z(n33204) );
  AND U32906 ( .A(n463), .B(n33432), .Z(n33431) );
  AND U32907 ( .A(n33394), .B(n33383), .Z(n33423) );
  XNOR U32908 ( .A(n33433), .B(n33434), .Z(n33383) );
  AND U32909 ( .A(n447), .B(n33365), .Z(n33434) );
  XNOR U32910 ( .A(n33363), .B(n33433), .Z(n33365) );
  XNOR U32911 ( .A(n33435), .B(n33436), .Z(n447) );
  AND U32912 ( .A(n33437), .B(n33438), .Z(n33436) );
  XNOR U32913 ( .A(n33435), .B(n33257), .Z(n33438) );
  IV U32914 ( .A(n33261), .Z(n33257) );
  XOR U32915 ( .A(n33439), .B(n33440), .Z(n33261) );
  AND U32916 ( .A(n451), .B(n33441), .Z(n33440) );
  XOR U32917 ( .A(n33442), .B(n33439), .Z(n33441) );
  XNOR U32918 ( .A(n33435), .B(n33370), .Z(n33437) );
  XOR U32919 ( .A(n33443), .B(n33444), .Z(n33370) );
  AND U32920 ( .A(n459), .B(n33405), .Z(n33444) );
  XOR U32921 ( .A(n33403), .B(n33443), .Z(n33405) );
  XOR U32922 ( .A(n33445), .B(n33446), .Z(n33435) );
  AND U32923 ( .A(n33447), .B(n33448), .Z(n33446) );
  XNOR U32924 ( .A(n33445), .B(n33273), .Z(n33448) );
  IV U32925 ( .A(n33276), .Z(n33273) );
  XOR U32926 ( .A(n33449), .B(n33450), .Z(n33276) );
  AND U32927 ( .A(n451), .B(n33451), .Z(n33450) );
  XOR U32928 ( .A(n33452), .B(n33449), .Z(n33451) );
  XOR U32929 ( .A(n33277), .B(n33445), .Z(n33447) );
  XOR U32930 ( .A(n33453), .B(n33454), .Z(n33277) );
  AND U32931 ( .A(n459), .B(n33413), .Z(n33454) );
  XOR U32932 ( .A(n33453), .B(n33411), .Z(n33413) );
  XOR U32933 ( .A(n33455), .B(n33456), .Z(n33445) );
  AND U32934 ( .A(n33457), .B(n33458), .Z(n33456) );
  XNOR U32935 ( .A(n33455), .B(n33301), .Z(n33458) );
  IV U32936 ( .A(n33304), .Z(n33301) );
  XOR U32937 ( .A(n33459), .B(n33460), .Z(n33304) );
  AND U32938 ( .A(n451), .B(n33461), .Z(n33460) );
  XNOR U32939 ( .A(n33462), .B(n33459), .Z(n33461) );
  XOR U32940 ( .A(n33305), .B(n33455), .Z(n33457) );
  XOR U32941 ( .A(n33463), .B(n33464), .Z(n33305) );
  AND U32942 ( .A(n459), .B(n33422), .Z(n33464) );
  XOR U32943 ( .A(n33463), .B(n33420), .Z(n33422) );
  XOR U32944 ( .A(n33379), .B(n33465), .Z(n33455) );
  AND U32945 ( .A(n33381), .B(n33466), .Z(n33465) );
  XNOR U32946 ( .A(n33379), .B(n33350), .Z(n33466) );
  IV U32947 ( .A(n33353), .Z(n33350) );
  XOR U32948 ( .A(n33467), .B(n33468), .Z(n33353) );
  AND U32949 ( .A(n451), .B(n33469), .Z(n33468) );
  XOR U32950 ( .A(n33470), .B(n33467), .Z(n33469) );
  XOR U32951 ( .A(n33354), .B(n33379), .Z(n33381) );
  XOR U32952 ( .A(n33471), .B(n33472), .Z(n33354) );
  AND U32953 ( .A(n459), .B(n33432), .Z(n33472) );
  XOR U32954 ( .A(n33471), .B(n33430), .Z(n33432) );
  AND U32955 ( .A(n33433), .B(n33363), .Z(n33379) );
  XNOR U32956 ( .A(n33473), .B(n33474), .Z(n33363) );
  AND U32957 ( .A(n451), .B(n33475), .Z(n33474) );
  XNOR U32958 ( .A(n33476), .B(n33473), .Z(n33475) );
  XNOR U32959 ( .A(n33477), .B(n33478), .Z(n451) );
  AND U32960 ( .A(n33479), .B(n33480), .Z(n33478) );
  XOR U32961 ( .A(n33442), .B(n33477), .Z(n33480) );
  AND U32962 ( .A(n33481), .B(n33482), .Z(n33442) );
  XNOR U32963 ( .A(n33439), .B(n33477), .Z(n33479) );
  XNOR U32964 ( .A(n33483), .B(n33484), .Z(n33439) );
  AND U32965 ( .A(n455), .B(n33485), .Z(n33484) );
  XNOR U32966 ( .A(n33486), .B(n33487), .Z(n33485) );
  XOR U32967 ( .A(n33488), .B(n33489), .Z(n33477) );
  AND U32968 ( .A(n33490), .B(n33491), .Z(n33489) );
  XNOR U32969 ( .A(n33488), .B(n33481), .Z(n33491) );
  IV U32970 ( .A(n33452), .Z(n33481) );
  XOR U32971 ( .A(n33492), .B(n33493), .Z(n33452) );
  XOR U32972 ( .A(n33494), .B(n33482), .Z(n33493) );
  AND U32973 ( .A(n33462), .B(n33495), .Z(n33482) );
  AND U32974 ( .A(n33496), .B(n33497), .Z(n33494) );
  XOR U32975 ( .A(n33498), .B(n33492), .Z(n33496) );
  XNOR U32976 ( .A(n33449), .B(n33488), .Z(n33490) );
  XNOR U32977 ( .A(n33499), .B(n33500), .Z(n33449) );
  AND U32978 ( .A(n455), .B(n33501), .Z(n33500) );
  XNOR U32979 ( .A(n33502), .B(n33503), .Z(n33501) );
  XOR U32980 ( .A(n33504), .B(n33505), .Z(n33488) );
  AND U32981 ( .A(n33506), .B(n33507), .Z(n33505) );
  XNOR U32982 ( .A(n33504), .B(n33462), .Z(n33507) );
  XOR U32983 ( .A(n33508), .B(n33497), .Z(n33462) );
  XNOR U32984 ( .A(n33509), .B(n33492), .Z(n33497) );
  XOR U32985 ( .A(n33510), .B(n33511), .Z(n33492) );
  AND U32986 ( .A(n33512), .B(n33513), .Z(n33511) );
  XOR U32987 ( .A(n33514), .B(n33510), .Z(n33512) );
  XNOR U32988 ( .A(n33515), .B(n33516), .Z(n33509) );
  AND U32989 ( .A(n33517), .B(n33518), .Z(n33516) );
  XOR U32990 ( .A(n33515), .B(n33519), .Z(n33517) );
  XNOR U32991 ( .A(n33498), .B(n33495), .Z(n33508) );
  AND U32992 ( .A(n33520), .B(n33521), .Z(n33495) );
  XOR U32993 ( .A(n33522), .B(n33523), .Z(n33498) );
  AND U32994 ( .A(n33524), .B(n33525), .Z(n33523) );
  XOR U32995 ( .A(n33522), .B(n33526), .Z(n33524) );
  XNOR U32996 ( .A(n33459), .B(n33504), .Z(n33506) );
  XNOR U32997 ( .A(n33527), .B(n33528), .Z(n33459) );
  AND U32998 ( .A(n455), .B(n33529), .Z(n33528) );
  XNOR U32999 ( .A(n33530), .B(n33531), .Z(n33529) );
  XOR U33000 ( .A(n33532), .B(n33533), .Z(n33504) );
  AND U33001 ( .A(n33534), .B(n33535), .Z(n33533) );
  XNOR U33002 ( .A(n33532), .B(n33520), .Z(n33535) );
  IV U33003 ( .A(n33470), .Z(n33520) );
  XNOR U33004 ( .A(n33536), .B(n33513), .Z(n33470) );
  XNOR U33005 ( .A(n33537), .B(n33519), .Z(n33513) );
  XOR U33006 ( .A(n33538), .B(n33539), .Z(n33519) );
  NOR U33007 ( .A(n33540), .B(n33541), .Z(n33539) );
  XNOR U33008 ( .A(n33538), .B(n33542), .Z(n33540) );
  XNOR U33009 ( .A(n33518), .B(n33510), .Z(n33537) );
  XOR U33010 ( .A(n33543), .B(n33544), .Z(n33510) );
  AND U33011 ( .A(n33545), .B(n33546), .Z(n33544) );
  XNOR U33012 ( .A(n33543), .B(n33547), .Z(n33545) );
  XNOR U33013 ( .A(n33548), .B(n33515), .Z(n33518) );
  XOR U33014 ( .A(n33549), .B(n33550), .Z(n33515) );
  AND U33015 ( .A(n33551), .B(n33552), .Z(n33550) );
  XOR U33016 ( .A(n33549), .B(n33553), .Z(n33551) );
  XNOR U33017 ( .A(n33554), .B(n33555), .Z(n33548) );
  NOR U33018 ( .A(n33556), .B(n33557), .Z(n33555) );
  XOR U33019 ( .A(n33554), .B(n33558), .Z(n33556) );
  XNOR U33020 ( .A(n33514), .B(n33521), .Z(n33536) );
  NOR U33021 ( .A(n33476), .B(n33559), .Z(n33521) );
  XOR U33022 ( .A(n33526), .B(n33525), .Z(n33514) );
  XNOR U33023 ( .A(n33560), .B(n33522), .Z(n33525) );
  XOR U33024 ( .A(n33561), .B(n33562), .Z(n33522) );
  AND U33025 ( .A(n33563), .B(n33564), .Z(n33562) );
  XOR U33026 ( .A(n33561), .B(n33565), .Z(n33563) );
  XNOR U33027 ( .A(n33566), .B(n33567), .Z(n33560) );
  NOR U33028 ( .A(n33568), .B(n33569), .Z(n33567) );
  XNOR U33029 ( .A(n33566), .B(n33570), .Z(n33568) );
  XOR U33030 ( .A(n33571), .B(n33572), .Z(n33526) );
  NOR U33031 ( .A(n33573), .B(n33574), .Z(n33572) );
  XNOR U33032 ( .A(n33571), .B(n33575), .Z(n33573) );
  XNOR U33033 ( .A(n33467), .B(n33532), .Z(n33534) );
  XNOR U33034 ( .A(n33576), .B(n33577), .Z(n33467) );
  AND U33035 ( .A(n455), .B(n33578), .Z(n33577) );
  XNOR U33036 ( .A(n33579), .B(n33580), .Z(n33578) );
  AND U33037 ( .A(n33473), .B(n33476), .Z(n33532) );
  XOR U33038 ( .A(n33581), .B(n33559), .Z(n33476) );
  XNOR U33039 ( .A(p_input[2048]), .B(p_input[320]), .Z(n33559) );
  XOR U33040 ( .A(n33547), .B(n33546), .Z(n33581) );
  XNOR U33041 ( .A(n33582), .B(n33553), .Z(n33546) );
  XNOR U33042 ( .A(n33542), .B(n33541), .Z(n33553) );
  XOR U33043 ( .A(n33583), .B(n33538), .Z(n33541) );
  XNOR U33044 ( .A(n29266), .B(p_input[330]), .Z(n33538) );
  XNOR U33045 ( .A(p_input[2059]), .B(p_input[331]), .Z(n33583) );
  XOR U33046 ( .A(p_input[2060]), .B(p_input[332]), .Z(n33542) );
  XNOR U33047 ( .A(n33552), .B(n33543), .Z(n33582) );
  XNOR U33048 ( .A(n29494), .B(p_input[321]), .Z(n33543) );
  XOR U33049 ( .A(n33584), .B(n33558), .Z(n33552) );
  XNOR U33050 ( .A(p_input[2063]), .B(p_input[335]), .Z(n33558) );
  XOR U33051 ( .A(n33549), .B(n33557), .Z(n33584) );
  XOR U33052 ( .A(n33585), .B(n33554), .Z(n33557) );
  XOR U33053 ( .A(p_input[2061]), .B(p_input[333]), .Z(n33554) );
  XNOR U33054 ( .A(p_input[2062]), .B(p_input[334]), .Z(n33585) );
  XNOR U33055 ( .A(n29036), .B(p_input[329]), .Z(n33549) );
  XNOR U33056 ( .A(n33565), .B(n33564), .Z(n33547) );
  XNOR U33057 ( .A(n33586), .B(n33570), .Z(n33564) );
  XOR U33058 ( .A(p_input[2056]), .B(p_input[328]), .Z(n33570) );
  XOR U33059 ( .A(n33561), .B(n33569), .Z(n33586) );
  XOR U33060 ( .A(n33587), .B(n33566), .Z(n33569) );
  XOR U33061 ( .A(p_input[2054]), .B(p_input[326]), .Z(n33566) );
  XNOR U33062 ( .A(p_input[2055]), .B(p_input[327]), .Z(n33587) );
  XNOR U33063 ( .A(n29039), .B(p_input[322]), .Z(n33561) );
  XNOR U33064 ( .A(n33575), .B(n33574), .Z(n33565) );
  XOR U33065 ( .A(n33588), .B(n33571), .Z(n33574) );
  XOR U33066 ( .A(p_input[2051]), .B(p_input[323]), .Z(n33571) );
  XNOR U33067 ( .A(p_input[2052]), .B(p_input[324]), .Z(n33588) );
  XOR U33068 ( .A(p_input[2053]), .B(p_input[325]), .Z(n33575) );
  XNOR U33069 ( .A(n33589), .B(n33590), .Z(n33473) );
  AND U33070 ( .A(n455), .B(n33591), .Z(n33590) );
  XNOR U33071 ( .A(n33592), .B(n33593), .Z(n455) );
  AND U33072 ( .A(n33594), .B(n33595), .Z(n33593) );
  XOR U33073 ( .A(n33487), .B(n33592), .Z(n33595) );
  XNOR U33074 ( .A(n33596), .B(n33592), .Z(n33594) );
  XOR U33075 ( .A(n33597), .B(n33598), .Z(n33592) );
  AND U33076 ( .A(n33599), .B(n33600), .Z(n33598) );
  XOR U33077 ( .A(n33502), .B(n33597), .Z(n33600) );
  XOR U33078 ( .A(n33597), .B(n33503), .Z(n33599) );
  XOR U33079 ( .A(n33601), .B(n33602), .Z(n33597) );
  AND U33080 ( .A(n33603), .B(n33604), .Z(n33602) );
  XOR U33081 ( .A(n33530), .B(n33601), .Z(n33604) );
  XOR U33082 ( .A(n33601), .B(n33531), .Z(n33603) );
  XOR U33083 ( .A(n33605), .B(n33606), .Z(n33601) );
  AND U33084 ( .A(n33607), .B(n33608), .Z(n33606) );
  XOR U33085 ( .A(n33605), .B(n33579), .Z(n33608) );
  XNOR U33086 ( .A(n33609), .B(n33610), .Z(n33433) );
  AND U33087 ( .A(n459), .B(n33611), .Z(n33610) );
  XNOR U33088 ( .A(n33612), .B(n33613), .Z(n459) );
  AND U33089 ( .A(n33614), .B(n33615), .Z(n33613) );
  XOR U33090 ( .A(n33612), .B(n33443), .Z(n33615) );
  XNOR U33091 ( .A(n33612), .B(n33403), .Z(n33614) );
  XOR U33092 ( .A(n33616), .B(n33617), .Z(n33612) );
  AND U33093 ( .A(n33618), .B(n33619), .Z(n33617) );
  XOR U33094 ( .A(n33616), .B(n33411), .Z(n33618) );
  XOR U33095 ( .A(n33620), .B(n33621), .Z(n33394) );
  AND U33096 ( .A(n463), .B(n33611), .Z(n33621) );
  XNOR U33097 ( .A(n33609), .B(n33620), .Z(n33611) );
  XNOR U33098 ( .A(n33622), .B(n33623), .Z(n463) );
  AND U33099 ( .A(n33624), .B(n33625), .Z(n33623) );
  XNOR U33100 ( .A(n33626), .B(n33622), .Z(n33625) );
  IV U33101 ( .A(n33443), .Z(n33626) );
  XOR U33102 ( .A(n33596), .B(n33627), .Z(n33443) );
  AND U33103 ( .A(n466), .B(n33628), .Z(n33627) );
  XOR U33104 ( .A(n33486), .B(n33483), .Z(n33628) );
  IV U33105 ( .A(n33596), .Z(n33486) );
  XNOR U33106 ( .A(n33403), .B(n33622), .Z(n33624) );
  XOR U33107 ( .A(n33629), .B(n33630), .Z(n33403) );
  AND U33108 ( .A(n482), .B(n33631), .Z(n33630) );
  XOR U33109 ( .A(n33616), .B(n33632), .Z(n33622) );
  AND U33110 ( .A(n33633), .B(n33619), .Z(n33632) );
  XNOR U33111 ( .A(n33453), .B(n33616), .Z(n33619) );
  XOR U33112 ( .A(n33503), .B(n33634), .Z(n33453) );
  AND U33113 ( .A(n466), .B(n33635), .Z(n33634) );
  XOR U33114 ( .A(n33499), .B(n33503), .Z(n33635) );
  XNOR U33115 ( .A(n33636), .B(n33616), .Z(n33633) );
  IV U33116 ( .A(n33411), .Z(n33636) );
  XOR U33117 ( .A(n33637), .B(n33638), .Z(n33411) );
  AND U33118 ( .A(n482), .B(n33639), .Z(n33638) );
  XOR U33119 ( .A(n33640), .B(n33641), .Z(n33616) );
  AND U33120 ( .A(n33642), .B(n33643), .Z(n33641) );
  XNOR U33121 ( .A(n33463), .B(n33640), .Z(n33643) );
  XOR U33122 ( .A(n33531), .B(n33644), .Z(n33463) );
  AND U33123 ( .A(n466), .B(n33645), .Z(n33644) );
  XOR U33124 ( .A(n33527), .B(n33531), .Z(n33645) );
  XOR U33125 ( .A(n33640), .B(n33420), .Z(n33642) );
  XOR U33126 ( .A(n33646), .B(n33647), .Z(n33420) );
  AND U33127 ( .A(n482), .B(n33648), .Z(n33647) );
  XOR U33128 ( .A(n33649), .B(n33650), .Z(n33640) );
  AND U33129 ( .A(n33651), .B(n33652), .Z(n33650) );
  XNOR U33130 ( .A(n33649), .B(n33471), .Z(n33652) );
  XOR U33131 ( .A(n33580), .B(n33653), .Z(n33471) );
  AND U33132 ( .A(n466), .B(n33654), .Z(n33653) );
  XOR U33133 ( .A(n33576), .B(n33580), .Z(n33654) );
  XNOR U33134 ( .A(n33655), .B(n33649), .Z(n33651) );
  IV U33135 ( .A(n33430), .Z(n33655) );
  XOR U33136 ( .A(n33656), .B(n33657), .Z(n33430) );
  AND U33137 ( .A(n482), .B(n33658), .Z(n33657) );
  AND U33138 ( .A(n33620), .B(n33609), .Z(n33649) );
  XNOR U33139 ( .A(n33659), .B(n33660), .Z(n33609) );
  AND U33140 ( .A(n466), .B(n33591), .Z(n33660) );
  XNOR U33141 ( .A(n33589), .B(n33659), .Z(n33591) );
  XNOR U33142 ( .A(n33661), .B(n33662), .Z(n466) );
  AND U33143 ( .A(n33663), .B(n33664), .Z(n33662) );
  XNOR U33144 ( .A(n33661), .B(n33483), .Z(n33664) );
  IV U33145 ( .A(n33487), .Z(n33483) );
  XOR U33146 ( .A(n33665), .B(n33666), .Z(n33487) );
  AND U33147 ( .A(n470), .B(n33667), .Z(n33666) );
  XOR U33148 ( .A(n33668), .B(n33665), .Z(n33667) );
  XNOR U33149 ( .A(n33661), .B(n33596), .Z(n33663) );
  XOR U33150 ( .A(n33669), .B(n33670), .Z(n33596) );
  AND U33151 ( .A(n478), .B(n33631), .Z(n33670) );
  XOR U33152 ( .A(n33629), .B(n33669), .Z(n33631) );
  XOR U33153 ( .A(n33671), .B(n33672), .Z(n33661) );
  AND U33154 ( .A(n33673), .B(n33674), .Z(n33672) );
  XNOR U33155 ( .A(n33671), .B(n33499), .Z(n33674) );
  IV U33156 ( .A(n33502), .Z(n33499) );
  XOR U33157 ( .A(n33675), .B(n33676), .Z(n33502) );
  AND U33158 ( .A(n470), .B(n33677), .Z(n33676) );
  XOR U33159 ( .A(n33678), .B(n33675), .Z(n33677) );
  XOR U33160 ( .A(n33503), .B(n33671), .Z(n33673) );
  XOR U33161 ( .A(n33679), .B(n33680), .Z(n33503) );
  AND U33162 ( .A(n478), .B(n33639), .Z(n33680) );
  XOR U33163 ( .A(n33679), .B(n33637), .Z(n33639) );
  XOR U33164 ( .A(n33681), .B(n33682), .Z(n33671) );
  AND U33165 ( .A(n33683), .B(n33684), .Z(n33682) );
  XNOR U33166 ( .A(n33681), .B(n33527), .Z(n33684) );
  IV U33167 ( .A(n33530), .Z(n33527) );
  XOR U33168 ( .A(n33685), .B(n33686), .Z(n33530) );
  AND U33169 ( .A(n470), .B(n33687), .Z(n33686) );
  XNOR U33170 ( .A(n33688), .B(n33685), .Z(n33687) );
  XOR U33171 ( .A(n33531), .B(n33681), .Z(n33683) );
  XOR U33172 ( .A(n33689), .B(n33690), .Z(n33531) );
  AND U33173 ( .A(n478), .B(n33648), .Z(n33690) );
  XOR U33174 ( .A(n33689), .B(n33646), .Z(n33648) );
  XOR U33175 ( .A(n33605), .B(n33691), .Z(n33681) );
  AND U33176 ( .A(n33607), .B(n33692), .Z(n33691) );
  XNOR U33177 ( .A(n33605), .B(n33576), .Z(n33692) );
  IV U33178 ( .A(n33579), .Z(n33576) );
  XOR U33179 ( .A(n33693), .B(n33694), .Z(n33579) );
  AND U33180 ( .A(n470), .B(n33695), .Z(n33694) );
  XOR U33181 ( .A(n33696), .B(n33693), .Z(n33695) );
  XOR U33182 ( .A(n33580), .B(n33605), .Z(n33607) );
  XOR U33183 ( .A(n33697), .B(n33698), .Z(n33580) );
  AND U33184 ( .A(n478), .B(n33658), .Z(n33698) );
  XOR U33185 ( .A(n33697), .B(n33656), .Z(n33658) );
  AND U33186 ( .A(n33659), .B(n33589), .Z(n33605) );
  XNOR U33187 ( .A(n33699), .B(n33700), .Z(n33589) );
  AND U33188 ( .A(n470), .B(n33701), .Z(n33700) );
  XNOR U33189 ( .A(n33702), .B(n33699), .Z(n33701) );
  XNOR U33190 ( .A(n33703), .B(n33704), .Z(n470) );
  AND U33191 ( .A(n33705), .B(n33706), .Z(n33704) );
  XOR U33192 ( .A(n33668), .B(n33703), .Z(n33706) );
  AND U33193 ( .A(n33707), .B(n33708), .Z(n33668) );
  XNOR U33194 ( .A(n33665), .B(n33703), .Z(n33705) );
  XNOR U33195 ( .A(n33709), .B(n33710), .Z(n33665) );
  AND U33196 ( .A(n474), .B(n33711), .Z(n33710) );
  XNOR U33197 ( .A(n33712), .B(n33713), .Z(n33711) );
  XOR U33198 ( .A(n33714), .B(n33715), .Z(n33703) );
  AND U33199 ( .A(n33716), .B(n33717), .Z(n33715) );
  XNOR U33200 ( .A(n33714), .B(n33707), .Z(n33717) );
  IV U33201 ( .A(n33678), .Z(n33707) );
  XOR U33202 ( .A(n33718), .B(n33719), .Z(n33678) );
  XOR U33203 ( .A(n33720), .B(n33708), .Z(n33719) );
  AND U33204 ( .A(n33688), .B(n33721), .Z(n33708) );
  AND U33205 ( .A(n33722), .B(n33723), .Z(n33720) );
  XOR U33206 ( .A(n33724), .B(n33718), .Z(n33722) );
  XNOR U33207 ( .A(n33675), .B(n33714), .Z(n33716) );
  XNOR U33208 ( .A(n33725), .B(n33726), .Z(n33675) );
  AND U33209 ( .A(n474), .B(n33727), .Z(n33726) );
  XNOR U33210 ( .A(n33728), .B(n33729), .Z(n33727) );
  XOR U33211 ( .A(n33730), .B(n33731), .Z(n33714) );
  AND U33212 ( .A(n33732), .B(n33733), .Z(n33731) );
  XNOR U33213 ( .A(n33730), .B(n33688), .Z(n33733) );
  XOR U33214 ( .A(n33734), .B(n33723), .Z(n33688) );
  XNOR U33215 ( .A(n33735), .B(n33718), .Z(n33723) );
  XOR U33216 ( .A(n33736), .B(n33737), .Z(n33718) );
  AND U33217 ( .A(n33738), .B(n33739), .Z(n33737) );
  XOR U33218 ( .A(n33740), .B(n33736), .Z(n33738) );
  XNOR U33219 ( .A(n33741), .B(n33742), .Z(n33735) );
  AND U33220 ( .A(n33743), .B(n33744), .Z(n33742) );
  XOR U33221 ( .A(n33741), .B(n33745), .Z(n33743) );
  XNOR U33222 ( .A(n33724), .B(n33721), .Z(n33734) );
  AND U33223 ( .A(n33746), .B(n33747), .Z(n33721) );
  XOR U33224 ( .A(n33748), .B(n33749), .Z(n33724) );
  AND U33225 ( .A(n33750), .B(n33751), .Z(n33749) );
  XOR U33226 ( .A(n33748), .B(n33752), .Z(n33750) );
  XNOR U33227 ( .A(n33685), .B(n33730), .Z(n33732) );
  XNOR U33228 ( .A(n33753), .B(n33754), .Z(n33685) );
  AND U33229 ( .A(n474), .B(n33755), .Z(n33754) );
  XNOR U33230 ( .A(n33756), .B(n33757), .Z(n33755) );
  XOR U33231 ( .A(n33758), .B(n33759), .Z(n33730) );
  AND U33232 ( .A(n33760), .B(n33761), .Z(n33759) );
  XNOR U33233 ( .A(n33758), .B(n33746), .Z(n33761) );
  IV U33234 ( .A(n33696), .Z(n33746) );
  XNOR U33235 ( .A(n33762), .B(n33739), .Z(n33696) );
  XNOR U33236 ( .A(n33763), .B(n33745), .Z(n33739) );
  XOR U33237 ( .A(n33764), .B(n33765), .Z(n33745) );
  NOR U33238 ( .A(n33766), .B(n33767), .Z(n33765) );
  XNOR U33239 ( .A(n33764), .B(n33768), .Z(n33766) );
  XNOR U33240 ( .A(n33744), .B(n33736), .Z(n33763) );
  XOR U33241 ( .A(n33769), .B(n33770), .Z(n33736) );
  AND U33242 ( .A(n33771), .B(n33772), .Z(n33770) );
  XNOR U33243 ( .A(n33769), .B(n33773), .Z(n33771) );
  XNOR U33244 ( .A(n33774), .B(n33741), .Z(n33744) );
  XOR U33245 ( .A(n33775), .B(n33776), .Z(n33741) );
  AND U33246 ( .A(n33777), .B(n33778), .Z(n33776) );
  XOR U33247 ( .A(n33775), .B(n33779), .Z(n33777) );
  XNOR U33248 ( .A(n33780), .B(n33781), .Z(n33774) );
  NOR U33249 ( .A(n33782), .B(n33783), .Z(n33781) );
  XOR U33250 ( .A(n33780), .B(n33784), .Z(n33782) );
  XNOR U33251 ( .A(n33740), .B(n33747), .Z(n33762) );
  NOR U33252 ( .A(n33702), .B(n33785), .Z(n33747) );
  XOR U33253 ( .A(n33752), .B(n33751), .Z(n33740) );
  XNOR U33254 ( .A(n33786), .B(n33748), .Z(n33751) );
  XOR U33255 ( .A(n33787), .B(n33788), .Z(n33748) );
  AND U33256 ( .A(n33789), .B(n33790), .Z(n33788) );
  XOR U33257 ( .A(n33787), .B(n33791), .Z(n33789) );
  XNOR U33258 ( .A(n33792), .B(n33793), .Z(n33786) );
  NOR U33259 ( .A(n33794), .B(n33795), .Z(n33793) );
  XNOR U33260 ( .A(n33792), .B(n33796), .Z(n33794) );
  XOR U33261 ( .A(n33797), .B(n33798), .Z(n33752) );
  NOR U33262 ( .A(n33799), .B(n33800), .Z(n33798) );
  XNOR U33263 ( .A(n33797), .B(n33801), .Z(n33799) );
  XNOR U33264 ( .A(n33693), .B(n33758), .Z(n33760) );
  XNOR U33265 ( .A(n33802), .B(n33803), .Z(n33693) );
  AND U33266 ( .A(n474), .B(n33804), .Z(n33803) );
  XNOR U33267 ( .A(n33805), .B(n33806), .Z(n33804) );
  AND U33268 ( .A(n33699), .B(n33702), .Z(n33758) );
  XOR U33269 ( .A(n33807), .B(n33785), .Z(n33702) );
  XNOR U33270 ( .A(p_input[2048]), .B(p_input[336]), .Z(n33785) );
  XOR U33271 ( .A(n33773), .B(n33772), .Z(n33807) );
  XNOR U33272 ( .A(n33808), .B(n33779), .Z(n33772) );
  XNOR U33273 ( .A(n33768), .B(n33767), .Z(n33779) );
  XOR U33274 ( .A(n33809), .B(n33764), .Z(n33767) );
  XNOR U33275 ( .A(n29266), .B(p_input[346]), .Z(n33764) );
  XNOR U33276 ( .A(p_input[2059]), .B(p_input[347]), .Z(n33809) );
  XOR U33277 ( .A(p_input[2060]), .B(p_input[348]), .Z(n33768) );
  XNOR U33278 ( .A(n33778), .B(n33769), .Z(n33808) );
  XNOR U33279 ( .A(n29494), .B(p_input[337]), .Z(n33769) );
  XOR U33280 ( .A(n33810), .B(n33784), .Z(n33778) );
  XNOR U33281 ( .A(p_input[2063]), .B(p_input[351]), .Z(n33784) );
  XOR U33282 ( .A(n33775), .B(n33783), .Z(n33810) );
  XOR U33283 ( .A(n33811), .B(n33780), .Z(n33783) );
  XOR U33284 ( .A(p_input[2061]), .B(p_input[349]), .Z(n33780) );
  XNOR U33285 ( .A(p_input[2062]), .B(p_input[350]), .Z(n33811) );
  XNOR U33286 ( .A(n29036), .B(p_input[345]), .Z(n33775) );
  XNOR U33287 ( .A(n33791), .B(n33790), .Z(n33773) );
  XNOR U33288 ( .A(n33812), .B(n33796), .Z(n33790) );
  XOR U33289 ( .A(p_input[2056]), .B(p_input[344]), .Z(n33796) );
  XOR U33290 ( .A(n33787), .B(n33795), .Z(n33812) );
  XOR U33291 ( .A(n33813), .B(n33792), .Z(n33795) );
  XOR U33292 ( .A(p_input[2054]), .B(p_input[342]), .Z(n33792) );
  XNOR U33293 ( .A(p_input[2055]), .B(p_input[343]), .Z(n33813) );
  XNOR U33294 ( .A(n29039), .B(p_input[338]), .Z(n33787) );
  XNOR U33295 ( .A(n33801), .B(n33800), .Z(n33791) );
  XOR U33296 ( .A(n33814), .B(n33797), .Z(n33800) );
  XOR U33297 ( .A(p_input[2051]), .B(p_input[339]), .Z(n33797) );
  XNOR U33298 ( .A(p_input[2052]), .B(p_input[340]), .Z(n33814) );
  XOR U33299 ( .A(p_input[2053]), .B(p_input[341]), .Z(n33801) );
  XNOR U33300 ( .A(n33815), .B(n33816), .Z(n33699) );
  AND U33301 ( .A(n474), .B(n33817), .Z(n33816) );
  XNOR U33302 ( .A(n33818), .B(n33819), .Z(n474) );
  AND U33303 ( .A(n33820), .B(n33821), .Z(n33819) );
  XOR U33304 ( .A(n33713), .B(n33818), .Z(n33821) );
  XNOR U33305 ( .A(n33822), .B(n33818), .Z(n33820) );
  XOR U33306 ( .A(n33823), .B(n33824), .Z(n33818) );
  AND U33307 ( .A(n33825), .B(n33826), .Z(n33824) );
  XOR U33308 ( .A(n33728), .B(n33823), .Z(n33826) );
  XOR U33309 ( .A(n33823), .B(n33729), .Z(n33825) );
  XOR U33310 ( .A(n33827), .B(n33828), .Z(n33823) );
  AND U33311 ( .A(n33829), .B(n33830), .Z(n33828) );
  XOR U33312 ( .A(n33756), .B(n33827), .Z(n33830) );
  XOR U33313 ( .A(n33827), .B(n33757), .Z(n33829) );
  XOR U33314 ( .A(n33831), .B(n33832), .Z(n33827) );
  AND U33315 ( .A(n33833), .B(n33834), .Z(n33832) );
  XOR U33316 ( .A(n33831), .B(n33805), .Z(n33834) );
  XNOR U33317 ( .A(n33835), .B(n33836), .Z(n33659) );
  AND U33318 ( .A(n478), .B(n33837), .Z(n33836) );
  XNOR U33319 ( .A(n33838), .B(n33839), .Z(n478) );
  AND U33320 ( .A(n33840), .B(n33841), .Z(n33839) );
  XOR U33321 ( .A(n33838), .B(n33669), .Z(n33841) );
  XNOR U33322 ( .A(n33838), .B(n33629), .Z(n33840) );
  XOR U33323 ( .A(n33842), .B(n33843), .Z(n33838) );
  AND U33324 ( .A(n33844), .B(n33845), .Z(n33843) );
  XOR U33325 ( .A(n33842), .B(n33637), .Z(n33844) );
  XOR U33326 ( .A(n33846), .B(n33847), .Z(n33620) );
  AND U33327 ( .A(n482), .B(n33837), .Z(n33847) );
  XNOR U33328 ( .A(n33835), .B(n33846), .Z(n33837) );
  XNOR U33329 ( .A(n33848), .B(n33849), .Z(n482) );
  AND U33330 ( .A(n33850), .B(n33851), .Z(n33849) );
  XNOR U33331 ( .A(n33852), .B(n33848), .Z(n33851) );
  IV U33332 ( .A(n33669), .Z(n33852) );
  XOR U33333 ( .A(n33822), .B(n33853), .Z(n33669) );
  AND U33334 ( .A(n485), .B(n33854), .Z(n33853) );
  XOR U33335 ( .A(n33712), .B(n33709), .Z(n33854) );
  IV U33336 ( .A(n33822), .Z(n33712) );
  XNOR U33337 ( .A(n33629), .B(n33848), .Z(n33850) );
  XOR U33338 ( .A(n33855), .B(n33856), .Z(n33629) );
  AND U33339 ( .A(n501), .B(n33857), .Z(n33856) );
  XOR U33340 ( .A(n33842), .B(n33858), .Z(n33848) );
  AND U33341 ( .A(n33859), .B(n33845), .Z(n33858) );
  XNOR U33342 ( .A(n33679), .B(n33842), .Z(n33845) );
  XOR U33343 ( .A(n33729), .B(n33860), .Z(n33679) );
  AND U33344 ( .A(n485), .B(n33861), .Z(n33860) );
  XOR U33345 ( .A(n33725), .B(n33729), .Z(n33861) );
  XNOR U33346 ( .A(n33862), .B(n33842), .Z(n33859) );
  IV U33347 ( .A(n33637), .Z(n33862) );
  XOR U33348 ( .A(n33863), .B(n33864), .Z(n33637) );
  AND U33349 ( .A(n501), .B(n33865), .Z(n33864) );
  XOR U33350 ( .A(n33866), .B(n33867), .Z(n33842) );
  AND U33351 ( .A(n33868), .B(n33869), .Z(n33867) );
  XNOR U33352 ( .A(n33689), .B(n33866), .Z(n33869) );
  XOR U33353 ( .A(n33757), .B(n33870), .Z(n33689) );
  AND U33354 ( .A(n485), .B(n33871), .Z(n33870) );
  XOR U33355 ( .A(n33753), .B(n33757), .Z(n33871) );
  XOR U33356 ( .A(n33866), .B(n33646), .Z(n33868) );
  XOR U33357 ( .A(n33872), .B(n33873), .Z(n33646) );
  AND U33358 ( .A(n501), .B(n33874), .Z(n33873) );
  XOR U33359 ( .A(n33875), .B(n33876), .Z(n33866) );
  AND U33360 ( .A(n33877), .B(n33878), .Z(n33876) );
  XNOR U33361 ( .A(n33875), .B(n33697), .Z(n33878) );
  XOR U33362 ( .A(n33806), .B(n33879), .Z(n33697) );
  AND U33363 ( .A(n485), .B(n33880), .Z(n33879) );
  XOR U33364 ( .A(n33802), .B(n33806), .Z(n33880) );
  XNOR U33365 ( .A(n33881), .B(n33875), .Z(n33877) );
  IV U33366 ( .A(n33656), .Z(n33881) );
  XOR U33367 ( .A(n33882), .B(n33883), .Z(n33656) );
  AND U33368 ( .A(n501), .B(n33884), .Z(n33883) );
  AND U33369 ( .A(n33846), .B(n33835), .Z(n33875) );
  XNOR U33370 ( .A(n33885), .B(n33886), .Z(n33835) );
  AND U33371 ( .A(n485), .B(n33817), .Z(n33886) );
  XNOR U33372 ( .A(n33815), .B(n33885), .Z(n33817) );
  XNOR U33373 ( .A(n33887), .B(n33888), .Z(n485) );
  AND U33374 ( .A(n33889), .B(n33890), .Z(n33888) );
  XNOR U33375 ( .A(n33887), .B(n33709), .Z(n33890) );
  IV U33376 ( .A(n33713), .Z(n33709) );
  XOR U33377 ( .A(n33891), .B(n33892), .Z(n33713) );
  AND U33378 ( .A(n489), .B(n33893), .Z(n33892) );
  XOR U33379 ( .A(n33894), .B(n33891), .Z(n33893) );
  XNOR U33380 ( .A(n33887), .B(n33822), .Z(n33889) );
  XOR U33381 ( .A(n33895), .B(n33896), .Z(n33822) );
  AND U33382 ( .A(n497), .B(n33857), .Z(n33896) );
  XOR U33383 ( .A(n33855), .B(n33895), .Z(n33857) );
  XOR U33384 ( .A(n33897), .B(n33898), .Z(n33887) );
  AND U33385 ( .A(n33899), .B(n33900), .Z(n33898) );
  XNOR U33386 ( .A(n33897), .B(n33725), .Z(n33900) );
  IV U33387 ( .A(n33728), .Z(n33725) );
  XOR U33388 ( .A(n33901), .B(n33902), .Z(n33728) );
  AND U33389 ( .A(n489), .B(n33903), .Z(n33902) );
  XOR U33390 ( .A(n33904), .B(n33901), .Z(n33903) );
  XOR U33391 ( .A(n33729), .B(n33897), .Z(n33899) );
  XOR U33392 ( .A(n33905), .B(n33906), .Z(n33729) );
  AND U33393 ( .A(n497), .B(n33865), .Z(n33906) );
  XOR U33394 ( .A(n33905), .B(n33863), .Z(n33865) );
  XOR U33395 ( .A(n33907), .B(n33908), .Z(n33897) );
  AND U33396 ( .A(n33909), .B(n33910), .Z(n33908) );
  XNOR U33397 ( .A(n33907), .B(n33753), .Z(n33910) );
  IV U33398 ( .A(n33756), .Z(n33753) );
  XOR U33399 ( .A(n33911), .B(n33912), .Z(n33756) );
  AND U33400 ( .A(n489), .B(n33913), .Z(n33912) );
  XNOR U33401 ( .A(n33914), .B(n33911), .Z(n33913) );
  XOR U33402 ( .A(n33757), .B(n33907), .Z(n33909) );
  XOR U33403 ( .A(n33915), .B(n33916), .Z(n33757) );
  AND U33404 ( .A(n497), .B(n33874), .Z(n33916) );
  XOR U33405 ( .A(n33915), .B(n33872), .Z(n33874) );
  XOR U33406 ( .A(n33831), .B(n33917), .Z(n33907) );
  AND U33407 ( .A(n33833), .B(n33918), .Z(n33917) );
  XNOR U33408 ( .A(n33831), .B(n33802), .Z(n33918) );
  IV U33409 ( .A(n33805), .Z(n33802) );
  XOR U33410 ( .A(n33919), .B(n33920), .Z(n33805) );
  AND U33411 ( .A(n489), .B(n33921), .Z(n33920) );
  XOR U33412 ( .A(n33922), .B(n33919), .Z(n33921) );
  XOR U33413 ( .A(n33806), .B(n33831), .Z(n33833) );
  XOR U33414 ( .A(n33923), .B(n33924), .Z(n33806) );
  AND U33415 ( .A(n497), .B(n33884), .Z(n33924) );
  XOR U33416 ( .A(n33923), .B(n33882), .Z(n33884) );
  AND U33417 ( .A(n33885), .B(n33815), .Z(n33831) );
  XNOR U33418 ( .A(n33925), .B(n33926), .Z(n33815) );
  AND U33419 ( .A(n489), .B(n33927), .Z(n33926) );
  XNOR U33420 ( .A(n33928), .B(n33925), .Z(n33927) );
  XNOR U33421 ( .A(n33929), .B(n33930), .Z(n489) );
  AND U33422 ( .A(n33931), .B(n33932), .Z(n33930) );
  XOR U33423 ( .A(n33894), .B(n33929), .Z(n33932) );
  AND U33424 ( .A(n33933), .B(n33934), .Z(n33894) );
  XNOR U33425 ( .A(n33891), .B(n33929), .Z(n33931) );
  XNOR U33426 ( .A(n33935), .B(n33936), .Z(n33891) );
  AND U33427 ( .A(n493), .B(n33937), .Z(n33936) );
  XNOR U33428 ( .A(n33938), .B(n33939), .Z(n33937) );
  XOR U33429 ( .A(n33940), .B(n33941), .Z(n33929) );
  AND U33430 ( .A(n33942), .B(n33943), .Z(n33941) );
  XNOR U33431 ( .A(n33940), .B(n33933), .Z(n33943) );
  IV U33432 ( .A(n33904), .Z(n33933) );
  XOR U33433 ( .A(n33944), .B(n33945), .Z(n33904) );
  XOR U33434 ( .A(n33946), .B(n33934), .Z(n33945) );
  AND U33435 ( .A(n33914), .B(n33947), .Z(n33934) );
  AND U33436 ( .A(n33948), .B(n33949), .Z(n33946) );
  XOR U33437 ( .A(n33950), .B(n33944), .Z(n33948) );
  XNOR U33438 ( .A(n33901), .B(n33940), .Z(n33942) );
  XNOR U33439 ( .A(n33951), .B(n33952), .Z(n33901) );
  AND U33440 ( .A(n493), .B(n33953), .Z(n33952) );
  XNOR U33441 ( .A(n33954), .B(n33955), .Z(n33953) );
  XOR U33442 ( .A(n33956), .B(n33957), .Z(n33940) );
  AND U33443 ( .A(n33958), .B(n33959), .Z(n33957) );
  XNOR U33444 ( .A(n33956), .B(n33914), .Z(n33959) );
  XOR U33445 ( .A(n33960), .B(n33949), .Z(n33914) );
  XNOR U33446 ( .A(n33961), .B(n33944), .Z(n33949) );
  XOR U33447 ( .A(n33962), .B(n33963), .Z(n33944) );
  AND U33448 ( .A(n33964), .B(n33965), .Z(n33963) );
  XOR U33449 ( .A(n33966), .B(n33962), .Z(n33964) );
  XNOR U33450 ( .A(n33967), .B(n33968), .Z(n33961) );
  AND U33451 ( .A(n33969), .B(n33970), .Z(n33968) );
  XOR U33452 ( .A(n33967), .B(n33971), .Z(n33969) );
  XNOR U33453 ( .A(n33950), .B(n33947), .Z(n33960) );
  AND U33454 ( .A(n33972), .B(n33973), .Z(n33947) );
  XOR U33455 ( .A(n33974), .B(n33975), .Z(n33950) );
  AND U33456 ( .A(n33976), .B(n33977), .Z(n33975) );
  XOR U33457 ( .A(n33974), .B(n33978), .Z(n33976) );
  XNOR U33458 ( .A(n33911), .B(n33956), .Z(n33958) );
  XNOR U33459 ( .A(n33979), .B(n33980), .Z(n33911) );
  AND U33460 ( .A(n493), .B(n33981), .Z(n33980) );
  XNOR U33461 ( .A(n33982), .B(n33983), .Z(n33981) );
  XOR U33462 ( .A(n33984), .B(n33985), .Z(n33956) );
  AND U33463 ( .A(n33986), .B(n33987), .Z(n33985) );
  XNOR U33464 ( .A(n33984), .B(n33972), .Z(n33987) );
  IV U33465 ( .A(n33922), .Z(n33972) );
  XNOR U33466 ( .A(n33988), .B(n33965), .Z(n33922) );
  XNOR U33467 ( .A(n33989), .B(n33971), .Z(n33965) );
  XOR U33468 ( .A(n33990), .B(n33991), .Z(n33971) );
  NOR U33469 ( .A(n33992), .B(n33993), .Z(n33991) );
  XNOR U33470 ( .A(n33990), .B(n33994), .Z(n33992) );
  XNOR U33471 ( .A(n33970), .B(n33962), .Z(n33989) );
  XOR U33472 ( .A(n33995), .B(n33996), .Z(n33962) );
  AND U33473 ( .A(n33997), .B(n33998), .Z(n33996) );
  XNOR U33474 ( .A(n33995), .B(n33999), .Z(n33997) );
  XNOR U33475 ( .A(n34000), .B(n33967), .Z(n33970) );
  XOR U33476 ( .A(n34001), .B(n34002), .Z(n33967) );
  AND U33477 ( .A(n34003), .B(n34004), .Z(n34002) );
  XOR U33478 ( .A(n34001), .B(n34005), .Z(n34003) );
  XNOR U33479 ( .A(n34006), .B(n34007), .Z(n34000) );
  NOR U33480 ( .A(n34008), .B(n34009), .Z(n34007) );
  XOR U33481 ( .A(n34006), .B(n34010), .Z(n34008) );
  XNOR U33482 ( .A(n33966), .B(n33973), .Z(n33988) );
  NOR U33483 ( .A(n33928), .B(n34011), .Z(n33973) );
  XOR U33484 ( .A(n33978), .B(n33977), .Z(n33966) );
  XNOR U33485 ( .A(n34012), .B(n33974), .Z(n33977) );
  XOR U33486 ( .A(n34013), .B(n34014), .Z(n33974) );
  AND U33487 ( .A(n34015), .B(n34016), .Z(n34014) );
  XOR U33488 ( .A(n34013), .B(n34017), .Z(n34015) );
  XNOR U33489 ( .A(n34018), .B(n34019), .Z(n34012) );
  NOR U33490 ( .A(n34020), .B(n34021), .Z(n34019) );
  XNOR U33491 ( .A(n34018), .B(n34022), .Z(n34020) );
  XOR U33492 ( .A(n34023), .B(n34024), .Z(n33978) );
  NOR U33493 ( .A(n34025), .B(n34026), .Z(n34024) );
  XNOR U33494 ( .A(n34023), .B(n34027), .Z(n34025) );
  XNOR U33495 ( .A(n33919), .B(n33984), .Z(n33986) );
  XNOR U33496 ( .A(n34028), .B(n34029), .Z(n33919) );
  AND U33497 ( .A(n493), .B(n34030), .Z(n34029) );
  XNOR U33498 ( .A(n34031), .B(n34032), .Z(n34030) );
  AND U33499 ( .A(n33925), .B(n33928), .Z(n33984) );
  XOR U33500 ( .A(n34033), .B(n34011), .Z(n33928) );
  XNOR U33501 ( .A(p_input[2048]), .B(p_input[352]), .Z(n34011) );
  XOR U33502 ( .A(n33999), .B(n33998), .Z(n34033) );
  XNOR U33503 ( .A(n34034), .B(n34005), .Z(n33998) );
  XNOR U33504 ( .A(n33994), .B(n33993), .Z(n34005) );
  XOR U33505 ( .A(n34035), .B(n33990), .Z(n33993) );
  XNOR U33506 ( .A(n29266), .B(p_input[362]), .Z(n33990) );
  XNOR U33507 ( .A(p_input[2059]), .B(p_input[363]), .Z(n34035) );
  XOR U33508 ( .A(p_input[2060]), .B(p_input[364]), .Z(n33994) );
  XNOR U33509 ( .A(n34004), .B(n33995), .Z(n34034) );
  XNOR U33510 ( .A(n29494), .B(p_input[353]), .Z(n33995) );
  XOR U33511 ( .A(n34036), .B(n34010), .Z(n34004) );
  XNOR U33512 ( .A(p_input[2063]), .B(p_input[367]), .Z(n34010) );
  XOR U33513 ( .A(n34001), .B(n34009), .Z(n34036) );
  XOR U33514 ( .A(n34037), .B(n34006), .Z(n34009) );
  XOR U33515 ( .A(p_input[2061]), .B(p_input[365]), .Z(n34006) );
  XNOR U33516 ( .A(p_input[2062]), .B(p_input[366]), .Z(n34037) );
  XNOR U33517 ( .A(n29036), .B(p_input[361]), .Z(n34001) );
  XNOR U33518 ( .A(n34017), .B(n34016), .Z(n33999) );
  XNOR U33519 ( .A(n34038), .B(n34022), .Z(n34016) );
  XOR U33520 ( .A(p_input[2056]), .B(p_input[360]), .Z(n34022) );
  XOR U33521 ( .A(n34013), .B(n34021), .Z(n34038) );
  XOR U33522 ( .A(n34039), .B(n34018), .Z(n34021) );
  XOR U33523 ( .A(p_input[2054]), .B(p_input[358]), .Z(n34018) );
  XNOR U33524 ( .A(p_input[2055]), .B(p_input[359]), .Z(n34039) );
  XNOR U33525 ( .A(n29039), .B(p_input[354]), .Z(n34013) );
  XNOR U33526 ( .A(n34027), .B(n34026), .Z(n34017) );
  XOR U33527 ( .A(n34040), .B(n34023), .Z(n34026) );
  XOR U33528 ( .A(p_input[2051]), .B(p_input[355]), .Z(n34023) );
  XNOR U33529 ( .A(p_input[2052]), .B(p_input[356]), .Z(n34040) );
  XOR U33530 ( .A(p_input[2053]), .B(p_input[357]), .Z(n34027) );
  XNOR U33531 ( .A(n34041), .B(n34042), .Z(n33925) );
  AND U33532 ( .A(n493), .B(n34043), .Z(n34042) );
  XNOR U33533 ( .A(n34044), .B(n34045), .Z(n493) );
  AND U33534 ( .A(n34046), .B(n34047), .Z(n34045) );
  XOR U33535 ( .A(n33939), .B(n34044), .Z(n34047) );
  XNOR U33536 ( .A(n34048), .B(n34044), .Z(n34046) );
  XOR U33537 ( .A(n34049), .B(n34050), .Z(n34044) );
  AND U33538 ( .A(n34051), .B(n34052), .Z(n34050) );
  XOR U33539 ( .A(n33954), .B(n34049), .Z(n34052) );
  XOR U33540 ( .A(n34049), .B(n33955), .Z(n34051) );
  XOR U33541 ( .A(n34053), .B(n34054), .Z(n34049) );
  AND U33542 ( .A(n34055), .B(n34056), .Z(n34054) );
  XOR U33543 ( .A(n33982), .B(n34053), .Z(n34056) );
  XOR U33544 ( .A(n34053), .B(n33983), .Z(n34055) );
  XOR U33545 ( .A(n34057), .B(n34058), .Z(n34053) );
  AND U33546 ( .A(n34059), .B(n34060), .Z(n34058) );
  XOR U33547 ( .A(n34057), .B(n34031), .Z(n34060) );
  XNOR U33548 ( .A(n34061), .B(n34062), .Z(n33885) );
  AND U33549 ( .A(n497), .B(n34063), .Z(n34062) );
  XNOR U33550 ( .A(n34064), .B(n34065), .Z(n497) );
  AND U33551 ( .A(n34066), .B(n34067), .Z(n34065) );
  XOR U33552 ( .A(n34064), .B(n33895), .Z(n34067) );
  XNOR U33553 ( .A(n34064), .B(n33855), .Z(n34066) );
  XOR U33554 ( .A(n34068), .B(n34069), .Z(n34064) );
  AND U33555 ( .A(n34070), .B(n34071), .Z(n34069) );
  XOR U33556 ( .A(n34068), .B(n33863), .Z(n34070) );
  XOR U33557 ( .A(n34072), .B(n34073), .Z(n33846) );
  AND U33558 ( .A(n501), .B(n34063), .Z(n34073) );
  XNOR U33559 ( .A(n34061), .B(n34072), .Z(n34063) );
  XNOR U33560 ( .A(n34074), .B(n34075), .Z(n501) );
  AND U33561 ( .A(n34076), .B(n34077), .Z(n34075) );
  XNOR U33562 ( .A(n34078), .B(n34074), .Z(n34077) );
  IV U33563 ( .A(n33895), .Z(n34078) );
  XOR U33564 ( .A(n34048), .B(n34079), .Z(n33895) );
  AND U33565 ( .A(n504), .B(n34080), .Z(n34079) );
  XOR U33566 ( .A(n33938), .B(n33935), .Z(n34080) );
  IV U33567 ( .A(n34048), .Z(n33938) );
  XNOR U33568 ( .A(n33855), .B(n34074), .Z(n34076) );
  XOR U33569 ( .A(n34081), .B(n34082), .Z(n33855) );
  AND U33570 ( .A(n520), .B(n34083), .Z(n34082) );
  XOR U33571 ( .A(n34068), .B(n34084), .Z(n34074) );
  AND U33572 ( .A(n34085), .B(n34071), .Z(n34084) );
  XNOR U33573 ( .A(n33905), .B(n34068), .Z(n34071) );
  XOR U33574 ( .A(n33955), .B(n34086), .Z(n33905) );
  AND U33575 ( .A(n504), .B(n34087), .Z(n34086) );
  XOR U33576 ( .A(n33951), .B(n33955), .Z(n34087) );
  XNOR U33577 ( .A(n34088), .B(n34068), .Z(n34085) );
  IV U33578 ( .A(n33863), .Z(n34088) );
  XOR U33579 ( .A(n34089), .B(n34090), .Z(n33863) );
  AND U33580 ( .A(n520), .B(n34091), .Z(n34090) );
  XOR U33581 ( .A(n34092), .B(n34093), .Z(n34068) );
  AND U33582 ( .A(n34094), .B(n34095), .Z(n34093) );
  XNOR U33583 ( .A(n33915), .B(n34092), .Z(n34095) );
  XOR U33584 ( .A(n33983), .B(n34096), .Z(n33915) );
  AND U33585 ( .A(n504), .B(n34097), .Z(n34096) );
  XOR U33586 ( .A(n33979), .B(n33983), .Z(n34097) );
  XOR U33587 ( .A(n34092), .B(n33872), .Z(n34094) );
  XOR U33588 ( .A(n34098), .B(n34099), .Z(n33872) );
  AND U33589 ( .A(n520), .B(n34100), .Z(n34099) );
  XOR U33590 ( .A(n34101), .B(n34102), .Z(n34092) );
  AND U33591 ( .A(n34103), .B(n34104), .Z(n34102) );
  XNOR U33592 ( .A(n34101), .B(n33923), .Z(n34104) );
  XOR U33593 ( .A(n34032), .B(n34105), .Z(n33923) );
  AND U33594 ( .A(n504), .B(n34106), .Z(n34105) );
  XOR U33595 ( .A(n34028), .B(n34032), .Z(n34106) );
  XNOR U33596 ( .A(n34107), .B(n34101), .Z(n34103) );
  IV U33597 ( .A(n33882), .Z(n34107) );
  XOR U33598 ( .A(n34108), .B(n34109), .Z(n33882) );
  AND U33599 ( .A(n520), .B(n34110), .Z(n34109) );
  AND U33600 ( .A(n34072), .B(n34061), .Z(n34101) );
  XNOR U33601 ( .A(n34111), .B(n34112), .Z(n34061) );
  AND U33602 ( .A(n504), .B(n34043), .Z(n34112) );
  XNOR U33603 ( .A(n34041), .B(n34111), .Z(n34043) );
  XNOR U33604 ( .A(n34113), .B(n34114), .Z(n504) );
  AND U33605 ( .A(n34115), .B(n34116), .Z(n34114) );
  XNOR U33606 ( .A(n34113), .B(n33935), .Z(n34116) );
  IV U33607 ( .A(n33939), .Z(n33935) );
  XOR U33608 ( .A(n34117), .B(n34118), .Z(n33939) );
  AND U33609 ( .A(n508), .B(n34119), .Z(n34118) );
  XOR U33610 ( .A(n34120), .B(n34117), .Z(n34119) );
  XNOR U33611 ( .A(n34113), .B(n34048), .Z(n34115) );
  XOR U33612 ( .A(n34121), .B(n34122), .Z(n34048) );
  AND U33613 ( .A(n516), .B(n34083), .Z(n34122) );
  XOR U33614 ( .A(n34081), .B(n34121), .Z(n34083) );
  XOR U33615 ( .A(n34123), .B(n34124), .Z(n34113) );
  AND U33616 ( .A(n34125), .B(n34126), .Z(n34124) );
  XNOR U33617 ( .A(n34123), .B(n33951), .Z(n34126) );
  IV U33618 ( .A(n33954), .Z(n33951) );
  XOR U33619 ( .A(n34127), .B(n34128), .Z(n33954) );
  AND U33620 ( .A(n508), .B(n34129), .Z(n34128) );
  XOR U33621 ( .A(n34130), .B(n34127), .Z(n34129) );
  XOR U33622 ( .A(n33955), .B(n34123), .Z(n34125) );
  XOR U33623 ( .A(n34131), .B(n34132), .Z(n33955) );
  AND U33624 ( .A(n516), .B(n34091), .Z(n34132) );
  XOR U33625 ( .A(n34131), .B(n34089), .Z(n34091) );
  XOR U33626 ( .A(n34133), .B(n34134), .Z(n34123) );
  AND U33627 ( .A(n34135), .B(n34136), .Z(n34134) );
  XNOR U33628 ( .A(n34133), .B(n33979), .Z(n34136) );
  IV U33629 ( .A(n33982), .Z(n33979) );
  XOR U33630 ( .A(n34137), .B(n34138), .Z(n33982) );
  AND U33631 ( .A(n508), .B(n34139), .Z(n34138) );
  XNOR U33632 ( .A(n34140), .B(n34137), .Z(n34139) );
  XOR U33633 ( .A(n33983), .B(n34133), .Z(n34135) );
  XOR U33634 ( .A(n34141), .B(n34142), .Z(n33983) );
  AND U33635 ( .A(n516), .B(n34100), .Z(n34142) );
  XOR U33636 ( .A(n34141), .B(n34098), .Z(n34100) );
  XOR U33637 ( .A(n34057), .B(n34143), .Z(n34133) );
  AND U33638 ( .A(n34059), .B(n34144), .Z(n34143) );
  XNOR U33639 ( .A(n34057), .B(n34028), .Z(n34144) );
  IV U33640 ( .A(n34031), .Z(n34028) );
  XOR U33641 ( .A(n34145), .B(n34146), .Z(n34031) );
  AND U33642 ( .A(n508), .B(n34147), .Z(n34146) );
  XOR U33643 ( .A(n34148), .B(n34145), .Z(n34147) );
  XOR U33644 ( .A(n34032), .B(n34057), .Z(n34059) );
  XOR U33645 ( .A(n34149), .B(n34150), .Z(n34032) );
  AND U33646 ( .A(n516), .B(n34110), .Z(n34150) );
  XOR U33647 ( .A(n34149), .B(n34108), .Z(n34110) );
  AND U33648 ( .A(n34111), .B(n34041), .Z(n34057) );
  XNOR U33649 ( .A(n34151), .B(n34152), .Z(n34041) );
  AND U33650 ( .A(n508), .B(n34153), .Z(n34152) );
  XNOR U33651 ( .A(n34154), .B(n34151), .Z(n34153) );
  XNOR U33652 ( .A(n34155), .B(n34156), .Z(n508) );
  AND U33653 ( .A(n34157), .B(n34158), .Z(n34156) );
  XOR U33654 ( .A(n34120), .B(n34155), .Z(n34158) );
  AND U33655 ( .A(n34159), .B(n34160), .Z(n34120) );
  XNOR U33656 ( .A(n34117), .B(n34155), .Z(n34157) );
  XNOR U33657 ( .A(n34161), .B(n34162), .Z(n34117) );
  AND U33658 ( .A(n512), .B(n34163), .Z(n34162) );
  XNOR U33659 ( .A(n34164), .B(n34165), .Z(n34163) );
  XOR U33660 ( .A(n34166), .B(n34167), .Z(n34155) );
  AND U33661 ( .A(n34168), .B(n34169), .Z(n34167) );
  XNOR U33662 ( .A(n34166), .B(n34159), .Z(n34169) );
  IV U33663 ( .A(n34130), .Z(n34159) );
  XOR U33664 ( .A(n34170), .B(n34171), .Z(n34130) );
  XOR U33665 ( .A(n34172), .B(n34160), .Z(n34171) );
  AND U33666 ( .A(n34140), .B(n34173), .Z(n34160) );
  AND U33667 ( .A(n34174), .B(n34175), .Z(n34172) );
  XOR U33668 ( .A(n34176), .B(n34170), .Z(n34174) );
  XNOR U33669 ( .A(n34127), .B(n34166), .Z(n34168) );
  XNOR U33670 ( .A(n34177), .B(n34178), .Z(n34127) );
  AND U33671 ( .A(n512), .B(n34179), .Z(n34178) );
  XNOR U33672 ( .A(n34180), .B(n34181), .Z(n34179) );
  XOR U33673 ( .A(n34182), .B(n34183), .Z(n34166) );
  AND U33674 ( .A(n34184), .B(n34185), .Z(n34183) );
  XNOR U33675 ( .A(n34182), .B(n34140), .Z(n34185) );
  XOR U33676 ( .A(n34186), .B(n34175), .Z(n34140) );
  XNOR U33677 ( .A(n34187), .B(n34170), .Z(n34175) );
  XOR U33678 ( .A(n34188), .B(n34189), .Z(n34170) );
  AND U33679 ( .A(n34190), .B(n34191), .Z(n34189) );
  XOR U33680 ( .A(n34192), .B(n34188), .Z(n34190) );
  XNOR U33681 ( .A(n34193), .B(n34194), .Z(n34187) );
  AND U33682 ( .A(n34195), .B(n34196), .Z(n34194) );
  XOR U33683 ( .A(n34193), .B(n34197), .Z(n34195) );
  XNOR U33684 ( .A(n34176), .B(n34173), .Z(n34186) );
  AND U33685 ( .A(n34198), .B(n34199), .Z(n34173) );
  XOR U33686 ( .A(n34200), .B(n34201), .Z(n34176) );
  AND U33687 ( .A(n34202), .B(n34203), .Z(n34201) );
  XOR U33688 ( .A(n34200), .B(n34204), .Z(n34202) );
  XNOR U33689 ( .A(n34137), .B(n34182), .Z(n34184) );
  XNOR U33690 ( .A(n34205), .B(n34206), .Z(n34137) );
  AND U33691 ( .A(n512), .B(n34207), .Z(n34206) );
  XNOR U33692 ( .A(n34208), .B(n34209), .Z(n34207) );
  XOR U33693 ( .A(n34210), .B(n34211), .Z(n34182) );
  AND U33694 ( .A(n34212), .B(n34213), .Z(n34211) );
  XNOR U33695 ( .A(n34210), .B(n34198), .Z(n34213) );
  IV U33696 ( .A(n34148), .Z(n34198) );
  XNOR U33697 ( .A(n34214), .B(n34191), .Z(n34148) );
  XNOR U33698 ( .A(n34215), .B(n34197), .Z(n34191) );
  XOR U33699 ( .A(n34216), .B(n34217), .Z(n34197) );
  NOR U33700 ( .A(n34218), .B(n34219), .Z(n34217) );
  XNOR U33701 ( .A(n34216), .B(n34220), .Z(n34218) );
  XNOR U33702 ( .A(n34196), .B(n34188), .Z(n34215) );
  XOR U33703 ( .A(n34221), .B(n34222), .Z(n34188) );
  AND U33704 ( .A(n34223), .B(n34224), .Z(n34222) );
  XNOR U33705 ( .A(n34221), .B(n34225), .Z(n34223) );
  XNOR U33706 ( .A(n34226), .B(n34193), .Z(n34196) );
  XOR U33707 ( .A(n34227), .B(n34228), .Z(n34193) );
  AND U33708 ( .A(n34229), .B(n34230), .Z(n34228) );
  XOR U33709 ( .A(n34227), .B(n34231), .Z(n34229) );
  XNOR U33710 ( .A(n34232), .B(n34233), .Z(n34226) );
  NOR U33711 ( .A(n34234), .B(n34235), .Z(n34233) );
  XOR U33712 ( .A(n34232), .B(n34236), .Z(n34234) );
  XNOR U33713 ( .A(n34192), .B(n34199), .Z(n34214) );
  NOR U33714 ( .A(n34154), .B(n34237), .Z(n34199) );
  XOR U33715 ( .A(n34204), .B(n34203), .Z(n34192) );
  XNOR U33716 ( .A(n34238), .B(n34200), .Z(n34203) );
  XOR U33717 ( .A(n34239), .B(n34240), .Z(n34200) );
  AND U33718 ( .A(n34241), .B(n34242), .Z(n34240) );
  XOR U33719 ( .A(n34239), .B(n34243), .Z(n34241) );
  XNOR U33720 ( .A(n34244), .B(n34245), .Z(n34238) );
  NOR U33721 ( .A(n34246), .B(n34247), .Z(n34245) );
  XNOR U33722 ( .A(n34244), .B(n34248), .Z(n34246) );
  XOR U33723 ( .A(n34249), .B(n34250), .Z(n34204) );
  NOR U33724 ( .A(n34251), .B(n34252), .Z(n34250) );
  XNOR U33725 ( .A(n34249), .B(n34253), .Z(n34251) );
  XNOR U33726 ( .A(n34145), .B(n34210), .Z(n34212) );
  XNOR U33727 ( .A(n34254), .B(n34255), .Z(n34145) );
  AND U33728 ( .A(n512), .B(n34256), .Z(n34255) );
  XNOR U33729 ( .A(n34257), .B(n34258), .Z(n34256) );
  AND U33730 ( .A(n34151), .B(n34154), .Z(n34210) );
  XOR U33731 ( .A(n34259), .B(n34237), .Z(n34154) );
  XNOR U33732 ( .A(p_input[2048]), .B(p_input[368]), .Z(n34237) );
  XOR U33733 ( .A(n34225), .B(n34224), .Z(n34259) );
  XNOR U33734 ( .A(n34260), .B(n34231), .Z(n34224) );
  XNOR U33735 ( .A(n34220), .B(n34219), .Z(n34231) );
  XOR U33736 ( .A(n34261), .B(n34216), .Z(n34219) );
  XNOR U33737 ( .A(n29266), .B(p_input[378]), .Z(n34216) );
  XNOR U33738 ( .A(p_input[2059]), .B(p_input[379]), .Z(n34261) );
  XOR U33739 ( .A(p_input[2060]), .B(p_input[380]), .Z(n34220) );
  XNOR U33740 ( .A(n34230), .B(n34221), .Z(n34260) );
  XNOR U33741 ( .A(n29494), .B(p_input[369]), .Z(n34221) );
  XOR U33742 ( .A(n34262), .B(n34236), .Z(n34230) );
  XNOR U33743 ( .A(p_input[2063]), .B(p_input[383]), .Z(n34236) );
  XOR U33744 ( .A(n34227), .B(n34235), .Z(n34262) );
  XOR U33745 ( .A(n34263), .B(n34232), .Z(n34235) );
  XOR U33746 ( .A(p_input[2061]), .B(p_input[381]), .Z(n34232) );
  XNOR U33747 ( .A(p_input[2062]), .B(p_input[382]), .Z(n34263) );
  XNOR U33748 ( .A(n29036), .B(p_input[377]), .Z(n34227) );
  XNOR U33749 ( .A(n34243), .B(n34242), .Z(n34225) );
  XNOR U33750 ( .A(n34264), .B(n34248), .Z(n34242) );
  XOR U33751 ( .A(p_input[2056]), .B(p_input[376]), .Z(n34248) );
  XOR U33752 ( .A(n34239), .B(n34247), .Z(n34264) );
  XOR U33753 ( .A(n34265), .B(n34244), .Z(n34247) );
  XOR U33754 ( .A(p_input[2054]), .B(p_input[374]), .Z(n34244) );
  XNOR U33755 ( .A(p_input[2055]), .B(p_input[375]), .Z(n34265) );
  XNOR U33756 ( .A(n29039), .B(p_input[370]), .Z(n34239) );
  XNOR U33757 ( .A(n34253), .B(n34252), .Z(n34243) );
  XOR U33758 ( .A(n34266), .B(n34249), .Z(n34252) );
  XOR U33759 ( .A(p_input[2051]), .B(p_input[371]), .Z(n34249) );
  XNOR U33760 ( .A(p_input[2052]), .B(p_input[372]), .Z(n34266) );
  XOR U33761 ( .A(p_input[2053]), .B(p_input[373]), .Z(n34253) );
  XNOR U33762 ( .A(n34267), .B(n34268), .Z(n34151) );
  AND U33763 ( .A(n512), .B(n34269), .Z(n34268) );
  XNOR U33764 ( .A(n34270), .B(n34271), .Z(n512) );
  AND U33765 ( .A(n34272), .B(n34273), .Z(n34271) );
  XOR U33766 ( .A(n34165), .B(n34270), .Z(n34273) );
  XNOR U33767 ( .A(n34274), .B(n34270), .Z(n34272) );
  XOR U33768 ( .A(n34275), .B(n34276), .Z(n34270) );
  AND U33769 ( .A(n34277), .B(n34278), .Z(n34276) );
  XOR U33770 ( .A(n34180), .B(n34275), .Z(n34278) );
  XOR U33771 ( .A(n34275), .B(n34181), .Z(n34277) );
  XOR U33772 ( .A(n34279), .B(n34280), .Z(n34275) );
  AND U33773 ( .A(n34281), .B(n34282), .Z(n34280) );
  XOR U33774 ( .A(n34208), .B(n34279), .Z(n34282) );
  XOR U33775 ( .A(n34279), .B(n34209), .Z(n34281) );
  XOR U33776 ( .A(n34283), .B(n34284), .Z(n34279) );
  AND U33777 ( .A(n34285), .B(n34286), .Z(n34284) );
  XOR U33778 ( .A(n34283), .B(n34257), .Z(n34286) );
  XNOR U33779 ( .A(n34287), .B(n34288), .Z(n34111) );
  AND U33780 ( .A(n516), .B(n34289), .Z(n34288) );
  XNOR U33781 ( .A(n34290), .B(n34291), .Z(n516) );
  AND U33782 ( .A(n34292), .B(n34293), .Z(n34291) );
  XOR U33783 ( .A(n34290), .B(n34121), .Z(n34293) );
  XNOR U33784 ( .A(n34290), .B(n34081), .Z(n34292) );
  XOR U33785 ( .A(n34294), .B(n34295), .Z(n34290) );
  AND U33786 ( .A(n34296), .B(n34297), .Z(n34295) );
  XOR U33787 ( .A(n34294), .B(n34089), .Z(n34296) );
  XOR U33788 ( .A(n34298), .B(n34299), .Z(n34072) );
  AND U33789 ( .A(n520), .B(n34289), .Z(n34299) );
  XNOR U33790 ( .A(n34287), .B(n34298), .Z(n34289) );
  XNOR U33791 ( .A(n34300), .B(n34301), .Z(n520) );
  AND U33792 ( .A(n34302), .B(n34303), .Z(n34301) );
  XNOR U33793 ( .A(n34304), .B(n34300), .Z(n34303) );
  IV U33794 ( .A(n34121), .Z(n34304) );
  XOR U33795 ( .A(n34274), .B(n34305), .Z(n34121) );
  AND U33796 ( .A(n523), .B(n34306), .Z(n34305) );
  XOR U33797 ( .A(n34164), .B(n34161), .Z(n34306) );
  IV U33798 ( .A(n34274), .Z(n34164) );
  XNOR U33799 ( .A(n34081), .B(n34300), .Z(n34302) );
  XOR U33800 ( .A(n34307), .B(n34308), .Z(n34081) );
  AND U33801 ( .A(n539), .B(n34309), .Z(n34308) );
  XOR U33802 ( .A(n34294), .B(n34310), .Z(n34300) );
  AND U33803 ( .A(n34311), .B(n34297), .Z(n34310) );
  XNOR U33804 ( .A(n34131), .B(n34294), .Z(n34297) );
  XOR U33805 ( .A(n34181), .B(n34312), .Z(n34131) );
  AND U33806 ( .A(n523), .B(n34313), .Z(n34312) );
  XOR U33807 ( .A(n34177), .B(n34181), .Z(n34313) );
  XNOR U33808 ( .A(n34314), .B(n34294), .Z(n34311) );
  IV U33809 ( .A(n34089), .Z(n34314) );
  XOR U33810 ( .A(n34315), .B(n34316), .Z(n34089) );
  AND U33811 ( .A(n539), .B(n34317), .Z(n34316) );
  XOR U33812 ( .A(n34318), .B(n34319), .Z(n34294) );
  AND U33813 ( .A(n34320), .B(n34321), .Z(n34319) );
  XNOR U33814 ( .A(n34141), .B(n34318), .Z(n34321) );
  XOR U33815 ( .A(n34209), .B(n34322), .Z(n34141) );
  AND U33816 ( .A(n523), .B(n34323), .Z(n34322) );
  XOR U33817 ( .A(n34205), .B(n34209), .Z(n34323) );
  XOR U33818 ( .A(n34318), .B(n34098), .Z(n34320) );
  XOR U33819 ( .A(n34324), .B(n34325), .Z(n34098) );
  AND U33820 ( .A(n539), .B(n34326), .Z(n34325) );
  XOR U33821 ( .A(n34327), .B(n34328), .Z(n34318) );
  AND U33822 ( .A(n34329), .B(n34330), .Z(n34328) );
  XNOR U33823 ( .A(n34327), .B(n34149), .Z(n34330) );
  XOR U33824 ( .A(n34258), .B(n34331), .Z(n34149) );
  AND U33825 ( .A(n523), .B(n34332), .Z(n34331) );
  XOR U33826 ( .A(n34254), .B(n34258), .Z(n34332) );
  XNOR U33827 ( .A(n34333), .B(n34327), .Z(n34329) );
  IV U33828 ( .A(n34108), .Z(n34333) );
  XOR U33829 ( .A(n34334), .B(n34335), .Z(n34108) );
  AND U33830 ( .A(n539), .B(n34336), .Z(n34335) );
  AND U33831 ( .A(n34298), .B(n34287), .Z(n34327) );
  XNOR U33832 ( .A(n34337), .B(n34338), .Z(n34287) );
  AND U33833 ( .A(n523), .B(n34269), .Z(n34338) );
  XNOR U33834 ( .A(n34267), .B(n34337), .Z(n34269) );
  XNOR U33835 ( .A(n34339), .B(n34340), .Z(n523) );
  AND U33836 ( .A(n34341), .B(n34342), .Z(n34340) );
  XNOR U33837 ( .A(n34339), .B(n34161), .Z(n34342) );
  IV U33838 ( .A(n34165), .Z(n34161) );
  XOR U33839 ( .A(n34343), .B(n34344), .Z(n34165) );
  AND U33840 ( .A(n527), .B(n34345), .Z(n34344) );
  XOR U33841 ( .A(n34346), .B(n34343), .Z(n34345) );
  XNOR U33842 ( .A(n34339), .B(n34274), .Z(n34341) );
  XOR U33843 ( .A(n34347), .B(n34348), .Z(n34274) );
  AND U33844 ( .A(n535), .B(n34309), .Z(n34348) );
  XOR U33845 ( .A(n34307), .B(n34347), .Z(n34309) );
  XOR U33846 ( .A(n34349), .B(n34350), .Z(n34339) );
  AND U33847 ( .A(n34351), .B(n34352), .Z(n34350) );
  XNOR U33848 ( .A(n34349), .B(n34177), .Z(n34352) );
  IV U33849 ( .A(n34180), .Z(n34177) );
  XOR U33850 ( .A(n34353), .B(n34354), .Z(n34180) );
  AND U33851 ( .A(n527), .B(n34355), .Z(n34354) );
  XOR U33852 ( .A(n34356), .B(n34353), .Z(n34355) );
  XOR U33853 ( .A(n34181), .B(n34349), .Z(n34351) );
  XOR U33854 ( .A(n34357), .B(n34358), .Z(n34181) );
  AND U33855 ( .A(n535), .B(n34317), .Z(n34358) );
  XOR U33856 ( .A(n34357), .B(n34315), .Z(n34317) );
  XOR U33857 ( .A(n34359), .B(n34360), .Z(n34349) );
  AND U33858 ( .A(n34361), .B(n34362), .Z(n34360) );
  XNOR U33859 ( .A(n34359), .B(n34205), .Z(n34362) );
  IV U33860 ( .A(n34208), .Z(n34205) );
  XOR U33861 ( .A(n34363), .B(n34364), .Z(n34208) );
  AND U33862 ( .A(n527), .B(n34365), .Z(n34364) );
  XNOR U33863 ( .A(n34366), .B(n34363), .Z(n34365) );
  XOR U33864 ( .A(n34209), .B(n34359), .Z(n34361) );
  XOR U33865 ( .A(n34367), .B(n34368), .Z(n34209) );
  AND U33866 ( .A(n535), .B(n34326), .Z(n34368) );
  XOR U33867 ( .A(n34367), .B(n34324), .Z(n34326) );
  XOR U33868 ( .A(n34283), .B(n34369), .Z(n34359) );
  AND U33869 ( .A(n34285), .B(n34370), .Z(n34369) );
  XNOR U33870 ( .A(n34283), .B(n34254), .Z(n34370) );
  IV U33871 ( .A(n34257), .Z(n34254) );
  XOR U33872 ( .A(n34371), .B(n34372), .Z(n34257) );
  AND U33873 ( .A(n527), .B(n34373), .Z(n34372) );
  XOR U33874 ( .A(n34374), .B(n34371), .Z(n34373) );
  XOR U33875 ( .A(n34258), .B(n34283), .Z(n34285) );
  XOR U33876 ( .A(n34375), .B(n34376), .Z(n34258) );
  AND U33877 ( .A(n535), .B(n34336), .Z(n34376) );
  XOR U33878 ( .A(n34375), .B(n34334), .Z(n34336) );
  AND U33879 ( .A(n34337), .B(n34267), .Z(n34283) );
  XNOR U33880 ( .A(n34377), .B(n34378), .Z(n34267) );
  AND U33881 ( .A(n527), .B(n34379), .Z(n34378) );
  XNOR U33882 ( .A(n34380), .B(n34377), .Z(n34379) );
  XNOR U33883 ( .A(n34381), .B(n34382), .Z(n527) );
  AND U33884 ( .A(n34383), .B(n34384), .Z(n34382) );
  XOR U33885 ( .A(n34346), .B(n34381), .Z(n34384) );
  AND U33886 ( .A(n34385), .B(n34386), .Z(n34346) );
  XNOR U33887 ( .A(n34343), .B(n34381), .Z(n34383) );
  XNOR U33888 ( .A(n34387), .B(n34388), .Z(n34343) );
  AND U33889 ( .A(n531), .B(n34389), .Z(n34388) );
  XNOR U33890 ( .A(n34390), .B(n34391), .Z(n34389) );
  XOR U33891 ( .A(n34392), .B(n34393), .Z(n34381) );
  AND U33892 ( .A(n34394), .B(n34395), .Z(n34393) );
  XNOR U33893 ( .A(n34392), .B(n34385), .Z(n34395) );
  IV U33894 ( .A(n34356), .Z(n34385) );
  XOR U33895 ( .A(n34396), .B(n34397), .Z(n34356) );
  XOR U33896 ( .A(n34398), .B(n34386), .Z(n34397) );
  AND U33897 ( .A(n34366), .B(n34399), .Z(n34386) );
  AND U33898 ( .A(n34400), .B(n34401), .Z(n34398) );
  XOR U33899 ( .A(n34402), .B(n34396), .Z(n34400) );
  XNOR U33900 ( .A(n34353), .B(n34392), .Z(n34394) );
  XNOR U33901 ( .A(n34403), .B(n34404), .Z(n34353) );
  AND U33902 ( .A(n531), .B(n34405), .Z(n34404) );
  XNOR U33903 ( .A(n34406), .B(n34407), .Z(n34405) );
  XOR U33904 ( .A(n34408), .B(n34409), .Z(n34392) );
  AND U33905 ( .A(n34410), .B(n34411), .Z(n34409) );
  XNOR U33906 ( .A(n34408), .B(n34366), .Z(n34411) );
  XOR U33907 ( .A(n34412), .B(n34401), .Z(n34366) );
  XNOR U33908 ( .A(n34413), .B(n34396), .Z(n34401) );
  XOR U33909 ( .A(n34414), .B(n34415), .Z(n34396) );
  AND U33910 ( .A(n34416), .B(n34417), .Z(n34415) );
  XOR U33911 ( .A(n34418), .B(n34414), .Z(n34416) );
  XNOR U33912 ( .A(n34419), .B(n34420), .Z(n34413) );
  AND U33913 ( .A(n34421), .B(n34422), .Z(n34420) );
  XOR U33914 ( .A(n34419), .B(n34423), .Z(n34421) );
  XNOR U33915 ( .A(n34402), .B(n34399), .Z(n34412) );
  AND U33916 ( .A(n34424), .B(n34425), .Z(n34399) );
  XOR U33917 ( .A(n34426), .B(n34427), .Z(n34402) );
  AND U33918 ( .A(n34428), .B(n34429), .Z(n34427) );
  XOR U33919 ( .A(n34426), .B(n34430), .Z(n34428) );
  XNOR U33920 ( .A(n34363), .B(n34408), .Z(n34410) );
  XNOR U33921 ( .A(n34431), .B(n34432), .Z(n34363) );
  AND U33922 ( .A(n531), .B(n34433), .Z(n34432) );
  XNOR U33923 ( .A(n34434), .B(n34435), .Z(n34433) );
  XOR U33924 ( .A(n34436), .B(n34437), .Z(n34408) );
  AND U33925 ( .A(n34438), .B(n34439), .Z(n34437) );
  XNOR U33926 ( .A(n34436), .B(n34424), .Z(n34439) );
  IV U33927 ( .A(n34374), .Z(n34424) );
  XNOR U33928 ( .A(n34440), .B(n34417), .Z(n34374) );
  XNOR U33929 ( .A(n34441), .B(n34423), .Z(n34417) );
  XOR U33930 ( .A(n34442), .B(n34443), .Z(n34423) );
  NOR U33931 ( .A(n34444), .B(n34445), .Z(n34443) );
  XNOR U33932 ( .A(n34442), .B(n34446), .Z(n34444) );
  XNOR U33933 ( .A(n34422), .B(n34414), .Z(n34441) );
  XOR U33934 ( .A(n34447), .B(n34448), .Z(n34414) );
  AND U33935 ( .A(n34449), .B(n34450), .Z(n34448) );
  XNOR U33936 ( .A(n34447), .B(n34451), .Z(n34449) );
  XNOR U33937 ( .A(n34452), .B(n34419), .Z(n34422) );
  XOR U33938 ( .A(n34453), .B(n34454), .Z(n34419) );
  AND U33939 ( .A(n34455), .B(n34456), .Z(n34454) );
  XOR U33940 ( .A(n34453), .B(n34457), .Z(n34455) );
  XNOR U33941 ( .A(n34458), .B(n34459), .Z(n34452) );
  NOR U33942 ( .A(n34460), .B(n34461), .Z(n34459) );
  XOR U33943 ( .A(n34458), .B(n34462), .Z(n34460) );
  XNOR U33944 ( .A(n34418), .B(n34425), .Z(n34440) );
  NOR U33945 ( .A(n34380), .B(n34463), .Z(n34425) );
  XOR U33946 ( .A(n34430), .B(n34429), .Z(n34418) );
  XNOR U33947 ( .A(n34464), .B(n34426), .Z(n34429) );
  XOR U33948 ( .A(n34465), .B(n34466), .Z(n34426) );
  AND U33949 ( .A(n34467), .B(n34468), .Z(n34466) );
  XOR U33950 ( .A(n34465), .B(n34469), .Z(n34467) );
  XNOR U33951 ( .A(n34470), .B(n34471), .Z(n34464) );
  NOR U33952 ( .A(n34472), .B(n34473), .Z(n34471) );
  XNOR U33953 ( .A(n34470), .B(n34474), .Z(n34472) );
  XOR U33954 ( .A(n34475), .B(n34476), .Z(n34430) );
  NOR U33955 ( .A(n34477), .B(n34478), .Z(n34476) );
  XNOR U33956 ( .A(n34475), .B(n34479), .Z(n34477) );
  XNOR U33957 ( .A(n34371), .B(n34436), .Z(n34438) );
  XNOR U33958 ( .A(n34480), .B(n34481), .Z(n34371) );
  AND U33959 ( .A(n531), .B(n34482), .Z(n34481) );
  XNOR U33960 ( .A(n34483), .B(n34484), .Z(n34482) );
  AND U33961 ( .A(n34377), .B(n34380), .Z(n34436) );
  XOR U33962 ( .A(n34485), .B(n34463), .Z(n34380) );
  XNOR U33963 ( .A(p_input[2048]), .B(p_input[384]), .Z(n34463) );
  XOR U33964 ( .A(n34451), .B(n34450), .Z(n34485) );
  XNOR U33965 ( .A(n34486), .B(n34457), .Z(n34450) );
  XNOR U33966 ( .A(n34446), .B(n34445), .Z(n34457) );
  XOR U33967 ( .A(n34487), .B(n34442), .Z(n34445) );
  XNOR U33968 ( .A(n29266), .B(p_input[394]), .Z(n34442) );
  XNOR U33969 ( .A(p_input[2059]), .B(p_input[395]), .Z(n34487) );
  XOR U33970 ( .A(p_input[2060]), .B(p_input[396]), .Z(n34446) );
  XNOR U33971 ( .A(n34456), .B(n34447), .Z(n34486) );
  XNOR U33972 ( .A(n29494), .B(p_input[385]), .Z(n34447) );
  XOR U33973 ( .A(n34488), .B(n34462), .Z(n34456) );
  XNOR U33974 ( .A(p_input[2063]), .B(p_input[399]), .Z(n34462) );
  XOR U33975 ( .A(n34453), .B(n34461), .Z(n34488) );
  XOR U33976 ( .A(n34489), .B(n34458), .Z(n34461) );
  XOR U33977 ( .A(p_input[2061]), .B(p_input[397]), .Z(n34458) );
  XNOR U33978 ( .A(p_input[2062]), .B(p_input[398]), .Z(n34489) );
  XNOR U33979 ( .A(n29036), .B(p_input[393]), .Z(n34453) );
  XNOR U33980 ( .A(n34469), .B(n34468), .Z(n34451) );
  XNOR U33981 ( .A(n34490), .B(n34474), .Z(n34468) );
  XOR U33982 ( .A(p_input[2056]), .B(p_input[392]), .Z(n34474) );
  XOR U33983 ( .A(n34465), .B(n34473), .Z(n34490) );
  XOR U33984 ( .A(n34491), .B(n34470), .Z(n34473) );
  XOR U33985 ( .A(p_input[2054]), .B(p_input[390]), .Z(n34470) );
  XNOR U33986 ( .A(p_input[2055]), .B(p_input[391]), .Z(n34491) );
  XNOR U33987 ( .A(n29039), .B(p_input[386]), .Z(n34465) );
  XNOR U33988 ( .A(n34479), .B(n34478), .Z(n34469) );
  XOR U33989 ( .A(n34492), .B(n34475), .Z(n34478) );
  XOR U33990 ( .A(p_input[2051]), .B(p_input[387]), .Z(n34475) );
  XNOR U33991 ( .A(p_input[2052]), .B(p_input[388]), .Z(n34492) );
  XOR U33992 ( .A(p_input[2053]), .B(p_input[389]), .Z(n34479) );
  XNOR U33993 ( .A(n34493), .B(n34494), .Z(n34377) );
  AND U33994 ( .A(n531), .B(n34495), .Z(n34494) );
  XNOR U33995 ( .A(n34496), .B(n34497), .Z(n531) );
  AND U33996 ( .A(n34498), .B(n34499), .Z(n34497) );
  XOR U33997 ( .A(n34391), .B(n34496), .Z(n34499) );
  XNOR U33998 ( .A(n34500), .B(n34496), .Z(n34498) );
  XOR U33999 ( .A(n34501), .B(n34502), .Z(n34496) );
  AND U34000 ( .A(n34503), .B(n34504), .Z(n34502) );
  XOR U34001 ( .A(n34406), .B(n34501), .Z(n34504) );
  XOR U34002 ( .A(n34501), .B(n34407), .Z(n34503) );
  XOR U34003 ( .A(n34505), .B(n34506), .Z(n34501) );
  AND U34004 ( .A(n34507), .B(n34508), .Z(n34506) );
  XOR U34005 ( .A(n34434), .B(n34505), .Z(n34508) );
  XOR U34006 ( .A(n34505), .B(n34435), .Z(n34507) );
  XOR U34007 ( .A(n34509), .B(n34510), .Z(n34505) );
  AND U34008 ( .A(n34511), .B(n34512), .Z(n34510) );
  XOR U34009 ( .A(n34509), .B(n34483), .Z(n34512) );
  XNOR U34010 ( .A(n34513), .B(n34514), .Z(n34337) );
  AND U34011 ( .A(n535), .B(n34515), .Z(n34514) );
  XNOR U34012 ( .A(n34516), .B(n34517), .Z(n535) );
  AND U34013 ( .A(n34518), .B(n34519), .Z(n34517) );
  XOR U34014 ( .A(n34516), .B(n34347), .Z(n34519) );
  XNOR U34015 ( .A(n34516), .B(n34307), .Z(n34518) );
  XOR U34016 ( .A(n34520), .B(n34521), .Z(n34516) );
  AND U34017 ( .A(n34522), .B(n34523), .Z(n34521) );
  XOR U34018 ( .A(n34520), .B(n34315), .Z(n34522) );
  XOR U34019 ( .A(n34524), .B(n34525), .Z(n34298) );
  AND U34020 ( .A(n539), .B(n34515), .Z(n34525) );
  XNOR U34021 ( .A(n34513), .B(n34524), .Z(n34515) );
  XNOR U34022 ( .A(n34526), .B(n34527), .Z(n539) );
  AND U34023 ( .A(n34528), .B(n34529), .Z(n34527) );
  XNOR U34024 ( .A(n34530), .B(n34526), .Z(n34529) );
  IV U34025 ( .A(n34347), .Z(n34530) );
  XOR U34026 ( .A(n34500), .B(n34531), .Z(n34347) );
  AND U34027 ( .A(n542), .B(n34532), .Z(n34531) );
  XOR U34028 ( .A(n34390), .B(n34387), .Z(n34532) );
  IV U34029 ( .A(n34500), .Z(n34390) );
  XNOR U34030 ( .A(n34307), .B(n34526), .Z(n34528) );
  XOR U34031 ( .A(n34533), .B(n34534), .Z(n34307) );
  AND U34032 ( .A(n558), .B(n34535), .Z(n34534) );
  XOR U34033 ( .A(n34520), .B(n34536), .Z(n34526) );
  AND U34034 ( .A(n34537), .B(n34523), .Z(n34536) );
  XNOR U34035 ( .A(n34357), .B(n34520), .Z(n34523) );
  XOR U34036 ( .A(n34407), .B(n34538), .Z(n34357) );
  AND U34037 ( .A(n542), .B(n34539), .Z(n34538) );
  XOR U34038 ( .A(n34403), .B(n34407), .Z(n34539) );
  XNOR U34039 ( .A(n34540), .B(n34520), .Z(n34537) );
  IV U34040 ( .A(n34315), .Z(n34540) );
  XOR U34041 ( .A(n34541), .B(n34542), .Z(n34315) );
  AND U34042 ( .A(n558), .B(n34543), .Z(n34542) );
  XOR U34043 ( .A(n34544), .B(n34545), .Z(n34520) );
  AND U34044 ( .A(n34546), .B(n34547), .Z(n34545) );
  XNOR U34045 ( .A(n34367), .B(n34544), .Z(n34547) );
  XOR U34046 ( .A(n34435), .B(n34548), .Z(n34367) );
  AND U34047 ( .A(n542), .B(n34549), .Z(n34548) );
  XOR U34048 ( .A(n34431), .B(n34435), .Z(n34549) );
  XOR U34049 ( .A(n34544), .B(n34324), .Z(n34546) );
  XOR U34050 ( .A(n34550), .B(n34551), .Z(n34324) );
  AND U34051 ( .A(n558), .B(n34552), .Z(n34551) );
  XOR U34052 ( .A(n34553), .B(n34554), .Z(n34544) );
  AND U34053 ( .A(n34555), .B(n34556), .Z(n34554) );
  XNOR U34054 ( .A(n34553), .B(n34375), .Z(n34556) );
  XOR U34055 ( .A(n34484), .B(n34557), .Z(n34375) );
  AND U34056 ( .A(n542), .B(n34558), .Z(n34557) );
  XOR U34057 ( .A(n34480), .B(n34484), .Z(n34558) );
  XNOR U34058 ( .A(n34559), .B(n34553), .Z(n34555) );
  IV U34059 ( .A(n34334), .Z(n34559) );
  XOR U34060 ( .A(n34560), .B(n34561), .Z(n34334) );
  AND U34061 ( .A(n558), .B(n34562), .Z(n34561) );
  AND U34062 ( .A(n34524), .B(n34513), .Z(n34553) );
  XNOR U34063 ( .A(n34563), .B(n34564), .Z(n34513) );
  AND U34064 ( .A(n542), .B(n34495), .Z(n34564) );
  XNOR U34065 ( .A(n34493), .B(n34563), .Z(n34495) );
  XNOR U34066 ( .A(n34565), .B(n34566), .Z(n542) );
  AND U34067 ( .A(n34567), .B(n34568), .Z(n34566) );
  XNOR U34068 ( .A(n34565), .B(n34387), .Z(n34568) );
  IV U34069 ( .A(n34391), .Z(n34387) );
  XOR U34070 ( .A(n34569), .B(n34570), .Z(n34391) );
  AND U34071 ( .A(n546), .B(n34571), .Z(n34570) );
  XOR U34072 ( .A(n34572), .B(n34569), .Z(n34571) );
  XNOR U34073 ( .A(n34565), .B(n34500), .Z(n34567) );
  XOR U34074 ( .A(n34573), .B(n34574), .Z(n34500) );
  AND U34075 ( .A(n554), .B(n34535), .Z(n34574) );
  XOR U34076 ( .A(n34533), .B(n34573), .Z(n34535) );
  XOR U34077 ( .A(n34575), .B(n34576), .Z(n34565) );
  AND U34078 ( .A(n34577), .B(n34578), .Z(n34576) );
  XNOR U34079 ( .A(n34575), .B(n34403), .Z(n34578) );
  IV U34080 ( .A(n34406), .Z(n34403) );
  XOR U34081 ( .A(n34579), .B(n34580), .Z(n34406) );
  AND U34082 ( .A(n546), .B(n34581), .Z(n34580) );
  XOR U34083 ( .A(n34582), .B(n34579), .Z(n34581) );
  XOR U34084 ( .A(n34407), .B(n34575), .Z(n34577) );
  XOR U34085 ( .A(n34583), .B(n34584), .Z(n34407) );
  AND U34086 ( .A(n554), .B(n34543), .Z(n34584) );
  XOR U34087 ( .A(n34583), .B(n34541), .Z(n34543) );
  XOR U34088 ( .A(n34585), .B(n34586), .Z(n34575) );
  AND U34089 ( .A(n34587), .B(n34588), .Z(n34586) );
  XNOR U34090 ( .A(n34585), .B(n34431), .Z(n34588) );
  IV U34091 ( .A(n34434), .Z(n34431) );
  XOR U34092 ( .A(n34589), .B(n34590), .Z(n34434) );
  AND U34093 ( .A(n546), .B(n34591), .Z(n34590) );
  XNOR U34094 ( .A(n34592), .B(n34589), .Z(n34591) );
  XOR U34095 ( .A(n34435), .B(n34585), .Z(n34587) );
  XOR U34096 ( .A(n34593), .B(n34594), .Z(n34435) );
  AND U34097 ( .A(n554), .B(n34552), .Z(n34594) );
  XOR U34098 ( .A(n34593), .B(n34550), .Z(n34552) );
  XOR U34099 ( .A(n34509), .B(n34595), .Z(n34585) );
  AND U34100 ( .A(n34511), .B(n34596), .Z(n34595) );
  XNOR U34101 ( .A(n34509), .B(n34480), .Z(n34596) );
  IV U34102 ( .A(n34483), .Z(n34480) );
  XOR U34103 ( .A(n34597), .B(n34598), .Z(n34483) );
  AND U34104 ( .A(n546), .B(n34599), .Z(n34598) );
  XOR U34105 ( .A(n34600), .B(n34597), .Z(n34599) );
  XOR U34106 ( .A(n34484), .B(n34509), .Z(n34511) );
  XOR U34107 ( .A(n34601), .B(n34602), .Z(n34484) );
  AND U34108 ( .A(n554), .B(n34562), .Z(n34602) );
  XOR U34109 ( .A(n34601), .B(n34560), .Z(n34562) );
  AND U34110 ( .A(n34563), .B(n34493), .Z(n34509) );
  XNOR U34111 ( .A(n34603), .B(n34604), .Z(n34493) );
  AND U34112 ( .A(n546), .B(n34605), .Z(n34604) );
  XNOR U34113 ( .A(n34606), .B(n34603), .Z(n34605) );
  XNOR U34114 ( .A(n34607), .B(n34608), .Z(n546) );
  AND U34115 ( .A(n34609), .B(n34610), .Z(n34608) );
  XOR U34116 ( .A(n34572), .B(n34607), .Z(n34610) );
  AND U34117 ( .A(n34611), .B(n34612), .Z(n34572) );
  XNOR U34118 ( .A(n34569), .B(n34607), .Z(n34609) );
  XNOR U34119 ( .A(n34613), .B(n34614), .Z(n34569) );
  AND U34120 ( .A(n550), .B(n34615), .Z(n34614) );
  XNOR U34121 ( .A(n34616), .B(n34617), .Z(n34615) );
  XOR U34122 ( .A(n34618), .B(n34619), .Z(n34607) );
  AND U34123 ( .A(n34620), .B(n34621), .Z(n34619) );
  XNOR U34124 ( .A(n34618), .B(n34611), .Z(n34621) );
  IV U34125 ( .A(n34582), .Z(n34611) );
  XOR U34126 ( .A(n34622), .B(n34623), .Z(n34582) );
  XOR U34127 ( .A(n34624), .B(n34612), .Z(n34623) );
  AND U34128 ( .A(n34592), .B(n34625), .Z(n34612) );
  AND U34129 ( .A(n34626), .B(n34627), .Z(n34624) );
  XOR U34130 ( .A(n34628), .B(n34622), .Z(n34626) );
  XNOR U34131 ( .A(n34579), .B(n34618), .Z(n34620) );
  XNOR U34132 ( .A(n34629), .B(n34630), .Z(n34579) );
  AND U34133 ( .A(n550), .B(n34631), .Z(n34630) );
  XNOR U34134 ( .A(n34632), .B(n34633), .Z(n34631) );
  XOR U34135 ( .A(n34634), .B(n34635), .Z(n34618) );
  AND U34136 ( .A(n34636), .B(n34637), .Z(n34635) );
  XNOR U34137 ( .A(n34634), .B(n34592), .Z(n34637) );
  XOR U34138 ( .A(n34638), .B(n34627), .Z(n34592) );
  XNOR U34139 ( .A(n34639), .B(n34622), .Z(n34627) );
  XOR U34140 ( .A(n34640), .B(n34641), .Z(n34622) );
  AND U34141 ( .A(n34642), .B(n34643), .Z(n34641) );
  XOR U34142 ( .A(n34644), .B(n34640), .Z(n34642) );
  XNOR U34143 ( .A(n34645), .B(n34646), .Z(n34639) );
  AND U34144 ( .A(n34647), .B(n34648), .Z(n34646) );
  XOR U34145 ( .A(n34645), .B(n34649), .Z(n34647) );
  XNOR U34146 ( .A(n34628), .B(n34625), .Z(n34638) );
  AND U34147 ( .A(n34650), .B(n34651), .Z(n34625) );
  XOR U34148 ( .A(n34652), .B(n34653), .Z(n34628) );
  AND U34149 ( .A(n34654), .B(n34655), .Z(n34653) );
  XOR U34150 ( .A(n34652), .B(n34656), .Z(n34654) );
  XNOR U34151 ( .A(n34589), .B(n34634), .Z(n34636) );
  XNOR U34152 ( .A(n34657), .B(n34658), .Z(n34589) );
  AND U34153 ( .A(n550), .B(n34659), .Z(n34658) );
  XNOR U34154 ( .A(n34660), .B(n34661), .Z(n34659) );
  XOR U34155 ( .A(n34662), .B(n34663), .Z(n34634) );
  AND U34156 ( .A(n34664), .B(n34665), .Z(n34663) );
  XNOR U34157 ( .A(n34662), .B(n34650), .Z(n34665) );
  IV U34158 ( .A(n34600), .Z(n34650) );
  XNOR U34159 ( .A(n34666), .B(n34643), .Z(n34600) );
  XNOR U34160 ( .A(n34667), .B(n34649), .Z(n34643) );
  XOR U34161 ( .A(n34668), .B(n34669), .Z(n34649) );
  NOR U34162 ( .A(n34670), .B(n34671), .Z(n34669) );
  XNOR U34163 ( .A(n34668), .B(n34672), .Z(n34670) );
  XNOR U34164 ( .A(n34648), .B(n34640), .Z(n34667) );
  XOR U34165 ( .A(n34673), .B(n34674), .Z(n34640) );
  AND U34166 ( .A(n34675), .B(n34676), .Z(n34674) );
  XNOR U34167 ( .A(n34673), .B(n34677), .Z(n34675) );
  XNOR U34168 ( .A(n34678), .B(n34645), .Z(n34648) );
  XOR U34169 ( .A(n34679), .B(n34680), .Z(n34645) );
  AND U34170 ( .A(n34681), .B(n34682), .Z(n34680) );
  XOR U34171 ( .A(n34679), .B(n34683), .Z(n34681) );
  XNOR U34172 ( .A(n34684), .B(n34685), .Z(n34678) );
  NOR U34173 ( .A(n34686), .B(n34687), .Z(n34685) );
  XOR U34174 ( .A(n34684), .B(n34688), .Z(n34686) );
  XNOR U34175 ( .A(n34644), .B(n34651), .Z(n34666) );
  NOR U34176 ( .A(n34606), .B(n34689), .Z(n34651) );
  XOR U34177 ( .A(n34656), .B(n34655), .Z(n34644) );
  XNOR U34178 ( .A(n34690), .B(n34652), .Z(n34655) );
  XOR U34179 ( .A(n34691), .B(n34692), .Z(n34652) );
  AND U34180 ( .A(n34693), .B(n34694), .Z(n34692) );
  XOR U34181 ( .A(n34691), .B(n34695), .Z(n34693) );
  XNOR U34182 ( .A(n34696), .B(n34697), .Z(n34690) );
  NOR U34183 ( .A(n34698), .B(n34699), .Z(n34697) );
  XNOR U34184 ( .A(n34696), .B(n34700), .Z(n34698) );
  XOR U34185 ( .A(n34701), .B(n34702), .Z(n34656) );
  NOR U34186 ( .A(n34703), .B(n34704), .Z(n34702) );
  XNOR U34187 ( .A(n34701), .B(n34705), .Z(n34703) );
  XNOR U34188 ( .A(n34597), .B(n34662), .Z(n34664) );
  XNOR U34189 ( .A(n34706), .B(n34707), .Z(n34597) );
  AND U34190 ( .A(n550), .B(n34708), .Z(n34707) );
  XNOR U34191 ( .A(n34709), .B(n34710), .Z(n34708) );
  AND U34192 ( .A(n34603), .B(n34606), .Z(n34662) );
  XOR U34193 ( .A(n34711), .B(n34689), .Z(n34606) );
  XNOR U34194 ( .A(p_input[2048]), .B(p_input[400]), .Z(n34689) );
  XOR U34195 ( .A(n34677), .B(n34676), .Z(n34711) );
  XNOR U34196 ( .A(n34712), .B(n34683), .Z(n34676) );
  XNOR U34197 ( .A(n34672), .B(n34671), .Z(n34683) );
  XOR U34198 ( .A(n34713), .B(n34668), .Z(n34671) );
  XNOR U34199 ( .A(n29266), .B(p_input[410]), .Z(n34668) );
  XNOR U34200 ( .A(p_input[2059]), .B(p_input[411]), .Z(n34713) );
  XOR U34201 ( .A(p_input[2060]), .B(p_input[412]), .Z(n34672) );
  XNOR U34202 ( .A(n34682), .B(n34673), .Z(n34712) );
  XNOR U34203 ( .A(n29494), .B(p_input[401]), .Z(n34673) );
  XOR U34204 ( .A(n34714), .B(n34688), .Z(n34682) );
  XNOR U34205 ( .A(p_input[2063]), .B(p_input[415]), .Z(n34688) );
  XOR U34206 ( .A(n34679), .B(n34687), .Z(n34714) );
  XOR U34207 ( .A(n34715), .B(n34684), .Z(n34687) );
  XOR U34208 ( .A(p_input[2061]), .B(p_input[413]), .Z(n34684) );
  XNOR U34209 ( .A(p_input[2062]), .B(p_input[414]), .Z(n34715) );
  XNOR U34210 ( .A(n29036), .B(p_input[409]), .Z(n34679) );
  XNOR U34211 ( .A(n34695), .B(n34694), .Z(n34677) );
  XNOR U34212 ( .A(n34716), .B(n34700), .Z(n34694) );
  XOR U34213 ( .A(p_input[2056]), .B(p_input[408]), .Z(n34700) );
  XOR U34214 ( .A(n34691), .B(n34699), .Z(n34716) );
  XOR U34215 ( .A(n34717), .B(n34696), .Z(n34699) );
  XOR U34216 ( .A(p_input[2054]), .B(p_input[406]), .Z(n34696) );
  XNOR U34217 ( .A(p_input[2055]), .B(p_input[407]), .Z(n34717) );
  XNOR U34218 ( .A(n29039), .B(p_input[402]), .Z(n34691) );
  XNOR U34219 ( .A(n34705), .B(n34704), .Z(n34695) );
  XOR U34220 ( .A(n34718), .B(n34701), .Z(n34704) );
  XOR U34221 ( .A(p_input[2051]), .B(p_input[403]), .Z(n34701) );
  XNOR U34222 ( .A(p_input[2052]), .B(p_input[404]), .Z(n34718) );
  XOR U34223 ( .A(p_input[2053]), .B(p_input[405]), .Z(n34705) );
  XNOR U34224 ( .A(n34719), .B(n34720), .Z(n34603) );
  AND U34225 ( .A(n550), .B(n34721), .Z(n34720) );
  XNOR U34226 ( .A(n34722), .B(n34723), .Z(n550) );
  AND U34227 ( .A(n34724), .B(n34725), .Z(n34723) );
  XOR U34228 ( .A(n34617), .B(n34722), .Z(n34725) );
  XNOR U34229 ( .A(n34726), .B(n34722), .Z(n34724) );
  XOR U34230 ( .A(n34727), .B(n34728), .Z(n34722) );
  AND U34231 ( .A(n34729), .B(n34730), .Z(n34728) );
  XOR U34232 ( .A(n34632), .B(n34727), .Z(n34730) );
  XOR U34233 ( .A(n34727), .B(n34633), .Z(n34729) );
  XOR U34234 ( .A(n34731), .B(n34732), .Z(n34727) );
  AND U34235 ( .A(n34733), .B(n34734), .Z(n34732) );
  XOR U34236 ( .A(n34660), .B(n34731), .Z(n34734) );
  XOR U34237 ( .A(n34731), .B(n34661), .Z(n34733) );
  XOR U34238 ( .A(n34735), .B(n34736), .Z(n34731) );
  AND U34239 ( .A(n34737), .B(n34738), .Z(n34736) );
  XOR U34240 ( .A(n34735), .B(n34709), .Z(n34738) );
  XNOR U34241 ( .A(n34739), .B(n34740), .Z(n34563) );
  AND U34242 ( .A(n554), .B(n34741), .Z(n34740) );
  XNOR U34243 ( .A(n34742), .B(n34743), .Z(n554) );
  AND U34244 ( .A(n34744), .B(n34745), .Z(n34743) );
  XOR U34245 ( .A(n34742), .B(n34573), .Z(n34745) );
  XNOR U34246 ( .A(n34742), .B(n34533), .Z(n34744) );
  XOR U34247 ( .A(n34746), .B(n34747), .Z(n34742) );
  AND U34248 ( .A(n34748), .B(n34749), .Z(n34747) );
  XOR U34249 ( .A(n34746), .B(n34541), .Z(n34748) );
  XOR U34250 ( .A(n34750), .B(n34751), .Z(n34524) );
  AND U34251 ( .A(n558), .B(n34741), .Z(n34751) );
  XNOR U34252 ( .A(n34739), .B(n34750), .Z(n34741) );
  XNOR U34253 ( .A(n34752), .B(n34753), .Z(n558) );
  AND U34254 ( .A(n34754), .B(n34755), .Z(n34753) );
  XNOR U34255 ( .A(n34756), .B(n34752), .Z(n34755) );
  IV U34256 ( .A(n34573), .Z(n34756) );
  XOR U34257 ( .A(n34726), .B(n34757), .Z(n34573) );
  AND U34258 ( .A(n561), .B(n34758), .Z(n34757) );
  XOR U34259 ( .A(n34616), .B(n34613), .Z(n34758) );
  IV U34260 ( .A(n34726), .Z(n34616) );
  XNOR U34261 ( .A(n34533), .B(n34752), .Z(n34754) );
  XOR U34262 ( .A(n34759), .B(n34760), .Z(n34533) );
  AND U34263 ( .A(n577), .B(n34761), .Z(n34760) );
  XOR U34264 ( .A(n34746), .B(n34762), .Z(n34752) );
  AND U34265 ( .A(n34763), .B(n34749), .Z(n34762) );
  XNOR U34266 ( .A(n34583), .B(n34746), .Z(n34749) );
  XOR U34267 ( .A(n34633), .B(n34764), .Z(n34583) );
  AND U34268 ( .A(n561), .B(n34765), .Z(n34764) );
  XOR U34269 ( .A(n34629), .B(n34633), .Z(n34765) );
  XNOR U34270 ( .A(n34766), .B(n34746), .Z(n34763) );
  IV U34271 ( .A(n34541), .Z(n34766) );
  XOR U34272 ( .A(n34767), .B(n34768), .Z(n34541) );
  AND U34273 ( .A(n577), .B(n34769), .Z(n34768) );
  XOR U34274 ( .A(n34770), .B(n34771), .Z(n34746) );
  AND U34275 ( .A(n34772), .B(n34773), .Z(n34771) );
  XNOR U34276 ( .A(n34593), .B(n34770), .Z(n34773) );
  XOR U34277 ( .A(n34661), .B(n34774), .Z(n34593) );
  AND U34278 ( .A(n561), .B(n34775), .Z(n34774) );
  XOR U34279 ( .A(n34657), .B(n34661), .Z(n34775) );
  XOR U34280 ( .A(n34770), .B(n34550), .Z(n34772) );
  XOR U34281 ( .A(n34776), .B(n34777), .Z(n34550) );
  AND U34282 ( .A(n577), .B(n34778), .Z(n34777) );
  XOR U34283 ( .A(n34779), .B(n34780), .Z(n34770) );
  AND U34284 ( .A(n34781), .B(n34782), .Z(n34780) );
  XNOR U34285 ( .A(n34779), .B(n34601), .Z(n34782) );
  XOR U34286 ( .A(n34710), .B(n34783), .Z(n34601) );
  AND U34287 ( .A(n561), .B(n34784), .Z(n34783) );
  XOR U34288 ( .A(n34706), .B(n34710), .Z(n34784) );
  XNOR U34289 ( .A(n34785), .B(n34779), .Z(n34781) );
  IV U34290 ( .A(n34560), .Z(n34785) );
  XOR U34291 ( .A(n34786), .B(n34787), .Z(n34560) );
  AND U34292 ( .A(n577), .B(n34788), .Z(n34787) );
  AND U34293 ( .A(n34750), .B(n34739), .Z(n34779) );
  XNOR U34294 ( .A(n34789), .B(n34790), .Z(n34739) );
  AND U34295 ( .A(n561), .B(n34721), .Z(n34790) );
  XNOR U34296 ( .A(n34719), .B(n34789), .Z(n34721) );
  XNOR U34297 ( .A(n34791), .B(n34792), .Z(n561) );
  AND U34298 ( .A(n34793), .B(n34794), .Z(n34792) );
  XNOR U34299 ( .A(n34791), .B(n34613), .Z(n34794) );
  IV U34300 ( .A(n34617), .Z(n34613) );
  XOR U34301 ( .A(n34795), .B(n34796), .Z(n34617) );
  AND U34302 ( .A(n565), .B(n34797), .Z(n34796) );
  XOR U34303 ( .A(n34798), .B(n34795), .Z(n34797) );
  XNOR U34304 ( .A(n34791), .B(n34726), .Z(n34793) );
  XOR U34305 ( .A(n34799), .B(n34800), .Z(n34726) );
  AND U34306 ( .A(n573), .B(n34761), .Z(n34800) );
  XOR U34307 ( .A(n34759), .B(n34799), .Z(n34761) );
  XOR U34308 ( .A(n34801), .B(n34802), .Z(n34791) );
  AND U34309 ( .A(n34803), .B(n34804), .Z(n34802) );
  XNOR U34310 ( .A(n34801), .B(n34629), .Z(n34804) );
  IV U34311 ( .A(n34632), .Z(n34629) );
  XOR U34312 ( .A(n34805), .B(n34806), .Z(n34632) );
  AND U34313 ( .A(n565), .B(n34807), .Z(n34806) );
  XOR U34314 ( .A(n34808), .B(n34805), .Z(n34807) );
  XOR U34315 ( .A(n34633), .B(n34801), .Z(n34803) );
  XOR U34316 ( .A(n34809), .B(n34810), .Z(n34633) );
  AND U34317 ( .A(n573), .B(n34769), .Z(n34810) );
  XOR U34318 ( .A(n34809), .B(n34767), .Z(n34769) );
  XOR U34319 ( .A(n34811), .B(n34812), .Z(n34801) );
  AND U34320 ( .A(n34813), .B(n34814), .Z(n34812) );
  XNOR U34321 ( .A(n34811), .B(n34657), .Z(n34814) );
  IV U34322 ( .A(n34660), .Z(n34657) );
  XOR U34323 ( .A(n34815), .B(n34816), .Z(n34660) );
  AND U34324 ( .A(n565), .B(n34817), .Z(n34816) );
  XNOR U34325 ( .A(n34818), .B(n34815), .Z(n34817) );
  XOR U34326 ( .A(n34661), .B(n34811), .Z(n34813) );
  XOR U34327 ( .A(n34819), .B(n34820), .Z(n34661) );
  AND U34328 ( .A(n573), .B(n34778), .Z(n34820) );
  XOR U34329 ( .A(n34819), .B(n34776), .Z(n34778) );
  XOR U34330 ( .A(n34735), .B(n34821), .Z(n34811) );
  AND U34331 ( .A(n34737), .B(n34822), .Z(n34821) );
  XNOR U34332 ( .A(n34735), .B(n34706), .Z(n34822) );
  IV U34333 ( .A(n34709), .Z(n34706) );
  XOR U34334 ( .A(n34823), .B(n34824), .Z(n34709) );
  AND U34335 ( .A(n565), .B(n34825), .Z(n34824) );
  XOR U34336 ( .A(n34826), .B(n34823), .Z(n34825) );
  XOR U34337 ( .A(n34710), .B(n34735), .Z(n34737) );
  XOR U34338 ( .A(n34827), .B(n34828), .Z(n34710) );
  AND U34339 ( .A(n573), .B(n34788), .Z(n34828) );
  XOR U34340 ( .A(n34827), .B(n34786), .Z(n34788) );
  AND U34341 ( .A(n34789), .B(n34719), .Z(n34735) );
  XNOR U34342 ( .A(n34829), .B(n34830), .Z(n34719) );
  AND U34343 ( .A(n565), .B(n34831), .Z(n34830) );
  XNOR U34344 ( .A(n34832), .B(n34829), .Z(n34831) );
  XNOR U34345 ( .A(n34833), .B(n34834), .Z(n565) );
  AND U34346 ( .A(n34835), .B(n34836), .Z(n34834) );
  XOR U34347 ( .A(n34798), .B(n34833), .Z(n34836) );
  AND U34348 ( .A(n34837), .B(n34838), .Z(n34798) );
  XNOR U34349 ( .A(n34795), .B(n34833), .Z(n34835) );
  XNOR U34350 ( .A(n34839), .B(n34840), .Z(n34795) );
  AND U34351 ( .A(n569), .B(n34841), .Z(n34840) );
  XNOR U34352 ( .A(n34842), .B(n34843), .Z(n34841) );
  XOR U34353 ( .A(n34844), .B(n34845), .Z(n34833) );
  AND U34354 ( .A(n34846), .B(n34847), .Z(n34845) );
  XNOR U34355 ( .A(n34844), .B(n34837), .Z(n34847) );
  IV U34356 ( .A(n34808), .Z(n34837) );
  XOR U34357 ( .A(n34848), .B(n34849), .Z(n34808) );
  XOR U34358 ( .A(n34850), .B(n34838), .Z(n34849) );
  AND U34359 ( .A(n34818), .B(n34851), .Z(n34838) );
  AND U34360 ( .A(n34852), .B(n34853), .Z(n34850) );
  XOR U34361 ( .A(n34854), .B(n34848), .Z(n34852) );
  XNOR U34362 ( .A(n34805), .B(n34844), .Z(n34846) );
  XNOR U34363 ( .A(n34855), .B(n34856), .Z(n34805) );
  AND U34364 ( .A(n569), .B(n34857), .Z(n34856) );
  XNOR U34365 ( .A(n34858), .B(n34859), .Z(n34857) );
  XOR U34366 ( .A(n34860), .B(n34861), .Z(n34844) );
  AND U34367 ( .A(n34862), .B(n34863), .Z(n34861) );
  XNOR U34368 ( .A(n34860), .B(n34818), .Z(n34863) );
  XOR U34369 ( .A(n34864), .B(n34853), .Z(n34818) );
  XNOR U34370 ( .A(n34865), .B(n34848), .Z(n34853) );
  XOR U34371 ( .A(n34866), .B(n34867), .Z(n34848) );
  AND U34372 ( .A(n34868), .B(n34869), .Z(n34867) );
  XOR U34373 ( .A(n34870), .B(n34866), .Z(n34868) );
  XNOR U34374 ( .A(n34871), .B(n34872), .Z(n34865) );
  AND U34375 ( .A(n34873), .B(n34874), .Z(n34872) );
  XOR U34376 ( .A(n34871), .B(n34875), .Z(n34873) );
  XNOR U34377 ( .A(n34854), .B(n34851), .Z(n34864) );
  AND U34378 ( .A(n34876), .B(n34877), .Z(n34851) );
  XOR U34379 ( .A(n34878), .B(n34879), .Z(n34854) );
  AND U34380 ( .A(n34880), .B(n34881), .Z(n34879) );
  XOR U34381 ( .A(n34878), .B(n34882), .Z(n34880) );
  XNOR U34382 ( .A(n34815), .B(n34860), .Z(n34862) );
  XNOR U34383 ( .A(n34883), .B(n34884), .Z(n34815) );
  AND U34384 ( .A(n569), .B(n34885), .Z(n34884) );
  XNOR U34385 ( .A(n34886), .B(n34887), .Z(n34885) );
  XOR U34386 ( .A(n34888), .B(n34889), .Z(n34860) );
  AND U34387 ( .A(n34890), .B(n34891), .Z(n34889) );
  XNOR U34388 ( .A(n34888), .B(n34876), .Z(n34891) );
  IV U34389 ( .A(n34826), .Z(n34876) );
  XNOR U34390 ( .A(n34892), .B(n34869), .Z(n34826) );
  XNOR U34391 ( .A(n34893), .B(n34875), .Z(n34869) );
  XOR U34392 ( .A(n34894), .B(n34895), .Z(n34875) );
  NOR U34393 ( .A(n34896), .B(n34897), .Z(n34895) );
  XNOR U34394 ( .A(n34894), .B(n34898), .Z(n34896) );
  XNOR U34395 ( .A(n34874), .B(n34866), .Z(n34893) );
  XOR U34396 ( .A(n34899), .B(n34900), .Z(n34866) );
  AND U34397 ( .A(n34901), .B(n34902), .Z(n34900) );
  XNOR U34398 ( .A(n34899), .B(n34903), .Z(n34901) );
  XNOR U34399 ( .A(n34904), .B(n34871), .Z(n34874) );
  XOR U34400 ( .A(n34905), .B(n34906), .Z(n34871) );
  AND U34401 ( .A(n34907), .B(n34908), .Z(n34906) );
  XOR U34402 ( .A(n34905), .B(n34909), .Z(n34907) );
  XNOR U34403 ( .A(n34910), .B(n34911), .Z(n34904) );
  NOR U34404 ( .A(n34912), .B(n34913), .Z(n34911) );
  XOR U34405 ( .A(n34910), .B(n34914), .Z(n34912) );
  XNOR U34406 ( .A(n34870), .B(n34877), .Z(n34892) );
  NOR U34407 ( .A(n34832), .B(n34915), .Z(n34877) );
  XOR U34408 ( .A(n34882), .B(n34881), .Z(n34870) );
  XNOR U34409 ( .A(n34916), .B(n34878), .Z(n34881) );
  XOR U34410 ( .A(n34917), .B(n34918), .Z(n34878) );
  AND U34411 ( .A(n34919), .B(n34920), .Z(n34918) );
  XOR U34412 ( .A(n34917), .B(n34921), .Z(n34919) );
  XNOR U34413 ( .A(n34922), .B(n34923), .Z(n34916) );
  NOR U34414 ( .A(n34924), .B(n34925), .Z(n34923) );
  XNOR U34415 ( .A(n34922), .B(n34926), .Z(n34924) );
  XOR U34416 ( .A(n34927), .B(n34928), .Z(n34882) );
  NOR U34417 ( .A(n34929), .B(n34930), .Z(n34928) );
  XNOR U34418 ( .A(n34927), .B(n34931), .Z(n34929) );
  XNOR U34419 ( .A(n34823), .B(n34888), .Z(n34890) );
  XNOR U34420 ( .A(n34932), .B(n34933), .Z(n34823) );
  AND U34421 ( .A(n569), .B(n34934), .Z(n34933) );
  XNOR U34422 ( .A(n34935), .B(n34936), .Z(n34934) );
  AND U34423 ( .A(n34829), .B(n34832), .Z(n34888) );
  XOR U34424 ( .A(n34937), .B(n34915), .Z(n34832) );
  XNOR U34425 ( .A(p_input[2048]), .B(p_input[416]), .Z(n34915) );
  XOR U34426 ( .A(n34903), .B(n34902), .Z(n34937) );
  XNOR U34427 ( .A(n34938), .B(n34909), .Z(n34902) );
  XNOR U34428 ( .A(n34898), .B(n34897), .Z(n34909) );
  XOR U34429 ( .A(n34939), .B(n34894), .Z(n34897) );
  XNOR U34430 ( .A(n29266), .B(p_input[426]), .Z(n34894) );
  XNOR U34431 ( .A(p_input[2059]), .B(p_input[427]), .Z(n34939) );
  XOR U34432 ( .A(p_input[2060]), .B(p_input[428]), .Z(n34898) );
  XNOR U34433 ( .A(n34908), .B(n34899), .Z(n34938) );
  XNOR U34434 ( .A(n29494), .B(p_input[417]), .Z(n34899) );
  XOR U34435 ( .A(n34940), .B(n34914), .Z(n34908) );
  XNOR U34436 ( .A(p_input[2063]), .B(p_input[431]), .Z(n34914) );
  XOR U34437 ( .A(n34905), .B(n34913), .Z(n34940) );
  XOR U34438 ( .A(n34941), .B(n34910), .Z(n34913) );
  XOR U34439 ( .A(p_input[2061]), .B(p_input[429]), .Z(n34910) );
  XNOR U34440 ( .A(p_input[2062]), .B(p_input[430]), .Z(n34941) );
  XNOR U34441 ( .A(n29036), .B(p_input[425]), .Z(n34905) );
  XNOR U34442 ( .A(n34921), .B(n34920), .Z(n34903) );
  XNOR U34443 ( .A(n34942), .B(n34926), .Z(n34920) );
  XOR U34444 ( .A(p_input[2056]), .B(p_input[424]), .Z(n34926) );
  XOR U34445 ( .A(n34917), .B(n34925), .Z(n34942) );
  XOR U34446 ( .A(n34943), .B(n34922), .Z(n34925) );
  XOR U34447 ( .A(p_input[2054]), .B(p_input[422]), .Z(n34922) );
  XNOR U34448 ( .A(p_input[2055]), .B(p_input[423]), .Z(n34943) );
  XNOR U34449 ( .A(n29039), .B(p_input[418]), .Z(n34917) );
  XNOR U34450 ( .A(n34931), .B(n34930), .Z(n34921) );
  XOR U34451 ( .A(n34944), .B(n34927), .Z(n34930) );
  XOR U34452 ( .A(p_input[2051]), .B(p_input[419]), .Z(n34927) );
  XNOR U34453 ( .A(p_input[2052]), .B(p_input[420]), .Z(n34944) );
  XOR U34454 ( .A(p_input[2053]), .B(p_input[421]), .Z(n34931) );
  XNOR U34455 ( .A(n34945), .B(n34946), .Z(n34829) );
  AND U34456 ( .A(n569), .B(n34947), .Z(n34946) );
  XNOR U34457 ( .A(n34948), .B(n34949), .Z(n569) );
  AND U34458 ( .A(n34950), .B(n34951), .Z(n34949) );
  XOR U34459 ( .A(n34843), .B(n34948), .Z(n34951) );
  XNOR U34460 ( .A(n34952), .B(n34948), .Z(n34950) );
  XOR U34461 ( .A(n34953), .B(n34954), .Z(n34948) );
  AND U34462 ( .A(n34955), .B(n34956), .Z(n34954) );
  XOR U34463 ( .A(n34858), .B(n34953), .Z(n34956) );
  XOR U34464 ( .A(n34953), .B(n34859), .Z(n34955) );
  XOR U34465 ( .A(n34957), .B(n34958), .Z(n34953) );
  AND U34466 ( .A(n34959), .B(n34960), .Z(n34958) );
  XOR U34467 ( .A(n34886), .B(n34957), .Z(n34960) );
  XOR U34468 ( .A(n34957), .B(n34887), .Z(n34959) );
  XOR U34469 ( .A(n34961), .B(n34962), .Z(n34957) );
  AND U34470 ( .A(n34963), .B(n34964), .Z(n34962) );
  XOR U34471 ( .A(n34961), .B(n34935), .Z(n34964) );
  XNOR U34472 ( .A(n34965), .B(n34966), .Z(n34789) );
  AND U34473 ( .A(n573), .B(n34967), .Z(n34966) );
  XNOR U34474 ( .A(n34968), .B(n34969), .Z(n573) );
  AND U34475 ( .A(n34970), .B(n34971), .Z(n34969) );
  XOR U34476 ( .A(n34968), .B(n34799), .Z(n34971) );
  XNOR U34477 ( .A(n34968), .B(n34759), .Z(n34970) );
  XOR U34478 ( .A(n34972), .B(n34973), .Z(n34968) );
  AND U34479 ( .A(n34974), .B(n34975), .Z(n34973) );
  XOR U34480 ( .A(n34972), .B(n34767), .Z(n34974) );
  XOR U34481 ( .A(n34976), .B(n34977), .Z(n34750) );
  AND U34482 ( .A(n577), .B(n34967), .Z(n34977) );
  XNOR U34483 ( .A(n34965), .B(n34976), .Z(n34967) );
  XNOR U34484 ( .A(n34978), .B(n34979), .Z(n577) );
  AND U34485 ( .A(n34980), .B(n34981), .Z(n34979) );
  XNOR U34486 ( .A(n34982), .B(n34978), .Z(n34981) );
  IV U34487 ( .A(n34799), .Z(n34982) );
  XOR U34488 ( .A(n34952), .B(n34983), .Z(n34799) );
  AND U34489 ( .A(n580), .B(n34984), .Z(n34983) );
  XOR U34490 ( .A(n34842), .B(n34839), .Z(n34984) );
  IV U34491 ( .A(n34952), .Z(n34842) );
  XNOR U34492 ( .A(n34759), .B(n34978), .Z(n34980) );
  XOR U34493 ( .A(n34985), .B(n34986), .Z(n34759) );
  AND U34494 ( .A(n596), .B(n34987), .Z(n34986) );
  XOR U34495 ( .A(n34972), .B(n34988), .Z(n34978) );
  AND U34496 ( .A(n34989), .B(n34975), .Z(n34988) );
  XNOR U34497 ( .A(n34809), .B(n34972), .Z(n34975) );
  XOR U34498 ( .A(n34859), .B(n34990), .Z(n34809) );
  AND U34499 ( .A(n580), .B(n34991), .Z(n34990) );
  XOR U34500 ( .A(n34855), .B(n34859), .Z(n34991) );
  XNOR U34501 ( .A(n34992), .B(n34972), .Z(n34989) );
  IV U34502 ( .A(n34767), .Z(n34992) );
  XOR U34503 ( .A(n34993), .B(n34994), .Z(n34767) );
  AND U34504 ( .A(n596), .B(n34995), .Z(n34994) );
  XOR U34505 ( .A(n34996), .B(n34997), .Z(n34972) );
  AND U34506 ( .A(n34998), .B(n34999), .Z(n34997) );
  XNOR U34507 ( .A(n34819), .B(n34996), .Z(n34999) );
  XOR U34508 ( .A(n34887), .B(n35000), .Z(n34819) );
  AND U34509 ( .A(n580), .B(n35001), .Z(n35000) );
  XOR U34510 ( .A(n34883), .B(n34887), .Z(n35001) );
  XOR U34511 ( .A(n34996), .B(n34776), .Z(n34998) );
  XOR U34512 ( .A(n35002), .B(n35003), .Z(n34776) );
  AND U34513 ( .A(n596), .B(n35004), .Z(n35003) );
  XOR U34514 ( .A(n35005), .B(n35006), .Z(n34996) );
  AND U34515 ( .A(n35007), .B(n35008), .Z(n35006) );
  XNOR U34516 ( .A(n35005), .B(n34827), .Z(n35008) );
  XOR U34517 ( .A(n34936), .B(n35009), .Z(n34827) );
  AND U34518 ( .A(n580), .B(n35010), .Z(n35009) );
  XOR U34519 ( .A(n34932), .B(n34936), .Z(n35010) );
  XNOR U34520 ( .A(n35011), .B(n35005), .Z(n35007) );
  IV U34521 ( .A(n34786), .Z(n35011) );
  XOR U34522 ( .A(n35012), .B(n35013), .Z(n34786) );
  AND U34523 ( .A(n596), .B(n35014), .Z(n35013) );
  AND U34524 ( .A(n34976), .B(n34965), .Z(n35005) );
  XNOR U34525 ( .A(n35015), .B(n35016), .Z(n34965) );
  AND U34526 ( .A(n580), .B(n34947), .Z(n35016) );
  XNOR U34527 ( .A(n34945), .B(n35015), .Z(n34947) );
  XNOR U34528 ( .A(n35017), .B(n35018), .Z(n580) );
  AND U34529 ( .A(n35019), .B(n35020), .Z(n35018) );
  XNOR U34530 ( .A(n35017), .B(n34839), .Z(n35020) );
  IV U34531 ( .A(n34843), .Z(n34839) );
  XOR U34532 ( .A(n35021), .B(n35022), .Z(n34843) );
  AND U34533 ( .A(n584), .B(n35023), .Z(n35022) );
  XOR U34534 ( .A(n35024), .B(n35021), .Z(n35023) );
  XNOR U34535 ( .A(n35017), .B(n34952), .Z(n35019) );
  XOR U34536 ( .A(n35025), .B(n35026), .Z(n34952) );
  AND U34537 ( .A(n592), .B(n34987), .Z(n35026) );
  XOR U34538 ( .A(n34985), .B(n35025), .Z(n34987) );
  XOR U34539 ( .A(n35027), .B(n35028), .Z(n35017) );
  AND U34540 ( .A(n35029), .B(n35030), .Z(n35028) );
  XNOR U34541 ( .A(n35027), .B(n34855), .Z(n35030) );
  IV U34542 ( .A(n34858), .Z(n34855) );
  XOR U34543 ( .A(n35031), .B(n35032), .Z(n34858) );
  AND U34544 ( .A(n584), .B(n35033), .Z(n35032) );
  XOR U34545 ( .A(n35034), .B(n35031), .Z(n35033) );
  XOR U34546 ( .A(n34859), .B(n35027), .Z(n35029) );
  XOR U34547 ( .A(n35035), .B(n35036), .Z(n34859) );
  AND U34548 ( .A(n592), .B(n34995), .Z(n35036) );
  XOR U34549 ( .A(n35035), .B(n34993), .Z(n34995) );
  XOR U34550 ( .A(n35037), .B(n35038), .Z(n35027) );
  AND U34551 ( .A(n35039), .B(n35040), .Z(n35038) );
  XNOR U34552 ( .A(n35037), .B(n34883), .Z(n35040) );
  IV U34553 ( .A(n34886), .Z(n34883) );
  XOR U34554 ( .A(n35041), .B(n35042), .Z(n34886) );
  AND U34555 ( .A(n584), .B(n35043), .Z(n35042) );
  XNOR U34556 ( .A(n35044), .B(n35041), .Z(n35043) );
  XOR U34557 ( .A(n34887), .B(n35037), .Z(n35039) );
  XOR U34558 ( .A(n35045), .B(n35046), .Z(n34887) );
  AND U34559 ( .A(n592), .B(n35004), .Z(n35046) );
  XOR U34560 ( .A(n35045), .B(n35002), .Z(n35004) );
  XOR U34561 ( .A(n34961), .B(n35047), .Z(n35037) );
  AND U34562 ( .A(n34963), .B(n35048), .Z(n35047) );
  XNOR U34563 ( .A(n34961), .B(n34932), .Z(n35048) );
  IV U34564 ( .A(n34935), .Z(n34932) );
  XOR U34565 ( .A(n35049), .B(n35050), .Z(n34935) );
  AND U34566 ( .A(n584), .B(n35051), .Z(n35050) );
  XOR U34567 ( .A(n35052), .B(n35049), .Z(n35051) );
  XOR U34568 ( .A(n34936), .B(n34961), .Z(n34963) );
  XOR U34569 ( .A(n35053), .B(n35054), .Z(n34936) );
  AND U34570 ( .A(n592), .B(n35014), .Z(n35054) );
  XOR U34571 ( .A(n35053), .B(n35012), .Z(n35014) );
  AND U34572 ( .A(n35015), .B(n34945), .Z(n34961) );
  XNOR U34573 ( .A(n35055), .B(n35056), .Z(n34945) );
  AND U34574 ( .A(n584), .B(n35057), .Z(n35056) );
  XNOR U34575 ( .A(n35058), .B(n35055), .Z(n35057) );
  XNOR U34576 ( .A(n35059), .B(n35060), .Z(n584) );
  AND U34577 ( .A(n35061), .B(n35062), .Z(n35060) );
  XOR U34578 ( .A(n35024), .B(n35059), .Z(n35062) );
  AND U34579 ( .A(n35063), .B(n35064), .Z(n35024) );
  XNOR U34580 ( .A(n35021), .B(n35059), .Z(n35061) );
  XNOR U34581 ( .A(n35065), .B(n35066), .Z(n35021) );
  AND U34582 ( .A(n588), .B(n35067), .Z(n35066) );
  XNOR U34583 ( .A(n35068), .B(n35069), .Z(n35067) );
  XOR U34584 ( .A(n35070), .B(n35071), .Z(n35059) );
  AND U34585 ( .A(n35072), .B(n35073), .Z(n35071) );
  XNOR U34586 ( .A(n35070), .B(n35063), .Z(n35073) );
  IV U34587 ( .A(n35034), .Z(n35063) );
  XOR U34588 ( .A(n35074), .B(n35075), .Z(n35034) );
  XOR U34589 ( .A(n35076), .B(n35064), .Z(n35075) );
  AND U34590 ( .A(n35044), .B(n35077), .Z(n35064) );
  AND U34591 ( .A(n35078), .B(n35079), .Z(n35076) );
  XOR U34592 ( .A(n35080), .B(n35074), .Z(n35078) );
  XNOR U34593 ( .A(n35031), .B(n35070), .Z(n35072) );
  XNOR U34594 ( .A(n35081), .B(n35082), .Z(n35031) );
  AND U34595 ( .A(n588), .B(n35083), .Z(n35082) );
  XNOR U34596 ( .A(n35084), .B(n35085), .Z(n35083) );
  XOR U34597 ( .A(n35086), .B(n35087), .Z(n35070) );
  AND U34598 ( .A(n35088), .B(n35089), .Z(n35087) );
  XNOR U34599 ( .A(n35086), .B(n35044), .Z(n35089) );
  XOR U34600 ( .A(n35090), .B(n35079), .Z(n35044) );
  XNOR U34601 ( .A(n35091), .B(n35074), .Z(n35079) );
  XOR U34602 ( .A(n35092), .B(n35093), .Z(n35074) );
  AND U34603 ( .A(n35094), .B(n35095), .Z(n35093) );
  XOR U34604 ( .A(n35096), .B(n35092), .Z(n35094) );
  XNOR U34605 ( .A(n35097), .B(n35098), .Z(n35091) );
  AND U34606 ( .A(n35099), .B(n35100), .Z(n35098) );
  XOR U34607 ( .A(n35097), .B(n35101), .Z(n35099) );
  XNOR U34608 ( .A(n35080), .B(n35077), .Z(n35090) );
  AND U34609 ( .A(n35102), .B(n35103), .Z(n35077) );
  XOR U34610 ( .A(n35104), .B(n35105), .Z(n35080) );
  AND U34611 ( .A(n35106), .B(n35107), .Z(n35105) );
  XOR U34612 ( .A(n35104), .B(n35108), .Z(n35106) );
  XNOR U34613 ( .A(n35041), .B(n35086), .Z(n35088) );
  XNOR U34614 ( .A(n35109), .B(n35110), .Z(n35041) );
  AND U34615 ( .A(n588), .B(n35111), .Z(n35110) );
  XNOR U34616 ( .A(n35112), .B(n35113), .Z(n35111) );
  XOR U34617 ( .A(n35114), .B(n35115), .Z(n35086) );
  AND U34618 ( .A(n35116), .B(n35117), .Z(n35115) );
  XNOR U34619 ( .A(n35114), .B(n35102), .Z(n35117) );
  IV U34620 ( .A(n35052), .Z(n35102) );
  XNOR U34621 ( .A(n35118), .B(n35095), .Z(n35052) );
  XNOR U34622 ( .A(n35119), .B(n35101), .Z(n35095) );
  XOR U34623 ( .A(n35120), .B(n35121), .Z(n35101) );
  NOR U34624 ( .A(n35122), .B(n35123), .Z(n35121) );
  XNOR U34625 ( .A(n35120), .B(n35124), .Z(n35122) );
  XNOR U34626 ( .A(n35100), .B(n35092), .Z(n35119) );
  XOR U34627 ( .A(n35125), .B(n35126), .Z(n35092) );
  AND U34628 ( .A(n35127), .B(n35128), .Z(n35126) );
  XNOR U34629 ( .A(n35125), .B(n35129), .Z(n35127) );
  XNOR U34630 ( .A(n35130), .B(n35097), .Z(n35100) );
  XOR U34631 ( .A(n35131), .B(n35132), .Z(n35097) );
  AND U34632 ( .A(n35133), .B(n35134), .Z(n35132) );
  XOR U34633 ( .A(n35131), .B(n35135), .Z(n35133) );
  XNOR U34634 ( .A(n35136), .B(n35137), .Z(n35130) );
  NOR U34635 ( .A(n35138), .B(n35139), .Z(n35137) );
  XOR U34636 ( .A(n35136), .B(n35140), .Z(n35138) );
  XNOR U34637 ( .A(n35096), .B(n35103), .Z(n35118) );
  NOR U34638 ( .A(n35058), .B(n35141), .Z(n35103) );
  XOR U34639 ( .A(n35108), .B(n35107), .Z(n35096) );
  XNOR U34640 ( .A(n35142), .B(n35104), .Z(n35107) );
  XOR U34641 ( .A(n35143), .B(n35144), .Z(n35104) );
  AND U34642 ( .A(n35145), .B(n35146), .Z(n35144) );
  XOR U34643 ( .A(n35143), .B(n35147), .Z(n35145) );
  XNOR U34644 ( .A(n35148), .B(n35149), .Z(n35142) );
  NOR U34645 ( .A(n35150), .B(n35151), .Z(n35149) );
  XNOR U34646 ( .A(n35148), .B(n35152), .Z(n35150) );
  XOR U34647 ( .A(n35153), .B(n35154), .Z(n35108) );
  NOR U34648 ( .A(n35155), .B(n35156), .Z(n35154) );
  XNOR U34649 ( .A(n35153), .B(n35157), .Z(n35155) );
  XNOR U34650 ( .A(n35049), .B(n35114), .Z(n35116) );
  XNOR U34651 ( .A(n35158), .B(n35159), .Z(n35049) );
  AND U34652 ( .A(n588), .B(n35160), .Z(n35159) );
  XNOR U34653 ( .A(n35161), .B(n35162), .Z(n35160) );
  AND U34654 ( .A(n35055), .B(n35058), .Z(n35114) );
  XOR U34655 ( .A(n35163), .B(n35141), .Z(n35058) );
  XNOR U34656 ( .A(p_input[2048]), .B(p_input[432]), .Z(n35141) );
  XOR U34657 ( .A(n35129), .B(n35128), .Z(n35163) );
  XNOR U34658 ( .A(n35164), .B(n35135), .Z(n35128) );
  XNOR U34659 ( .A(n35124), .B(n35123), .Z(n35135) );
  XOR U34660 ( .A(n35165), .B(n35120), .Z(n35123) );
  XNOR U34661 ( .A(n29266), .B(p_input[442]), .Z(n35120) );
  XNOR U34662 ( .A(p_input[2059]), .B(p_input[443]), .Z(n35165) );
  XOR U34663 ( .A(p_input[2060]), .B(p_input[444]), .Z(n35124) );
  XNOR U34664 ( .A(n35134), .B(n35125), .Z(n35164) );
  XNOR U34665 ( .A(n29494), .B(p_input[433]), .Z(n35125) );
  XOR U34666 ( .A(n35166), .B(n35140), .Z(n35134) );
  XNOR U34667 ( .A(p_input[2063]), .B(p_input[447]), .Z(n35140) );
  XOR U34668 ( .A(n35131), .B(n35139), .Z(n35166) );
  XOR U34669 ( .A(n35167), .B(n35136), .Z(n35139) );
  XOR U34670 ( .A(p_input[2061]), .B(p_input[445]), .Z(n35136) );
  XNOR U34671 ( .A(p_input[2062]), .B(p_input[446]), .Z(n35167) );
  XNOR U34672 ( .A(n29036), .B(p_input[441]), .Z(n35131) );
  XNOR U34673 ( .A(n35147), .B(n35146), .Z(n35129) );
  XNOR U34674 ( .A(n35168), .B(n35152), .Z(n35146) );
  XOR U34675 ( .A(p_input[2056]), .B(p_input[440]), .Z(n35152) );
  XOR U34676 ( .A(n35143), .B(n35151), .Z(n35168) );
  XOR U34677 ( .A(n35169), .B(n35148), .Z(n35151) );
  XOR U34678 ( .A(p_input[2054]), .B(p_input[438]), .Z(n35148) );
  XNOR U34679 ( .A(p_input[2055]), .B(p_input[439]), .Z(n35169) );
  XNOR U34680 ( .A(n29039), .B(p_input[434]), .Z(n35143) );
  XNOR U34681 ( .A(n35157), .B(n35156), .Z(n35147) );
  XOR U34682 ( .A(n35170), .B(n35153), .Z(n35156) );
  XOR U34683 ( .A(p_input[2051]), .B(p_input[435]), .Z(n35153) );
  XNOR U34684 ( .A(p_input[2052]), .B(p_input[436]), .Z(n35170) );
  XOR U34685 ( .A(p_input[2053]), .B(p_input[437]), .Z(n35157) );
  XNOR U34686 ( .A(n35171), .B(n35172), .Z(n35055) );
  AND U34687 ( .A(n588), .B(n35173), .Z(n35172) );
  XNOR U34688 ( .A(n35174), .B(n35175), .Z(n588) );
  AND U34689 ( .A(n35176), .B(n35177), .Z(n35175) );
  XOR U34690 ( .A(n35069), .B(n35174), .Z(n35177) );
  XNOR U34691 ( .A(n35178), .B(n35174), .Z(n35176) );
  XOR U34692 ( .A(n35179), .B(n35180), .Z(n35174) );
  AND U34693 ( .A(n35181), .B(n35182), .Z(n35180) );
  XOR U34694 ( .A(n35084), .B(n35179), .Z(n35182) );
  XOR U34695 ( .A(n35179), .B(n35085), .Z(n35181) );
  XOR U34696 ( .A(n35183), .B(n35184), .Z(n35179) );
  AND U34697 ( .A(n35185), .B(n35186), .Z(n35184) );
  XOR U34698 ( .A(n35112), .B(n35183), .Z(n35186) );
  XOR U34699 ( .A(n35183), .B(n35113), .Z(n35185) );
  XOR U34700 ( .A(n35187), .B(n35188), .Z(n35183) );
  AND U34701 ( .A(n35189), .B(n35190), .Z(n35188) );
  XOR U34702 ( .A(n35187), .B(n35161), .Z(n35190) );
  XNOR U34703 ( .A(n35191), .B(n35192), .Z(n35015) );
  AND U34704 ( .A(n592), .B(n35193), .Z(n35192) );
  XNOR U34705 ( .A(n35194), .B(n35195), .Z(n592) );
  AND U34706 ( .A(n35196), .B(n35197), .Z(n35195) );
  XOR U34707 ( .A(n35194), .B(n35025), .Z(n35197) );
  XNOR U34708 ( .A(n35194), .B(n34985), .Z(n35196) );
  XOR U34709 ( .A(n35198), .B(n35199), .Z(n35194) );
  AND U34710 ( .A(n35200), .B(n35201), .Z(n35199) );
  XOR U34711 ( .A(n35198), .B(n34993), .Z(n35200) );
  XOR U34712 ( .A(n35202), .B(n35203), .Z(n34976) );
  AND U34713 ( .A(n596), .B(n35193), .Z(n35203) );
  XNOR U34714 ( .A(n35191), .B(n35202), .Z(n35193) );
  XNOR U34715 ( .A(n35204), .B(n35205), .Z(n596) );
  AND U34716 ( .A(n35206), .B(n35207), .Z(n35205) );
  XNOR U34717 ( .A(n35208), .B(n35204), .Z(n35207) );
  IV U34718 ( .A(n35025), .Z(n35208) );
  XOR U34719 ( .A(n35178), .B(n35209), .Z(n35025) );
  AND U34720 ( .A(n599), .B(n35210), .Z(n35209) );
  XOR U34721 ( .A(n35068), .B(n35065), .Z(n35210) );
  IV U34722 ( .A(n35178), .Z(n35068) );
  XNOR U34723 ( .A(n34985), .B(n35204), .Z(n35206) );
  XOR U34724 ( .A(n35211), .B(n35212), .Z(n34985) );
  AND U34725 ( .A(n615), .B(n35213), .Z(n35212) );
  XOR U34726 ( .A(n35198), .B(n35214), .Z(n35204) );
  AND U34727 ( .A(n35215), .B(n35201), .Z(n35214) );
  XNOR U34728 ( .A(n35035), .B(n35198), .Z(n35201) );
  XOR U34729 ( .A(n35085), .B(n35216), .Z(n35035) );
  AND U34730 ( .A(n599), .B(n35217), .Z(n35216) );
  XOR U34731 ( .A(n35081), .B(n35085), .Z(n35217) );
  XNOR U34732 ( .A(n35218), .B(n35198), .Z(n35215) );
  IV U34733 ( .A(n34993), .Z(n35218) );
  XOR U34734 ( .A(n35219), .B(n35220), .Z(n34993) );
  AND U34735 ( .A(n615), .B(n35221), .Z(n35220) );
  XOR U34736 ( .A(n35222), .B(n35223), .Z(n35198) );
  AND U34737 ( .A(n35224), .B(n35225), .Z(n35223) );
  XNOR U34738 ( .A(n35045), .B(n35222), .Z(n35225) );
  XOR U34739 ( .A(n35113), .B(n35226), .Z(n35045) );
  AND U34740 ( .A(n599), .B(n35227), .Z(n35226) );
  XOR U34741 ( .A(n35109), .B(n35113), .Z(n35227) );
  XOR U34742 ( .A(n35222), .B(n35002), .Z(n35224) );
  XOR U34743 ( .A(n35228), .B(n35229), .Z(n35002) );
  AND U34744 ( .A(n615), .B(n35230), .Z(n35229) );
  XOR U34745 ( .A(n35231), .B(n35232), .Z(n35222) );
  AND U34746 ( .A(n35233), .B(n35234), .Z(n35232) );
  XNOR U34747 ( .A(n35231), .B(n35053), .Z(n35234) );
  XOR U34748 ( .A(n35162), .B(n35235), .Z(n35053) );
  AND U34749 ( .A(n599), .B(n35236), .Z(n35235) );
  XOR U34750 ( .A(n35158), .B(n35162), .Z(n35236) );
  XNOR U34751 ( .A(n35237), .B(n35231), .Z(n35233) );
  IV U34752 ( .A(n35012), .Z(n35237) );
  XOR U34753 ( .A(n35238), .B(n35239), .Z(n35012) );
  AND U34754 ( .A(n615), .B(n35240), .Z(n35239) );
  AND U34755 ( .A(n35202), .B(n35191), .Z(n35231) );
  XNOR U34756 ( .A(n35241), .B(n35242), .Z(n35191) );
  AND U34757 ( .A(n599), .B(n35173), .Z(n35242) );
  XNOR U34758 ( .A(n35171), .B(n35241), .Z(n35173) );
  XNOR U34759 ( .A(n35243), .B(n35244), .Z(n599) );
  AND U34760 ( .A(n35245), .B(n35246), .Z(n35244) );
  XNOR U34761 ( .A(n35243), .B(n35065), .Z(n35246) );
  IV U34762 ( .A(n35069), .Z(n35065) );
  XOR U34763 ( .A(n35247), .B(n35248), .Z(n35069) );
  AND U34764 ( .A(n603), .B(n35249), .Z(n35248) );
  XOR U34765 ( .A(n35250), .B(n35247), .Z(n35249) );
  XNOR U34766 ( .A(n35243), .B(n35178), .Z(n35245) );
  XOR U34767 ( .A(n35251), .B(n35252), .Z(n35178) );
  AND U34768 ( .A(n611), .B(n35213), .Z(n35252) );
  XOR U34769 ( .A(n35211), .B(n35251), .Z(n35213) );
  XOR U34770 ( .A(n35253), .B(n35254), .Z(n35243) );
  AND U34771 ( .A(n35255), .B(n35256), .Z(n35254) );
  XNOR U34772 ( .A(n35253), .B(n35081), .Z(n35256) );
  IV U34773 ( .A(n35084), .Z(n35081) );
  XOR U34774 ( .A(n35257), .B(n35258), .Z(n35084) );
  AND U34775 ( .A(n603), .B(n35259), .Z(n35258) );
  XOR U34776 ( .A(n35260), .B(n35257), .Z(n35259) );
  XOR U34777 ( .A(n35085), .B(n35253), .Z(n35255) );
  XOR U34778 ( .A(n35261), .B(n35262), .Z(n35085) );
  AND U34779 ( .A(n611), .B(n35221), .Z(n35262) );
  XOR U34780 ( .A(n35261), .B(n35219), .Z(n35221) );
  XOR U34781 ( .A(n35263), .B(n35264), .Z(n35253) );
  AND U34782 ( .A(n35265), .B(n35266), .Z(n35264) );
  XNOR U34783 ( .A(n35263), .B(n35109), .Z(n35266) );
  IV U34784 ( .A(n35112), .Z(n35109) );
  XOR U34785 ( .A(n35267), .B(n35268), .Z(n35112) );
  AND U34786 ( .A(n603), .B(n35269), .Z(n35268) );
  XNOR U34787 ( .A(n35270), .B(n35267), .Z(n35269) );
  XOR U34788 ( .A(n35113), .B(n35263), .Z(n35265) );
  XOR U34789 ( .A(n35271), .B(n35272), .Z(n35113) );
  AND U34790 ( .A(n611), .B(n35230), .Z(n35272) );
  XOR U34791 ( .A(n35271), .B(n35228), .Z(n35230) );
  XOR U34792 ( .A(n35187), .B(n35273), .Z(n35263) );
  AND U34793 ( .A(n35189), .B(n35274), .Z(n35273) );
  XNOR U34794 ( .A(n35187), .B(n35158), .Z(n35274) );
  IV U34795 ( .A(n35161), .Z(n35158) );
  XOR U34796 ( .A(n35275), .B(n35276), .Z(n35161) );
  AND U34797 ( .A(n603), .B(n35277), .Z(n35276) );
  XOR U34798 ( .A(n35278), .B(n35275), .Z(n35277) );
  XOR U34799 ( .A(n35162), .B(n35187), .Z(n35189) );
  XOR U34800 ( .A(n35279), .B(n35280), .Z(n35162) );
  AND U34801 ( .A(n611), .B(n35240), .Z(n35280) );
  XOR U34802 ( .A(n35279), .B(n35238), .Z(n35240) );
  AND U34803 ( .A(n35241), .B(n35171), .Z(n35187) );
  XNOR U34804 ( .A(n35281), .B(n35282), .Z(n35171) );
  AND U34805 ( .A(n603), .B(n35283), .Z(n35282) );
  XNOR U34806 ( .A(n35284), .B(n35281), .Z(n35283) );
  XNOR U34807 ( .A(n35285), .B(n35286), .Z(n603) );
  AND U34808 ( .A(n35287), .B(n35288), .Z(n35286) );
  XOR U34809 ( .A(n35250), .B(n35285), .Z(n35288) );
  AND U34810 ( .A(n35289), .B(n35290), .Z(n35250) );
  XNOR U34811 ( .A(n35247), .B(n35285), .Z(n35287) );
  XNOR U34812 ( .A(n35291), .B(n35292), .Z(n35247) );
  AND U34813 ( .A(n607), .B(n35293), .Z(n35292) );
  XNOR U34814 ( .A(n35294), .B(n35295), .Z(n35293) );
  XOR U34815 ( .A(n35296), .B(n35297), .Z(n35285) );
  AND U34816 ( .A(n35298), .B(n35299), .Z(n35297) );
  XNOR U34817 ( .A(n35296), .B(n35289), .Z(n35299) );
  IV U34818 ( .A(n35260), .Z(n35289) );
  XOR U34819 ( .A(n35300), .B(n35301), .Z(n35260) );
  XOR U34820 ( .A(n35302), .B(n35290), .Z(n35301) );
  AND U34821 ( .A(n35270), .B(n35303), .Z(n35290) );
  AND U34822 ( .A(n35304), .B(n35305), .Z(n35302) );
  XOR U34823 ( .A(n35306), .B(n35300), .Z(n35304) );
  XNOR U34824 ( .A(n35257), .B(n35296), .Z(n35298) );
  XNOR U34825 ( .A(n35307), .B(n35308), .Z(n35257) );
  AND U34826 ( .A(n607), .B(n35309), .Z(n35308) );
  XNOR U34827 ( .A(n35310), .B(n35311), .Z(n35309) );
  XOR U34828 ( .A(n35312), .B(n35313), .Z(n35296) );
  AND U34829 ( .A(n35314), .B(n35315), .Z(n35313) );
  XNOR U34830 ( .A(n35312), .B(n35270), .Z(n35315) );
  XOR U34831 ( .A(n35316), .B(n35305), .Z(n35270) );
  XNOR U34832 ( .A(n35317), .B(n35300), .Z(n35305) );
  XOR U34833 ( .A(n35318), .B(n35319), .Z(n35300) );
  AND U34834 ( .A(n35320), .B(n35321), .Z(n35319) );
  XOR U34835 ( .A(n35322), .B(n35318), .Z(n35320) );
  XNOR U34836 ( .A(n35323), .B(n35324), .Z(n35317) );
  AND U34837 ( .A(n35325), .B(n35326), .Z(n35324) );
  XOR U34838 ( .A(n35323), .B(n35327), .Z(n35325) );
  XNOR U34839 ( .A(n35306), .B(n35303), .Z(n35316) );
  AND U34840 ( .A(n35328), .B(n35329), .Z(n35303) );
  XOR U34841 ( .A(n35330), .B(n35331), .Z(n35306) );
  AND U34842 ( .A(n35332), .B(n35333), .Z(n35331) );
  XOR U34843 ( .A(n35330), .B(n35334), .Z(n35332) );
  XNOR U34844 ( .A(n35267), .B(n35312), .Z(n35314) );
  XNOR U34845 ( .A(n35335), .B(n35336), .Z(n35267) );
  AND U34846 ( .A(n607), .B(n35337), .Z(n35336) );
  XNOR U34847 ( .A(n35338), .B(n35339), .Z(n35337) );
  XOR U34848 ( .A(n35340), .B(n35341), .Z(n35312) );
  AND U34849 ( .A(n35342), .B(n35343), .Z(n35341) );
  XNOR U34850 ( .A(n35340), .B(n35328), .Z(n35343) );
  IV U34851 ( .A(n35278), .Z(n35328) );
  XNOR U34852 ( .A(n35344), .B(n35321), .Z(n35278) );
  XNOR U34853 ( .A(n35345), .B(n35327), .Z(n35321) );
  XOR U34854 ( .A(n35346), .B(n35347), .Z(n35327) );
  NOR U34855 ( .A(n35348), .B(n35349), .Z(n35347) );
  XNOR U34856 ( .A(n35346), .B(n35350), .Z(n35348) );
  XNOR U34857 ( .A(n35326), .B(n35318), .Z(n35345) );
  XOR U34858 ( .A(n35351), .B(n35352), .Z(n35318) );
  AND U34859 ( .A(n35353), .B(n35354), .Z(n35352) );
  XNOR U34860 ( .A(n35351), .B(n35355), .Z(n35353) );
  XNOR U34861 ( .A(n35356), .B(n35323), .Z(n35326) );
  XOR U34862 ( .A(n35357), .B(n35358), .Z(n35323) );
  AND U34863 ( .A(n35359), .B(n35360), .Z(n35358) );
  XOR U34864 ( .A(n35357), .B(n35361), .Z(n35359) );
  XNOR U34865 ( .A(n35362), .B(n35363), .Z(n35356) );
  NOR U34866 ( .A(n35364), .B(n35365), .Z(n35363) );
  XOR U34867 ( .A(n35362), .B(n35366), .Z(n35364) );
  XNOR U34868 ( .A(n35322), .B(n35329), .Z(n35344) );
  NOR U34869 ( .A(n35284), .B(n35367), .Z(n35329) );
  XOR U34870 ( .A(n35334), .B(n35333), .Z(n35322) );
  XNOR U34871 ( .A(n35368), .B(n35330), .Z(n35333) );
  XOR U34872 ( .A(n35369), .B(n35370), .Z(n35330) );
  AND U34873 ( .A(n35371), .B(n35372), .Z(n35370) );
  XOR U34874 ( .A(n35369), .B(n35373), .Z(n35371) );
  XNOR U34875 ( .A(n35374), .B(n35375), .Z(n35368) );
  NOR U34876 ( .A(n35376), .B(n35377), .Z(n35375) );
  XNOR U34877 ( .A(n35374), .B(n35378), .Z(n35376) );
  XOR U34878 ( .A(n35379), .B(n35380), .Z(n35334) );
  NOR U34879 ( .A(n35381), .B(n35382), .Z(n35380) );
  XNOR U34880 ( .A(n35379), .B(n35383), .Z(n35381) );
  XNOR U34881 ( .A(n35275), .B(n35340), .Z(n35342) );
  XNOR U34882 ( .A(n35384), .B(n35385), .Z(n35275) );
  AND U34883 ( .A(n607), .B(n35386), .Z(n35385) );
  XNOR U34884 ( .A(n35387), .B(n35388), .Z(n35386) );
  AND U34885 ( .A(n35281), .B(n35284), .Z(n35340) );
  XOR U34886 ( .A(n35389), .B(n35367), .Z(n35284) );
  XNOR U34887 ( .A(p_input[2048]), .B(p_input[448]), .Z(n35367) );
  XOR U34888 ( .A(n35355), .B(n35354), .Z(n35389) );
  XNOR U34889 ( .A(n35390), .B(n35361), .Z(n35354) );
  XNOR U34890 ( .A(n35350), .B(n35349), .Z(n35361) );
  XOR U34891 ( .A(n35391), .B(n35346), .Z(n35349) );
  XNOR U34892 ( .A(n29266), .B(p_input[458]), .Z(n35346) );
  XNOR U34893 ( .A(p_input[2059]), .B(p_input[459]), .Z(n35391) );
  XOR U34894 ( .A(p_input[2060]), .B(p_input[460]), .Z(n35350) );
  XNOR U34895 ( .A(n35360), .B(n35351), .Z(n35390) );
  XNOR U34896 ( .A(n29494), .B(p_input[449]), .Z(n35351) );
  XOR U34897 ( .A(n35392), .B(n35366), .Z(n35360) );
  XNOR U34898 ( .A(p_input[2063]), .B(p_input[463]), .Z(n35366) );
  XOR U34899 ( .A(n35357), .B(n35365), .Z(n35392) );
  XOR U34900 ( .A(n35393), .B(n35362), .Z(n35365) );
  XOR U34901 ( .A(p_input[2061]), .B(p_input[461]), .Z(n35362) );
  XNOR U34902 ( .A(p_input[2062]), .B(p_input[462]), .Z(n35393) );
  XNOR U34903 ( .A(n29036), .B(p_input[457]), .Z(n35357) );
  XNOR U34904 ( .A(n35373), .B(n35372), .Z(n35355) );
  XNOR U34905 ( .A(n35394), .B(n35378), .Z(n35372) );
  XOR U34906 ( .A(p_input[2056]), .B(p_input[456]), .Z(n35378) );
  XOR U34907 ( .A(n35369), .B(n35377), .Z(n35394) );
  XOR U34908 ( .A(n35395), .B(n35374), .Z(n35377) );
  XOR U34909 ( .A(p_input[2054]), .B(p_input[454]), .Z(n35374) );
  XNOR U34910 ( .A(p_input[2055]), .B(p_input[455]), .Z(n35395) );
  XNOR U34911 ( .A(n29039), .B(p_input[450]), .Z(n35369) );
  XNOR U34912 ( .A(n35383), .B(n35382), .Z(n35373) );
  XOR U34913 ( .A(n35396), .B(n35379), .Z(n35382) );
  XOR U34914 ( .A(p_input[2051]), .B(p_input[451]), .Z(n35379) );
  XNOR U34915 ( .A(p_input[2052]), .B(p_input[452]), .Z(n35396) );
  XOR U34916 ( .A(p_input[2053]), .B(p_input[453]), .Z(n35383) );
  XNOR U34917 ( .A(n35397), .B(n35398), .Z(n35281) );
  AND U34918 ( .A(n607), .B(n35399), .Z(n35398) );
  XNOR U34919 ( .A(n35400), .B(n35401), .Z(n607) );
  AND U34920 ( .A(n35402), .B(n35403), .Z(n35401) );
  XOR U34921 ( .A(n35295), .B(n35400), .Z(n35403) );
  XNOR U34922 ( .A(n35404), .B(n35400), .Z(n35402) );
  XOR U34923 ( .A(n35405), .B(n35406), .Z(n35400) );
  AND U34924 ( .A(n35407), .B(n35408), .Z(n35406) );
  XOR U34925 ( .A(n35310), .B(n35405), .Z(n35408) );
  XOR U34926 ( .A(n35405), .B(n35311), .Z(n35407) );
  XOR U34927 ( .A(n35409), .B(n35410), .Z(n35405) );
  AND U34928 ( .A(n35411), .B(n35412), .Z(n35410) );
  XOR U34929 ( .A(n35338), .B(n35409), .Z(n35412) );
  XOR U34930 ( .A(n35409), .B(n35339), .Z(n35411) );
  XOR U34931 ( .A(n35413), .B(n35414), .Z(n35409) );
  AND U34932 ( .A(n35415), .B(n35416), .Z(n35414) );
  XOR U34933 ( .A(n35413), .B(n35387), .Z(n35416) );
  XNOR U34934 ( .A(n35417), .B(n35418), .Z(n35241) );
  AND U34935 ( .A(n611), .B(n35419), .Z(n35418) );
  XNOR U34936 ( .A(n35420), .B(n35421), .Z(n611) );
  AND U34937 ( .A(n35422), .B(n35423), .Z(n35421) );
  XOR U34938 ( .A(n35420), .B(n35251), .Z(n35423) );
  XNOR U34939 ( .A(n35420), .B(n35211), .Z(n35422) );
  XOR U34940 ( .A(n35424), .B(n35425), .Z(n35420) );
  AND U34941 ( .A(n35426), .B(n35427), .Z(n35425) );
  XOR U34942 ( .A(n35424), .B(n35219), .Z(n35426) );
  XOR U34943 ( .A(n35428), .B(n35429), .Z(n35202) );
  AND U34944 ( .A(n615), .B(n35419), .Z(n35429) );
  XNOR U34945 ( .A(n35417), .B(n35428), .Z(n35419) );
  XNOR U34946 ( .A(n35430), .B(n35431), .Z(n615) );
  AND U34947 ( .A(n35432), .B(n35433), .Z(n35431) );
  XNOR U34948 ( .A(n35434), .B(n35430), .Z(n35433) );
  IV U34949 ( .A(n35251), .Z(n35434) );
  XOR U34950 ( .A(n35404), .B(n35435), .Z(n35251) );
  AND U34951 ( .A(n618), .B(n35436), .Z(n35435) );
  XOR U34952 ( .A(n35294), .B(n35291), .Z(n35436) );
  IV U34953 ( .A(n35404), .Z(n35294) );
  XNOR U34954 ( .A(n35211), .B(n35430), .Z(n35432) );
  XOR U34955 ( .A(n35437), .B(n35438), .Z(n35211) );
  AND U34956 ( .A(n634), .B(n35439), .Z(n35438) );
  XOR U34957 ( .A(n35424), .B(n35440), .Z(n35430) );
  AND U34958 ( .A(n35441), .B(n35427), .Z(n35440) );
  XNOR U34959 ( .A(n35261), .B(n35424), .Z(n35427) );
  XOR U34960 ( .A(n35311), .B(n35442), .Z(n35261) );
  AND U34961 ( .A(n618), .B(n35443), .Z(n35442) );
  XOR U34962 ( .A(n35307), .B(n35311), .Z(n35443) );
  XNOR U34963 ( .A(n35444), .B(n35424), .Z(n35441) );
  IV U34964 ( .A(n35219), .Z(n35444) );
  XOR U34965 ( .A(n35445), .B(n35446), .Z(n35219) );
  AND U34966 ( .A(n634), .B(n35447), .Z(n35446) );
  XOR U34967 ( .A(n35448), .B(n35449), .Z(n35424) );
  AND U34968 ( .A(n35450), .B(n35451), .Z(n35449) );
  XNOR U34969 ( .A(n35271), .B(n35448), .Z(n35451) );
  XOR U34970 ( .A(n35339), .B(n35452), .Z(n35271) );
  AND U34971 ( .A(n618), .B(n35453), .Z(n35452) );
  XOR U34972 ( .A(n35335), .B(n35339), .Z(n35453) );
  XOR U34973 ( .A(n35448), .B(n35228), .Z(n35450) );
  XOR U34974 ( .A(n35454), .B(n35455), .Z(n35228) );
  AND U34975 ( .A(n634), .B(n35456), .Z(n35455) );
  XOR U34976 ( .A(n35457), .B(n35458), .Z(n35448) );
  AND U34977 ( .A(n35459), .B(n35460), .Z(n35458) );
  XNOR U34978 ( .A(n35457), .B(n35279), .Z(n35460) );
  XOR U34979 ( .A(n35388), .B(n35461), .Z(n35279) );
  AND U34980 ( .A(n618), .B(n35462), .Z(n35461) );
  XOR U34981 ( .A(n35384), .B(n35388), .Z(n35462) );
  XNOR U34982 ( .A(n35463), .B(n35457), .Z(n35459) );
  IV U34983 ( .A(n35238), .Z(n35463) );
  XOR U34984 ( .A(n35464), .B(n35465), .Z(n35238) );
  AND U34985 ( .A(n634), .B(n35466), .Z(n35465) );
  AND U34986 ( .A(n35428), .B(n35417), .Z(n35457) );
  XNOR U34987 ( .A(n35467), .B(n35468), .Z(n35417) );
  AND U34988 ( .A(n618), .B(n35399), .Z(n35468) );
  XNOR U34989 ( .A(n35397), .B(n35467), .Z(n35399) );
  XNOR U34990 ( .A(n35469), .B(n35470), .Z(n618) );
  AND U34991 ( .A(n35471), .B(n35472), .Z(n35470) );
  XNOR U34992 ( .A(n35469), .B(n35291), .Z(n35472) );
  IV U34993 ( .A(n35295), .Z(n35291) );
  XOR U34994 ( .A(n35473), .B(n35474), .Z(n35295) );
  AND U34995 ( .A(n622), .B(n35475), .Z(n35474) );
  XOR U34996 ( .A(n35476), .B(n35473), .Z(n35475) );
  XNOR U34997 ( .A(n35469), .B(n35404), .Z(n35471) );
  XOR U34998 ( .A(n35477), .B(n35478), .Z(n35404) );
  AND U34999 ( .A(n630), .B(n35439), .Z(n35478) );
  XOR U35000 ( .A(n35437), .B(n35477), .Z(n35439) );
  XOR U35001 ( .A(n35479), .B(n35480), .Z(n35469) );
  AND U35002 ( .A(n35481), .B(n35482), .Z(n35480) );
  XNOR U35003 ( .A(n35479), .B(n35307), .Z(n35482) );
  IV U35004 ( .A(n35310), .Z(n35307) );
  XOR U35005 ( .A(n35483), .B(n35484), .Z(n35310) );
  AND U35006 ( .A(n622), .B(n35485), .Z(n35484) );
  XOR U35007 ( .A(n35486), .B(n35483), .Z(n35485) );
  XOR U35008 ( .A(n35311), .B(n35479), .Z(n35481) );
  XOR U35009 ( .A(n35487), .B(n35488), .Z(n35311) );
  AND U35010 ( .A(n630), .B(n35447), .Z(n35488) );
  XOR U35011 ( .A(n35487), .B(n35445), .Z(n35447) );
  XOR U35012 ( .A(n35489), .B(n35490), .Z(n35479) );
  AND U35013 ( .A(n35491), .B(n35492), .Z(n35490) );
  XNOR U35014 ( .A(n35489), .B(n35335), .Z(n35492) );
  IV U35015 ( .A(n35338), .Z(n35335) );
  XOR U35016 ( .A(n35493), .B(n35494), .Z(n35338) );
  AND U35017 ( .A(n622), .B(n35495), .Z(n35494) );
  XNOR U35018 ( .A(n35496), .B(n35493), .Z(n35495) );
  XOR U35019 ( .A(n35339), .B(n35489), .Z(n35491) );
  XOR U35020 ( .A(n35497), .B(n35498), .Z(n35339) );
  AND U35021 ( .A(n630), .B(n35456), .Z(n35498) );
  XOR U35022 ( .A(n35497), .B(n35454), .Z(n35456) );
  XOR U35023 ( .A(n35413), .B(n35499), .Z(n35489) );
  AND U35024 ( .A(n35415), .B(n35500), .Z(n35499) );
  XNOR U35025 ( .A(n35413), .B(n35384), .Z(n35500) );
  IV U35026 ( .A(n35387), .Z(n35384) );
  XOR U35027 ( .A(n35501), .B(n35502), .Z(n35387) );
  AND U35028 ( .A(n622), .B(n35503), .Z(n35502) );
  XOR U35029 ( .A(n35504), .B(n35501), .Z(n35503) );
  XOR U35030 ( .A(n35388), .B(n35413), .Z(n35415) );
  XOR U35031 ( .A(n35505), .B(n35506), .Z(n35388) );
  AND U35032 ( .A(n630), .B(n35466), .Z(n35506) );
  XOR U35033 ( .A(n35505), .B(n35464), .Z(n35466) );
  AND U35034 ( .A(n35467), .B(n35397), .Z(n35413) );
  XNOR U35035 ( .A(n35507), .B(n35508), .Z(n35397) );
  AND U35036 ( .A(n622), .B(n35509), .Z(n35508) );
  XNOR U35037 ( .A(n35510), .B(n35507), .Z(n35509) );
  XNOR U35038 ( .A(n35511), .B(n35512), .Z(n622) );
  AND U35039 ( .A(n35513), .B(n35514), .Z(n35512) );
  XOR U35040 ( .A(n35476), .B(n35511), .Z(n35514) );
  AND U35041 ( .A(n35515), .B(n35516), .Z(n35476) );
  XNOR U35042 ( .A(n35473), .B(n35511), .Z(n35513) );
  XNOR U35043 ( .A(n35517), .B(n35518), .Z(n35473) );
  AND U35044 ( .A(n626), .B(n35519), .Z(n35518) );
  XNOR U35045 ( .A(n35520), .B(n35521), .Z(n35519) );
  XOR U35046 ( .A(n35522), .B(n35523), .Z(n35511) );
  AND U35047 ( .A(n35524), .B(n35525), .Z(n35523) );
  XNOR U35048 ( .A(n35522), .B(n35515), .Z(n35525) );
  IV U35049 ( .A(n35486), .Z(n35515) );
  XOR U35050 ( .A(n35526), .B(n35527), .Z(n35486) );
  XOR U35051 ( .A(n35528), .B(n35516), .Z(n35527) );
  AND U35052 ( .A(n35496), .B(n35529), .Z(n35516) );
  AND U35053 ( .A(n35530), .B(n35531), .Z(n35528) );
  XOR U35054 ( .A(n35532), .B(n35526), .Z(n35530) );
  XNOR U35055 ( .A(n35483), .B(n35522), .Z(n35524) );
  XNOR U35056 ( .A(n35533), .B(n35534), .Z(n35483) );
  AND U35057 ( .A(n626), .B(n35535), .Z(n35534) );
  XNOR U35058 ( .A(n35536), .B(n35537), .Z(n35535) );
  XOR U35059 ( .A(n35538), .B(n35539), .Z(n35522) );
  AND U35060 ( .A(n35540), .B(n35541), .Z(n35539) );
  XNOR U35061 ( .A(n35538), .B(n35496), .Z(n35541) );
  XOR U35062 ( .A(n35542), .B(n35531), .Z(n35496) );
  XNOR U35063 ( .A(n35543), .B(n35526), .Z(n35531) );
  XOR U35064 ( .A(n35544), .B(n35545), .Z(n35526) );
  AND U35065 ( .A(n35546), .B(n35547), .Z(n35545) );
  XOR U35066 ( .A(n35548), .B(n35544), .Z(n35546) );
  XNOR U35067 ( .A(n35549), .B(n35550), .Z(n35543) );
  AND U35068 ( .A(n35551), .B(n35552), .Z(n35550) );
  XOR U35069 ( .A(n35549), .B(n35553), .Z(n35551) );
  XNOR U35070 ( .A(n35532), .B(n35529), .Z(n35542) );
  AND U35071 ( .A(n35554), .B(n35555), .Z(n35529) );
  XOR U35072 ( .A(n35556), .B(n35557), .Z(n35532) );
  AND U35073 ( .A(n35558), .B(n35559), .Z(n35557) );
  XOR U35074 ( .A(n35556), .B(n35560), .Z(n35558) );
  XNOR U35075 ( .A(n35493), .B(n35538), .Z(n35540) );
  XNOR U35076 ( .A(n35561), .B(n35562), .Z(n35493) );
  AND U35077 ( .A(n626), .B(n35563), .Z(n35562) );
  XNOR U35078 ( .A(n35564), .B(n35565), .Z(n35563) );
  XOR U35079 ( .A(n35566), .B(n35567), .Z(n35538) );
  AND U35080 ( .A(n35568), .B(n35569), .Z(n35567) );
  XNOR U35081 ( .A(n35566), .B(n35554), .Z(n35569) );
  IV U35082 ( .A(n35504), .Z(n35554) );
  XNOR U35083 ( .A(n35570), .B(n35547), .Z(n35504) );
  XNOR U35084 ( .A(n35571), .B(n35553), .Z(n35547) );
  XOR U35085 ( .A(n35572), .B(n35573), .Z(n35553) );
  NOR U35086 ( .A(n35574), .B(n35575), .Z(n35573) );
  XNOR U35087 ( .A(n35572), .B(n35576), .Z(n35574) );
  XNOR U35088 ( .A(n35552), .B(n35544), .Z(n35571) );
  XOR U35089 ( .A(n35577), .B(n35578), .Z(n35544) );
  AND U35090 ( .A(n35579), .B(n35580), .Z(n35578) );
  XNOR U35091 ( .A(n35577), .B(n35581), .Z(n35579) );
  XNOR U35092 ( .A(n35582), .B(n35549), .Z(n35552) );
  XOR U35093 ( .A(n35583), .B(n35584), .Z(n35549) );
  AND U35094 ( .A(n35585), .B(n35586), .Z(n35584) );
  XOR U35095 ( .A(n35583), .B(n35587), .Z(n35585) );
  XNOR U35096 ( .A(n35588), .B(n35589), .Z(n35582) );
  NOR U35097 ( .A(n35590), .B(n35591), .Z(n35589) );
  XOR U35098 ( .A(n35588), .B(n35592), .Z(n35590) );
  XNOR U35099 ( .A(n35548), .B(n35555), .Z(n35570) );
  NOR U35100 ( .A(n35510), .B(n35593), .Z(n35555) );
  XOR U35101 ( .A(n35560), .B(n35559), .Z(n35548) );
  XNOR U35102 ( .A(n35594), .B(n35556), .Z(n35559) );
  XOR U35103 ( .A(n35595), .B(n35596), .Z(n35556) );
  AND U35104 ( .A(n35597), .B(n35598), .Z(n35596) );
  XOR U35105 ( .A(n35595), .B(n35599), .Z(n35597) );
  XNOR U35106 ( .A(n35600), .B(n35601), .Z(n35594) );
  NOR U35107 ( .A(n35602), .B(n35603), .Z(n35601) );
  XNOR U35108 ( .A(n35600), .B(n35604), .Z(n35602) );
  XOR U35109 ( .A(n35605), .B(n35606), .Z(n35560) );
  NOR U35110 ( .A(n35607), .B(n35608), .Z(n35606) );
  XNOR U35111 ( .A(n35605), .B(n35609), .Z(n35607) );
  XNOR U35112 ( .A(n35501), .B(n35566), .Z(n35568) );
  XNOR U35113 ( .A(n35610), .B(n35611), .Z(n35501) );
  AND U35114 ( .A(n626), .B(n35612), .Z(n35611) );
  XNOR U35115 ( .A(n35613), .B(n35614), .Z(n35612) );
  AND U35116 ( .A(n35507), .B(n35510), .Z(n35566) );
  XOR U35117 ( .A(n35615), .B(n35593), .Z(n35510) );
  XNOR U35118 ( .A(p_input[2048]), .B(p_input[464]), .Z(n35593) );
  XOR U35119 ( .A(n35581), .B(n35580), .Z(n35615) );
  XNOR U35120 ( .A(n35616), .B(n35587), .Z(n35580) );
  XNOR U35121 ( .A(n35576), .B(n35575), .Z(n35587) );
  XOR U35122 ( .A(n35617), .B(n35572), .Z(n35575) );
  XNOR U35123 ( .A(n29266), .B(p_input[474]), .Z(n35572) );
  XNOR U35124 ( .A(p_input[2059]), .B(p_input[475]), .Z(n35617) );
  XOR U35125 ( .A(p_input[2060]), .B(p_input[476]), .Z(n35576) );
  XNOR U35126 ( .A(n35586), .B(n35577), .Z(n35616) );
  XNOR U35127 ( .A(n29494), .B(p_input[465]), .Z(n35577) );
  XOR U35128 ( .A(n35618), .B(n35592), .Z(n35586) );
  XNOR U35129 ( .A(p_input[2063]), .B(p_input[479]), .Z(n35592) );
  XOR U35130 ( .A(n35583), .B(n35591), .Z(n35618) );
  XOR U35131 ( .A(n35619), .B(n35588), .Z(n35591) );
  XOR U35132 ( .A(p_input[2061]), .B(p_input[477]), .Z(n35588) );
  XNOR U35133 ( .A(p_input[2062]), .B(p_input[478]), .Z(n35619) );
  XNOR U35134 ( .A(n29036), .B(p_input[473]), .Z(n35583) );
  XNOR U35135 ( .A(n35599), .B(n35598), .Z(n35581) );
  XNOR U35136 ( .A(n35620), .B(n35604), .Z(n35598) );
  XOR U35137 ( .A(p_input[2056]), .B(p_input[472]), .Z(n35604) );
  XOR U35138 ( .A(n35595), .B(n35603), .Z(n35620) );
  XOR U35139 ( .A(n35621), .B(n35600), .Z(n35603) );
  XOR U35140 ( .A(p_input[2054]), .B(p_input[470]), .Z(n35600) );
  XNOR U35141 ( .A(p_input[2055]), .B(p_input[471]), .Z(n35621) );
  XNOR U35142 ( .A(n29039), .B(p_input[466]), .Z(n35595) );
  XNOR U35143 ( .A(n35609), .B(n35608), .Z(n35599) );
  XOR U35144 ( .A(n35622), .B(n35605), .Z(n35608) );
  XOR U35145 ( .A(p_input[2051]), .B(p_input[467]), .Z(n35605) );
  XNOR U35146 ( .A(p_input[2052]), .B(p_input[468]), .Z(n35622) );
  XOR U35147 ( .A(p_input[2053]), .B(p_input[469]), .Z(n35609) );
  XNOR U35148 ( .A(n35623), .B(n35624), .Z(n35507) );
  AND U35149 ( .A(n626), .B(n35625), .Z(n35624) );
  XNOR U35150 ( .A(n35626), .B(n35627), .Z(n626) );
  AND U35151 ( .A(n35628), .B(n35629), .Z(n35627) );
  XOR U35152 ( .A(n35521), .B(n35626), .Z(n35629) );
  XNOR U35153 ( .A(n35630), .B(n35626), .Z(n35628) );
  XOR U35154 ( .A(n35631), .B(n35632), .Z(n35626) );
  AND U35155 ( .A(n35633), .B(n35634), .Z(n35632) );
  XOR U35156 ( .A(n35536), .B(n35631), .Z(n35634) );
  XOR U35157 ( .A(n35631), .B(n35537), .Z(n35633) );
  XOR U35158 ( .A(n35635), .B(n35636), .Z(n35631) );
  AND U35159 ( .A(n35637), .B(n35638), .Z(n35636) );
  XOR U35160 ( .A(n35564), .B(n35635), .Z(n35638) );
  XOR U35161 ( .A(n35635), .B(n35565), .Z(n35637) );
  XOR U35162 ( .A(n35639), .B(n35640), .Z(n35635) );
  AND U35163 ( .A(n35641), .B(n35642), .Z(n35640) );
  XOR U35164 ( .A(n35639), .B(n35613), .Z(n35642) );
  XNOR U35165 ( .A(n35643), .B(n35644), .Z(n35467) );
  AND U35166 ( .A(n630), .B(n35645), .Z(n35644) );
  XNOR U35167 ( .A(n35646), .B(n35647), .Z(n630) );
  AND U35168 ( .A(n35648), .B(n35649), .Z(n35647) );
  XOR U35169 ( .A(n35646), .B(n35477), .Z(n35649) );
  XNOR U35170 ( .A(n35646), .B(n35437), .Z(n35648) );
  XOR U35171 ( .A(n35650), .B(n35651), .Z(n35646) );
  AND U35172 ( .A(n35652), .B(n35653), .Z(n35651) );
  XOR U35173 ( .A(n35650), .B(n35445), .Z(n35652) );
  XOR U35174 ( .A(n35654), .B(n35655), .Z(n35428) );
  AND U35175 ( .A(n634), .B(n35645), .Z(n35655) );
  XNOR U35176 ( .A(n35643), .B(n35654), .Z(n35645) );
  XNOR U35177 ( .A(n35656), .B(n35657), .Z(n634) );
  AND U35178 ( .A(n35658), .B(n35659), .Z(n35657) );
  XNOR U35179 ( .A(n35660), .B(n35656), .Z(n35659) );
  IV U35180 ( .A(n35477), .Z(n35660) );
  XOR U35181 ( .A(n35630), .B(n35661), .Z(n35477) );
  AND U35182 ( .A(n637), .B(n35662), .Z(n35661) );
  XOR U35183 ( .A(n35520), .B(n35517), .Z(n35662) );
  IV U35184 ( .A(n35630), .Z(n35520) );
  XNOR U35185 ( .A(n35437), .B(n35656), .Z(n35658) );
  XOR U35186 ( .A(n35663), .B(n35664), .Z(n35437) );
  AND U35187 ( .A(n653), .B(n35665), .Z(n35664) );
  XOR U35188 ( .A(n35650), .B(n35666), .Z(n35656) );
  AND U35189 ( .A(n35667), .B(n35653), .Z(n35666) );
  XNOR U35190 ( .A(n35487), .B(n35650), .Z(n35653) );
  XOR U35191 ( .A(n35537), .B(n35668), .Z(n35487) );
  AND U35192 ( .A(n637), .B(n35669), .Z(n35668) );
  XOR U35193 ( .A(n35533), .B(n35537), .Z(n35669) );
  XNOR U35194 ( .A(n35670), .B(n35650), .Z(n35667) );
  IV U35195 ( .A(n35445), .Z(n35670) );
  XOR U35196 ( .A(n35671), .B(n35672), .Z(n35445) );
  AND U35197 ( .A(n653), .B(n35673), .Z(n35672) );
  XOR U35198 ( .A(n35674), .B(n35675), .Z(n35650) );
  AND U35199 ( .A(n35676), .B(n35677), .Z(n35675) );
  XNOR U35200 ( .A(n35497), .B(n35674), .Z(n35677) );
  XOR U35201 ( .A(n35565), .B(n35678), .Z(n35497) );
  AND U35202 ( .A(n637), .B(n35679), .Z(n35678) );
  XOR U35203 ( .A(n35561), .B(n35565), .Z(n35679) );
  XOR U35204 ( .A(n35674), .B(n35454), .Z(n35676) );
  XOR U35205 ( .A(n35680), .B(n35681), .Z(n35454) );
  AND U35206 ( .A(n653), .B(n35682), .Z(n35681) );
  XOR U35207 ( .A(n35683), .B(n35684), .Z(n35674) );
  AND U35208 ( .A(n35685), .B(n35686), .Z(n35684) );
  XNOR U35209 ( .A(n35683), .B(n35505), .Z(n35686) );
  XOR U35210 ( .A(n35614), .B(n35687), .Z(n35505) );
  AND U35211 ( .A(n637), .B(n35688), .Z(n35687) );
  XOR U35212 ( .A(n35610), .B(n35614), .Z(n35688) );
  XNOR U35213 ( .A(n35689), .B(n35683), .Z(n35685) );
  IV U35214 ( .A(n35464), .Z(n35689) );
  XOR U35215 ( .A(n35690), .B(n35691), .Z(n35464) );
  AND U35216 ( .A(n653), .B(n35692), .Z(n35691) );
  AND U35217 ( .A(n35654), .B(n35643), .Z(n35683) );
  XNOR U35218 ( .A(n35693), .B(n35694), .Z(n35643) );
  AND U35219 ( .A(n637), .B(n35625), .Z(n35694) );
  XNOR U35220 ( .A(n35623), .B(n35693), .Z(n35625) );
  XNOR U35221 ( .A(n35695), .B(n35696), .Z(n637) );
  AND U35222 ( .A(n35697), .B(n35698), .Z(n35696) );
  XNOR U35223 ( .A(n35695), .B(n35517), .Z(n35698) );
  IV U35224 ( .A(n35521), .Z(n35517) );
  XOR U35225 ( .A(n35699), .B(n35700), .Z(n35521) );
  AND U35226 ( .A(n641), .B(n35701), .Z(n35700) );
  XOR U35227 ( .A(n35702), .B(n35699), .Z(n35701) );
  XNOR U35228 ( .A(n35695), .B(n35630), .Z(n35697) );
  XOR U35229 ( .A(n35703), .B(n35704), .Z(n35630) );
  AND U35230 ( .A(n649), .B(n35665), .Z(n35704) );
  XOR U35231 ( .A(n35663), .B(n35703), .Z(n35665) );
  XOR U35232 ( .A(n35705), .B(n35706), .Z(n35695) );
  AND U35233 ( .A(n35707), .B(n35708), .Z(n35706) );
  XNOR U35234 ( .A(n35705), .B(n35533), .Z(n35708) );
  IV U35235 ( .A(n35536), .Z(n35533) );
  XOR U35236 ( .A(n35709), .B(n35710), .Z(n35536) );
  AND U35237 ( .A(n641), .B(n35711), .Z(n35710) );
  XOR U35238 ( .A(n35712), .B(n35709), .Z(n35711) );
  XOR U35239 ( .A(n35537), .B(n35705), .Z(n35707) );
  XOR U35240 ( .A(n35713), .B(n35714), .Z(n35537) );
  AND U35241 ( .A(n649), .B(n35673), .Z(n35714) );
  XOR U35242 ( .A(n35713), .B(n35671), .Z(n35673) );
  XOR U35243 ( .A(n35715), .B(n35716), .Z(n35705) );
  AND U35244 ( .A(n35717), .B(n35718), .Z(n35716) );
  XNOR U35245 ( .A(n35715), .B(n35561), .Z(n35718) );
  IV U35246 ( .A(n35564), .Z(n35561) );
  XOR U35247 ( .A(n35719), .B(n35720), .Z(n35564) );
  AND U35248 ( .A(n641), .B(n35721), .Z(n35720) );
  XNOR U35249 ( .A(n35722), .B(n35719), .Z(n35721) );
  XOR U35250 ( .A(n35565), .B(n35715), .Z(n35717) );
  XOR U35251 ( .A(n35723), .B(n35724), .Z(n35565) );
  AND U35252 ( .A(n649), .B(n35682), .Z(n35724) );
  XOR U35253 ( .A(n35723), .B(n35680), .Z(n35682) );
  XOR U35254 ( .A(n35639), .B(n35725), .Z(n35715) );
  AND U35255 ( .A(n35641), .B(n35726), .Z(n35725) );
  XNOR U35256 ( .A(n35639), .B(n35610), .Z(n35726) );
  IV U35257 ( .A(n35613), .Z(n35610) );
  XOR U35258 ( .A(n35727), .B(n35728), .Z(n35613) );
  AND U35259 ( .A(n641), .B(n35729), .Z(n35728) );
  XOR U35260 ( .A(n35730), .B(n35727), .Z(n35729) );
  XOR U35261 ( .A(n35614), .B(n35639), .Z(n35641) );
  XOR U35262 ( .A(n35731), .B(n35732), .Z(n35614) );
  AND U35263 ( .A(n649), .B(n35692), .Z(n35732) );
  XOR U35264 ( .A(n35731), .B(n35690), .Z(n35692) );
  AND U35265 ( .A(n35693), .B(n35623), .Z(n35639) );
  XNOR U35266 ( .A(n35733), .B(n35734), .Z(n35623) );
  AND U35267 ( .A(n641), .B(n35735), .Z(n35734) );
  XNOR U35268 ( .A(n35736), .B(n35733), .Z(n35735) );
  XNOR U35269 ( .A(n35737), .B(n35738), .Z(n641) );
  AND U35270 ( .A(n35739), .B(n35740), .Z(n35738) );
  XOR U35271 ( .A(n35702), .B(n35737), .Z(n35740) );
  AND U35272 ( .A(n35741), .B(n35742), .Z(n35702) );
  XNOR U35273 ( .A(n35699), .B(n35737), .Z(n35739) );
  XNOR U35274 ( .A(n35743), .B(n35744), .Z(n35699) );
  AND U35275 ( .A(n645), .B(n35745), .Z(n35744) );
  XNOR U35276 ( .A(n35746), .B(n35747), .Z(n35745) );
  XOR U35277 ( .A(n35748), .B(n35749), .Z(n35737) );
  AND U35278 ( .A(n35750), .B(n35751), .Z(n35749) );
  XNOR U35279 ( .A(n35748), .B(n35741), .Z(n35751) );
  IV U35280 ( .A(n35712), .Z(n35741) );
  XOR U35281 ( .A(n35752), .B(n35753), .Z(n35712) );
  XOR U35282 ( .A(n35754), .B(n35742), .Z(n35753) );
  AND U35283 ( .A(n35722), .B(n35755), .Z(n35742) );
  AND U35284 ( .A(n35756), .B(n35757), .Z(n35754) );
  XOR U35285 ( .A(n35758), .B(n35752), .Z(n35756) );
  XNOR U35286 ( .A(n35709), .B(n35748), .Z(n35750) );
  XNOR U35287 ( .A(n35759), .B(n35760), .Z(n35709) );
  AND U35288 ( .A(n645), .B(n35761), .Z(n35760) );
  XNOR U35289 ( .A(n35762), .B(n35763), .Z(n35761) );
  XOR U35290 ( .A(n35764), .B(n35765), .Z(n35748) );
  AND U35291 ( .A(n35766), .B(n35767), .Z(n35765) );
  XNOR U35292 ( .A(n35764), .B(n35722), .Z(n35767) );
  XOR U35293 ( .A(n35768), .B(n35757), .Z(n35722) );
  XNOR U35294 ( .A(n35769), .B(n35752), .Z(n35757) );
  XOR U35295 ( .A(n35770), .B(n35771), .Z(n35752) );
  AND U35296 ( .A(n35772), .B(n35773), .Z(n35771) );
  XOR U35297 ( .A(n35774), .B(n35770), .Z(n35772) );
  XNOR U35298 ( .A(n35775), .B(n35776), .Z(n35769) );
  AND U35299 ( .A(n35777), .B(n35778), .Z(n35776) );
  XOR U35300 ( .A(n35775), .B(n35779), .Z(n35777) );
  XNOR U35301 ( .A(n35758), .B(n35755), .Z(n35768) );
  AND U35302 ( .A(n35780), .B(n35781), .Z(n35755) );
  XOR U35303 ( .A(n35782), .B(n35783), .Z(n35758) );
  AND U35304 ( .A(n35784), .B(n35785), .Z(n35783) );
  XOR U35305 ( .A(n35782), .B(n35786), .Z(n35784) );
  XNOR U35306 ( .A(n35719), .B(n35764), .Z(n35766) );
  XNOR U35307 ( .A(n35787), .B(n35788), .Z(n35719) );
  AND U35308 ( .A(n645), .B(n35789), .Z(n35788) );
  XNOR U35309 ( .A(n35790), .B(n35791), .Z(n35789) );
  XOR U35310 ( .A(n35792), .B(n35793), .Z(n35764) );
  AND U35311 ( .A(n35794), .B(n35795), .Z(n35793) );
  XNOR U35312 ( .A(n35792), .B(n35780), .Z(n35795) );
  IV U35313 ( .A(n35730), .Z(n35780) );
  XNOR U35314 ( .A(n35796), .B(n35773), .Z(n35730) );
  XNOR U35315 ( .A(n35797), .B(n35779), .Z(n35773) );
  XOR U35316 ( .A(n35798), .B(n35799), .Z(n35779) );
  NOR U35317 ( .A(n35800), .B(n35801), .Z(n35799) );
  XNOR U35318 ( .A(n35798), .B(n35802), .Z(n35800) );
  XNOR U35319 ( .A(n35778), .B(n35770), .Z(n35797) );
  XOR U35320 ( .A(n35803), .B(n35804), .Z(n35770) );
  AND U35321 ( .A(n35805), .B(n35806), .Z(n35804) );
  XNOR U35322 ( .A(n35803), .B(n35807), .Z(n35805) );
  XNOR U35323 ( .A(n35808), .B(n35775), .Z(n35778) );
  XOR U35324 ( .A(n35809), .B(n35810), .Z(n35775) );
  AND U35325 ( .A(n35811), .B(n35812), .Z(n35810) );
  XOR U35326 ( .A(n35809), .B(n35813), .Z(n35811) );
  XNOR U35327 ( .A(n35814), .B(n35815), .Z(n35808) );
  NOR U35328 ( .A(n35816), .B(n35817), .Z(n35815) );
  XOR U35329 ( .A(n35814), .B(n35818), .Z(n35816) );
  XNOR U35330 ( .A(n35774), .B(n35781), .Z(n35796) );
  NOR U35331 ( .A(n35736), .B(n35819), .Z(n35781) );
  XOR U35332 ( .A(n35786), .B(n35785), .Z(n35774) );
  XNOR U35333 ( .A(n35820), .B(n35782), .Z(n35785) );
  XOR U35334 ( .A(n35821), .B(n35822), .Z(n35782) );
  AND U35335 ( .A(n35823), .B(n35824), .Z(n35822) );
  XOR U35336 ( .A(n35821), .B(n35825), .Z(n35823) );
  XNOR U35337 ( .A(n35826), .B(n35827), .Z(n35820) );
  NOR U35338 ( .A(n35828), .B(n35829), .Z(n35827) );
  XNOR U35339 ( .A(n35826), .B(n35830), .Z(n35828) );
  XOR U35340 ( .A(n35831), .B(n35832), .Z(n35786) );
  NOR U35341 ( .A(n35833), .B(n35834), .Z(n35832) );
  XNOR U35342 ( .A(n35831), .B(n35835), .Z(n35833) );
  XNOR U35343 ( .A(n35727), .B(n35792), .Z(n35794) );
  XNOR U35344 ( .A(n35836), .B(n35837), .Z(n35727) );
  AND U35345 ( .A(n645), .B(n35838), .Z(n35837) );
  XNOR U35346 ( .A(n35839), .B(n35840), .Z(n35838) );
  AND U35347 ( .A(n35733), .B(n35736), .Z(n35792) );
  XOR U35348 ( .A(n35841), .B(n35819), .Z(n35736) );
  XNOR U35349 ( .A(p_input[2048]), .B(p_input[480]), .Z(n35819) );
  XOR U35350 ( .A(n35807), .B(n35806), .Z(n35841) );
  XNOR U35351 ( .A(n35842), .B(n35813), .Z(n35806) );
  XNOR U35352 ( .A(n35802), .B(n35801), .Z(n35813) );
  XOR U35353 ( .A(n35843), .B(n35798), .Z(n35801) );
  XNOR U35354 ( .A(n29266), .B(p_input[490]), .Z(n35798) );
  XNOR U35355 ( .A(p_input[2059]), .B(p_input[491]), .Z(n35843) );
  XOR U35356 ( .A(p_input[2060]), .B(p_input[492]), .Z(n35802) );
  XNOR U35357 ( .A(n35812), .B(n35803), .Z(n35842) );
  XNOR U35358 ( .A(n29494), .B(p_input[481]), .Z(n35803) );
  XOR U35359 ( .A(n35844), .B(n35818), .Z(n35812) );
  XNOR U35360 ( .A(p_input[2063]), .B(p_input[495]), .Z(n35818) );
  XOR U35361 ( .A(n35809), .B(n35817), .Z(n35844) );
  XOR U35362 ( .A(n35845), .B(n35814), .Z(n35817) );
  XOR U35363 ( .A(p_input[2061]), .B(p_input[493]), .Z(n35814) );
  XNOR U35364 ( .A(p_input[2062]), .B(p_input[494]), .Z(n35845) );
  XNOR U35365 ( .A(n29036), .B(p_input[489]), .Z(n35809) );
  XNOR U35366 ( .A(n35825), .B(n35824), .Z(n35807) );
  XNOR U35367 ( .A(n35846), .B(n35830), .Z(n35824) );
  XOR U35368 ( .A(p_input[2056]), .B(p_input[488]), .Z(n35830) );
  XOR U35369 ( .A(n35821), .B(n35829), .Z(n35846) );
  XOR U35370 ( .A(n35847), .B(n35826), .Z(n35829) );
  XOR U35371 ( .A(p_input[2054]), .B(p_input[486]), .Z(n35826) );
  XNOR U35372 ( .A(p_input[2055]), .B(p_input[487]), .Z(n35847) );
  XNOR U35373 ( .A(n29039), .B(p_input[482]), .Z(n35821) );
  XNOR U35374 ( .A(n35835), .B(n35834), .Z(n35825) );
  XOR U35375 ( .A(n35848), .B(n35831), .Z(n35834) );
  XOR U35376 ( .A(p_input[2051]), .B(p_input[483]), .Z(n35831) );
  XNOR U35377 ( .A(p_input[2052]), .B(p_input[484]), .Z(n35848) );
  XOR U35378 ( .A(p_input[2053]), .B(p_input[485]), .Z(n35835) );
  XNOR U35379 ( .A(n35849), .B(n35850), .Z(n35733) );
  AND U35380 ( .A(n645), .B(n35851), .Z(n35850) );
  XNOR U35381 ( .A(n35852), .B(n35853), .Z(n645) );
  AND U35382 ( .A(n35854), .B(n35855), .Z(n35853) );
  XOR U35383 ( .A(n35747), .B(n35852), .Z(n35855) );
  XNOR U35384 ( .A(n35856), .B(n35852), .Z(n35854) );
  XOR U35385 ( .A(n35857), .B(n35858), .Z(n35852) );
  AND U35386 ( .A(n35859), .B(n35860), .Z(n35858) );
  XOR U35387 ( .A(n35762), .B(n35857), .Z(n35860) );
  XOR U35388 ( .A(n35857), .B(n35763), .Z(n35859) );
  XOR U35389 ( .A(n35861), .B(n35862), .Z(n35857) );
  AND U35390 ( .A(n35863), .B(n35864), .Z(n35862) );
  XOR U35391 ( .A(n35790), .B(n35861), .Z(n35864) );
  XOR U35392 ( .A(n35861), .B(n35791), .Z(n35863) );
  XOR U35393 ( .A(n35865), .B(n35866), .Z(n35861) );
  AND U35394 ( .A(n35867), .B(n35868), .Z(n35866) );
  XOR U35395 ( .A(n35865), .B(n35839), .Z(n35868) );
  XNOR U35396 ( .A(n35869), .B(n35870), .Z(n35693) );
  AND U35397 ( .A(n649), .B(n35871), .Z(n35870) );
  XNOR U35398 ( .A(n35872), .B(n35873), .Z(n649) );
  AND U35399 ( .A(n35874), .B(n35875), .Z(n35873) );
  XOR U35400 ( .A(n35872), .B(n35703), .Z(n35875) );
  XNOR U35401 ( .A(n35872), .B(n35663), .Z(n35874) );
  XOR U35402 ( .A(n35876), .B(n35877), .Z(n35872) );
  AND U35403 ( .A(n35878), .B(n35879), .Z(n35877) );
  XOR U35404 ( .A(n35876), .B(n35671), .Z(n35878) );
  XOR U35405 ( .A(n35880), .B(n35881), .Z(n35654) );
  AND U35406 ( .A(n653), .B(n35871), .Z(n35881) );
  XNOR U35407 ( .A(n35869), .B(n35880), .Z(n35871) );
  XNOR U35408 ( .A(n35882), .B(n35883), .Z(n653) );
  AND U35409 ( .A(n35884), .B(n35885), .Z(n35883) );
  XNOR U35410 ( .A(n35886), .B(n35882), .Z(n35885) );
  IV U35411 ( .A(n35703), .Z(n35886) );
  XOR U35412 ( .A(n35856), .B(n35887), .Z(n35703) );
  AND U35413 ( .A(n656), .B(n35888), .Z(n35887) );
  XOR U35414 ( .A(n35746), .B(n35743), .Z(n35888) );
  IV U35415 ( .A(n35856), .Z(n35746) );
  XNOR U35416 ( .A(n35663), .B(n35882), .Z(n35884) );
  XOR U35417 ( .A(n35889), .B(n35890), .Z(n35663) );
  AND U35418 ( .A(n672), .B(n35891), .Z(n35890) );
  XOR U35419 ( .A(n35876), .B(n35892), .Z(n35882) );
  AND U35420 ( .A(n35893), .B(n35879), .Z(n35892) );
  XNOR U35421 ( .A(n35713), .B(n35876), .Z(n35879) );
  XOR U35422 ( .A(n35763), .B(n35894), .Z(n35713) );
  AND U35423 ( .A(n656), .B(n35895), .Z(n35894) );
  XOR U35424 ( .A(n35759), .B(n35763), .Z(n35895) );
  XNOR U35425 ( .A(n35896), .B(n35876), .Z(n35893) );
  IV U35426 ( .A(n35671), .Z(n35896) );
  XOR U35427 ( .A(n35897), .B(n35898), .Z(n35671) );
  AND U35428 ( .A(n672), .B(n35899), .Z(n35898) );
  XOR U35429 ( .A(n35900), .B(n35901), .Z(n35876) );
  AND U35430 ( .A(n35902), .B(n35903), .Z(n35901) );
  XNOR U35431 ( .A(n35723), .B(n35900), .Z(n35903) );
  XOR U35432 ( .A(n35791), .B(n35904), .Z(n35723) );
  AND U35433 ( .A(n656), .B(n35905), .Z(n35904) );
  XOR U35434 ( .A(n35787), .B(n35791), .Z(n35905) );
  XOR U35435 ( .A(n35900), .B(n35680), .Z(n35902) );
  XOR U35436 ( .A(n35906), .B(n35907), .Z(n35680) );
  AND U35437 ( .A(n672), .B(n35908), .Z(n35907) );
  XOR U35438 ( .A(n35909), .B(n35910), .Z(n35900) );
  AND U35439 ( .A(n35911), .B(n35912), .Z(n35910) );
  XNOR U35440 ( .A(n35909), .B(n35731), .Z(n35912) );
  XOR U35441 ( .A(n35840), .B(n35913), .Z(n35731) );
  AND U35442 ( .A(n656), .B(n35914), .Z(n35913) );
  XOR U35443 ( .A(n35836), .B(n35840), .Z(n35914) );
  XNOR U35444 ( .A(n35915), .B(n35909), .Z(n35911) );
  IV U35445 ( .A(n35690), .Z(n35915) );
  XOR U35446 ( .A(n35916), .B(n35917), .Z(n35690) );
  AND U35447 ( .A(n672), .B(n35918), .Z(n35917) );
  AND U35448 ( .A(n35880), .B(n35869), .Z(n35909) );
  XNOR U35449 ( .A(n35919), .B(n35920), .Z(n35869) );
  AND U35450 ( .A(n656), .B(n35851), .Z(n35920) );
  XNOR U35451 ( .A(n35849), .B(n35919), .Z(n35851) );
  XNOR U35452 ( .A(n35921), .B(n35922), .Z(n656) );
  AND U35453 ( .A(n35923), .B(n35924), .Z(n35922) );
  XNOR U35454 ( .A(n35921), .B(n35743), .Z(n35924) );
  IV U35455 ( .A(n35747), .Z(n35743) );
  XOR U35456 ( .A(n35925), .B(n35926), .Z(n35747) );
  AND U35457 ( .A(n660), .B(n35927), .Z(n35926) );
  XOR U35458 ( .A(n35928), .B(n35925), .Z(n35927) );
  XNOR U35459 ( .A(n35921), .B(n35856), .Z(n35923) );
  XOR U35460 ( .A(n35929), .B(n35930), .Z(n35856) );
  AND U35461 ( .A(n668), .B(n35891), .Z(n35930) );
  XOR U35462 ( .A(n35889), .B(n35929), .Z(n35891) );
  XOR U35463 ( .A(n35931), .B(n35932), .Z(n35921) );
  AND U35464 ( .A(n35933), .B(n35934), .Z(n35932) );
  XNOR U35465 ( .A(n35931), .B(n35759), .Z(n35934) );
  IV U35466 ( .A(n35762), .Z(n35759) );
  XOR U35467 ( .A(n35935), .B(n35936), .Z(n35762) );
  AND U35468 ( .A(n660), .B(n35937), .Z(n35936) );
  XOR U35469 ( .A(n35938), .B(n35935), .Z(n35937) );
  XOR U35470 ( .A(n35763), .B(n35931), .Z(n35933) );
  XOR U35471 ( .A(n35939), .B(n35940), .Z(n35763) );
  AND U35472 ( .A(n668), .B(n35899), .Z(n35940) );
  XOR U35473 ( .A(n35939), .B(n35897), .Z(n35899) );
  XOR U35474 ( .A(n35941), .B(n35942), .Z(n35931) );
  AND U35475 ( .A(n35943), .B(n35944), .Z(n35942) );
  XNOR U35476 ( .A(n35941), .B(n35787), .Z(n35944) );
  IV U35477 ( .A(n35790), .Z(n35787) );
  XOR U35478 ( .A(n35945), .B(n35946), .Z(n35790) );
  AND U35479 ( .A(n660), .B(n35947), .Z(n35946) );
  XNOR U35480 ( .A(n35948), .B(n35945), .Z(n35947) );
  XOR U35481 ( .A(n35791), .B(n35941), .Z(n35943) );
  XOR U35482 ( .A(n35949), .B(n35950), .Z(n35791) );
  AND U35483 ( .A(n668), .B(n35908), .Z(n35950) );
  XOR U35484 ( .A(n35949), .B(n35906), .Z(n35908) );
  XOR U35485 ( .A(n35865), .B(n35951), .Z(n35941) );
  AND U35486 ( .A(n35867), .B(n35952), .Z(n35951) );
  XNOR U35487 ( .A(n35865), .B(n35836), .Z(n35952) );
  IV U35488 ( .A(n35839), .Z(n35836) );
  XOR U35489 ( .A(n35953), .B(n35954), .Z(n35839) );
  AND U35490 ( .A(n660), .B(n35955), .Z(n35954) );
  XOR U35491 ( .A(n35956), .B(n35953), .Z(n35955) );
  XOR U35492 ( .A(n35840), .B(n35865), .Z(n35867) );
  XOR U35493 ( .A(n35957), .B(n35958), .Z(n35840) );
  AND U35494 ( .A(n668), .B(n35918), .Z(n35958) );
  XOR U35495 ( .A(n35957), .B(n35916), .Z(n35918) );
  AND U35496 ( .A(n35919), .B(n35849), .Z(n35865) );
  XNOR U35497 ( .A(n35959), .B(n35960), .Z(n35849) );
  AND U35498 ( .A(n660), .B(n35961), .Z(n35960) );
  XNOR U35499 ( .A(n35962), .B(n35959), .Z(n35961) );
  XNOR U35500 ( .A(n35963), .B(n35964), .Z(n660) );
  AND U35501 ( .A(n35965), .B(n35966), .Z(n35964) );
  XOR U35502 ( .A(n35928), .B(n35963), .Z(n35966) );
  AND U35503 ( .A(n35967), .B(n35968), .Z(n35928) );
  XNOR U35504 ( .A(n35925), .B(n35963), .Z(n35965) );
  XNOR U35505 ( .A(n35969), .B(n35970), .Z(n35925) );
  AND U35506 ( .A(n664), .B(n35971), .Z(n35970) );
  XNOR U35507 ( .A(n35972), .B(n35973), .Z(n35971) );
  XOR U35508 ( .A(n35974), .B(n35975), .Z(n35963) );
  AND U35509 ( .A(n35976), .B(n35977), .Z(n35975) );
  XNOR U35510 ( .A(n35974), .B(n35967), .Z(n35977) );
  IV U35511 ( .A(n35938), .Z(n35967) );
  XOR U35512 ( .A(n35978), .B(n35979), .Z(n35938) );
  XOR U35513 ( .A(n35980), .B(n35968), .Z(n35979) );
  AND U35514 ( .A(n35948), .B(n35981), .Z(n35968) );
  AND U35515 ( .A(n35982), .B(n35983), .Z(n35980) );
  XOR U35516 ( .A(n35984), .B(n35978), .Z(n35982) );
  XNOR U35517 ( .A(n35935), .B(n35974), .Z(n35976) );
  XNOR U35518 ( .A(n35985), .B(n35986), .Z(n35935) );
  AND U35519 ( .A(n664), .B(n35987), .Z(n35986) );
  XNOR U35520 ( .A(n35988), .B(n35989), .Z(n35987) );
  XOR U35521 ( .A(n35990), .B(n35991), .Z(n35974) );
  AND U35522 ( .A(n35992), .B(n35993), .Z(n35991) );
  XNOR U35523 ( .A(n35990), .B(n35948), .Z(n35993) );
  XOR U35524 ( .A(n35994), .B(n35983), .Z(n35948) );
  XNOR U35525 ( .A(n35995), .B(n35978), .Z(n35983) );
  XOR U35526 ( .A(n35996), .B(n35997), .Z(n35978) );
  AND U35527 ( .A(n35998), .B(n35999), .Z(n35997) );
  XOR U35528 ( .A(n36000), .B(n35996), .Z(n35998) );
  XNOR U35529 ( .A(n36001), .B(n36002), .Z(n35995) );
  AND U35530 ( .A(n36003), .B(n36004), .Z(n36002) );
  XOR U35531 ( .A(n36001), .B(n36005), .Z(n36003) );
  XNOR U35532 ( .A(n35984), .B(n35981), .Z(n35994) );
  AND U35533 ( .A(n36006), .B(n36007), .Z(n35981) );
  XOR U35534 ( .A(n36008), .B(n36009), .Z(n35984) );
  AND U35535 ( .A(n36010), .B(n36011), .Z(n36009) );
  XOR U35536 ( .A(n36008), .B(n36012), .Z(n36010) );
  XNOR U35537 ( .A(n35945), .B(n35990), .Z(n35992) );
  XNOR U35538 ( .A(n36013), .B(n36014), .Z(n35945) );
  AND U35539 ( .A(n664), .B(n36015), .Z(n36014) );
  XNOR U35540 ( .A(n36016), .B(n36017), .Z(n36015) );
  XOR U35541 ( .A(n36018), .B(n36019), .Z(n35990) );
  AND U35542 ( .A(n36020), .B(n36021), .Z(n36019) );
  XNOR U35543 ( .A(n36018), .B(n36006), .Z(n36021) );
  IV U35544 ( .A(n35956), .Z(n36006) );
  XNOR U35545 ( .A(n36022), .B(n35999), .Z(n35956) );
  XNOR U35546 ( .A(n36023), .B(n36005), .Z(n35999) );
  XOR U35547 ( .A(n36024), .B(n36025), .Z(n36005) );
  NOR U35548 ( .A(n36026), .B(n36027), .Z(n36025) );
  XNOR U35549 ( .A(n36024), .B(n36028), .Z(n36026) );
  XNOR U35550 ( .A(n36004), .B(n35996), .Z(n36023) );
  XOR U35551 ( .A(n36029), .B(n36030), .Z(n35996) );
  AND U35552 ( .A(n36031), .B(n36032), .Z(n36030) );
  XNOR U35553 ( .A(n36029), .B(n36033), .Z(n36031) );
  XNOR U35554 ( .A(n36034), .B(n36001), .Z(n36004) );
  XOR U35555 ( .A(n36035), .B(n36036), .Z(n36001) );
  AND U35556 ( .A(n36037), .B(n36038), .Z(n36036) );
  XOR U35557 ( .A(n36035), .B(n36039), .Z(n36037) );
  XNOR U35558 ( .A(n36040), .B(n36041), .Z(n36034) );
  NOR U35559 ( .A(n36042), .B(n36043), .Z(n36041) );
  XOR U35560 ( .A(n36040), .B(n36044), .Z(n36042) );
  XNOR U35561 ( .A(n36000), .B(n36007), .Z(n36022) );
  NOR U35562 ( .A(n35962), .B(n36045), .Z(n36007) );
  XOR U35563 ( .A(n36012), .B(n36011), .Z(n36000) );
  XNOR U35564 ( .A(n36046), .B(n36008), .Z(n36011) );
  XOR U35565 ( .A(n36047), .B(n36048), .Z(n36008) );
  AND U35566 ( .A(n36049), .B(n36050), .Z(n36048) );
  XOR U35567 ( .A(n36047), .B(n36051), .Z(n36049) );
  XNOR U35568 ( .A(n36052), .B(n36053), .Z(n36046) );
  NOR U35569 ( .A(n36054), .B(n36055), .Z(n36053) );
  XNOR U35570 ( .A(n36052), .B(n36056), .Z(n36054) );
  XOR U35571 ( .A(n36057), .B(n36058), .Z(n36012) );
  NOR U35572 ( .A(n36059), .B(n36060), .Z(n36058) );
  XNOR U35573 ( .A(n36057), .B(n36061), .Z(n36059) );
  XNOR U35574 ( .A(n35953), .B(n36018), .Z(n36020) );
  XNOR U35575 ( .A(n36062), .B(n36063), .Z(n35953) );
  AND U35576 ( .A(n664), .B(n36064), .Z(n36063) );
  XNOR U35577 ( .A(n36065), .B(n36066), .Z(n36064) );
  AND U35578 ( .A(n35959), .B(n35962), .Z(n36018) );
  XOR U35579 ( .A(n36067), .B(n36045), .Z(n35962) );
  XNOR U35580 ( .A(p_input[2048]), .B(p_input[496]), .Z(n36045) );
  XOR U35581 ( .A(n36033), .B(n36032), .Z(n36067) );
  XNOR U35582 ( .A(n36068), .B(n36039), .Z(n36032) );
  XNOR U35583 ( .A(n36028), .B(n36027), .Z(n36039) );
  XOR U35584 ( .A(n36069), .B(n36024), .Z(n36027) );
  XNOR U35585 ( .A(n29266), .B(p_input[506]), .Z(n36024) );
  XNOR U35586 ( .A(p_input[2059]), .B(p_input[507]), .Z(n36069) );
  XOR U35587 ( .A(p_input[2060]), .B(p_input[508]), .Z(n36028) );
  XNOR U35588 ( .A(n36038), .B(n36029), .Z(n36068) );
  XNOR U35589 ( .A(n29494), .B(p_input[497]), .Z(n36029) );
  XOR U35590 ( .A(n36070), .B(n36044), .Z(n36038) );
  XNOR U35591 ( .A(p_input[2063]), .B(p_input[511]), .Z(n36044) );
  XOR U35592 ( .A(n36035), .B(n36043), .Z(n36070) );
  XOR U35593 ( .A(n36071), .B(n36040), .Z(n36043) );
  XOR U35594 ( .A(p_input[2061]), .B(p_input[509]), .Z(n36040) );
  XNOR U35595 ( .A(p_input[2062]), .B(p_input[510]), .Z(n36071) );
  XNOR U35596 ( .A(n29036), .B(p_input[505]), .Z(n36035) );
  XNOR U35597 ( .A(n36051), .B(n36050), .Z(n36033) );
  XNOR U35598 ( .A(n36072), .B(n36056), .Z(n36050) );
  XOR U35599 ( .A(p_input[2056]), .B(p_input[504]), .Z(n36056) );
  XOR U35600 ( .A(n36047), .B(n36055), .Z(n36072) );
  XOR U35601 ( .A(n36073), .B(n36052), .Z(n36055) );
  XOR U35602 ( .A(p_input[2054]), .B(p_input[502]), .Z(n36052) );
  XNOR U35603 ( .A(p_input[2055]), .B(p_input[503]), .Z(n36073) );
  XNOR U35604 ( .A(n29039), .B(p_input[498]), .Z(n36047) );
  XNOR U35605 ( .A(n36061), .B(n36060), .Z(n36051) );
  XOR U35606 ( .A(n36074), .B(n36057), .Z(n36060) );
  XOR U35607 ( .A(p_input[2051]), .B(p_input[499]), .Z(n36057) );
  XNOR U35608 ( .A(p_input[2052]), .B(p_input[500]), .Z(n36074) );
  XOR U35609 ( .A(p_input[2053]), .B(p_input[501]), .Z(n36061) );
  XNOR U35610 ( .A(n36075), .B(n36076), .Z(n35959) );
  AND U35611 ( .A(n664), .B(n36077), .Z(n36076) );
  XNOR U35612 ( .A(n36078), .B(n36079), .Z(n664) );
  AND U35613 ( .A(n36080), .B(n36081), .Z(n36079) );
  XOR U35614 ( .A(n35973), .B(n36078), .Z(n36081) );
  XNOR U35615 ( .A(n36082), .B(n36078), .Z(n36080) );
  XOR U35616 ( .A(n36083), .B(n36084), .Z(n36078) );
  AND U35617 ( .A(n36085), .B(n36086), .Z(n36084) );
  XOR U35618 ( .A(n35988), .B(n36083), .Z(n36086) );
  XOR U35619 ( .A(n36083), .B(n35989), .Z(n36085) );
  XOR U35620 ( .A(n36087), .B(n36088), .Z(n36083) );
  AND U35621 ( .A(n36089), .B(n36090), .Z(n36088) );
  XOR U35622 ( .A(n36016), .B(n36087), .Z(n36090) );
  XOR U35623 ( .A(n36087), .B(n36017), .Z(n36089) );
  XOR U35624 ( .A(n36091), .B(n36092), .Z(n36087) );
  AND U35625 ( .A(n36093), .B(n36094), .Z(n36092) );
  XOR U35626 ( .A(n36091), .B(n36065), .Z(n36094) );
  XNOR U35627 ( .A(n36095), .B(n36096), .Z(n35919) );
  AND U35628 ( .A(n668), .B(n36097), .Z(n36096) );
  XNOR U35629 ( .A(n36098), .B(n36099), .Z(n668) );
  AND U35630 ( .A(n36100), .B(n36101), .Z(n36099) );
  XOR U35631 ( .A(n36098), .B(n35929), .Z(n36101) );
  XNOR U35632 ( .A(n36098), .B(n35889), .Z(n36100) );
  XOR U35633 ( .A(n36102), .B(n36103), .Z(n36098) );
  AND U35634 ( .A(n36104), .B(n36105), .Z(n36103) );
  XOR U35635 ( .A(n36102), .B(n35897), .Z(n36104) );
  XOR U35636 ( .A(n36106), .B(n36107), .Z(n35880) );
  AND U35637 ( .A(n672), .B(n36097), .Z(n36107) );
  XNOR U35638 ( .A(n36095), .B(n36106), .Z(n36097) );
  XNOR U35639 ( .A(n36108), .B(n36109), .Z(n672) );
  AND U35640 ( .A(n36110), .B(n36111), .Z(n36109) );
  XNOR U35641 ( .A(n36112), .B(n36108), .Z(n36111) );
  IV U35642 ( .A(n35929), .Z(n36112) );
  XOR U35643 ( .A(n36082), .B(n36113), .Z(n35929) );
  AND U35644 ( .A(n675), .B(n36114), .Z(n36113) );
  XOR U35645 ( .A(n35972), .B(n35969), .Z(n36114) );
  IV U35646 ( .A(n36082), .Z(n35972) );
  XNOR U35647 ( .A(n35889), .B(n36108), .Z(n36110) );
  XOR U35648 ( .A(n36115), .B(n36116), .Z(n35889) );
  AND U35649 ( .A(n691), .B(n36117), .Z(n36116) );
  XOR U35650 ( .A(n36102), .B(n36118), .Z(n36108) );
  AND U35651 ( .A(n36119), .B(n36105), .Z(n36118) );
  XNOR U35652 ( .A(n35939), .B(n36102), .Z(n36105) );
  XOR U35653 ( .A(n35989), .B(n36120), .Z(n35939) );
  AND U35654 ( .A(n675), .B(n36121), .Z(n36120) );
  XOR U35655 ( .A(n35985), .B(n35989), .Z(n36121) );
  XNOR U35656 ( .A(n36122), .B(n36102), .Z(n36119) );
  IV U35657 ( .A(n35897), .Z(n36122) );
  XOR U35658 ( .A(n36123), .B(n36124), .Z(n35897) );
  AND U35659 ( .A(n691), .B(n36125), .Z(n36124) );
  XOR U35660 ( .A(n36126), .B(n36127), .Z(n36102) );
  AND U35661 ( .A(n36128), .B(n36129), .Z(n36127) );
  XNOR U35662 ( .A(n35949), .B(n36126), .Z(n36129) );
  XOR U35663 ( .A(n36017), .B(n36130), .Z(n35949) );
  AND U35664 ( .A(n675), .B(n36131), .Z(n36130) );
  XOR U35665 ( .A(n36013), .B(n36017), .Z(n36131) );
  XOR U35666 ( .A(n36126), .B(n35906), .Z(n36128) );
  XOR U35667 ( .A(n36132), .B(n36133), .Z(n35906) );
  AND U35668 ( .A(n691), .B(n36134), .Z(n36133) );
  XOR U35669 ( .A(n36135), .B(n36136), .Z(n36126) );
  AND U35670 ( .A(n36137), .B(n36138), .Z(n36136) );
  XNOR U35671 ( .A(n36135), .B(n35957), .Z(n36138) );
  XOR U35672 ( .A(n36066), .B(n36139), .Z(n35957) );
  AND U35673 ( .A(n675), .B(n36140), .Z(n36139) );
  XOR U35674 ( .A(n36062), .B(n36066), .Z(n36140) );
  XNOR U35675 ( .A(n36141), .B(n36135), .Z(n36137) );
  IV U35676 ( .A(n35916), .Z(n36141) );
  XOR U35677 ( .A(n36142), .B(n36143), .Z(n35916) );
  AND U35678 ( .A(n691), .B(n36144), .Z(n36143) );
  AND U35679 ( .A(n36106), .B(n36095), .Z(n36135) );
  XNOR U35680 ( .A(n36145), .B(n36146), .Z(n36095) );
  AND U35681 ( .A(n675), .B(n36077), .Z(n36146) );
  XNOR U35682 ( .A(n36075), .B(n36145), .Z(n36077) );
  XNOR U35683 ( .A(n36147), .B(n36148), .Z(n675) );
  AND U35684 ( .A(n36149), .B(n36150), .Z(n36148) );
  XNOR U35685 ( .A(n36147), .B(n35969), .Z(n36150) );
  IV U35686 ( .A(n35973), .Z(n35969) );
  XOR U35687 ( .A(n36151), .B(n36152), .Z(n35973) );
  AND U35688 ( .A(n679), .B(n36153), .Z(n36152) );
  XOR U35689 ( .A(n36154), .B(n36151), .Z(n36153) );
  XNOR U35690 ( .A(n36147), .B(n36082), .Z(n36149) );
  XOR U35691 ( .A(n36155), .B(n36156), .Z(n36082) );
  AND U35692 ( .A(n687), .B(n36117), .Z(n36156) );
  XOR U35693 ( .A(n36115), .B(n36155), .Z(n36117) );
  XOR U35694 ( .A(n36157), .B(n36158), .Z(n36147) );
  AND U35695 ( .A(n36159), .B(n36160), .Z(n36158) );
  XNOR U35696 ( .A(n36157), .B(n35985), .Z(n36160) );
  IV U35697 ( .A(n35988), .Z(n35985) );
  XOR U35698 ( .A(n36161), .B(n36162), .Z(n35988) );
  AND U35699 ( .A(n679), .B(n36163), .Z(n36162) );
  XOR U35700 ( .A(n36164), .B(n36161), .Z(n36163) );
  XOR U35701 ( .A(n35989), .B(n36157), .Z(n36159) );
  XOR U35702 ( .A(n36165), .B(n36166), .Z(n35989) );
  AND U35703 ( .A(n687), .B(n36125), .Z(n36166) );
  XOR U35704 ( .A(n36165), .B(n36123), .Z(n36125) );
  XOR U35705 ( .A(n36167), .B(n36168), .Z(n36157) );
  AND U35706 ( .A(n36169), .B(n36170), .Z(n36168) );
  XNOR U35707 ( .A(n36167), .B(n36013), .Z(n36170) );
  IV U35708 ( .A(n36016), .Z(n36013) );
  XOR U35709 ( .A(n36171), .B(n36172), .Z(n36016) );
  AND U35710 ( .A(n679), .B(n36173), .Z(n36172) );
  XNOR U35711 ( .A(n36174), .B(n36171), .Z(n36173) );
  XOR U35712 ( .A(n36017), .B(n36167), .Z(n36169) );
  XOR U35713 ( .A(n36175), .B(n36176), .Z(n36017) );
  AND U35714 ( .A(n687), .B(n36134), .Z(n36176) );
  XOR U35715 ( .A(n36175), .B(n36132), .Z(n36134) );
  XOR U35716 ( .A(n36091), .B(n36177), .Z(n36167) );
  AND U35717 ( .A(n36093), .B(n36178), .Z(n36177) );
  XNOR U35718 ( .A(n36091), .B(n36062), .Z(n36178) );
  IV U35719 ( .A(n36065), .Z(n36062) );
  XOR U35720 ( .A(n36179), .B(n36180), .Z(n36065) );
  AND U35721 ( .A(n679), .B(n36181), .Z(n36180) );
  XOR U35722 ( .A(n36182), .B(n36179), .Z(n36181) );
  XOR U35723 ( .A(n36066), .B(n36091), .Z(n36093) );
  XOR U35724 ( .A(n36183), .B(n36184), .Z(n36066) );
  AND U35725 ( .A(n687), .B(n36144), .Z(n36184) );
  XOR U35726 ( .A(n36183), .B(n36142), .Z(n36144) );
  AND U35727 ( .A(n36145), .B(n36075), .Z(n36091) );
  XNOR U35728 ( .A(n36185), .B(n36186), .Z(n36075) );
  AND U35729 ( .A(n679), .B(n36187), .Z(n36186) );
  XNOR U35730 ( .A(n36188), .B(n36185), .Z(n36187) );
  XNOR U35731 ( .A(n36189), .B(n36190), .Z(n679) );
  AND U35732 ( .A(n36191), .B(n36192), .Z(n36190) );
  XOR U35733 ( .A(n36154), .B(n36189), .Z(n36192) );
  AND U35734 ( .A(n36193), .B(n36194), .Z(n36154) );
  XNOR U35735 ( .A(n36151), .B(n36189), .Z(n36191) );
  XNOR U35736 ( .A(n36195), .B(n36196), .Z(n36151) );
  AND U35737 ( .A(n683), .B(n36197), .Z(n36196) );
  XNOR U35738 ( .A(n36198), .B(n36199), .Z(n36197) );
  XOR U35739 ( .A(n36200), .B(n36201), .Z(n36189) );
  AND U35740 ( .A(n36202), .B(n36203), .Z(n36201) );
  XNOR U35741 ( .A(n36200), .B(n36193), .Z(n36203) );
  IV U35742 ( .A(n36164), .Z(n36193) );
  XOR U35743 ( .A(n36204), .B(n36205), .Z(n36164) );
  XOR U35744 ( .A(n36206), .B(n36194), .Z(n36205) );
  AND U35745 ( .A(n36174), .B(n36207), .Z(n36194) );
  AND U35746 ( .A(n36208), .B(n36209), .Z(n36206) );
  XOR U35747 ( .A(n36210), .B(n36204), .Z(n36208) );
  XNOR U35748 ( .A(n36161), .B(n36200), .Z(n36202) );
  XNOR U35749 ( .A(n36211), .B(n36212), .Z(n36161) );
  AND U35750 ( .A(n683), .B(n36213), .Z(n36212) );
  XNOR U35751 ( .A(n36214), .B(n36215), .Z(n36213) );
  XOR U35752 ( .A(n36216), .B(n36217), .Z(n36200) );
  AND U35753 ( .A(n36218), .B(n36219), .Z(n36217) );
  XNOR U35754 ( .A(n36216), .B(n36174), .Z(n36219) );
  XOR U35755 ( .A(n36220), .B(n36209), .Z(n36174) );
  XNOR U35756 ( .A(n36221), .B(n36204), .Z(n36209) );
  XOR U35757 ( .A(n36222), .B(n36223), .Z(n36204) );
  AND U35758 ( .A(n36224), .B(n36225), .Z(n36223) );
  XOR U35759 ( .A(n36226), .B(n36222), .Z(n36224) );
  XNOR U35760 ( .A(n36227), .B(n36228), .Z(n36221) );
  AND U35761 ( .A(n36229), .B(n36230), .Z(n36228) );
  XOR U35762 ( .A(n36227), .B(n36231), .Z(n36229) );
  XNOR U35763 ( .A(n36210), .B(n36207), .Z(n36220) );
  AND U35764 ( .A(n36232), .B(n36233), .Z(n36207) );
  XOR U35765 ( .A(n36234), .B(n36235), .Z(n36210) );
  AND U35766 ( .A(n36236), .B(n36237), .Z(n36235) );
  XOR U35767 ( .A(n36234), .B(n36238), .Z(n36236) );
  XNOR U35768 ( .A(n36171), .B(n36216), .Z(n36218) );
  XNOR U35769 ( .A(n36239), .B(n36240), .Z(n36171) );
  AND U35770 ( .A(n683), .B(n36241), .Z(n36240) );
  XNOR U35771 ( .A(n36242), .B(n36243), .Z(n36241) );
  XOR U35772 ( .A(n36244), .B(n36245), .Z(n36216) );
  AND U35773 ( .A(n36246), .B(n36247), .Z(n36245) );
  XNOR U35774 ( .A(n36244), .B(n36232), .Z(n36247) );
  IV U35775 ( .A(n36182), .Z(n36232) );
  XNOR U35776 ( .A(n36248), .B(n36225), .Z(n36182) );
  XNOR U35777 ( .A(n36249), .B(n36231), .Z(n36225) );
  XOR U35778 ( .A(n36250), .B(n36251), .Z(n36231) );
  NOR U35779 ( .A(n36252), .B(n36253), .Z(n36251) );
  XNOR U35780 ( .A(n36250), .B(n36254), .Z(n36252) );
  XNOR U35781 ( .A(n36230), .B(n36222), .Z(n36249) );
  XOR U35782 ( .A(n36255), .B(n36256), .Z(n36222) );
  AND U35783 ( .A(n36257), .B(n36258), .Z(n36256) );
  XNOR U35784 ( .A(n36255), .B(n36259), .Z(n36257) );
  XNOR U35785 ( .A(n36260), .B(n36227), .Z(n36230) );
  XOR U35786 ( .A(n36261), .B(n36262), .Z(n36227) );
  AND U35787 ( .A(n36263), .B(n36264), .Z(n36262) );
  XOR U35788 ( .A(n36261), .B(n36265), .Z(n36263) );
  XNOR U35789 ( .A(n36266), .B(n36267), .Z(n36260) );
  NOR U35790 ( .A(n36268), .B(n36269), .Z(n36267) );
  XOR U35791 ( .A(n36266), .B(n36270), .Z(n36268) );
  XNOR U35792 ( .A(n36226), .B(n36233), .Z(n36248) );
  NOR U35793 ( .A(n36188), .B(n36271), .Z(n36233) );
  XOR U35794 ( .A(n36238), .B(n36237), .Z(n36226) );
  XNOR U35795 ( .A(n36272), .B(n36234), .Z(n36237) );
  XOR U35796 ( .A(n36273), .B(n36274), .Z(n36234) );
  AND U35797 ( .A(n36275), .B(n36276), .Z(n36274) );
  XOR U35798 ( .A(n36273), .B(n36277), .Z(n36275) );
  XNOR U35799 ( .A(n36278), .B(n36279), .Z(n36272) );
  NOR U35800 ( .A(n36280), .B(n36281), .Z(n36279) );
  XNOR U35801 ( .A(n36278), .B(n36282), .Z(n36280) );
  XOR U35802 ( .A(n36283), .B(n36284), .Z(n36238) );
  NOR U35803 ( .A(n36285), .B(n36286), .Z(n36284) );
  XNOR U35804 ( .A(n36283), .B(n36287), .Z(n36285) );
  XNOR U35805 ( .A(n36179), .B(n36244), .Z(n36246) );
  XNOR U35806 ( .A(n36288), .B(n36289), .Z(n36179) );
  AND U35807 ( .A(n683), .B(n36290), .Z(n36289) );
  XNOR U35808 ( .A(n36291), .B(n36292), .Z(n36290) );
  AND U35809 ( .A(n36185), .B(n36188), .Z(n36244) );
  XOR U35810 ( .A(n36293), .B(n36271), .Z(n36188) );
  XNOR U35811 ( .A(p_input[2048]), .B(p_input[512]), .Z(n36271) );
  XOR U35812 ( .A(n36259), .B(n36258), .Z(n36293) );
  XNOR U35813 ( .A(n36294), .B(n36265), .Z(n36258) );
  XNOR U35814 ( .A(n36254), .B(n36253), .Z(n36265) );
  XOR U35815 ( .A(n36295), .B(n36250), .Z(n36253) );
  XNOR U35816 ( .A(n29266), .B(p_input[522]), .Z(n36250) );
  XNOR U35817 ( .A(p_input[2059]), .B(p_input[523]), .Z(n36295) );
  XOR U35818 ( .A(p_input[2060]), .B(p_input[524]), .Z(n36254) );
  XNOR U35819 ( .A(n36264), .B(n36255), .Z(n36294) );
  XNOR U35820 ( .A(n29494), .B(p_input[513]), .Z(n36255) );
  XOR U35821 ( .A(n36296), .B(n36270), .Z(n36264) );
  XNOR U35822 ( .A(p_input[2063]), .B(p_input[527]), .Z(n36270) );
  XOR U35823 ( .A(n36261), .B(n36269), .Z(n36296) );
  XOR U35824 ( .A(n36297), .B(n36266), .Z(n36269) );
  XOR U35825 ( .A(p_input[2061]), .B(p_input[525]), .Z(n36266) );
  XNOR U35826 ( .A(p_input[2062]), .B(p_input[526]), .Z(n36297) );
  XNOR U35827 ( .A(n29036), .B(p_input[521]), .Z(n36261) );
  XNOR U35828 ( .A(n36277), .B(n36276), .Z(n36259) );
  XNOR U35829 ( .A(n36298), .B(n36282), .Z(n36276) );
  XOR U35830 ( .A(p_input[2056]), .B(p_input[520]), .Z(n36282) );
  XOR U35831 ( .A(n36273), .B(n36281), .Z(n36298) );
  XOR U35832 ( .A(n36299), .B(n36278), .Z(n36281) );
  XOR U35833 ( .A(p_input[2054]), .B(p_input[518]), .Z(n36278) );
  XNOR U35834 ( .A(p_input[2055]), .B(p_input[519]), .Z(n36299) );
  XNOR U35835 ( .A(n29039), .B(p_input[514]), .Z(n36273) );
  XNOR U35836 ( .A(n36287), .B(n36286), .Z(n36277) );
  XOR U35837 ( .A(n36300), .B(n36283), .Z(n36286) );
  XOR U35838 ( .A(p_input[2051]), .B(p_input[515]), .Z(n36283) );
  XNOR U35839 ( .A(p_input[2052]), .B(p_input[516]), .Z(n36300) );
  XOR U35840 ( .A(p_input[2053]), .B(p_input[517]), .Z(n36287) );
  XNOR U35841 ( .A(n36301), .B(n36302), .Z(n36185) );
  AND U35842 ( .A(n683), .B(n36303), .Z(n36302) );
  XNOR U35843 ( .A(n36304), .B(n36305), .Z(n683) );
  AND U35844 ( .A(n36306), .B(n36307), .Z(n36305) );
  XOR U35845 ( .A(n36199), .B(n36304), .Z(n36307) );
  XNOR U35846 ( .A(n36308), .B(n36304), .Z(n36306) );
  XOR U35847 ( .A(n36309), .B(n36310), .Z(n36304) );
  AND U35848 ( .A(n36311), .B(n36312), .Z(n36310) );
  XOR U35849 ( .A(n36214), .B(n36309), .Z(n36312) );
  XOR U35850 ( .A(n36309), .B(n36215), .Z(n36311) );
  XOR U35851 ( .A(n36313), .B(n36314), .Z(n36309) );
  AND U35852 ( .A(n36315), .B(n36316), .Z(n36314) );
  XOR U35853 ( .A(n36242), .B(n36313), .Z(n36316) );
  XOR U35854 ( .A(n36313), .B(n36243), .Z(n36315) );
  XOR U35855 ( .A(n36317), .B(n36318), .Z(n36313) );
  AND U35856 ( .A(n36319), .B(n36320), .Z(n36318) );
  XOR U35857 ( .A(n36317), .B(n36291), .Z(n36320) );
  XNOR U35858 ( .A(n36321), .B(n36322), .Z(n36145) );
  AND U35859 ( .A(n687), .B(n36323), .Z(n36322) );
  XNOR U35860 ( .A(n36324), .B(n36325), .Z(n687) );
  AND U35861 ( .A(n36326), .B(n36327), .Z(n36325) );
  XOR U35862 ( .A(n36324), .B(n36155), .Z(n36327) );
  XNOR U35863 ( .A(n36324), .B(n36115), .Z(n36326) );
  XOR U35864 ( .A(n36328), .B(n36329), .Z(n36324) );
  AND U35865 ( .A(n36330), .B(n36331), .Z(n36329) );
  XOR U35866 ( .A(n36328), .B(n36123), .Z(n36330) );
  XOR U35867 ( .A(n36332), .B(n36333), .Z(n36106) );
  AND U35868 ( .A(n691), .B(n36323), .Z(n36333) );
  XNOR U35869 ( .A(n36321), .B(n36332), .Z(n36323) );
  XNOR U35870 ( .A(n36334), .B(n36335), .Z(n691) );
  AND U35871 ( .A(n36336), .B(n36337), .Z(n36335) );
  XNOR U35872 ( .A(n36338), .B(n36334), .Z(n36337) );
  IV U35873 ( .A(n36155), .Z(n36338) );
  XOR U35874 ( .A(n36308), .B(n36339), .Z(n36155) );
  AND U35875 ( .A(n694), .B(n36340), .Z(n36339) );
  XOR U35876 ( .A(n36198), .B(n36195), .Z(n36340) );
  IV U35877 ( .A(n36308), .Z(n36198) );
  XNOR U35878 ( .A(n36115), .B(n36334), .Z(n36336) );
  XOR U35879 ( .A(n36341), .B(n36342), .Z(n36115) );
  AND U35880 ( .A(n710), .B(n36343), .Z(n36342) );
  XOR U35881 ( .A(n36328), .B(n36344), .Z(n36334) );
  AND U35882 ( .A(n36345), .B(n36331), .Z(n36344) );
  XNOR U35883 ( .A(n36165), .B(n36328), .Z(n36331) );
  XOR U35884 ( .A(n36215), .B(n36346), .Z(n36165) );
  AND U35885 ( .A(n694), .B(n36347), .Z(n36346) );
  XOR U35886 ( .A(n36211), .B(n36215), .Z(n36347) );
  XNOR U35887 ( .A(n36348), .B(n36328), .Z(n36345) );
  IV U35888 ( .A(n36123), .Z(n36348) );
  XOR U35889 ( .A(n36349), .B(n36350), .Z(n36123) );
  AND U35890 ( .A(n710), .B(n36351), .Z(n36350) );
  XOR U35891 ( .A(n36352), .B(n36353), .Z(n36328) );
  AND U35892 ( .A(n36354), .B(n36355), .Z(n36353) );
  XNOR U35893 ( .A(n36175), .B(n36352), .Z(n36355) );
  XOR U35894 ( .A(n36243), .B(n36356), .Z(n36175) );
  AND U35895 ( .A(n694), .B(n36357), .Z(n36356) );
  XOR U35896 ( .A(n36239), .B(n36243), .Z(n36357) );
  XOR U35897 ( .A(n36352), .B(n36132), .Z(n36354) );
  XOR U35898 ( .A(n36358), .B(n36359), .Z(n36132) );
  AND U35899 ( .A(n710), .B(n36360), .Z(n36359) );
  XOR U35900 ( .A(n36361), .B(n36362), .Z(n36352) );
  AND U35901 ( .A(n36363), .B(n36364), .Z(n36362) );
  XNOR U35902 ( .A(n36361), .B(n36183), .Z(n36364) );
  XOR U35903 ( .A(n36292), .B(n36365), .Z(n36183) );
  AND U35904 ( .A(n694), .B(n36366), .Z(n36365) );
  XOR U35905 ( .A(n36288), .B(n36292), .Z(n36366) );
  XNOR U35906 ( .A(n36367), .B(n36361), .Z(n36363) );
  IV U35907 ( .A(n36142), .Z(n36367) );
  XOR U35908 ( .A(n36368), .B(n36369), .Z(n36142) );
  AND U35909 ( .A(n710), .B(n36370), .Z(n36369) );
  AND U35910 ( .A(n36332), .B(n36321), .Z(n36361) );
  XNOR U35911 ( .A(n36371), .B(n36372), .Z(n36321) );
  AND U35912 ( .A(n694), .B(n36303), .Z(n36372) );
  XNOR U35913 ( .A(n36301), .B(n36371), .Z(n36303) );
  XNOR U35914 ( .A(n36373), .B(n36374), .Z(n694) );
  AND U35915 ( .A(n36375), .B(n36376), .Z(n36374) );
  XNOR U35916 ( .A(n36373), .B(n36195), .Z(n36376) );
  IV U35917 ( .A(n36199), .Z(n36195) );
  XOR U35918 ( .A(n36377), .B(n36378), .Z(n36199) );
  AND U35919 ( .A(n698), .B(n36379), .Z(n36378) );
  XOR U35920 ( .A(n36380), .B(n36377), .Z(n36379) );
  XNOR U35921 ( .A(n36373), .B(n36308), .Z(n36375) );
  XOR U35922 ( .A(n36381), .B(n36382), .Z(n36308) );
  AND U35923 ( .A(n706), .B(n36343), .Z(n36382) );
  XOR U35924 ( .A(n36341), .B(n36381), .Z(n36343) );
  XOR U35925 ( .A(n36383), .B(n36384), .Z(n36373) );
  AND U35926 ( .A(n36385), .B(n36386), .Z(n36384) );
  XNOR U35927 ( .A(n36383), .B(n36211), .Z(n36386) );
  IV U35928 ( .A(n36214), .Z(n36211) );
  XOR U35929 ( .A(n36387), .B(n36388), .Z(n36214) );
  AND U35930 ( .A(n698), .B(n36389), .Z(n36388) );
  XOR U35931 ( .A(n36390), .B(n36387), .Z(n36389) );
  XOR U35932 ( .A(n36215), .B(n36383), .Z(n36385) );
  XOR U35933 ( .A(n36391), .B(n36392), .Z(n36215) );
  AND U35934 ( .A(n706), .B(n36351), .Z(n36392) );
  XOR U35935 ( .A(n36391), .B(n36349), .Z(n36351) );
  XOR U35936 ( .A(n36393), .B(n36394), .Z(n36383) );
  AND U35937 ( .A(n36395), .B(n36396), .Z(n36394) );
  XNOR U35938 ( .A(n36393), .B(n36239), .Z(n36396) );
  IV U35939 ( .A(n36242), .Z(n36239) );
  XOR U35940 ( .A(n36397), .B(n36398), .Z(n36242) );
  AND U35941 ( .A(n698), .B(n36399), .Z(n36398) );
  XNOR U35942 ( .A(n36400), .B(n36397), .Z(n36399) );
  XOR U35943 ( .A(n36243), .B(n36393), .Z(n36395) );
  XOR U35944 ( .A(n36401), .B(n36402), .Z(n36243) );
  AND U35945 ( .A(n706), .B(n36360), .Z(n36402) );
  XOR U35946 ( .A(n36401), .B(n36358), .Z(n36360) );
  XOR U35947 ( .A(n36317), .B(n36403), .Z(n36393) );
  AND U35948 ( .A(n36319), .B(n36404), .Z(n36403) );
  XNOR U35949 ( .A(n36317), .B(n36288), .Z(n36404) );
  IV U35950 ( .A(n36291), .Z(n36288) );
  XOR U35951 ( .A(n36405), .B(n36406), .Z(n36291) );
  AND U35952 ( .A(n698), .B(n36407), .Z(n36406) );
  XOR U35953 ( .A(n36408), .B(n36405), .Z(n36407) );
  XOR U35954 ( .A(n36292), .B(n36317), .Z(n36319) );
  XOR U35955 ( .A(n36409), .B(n36410), .Z(n36292) );
  AND U35956 ( .A(n706), .B(n36370), .Z(n36410) );
  XOR U35957 ( .A(n36409), .B(n36368), .Z(n36370) );
  AND U35958 ( .A(n36371), .B(n36301), .Z(n36317) );
  XNOR U35959 ( .A(n36411), .B(n36412), .Z(n36301) );
  AND U35960 ( .A(n698), .B(n36413), .Z(n36412) );
  XNOR U35961 ( .A(n36414), .B(n36411), .Z(n36413) );
  XNOR U35962 ( .A(n36415), .B(n36416), .Z(n698) );
  AND U35963 ( .A(n36417), .B(n36418), .Z(n36416) );
  XOR U35964 ( .A(n36380), .B(n36415), .Z(n36418) );
  AND U35965 ( .A(n36419), .B(n36420), .Z(n36380) );
  XNOR U35966 ( .A(n36377), .B(n36415), .Z(n36417) );
  XNOR U35967 ( .A(n36421), .B(n36422), .Z(n36377) );
  AND U35968 ( .A(n702), .B(n36423), .Z(n36422) );
  XNOR U35969 ( .A(n36424), .B(n36425), .Z(n36423) );
  XOR U35970 ( .A(n36426), .B(n36427), .Z(n36415) );
  AND U35971 ( .A(n36428), .B(n36429), .Z(n36427) );
  XNOR U35972 ( .A(n36426), .B(n36419), .Z(n36429) );
  IV U35973 ( .A(n36390), .Z(n36419) );
  XOR U35974 ( .A(n36430), .B(n36431), .Z(n36390) );
  XOR U35975 ( .A(n36432), .B(n36420), .Z(n36431) );
  AND U35976 ( .A(n36400), .B(n36433), .Z(n36420) );
  AND U35977 ( .A(n36434), .B(n36435), .Z(n36432) );
  XOR U35978 ( .A(n36436), .B(n36430), .Z(n36434) );
  XNOR U35979 ( .A(n36387), .B(n36426), .Z(n36428) );
  XNOR U35980 ( .A(n36437), .B(n36438), .Z(n36387) );
  AND U35981 ( .A(n702), .B(n36439), .Z(n36438) );
  XNOR U35982 ( .A(n36440), .B(n36441), .Z(n36439) );
  XOR U35983 ( .A(n36442), .B(n36443), .Z(n36426) );
  AND U35984 ( .A(n36444), .B(n36445), .Z(n36443) );
  XNOR U35985 ( .A(n36442), .B(n36400), .Z(n36445) );
  XOR U35986 ( .A(n36446), .B(n36435), .Z(n36400) );
  XNOR U35987 ( .A(n36447), .B(n36430), .Z(n36435) );
  XOR U35988 ( .A(n36448), .B(n36449), .Z(n36430) );
  AND U35989 ( .A(n36450), .B(n36451), .Z(n36449) );
  XOR U35990 ( .A(n36452), .B(n36448), .Z(n36450) );
  XNOR U35991 ( .A(n36453), .B(n36454), .Z(n36447) );
  AND U35992 ( .A(n36455), .B(n36456), .Z(n36454) );
  XOR U35993 ( .A(n36453), .B(n36457), .Z(n36455) );
  XNOR U35994 ( .A(n36436), .B(n36433), .Z(n36446) );
  AND U35995 ( .A(n36458), .B(n36459), .Z(n36433) );
  XOR U35996 ( .A(n36460), .B(n36461), .Z(n36436) );
  AND U35997 ( .A(n36462), .B(n36463), .Z(n36461) );
  XOR U35998 ( .A(n36460), .B(n36464), .Z(n36462) );
  XNOR U35999 ( .A(n36397), .B(n36442), .Z(n36444) );
  XNOR U36000 ( .A(n36465), .B(n36466), .Z(n36397) );
  AND U36001 ( .A(n702), .B(n36467), .Z(n36466) );
  XNOR U36002 ( .A(n36468), .B(n36469), .Z(n36467) );
  XOR U36003 ( .A(n36470), .B(n36471), .Z(n36442) );
  AND U36004 ( .A(n36472), .B(n36473), .Z(n36471) );
  XNOR U36005 ( .A(n36470), .B(n36458), .Z(n36473) );
  IV U36006 ( .A(n36408), .Z(n36458) );
  XNOR U36007 ( .A(n36474), .B(n36451), .Z(n36408) );
  XNOR U36008 ( .A(n36475), .B(n36457), .Z(n36451) );
  XOR U36009 ( .A(n36476), .B(n36477), .Z(n36457) );
  NOR U36010 ( .A(n36478), .B(n36479), .Z(n36477) );
  XNOR U36011 ( .A(n36476), .B(n36480), .Z(n36478) );
  XNOR U36012 ( .A(n36456), .B(n36448), .Z(n36475) );
  XOR U36013 ( .A(n36481), .B(n36482), .Z(n36448) );
  AND U36014 ( .A(n36483), .B(n36484), .Z(n36482) );
  XNOR U36015 ( .A(n36481), .B(n36485), .Z(n36483) );
  XNOR U36016 ( .A(n36486), .B(n36453), .Z(n36456) );
  XOR U36017 ( .A(n36487), .B(n36488), .Z(n36453) );
  AND U36018 ( .A(n36489), .B(n36490), .Z(n36488) );
  XOR U36019 ( .A(n36487), .B(n36491), .Z(n36489) );
  XNOR U36020 ( .A(n36492), .B(n36493), .Z(n36486) );
  NOR U36021 ( .A(n36494), .B(n36495), .Z(n36493) );
  XOR U36022 ( .A(n36492), .B(n36496), .Z(n36494) );
  XNOR U36023 ( .A(n36452), .B(n36459), .Z(n36474) );
  NOR U36024 ( .A(n36414), .B(n36497), .Z(n36459) );
  XOR U36025 ( .A(n36464), .B(n36463), .Z(n36452) );
  XNOR U36026 ( .A(n36498), .B(n36460), .Z(n36463) );
  XOR U36027 ( .A(n36499), .B(n36500), .Z(n36460) );
  AND U36028 ( .A(n36501), .B(n36502), .Z(n36500) );
  XOR U36029 ( .A(n36499), .B(n36503), .Z(n36501) );
  XNOR U36030 ( .A(n36504), .B(n36505), .Z(n36498) );
  NOR U36031 ( .A(n36506), .B(n36507), .Z(n36505) );
  XNOR U36032 ( .A(n36504), .B(n36508), .Z(n36506) );
  XOR U36033 ( .A(n36509), .B(n36510), .Z(n36464) );
  NOR U36034 ( .A(n36511), .B(n36512), .Z(n36510) );
  XNOR U36035 ( .A(n36509), .B(n36513), .Z(n36511) );
  XNOR U36036 ( .A(n36405), .B(n36470), .Z(n36472) );
  XNOR U36037 ( .A(n36514), .B(n36515), .Z(n36405) );
  AND U36038 ( .A(n702), .B(n36516), .Z(n36515) );
  XNOR U36039 ( .A(n36517), .B(n36518), .Z(n36516) );
  AND U36040 ( .A(n36411), .B(n36414), .Z(n36470) );
  XOR U36041 ( .A(n36519), .B(n36497), .Z(n36414) );
  XNOR U36042 ( .A(p_input[2048]), .B(p_input[528]), .Z(n36497) );
  XOR U36043 ( .A(n36485), .B(n36484), .Z(n36519) );
  XNOR U36044 ( .A(n36520), .B(n36491), .Z(n36484) );
  XNOR U36045 ( .A(n36480), .B(n36479), .Z(n36491) );
  XOR U36046 ( .A(n36521), .B(n36476), .Z(n36479) );
  XNOR U36047 ( .A(n29266), .B(p_input[538]), .Z(n36476) );
  XNOR U36048 ( .A(p_input[2059]), .B(p_input[539]), .Z(n36521) );
  XOR U36049 ( .A(p_input[2060]), .B(p_input[540]), .Z(n36480) );
  XNOR U36050 ( .A(n36490), .B(n36481), .Z(n36520) );
  XNOR U36051 ( .A(n29494), .B(p_input[529]), .Z(n36481) );
  XOR U36052 ( .A(n36522), .B(n36496), .Z(n36490) );
  XNOR U36053 ( .A(p_input[2063]), .B(p_input[543]), .Z(n36496) );
  XOR U36054 ( .A(n36487), .B(n36495), .Z(n36522) );
  XOR U36055 ( .A(n36523), .B(n36492), .Z(n36495) );
  XOR U36056 ( .A(p_input[2061]), .B(p_input[541]), .Z(n36492) );
  XNOR U36057 ( .A(p_input[2062]), .B(p_input[542]), .Z(n36523) );
  XNOR U36058 ( .A(n29036), .B(p_input[537]), .Z(n36487) );
  XNOR U36059 ( .A(n36503), .B(n36502), .Z(n36485) );
  XNOR U36060 ( .A(n36524), .B(n36508), .Z(n36502) );
  XOR U36061 ( .A(p_input[2056]), .B(p_input[536]), .Z(n36508) );
  XOR U36062 ( .A(n36499), .B(n36507), .Z(n36524) );
  XOR U36063 ( .A(n36525), .B(n36504), .Z(n36507) );
  XOR U36064 ( .A(p_input[2054]), .B(p_input[534]), .Z(n36504) );
  XNOR U36065 ( .A(p_input[2055]), .B(p_input[535]), .Z(n36525) );
  XNOR U36066 ( .A(n29039), .B(p_input[530]), .Z(n36499) );
  XNOR U36067 ( .A(n36513), .B(n36512), .Z(n36503) );
  XOR U36068 ( .A(n36526), .B(n36509), .Z(n36512) );
  XOR U36069 ( .A(p_input[2051]), .B(p_input[531]), .Z(n36509) );
  XNOR U36070 ( .A(p_input[2052]), .B(p_input[532]), .Z(n36526) );
  XOR U36071 ( .A(p_input[2053]), .B(p_input[533]), .Z(n36513) );
  XNOR U36072 ( .A(n36527), .B(n36528), .Z(n36411) );
  AND U36073 ( .A(n702), .B(n36529), .Z(n36528) );
  XNOR U36074 ( .A(n36530), .B(n36531), .Z(n702) );
  AND U36075 ( .A(n36532), .B(n36533), .Z(n36531) );
  XOR U36076 ( .A(n36425), .B(n36530), .Z(n36533) );
  XNOR U36077 ( .A(n36534), .B(n36530), .Z(n36532) );
  XOR U36078 ( .A(n36535), .B(n36536), .Z(n36530) );
  AND U36079 ( .A(n36537), .B(n36538), .Z(n36536) );
  XOR U36080 ( .A(n36440), .B(n36535), .Z(n36538) );
  XOR U36081 ( .A(n36535), .B(n36441), .Z(n36537) );
  XOR U36082 ( .A(n36539), .B(n36540), .Z(n36535) );
  AND U36083 ( .A(n36541), .B(n36542), .Z(n36540) );
  XOR U36084 ( .A(n36468), .B(n36539), .Z(n36542) );
  XOR U36085 ( .A(n36539), .B(n36469), .Z(n36541) );
  XOR U36086 ( .A(n36543), .B(n36544), .Z(n36539) );
  AND U36087 ( .A(n36545), .B(n36546), .Z(n36544) );
  XOR U36088 ( .A(n36543), .B(n36517), .Z(n36546) );
  XNOR U36089 ( .A(n36547), .B(n36548), .Z(n36371) );
  AND U36090 ( .A(n706), .B(n36549), .Z(n36548) );
  XNOR U36091 ( .A(n36550), .B(n36551), .Z(n706) );
  AND U36092 ( .A(n36552), .B(n36553), .Z(n36551) );
  XOR U36093 ( .A(n36550), .B(n36381), .Z(n36553) );
  XNOR U36094 ( .A(n36550), .B(n36341), .Z(n36552) );
  XOR U36095 ( .A(n36554), .B(n36555), .Z(n36550) );
  AND U36096 ( .A(n36556), .B(n36557), .Z(n36555) );
  XOR U36097 ( .A(n36554), .B(n36349), .Z(n36556) );
  XOR U36098 ( .A(n36558), .B(n36559), .Z(n36332) );
  AND U36099 ( .A(n710), .B(n36549), .Z(n36559) );
  XNOR U36100 ( .A(n36547), .B(n36558), .Z(n36549) );
  XNOR U36101 ( .A(n36560), .B(n36561), .Z(n710) );
  AND U36102 ( .A(n36562), .B(n36563), .Z(n36561) );
  XNOR U36103 ( .A(n36564), .B(n36560), .Z(n36563) );
  IV U36104 ( .A(n36381), .Z(n36564) );
  XOR U36105 ( .A(n36534), .B(n36565), .Z(n36381) );
  AND U36106 ( .A(n713), .B(n36566), .Z(n36565) );
  XOR U36107 ( .A(n36424), .B(n36421), .Z(n36566) );
  IV U36108 ( .A(n36534), .Z(n36424) );
  XNOR U36109 ( .A(n36341), .B(n36560), .Z(n36562) );
  XOR U36110 ( .A(n36567), .B(n36568), .Z(n36341) );
  AND U36111 ( .A(n729), .B(n36569), .Z(n36568) );
  XOR U36112 ( .A(n36554), .B(n36570), .Z(n36560) );
  AND U36113 ( .A(n36571), .B(n36557), .Z(n36570) );
  XNOR U36114 ( .A(n36391), .B(n36554), .Z(n36557) );
  XOR U36115 ( .A(n36441), .B(n36572), .Z(n36391) );
  AND U36116 ( .A(n713), .B(n36573), .Z(n36572) );
  XOR U36117 ( .A(n36437), .B(n36441), .Z(n36573) );
  XNOR U36118 ( .A(n36574), .B(n36554), .Z(n36571) );
  IV U36119 ( .A(n36349), .Z(n36574) );
  XOR U36120 ( .A(n36575), .B(n36576), .Z(n36349) );
  AND U36121 ( .A(n729), .B(n36577), .Z(n36576) );
  XOR U36122 ( .A(n36578), .B(n36579), .Z(n36554) );
  AND U36123 ( .A(n36580), .B(n36581), .Z(n36579) );
  XNOR U36124 ( .A(n36401), .B(n36578), .Z(n36581) );
  XOR U36125 ( .A(n36469), .B(n36582), .Z(n36401) );
  AND U36126 ( .A(n713), .B(n36583), .Z(n36582) );
  XOR U36127 ( .A(n36465), .B(n36469), .Z(n36583) );
  XOR U36128 ( .A(n36578), .B(n36358), .Z(n36580) );
  XOR U36129 ( .A(n36584), .B(n36585), .Z(n36358) );
  AND U36130 ( .A(n729), .B(n36586), .Z(n36585) );
  XOR U36131 ( .A(n36587), .B(n36588), .Z(n36578) );
  AND U36132 ( .A(n36589), .B(n36590), .Z(n36588) );
  XNOR U36133 ( .A(n36587), .B(n36409), .Z(n36590) );
  XOR U36134 ( .A(n36518), .B(n36591), .Z(n36409) );
  AND U36135 ( .A(n713), .B(n36592), .Z(n36591) );
  XOR U36136 ( .A(n36514), .B(n36518), .Z(n36592) );
  XNOR U36137 ( .A(n36593), .B(n36587), .Z(n36589) );
  IV U36138 ( .A(n36368), .Z(n36593) );
  XOR U36139 ( .A(n36594), .B(n36595), .Z(n36368) );
  AND U36140 ( .A(n729), .B(n36596), .Z(n36595) );
  AND U36141 ( .A(n36558), .B(n36547), .Z(n36587) );
  XNOR U36142 ( .A(n36597), .B(n36598), .Z(n36547) );
  AND U36143 ( .A(n713), .B(n36529), .Z(n36598) );
  XNOR U36144 ( .A(n36527), .B(n36597), .Z(n36529) );
  XNOR U36145 ( .A(n36599), .B(n36600), .Z(n713) );
  AND U36146 ( .A(n36601), .B(n36602), .Z(n36600) );
  XNOR U36147 ( .A(n36599), .B(n36421), .Z(n36602) );
  IV U36148 ( .A(n36425), .Z(n36421) );
  XOR U36149 ( .A(n36603), .B(n36604), .Z(n36425) );
  AND U36150 ( .A(n717), .B(n36605), .Z(n36604) );
  XOR U36151 ( .A(n36606), .B(n36603), .Z(n36605) );
  XNOR U36152 ( .A(n36599), .B(n36534), .Z(n36601) );
  XOR U36153 ( .A(n36607), .B(n36608), .Z(n36534) );
  AND U36154 ( .A(n725), .B(n36569), .Z(n36608) );
  XOR U36155 ( .A(n36567), .B(n36607), .Z(n36569) );
  XOR U36156 ( .A(n36609), .B(n36610), .Z(n36599) );
  AND U36157 ( .A(n36611), .B(n36612), .Z(n36610) );
  XNOR U36158 ( .A(n36609), .B(n36437), .Z(n36612) );
  IV U36159 ( .A(n36440), .Z(n36437) );
  XOR U36160 ( .A(n36613), .B(n36614), .Z(n36440) );
  AND U36161 ( .A(n717), .B(n36615), .Z(n36614) );
  XOR U36162 ( .A(n36616), .B(n36613), .Z(n36615) );
  XOR U36163 ( .A(n36441), .B(n36609), .Z(n36611) );
  XOR U36164 ( .A(n36617), .B(n36618), .Z(n36441) );
  AND U36165 ( .A(n725), .B(n36577), .Z(n36618) );
  XOR U36166 ( .A(n36617), .B(n36575), .Z(n36577) );
  XOR U36167 ( .A(n36619), .B(n36620), .Z(n36609) );
  AND U36168 ( .A(n36621), .B(n36622), .Z(n36620) );
  XNOR U36169 ( .A(n36619), .B(n36465), .Z(n36622) );
  IV U36170 ( .A(n36468), .Z(n36465) );
  XOR U36171 ( .A(n36623), .B(n36624), .Z(n36468) );
  AND U36172 ( .A(n717), .B(n36625), .Z(n36624) );
  XNOR U36173 ( .A(n36626), .B(n36623), .Z(n36625) );
  XOR U36174 ( .A(n36469), .B(n36619), .Z(n36621) );
  XOR U36175 ( .A(n36627), .B(n36628), .Z(n36469) );
  AND U36176 ( .A(n725), .B(n36586), .Z(n36628) );
  XOR U36177 ( .A(n36627), .B(n36584), .Z(n36586) );
  XOR U36178 ( .A(n36543), .B(n36629), .Z(n36619) );
  AND U36179 ( .A(n36545), .B(n36630), .Z(n36629) );
  XNOR U36180 ( .A(n36543), .B(n36514), .Z(n36630) );
  IV U36181 ( .A(n36517), .Z(n36514) );
  XOR U36182 ( .A(n36631), .B(n36632), .Z(n36517) );
  AND U36183 ( .A(n717), .B(n36633), .Z(n36632) );
  XOR U36184 ( .A(n36634), .B(n36631), .Z(n36633) );
  XOR U36185 ( .A(n36518), .B(n36543), .Z(n36545) );
  XOR U36186 ( .A(n36635), .B(n36636), .Z(n36518) );
  AND U36187 ( .A(n725), .B(n36596), .Z(n36636) );
  XOR U36188 ( .A(n36635), .B(n36594), .Z(n36596) );
  AND U36189 ( .A(n36597), .B(n36527), .Z(n36543) );
  XNOR U36190 ( .A(n36637), .B(n36638), .Z(n36527) );
  AND U36191 ( .A(n717), .B(n36639), .Z(n36638) );
  XNOR U36192 ( .A(n36640), .B(n36637), .Z(n36639) );
  XNOR U36193 ( .A(n36641), .B(n36642), .Z(n717) );
  AND U36194 ( .A(n36643), .B(n36644), .Z(n36642) );
  XOR U36195 ( .A(n36606), .B(n36641), .Z(n36644) );
  AND U36196 ( .A(n36645), .B(n36646), .Z(n36606) );
  XNOR U36197 ( .A(n36603), .B(n36641), .Z(n36643) );
  XNOR U36198 ( .A(n36647), .B(n36648), .Z(n36603) );
  AND U36199 ( .A(n721), .B(n36649), .Z(n36648) );
  XNOR U36200 ( .A(n36650), .B(n36651), .Z(n36649) );
  XOR U36201 ( .A(n36652), .B(n36653), .Z(n36641) );
  AND U36202 ( .A(n36654), .B(n36655), .Z(n36653) );
  XNOR U36203 ( .A(n36652), .B(n36645), .Z(n36655) );
  IV U36204 ( .A(n36616), .Z(n36645) );
  XOR U36205 ( .A(n36656), .B(n36657), .Z(n36616) );
  XOR U36206 ( .A(n36658), .B(n36646), .Z(n36657) );
  AND U36207 ( .A(n36626), .B(n36659), .Z(n36646) );
  AND U36208 ( .A(n36660), .B(n36661), .Z(n36658) );
  XOR U36209 ( .A(n36662), .B(n36656), .Z(n36660) );
  XNOR U36210 ( .A(n36613), .B(n36652), .Z(n36654) );
  XNOR U36211 ( .A(n36663), .B(n36664), .Z(n36613) );
  AND U36212 ( .A(n721), .B(n36665), .Z(n36664) );
  XNOR U36213 ( .A(n36666), .B(n36667), .Z(n36665) );
  XOR U36214 ( .A(n36668), .B(n36669), .Z(n36652) );
  AND U36215 ( .A(n36670), .B(n36671), .Z(n36669) );
  XNOR U36216 ( .A(n36668), .B(n36626), .Z(n36671) );
  XOR U36217 ( .A(n36672), .B(n36661), .Z(n36626) );
  XNOR U36218 ( .A(n36673), .B(n36656), .Z(n36661) );
  XOR U36219 ( .A(n36674), .B(n36675), .Z(n36656) );
  AND U36220 ( .A(n36676), .B(n36677), .Z(n36675) );
  XOR U36221 ( .A(n36678), .B(n36674), .Z(n36676) );
  XNOR U36222 ( .A(n36679), .B(n36680), .Z(n36673) );
  AND U36223 ( .A(n36681), .B(n36682), .Z(n36680) );
  XOR U36224 ( .A(n36679), .B(n36683), .Z(n36681) );
  XNOR U36225 ( .A(n36662), .B(n36659), .Z(n36672) );
  AND U36226 ( .A(n36684), .B(n36685), .Z(n36659) );
  XOR U36227 ( .A(n36686), .B(n36687), .Z(n36662) );
  AND U36228 ( .A(n36688), .B(n36689), .Z(n36687) );
  XOR U36229 ( .A(n36686), .B(n36690), .Z(n36688) );
  XNOR U36230 ( .A(n36623), .B(n36668), .Z(n36670) );
  XNOR U36231 ( .A(n36691), .B(n36692), .Z(n36623) );
  AND U36232 ( .A(n721), .B(n36693), .Z(n36692) );
  XNOR U36233 ( .A(n36694), .B(n36695), .Z(n36693) );
  XOR U36234 ( .A(n36696), .B(n36697), .Z(n36668) );
  AND U36235 ( .A(n36698), .B(n36699), .Z(n36697) );
  XNOR U36236 ( .A(n36696), .B(n36684), .Z(n36699) );
  IV U36237 ( .A(n36634), .Z(n36684) );
  XNOR U36238 ( .A(n36700), .B(n36677), .Z(n36634) );
  XNOR U36239 ( .A(n36701), .B(n36683), .Z(n36677) );
  XOR U36240 ( .A(n36702), .B(n36703), .Z(n36683) );
  NOR U36241 ( .A(n36704), .B(n36705), .Z(n36703) );
  XNOR U36242 ( .A(n36702), .B(n36706), .Z(n36704) );
  XNOR U36243 ( .A(n36682), .B(n36674), .Z(n36701) );
  XOR U36244 ( .A(n36707), .B(n36708), .Z(n36674) );
  AND U36245 ( .A(n36709), .B(n36710), .Z(n36708) );
  XNOR U36246 ( .A(n36707), .B(n36711), .Z(n36709) );
  XNOR U36247 ( .A(n36712), .B(n36679), .Z(n36682) );
  XOR U36248 ( .A(n36713), .B(n36714), .Z(n36679) );
  AND U36249 ( .A(n36715), .B(n36716), .Z(n36714) );
  XOR U36250 ( .A(n36713), .B(n36717), .Z(n36715) );
  XNOR U36251 ( .A(n36718), .B(n36719), .Z(n36712) );
  NOR U36252 ( .A(n36720), .B(n36721), .Z(n36719) );
  XOR U36253 ( .A(n36718), .B(n36722), .Z(n36720) );
  XNOR U36254 ( .A(n36678), .B(n36685), .Z(n36700) );
  NOR U36255 ( .A(n36640), .B(n36723), .Z(n36685) );
  XOR U36256 ( .A(n36690), .B(n36689), .Z(n36678) );
  XNOR U36257 ( .A(n36724), .B(n36686), .Z(n36689) );
  XOR U36258 ( .A(n36725), .B(n36726), .Z(n36686) );
  AND U36259 ( .A(n36727), .B(n36728), .Z(n36726) );
  XOR U36260 ( .A(n36725), .B(n36729), .Z(n36727) );
  XNOR U36261 ( .A(n36730), .B(n36731), .Z(n36724) );
  NOR U36262 ( .A(n36732), .B(n36733), .Z(n36731) );
  XNOR U36263 ( .A(n36730), .B(n36734), .Z(n36732) );
  XOR U36264 ( .A(n36735), .B(n36736), .Z(n36690) );
  NOR U36265 ( .A(n36737), .B(n36738), .Z(n36736) );
  XNOR U36266 ( .A(n36735), .B(n36739), .Z(n36737) );
  XNOR U36267 ( .A(n36631), .B(n36696), .Z(n36698) );
  XNOR U36268 ( .A(n36740), .B(n36741), .Z(n36631) );
  AND U36269 ( .A(n721), .B(n36742), .Z(n36741) );
  XNOR U36270 ( .A(n36743), .B(n36744), .Z(n36742) );
  AND U36271 ( .A(n36637), .B(n36640), .Z(n36696) );
  XOR U36272 ( .A(n36745), .B(n36723), .Z(n36640) );
  XNOR U36273 ( .A(p_input[2048]), .B(p_input[544]), .Z(n36723) );
  XOR U36274 ( .A(n36711), .B(n36710), .Z(n36745) );
  XNOR U36275 ( .A(n36746), .B(n36717), .Z(n36710) );
  XNOR U36276 ( .A(n36706), .B(n36705), .Z(n36717) );
  XOR U36277 ( .A(n36747), .B(n36702), .Z(n36705) );
  XNOR U36278 ( .A(n29266), .B(p_input[554]), .Z(n36702) );
  XNOR U36279 ( .A(p_input[2059]), .B(p_input[555]), .Z(n36747) );
  XOR U36280 ( .A(p_input[2060]), .B(p_input[556]), .Z(n36706) );
  XNOR U36281 ( .A(n36716), .B(n36707), .Z(n36746) );
  XNOR U36282 ( .A(n29494), .B(p_input[545]), .Z(n36707) );
  XOR U36283 ( .A(n36748), .B(n36722), .Z(n36716) );
  XNOR U36284 ( .A(p_input[2063]), .B(p_input[559]), .Z(n36722) );
  XOR U36285 ( .A(n36713), .B(n36721), .Z(n36748) );
  XOR U36286 ( .A(n36749), .B(n36718), .Z(n36721) );
  XOR U36287 ( .A(p_input[2061]), .B(p_input[557]), .Z(n36718) );
  XNOR U36288 ( .A(p_input[2062]), .B(p_input[558]), .Z(n36749) );
  XNOR U36289 ( .A(n29036), .B(p_input[553]), .Z(n36713) );
  XNOR U36290 ( .A(n36729), .B(n36728), .Z(n36711) );
  XNOR U36291 ( .A(n36750), .B(n36734), .Z(n36728) );
  XOR U36292 ( .A(p_input[2056]), .B(p_input[552]), .Z(n36734) );
  XOR U36293 ( .A(n36725), .B(n36733), .Z(n36750) );
  XOR U36294 ( .A(n36751), .B(n36730), .Z(n36733) );
  XOR U36295 ( .A(p_input[2054]), .B(p_input[550]), .Z(n36730) );
  XNOR U36296 ( .A(p_input[2055]), .B(p_input[551]), .Z(n36751) );
  XNOR U36297 ( .A(n29039), .B(p_input[546]), .Z(n36725) );
  XNOR U36298 ( .A(n36739), .B(n36738), .Z(n36729) );
  XOR U36299 ( .A(n36752), .B(n36735), .Z(n36738) );
  XOR U36300 ( .A(p_input[2051]), .B(p_input[547]), .Z(n36735) );
  XNOR U36301 ( .A(p_input[2052]), .B(p_input[548]), .Z(n36752) );
  XOR U36302 ( .A(p_input[2053]), .B(p_input[549]), .Z(n36739) );
  XNOR U36303 ( .A(n36753), .B(n36754), .Z(n36637) );
  AND U36304 ( .A(n721), .B(n36755), .Z(n36754) );
  XNOR U36305 ( .A(n36756), .B(n36757), .Z(n721) );
  AND U36306 ( .A(n36758), .B(n36759), .Z(n36757) );
  XOR U36307 ( .A(n36651), .B(n36756), .Z(n36759) );
  XNOR U36308 ( .A(n36760), .B(n36756), .Z(n36758) );
  XOR U36309 ( .A(n36761), .B(n36762), .Z(n36756) );
  AND U36310 ( .A(n36763), .B(n36764), .Z(n36762) );
  XOR U36311 ( .A(n36666), .B(n36761), .Z(n36764) );
  XOR U36312 ( .A(n36761), .B(n36667), .Z(n36763) );
  XOR U36313 ( .A(n36765), .B(n36766), .Z(n36761) );
  AND U36314 ( .A(n36767), .B(n36768), .Z(n36766) );
  XOR U36315 ( .A(n36694), .B(n36765), .Z(n36768) );
  XOR U36316 ( .A(n36765), .B(n36695), .Z(n36767) );
  XOR U36317 ( .A(n36769), .B(n36770), .Z(n36765) );
  AND U36318 ( .A(n36771), .B(n36772), .Z(n36770) );
  XOR U36319 ( .A(n36769), .B(n36743), .Z(n36772) );
  XNOR U36320 ( .A(n36773), .B(n36774), .Z(n36597) );
  AND U36321 ( .A(n725), .B(n36775), .Z(n36774) );
  XNOR U36322 ( .A(n36776), .B(n36777), .Z(n725) );
  AND U36323 ( .A(n36778), .B(n36779), .Z(n36777) );
  XOR U36324 ( .A(n36776), .B(n36607), .Z(n36779) );
  XNOR U36325 ( .A(n36776), .B(n36567), .Z(n36778) );
  XOR U36326 ( .A(n36780), .B(n36781), .Z(n36776) );
  AND U36327 ( .A(n36782), .B(n36783), .Z(n36781) );
  XOR U36328 ( .A(n36780), .B(n36575), .Z(n36782) );
  XOR U36329 ( .A(n36784), .B(n36785), .Z(n36558) );
  AND U36330 ( .A(n729), .B(n36775), .Z(n36785) );
  XNOR U36331 ( .A(n36773), .B(n36784), .Z(n36775) );
  XNOR U36332 ( .A(n36786), .B(n36787), .Z(n729) );
  AND U36333 ( .A(n36788), .B(n36789), .Z(n36787) );
  XNOR U36334 ( .A(n36790), .B(n36786), .Z(n36789) );
  IV U36335 ( .A(n36607), .Z(n36790) );
  XOR U36336 ( .A(n36760), .B(n36791), .Z(n36607) );
  AND U36337 ( .A(n732), .B(n36792), .Z(n36791) );
  XOR U36338 ( .A(n36650), .B(n36647), .Z(n36792) );
  IV U36339 ( .A(n36760), .Z(n36650) );
  XNOR U36340 ( .A(n36567), .B(n36786), .Z(n36788) );
  XOR U36341 ( .A(n36793), .B(n36794), .Z(n36567) );
  AND U36342 ( .A(n748), .B(n36795), .Z(n36794) );
  XOR U36343 ( .A(n36780), .B(n36796), .Z(n36786) );
  AND U36344 ( .A(n36797), .B(n36783), .Z(n36796) );
  XNOR U36345 ( .A(n36617), .B(n36780), .Z(n36783) );
  XOR U36346 ( .A(n36667), .B(n36798), .Z(n36617) );
  AND U36347 ( .A(n732), .B(n36799), .Z(n36798) );
  XOR U36348 ( .A(n36663), .B(n36667), .Z(n36799) );
  XNOR U36349 ( .A(n36800), .B(n36780), .Z(n36797) );
  IV U36350 ( .A(n36575), .Z(n36800) );
  XOR U36351 ( .A(n36801), .B(n36802), .Z(n36575) );
  AND U36352 ( .A(n748), .B(n36803), .Z(n36802) );
  XOR U36353 ( .A(n36804), .B(n36805), .Z(n36780) );
  AND U36354 ( .A(n36806), .B(n36807), .Z(n36805) );
  XNOR U36355 ( .A(n36627), .B(n36804), .Z(n36807) );
  XOR U36356 ( .A(n36695), .B(n36808), .Z(n36627) );
  AND U36357 ( .A(n732), .B(n36809), .Z(n36808) );
  XOR U36358 ( .A(n36691), .B(n36695), .Z(n36809) );
  XOR U36359 ( .A(n36804), .B(n36584), .Z(n36806) );
  XOR U36360 ( .A(n36810), .B(n36811), .Z(n36584) );
  AND U36361 ( .A(n748), .B(n36812), .Z(n36811) );
  XOR U36362 ( .A(n36813), .B(n36814), .Z(n36804) );
  AND U36363 ( .A(n36815), .B(n36816), .Z(n36814) );
  XNOR U36364 ( .A(n36813), .B(n36635), .Z(n36816) );
  XOR U36365 ( .A(n36744), .B(n36817), .Z(n36635) );
  AND U36366 ( .A(n732), .B(n36818), .Z(n36817) );
  XOR U36367 ( .A(n36740), .B(n36744), .Z(n36818) );
  XNOR U36368 ( .A(n36819), .B(n36813), .Z(n36815) );
  IV U36369 ( .A(n36594), .Z(n36819) );
  XOR U36370 ( .A(n36820), .B(n36821), .Z(n36594) );
  AND U36371 ( .A(n748), .B(n36822), .Z(n36821) );
  AND U36372 ( .A(n36784), .B(n36773), .Z(n36813) );
  XNOR U36373 ( .A(n36823), .B(n36824), .Z(n36773) );
  AND U36374 ( .A(n732), .B(n36755), .Z(n36824) );
  XNOR U36375 ( .A(n36753), .B(n36823), .Z(n36755) );
  XNOR U36376 ( .A(n36825), .B(n36826), .Z(n732) );
  AND U36377 ( .A(n36827), .B(n36828), .Z(n36826) );
  XNOR U36378 ( .A(n36825), .B(n36647), .Z(n36828) );
  IV U36379 ( .A(n36651), .Z(n36647) );
  XOR U36380 ( .A(n36829), .B(n36830), .Z(n36651) );
  AND U36381 ( .A(n736), .B(n36831), .Z(n36830) );
  XOR U36382 ( .A(n36832), .B(n36829), .Z(n36831) );
  XNOR U36383 ( .A(n36825), .B(n36760), .Z(n36827) );
  XOR U36384 ( .A(n36833), .B(n36834), .Z(n36760) );
  AND U36385 ( .A(n744), .B(n36795), .Z(n36834) );
  XOR U36386 ( .A(n36793), .B(n36833), .Z(n36795) );
  XOR U36387 ( .A(n36835), .B(n36836), .Z(n36825) );
  AND U36388 ( .A(n36837), .B(n36838), .Z(n36836) );
  XNOR U36389 ( .A(n36835), .B(n36663), .Z(n36838) );
  IV U36390 ( .A(n36666), .Z(n36663) );
  XOR U36391 ( .A(n36839), .B(n36840), .Z(n36666) );
  AND U36392 ( .A(n736), .B(n36841), .Z(n36840) );
  XOR U36393 ( .A(n36842), .B(n36839), .Z(n36841) );
  XOR U36394 ( .A(n36667), .B(n36835), .Z(n36837) );
  XOR U36395 ( .A(n36843), .B(n36844), .Z(n36667) );
  AND U36396 ( .A(n744), .B(n36803), .Z(n36844) );
  XOR U36397 ( .A(n36843), .B(n36801), .Z(n36803) );
  XOR U36398 ( .A(n36845), .B(n36846), .Z(n36835) );
  AND U36399 ( .A(n36847), .B(n36848), .Z(n36846) );
  XNOR U36400 ( .A(n36845), .B(n36691), .Z(n36848) );
  IV U36401 ( .A(n36694), .Z(n36691) );
  XOR U36402 ( .A(n36849), .B(n36850), .Z(n36694) );
  AND U36403 ( .A(n736), .B(n36851), .Z(n36850) );
  XNOR U36404 ( .A(n36852), .B(n36849), .Z(n36851) );
  XOR U36405 ( .A(n36695), .B(n36845), .Z(n36847) );
  XOR U36406 ( .A(n36853), .B(n36854), .Z(n36695) );
  AND U36407 ( .A(n744), .B(n36812), .Z(n36854) );
  XOR U36408 ( .A(n36853), .B(n36810), .Z(n36812) );
  XOR U36409 ( .A(n36769), .B(n36855), .Z(n36845) );
  AND U36410 ( .A(n36771), .B(n36856), .Z(n36855) );
  XNOR U36411 ( .A(n36769), .B(n36740), .Z(n36856) );
  IV U36412 ( .A(n36743), .Z(n36740) );
  XOR U36413 ( .A(n36857), .B(n36858), .Z(n36743) );
  AND U36414 ( .A(n736), .B(n36859), .Z(n36858) );
  XOR U36415 ( .A(n36860), .B(n36857), .Z(n36859) );
  XOR U36416 ( .A(n36744), .B(n36769), .Z(n36771) );
  XOR U36417 ( .A(n36861), .B(n36862), .Z(n36744) );
  AND U36418 ( .A(n744), .B(n36822), .Z(n36862) );
  XOR U36419 ( .A(n36861), .B(n36820), .Z(n36822) );
  AND U36420 ( .A(n36823), .B(n36753), .Z(n36769) );
  XNOR U36421 ( .A(n36863), .B(n36864), .Z(n36753) );
  AND U36422 ( .A(n736), .B(n36865), .Z(n36864) );
  XNOR U36423 ( .A(n36866), .B(n36863), .Z(n36865) );
  XNOR U36424 ( .A(n36867), .B(n36868), .Z(n736) );
  AND U36425 ( .A(n36869), .B(n36870), .Z(n36868) );
  XOR U36426 ( .A(n36832), .B(n36867), .Z(n36870) );
  AND U36427 ( .A(n36871), .B(n36872), .Z(n36832) );
  XNOR U36428 ( .A(n36829), .B(n36867), .Z(n36869) );
  XNOR U36429 ( .A(n36873), .B(n36874), .Z(n36829) );
  AND U36430 ( .A(n740), .B(n36875), .Z(n36874) );
  XNOR U36431 ( .A(n36876), .B(n36877), .Z(n36875) );
  XOR U36432 ( .A(n36878), .B(n36879), .Z(n36867) );
  AND U36433 ( .A(n36880), .B(n36881), .Z(n36879) );
  XNOR U36434 ( .A(n36878), .B(n36871), .Z(n36881) );
  IV U36435 ( .A(n36842), .Z(n36871) );
  XOR U36436 ( .A(n36882), .B(n36883), .Z(n36842) );
  XOR U36437 ( .A(n36884), .B(n36872), .Z(n36883) );
  AND U36438 ( .A(n36852), .B(n36885), .Z(n36872) );
  AND U36439 ( .A(n36886), .B(n36887), .Z(n36884) );
  XOR U36440 ( .A(n36888), .B(n36882), .Z(n36886) );
  XNOR U36441 ( .A(n36839), .B(n36878), .Z(n36880) );
  XNOR U36442 ( .A(n36889), .B(n36890), .Z(n36839) );
  AND U36443 ( .A(n740), .B(n36891), .Z(n36890) );
  XNOR U36444 ( .A(n36892), .B(n36893), .Z(n36891) );
  XOR U36445 ( .A(n36894), .B(n36895), .Z(n36878) );
  AND U36446 ( .A(n36896), .B(n36897), .Z(n36895) );
  XNOR U36447 ( .A(n36894), .B(n36852), .Z(n36897) );
  XOR U36448 ( .A(n36898), .B(n36887), .Z(n36852) );
  XNOR U36449 ( .A(n36899), .B(n36882), .Z(n36887) );
  XOR U36450 ( .A(n36900), .B(n36901), .Z(n36882) );
  AND U36451 ( .A(n36902), .B(n36903), .Z(n36901) );
  XOR U36452 ( .A(n36904), .B(n36900), .Z(n36902) );
  XNOR U36453 ( .A(n36905), .B(n36906), .Z(n36899) );
  AND U36454 ( .A(n36907), .B(n36908), .Z(n36906) );
  XOR U36455 ( .A(n36905), .B(n36909), .Z(n36907) );
  XNOR U36456 ( .A(n36888), .B(n36885), .Z(n36898) );
  AND U36457 ( .A(n36910), .B(n36911), .Z(n36885) );
  XOR U36458 ( .A(n36912), .B(n36913), .Z(n36888) );
  AND U36459 ( .A(n36914), .B(n36915), .Z(n36913) );
  XOR U36460 ( .A(n36912), .B(n36916), .Z(n36914) );
  XNOR U36461 ( .A(n36849), .B(n36894), .Z(n36896) );
  XNOR U36462 ( .A(n36917), .B(n36918), .Z(n36849) );
  AND U36463 ( .A(n740), .B(n36919), .Z(n36918) );
  XNOR U36464 ( .A(n36920), .B(n36921), .Z(n36919) );
  XOR U36465 ( .A(n36922), .B(n36923), .Z(n36894) );
  AND U36466 ( .A(n36924), .B(n36925), .Z(n36923) );
  XNOR U36467 ( .A(n36922), .B(n36910), .Z(n36925) );
  IV U36468 ( .A(n36860), .Z(n36910) );
  XNOR U36469 ( .A(n36926), .B(n36903), .Z(n36860) );
  XNOR U36470 ( .A(n36927), .B(n36909), .Z(n36903) );
  XOR U36471 ( .A(n36928), .B(n36929), .Z(n36909) );
  NOR U36472 ( .A(n36930), .B(n36931), .Z(n36929) );
  XNOR U36473 ( .A(n36928), .B(n36932), .Z(n36930) );
  XNOR U36474 ( .A(n36908), .B(n36900), .Z(n36927) );
  XOR U36475 ( .A(n36933), .B(n36934), .Z(n36900) );
  AND U36476 ( .A(n36935), .B(n36936), .Z(n36934) );
  XNOR U36477 ( .A(n36933), .B(n36937), .Z(n36935) );
  XNOR U36478 ( .A(n36938), .B(n36905), .Z(n36908) );
  XOR U36479 ( .A(n36939), .B(n36940), .Z(n36905) );
  AND U36480 ( .A(n36941), .B(n36942), .Z(n36940) );
  XOR U36481 ( .A(n36939), .B(n36943), .Z(n36941) );
  XNOR U36482 ( .A(n36944), .B(n36945), .Z(n36938) );
  NOR U36483 ( .A(n36946), .B(n36947), .Z(n36945) );
  XOR U36484 ( .A(n36944), .B(n36948), .Z(n36946) );
  XNOR U36485 ( .A(n36904), .B(n36911), .Z(n36926) );
  NOR U36486 ( .A(n36866), .B(n36949), .Z(n36911) );
  XOR U36487 ( .A(n36916), .B(n36915), .Z(n36904) );
  XNOR U36488 ( .A(n36950), .B(n36912), .Z(n36915) );
  XOR U36489 ( .A(n36951), .B(n36952), .Z(n36912) );
  AND U36490 ( .A(n36953), .B(n36954), .Z(n36952) );
  XOR U36491 ( .A(n36951), .B(n36955), .Z(n36953) );
  XNOR U36492 ( .A(n36956), .B(n36957), .Z(n36950) );
  NOR U36493 ( .A(n36958), .B(n36959), .Z(n36957) );
  XNOR U36494 ( .A(n36956), .B(n36960), .Z(n36958) );
  XOR U36495 ( .A(n36961), .B(n36962), .Z(n36916) );
  NOR U36496 ( .A(n36963), .B(n36964), .Z(n36962) );
  XNOR U36497 ( .A(n36961), .B(n36965), .Z(n36963) );
  XNOR U36498 ( .A(n36857), .B(n36922), .Z(n36924) );
  XNOR U36499 ( .A(n36966), .B(n36967), .Z(n36857) );
  AND U36500 ( .A(n740), .B(n36968), .Z(n36967) );
  XNOR U36501 ( .A(n36969), .B(n36970), .Z(n36968) );
  AND U36502 ( .A(n36863), .B(n36866), .Z(n36922) );
  XOR U36503 ( .A(n36971), .B(n36949), .Z(n36866) );
  XNOR U36504 ( .A(p_input[2048]), .B(p_input[560]), .Z(n36949) );
  XOR U36505 ( .A(n36937), .B(n36936), .Z(n36971) );
  XNOR U36506 ( .A(n36972), .B(n36943), .Z(n36936) );
  XNOR U36507 ( .A(n36932), .B(n36931), .Z(n36943) );
  XOR U36508 ( .A(n36973), .B(n36928), .Z(n36931) );
  XNOR U36509 ( .A(n29266), .B(p_input[570]), .Z(n36928) );
  XNOR U36510 ( .A(p_input[2059]), .B(p_input[571]), .Z(n36973) );
  XOR U36511 ( .A(p_input[2060]), .B(p_input[572]), .Z(n36932) );
  XNOR U36512 ( .A(n36942), .B(n36933), .Z(n36972) );
  XNOR U36513 ( .A(n29494), .B(p_input[561]), .Z(n36933) );
  XOR U36514 ( .A(n36974), .B(n36948), .Z(n36942) );
  XNOR U36515 ( .A(p_input[2063]), .B(p_input[575]), .Z(n36948) );
  XOR U36516 ( .A(n36939), .B(n36947), .Z(n36974) );
  XOR U36517 ( .A(n36975), .B(n36944), .Z(n36947) );
  XOR U36518 ( .A(p_input[2061]), .B(p_input[573]), .Z(n36944) );
  XNOR U36519 ( .A(p_input[2062]), .B(p_input[574]), .Z(n36975) );
  XNOR U36520 ( .A(n29036), .B(p_input[569]), .Z(n36939) );
  XNOR U36521 ( .A(n36955), .B(n36954), .Z(n36937) );
  XNOR U36522 ( .A(n36976), .B(n36960), .Z(n36954) );
  XOR U36523 ( .A(p_input[2056]), .B(p_input[568]), .Z(n36960) );
  XOR U36524 ( .A(n36951), .B(n36959), .Z(n36976) );
  XOR U36525 ( .A(n36977), .B(n36956), .Z(n36959) );
  XOR U36526 ( .A(p_input[2054]), .B(p_input[566]), .Z(n36956) );
  XNOR U36527 ( .A(p_input[2055]), .B(p_input[567]), .Z(n36977) );
  XNOR U36528 ( .A(n29039), .B(p_input[562]), .Z(n36951) );
  XNOR U36529 ( .A(n36965), .B(n36964), .Z(n36955) );
  XOR U36530 ( .A(n36978), .B(n36961), .Z(n36964) );
  XOR U36531 ( .A(p_input[2051]), .B(p_input[563]), .Z(n36961) );
  XNOR U36532 ( .A(p_input[2052]), .B(p_input[564]), .Z(n36978) );
  XOR U36533 ( .A(p_input[2053]), .B(p_input[565]), .Z(n36965) );
  XNOR U36534 ( .A(n36979), .B(n36980), .Z(n36863) );
  AND U36535 ( .A(n740), .B(n36981), .Z(n36980) );
  XNOR U36536 ( .A(n36982), .B(n36983), .Z(n740) );
  AND U36537 ( .A(n36984), .B(n36985), .Z(n36983) );
  XOR U36538 ( .A(n36877), .B(n36982), .Z(n36985) );
  XNOR U36539 ( .A(n36986), .B(n36982), .Z(n36984) );
  XOR U36540 ( .A(n36987), .B(n36988), .Z(n36982) );
  AND U36541 ( .A(n36989), .B(n36990), .Z(n36988) );
  XOR U36542 ( .A(n36892), .B(n36987), .Z(n36990) );
  XOR U36543 ( .A(n36987), .B(n36893), .Z(n36989) );
  XOR U36544 ( .A(n36991), .B(n36992), .Z(n36987) );
  AND U36545 ( .A(n36993), .B(n36994), .Z(n36992) );
  XOR U36546 ( .A(n36920), .B(n36991), .Z(n36994) );
  XOR U36547 ( .A(n36991), .B(n36921), .Z(n36993) );
  XOR U36548 ( .A(n36995), .B(n36996), .Z(n36991) );
  AND U36549 ( .A(n36997), .B(n36998), .Z(n36996) );
  XOR U36550 ( .A(n36995), .B(n36969), .Z(n36998) );
  XNOR U36551 ( .A(n36999), .B(n37000), .Z(n36823) );
  AND U36552 ( .A(n744), .B(n37001), .Z(n37000) );
  XNOR U36553 ( .A(n37002), .B(n37003), .Z(n744) );
  AND U36554 ( .A(n37004), .B(n37005), .Z(n37003) );
  XOR U36555 ( .A(n37002), .B(n36833), .Z(n37005) );
  XNOR U36556 ( .A(n37002), .B(n36793), .Z(n37004) );
  XOR U36557 ( .A(n37006), .B(n37007), .Z(n37002) );
  AND U36558 ( .A(n37008), .B(n37009), .Z(n37007) );
  XOR U36559 ( .A(n37006), .B(n36801), .Z(n37008) );
  XOR U36560 ( .A(n37010), .B(n37011), .Z(n36784) );
  AND U36561 ( .A(n748), .B(n37001), .Z(n37011) );
  XNOR U36562 ( .A(n36999), .B(n37010), .Z(n37001) );
  XNOR U36563 ( .A(n37012), .B(n37013), .Z(n748) );
  AND U36564 ( .A(n37014), .B(n37015), .Z(n37013) );
  XNOR U36565 ( .A(n37016), .B(n37012), .Z(n37015) );
  IV U36566 ( .A(n36833), .Z(n37016) );
  XOR U36567 ( .A(n36986), .B(n37017), .Z(n36833) );
  AND U36568 ( .A(n751), .B(n37018), .Z(n37017) );
  XOR U36569 ( .A(n36876), .B(n36873), .Z(n37018) );
  IV U36570 ( .A(n36986), .Z(n36876) );
  XNOR U36571 ( .A(n36793), .B(n37012), .Z(n37014) );
  XOR U36572 ( .A(n37019), .B(n37020), .Z(n36793) );
  AND U36573 ( .A(n767), .B(n37021), .Z(n37020) );
  XOR U36574 ( .A(n37006), .B(n37022), .Z(n37012) );
  AND U36575 ( .A(n37023), .B(n37009), .Z(n37022) );
  XNOR U36576 ( .A(n36843), .B(n37006), .Z(n37009) );
  XOR U36577 ( .A(n36893), .B(n37024), .Z(n36843) );
  AND U36578 ( .A(n751), .B(n37025), .Z(n37024) );
  XOR U36579 ( .A(n36889), .B(n36893), .Z(n37025) );
  XNOR U36580 ( .A(n37026), .B(n37006), .Z(n37023) );
  IV U36581 ( .A(n36801), .Z(n37026) );
  XOR U36582 ( .A(n37027), .B(n37028), .Z(n36801) );
  AND U36583 ( .A(n767), .B(n37029), .Z(n37028) );
  XOR U36584 ( .A(n37030), .B(n37031), .Z(n37006) );
  AND U36585 ( .A(n37032), .B(n37033), .Z(n37031) );
  XNOR U36586 ( .A(n36853), .B(n37030), .Z(n37033) );
  XOR U36587 ( .A(n36921), .B(n37034), .Z(n36853) );
  AND U36588 ( .A(n751), .B(n37035), .Z(n37034) );
  XOR U36589 ( .A(n36917), .B(n36921), .Z(n37035) );
  XOR U36590 ( .A(n37030), .B(n36810), .Z(n37032) );
  XOR U36591 ( .A(n37036), .B(n37037), .Z(n36810) );
  AND U36592 ( .A(n767), .B(n37038), .Z(n37037) );
  XOR U36593 ( .A(n37039), .B(n37040), .Z(n37030) );
  AND U36594 ( .A(n37041), .B(n37042), .Z(n37040) );
  XNOR U36595 ( .A(n37039), .B(n36861), .Z(n37042) );
  XOR U36596 ( .A(n36970), .B(n37043), .Z(n36861) );
  AND U36597 ( .A(n751), .B(n37044), .Z(n37043) );
  XOR U36598 ( .A(n36966), .B(n36970), .Z(n37044) );
  XNOR U36599 ( .A(n37045), .B(n37039), .Z(n37041) );
  IV U36600 ( .A(n36820), .Z(n37045) );
  XOR U36601 ( .A(n37046), .B(n37047), .Z(n36820) );
  AND U36602 ( .A(n767), .B(n37048), .Z(n37047) );
  AND U36603 ( .A(n37010), .B(n36999), .Z(n37039) );
  XNOR U36604 ( .A(n37049), .B(n37050), .Z(n36999) );
  AND U36605 ( .A(n751), .B(n36981), .Z(n37050) );
  XNOR U36606 ( .A(n36979), .B(n37049), .Z(n36981) );
  XNOR U36607 ( .A(n37051), .B(n37052), .Z(n751) );
  AND U36608 ( .A(n37053), .B(n37054), .Z(n37052) );
  XNOR U36609 ( .A(n37051), .B(n36873), .Z(n37054) );
  IV U36610 ( .A(n36877), .Z(n36873) );
  XOR U36611 ( .A(n37055), .B(n37056), .Z(n36877) );
  AND U36612 ( .A(n755), .B(n37057), .Z(n37056) );
  XOR U36613 ( .A(n37058), .B(n37055), .Z(n37057) );
  XNOR U36614 ( .A(n37051), .B(n36986), .Z(n37053) );
  XOR U36615 ( .A(n37059), .B(n37060), .Z(n36986) );
  AND U36616 ( .A(n763), .B(n37021), .Z(n37060) );
  XOR U36617 ( .A(n37019), .B(n37059), .Z(n37021) );
  XOR U36618 ( .A(n37061), .B(n37062), .Z(n37051) );
  AND U36619 ( .A(n37063), .B(n37064), .Z(n37062) );
  XNOR U36620 ( .A(n37061), .B(n36889), .Z(n37064) );
  IV U36621 ( .A(n36892), .Z(n36889) );
  XOR U36622 ( .A(n37065), .B(n37066), .Z(n36892) );
  AND U36623 ( .A(n755), .B(n37067), .Z(n37066) );
  XOR U36624 ( .A(n37068), .B(n37065), .Z(n37067) );
  XOR U36625 ( .A(n36893), .B(n37061), .Z(n37063) );
  XOR U36626 ( .A(n37069), .B(n37070), .Z(n36893) );
  AND U36627 ( .A(n763), .B(n37029), .Z(n37070) );
  XOR U36628 ( .A(n37069), .B(n37027), .Z(n37029) );
  XOR U36629 ( .A(n37071), .B(n37072), .Z(n37061) );
  AND U36630 ( .A(n37073), .B(n37074), .Z(n37072) );
  XNOR U36631 ( .A(n37071), .B(n36917), .Z(n37074) );
  IV U36632 ( .A(n36920), .Z(n36917) );
  XOR U36633 ( .A(n37075), .B(n37076), .Z(n36920) );
  AND U36634 ( .A(n755), .B(n37077), .Z(n37076) );
  XNOR U36635 ( .A(n37078), .B(n37075), .Z(n37077) );
  XOR U36636 ( .A(n36921), .B(n37071), .Z(n37073) );
  XOR U36637 ( .A(n37079), .B(n37080), .Z(n36921) );
  AND U36638 ( .A(n763), .B(n37038), .Z(n37080) );
  XOR U36639 ( .A(n37079), .B(n37036), .Z(n37038) );
  XOR U36640 ( .A(n36995), .B(n37081), .Z(n37071) );
  AND U36641 ( .A(n36997), .B(n37082), .Z(n37081) );
  XNOR U36642 ( .A(n36995), .B(n36966), .Z(n37082) );
  IV U36643 ( .A(n36969), .Z(n36966) );
  XOR U36644 ( .A(n37083), .B(n37084), .Z(n36969) );
  AND U36645 ( .A(n755), .B(n37085), .Z(n37084) );
  XOR U36646 ( .A(n37086), .B(n37083), .Z(n37085) );
  XOR U36647 ( .A(n36970), .B(n36995), .Z(n36997) );
  XOR U36648 ( .A(n37087), .B(n37088), .Z(n36970) );
  AND U36649 ( .A(n763), .B(n37048), .Z(n37088) );
  XOR U36650 ( .A(n37087), .B(n37046), .Z(n37048) );
  AND U36651 ( .A(n37049), .B(n36979), .Z(n36995) );
  XNOR U36652 ( .A(n37089), .B(n37090), .Z(n36979) );
  AND U36653 ( .A(n755), .B(n37091), .Z(n37090) );
  XNOR U36654 ( .A(n37092), .B(n37089), .Z(n37091) );
  XNOR U36655 ( .A(n37093), .B(n37094), .Z(n755) );
  AND U36656 ( .A(n37095), .B(n37096), .Z(n37094) );
  XOR U36657 ( .A(n37058), .B(n37093), .Z(n37096) );
  AND U36658 ( .A(n37097), .B(n37098), .Z(n37058) );
  XNOR U36659 ( .A(n37055), .B(n37093), .Z(n37095) );
  XNOR U36660 ( .A(n37099), .B(n37100), .Z(n37055) );
  AND U36661 ( .A(n759), .B(n37101), .Z(n37100) );
  XNOR U36662 ( .A(n37102), .B(n37103), .Z(n37101) );
  XOR U36663 ( .A(n37104), .B(n37105), .Z(n37093) );
  AND U36664 ( .A(n37106), .B(n37107), .Z(n37105) );
  XNOR U36665 ( .A(n37104), .B(n37097), .Z(n37107) );
  IV U36666 ( .A(n37068), .Z(n37097) );
  XOR U36667 ( .A(n37108), .B(n37109), .Z(n37068) );
  XOR U36668 ( .A(n37110), .B(n37098), .Z(n37109) );
  AND U36669 ( .A(n37078), .B(n37111), .Z(n37098) );
  AND U36670 ( .A(n37112), .B(n37113), .Z(n37110) );
  XOR U36671 ( .A(n37114), .B(n37108), .Z(n37112) );
  XNOR U36672 ( .A(n37065), .B(n37104), .Z(n37106) );
  XNOR U36673 ( .A(n37115), .B(n37116), .Z(n37065) );
  AND U36674 ( .A(n759), .B(n37117), .Z(n37116) );
  XNOR U36675 ( .A(n37118), .B(n37119), .Z(n37117) );
  XOR U36676 ( .A(n37120), .B(n37121), .Z(n37104) );
  AND U36677 ( .A(n37122), .B(n37123), .Z(n37121) );
  XNOR U36678 ( .A(n37120), .B(n37078), .Z(n37123) );
  XOR U36679 ( .A(n37124), .B(n37113), .Z(n37078) );
  XNOR U36680 ( .A(n37125), .B(n37108), .Z(n37113) );
  XOR U36681 ( .A(n37126), .B(n37127), .Z(n37108) );
  AND U36682 ( .A(n37128), .B(n37129), .Z(n37127) );
  XOR U36683 ( .A(n37130), .B(n37126), .Z(n37128) );
  XNOR U36684 ( .A(n37131), .B(n37132), .Z(n37125) );
  AND U36685 ( .A(n37133), .B(n37134), .Z(n37132) );
  XOR U36686 ( .A(n37131), .B(n37135), .Z(n37133) );
  XNOR U36687 ( .A(n37114), .B(n37111), .Z(n37124) );
  AND U36688 ( .A(n37136), .B(n37137), .Z(n37111) );
  XOR U36689 ( .A(n37138), .B(n37139), .Z(n37114) );
  AND U36690 ( .A(n37140), .B(n37141), .Z(n37139) );
  XOR U36691 ( .A(n37138), .B(n37142), .Z(n37140) );
  XNOR U36692 ( .A(n37075), .B(n37120), .Z(n37122) );
  XNOR U36693 ( .A(n37143), .B(n37144), .Z(n37075) );
  AND U36694 ( .A(n759), .B(n37145), .Z(n37144) );
  XNOR U36695 ( .A(n37146), .B(n37147), .Z(n37145) );
  XOR U36696 ( .A(n37148), .B(n37149), .Z(n37120) );
  AND U36697 ( .A(n37150), .B(n37151), .Z(n37149) );
  XNOR U36698 ( .A(n37148), .B(n37136), .Z(n37151) );
  IV U36699 ( .A(n37086), .Z(n37136) );
  XNOR U36700 ( .A(n37152), .B(n37129), .Z(n37086) );
  XNOR U36701 ( .A(n37153), .B(n37135), .Z(n37129) );
  XOR U36702 ( .A(n37154), .B(n37155), .Z(n37135) );
  NOR U36703 ( .A(n37156), .B(n37157), .Z(n37155) );
  XNOR U36704 ( .A(n37154), .B(n37158), .Z(n37156) );
  XNOR U36705 ( .A(n37134), .B(n37126), .Z(n37153) );
  XOR U36706 ( .A(n37159), .B(n37160), .Z(n37126) );
  AND U36707 ( .A(n37161), .B(n37162), .Z(n37160) );
  XNOR U36708 ( .A(n37159), .B(n37163), .Z(n37161) );
  XNOR U36709 ( .A(n37164), .B(n37131), .Z(n37134) );
  XOR U36710 ( .A(n37165), .B(n37166), .Z(n37131) );
  AND U36711 ( .A(n37167), .B(n37168), .Z(n37166) );
  XOR U36712 ( .A(n37165), .B(n37169), .Z(n37167) );
  XNOR U36713 ( .A(n37170), .B(n37171), .Z(n37164) );
  NOR U36714 ( .A(n37172), .B(n37173), .Z(n37171) );
  XOR U36715 ( .A(n37170), .B(n37174), .Z(n37172) );
  XNOR U36716 ( .A(n37130), .B(n37137), .Z(n37152) );
  NOR U36717 ( .A(n37092), .B(n37175), .Z(n37137) );
  XOR U36718 ( .A(n37142), .B(n37141), .Z(n37130) );
  XNOR U36719 ( .A(n37176), .B(n37138), .Z(n37141) );
  XOR U36720 ( .A(n37177), .B(n37178), .Z(n37138) );
  AND U36721 ( .A(n37179), .B(n37180), .Z(n37178) );
  XOR U36722 ( .A(n37177), .B(n37181), .Z(n37179) );
  XNOR U36723 ( .A(n37182), .B(n37183), .Z(n37176) );
  NOR U36724 ( .A(n37184), .B(n37185), .Z(n37183) );
  XNOR U36725 ( .A(n37182), .B(n37186), .Z(n37184) );
  XOR U36726 ( .A(n37187), .B(n37188), .Z(n37142) );
  NOR U36727 ( .A(n37189), .B(n37190), .Z(n37188) );
  XNOR U36728 ( .A(n37187), .B(n37191), .Z(n37189) );
  XNOR U36729 ( .A(n37083), .B(n37148), .Z(n37150) );
  XNOR U36730 ( .A(n37192), .B(n37193), .Z(n37083) );
  AND U36731 ( .A(n759), .B(n37194), .Z(n37193) );
  XNOR U36732 ( .A(n37195), .B(n37196), .Z(n37194) );
  AND U36733 ( .A(n37089), .B(n37092), .Z(n37148) );
  XOR U36734 ( .A(n37197), .B(n37175), .Z(n37092) );
  XNOR U36735 ( .A(p_input[2048]), .B(p_input[576]), .Z(n37175) );
  XOR U36736 ( .A(n37163), .B(n37162), .Z(n37197) );
  XNOR U36737 ( .A(n37198), .B(n37169), .Z(n37162) );
  XNOR U36738 ( .A(n37158), .B(n37157), .Z(n37169) );
  XOR U36739 ( .A(n37199), .B(n37154), .Z(n37157) );
  XNOR U36740 ( .A(n29266), .B(p_input[586]), .Z(n37154) );
  XNOR U36741 ( .A(p_input[2059]), .B(p_input[587]), .Z(n37199) );
  XOR U36742 ( .A(p_input[2060]), .B(p_input[588]), .Z(n37158) );
  XNOR U36743 ( .A(n37168), .B(n37159), .Z(n37198) );
  XNOR U36744 ( .A(n29494), .B(p_input[577]), .Z(n37159) );
  XOR U36745 ( .A(n37200), .B(n37174), .Z(n37168) );
  XNOR U36746 ( .A(p_input[2063]), .B(p_input[591]), .Z(n37174) );
  XOR U36747 ( .A(n37165), .B(n37173), .Z(n37200) );
  XOR U36748 ( .A(n37201), .B(n37170), .Z(n37173) );
  XOR U36749 ( .A(p_input[2061]), .B(p_input[589]), .Z(n37170) );
  XNOR U36750 ( .A(p_input[2062]), .B(p_input[590]), .Z(n37201) );
  XNOR U36751 ( .A(n29036), .B(p_input[585]), .Z(n37165) );
  XNOR U36752 ( .A(n37181), .B(n37180), .Z(n37163) );
  XNOR U36753 ( .A(n37202), .B(n37186), .Z(n37180) );
  XOR U36754 ( .A(p_input[2056]), .B(p_input[584]), .Z(n37186) );
  XOR U36755 ( .A(n37177), .B(n37185), .Z(n37202) );
  XOR U36756 ( .A(n37203), .B(n37182), .Z(n37185) );
  XOR U36757 ( .A(p_input[2054]), .B(p_input[582]), .Z(n37182) );
  XNOR U36758 ( .A(p_input[2055]), .B(p_input[583]), .Z(n37203) );
  XNOR U36759 ( .A(n29039), .B(p_input[578]), .Z(n37177) );
  XNOR U36760 ( .A(n37191), .B(n37190), .Z(n37181) );
  XOR U36761 ( .A(n37204), .B(n37187), .Z(n37190) );
  XOR U36762 ( .A(p_input[2051]), .B(p_input[579]), .Z(n37187) );
  XNOR U36763 ( .A(p_input[2052]), .B(p_input[580]), .Z(n37204) );
  XOR U36764 ( .A(p_input[2053]), .B(p_input[581]), .Z(n37191) );
  XNOR U36765 ( .A(n37205), .B(n37206), .Z(n37089) );
  AND U36766 ( .A(n759), .B(n37207), .Z(n37206) );
  XNOR U36767 ( .A(n37208), .B(n37209), .Z(n759) );
  AND U36768 ( .A(n37210), .B(n37211), .Z(n37209) );
  XOR U36769 ( .A(n37103), .B(n37208), .Z(n37211) );
  XNOR U36770 ( .A(n37212), .B(n37208), .Z(n37210) );
  XOR U36771 ( .A(n37213), .B(n37214), .Z(n37208) );
  AND U36772 ( .A(n37215), .B(n37216), .Z(n37214) );
  XOR U36773 ( .A(n37118), .B(n37213), .Z(n37216) );
  XOR U36774 ( .A(n37213), .B(n37119), .Z(n37215) );
  XOR U36775 ( .A(n37217), .B(n37218), .Z(n37213) );
  AND U36776 ( .A(n37219), .B(n37220), .Z(n37218) );
  XOR U36777 ( .A(n37146), .B(n37217), .Z(n37220) );
  XOR U36778 ( .A(n37217), .B(n37147), .Z(n37219) );
  XOR U36779 ( .A(n37221), .B(n37222), .Z(n37217) );
  AND U36780 ( .A(n37223), .B(n37224), .Z(n37222) );
  XOR U36781 ( .A(n37221), .B(n37195), .Z(n37224) );
  XNOR U36782 ( .A(n37225), .B(n37226), .Z(n37049) );
  AND U36783 ( .A(n763), .B(n37227), .Z(n37226) );
  XNOR U36784 ( .A(n37228), .B(n37229), .Z(n763) );
  AND U36785 ( .A(n37230), .B(n37231), .Z(n37229) );
  XOR U36786 ( .A(n37228), .B(n37059), .Z(n37231) );
  XNOR U36787 ( .A(n37228), .B(n37019), .Z(n37230) );
  XOR U36788 ( .A(n37232), .B(n37233), .Z(n37228) );
  AND U36789 ( .A(n37234), .B(n37235), .Z(n37233) );
  XOR U36790 ( .A(n37232), .B(n37027), .Z(n37234) );
  XOR U36791 ( .A(n37236), .B(n37237), .Z(n37010) );
  AND U36792 ( .A(n767), .B(n37227), .Z(n37237) );
  XNOR U36793 ( .A(n37225), .B(n37236), .Z(n37227) );
  XNOR U36794 ( .A(n37238), .B(n37239), .Z(n767) );
  AND U36795 ( .A(n37240), .B(n37241), .Z(n37239) );
  XNOR U36796 ( .A(n37242), .B(n37238), .Z(n37241) );
  IV U36797 ( .A(n37059), .Z(n37242) );
  XOR U36798 ( .A(n37212), .B(n37243), .Z(n37059) );
  AND U36799 ( .A(n770), .B(n37244), .Z(n37243) );
  XOR U36800 ( .A(n37102), .B(n37099), .Z(n37244) );
  IV U36801 ( .A(n37212), .Z(n37102) );
  XNOR U36802 ( .A(n37019), .B(n37238), .Z(n37240) );
  XOR U36803 ( .A(n37245), .B(n37246), .Z(n37019) );
  AND U36804 ( .A(n786), .B(n37247), .Z(n37246) );
  XOR U36805 ( .A(n37232), .B(n37248), .Z(n37238) );
  AND U36806 ( .A(n37249), .B(n37235), .Z(n37248) );
  XNOR U36807 ( .A(n37069), .B(n37232), .Z(n37235) );
  XOR U36808 ( .A(n37119), .B(n37250), .Z(n37069) );
  AND U36809 ( .A(n770), .B(n37251), .Z(n37250) );
  XOR U36810 ( .A(n37115), .B(n37119), .Z(n37251) );
  XNOR U36811 ( .A(n37252), .B(n37232), .Z(n37249) );
  IV U36812 ( .A(n37027), .Z(n37252) );
  XOR U36813 ( .A(n37253), .B(n37254), .Z(n37027) );
  AND U36814 ( .A(n786), .B(n37255), .Z(n37254) );
  XOR U36815 ( .A(n37256), .B(n37257), .Z(n37232) );
  AND U36816 ( .A(n37258), .B(n37259), .Z(n37257) );
  XNOR U36817 ( .A(n37079), .B(n37256), .Z(n37259) );
  XOR U36818 ( .A(n37147), .B(n37260), .Z(n37079) );
  AND U36819 ( .A(n770), .B(n37261), .Z(n37260) );
  XOR U36820 ( .A(n37143), .B(n37147), .Z(n37261) );
  XOR U36821 ( .A(n37256), .B(n37036), .Z(n37258) );
  XOR U36822 ( .A(n37262), .B(n37263), .Z(n37036) );
  AND U36823 ( .A(n786), .B(n37264), .Z(n37263) );
  XOR U36824 ( .A(n37265), .B(n37266), .Z(n37256) );
  AND U36825 ( .A(n37267), .B(n37268), .Z(n37266) );
  XNOR U36826 ( .A(n37265), .B(n37087), .Z(n37268) );
  XOR U36827 ( .A(n37196), .B(n37269), .Z(n37087) );
  AND U36828 ( .A(n770), .B(n37270), .Z(n37269) );
  XOR U36829 ( .A(n37192), .B(n37196), .Z(n37270) );
  XNOR U36830 ( .A(n37271), .B(n37265), .Z(n37267) );
  IV U36831 ( .A(n37046), .Z(n37271) );
  XOR U36832 ( .A(n37272), .B(n37273), .Z(n37046) );
  AND U36833 ( .A(n786), .B(n37274), .Z(n37273) );
  AND U36834 ( .A(n37236), .B(n37225), .Z(n37265) );
  XNOR U36835 ( .A(n37275), .B(n37276), .Z(n37225) );
  AND U36836 ( .A(n770), .B(n37207), .Z(n37276) );
  XNOR U36837 ( .A(n37205), .B(n37275), .Z(n37207) );
  XNOR U36838 ( .A(n37277), .B(n37278), .Z(n770) );
  AND U36839 ( .A(n37279), .B(n37280), .Z(n37278) );
  XNOR U36840 ( .A(n37277), .B(n37099), .Z(n37280) );
  IV U36841 ( .A(n37103), .Z(n37099) );
  XOR U36842 ( .A(n37281), .B(n37282), .Z(n37103) );
  AND U36843 ( .A(n774), .B(n37283), .Z(n37282) );
  XOR U36844 ( .A(n37284), .B(n37281), .Z(n37283) );
  XNOR U36845 ( .A(n37277), .B(n37212), .Z(n37279) );
  XOR U36846 ( .A(n37285), .B(n37286), .Z(n37212) );
  AND U36847 ( .A(n782), .B(n37247), .Z(n37286) );
  XOR U36848 ( .A(n37245), .B(n37285), .Z(n37247) );
  XOR U36849 ( .A(n37287), .B(n37288), .Z(n37277) );
  AND U36850 ( .A(n37289), .B(n37290), .Z(n37288) );
  XNOR U36851 ( .A(n37287), .B(n37115), .Z(n37290) );
  IV U36852 ( .A(n37118), .Z(n37115) );
  XOR U36853 ( .A(n37291), .B(n37292), .Z(n37118) );
  AND U36854 ( .A(n774), .B(n37293), .Z(n37292) );
  XOR U36855 ( .A(n37294), .B(n37291), .Z(n37293) );
  XOR U36856 ( .A(n37119), .B(n37287), .Z(n37289) );
  XOR U36857 ( .A(n37295), .B(n37296), .Z(n37119) );
  AND U36858 ( .A(n782), .B(n37255), .Z(n37296) );
  XOR U36859 ( .A(n37295), .B(n37253), .Z(n37255) );
  XOR U36860 ( .A(n37297), .B(n37298), .Z(n37287) );
  AND U36861 ( .A(n37299), .B(n37300), .Z(n37298) );
  XNOR U36862 ( .A(n37297), .B(n37143), .Z(n37300) );
  IV U36863 ( .A(n37146), .Z(n37143) );
  XOR U36864 ( .A(n37301), .B(n37302), .Z(n37146) );
  AND U36865 ( .A(n774), .B(n37303), .Z(n37302) );
  XNOR U36866 ( .A(n37304), .B(n37301), .Z(n37303) );
  XOR U36867 ( .A(n37147), .B(n37297), .Z(n37299) );
  XOR U36868 ( .A(n37305), .B(n37306), .Z(n37147) );
  AND U36869 ( .A(n782), .B(n37264), .Z(n37306) );
  XOR U36870 ( .A(n37305), .B(n37262), .Z(n37264) );
  XOR U36871 ( .A(n37221), .B(n37307), .Z(n37297) );
  AND U36872 ( .A(n37223), .B(n37308), .Z(n37307) );
  XNOR U36873 ( .A(n37221), .B(n37192), .Z(n37308) );
  IV U36874 ( .A(n37195), .Z(n37192) );
  XOR U36875 ( .A(n37309), .B(n37310), .Z(n37195) );
  AND U36876 ( .A(n774), .B(n37311), .Z(n37310) );
  XOR U36877 ( .A(n37312), .B(n37309), .Z(n37311) );
  XOR U36878 ( .A(n37196), .B(n37221), .Z(n37223) );
  XOR U36879 ( .A(n37313), .B(n37314), .Z(n37196) );
  AND U36880 ( .A(n782), .B(n37274), .Z(n37314) );
  XOR U36881 ( .A(n37313), .B(n37272), .Z(n37274) );
  AND U36882 ( .A(n37275), .B(n37205), .Z(n37221) );
  XNOR U36883 ( .A(n37315), .B(n37316), .Z(n37205) );
  AND U36884 ( .A(n774), .B(n37317), .Z(n37316) );
  XNOR U36885 ( .A(n37318), .B(n37315), .Z(n37317) );
  XNOR U36886 ( .A(n37319), .B(n37320), .Z(n774) );
  AND U36887 ( .A(n37321), .B(n37322), .Z(n37320) );
  XOR U36888 ( .A(n37284), .B(n37319), .Z(n37322) );
  AND U36889 ( .A(n37323), .B(n37324), .Z(n37284) );
  XNOR U36890 ( .A(n37281), .B(n37319), .Z(n37321) );
  XNOR U36891 ( .A(n37325), .B(n37326), .Z(n37281) );
  AND U36892 ( .A(n778), .B(n37327), .Z(n37326) );
  XNOR U36893 ( .A(n37328), .B(n37329), .Z(n37327) );
  XOR U36894 ( .A(n37330), .B(n37331), .Z(n37319) );
  AND U36895 ( .A(n37332), .B(n37333), .Z(n37331) );
  XNOR U36896 ( .A(n37330), .B(n37323), .Z(n37333) );
  IV U36897 ( .A(n37294), .Z(n37323) );
  XOR U36898 ( .A(n37334), .B(n37335), .Z(n37294) );
  XOR U36899 ( .A(n37336), .B(n37324), .Z(n37335) );
  AND U36900 ( .A(n37304), .B(n37337), .Z(n37324) );
  AND U36901 ( .A(n37338), .B(n37339), .Z(n37336) );
  XOR U36902 ( .A(n37340), .B(n37334), .Z(n37338) );
  XNOR U36903 ( .A(n37291), .B(n37330), .Z(n37332) );
  XNOR U36904 ( .A(n37341), .B(n37342), .Z(n37291) );
  AND U36905 ( .A(n778), .B(n37343), .Z(n37342) );
  XNOR U36906 ( .A(n37344), .B(n37345), .Z(n37343) );
  XOR U36907 ( .A(n37346), .B(n37347), .Z(n37330) );
  AND U36908 ( .A(n37348), .B(n37349), .Z(n37347) );
  XNOR U36909 ( .A(n37346), .B(n37304), .Z(n37349) );
  XOR U36910 ( .A(n37350), .B(n37339), .Z(n37304) );
  XNOR U36911 ( .A(n37351), .B(n37334), .Z(n37339) );
  XOR U36912 ( .A(n37352), .B(n37353), .Z(n37334) );
  AND U36913 ( .A(n37354), .B(n37355), .Z(n37353) );
  XOR U36914 ( .A(n37356), .B(n37352), .Z(n37354) );
  XNOR U36915 ( .A(n37357), .B(n37358), .Z(n37351) );
  AND U36916 ( .A(n37359), .B(n37360), .Z(n37358) );
  XOR U36917 ( .A(n37357), .B(n37361), .Z(n37359) );
  XNOR U36918 ( .A(n37340), .B(n37337), .Z(n37350) );
  AND U36919 ( .A(n37362), .B(n37363), .Z(n37337) );
  XOR U36920 ( .A(n37364), .B(n37365), .Z(n37340) );
  AND U36921 ( .A(n37366), .B(n37367), .Z(n37365) );
  XOR U36922 ( .A(n37364), .B(n37368), .Z(n37366) );
  XNOR U36923 ( .A(n37301), .B(n37346), .Z(n37348) );
  XNOR U36924 ( .A(n37369), .B(n37370), .Z(n37301) );
  AND U36925 ( .A(n778), .B(n37371), .Z(n37370) );
  XNOR U36926 ( .A(n37372), .B(n37373), .Z(n37371) );
  XOR U36927 ( .A(n37374), .B(n37375), .Z(n37346) );
  AND U36928 ( .A(n37376), .B(n37377), .Z(n37375) );
  XNOR U36929 ( .A(n37374), .B(n37362), .Z(n37377) );
  IV U36930 ( .A(n37312), .Z(n37362) );
  XNOR U36931 ( .A(n37378), .B(n37355), .Z(n37312) );
  XNOR U36932 ( .A(n37379), .B(n37361), .Z(n37355) );
  XOR U36933 ( .A(n37380), .B(n37381), .Z(n37361) );
  NOR U36934 ( .A(n37382), .B(n37383), .Z(n37381) );
  XNOR U36935 ( .A(n37380), .B(n37384), .Z(n37382) );
  XNOR U36936 ( .A(n37360), .B(n37352), .Z(n37379) );
  XOR U36937 ( .A(n37385), .B(n37386), .Z(n37352) );
  AND U36938 ( .A(n37387), .B(n37388), .Z(n37386) );
  XNOR U36939 ( .A(n37385), .B(n37389), .Z(n37387) );
  XNOR U36940 ( .A(n37390), .B(n37357), .Z(n37360) );
  XOR U36941 ( .A(n37391), .B(n37392), .Z(n37357) );
  AND U36942 ( .A(n37393), .B(n37394), .Z(n37392) );
  XOR U36943 ( .A(n37391), .B(n37395), .Z(n37393) );
  XNOR U36944 ( .A(n37396), .B(n37397), .Z(n37390) );
  NOR U36945 ( .A(n37398), .B(n37399), .Z(n37397) );
  XOR U36946 ( .A(n37396), .B(n37400), .Z(n37398) );
  XNOR U36947 ( .A(n37356), .B(n37363), .Z(n37378) );
  NOR U36948 ( .A(n37318), .B(n37401), .Z(n37363) );
  XOR U36949 ( .A(n37368), .B(n37367), .Z(n37356) );
  XNOR U36950 ( .A(n37402), .B(n37364), .Z(n37367) );
  XOR U36951 ( .A(n37403), .B(n37404), .Z(n37364) );
  AND U36952 ( .A(n37405), .B(n37406), .Z(n37404) );
  XOR U36953 ( .A(n37403), .B(n37407), .Z(n37405) );
  XNOR U36954 ( .A(n37408), .B(n37409), .Z(n37402) );
  NOR U36955 ( .A(n37410), .B(n37411), .Z(n37409) );
  XNOR U36956 ( .A(n37408), .B(n37412), .Z(n37410) );
  XOR U36957 ( .A(n37413), .B(n37414), .Z(n37368) );
  NOR U36958 ( .A(n37415), .B(n37416), .Z(n37414) );
  XNOR U36959 ( .A(n37413), .B(n37417), .Z(n37415) );
  XNOR U36960 ( .A(n37309), .B(n37374), .Z(n37376) );
  XNOR U36961 ( .A(n37418), .B(n37419), .Z(n37309) );
  AND U36962 ( .A(n778), .B(n37420), .Z(n37419) );
  XNOR U36963 ( .A(n37421), .B(n37422), .Z(n37420) );
  AND U36964 ( .A(n37315), .B(n37318), .Z(n37374) );
  XOR U36965 ( .A(n37423), .B(n37401), .Z(n37318) );
  XNOR U36966 ( .A(p_input[2048]), .B(p_input[592]), .Z(n37401) );
  XOR U36967 ( .A(n37389), .B(n37388), .Z(n37423) );
  XNOR U36968 ( .A(n37424), .B(n37395), .Z(n37388) );
  XNOR U36969 ( .A(n37384), .B(n37383), .Z(n37395) );
  XOR U36970 ( .A(n37425), .B(n37380), .Z(n37383) );
  XNOR U36971 ( .A(n29266), .B(p_input[602]), .Z(n37380) );
  XNOR U36972 ( .A(p_input[2059]), .B(p_input[603]), .Z(n37425) );
  XOR U36973 ( .A(p_input[2060]), .B(p_input[604]), .Z(n37384) );
  XNOR U36974 ( .A(n37394), .B(n37385), .Z(n37424) );
  XNOR U36975 ( .A(n29494), .B(p_input[593]), .Z(n37385) );
  XOR U36976 ( .A(n37426), .B(n37400), .Z(n37394) );
  XNOR U36977 ( .A(p_input[2063]), .B(p_input[607]), .Z(n37400) );
  XOR U36978 ( .A(n37391), .B(n37399), .Z(n37426) );
  XOR U36979 ( .A(n37427), .B(n37396), .Z(n37399) );
  XOR U36980 ( .A(p_input[2061]), .B(p_input[605]), .Z(n37396) );
  XNOR U36981 ( .A(p_input[2062]), .B(p_input[606]), .Z(n37427) );
  XNOR U36982 ( .A(n29036), .B(p_input[601]), .Z(n37391) );
  XNOR U36983 ( .A(n37407), .B(n37406), .Z(n37389) );
  XNOR U36984 ( .A(n37428), .B(n37412), .Z(n37406) );
  XOR U36985 ( .A(p_input[2056]), .B(p_input[600]), .Z(n37412) );
  XOR U36986 ( .A(n37403), .B(n37411), .Z(n37428) );
  XOR U36987 ( .A(n37429), .B(n37408), .Z(n37411) );
  XOR U36988 ( .A(p_input[2054]), .B(p_input[598]), .Z(n37408) );
  XNOR U36989 ( .A(p_input[2055]), .B(p_input[599]), .Z(n37429) );
  XNOR U36990 ( .A(n29039), .B(p_input[594]), .Z(n37403) );
  XNOR U36991 ( .A(n37417), .B(n37416), .Z(n37407) );
  XOR U36992 ( .A(n37430), .B(n37413), .Z(n37416) );
  XOR U36993 ( .A(p_input[2051]), .B(p_input[595]), .Z(n37413) );
  XNOR U36994 ( .A(p_input[2052]), .B(p_input[596]), .Z(n37430) );
  XOR U36995 ( .A(p_input[2053]), .B(p_input[597]), .Z(n37417) );
  XNOR U36996 ( .A(n37431), .B(n37432), .Z(n37315) );
  AND U36997 ( .A(n778), .B(n37433), .Z(n37432) );
  XNOR U36998 ( .A(n37434), .B(n37435), .Z(n778) );
  AND U36999 ( .A(n37436), .B(n37437), .Z(n37435) );
  XOR U37000 ( .A(n37329), .B(n37434), .Z(n37437) );
  XNOR U37001 ( .A(n37438), .B(n37434), .Z(n37436) );
  XOR U37002 ( .A(n37439), .B(n37440), .Z(n37434) );
  AND U37003 ( .A(n37441), .B(n37442), .Z(n37440) );
  XOR U37004 ( .A(n37344), .B(n37439), .Z(n37442) );
  XOR U37005 ( .A(n37439), .B(n37345), .Z(n37441) );
  XOR U37006 ( .A(n37443), .B(n37444), .Z(n37439) );
  AND U37007 ( .A(n37445), .B(n37446), .Z(n37444) );
  XOR U37008 ( .A(n37372), .B(n37443), .Z(n37446) );
  XOR U37009 ( .A(n37443), .B(n37373), .Z(n37445) );
  XOR U37010 ( .A(n37447), .B(n37448), .Z(n37443) );
  AND U37011 ( .A(n37449), .B(n37450), .Z(n37448) );
  XOR U37012 ( .A(n37447), .B(n37421), .Z(n37450) );
  XNOR U37013 ( .A(n37451), .B(n37452), .Z(n37275) );
  AND U37014 ( .A(n782), .B(n37453), .Z(n37452) );
  XNOR U37015 ( .A(n37454), .B(n37455), .Z(n782) );
  AND U37016 ( .A(n37456), .B(n37457), .Z(n37455) );
  XOR U37017 ( .A(n37454), .B(n37285), .Z(n37457) );
  XNOR U37018 ( .A(n37454), .B(n37245), .Z(n37456) );
  XOR U37019 ( .A(n37458), .B(n37459), .Z(n37454) );
  AND U37020 ( .A(n37460), .B(n37461), .Z(n37459) );
  XOR U37021 ( .A(n37458), .B(n37253), .Z(n37460) );
  XOR U37022 ( .A(n37462), .B(n37463), .Z(n37236) );
  AND U37023 ( .A(n786), .B(n37453), .Z(n37463) );
  XNOR U37024 ( .A(n37451), .B(n37462), .Z(n37453) );
  XNOR U37025 ( .A(n37464), .B(n37465), .Z(n786) );
  AND U37026 ( .A(n37466), .B(n37467), .Z(n37465) );
  XNOR U37027 ( .A(n37468), .B(n37464), .Z(n37467) );
  IV U37028 ( .A(n37285), .Z(n37468) );
  XOR U37029 ( .A(n37438), .B(n37469), .Z(n37285) );
  AND U37030 ( .A(n789), .B(n37470), .Z(n37469) );
  XOR U37031 ( .A(n37328), .B(n37325), .Z(n37470) );
  IV U37032 ( .A(n37438), .Z(n37328) );
  XNOR U37033 ( .A(n37245), .B(n37464), .Z(n37466) );
  XOR U37034 ( .A(n37471), .B(n37472), .Z(n37245) );
  AND U37035 ( .A(n805), .B(n37473), .Z(n37472) );
  XOR U37036 ( .A(n37458), .B(n37474), .Z(n37464) );
  AND U37037 ( .A(n37475), .B(n37461), .Z(n37474) );
  XNOR U37038 ( .A(n37295), .B(n37458), .Z(n37461) );
  XOR U37039 ( .A(n37345), .B(n37476), .Z(n37295) );
  AND U37040 ( .A(n789), .B(n37477), .Z(n37476) );
  XOR U37041 ( .A(n37341), .B(n37345), .Z(n37477) );
  XNOR U37042 ( .A(n37478), .B(n37458), .Z(n37475) );
  IV U37043 ( .A(n37253), .Z(n37478) );
  XOR U37044 ( .A(n37479), .B(n37480), .Z(n37253) );
  AND U37045 ( .A(n805), .B(n37481), .Z(n37480) );
  XOR U37046 ( .A(n37482), .B(n37483), .Z(n37458) );
  AND U37047 ( .A(n37484), .B(n37485), .Z(n37483) );
  XNOR U37048 ( .A(n37305), .B(n37482), .Z(n37485) );
  XOR U37049 ( .A(n37373), .B(n37486), .Z(n37305) );
  AND U37050 ( .A(n789), .B(n37487), .Z(n37486) );
  XOR U37051 ( .A(n37369), .B(n37373), .Z(n37487) );
  XOR U37052 ( .A(n37482), .B(n37262), .Z(n37484) );
  XOR U37053 ( .A(n37488), .B(n37489), .Z(n37262) );
  AND U37054 ( .A(n805), .B(n37490), .Z(n37489) );
  XOR U37055 ( .A(n37491), .B(n37492), .Z(n37482) );
  AND U37056 ( .A(n37493), .B(n37494), .Z(n37492) );
  XNOR U37057 ( .A(n37491), .B(n37313), .Z(n37494) );
  XOR U37058 ( .A(n37422), .B(n37495), .Z(n37313) );
  AND U37059 ( .A(n789), .B(n37496), .Z(n37495) );
  XOR U37060 ( .A(n37418), .B(n37422), .Z(n37496) );
  XNOR U37061 ( .A(n37497), .B(n37491), .Z(n37493) );
  IV U37062 ( .A(n37272), .Z(n37497) );
  XOR U37063 ( .A(n37498), .B(n37499), .Z(n37272) );
  AND U37064 ( .A(n805), .B(n37500), .Z(n37499) );
  AND U37065 ( .A(n37462), .B(n37451), .Z(n37491) );
  XNOR U37066 ( .A(n37501), .B(n37502), .Z(n37451) );
  AND U37067 ( .A(n789), .B(n37433), .Z(n37502) );
  XNOR U37068 ( .A(n37431), .B(n37501), .Z(n37433) );
  XNOR U37069 ( .A(n37503), .B(n37504), .Z(n789) );
  AND U37070 ( .A(n37505), .B(n37506), .Z(n37504) );
  XNOR U37071 ( .A(n37503), .B(n37325), .Z(n37506) );
  IV U37072 ( .A(n37329), .Z(n37325) );
  XOR U37073 ( .A(n37507), .B(n37508), .Z(n37329) );
  AND U37074 ( .A(n793), .B(n37509), .Z(n37508) );
  XOR U37075 ( .A(n37510), .B(n37507), .Z(n37509) );
  XNOR U37076 ( .A(n37503), .B(n37438), .Z(n37505) );
  XOR U37077 ( .A(n37511), .B(n37512), .Z(n37438) );
  AND U37078 ( .A(n801), .B(n37473), .Z(n37512) );
  XOR U37079 ( .A(n37471), .B(n37511), .Z(n37473) );
  XOR U37080 ( .A(n37513), .B(n37514), .Z(n37503) );
  AND U37081 ( .A(n37515), .B(n37516), .Z(n37514) );
  XNOR U37082 ( .A(n37513), .B(n37341), .Z(n37516) );
  IV U37083 ( .A(n37344), .Z(n37341) );
  XOR U37084 ( .A(n37517), .B(n37518), .Z(n37344) );
  AND U37085 ( .A(n793), .B(n37519), .Z(n37518) );
  XOR U37086 ( .A(n37520), .B(n37517), .Z(n37519) );
  XOR U37087 ( .A(n37345), .B(n37513), .Z(n37515) );
  XOR U37088 ( .A(n37521), .B(n37522), .Z(n37345) );
  AND U37089 ( .A(n801), .B(n37481), .Z(n37522) );
  XOR U37090 ( .A(n37521), .B(n37479), .Z(n37481) );
  XOR U37091 ( .A(n37523), .B(n37524), .Z(n37513) );
  AND U37092 ( .A(n37525), .B(n37526), .Z(n37524) );
  XNOR U37093 ( .A(n37523), .B(n37369), .Z(n37526) );
  IV U37094 ( .A(n37372), .Z(n37369) );
  XOR U37095 ( .A(n37527), .B(n37528), .Z(n37372) );
  AND U37096 ( .A(n793), .B(n37529), .Z(n37528) );
  XNOR U37097 ( .A(n37530), .B(n37527), .Z(n37529) );
  XOR U37098 ( .A(n37373), .B(n37523), .Z(n37525) );
  XOR U37099 ( .A(n37531), .B(n37532), .Z(n37373) );
  AND U37100 ( .A(n801), .B(n37490), .Z(n37532) );
  XOR U37101 ( .A(n37531), .B(n37488), .Z(n37490) );
  XOR U37102 ( .A(n37447), .B(n37533), .Z(n37523) );
  AND U37103 ( .A(n37449), .B(n37534), .Z(n37533) );
  XNOR U37104 ( .A(n37447), .B(n37418), .Z(n37534) );
  IV U37105 ( .A(n37421), .Z(n37418) );
  XOR U37106 ( .A(n37535), .B(n37536), .Z(n37421) );
  AND U37107 ( .A(n793), .B(n37537), .Z(n37536) );
  XOR U37108 ( .A(n37538), .B(n37535), .Z(n37537) );
  XOR U37109 ( .A(n37422), .B(n37447), .Z(n37449) );
  XOR U37110 ( .A(n37539), .B(n37540), .Z(n37422) );
  AND U37111 ( .A(n801), .B(n37500), .Z(n37540) );
  XOR U37112 ( .A(n37539), .B(n37498), .Z(n37500) );
  AND U37113 ( .A(n37501), .B(n37431), .Z(n37447) );
  XNOR U37114 ( .A(n37541), .B(n37542), .Z(n37431) );
  AND U37115 ( .A(n793), .B(n37543), .Z(n37542) );
  XNOR U37116 ( .A(n37544), .B(n37541), .Z(n37543) );
  XNOR U37117 ( .A(n37545), .B(n37546), .Z(n793) );
  AND U37118 ( .A(n37547), .B(n37548), .Z(n37546) );
  XOR U37119 ( .A(n37510), .B(n37545), .Z(n37548) );
  AND U37120 ( .A(n37549), .B(n37550), .Z(n37510) );
  XNOR U37121 ( .A(n37507), .B(n37545), .Z(n37547) );
  XNOR U37122 ( .A(n37551), .B(n37552), .Z(n37507) );
  AND U37123 ( .A(n797), .B(n37553), .Z(n37552) );
  XNOR U37124 ( .A(n37554), .B(n37555), .Z(n37553) );
  XOR U37125 ( .A(n37556), .B(n37557), .Z(n37545) );
  AND U37126 ( .A(n37558), .B(n37559), .Z(n37557) );
  XNOR U37127 ( .A(n37556), .B(n37549), .Z(n37559) );
  IV U37128 ( .A(n37520), .Z(n37549) );
  XOR U37129 ( .A(n37560), .B(n37561), .Z(n37520) );
  XOR U37130 ( .A(n37562), .B(n37550), .Z(n37561) );
  AND U37131 ( .A(n37530), .B(n37563), .Z(n37550) );
  AND U37132 ( .A(n37564), .B(n37565), .Z(n37562) );
  XOR U37133 ( .A(n37566), .B(n37560), .Z(n37564) );
  XNOR U37134 ( .A(n37517), .B(n37556), .Z(n37558) );
  XNOR U37135 ( .A(n37567), .B(n37568), .Z(n37517) );
  AND U37136 ( .A(n797), .B(n37569), .Z(n37568) );
  XNOR U37137 ( .A(n37570), .B(n37571), .Z(n37569) );
  XOR U37138 ( .A(n37572), .B(n37573), .Z(n37556) );
  AND U37139 ( .A(n37574), .B(n37575), .Z(n37573) );
  XNOR U37140 ( .A(n37572), .B(n37530), .Z(n37575) );
  XOR U37141 ( .A(n37576), .B(n37565), .Z(n37530) );
  XNOR U37142 ( .A(n37577), .B(n37560), .Z(n37565) );
  XOR U37143 ( .A(n37578), .B(n37579), .Z(n37560) );
  AND U37144 ( .A(n37580), .B(n37581), .Z(n37579) );
  XOR U37145 ( .A(n37582), .B(n37578), .Z(n37580) );
  XNOR U37146 ( .A(n37583), .B(n37584), .Z(n37577) );
  AND U37147 ( .A(n37585), .B(n37586), .Z(n37584) );
  XOR U37148 ( .A(n37583), .B(n37587), .Z(n37585) );
  XNOR U37149 ( .A(n37566), .B(n37563), .Z(n37576) );
  AND U37150 ( .A(n37588), .B(n37589), .Z(n37563) );
  XOR U37151 ( .A(n37590), .B(n37591), .Z(n37566) );
  AND U37152 ( .A(n37592), .B(n37593), .Z(n37591) );
  XOR U37153 ( .A(n37590), .B(n37594), .Z(n37592) );
  XNOR U37154 ( .A(n37527), .B(n37572), .Z(n37574) );
  XNOR U37155 ( .A(n37595), .B(n37596), .Z(n37527) );
  AND U37156 ( .A(n797), .B(n37597), .Z(n37596) );
  XNOR U37157 ( .A(n37598), .B(n37599), .Z(n37597) );
  XOR U37158 ( .A(n37600), .B(n37601), .Z(n37572) );
  AND U37159 ( .A(n37602), .B(n37603), .Z(n37601) );
  XNOR U37160 ( .A(n37600), .B(n37588), .Z(n37603) );
  IV U37161 ( .A(n37538), .Z(n37588) );
  XNOR U37162 ( .A(n37604), .B(n37581), .Z(n37538) );
  XNOR U37163 ( .A(n37605), .B(n37587), .Z(n37581) );
  XOR U37164 ( .A(n37606), .B(n37607), .Z(n37587) );
  NOR U37165 ( .A(n37608), .B(n37609), .Z(n37607) );
  XNOR U37166 ( .A(n37606), .B(n37610), .Z(n37608) );
  XNOR U37167 ( .A(n37586), .B(n37578), .Z(n37605) );
  XOR U37168 ( .A(n37611), .B(n37612), .Z(n37578) );
  AND U37169 ( .A(n37613), .B(n37614), .Z(n37612) );
  XNOR U37170 ( .A(n37611), .B(n37615), .Z(n37613) );
  XNOR U37171 ( .A(n37616), .B(n37583), .Z(n37586) );
  XOR U37172 ( .A(n37617), .B(n37618), .Z(n37583) );
  AND U37173 ( .A(n37619), .B(n37620), .Z(n37618) );
  XOR U37174 ( .A(n37617), .B(n37621), .Z(n37619) );
  XNOR U37175 ( .A(n37622), .B(n37623), .Z(n37616) );
  NOR U37176 ( .A(n37624), .B(n37625), .Z(n37623) );
  XOR U37177 ( .A(n37622), .B(n37626), .Z(n37624) );
  XNOR U37178 ( .A(n37582), .B(n37589), .Z(n37604) );
  NOR U37179 ( .A(n37544), .B(n37627), .Z(n37589) );
  XOR U37180 ( .A(n37594), .B(n37593), .Z(n37582) );
  XNOR U37181 ( .A(n37628), .B(n37590), .Z(n37593) );
  XOR U37182 ( .A(n37629), .B(n37630), .Z(n37590) );
  AND U37183 ( .A(n37631), .B(n37632), .Z(n37630) );
  XOR U37184 ( .A(n37629), .B(n37633), .Z(n37631) );
  XNOR U37185 ( .A(n37634), .B(n37635), .Z(n37628) );
  NOR U37186 ( .A(n37636), .B(n37637), .Z(n37635) );
  XNOR U37187 ( .A(n37634), .B(n37638), .Z(n37636) );
  XOR U37188 ( .A(n37639), .B(n37640), .Z(n37594) );
  NOR U37189 ( .A(n37641), .B(n37642), .Z(n37640) );
  XNOR U37190 ( .A(n37639), .B(n37643), .Z(n37641) );
  XNOR U37191 ( .A(n37535), .B(n37600), .Z(n37602) );
  XNOR U37192 ( .A(n37644), .B(n37645), .Z(n37535) );
  AND U37193 ( .A(n797), .B(n37646), .Z(n37645) );
  XNOR U37194 ( .A(n37647), .B(n37648), .Z(n37646) );
  AND U37195 ( .A(n37541), .B(n37544), .Z(n37600) );
  XOR U37196 ( .A(n37649), .B(n37627), .Z(n37544) );
  XNOR U37197 ( .A(p_input[2048]), .B(p_input[608]), .Z(n37627) );
  XOR U37198 ( .A(n37615), .B(n37614), .Z(n37649) );
  XNOR U37199 ( .A(n37650), .B(n37621), .Z(n37614) );
  XNOR U37200 ( .A(n37610), .B(n37609), .Z(n37621) );
  XOR U37201 ( .A(n37651), .B(n37606), .Z(n37609) );
  XNOR U37202 ( .A(n29266), .B(p_input[618]), .Z(n37606) );
  XNOR U37203 ( .A(p_input[2059]), .B(p_input[619]), .Z(n37651) );
  XOR U37204 ( .A(p_input[2060]), .B(p_input[620]), .Z(n37610) );
  XNOR U37205 ( .A(n37620), .B(n37611), .Z(n37650) );
  XNOR U37206 ( .A(n29494), .B(p_input[609]), .Z(n37611) );
  XOR U37207 ( .A(n37652), .B(n37626), .Z(n37620) );
  XNOR U37208 ( .A(p_input[2063]), .B(p_input[623]), .Z(n37626) );
  XOR U37209 ( .A(n37617), .B(n37625), .Z(n37652) );
  XOR U37210 ( .A(n37653), .B(n37622), .Z(n37625) );
  XOR U37211 ( .A(p_input[2061]), .B(p_input[621]), .Z(n37622) );
  XNOR U37212 ( .A(p_input[2062]), .B(p_input[622]), .Z(n37653) );
  XNOR U37213 ( .A(n29036), .B(p_input[617]), .Z(n37617) );
  XNOR U37214 ( .A(n37633), .B(n37632), .Z(n37615) );
  XNOR U37215 ( .A(n37654), .B(n37638), .Z(n37632) );
  XOR U37216 ( .A(p_input[2056]), .B(p_input[616]), .Z(n37638) );
  XOR U37217 ( .A(n37629), .B(n37637), .Z(n37654) );
  XOR U37218 ( .A(n37655), .B(n37634), .Z(n37637) );
  XOR U37219 ( .A(p_input[2054]), .B(p_input[614]), .Z(n37634) );
  XNOR U37220 ( .A(p_input[2055]), .B(p_input[615]), .Z(n37655) );
  XNOR U37221 ( .A(n29039), .B(p_input[610]), .Z(n37629) );
  XNOR U37222 ( .A(n37643), .B(n37642), .Z(n37633) );
  XOR U37223 ( .A(n37656), .B(n37639), .Z(n37642) );
  XOR U37224 ( .A(p_input[2051]), .B(p_input[611]), .Z(n37639) );
  XNOR U37225 ( .A(p_input[2052]), .B(p_input[612]), .Z(n37656) );
  XOR U37226 ( .A(p_input[2053]), .B(p_input[613]), .Z(n37643) );
  XNOR U37227 ( .A(n37657), .B(n37658), .Z(n37541) );
  AND U37228 ( .A(n797), .B(n37659), .Z(n37658) );
  XNOR U37229 ( .A(n37660), .B(n37661), .Z(n797) );
  AND U37230 ( .A(n37662), .B(n37663), .Z(n37661) );
  XOR U37231 ( .A(n37555), .B(n37660), .Z(n37663) );
  XNOR U37232 ( .A(n37664), .B(n37660), .Z(n37662) );
  XOR U37233 ( .A(n37665), .B(n37666), .Z(n37660) );
  AND U37234 ( .A(n37667), .B(n37668), .Z(n37666) );
  XOR U37235 ( .A(n37570), .B(n37665), .Z(n37668) );
  XOR U37236 ( .A(n37665), .B(n37571), .Z(n37667) );
  XOR U37237 ( .A(n37669), .B(n37670), .Z(n37665) );
  AND U37238 ( .A(n37671), .B(n37672), .Z(n37670) );
  XOR U37239 ( .A(n37598), .B(n37669), .Z(n37672) );
  XOR U37240 ( .A(n37669), .B(n37599), .Z(n37671) );
  XOR U37241 ( .A(n37673), .B(n37674), .Z(n37669) );
  AND U37242 ( .A(n37675), .B(n37676), .Z(n37674) );
  XOR U37243 ( .A(n37673), .B(n37647), .Z(n37676) );
  XNOR U37244 ( .A(n37677), .B(n37678), .Z(n37501) );
  AND U37245 ( .A(n801), .B(n37679), .Z(n37678) );
  XNOR U37246 ( .A(n37680), .B(n37681), .Z(n801) );
  AND U37247 ( .A(n37682), .B(n37683), .Z(n37681) );
  XOR U37248 ( .A(n37680), .B(n37511), .Z(n37683) );
  XNOR U37249 ( .A(n37680), .B(n37471), .Z(n37682) );
  XOR U37250 ( .A(n37684), .B(n37685), .Z(n37680) );
  AND U37251 ( .A(n37686), .B(n37687), .Z(n37685) );
  XOR U37252 ( .A(n37684), .B(n37479), .Z(n37686) );
  XOR U37253 ( .A(n37688), .B(n37689), .Z(n37462) );
  AND U37254 ( .A(n805), .B(n37679), .Z(n37689) );
  XNOR U37255 ( .A(n37677), .B(n37688), .Z(n37679) );
  XNOR U37256 ( .A(n37690), .B(n37691), .Z(n805) );
  AND U37257 ( .A(n37692), .B(n37693), .Z(n37691) );
  XNOR U37258 ( .A(n37694), .B(n37690), .Z(n37693) );
  IV U37259 ( .A(n37511), .Z(n37694) );
  XOR U37260 ( .A(n37664), .B(n37695), .Z(n37511) );
  AND U37261 ( .A(n808), .B(n37696), .Z(n37695) );
  XOR U37262 ( .A(n37554), .B(n37551), .Z(n37696) );
  IV U37263 ( .A(n37664), .Z(n37554) );
  XNOR U37264 ( .A(n37471), .B(n37690), .Z(n37692) );
  XOR U37265 ( .A(n37697), .B(n37698), .Z(n37471) );
  AND U37266 ( .A(n824), .B(n37699), .Z(n37698) );
  XOR U37267 ( .A(n37684), .B(n37700), .Z(n37690) );
  AND U37268 ( .A(n37701), .B(n37687), .Z(n37700) );
  XNOR U37269 ( .A(n37521), .B(n37684), .Z(n37687) );
  XOR U37270 ( .A(n37571), .B(n37702), .Z(n37521) );
  AND U37271 ( .A(n808), .B(n37703), .Z(n37702) );
  XOR U37272 ( .A(n37567), .B(n37571), .Z(n37703) );
  XNOR U37273 ( .A(n37704), .B(n37684), .Z(n37701) );
  IV U37274 ( .A(n37479), .Z(n37704) );
  XOR U37275 ( .A(n37705), .B(n37706), .Z(n37479) );
  AND U37276 ( .A(n824), .B(n37707), .Z(n37706) );
  XOR U37277 ( .A(n37708), .B(n37709), .Z(n37684) );
  AND U37278 ( .A(n37710), .B(n37711), .Z(n37709) );
  XNOR U37279 ( .A(n37531), .B(n37708), .Z(n37711) );
  XOR U37280 ( .A(n37599), .B(n37712), .Z(n37531) );
  AND U37281 ( .A(n808), .B(n37713), .Z(n37712) );
  XOR U37282 ( .A(n37595), .B(n37599), .Z(n37713) );
  XOR U37283 ( .A(n37708), .B(n37488), .Z(n37710) );
  XOR U37284 ( .A(n37714), .B(n37715), .Z(n37488) );
  AND U37285 ( .A(n824), .B(n37716), .Z(n37715) );
  XOR U37286 ( .A(n37717), .B(n37718), .Z(n37708) );
  AND U37287 ( .A(n37719), .B(n37720), .Z(n37718) );
  XNOR U37288 ( .A(n37717), .B(n37539), .Z(n37720) );
  XOR U37289 ( .A(n37648), .B(n37721), .Z(n37539) );
  AND U37290 ( .A(n808), .B(n37722), .Z(n37721) );
  XOR U37291 ( .A(n37644), .B(n37648), .Z(n37722) );
  XNOR U37292 ( .A(n37723), .B(n37717), .Z(n37719) );
  IV U37293 ( .A(n37498), .Z(n37723) );
  XOR U37294 ( .A(n37724), .B(n37725), .Z(n37498) );
  AND U37295 ( .A(n824), .B(n37726), .Z(n37725) );
  AND U37296 ( .A(n37688), .B(n37677), .Z(n37717) );
  XNOR U37297 ( .A(n37727), .B(n37728), .Z(n37677) );
  AND U37298 ( .A(n808), .B(n37659), .Z(n37728) );
  XNOR U37299 ( .A(n37657), .B(n37727), .Z(n37659) );
  XNOR U37300 ( .A(n37729), .B(n37730), .Z(n808) );
  AND U37301 ( .A(n37731), .B(n37732), .Z(n37730) );
  XNOR U37302 ( .A(n37729), .B(n37551), .Z(n37732) );
  IV U37303 ( .A(n37555), .Z(n37551) );
  XOR U37304 ( .A(n37733), .B(n37734), .Z(n37555) );
  AND U37305 ( .A(n812), .B(n37735), .Z(n37734) );
  XOR U37306 ( .A(n37736), .B(n37733), .Z(n37735) );
  XNOR U37307 ( .A(n37729), .B(n37664), .Z(n37731) );
  XOR U37308 ( .A(n37737), .B(n37738), .Z(n37664) );
  AND U37309 ( .A(n820), .B(n37699), .Z(n37738) );
  XOR U37310 ( .A(n37697), .B(n37737), .Z(n37699) );
  XOR U37311 ( .A(n37739), .B(n37740), .Z(n37729) );
  AND U37312 ( .A(n37741), .B(n37742), .Z(n37740) );
  XNOR U37313 ( .A(n37739), .B(n37567), .Z(n37742) );
  IV U37314 ( .A(n37570), .Z(n37567) );
  XOR U37315 ( .A(n37743), .B(n37744), .Z(n37570) );
  AND U37316 ( .A(n812), .B(n37745), .Z(n37744) );
  XOR U37317 ( .A(n37746), .B(n37743), .Z(n37745) );
  XOR U37318 ( .A(n37571), .B(n37739), .Z(n37741) );
  XOR U37319 ( .A(n37747), .B(n37748), .Z(n37571) );
  AND U37320 ( .A(n820), .B(n37707), .Z(n37748) );
  XOR U37321 ( .A(n37747), .B(n37705), .Z(n37707) );
  XOR U37322 ( .A(n37749), .B(n37750), .Z(n37739) );
  AND U37323 ( .A(n37751), .B(n37752), .Z(n37750) );
  XNOR U37324 ( .A(n37749), .B(n37595), .Z(n37752) );
  IV U37325 ( .A(n37598), .Z(n37595) );
  XOR U37326 ( .A(n37753), .B(n37754), .Z(n37598) );
  AND U37327 ( .A(n812), .B(n37755), .Z(n37754) );
  XNOR U37328 ( .A(n37756), .B(n37753), .Z(n37755) );
  XOR U37329 ( .A(n37599), .B(n37749), .Z(n37751) );
  XOR U37330 ( .A(n37757), .B(n37758), .Z(n37599) );
  AND U37331 ( .A(n820), .B(n37716), .Z(n37758) );
  XOR U37332 ( .A(n37757), .B(n37714), .Z(n37716) );
  XOR U37333 ( .A(n37673), .B(n37759), .Z(n37749) );
  AND U37334 ( .A(n37675), .B(n37760), .Z(n37759) );
  XNOR U37335 ( .A(n37673), .B(n37644), .Z(n37760) );
  IV U37336 ( .A(n37647), .Z(n37644) );
  XOR U37337 ( .A(n37761), .B(n37762), .Z(n37647) );
  AND U37338 ( .A(n812), .B(n37763), .Z(n37762) );
  XOR U37339 ( .A(n37764), .B(n37761), .Z(n37763) );
  XOR U37340 ( .A(n37648), .B(n37673), .Z(n37675) );
  XOR U37341 ( .A(n37765), .B(n37766), .Z(n37648) );
  AND U37342 ( .A(n820), .B(n37726), .Z(n37766) );
  XOR U37343 ( .A(n37765), .B(n37724), .Z(n37726) );
  AND U37344 ( .A(n37727), .B(n37657), .Z(n37673) );
  XNOR U37345 ( .A(n37767), .B(n37768), .Z(n37657) );
  AND U37346 ( .A(n812), .B(n37769), .Z(n37768) );
  XNOR U37347 ( .A(n37770), .B(n37767), .Z(n37769) );
  XNOR U37348 ( .A(n37771), .B(n37772), .Z(n812) );
  AND U37349 ( .A(n37773), .B(n37774), .Z(n37772) );
  XOR U37350 ( .A(n37736), .B(n37771), .Z(n37774) );
  AND U37351 ( .A(n37775), .B(n37776), .Z(n37736) );
  XNOR U37352 ( .A(n37733), .B(n37771), .Z(n37773) );
  XNOR U37353 ( .A(n37777), .B(n37778), .Z(n37733) );
  AND U37354 ( .A(n816), .B(n37779), .Z(n37778) );
  XNOR U37355 ( .A(n37780), .B(n37781), .Z(n37779) );
  XOR U37356 ( .A(n37782), .B(n37783), .Z(n37771) );
  AND U37357 ( .A(n37784), .B(n37785), .Z(n37783) );
  XNOR U37358 ( .A(n37782), .B(n37775), .Z(n37785) );
  IV U37359 ( .A(n37746), .Z(n37775) );
  XOR U37360 ( .A(n37786), .B(n37787), .Z(n37746) );
  XOR U37361 ( .A(n37788), .B(n37776), .Z(n37787) );
  AND U37362 ( .A(n37756), .B(n37789), .Z(n37776) );
  AND U37363 ( .A(n37790), .B(n37791), .Z(n37788) );
  XOR U37364 ( .A(n37792), .B(n37786), .Z(n37790) );
  XNOR U37365 ( .A(n37743), .B(n37782), .Z(n37784) );
  XNOR U37366 ( .A(n37793), .B(n37794), .Z(n37743) );
  AND U37367 ( .A(n816), .B(n37795), .Z(n37794) );
  XNOR U37368 ( .A(n37796), .B(n37797), .Z(n37795) );
  XOR U37369 ( .A(n37798), .B(n37799), .Z(n37782) );
  AND U37370 ( .A(n37800), .B(n37801), .Z(n37799) );
  XNOR U37371 ( .A(n37798), .B(n37756), .Z(n37801) );
  XOR U37372 ( .A(n37802), .B(n37791), .Z(n37756) );
  XNOR U37373 ( .A(n37803), .B(n37786), .Z(n37791) );
  XOR U37374 ( .A(n37804), .B(n37805), .Z(n37786) );
  AND U37375 ( .A(n37806), .B(n37807), .Z(n37805) );
  XOR U37376 ( .A(n37808), .B(n37804), .Z(n37806) );
  XNOR U37377 ( .A(n37809), .B(n37810), .Z(n37803) );
  AND U37378 ( .A(n37811), .B(n37812), .Z(n37810) );
  XOR U37379 ( .A(n37809), .B(n37813), .Z(n37811) );
  XNOR U37380 ( .A(n37792), .B(n37789), .Z(n37802) );
  AND U37381 ( .A(n37814), .B(n37815), .Z(n37789) );
  XOR U37382 ( .A(n37816), .B(n37817), .Z(n37792) );
  AND U37383 ( .A(n37818), .B(n37819), .Z(n37817) );
  XOR U37384 ( .A(n37816), .B(n37820), .Z(n37818) );
  XNOR U37385 ( .A(n37753), .B(n37798), .Z(n37800) );
  XNOR U37386 ( .A(n37821), .B(n37822), .Z(n37753) );
  AND U37387 ( .A(n816), .B(n37823), .Z(n37822) );
  XNOR U37388 ( .A(n37824), .B(n37825), .Z(n37823) );
  XOR U37389 ( .A(n37826), .B(n37827), .Z(n37798) );
  AND U37390 ( .A(n37828), .B(n37829), .Z(n37827) );
  XNOR U37391 ( .A(n37826), .B(n37814), .Z(n37829) );
  IV U37392 ( .A(n37764), .Z(n37814) );
  XNOR U37393 ( .A(n37830), .B(n37807), .Z(n37764) );
  XNOR U37394 ( .A(n37831), .B(n37813), .Z(n37807) );
  XOR U37395 ( .A(n37832), .B(n37833), .Z(n37813) );
  NOR U37396 ( .A(n37834), .B(n37835), .Z(n37833) );
  XNOR U37397 ( .A(n37832), .B(n37836), .Z(n37834) );
  XNOR U37398 ( .A(n37812), .B(n37804), .Z(n37831) );
  XOR U37399 ( .A(n37837), .B(n37838), .Z(n37804) );
  AND U37400 ( .A(n37839), .B(n37840), .Z(n37838) );
  XNOR U37401 ( .A(n37837), .B(n37841), .Z(n37839) );
  XNOR U37402 ( .A(n37842), .B(n37809), .Z(n37812) );
  XOR U37403 ( .A(n37843), .B(n37844), .Z(n37809) );
  AND U37404 ( .A(n37845), .B(n37846), .Z(n37844) );
  XOR U37405 ( .A(n37843), .B(n37847), .Z(n37845) );
  XNOR U37406 ( .A(n37848), .B(n37849), .Z(n37842) );
  NOR U37407 ( .A(n37850), .B(n37851), .Z(n37849) );
  XOR U37408 ( .A(n37848), .B(n37852), .Z(n37850) );
  XNOR U37409 ( .A(n37808), .B(n37815), .Z(n37830) );
  NOR U37410 ( .A(n37770), .B(n37853), .Z(n37815) );
  XOR U37411 ( .A(n37820), .B(n37819), .Z(n37808) );
  XNOR U37412 ( .A(n37854), .B(n37816), .Z(n37819) );
  XOR U37413 ( .A(n37855), .B(n37856), .Z(n37816) );
  AND U37414 ( .A(n37857), .B(n37858), .Z(n37856) );
  XOR U37415 ( .A(n37855), .B(n37859), .Z(n37857) );
  XNOR U37416 ( .A(n37860), .B(n37861), .Z(n37854) );
  NOR U37417 ( .A(n37862), .B(n37863), .Z(n37861) );
  XNOR U37418 ( .A(n37860), .B(n37864), .Z(n37862) );
  XOR U37419 ( .A(n37865), .B(n37866), .Z(n37820) );
  NOR U37420 ( .A(n37867), .B(n37868), .Z(n37866) );
  XNOR U37421 ( .A(n37865), .B(n37869), .Z(n37867) );
  XNOR U37422 ( .A(n37761), .B(n37826), .Z(n37828) );
  XNOR U37423 ( .A(n37870), .B(n37871), .Z(n37761) );
  AND U37424 ( .A(n816), .B(n37872), .Z(n37871) );
  XNOR U37425 ( .A(n37873), .B(n37874), .Z(n37872) );
  AND U37426 ( .A(n37767), .B(n37770), .Z(n37826) );
  XOR U37427 ( .A(n37875), .B(n37853), .Z(n37770) );
  XNOR U37428 ( .A(p_input[2048]), .B(p_input[624]), .Z(n37853) );
  XOR U37429 ( .A(n37841), .B(n37840), .Z(n37875) );
  XNOR U37430 ( .A(n37876), .B(n37847), .Z(n37840) );
  XNOR U37431 ( .A(n37836), .B(n37835), .Z(n37847) );
  XOR U37432 ( .A(n37877), .B(n37832), .Z(n37835) );
  XNOR U37433 ( .A(n29266), .B(p_input[634]), .Z(n37832) );
  XNOR U37434 ( .A(p_input[2059]), .B(p_input[635]), .Z(n37877) );
  XOR U37435 ( .A(p_input[2060]), .B(p_input[636]), .Z(n37836) );
  XNOR U37436 ( .A(n37846), .B(n37837), .Z(n37876) );
  XNOR U37437 ( .A(n29494), .B(p_input[625]), .Z(n37837) );
  XOR U37438 ( .A(n37878), .B(n37852), .Z(n37846) );
  XNOR U37439 ( .A(p_input[2063]), .B(p_input[639]), .Z(n37852) );
  XOR U37440 ( .A(n37843), .B(n37851), .Z(n37878) );
  XOR U37441 ( .A(n37879), .B(n37848), .Z(n37851) );
  XOR U37442 ( .A(p_input[2061]), .B(p_input[637]), .Z(n37848) );
  XNOR U37443 ( .A(p_input[2062]), .B(p_input[638]), .Z(n37879) );
  XNOR U37444 ( .A(n29036), .B(p_input[633]), .Z(n37843) );
  XNOR U37445 ( .A(n37859), .B(n37858), .Z(n37841) );
  XNOR U37446 ( .A(n37880), .B(n37864), .Z(n37858) );
  XOR U37447 ( .A(p_input[2056]), .B(p_input[632]), .Z(n37864) );
  XOR U37448 ( .A(n37855), .B(n37863), .Z(n37880) );
  XOR U37449 ( .A(n37881), .B(n37860), .Z(n37863) );
  XOR U37450 ( .A(p_input[2054]), .B(p_input[630]), .Z(n37860) );
  XNOR U37451 ( .A(p_input[2055]), .B(p_input[631]), .Z(n37881) );
  XNOR U37452 ( .A(n29039), .B(p_input[626]), .Z(n37855) );
  XNOR U37453 ( .A(n37869), .B(n37868), .Z(n37859) );
  XOR U37454 ( .A(n37882), .B(n37865), .Z(n37868) );
  XOR U37455 ( .A(p_input[2051]), .B(p_input[627]), .Z(n37865) );
  XNOR U37456 ( .A(p_input[2052]), .B(p_input[628]), .Z(n37882) );
  XOR U37457 ( .A(p_input[2053]), .B(p_input[629]), .Z(n37869) );
  XNOR U37458 ( .A(n37883), .B(n37884), .Z(n37767) );
  AND U37459 ( .A(n816), .B(n37885), .Z(n37884) );
  XNOR U37460 ( .A(n37886), .B(n37887), .Z(n816) );
  AND U37461 ( .A(n37888), .B(n37889), .Z(n37887) );
  XOR U37462 ( .A(n37781), .B(n37886), .Z(n37889) );
  XNOR U37463 ( .A(n37890), .B(n37886), .Z(n37888) );
  XOR U37464 ( .A(n37891), .B(n37892), .Z(n37886) );
  AND U37465 ( .A(n37893), .B(n37894), .Z(n37892) );
  XOR U37466 ( .A(n37796), .B(n37891), .Z(n37894) );
  XOR U37467 ( .A(n37891), .B(n37797), .Z(n37893) );
  XOR U37468 ( .A(n37895), .B(n37896), .Z(n37891) );
  AND U37469 ( .A(n37897), .B(n37898), .Z(n37896) );
  XOR U37470 ( .A(n37824), .B(n37895), .Z(n37898) );
  XOR U37471 ( .A(n37895), .B(n37825), .Z(n37897) );
  XOR U37472 ( .A(n37899), .B(n37900), .Z(n37895) );
  AND U37473 ( .A(n37901), .B(n37902), .Z(n37900) );
  XOR U37474 ( .A(n37899), .B(n37873), .Z(n37902) );
  XNOR U37475 ( .A(n37903), .B(n37904), .Z(n37727) );
  AND U37476 ( .A(n820), .B(n37905), .Z(n37904) );
  XNOR U37477 ( .A(n37906), .B(n37907), .Z(n820) );
  AND U37478 ( .A(n37908), .B(n37909), .Z(n37907) );
  XOR U37479 ( .A(n37906), .B(n37737), .Z(n37909) );
  XNOR U37480 ( .A(n37906), .B(n37697), .Z(n37908) );
  XOR U37481 ( .A(n37910), .B(n37911), .Z(n37906) );
  AND U37482 ( .A(n37912), .B(n37913), .Z(n37911) );
  XOR U37483 ( .A(n37910), .B(n37705), .Z(n37912) );
  XOR U37484 ( .A(n37914), .B(n37915), .Z(n37688) );
  AND U37485 ( .A(n824), .B(n37905), .Z(n37915) );
  XNOR U37486 ( .A(n37903), .B(n37914), .Z(n37905) );
  XNOR U37487 ( .A(n37916), .B(n37917), .Z(n824) );
  AND U37488 ( .A(n37918), .B(n37919), .Z(n37917) );
  XNOR U37489 ( .A(n37920), .B(n37916), .Z(n37919) );
  IV U37490 ( .A(n37737), .Z(n37920) );
  XOR U37491 ( .A(n37890), .B(n37921), .Z(n37737) );
  AND U37492 ( .A(n827), .B(n37922), .Z(n37921) );
  XOR U37493 ( .A(n37780), .B(n37777), .Z(n37922) );
  IV U37494 ( .A(n37890), .Z(n37780) );
  XNOR U37495 ( .A(n37697), .B(n37916), .Z(n37918) );
  XOR U37496 ( .A(n37923), .B(n37924), .Z(n37697) );
  AND U37497 ( .A(n843), .B(n37925), .Z(n37924) );
  XOR U37498 ( .A(n37910), .B(n37926), .Z(n37916) );
  AND U37499 ( .A(n37927), .B(n37913), .Z(n37926) );
  XNOR U37500 ( .A(n37747), .B(n37910), .Z(n37913) );
  XOR U37501 ( .A(n37797), .B(n37928), .Z(n37747) );
  AND U37502 ( .A(n827), .B(n37929), .Z(n37928) );
  XOR U37503 ( .A(n37793), .B(n37797), .Z(n37929) );
  XNOR U37504 ( .A(n37930), .B(n37910), .Z(n37927) );
  IV U37505 ( .A(n37705), .Z(n37930) );
  XOR U37506 ( .A(n37931), .B(n37932), .Z(n37705) );
  AND U37507 ( .A(n843), .B(n37933), .Z(n37932) );
  XOR U37508 ( .A(n37934), .B(n37935), .Z(n37910) );
  AND U37509 ( .A(n37936), .B(n37937), .Z(n37935) );
  XNOR U37510 ( .A(n37757), .B(n37934), .Z(n37937) );
  XOR U37511 ( .A(n37825), .B(n37938), .Z(n37757) );
  AND U37512 ( .A(n827), .B(n37939), .Z(n37938) );
  XOR U37513 ( .A(n37821), .B(n37825), .Z(n37939) );
  XOR U37514 ( .A(n37934), .B(n37714), .Z(n37936) );
  XOR U37515 ( .A(n37940), .B(n37941), .Z(n37714) );
  AND U37516 ( .A(n843), .B(n37942), .Z(n37941) );
  XOR U37517 ( .A(n37943), .B(n37944), .Z(n37934) );
  AND U37518 ( .A(n37945), .B(n37946), .Z(n37944) );
  XNOR U37519 ( .A(n37943), .B(n37765), .Z(n37946) );
  XOR U37520 ( .A(n37874), .B(n37947), .Z(n37765) );
  AND U37521 ( .A(n827), .B(n37948), .Z(n37947) );
  XOR U37522 ( .A(n37870), .B(n37874), .Z(n37948) );
  XNOR U37523 ( .A(n37949), .B(n37943), .Z(n37945) );
  IV U37524 ( .A(n37724), .Z(n37949) );
  XOR U37525 ( .A(n37950), .B(n37951), .Z(n37724) );
  AND U37526 ( .A(n843), .B(n37952), .Z(n37951) );
  AND U37527 ( .A(n37914), .B(n37903), .Z(n37943) );
  XNOR U37528 ( .A(n37953), .B(n37954), .Z(n37903) );
  AND U37529 ( .A(n827), .B(n37885), .Z(n37954) );
  XNOR U37530 ( .A(n37883), .B(n37953), .Z(n37885) );
  XNOR U37531 ( .A(n37955), .B(n37956), .Z(n827) );
  AND U37532 ( .A(n37957), .B(n37958), .Z(n37956) );
  XNOR U37533 ( .A(n37955), .B(n37777), .Z(n37958) );
  IV U37534 ( .A(n37781), .Z(n37777) );
  XOR U37535 ( .A(n37959), .B(n37960), .Z(n37781) );
  AND U37536 ( .A(n831), .B(n37961), .Z(n37960) );
  XOR U37537 ( .A(n37962), .B(n37959), .Z(n37961) );
  XNOR U37538 ( .A(n37955), .B(n37890), .Z(n37957) );
  XOR U37539 ( .A(n37963), .B(n37964), .Z(n37890) );
  AND U37540 ( .A(n839), .B(n37925), .Z(n37964) );
  XOR U37541 ( .A(n37923), .B(n37963), .Z(n37925) );
  XOR U37542 ( .A(n37965), .B(n37966), .Z(n37955) );
  AND U37543 ( .A(n37967), .B(n37968), .Z(n37966) );
  XNOR U37544 ( .A(n37965), .B(n37793), .Z(n37968) );
  IV U37545 ( .A(n37796), .Z(n37793) );
  XOR U37546 ( .A(n37969), .B(n37970), .Z(n37796) );
  AND U37547 ( .A(n831), .B(n37971), .Z(n37970) );
  XOR U37548 ( .A(n37972), .B(n37969), .Z(n37971) );
  XOR U37549 ( .A(n37797), .B(n37965), .Z(n37967) );
  XOR U37550 ( .A(n37973), .B(n37974), .Z(n37797) );
  AND U37551 ( .A(n839), .B(n37933), .Z(n37974) );
  XOR U37552 ( .A(n37973), .B(n37931), .Z(n37933) );
  XOR U37553 ( .A(n37975), .B(n37976), .Z(n37965) );
  AND U37554 ( .A(n37977), .B(n37978), .Z(n37976) );
  XNOR U37555 ( .A(n37975), .B(n37821), .Z(n37978) );
  IV U37556 ( .A(n37824), .Z(n37821) );
  XOR U37557 ( .A(n37979), .B(n37980), .Z(n37824) );
  AND U37558 ( .A(n831), .B(n37981), .Z(n37980) );
  XNOR U37559 ( .A(n37982), .B(n37979), .Z(n37981) );
  XOR U37560 ( .A(n37825), .B(n37975), .Z(n37977) );
  XOR U37561 ( .A(n37983), .B(n37984), .Z(n37825) );
  AND U37562 ( .A(n839), .B(n37942), .Z(n37984) );
  XOR U37563 ( .A(n37983), .B(n37940), .Z(n37942) );
  XOR U37564 ( .A(n37899), .B(n37985), .Z(n37975) );
  AND U37565 ( .A(n37901), .B(n37986), .Z(n37985) );
  XNOR U37566 ( .A(n37899), .B(n37870), .Z(n37986) );
  IV U37567 ( .A(n37873), .Z(n37870) );
  XOR U37568 ( .A(n37987), .B(n37988), .Z(n37873) );
  AND U37569 ( .A(n831), .B(n37989), .Z(n37988) );
  XOR U37570 ( .A(n37990), .B(n37987), .Z(n37989) );
  XOR U37571 ( .A(n37874), .B(n37899), .Z(n37901) );
  XOR U37572 ( .A(n37991), .B(n37992), .Z(n37874) );
  AND U37573 ( .A(n839), .B(n37952), .Z(n37992) );
  XOR U37574 ( .A(n37991), .B(n37950), .Z(n37952) );
  AND U37575 ( .A(n37953), .B(n37883), .Z(n37899) );
  XNOR U37576 ( .A(n37993), .B(n37994), .Z(n37883) );
  AND U37577 ( .A(n831), .B(n37995), .Z(n37994) );
  XNOR U37578 ( .A(n37996), .B(n37993), .Z(n37995) );
  XNOR U37579 ( .A(n37997), .B(n37998), .Z(n831) );
  AND U37580 ( .A(n37999), .B(n38000), .Z(n37998) );
  XOR U37581 ( .A(n37962), .B(n37997), .Z(n38000) );
  AND U37582 ( .A(n38001), .B(n38002), .Z(n37962) );
  XNOR U37583 ( .A(n37959), .B(n37997), .Z(n37999) );
  XNOR U37584 ( .A(n38003), .B(n38004), .Z(n37959) );
  AND U37585 ( .A(n835), .B(n38005), .Z(n38004) );
  XNOR U37586 ( .A(n38006), .B(n38007), .Z(n38005) );
  XOR U37587 ( .A(n38008), .B(n38009), .Z(n37997) );
  AND U37588 ( .A(n38010), .B(n38011), .Z(n38009) );
  XNOR U37589 ( .A(n38008), .B(n38001), .Z(n38011) );
  IV U37590 ( .A(n37972), .Z(n38001) );
  XOR U37591 ( .A(n38012), .B(n38013), .Z(n37972) );
  XOR U37592 ( .A(n38014), .B(n38002), .Z(n38013) );
  AND U37593 ( .A(n37982), .B(n38015), .Z(n38002) );
  AND U37594 ( .A(n38016), .B(n38017), .Z(n38014) );
  XOR U37595 ( .A(n38018), .B(n38012), .Z(n38016) );
  XNOR U37596 ( .A(n37969), .B(n38008), .Z(n38010) );
  XNOR U37597 ( .A(n38019), .B(n38020), .Z(n37969) );
  AND U37598 ( .A(n835), .B(n38021), .Z(n38020) );
  XNOR U37599 ( .A(n38022), .B(n38023), .Z(n38021) );
  XOR U37600 ( .A(n38024), .B(n38025), .Z(n38008) );
  AND U37601 ( .A(n38026), .B(n38027), .Z(n38025) );
  XNOR U37602 ( .A(n38024), .B(n37982), .Z(n38027) );
  XOR U37603 ( .A(n38028), .B(n38017), .Z(n37982) );
  XNOR U37604 ( .A(n38029), .B(n38012), .Z(n38017) );
  XOR U37605 ( .A(n38030), .B(n38031), .Z(n38012) );
  AND U37606 ( .A(n38032), .B(n38033), .Z(n38031) );
  XOR U37607 ( .A(n38034), .B(n38030), .Z(n38032) );
  XNOR U37608 ( .A(n38035), .B(n38036), .Z(n38029) );
  AND U37609 ( .A(n38037), .B(n38038), .Z(n38036) );
  XOR U37610 ( .A(n38035), .B(n38039), .Z(n38037) );
  XNOR U37611 ( .A(n38018), .B(n38015), .Z(n38028) );
  AND U37612 ( .A(n38040), .B(n38041), .Z(n38015) );
  XOR U37613 ( .A(n38042), .B(n38043), .Z(n38018) );
  AND U37614 ( .A(n38044), .B(n38045), .Z(n38043) );
  XOR U37615 ( .A(n38042), .B(n38046), .Z(n38044) );
  XNOR U37616 ( .A(n37979), .B(n38024), .Z(n38026) );
  XNOR U37617 ( .A(n38047), .B(n38048), .Z(n37979) );
  AND U37618 ( .A(n835), .B(n38049), .Z(n38048) );
  XNOR U37619 ( .A(n38050), .B(n38051), .Z(n38049) );
  XOR U37620 ( .A(n38052), .B(n38053), .Z(n38024) );
  AND U37621 ( .A(n38054), .B(n38055), .Z(n38053) );
  XNOR U37622 ( .A(n38052), .B(n38040), .Z(n38055) );
  IV U37623 ( .A(n37990), .Z(n38040) );
  XNOR U37624 ( .A(n38056), .B(n38033), .Z(n37990) );
  XNOR U37625 ( .A(n38057), .B(n38039), .Z(n38033) );
  XOR U37626 ( .A(n38058), .B(n38059), .Z(n38039) );
  NOR U37627 ( .A(n38060), .B(n38061), .Z(n38059) );
  XNOR U37628 ( .A(n38058), .B(n38062), .Z(n38060) );
  XNOR U37629 ( .A(n38038), .B(n38030), .Z(n38057) );
  XOR U37630 ( .A(n38063), .B(n38064), .Z(n38030) );
  AND U37631 ( .A(n38065), .B(n38066), .Z(n38064) );
  XNOR U37632 ( .A(n38063), .B(n38067), .Z(n38065) );
  XNOR U37633 ( .A(n38068), .B(n38035), .Z(n38038) );
  XOR U37634 ( .A(n38069), .B(n38070), .Z(n38035) );
  AND U37635 ( .A(n38071), .B(n38072), .Z(n38070) );
  XOR U37636 ( .A(n38069), .B(n38073), .Z(n38071) );
  XNOR U37637 ( .A(n38074), .B(n38075), .Z(n38068) );
  NOR U37638 ( .A(n38076), .B(n38077), .Z(n38075) );
  XOR U37639 ( .A(n38074), .B(n38078), .Z(n38076) );
  XNOR U37640 ( .A(n38034), .B(n38041), .Z(n38056) );
  NOR U37641 ( .A(n37996), .B(n38079), .Z(n38041) );
  XOR U37642 ( .A(n38046), .B(n38045), .Z(n38034) );
  XNOR U37643 ( .A(n38080), .B(n38042), .Z(n38045) );
  XOR U37644 ( .A(n38081), .B(n38082), .Z(n38042) );
  AND U37645 ( .A(n38083), .B(n38084), .Z(n38082) );
  XOR U37646 ( .A(n38081), .B(n38085), .Z(n38083) );
  XNOR U37647 ( .A(n38086), .B(n38087), .Z(n38080) );
  NOR U37648 ( .A(n38088), .B(n38089), .Z(n38087) );
  XNOR U37649 ( .A(n38086), .B(n38090), .Z(n38088) );
  XOR U37650 ( .A(n38091), .B(n38092), .Z(n38046) );
  NOR U37651 ( .A(n38093), .B(n38094), .Z(n38092) );
  XNOR U37652 ( .A(n38091), .B(n38095), .Z(n38093) );
  XNOR U37653 ( .A(n37987), .B(n38052), .Z(n38054) );
  XNOR U37654 ( .A(n38096), .B(n38097), .Z(n37987) );
  AND U37655 ( .A(n835), .B(n38098), .Z(n38097) );
  XNOR U37656 ( .A(n38099), .B(n38100), .Z(n38098) );
  AND U37657 ( .A(n37993), .B(n37996), .Z(n38052) );
  XOR U37658 ( .A(n38101), .B(n38079), .Z(n37996) );
  XNOR U37659 ( .A(p_input[2048]), .B(p_input[640]), .Z(n38079) );
  XOR U37660 ( .A(n38067), .B(n38066), .Z(n38101) );
  XNOR U37661 ( .A(n38102), .B(n38073), .Z(n38066) );
  XNOR U37662 ( .A(n38062), .B(n38061), .Z(n38073) );
  XOR U37663 ( .A(n38103), .B(n38058), .Z(n38061) );
  XNOR U37664 ( .A(n29266), .B(p_input[650]), .Z(n38058) );
  XNOR U37665 ( .A(p_input[2059]), .B(p_input[651]), .Z(n38103) );
  XOR U37666 ( .A(p_input[2060]), .B(p_input[652]), .Z(n38062) );
  XNOR U37667 ( .A(n38072), .B(n38063), .Z(n38102) );
  XNOR U37668 ( .A(n29494), .B(p_input[641]), .Z(n38063) );
  XOR U37669 ( .A(n38104), .B(n38078), .Z(n38072) );
  XNOR U37670 ( .A(p_input[2063]), .B(p_input[655]), .Z(n38078) );
  XOR U37671 ( .A(n38069), .B(n38077), .Z(n38104) );
  XOR U37672 ( .A(n38105), .B(n38074), .Z(n38077) );
  XOR U37673 ( .A(p_input[2061]), .B(p_input[653]), .Z(n38074) );
  XNOR U37674 ( .A(p_input[2062]), .B(p_input[654]), .Z(n38105) );
  XNOR U37675 ( .A(n29036), .B(p_input[649]), .Z(n38069) );
  XNOR U37676 ( .A(n38085), .B(n38084), .Z(n38067) );
  XNOR U37677 ( .A(n38106), .B(n38090), .Z(n38084) );
  XOR U37678 ( .A(p_input[2056]), .B(p_input[648]), .Z(n38090) );
  XOR U37679 ( .A(n38081), .B(n38089), .Z(n38106) );
  XOR U37680 ( .A(n38107), .B(n38086), .Z(n38089) );
  XOR U37681 ( .A(p_input[2054]), .B(p_input[646]), .Z(n38086) );
  XNOR U37682 ( .A(p_input[2055]), .B(p_input[647]), .Z(n38107) );
  XNOR U37683 ( .A(n29039), .B(p_input[642]), .Z(n38081) );
  XNOR U37684 ( .A(n38095), .B(n38094), .Z(n38085) );
  XOR U37685 ( .A(n38108), .B(n38091), .Z(n38094) );
  XOR U37686 ( .A(p_input[2051]), .B(p_input[643]), .Z(n38091) );
  XNOR U37687 ( .A(p_input[2052]), .B(p_input[644]), .Z(n38108) );
  XOR U37688 ( .A(p_input[2053]), .B(p_input[645]), .Z(n38095) );
  XNOR U37689 ( .A(n38109), .B(n38110), .Z(n37993) );
  AND U37690 ( .A(n835), .B(n38111), .Z(n38110) );
  XNOR U37691 ( .A(n38112), .B(n38113), .Z(n835) );
  AND U37692 ( .A(n38114), .B(n38115), .Z(n38113) );
  XOR U37693 ( .A(n38007), .B(n38112), .Z(n38115) );
  XNOR U37694 ( .A(n38116), .B(n38112), .Z(n38114) );
  XOR U37695 ( .A(n38117), .B(n38118), .Z(n38112) );
  AND U37696 ( .A(n38119), .B(n38120), .Z(n38118) );
  XOR U37697 ( .A(n38022), .B(n38117), .Z(n38120) );
  XOR U37698 ( .A(n38117), .B(n38023), .Z(n38119) );
  XOR U37699 ( .A(n38121), .B(n38122), .Z(n38117) );
  AND U37700 ( .A(n38123), .B(n38124), .Z(n38122) );
  XOR U37701 ( .A(n38050), .B(n38121), .Z(n38124) );
  XOR U37702 ( .A(n38121), .B(n38051), .Z(n38123) );
  XOR U37703 ( .A(n38125), .B(n38126), .Z(n38121) );
  AND U37704 ( .A(n38127), .B(n38128), .Z(n38126) );
  XOR U37705 ( .A(n38125), .B(n38099), .Z(n38128) );
  XNOR U37706 ( .A(n38129), .B(n38130), .Z(n37953) );
  AND U37707 ( .A(n839), .B(n38131), .Z(n38130) );
  XNOR U37708 ( .A(n38132), .B(n38133), .Z(n839) );
  AND U37709 ( .A(n38134), .B(n38135), .Z(n38133) );
  XOR U37710 ( .A(n38132), .B(n37963), .Z(n38135) );
  XNOR U37711 ( .A(n38132), .B(n37923), .Z(n38134) );
  XOR U37712 ( .A(n38136), .B(n38137), .Z(n38132) );
  AND U37713 ( .A(n38138), .B(n38139), .Z(n38137) );
  XOR U37714 ( .A(n38136), .B(n37931), .Z(n38138) );
  XOR U37715 ( .A(n38140), .B(n38141), .Z(n37914) );
  AND U37716 ( .A(n843), .B(n38131), .Z(n38141) );
  XNOR U37717 ( .A(n38129), .B(n38140), .Z(n38131) );
  XNOR U37718 ( .A(n38142), .B(n38143), .Z(n843) );
  AND U37719 ( .A(n38144), .B(n38145), .Z(n38143) );
  XNOR U37720 ( .A(n38146), .B(n38142), .Z(n38145) );
  IV U37721 ( .A(n37963), .Z(n38146) );
  XOR U37722 ( .A(n38116), .B(n38147), .Z(n37963) );
  AND U37723 ( .A(n846), .B(n38148), .Z(n38147) );
  XOR U37724 ( .A(n38006), .B(n38003), .Z(n38148) );
  IV U37725 ( .A(n38116), .Z(n38006) );
  XNOR U37726 ( .A(n37923), .B(n38142), .Z(n38144) );
  XOR U37727 ( .A(n38149), .B(n38150), .Z(n37923) );
  AND U37728 ( .A(n862), .B(n38151), .Z(n38150) );
  XOR U37729 ( .A(n38136), .B(n38152), .Z(n38142) );
  AND U37730 ( .A(n38153), .B(n38139), .Z(n38152) );
  XNOR U37731 ( .A(n37973), .B(n38136), .Z(n38139) );
  XOR U37732 ( .A(n38023), .B(n38154), .Z(n37973) );
  AND U37733 ( .A(n846), .B(n38155), .Z(n38154) );
  XOR U37734 ( .A(n38019), .B(n38023), .Z(n38155) );
  XNOR U37735 ( .A(n38156), .B(n38136), .Z(n38153) );
  IV U37736 ( .A(n37931), .Z(n38156) );
  XOR U37737 ( .A(n38157), .B(n38158), .Z(n37931) );
  AND U37738 ( .A(n862), .B(n38159), .Z(n38158) );
  XOR U37739 ( .A(n38160), .B(n38161), .Z(n38136) );
  AND U37740 ( .A(n38162), .B(n38163), .Z(n38161) );
  XNOR U37741 ( .A(n37983), .B(n38160), .Z(n38163) );
  XOR U37742 ( .A(n38051), .B(n38164), .Z(n37983) );
  AND U37743 ( .A(n846), .B(n38165), .Z(n38164) );
  XOR U37744 ( .A(n38047), .B(n38051), .Z(n38165) );
  XOR U37745 ( .A(n38160), .B(n37940), .Z(n38162) );
  XOR U37746 ( .A(n38166), .B(n38167), .Z(n37940) );
  AND U37747 ( .A(n862), .B(n38168), .Z(n38167) );
  XOR U37748 ( .A(n38169), .B(n38170), .Z(n38160) );
  AND U37749 ( .A(n38171), .B(n38172), .Z(n38170) );
  XNOR U37750 ( .A(n38169), .B(n37991), .Z(n38172) );
  XOR U37751 ( .A(n38100), .B(n38173), .Z(n37991) );
  AND U37752 ( .A(n846), .B(n38174), .Z(n38173) );
  XOR U37753 ( .A(n38096), .B(n38100), .Z(n38174) );
  XNOR U37754 ( .A(n38175), .B(n38169), .Z(n38171) );
  IV U37755 ( .A(n37950), .Z(n38175) );
  XOR U37756 ( .A(n38176), .B(n38177), .Z(n37950) );
  AND U37757 ( .A(n862), .B(n38178), .Z(n38177) );
  AND U37758 ( .A(n38140), .B(n38129), .Z(n38169) );
  XNOR U37759 ( .A(n38179), .B(n38180), .Z(n38129) );
  AND U37760 ( .A(n846), .B(n38111), .Z(n38180) );
  XNOR U37761 ( .A(n38109), .B(n38179), .Z(n38111) );
  XNOR U37762 ( .A(n38181), .B(n38182), .Z(n846) );
  AND U37763 ( .A(n38183), .B(n38184), .Z(n38182) );
  XNOR U37764 ( .A(n38181), .B(n38003), .Z(n38184) );
  IV U37765 ( .A(n38007), .Z(n38003) );
  XOR U37766 ( .A(n38185), .B(n38186), .Z(n38007) );
  AND U37767 ( .A(n850), .B(n38187), .Z(n38186) );
  XOR U37768 ( .A(n38188), .B(n38185), .Z(n38187) );
  XNOR U37769 ( .A(n38181), .B(n38116), .Z(n38183) );
  XOR U37770 ( .A(n38189), .B(n38190), .Z(n38116) );
  AND U37771 ( .A(n858), .B(n38151), .Z(n38190) );
  XOR U37772 ( .A(n38149), .B(n38189), .Z(n38151) );
  XOR U37773 ( .A(n38191), .B(n38192), .Z(n38181) );
  AND U37774 ( .A(n38193), .B(n38194), .Z(n38192) );
  XNOR U37775 ( .A(n38191), .B(n38019), .Z(n38194) );
  IV U37776 ( .A(n38022), .Z(n38019) );
  XOR U37777 ( .A(n38195), .B(n38196), .Z(n38022) );
  AND U37778 ( .A(n850), .B(n38197), .Z(n38196) );
  XOR U37779 ( .A(n38198), .B(n38195), .Z(n38197) );
  XOR U37780 ( .A(n38023), .B(n38191), .Z(n38193) );
  XOR U37781 ( .A(n38199), .B(n38200), .Z(n38023) );
  AND U37782 ( .A(n858), .B(n38159), .Z(n38200) );
  XOR U37783 ( .A(n38199), .B(n38157), .Z(n38159) );
  XOR U37784 ( .A(n38201), .B(n38202), .Z(n38191) );
  AND U37785 ( .A(n38203), .B(n38204), .Z(n38202) );
  XNOR U37786 ( .A(n38201), .B(n38047), .Z(n38204) );
  IV U37787 ( .A(n38050), .Z(n38047) );
  XOR U37788 ( .A(n38205), .B(n38206), .Z(n38050) );
  AND U37789 ( .A(n850), .B(n38207), .Z(n38206) );
  XNOR U37790 ( .A(n38208), .B(n38205), .Z(n38207) );
  XOR U37791 ( .A(n38051), .B(n38201), .Z(n38203) );
  XOR U37792 ( .A(n38209), .B(n38210), .Z(n38051) );
  AND U37793 ( .A(n858), .B(n38168), .Z(n38210) );
  XOR U37794 ( .A(n38209), .B(n38166), .Z(n38168) );
  XOR U37795 ( .A(n38125), .B(n38211), .Z(n38201) );
  AND U37796 ( .A(n38127), .B(n38212), .Z(n38211) );
  XNOR U37797 ( .A(n38125), .B(n38096), .Z(n38212) );
  IV U37798 ( .A(n38099), .Z(n38096) );
  XOR U37799 ( .A(n38213), .B(n38214), .Z(n38099) );
  AND U37800 ( .A(n850), .B(n38215), .Z(n38214) );
  XOR U37801 ( .A(n38216), .B(n38213), .Z(n38215) );
  XOR U37802 ( .A(n38100), .B(n38125), .Z(n38127) );
  XOR U37803 ( .A(n38217), .B(n38218), .Z(n38100) );
  AND U37804 ( .A(n858), .B(n38178), .Z(n38218) );
  XOR U37805 ( .A(n38217), .B(n38176), .Z(n38178) );
  AND U37806 ( .A(n38179), .B(n38109), .Z(n38125) );
  XNOR U37807 ( .A(n38219), .B(n38220), .Z(n38109) );
  AND U37808 ( .A(n850), .B(n38221), .Z(n38220) );
  XNOR U37809 ( .A(n38222), .B(n38219), .Z(n38221) );
  XNOR U37810 ( .A(n38223), .B(n38224), .Z(n850) );
  AND U37811 ( .A(n38225), .B(n38226), .Z(n38224) );
  XOR U37812 ( .A(n38188), .B(n38223), .Z(n38226) );
  AND U37813 ( .A(n38227), .B(n38228), .Z(n38188) );
  XNOR U37814 ( .A(n38185), .B(n38223), .Z(n38225) );
  XNOR U37815 ( .A(n38229), .B(n38230), .Z(n38185) );
  AND U37816 ( .A(n854), .B(n38231), .Z(n38230) );
  XNOR U37817 ( .A(n38232), .B(n38233), .Z(n38231) );
  XOR U37818 ( .A(n38234), .B(n38235), .Z(n38223) );
  AND U37819 ( .A(n38236), .B(n38237), .Z(n38235) );
  XNOR U37820 ( .A(n38234), .B(n38227), .Z(n38237) );
  IV U37821 ( .A(n38198), .Z(n38227) );
  XOR U37822 ( .A(n38238), .B(n38239), .Z(n38198) );
  XOR U37823 ( .A(n38240), .B(n38228), .Z(n38239) );
  AND U37824 ( .A(n38208), .B(n38241), .Z(n38228) );
  AND U37825 ( .A(n38242), .B(n38243), .Z(n38240) );
  XOR U37826 ( .A(n38244), .B(n38238), .Z(n38242) );
  XNOR U37827 ( .A(n38195), .B(n38234), .Z(n38236) );
  XNOR U37828 ( .A(n38245), .B(n38246), .Z(n38195) );
  AND U37829 ( .A(n854), .B(n38247), .Z(n38246) );
  XNOR U37830 ( .A(n38248), .B(n38249), .Z(n38247) );
  XOR U37831 ( .A(n38250), .B(n38251), .Z(n38234) );
  AND U37832 ( .A(n38252), .B(n38253), .Z(n38251) );
  XNOR U37833 ( .A(n38250), .B(n38208), .Z(n38253) );
  XOR U37834 ( .A(n38254), .B(n38243), .Z(n38208) );
  XNOR U37835 ( .A(n38255), .B(n38238), .Z(n38243) );
  XOR U37836 ( .A(n38256), .B(n38257), .Z(n38238) );
  AND U37837 ( .A(n38258), .B(n38259), .Z(n38257) );
  XOR U37838 ( .A(n38260), .B(n38256), .Z(n38258) );
  XNOR U37839 ( .A(n38261), .B(n38262), .Z(n38255) );
  AND U37840 ( .A(n38263), .B(n38264), .Z(n38262) );
  XOR U37841 ( .A(n38261), .B(n38265), .Z(n38263) );
  XNOR U37842 ( .A(n38244), .B(n38241), .Z(n38254) );
  AND U37843 ( .A(n38266), .B(n38267), .Z(n38241) );
  XOR U37844 ( .A(n38268), .B(n38269), .Z(n38244) );
  AND U37845 ( .A(n38270), .B(n38271), .Z(n38269) );
  XOR U37846 ( .A(n38268), .B(n38272), .Z(n38270) );
  XNOR U37847 ( .A(n38205), .B(n38250), .Z(n38252) );
  XNOR U37848 ( .A(n38273), .B(n38274), .Z(n38205) );
  AND U37849 ( .A(n854), .B(n38275), .Z(n38274) );
  XNOR U37850 ( .A(n38276), .B(n38277), .Z(n38275) );
  XOR U37851 ( .A(n38278), .B(n38279), .Z(n38250) );
  AND U37852 ( .A(n38280), .B(n38281), .Z(n38279) );
  XNOR U37853 ( .A(n38278), .B(n38266), .Z(n38281) );
  IV U37854 ( .A(n38216), .Z(n38266) );
  XNOR U37855 ( .A(n38282), .B(n38259), .Z(n38216) );
  XNOR U37856 ( .A(n38283), .B(n38265), .Z(n38259) );
  XOR U37857 ( .A(n38284), .B(n38285), .Z(n38265) );
  NOR U37858 ( .A(n38286), .B(n38287), .Z(n38285) );
  XNOR U37859 ( .A(n38284), .B(n38288), .Z(n38286) );
  XNOR U37860 ( .A(n38264), .B(n38256), .Z(n38283) );
  XOR U37861 ( .A(n38289), .B(n38290), .Z(n38256) );
  AND U37862 ( .A(n38291), .B(n38292), .Z(n38290) );
  XNOR U37863 ( .A(n38289), .B(n38293), .Z(n38291) );
  XNOR U37864 ( .A(n38294), .B(n38261), .Z(n38264) );
  XOR U37865 ( .A(n38295), .B(n38296), .Z(n38261) );
  AND U37866 ( .A(n38297), .B(n38298), .Z(n38296) );
  XOR U37867 ( .A(n38295), .B(n38299), .Z(n38297) );
  XNOR U37868 ( .A(n38300), .B(n38301), .Z(n38294) );
  NOR U37869 ( .A(n38302), .B(n38303), .Z(n38301) );
  XOR U37870 ( .A(n38300), .B(n38304), .Z(n38302) );
  XNOR U37871 ( .A(n38260), .B(n38267), .Z(n38282) );
  NOR U37872 ( .A(n38222), .B(n38305), .Z(n38267) );
  XOR U37873 ( .A(n38272), .B(n38271), .Z(n38260) );
  XNOR U37874 ( .A(n38306), .B(n38268), .Z(n38271) );
  XOR U37875 ( .A(n38307), .B(n38308), .Z(n38268) );
  AND U37876 ( .A(n38309), .B(n38310), .Z(n38308) );
  XOR U37877 ( .A(n38307), .B(n38311), .Z(n38309) );
  XNOR U37878 ( .A(n38312), .B(n38313), .Z(n38306) );
  NOR U37879 ( .A(n38314), .B(n38315), .Z(n38313) );
  XNOR U37880 ( .A(n38312), .B(n38316), .Z(n38314) );
  XOR U37881 ( .A(n38317), .B(n38318), .Z(n38272) );
  NOR U37882 ( .A(n38319), .B(n38320), .Z(n38318) );
  XNOR U37883 ( .A(n38317), .B(n38321), .Z(n38319) );
  XNOR U37884 ( .A(n38213), .B(n38278), .Z(n38280) );
  XNOR U37885 ( .A(n38322), .B(n38323), .Z(n38213) );
  AND U37886 ( .A(n854), .B(n38324), .Z(n38323) );
  XNOR U37887 ( .A(n38325), .B(n38326), .Z(n38324) );
  AND U37888 ( .A(n38219), .B(n38222), .Z(n38278) );
  XOR U37889 ( .A(n38327), .B(n38305), .Z(n38222) );
  XNOR U37890 ( .A(p_input[2048]), .B(p_input[656]), .Z(n38305) );
  XOR U37891 ( .A(n38293), .B(n38292), .Z(n38327) );
  XNOR U37892 ( .A(n38328), .B(n38299), .Z(n38292) );
  XNOR U37893 ( .A(n38288), .B(n38287), .Z(n38299) );
  XOR U37894 ( .A(n38329), .B(n38284), .Z(n38287) );
  XNOR U37895 ( .A(n29266), .B(p_input[666]), .Z(n38284) );
  XNOR U37896 ( .A(p_input[2059]), .B(p_input[667]), .Z(n38329) );
  XOR U37897 ( .A(p_input[2060]), .B(p_input[668]), .Z(n38288) );
  XNOR U37898 ( .A(n38298), .B(n38289), .Z(n38328) );
  XNOR U37899 ( .A(n29494), .B(p_input[657]), .Z(n38289) );
  XOR U37900 ( .A(n38330), .B(n38304), .Z(n38298) );
  XNOR U37901 ( .A(p_input[2063]), .B(p_input[671]), .Z(n38304) );
  XOR U37902 ( .A(n38295), .B(n38303), .Z(n38330) );
  XOR U37903 ( .A(n38331), .B(n38300), .Z(n38303) );
  XOR U37904 ( .A(p_input[2061]), .B(p_input[669]), .Z(n38300) );
  XNOR U37905 ( .A(p_input[2062]), .B(p_input[670]), .Z(n38331) );
  XNOR U37906 ( .A(n29036), .B(p_input[665]), .Z(n38295) );
  XNOR U37907 ( .A(n38311), .B(n38310), .Z(n38293) );
  XNOR U37908 ( .A(n38332), .B(n38316), .Z(n38310) );
  XOR U37909 ( .A(p_input[2056]), .B(p_input[664]), .Z(n38316) );
  XOR U37910 ( .A(n38307), .B(n38315), .Z(n38332) );
  XOR U37911 ( .A(n38333), .B(n38312), .Z(n38315) );
  XOR U37912 ( .A(p_input[2054]), .B(p_input[662]), .Z(n38312) );
  XNOR U37913 ( .A(p_input[2055]), .B(p_input[663]), .Z(n38333) );
  XNOR U37914 ( .A(n29039), .B(p_input[658]), .Z(n38307) );
  XNOR U37915 ( .A(n38321), .B(n38320), .Z(n38311) );
  XOR U37916 ( .A(n38334), .B(n38317), .Z(n38320) );
  XOR U37917 ( .A(p_input[2051]), .B(p_input[659]), .Z(n38317) );
  XNOR U37918 ( .A(p_input[2052]), .B(p_input[660]), .Z(n38334) );
  XOR U37919 ( .A(p_input[2053]), .B(p_input[661]), .Z(n38321) );
  XNOR U37920 ( .A(n38335), .B(n38336), .Z(n38219) );
  AND U37921 ( .A(n854), .B(n38337), .Z(n38336) );
  XNOR U37922 ( .A(n38338), .B(n38339), .Z(n854) );
  AND U37923 ( .A(n38340), .B(n38341), .Z(n38339) );
  XOR U37924 ( .A(n38233), .B(n38338), .Z(n38341) );
  XNOR U37925 ( .A(n38342), .B(n38338), .Z(n38340) );
  XOR U37926 ( .A(n38343), .B(n38344), .Z(n38338) );
  AND U37927 ( .A(n38345), .B(n38346), .Z(n38344) );
  XOR U37928 ( .A(n38248), .B(n38343), .Z(n38346) );
  XOR U37929 ( .A(n38343), .B(n38249), .Z(n38345) );
  XOR U37930 ( .A(n38347), .B(n38348), .Z(n38343) );
  AND U37931 ( .A(n38349), .B(n38350), .Z(n38348) );
  XOR U37932 ( .A(n38276), .B(n38347), .Z(n38350) );
  XOR U37933 ( .A(n38347), .B(n38277), .Z(n38349) );
  XOR U37934 ( .A(n38351), .B(n38352), .Z(n38347) );
  AND U37935 ( .A(n38353), .B(n38354), .Z(n38352) );
  XOR U37936 ( .A(n38351), .B(n38325), .Z(n38354) );
  XNOR U37937 ( .A(n38355), .B(n38356), .Z(n38179) );
  AND U37938 ( .A(n858), .B(n38357), .Z(n38356) );
  XNOR U37939 ( .A(n38358), .B(n38359), .Z(n858) );
  AND U37940 ( .A(n38360), .B(n38361), .Z(n38359) );
  XOR U37941 ( .A(n38358), .B(n38189), .Z(n38361) );
  XNOR U37942 ( .A(n38358), .B(n38149), .Z(n38360) );
  XOR U37943 ( .A(n38362), .B(n38363), .Z(n38358) );
  AND U37944 ( .A(n38364), .B(n38365), .Z(n38363) );
  XOR U37945 ( .A(n38362), .B(n38157), .Z(n38364) );
  XOR U37946 ( .A(n38366), .B(n38367), .Z(n38140) );
  AND U37947 ( .A(n862), .B(n38357), .Z(n38367) );
  XNOR U37948 ( .A(n38355), .B(n38366), .Z(n38357) );
  XNOR U37949 ( .A(n38368), .B(n38369), .Z(n862) );
  AND U37950 ( .A(n38370), .B(n38371), .Z(n38369) );
  XNOR U37951 ( .A(n38372), .B(n38368), .Z(n38371) );
  IV U37952 ( .A(n38189), .Z(n38372) );
  XOR U37953 ( .A(n38342), .B(n38373), .Z(n38189) );
  AND U37954 ( .A(n865), .B(n38374), .Z(n38373) );
  XOR U37955 ( .A(n38232), .B(n38229), .Z(n38374) );
  IV U37956 ( .A(n38342), .Z(n38232) );
  XNOR U37957 ( .A(n38149), .B(n38368), .Z(n38370) );
  XOR U37958 ( .A(n38375), .B(n38376), .Z(n38149) );
  AND U37959 ( .A(n881), .B(n38377), .Z(n38376) );
  XOR U37960 ( .A(n38362), .B(n38378), .Z(n38368) );
  AND U37961 ( .A(n38379), .B(n38365), .Z(n38378) );
  XNOR U37962 ( .A(n38199), .B(n38362), .Z(n38365) );
  XOR U37963 ( .A(n38249), .B(n38380), .Z(n38199) );
  AND U37964 ( .A(n865), .B(n38381), .Z(n38380) );
  XOR U37965 ( .A(n38245), .B(n38249), .Z(n38381) );
  XNOR U37966 ( .A(n38382), .B(n38362), .Z(n38379) );
  IV U37967 ( .A(n38157), .Z(n38382) );
  XOR U37968 ( .A(n38383), .B(n38384), .Z(n38157) );
  AND U37969 ( .A(n881), .B(n38385), .Z(n38384) );
  XOR U37970 ( .A(n38386), .B(n38387), .Z(n38362) );
  AND U37971 ( .A(n38388), .B(n38389), .Z(n38387) );
  XNOR U37972 ( .A(n38209), .B(n38386), .Z(n38389) );
  XOR U37973 ( .A(n38277), .B(n38390), .Z(n38209) );
  AND U37974 ( .A(n865), .B(n38391), .Z(n38390) );
  XOR U37975 ( .A(n38273), .B(n38277), .Z(n38391) );
  XOR U37976 ( .A(n38386), .B(n38166), .Z(n38388) );
  XOR U37977 ( .A(n38392), .B(n38393), .Z(n38166) );
  AND U37978 ( .A(n881), .B(n38394), .Z(n38393) );
  XOR U37979 ( .A(n38395), .B(n38396), .Z(n38386) );
  AND U37980 ( .A(n38397), .B(n38398), .Z(n38396) );
  XNOR U37981 ( .A(n38395), .B(n38217), .Z(n38398) );
  XOR U37982 ( .A(n38326), .B(n38399), .Z(n38217) );
  AND U37983 ( .A(n865), .B(n38400), .Z(n38399) );
  XOR U37984 ( .A(n38322), .B(n38326), .Z(n38400) );
  XNOR U37985 ( .A(n38401), .B(n38395), .Z(n38397) );
  IV U37986 ( .A(n38176), .Z(n38401) );
  XOR U37987 ( .A(n38402), .B(n38403), .Z(n38176) );
  AND U37988 ( .A(n881), .B(n38404), .Z(n38403) );
  AND U37989 ( .A(n38366), .B(n38355), .Z(n38395) );
  XNOR U37990 ( .A(n38405), .B(n38406), .Z(n38355) );
  AND U37991 ( .A(n865), .B(n38337), .Z(n38406) );
  XNOR U37992 ( .A(n38335), .B(n38405), .Z(n38337) );
  XNOR U37993 ( .A(n38407), .B(n38408), .Z(n865) );
  AND U37994 ( .A(n38409), .B(n38410), .Z(n38408) );
  XNOR U37995 ( .A(n38407), .B(n38229), .Z(n38410) );
  IV U37996 ( .A(n38233), .Z(n38229) );
  XOR U37997 ( .A(n38411), .B(n38412), .Z(n38233) );
  AND U37998 ( .A(n869), .B(n38413), .Z(n38412) );
  XOR U37999 ( .A(n38414), .B(n38411), .Z(n38413) );
  XNOR U38000 ( .A(n38407), .B(n38342), .Z(n38409) );
  XOR U38001 ( .A(n38415), .B(n38416), .Z(n38342) );
  AND U38002 ( .A(n877), .B(n38377), .Z(n38416) );
  XOR U38003 ( .A(n38375), .B(n38415), .Z(n38377) );
  XOR U38004 ( .A(n38417), .B(n38418), .Z(n38407) );
  AND U38005 ( .A(n38419), .B(n38420), .Z(n38418) );
  XNOR U38006 ( .A(n38417), .B(n38245), .Z(n38420) );
  IV U38007 ( .A(n38248), .Z(n38245) );
  XOR U38008 ( .A(n38421), .B(n38422), .Z(n38248) );
  AND U38009 ( .A(n869), .B(n38423), .Z(n38422) );
  XOR U38010 ( .A(n38424), .B(n38421), .Z(n38423) );
  XOR U38011 ( .A(n38249), .B(n38417), .Z(n38419) );
  XOR U38012 ( .A(n38425), .B(n38426), .Z(n38249) );
  AND U38013 ( .A(n877), .B(n38385), .Z(n38426) );
  XOR U38014 ( .A(n38425), .B(n38383), .Z(n38385) );
  XOR U38015 ( .A(n38427), .B(n38428), .Z(n38417) );
  AND U38016 ( .A(n38429), .B(n38430), .Z(n38428) );
  XNOR U38017 ( .A(n38427), .B(n38273), .Z(n38430) );
  IV U38018 ( .A(n38276), .Z(n38273) );
  XOR U38019 ( .A(n38431), .B(n38432), .Z(n38276) );
  AND U38020 ( .A(n869), .B(n38433), .Z(n38432) );
  XNOR U38021 ( .A(n38434), .B(n38431), .Z(n38433) );
  XOR U38022 ( .A(n38277), .B(n38427), .Z(n38429) );
  XOR U38023 ( .A(n38435), .B(n38436), .Z(n38277) );
  AND U38024 ( .A(n877), .B(n38394), .Z(n38436) );
  XOR U38025 ( .A(n38435), .B(n38392), .Z(n38394) );
  XOR U38026 ( .A(n38351), .B(n38437), .Z(n38427) );
  AND U38027 ( .A(n38353), .B(n38438), .Z(n38437) );
  XNOR U38028 ( .A(n38351), .B(n38322), .Z(n38438) );
  IV U38029 ( .A(n38325), .Z(n38322) );
  XOR U38030 ( .A(n38439), .B(n38440), .Z(n38325) );
  AND U38031 ( .A(n869), .B(n38441), .Z(n38440) );
  XOR U38032 ( .A(n38442), .B(n38439), .Z(n38441) );
  XOR U38033 ( .A(n38326), .B(n38351), .Z(n38353) );
  XOR U38034 ( .A(n38443), .B(n38444), .Z(n38326) );
  AND U38035 ( .A(n877), .B(n38404), .Z(n38444) );
  XOR U38036 ( .A(n38443), .B(n38402), .Z(n38404) );
  AND U38037 ( .A(n38405), .B(n38335), .Z(n38351) );
  XNOR U38038 ( .A(n38445), .B(n38446), .Z(n38335) );
  AND U38039 ( .A(n869), .B(n38447), .Z(n38446) );
  XNOR U38040 ( .A(n38448), .B(n38445), .Z(n38447) );
  XNOR U38041 ( .A(n38449), .B(n38450), .Z(n869) );
  AND U38042 ( .A(n38451), .B(n38452), .Z(n38450) );
  XOR U38043 ( .A(n38414), .B(n38449), .Z(n38452) );
  AND U38044 ( .A(n38453), .B(n38454), .Z(n38414) );
  XNOR U38045 ( .A(n38411), .B(n38449), .Z(n38451) );
  XNOR U38046 ( .A(n38455), .B(n38456), .Z(n38411) );
  AND U38047 ( .A(n873), .B(n38457), .Z(n38456) );
  XNOR U38048 ( .A(n38458), .B(n38459), .Z(n38457) );
  XOR U38049 ( .A(n38460), .B(n38461), .Z(n38449) );
  AND U38050 ( .A(n38462), .B(n38463), .Z(n38461) );
  XNOR U38051 ( .A(n38460), .B(n38453), .Z(n38463) );
  IV U38052 ( .A(n38424), .Z(n38453) );
  XOR U38053 ( .A(n38464), .B(n38465), .Z(n38424) );
  XOR U38054 ( .A(n38466), .B(n38454), .Z(n38465) );
  AND U38055 ( .A(n38434), .B(n38467), .Z(n38454) );
  AND U38056 ( .A(n38468), .B(n38469), .Z(n38466) );
  XOR U38057 ( .A(n38470), .B(n38464), .Z(n38468) );
  XNOR U38058 ( .A(n38421), .B(n38460), .Z(n38462) );
  XNOR U38059 ( .A(n38471), .B(n38472), .Z(n38421) );
  AND U38060 ( .A(n873), .B(n38473), .Z(n38472) );
  XNOR U38061 ( .A(n38474), .B(n38475), .Z(n38473) );
  XOR U38062 ( .A(n38476), .B(n38477), .Z(n38460) );
  AND U38063 ( .A(n38478), .B(n38479), .Z(n38477) );
  XNOR U38064 ( .A(n38476), .B(n38434), .Z(n38479) );
  XOR U38065 ( .A(n38480), .B(n38469), .Z(n38434) );
  XNOR U38066 ( .A(n38481), .B(n38464), .Z(n38469) );
  XOR U38067 ( .A(n38482), .B(n38483), .Z(n38464) );
  AND U38068 ( .A(n38484), .B(n38485), .Z(n38483) );
  XOR U38069 ( .A(n38486), .B(n38482), .Z(n38484) );
  XNOR U38070 ( .A(n38487), .B(n38488), .Z(n38481) );
  AND U38071 ( .A(n38489), .B(n38490), .Z(n38488) );
  XOR U38072 ( .A(n38487), .B(n38491), .Z(n38489) );
  XNOR U38073 ( .A(n38470), .B(n38467), .Z(n38480) );
  AND U38074 ( .A(n38492), .B(n38493), .Z(n38467) );
  XOR U38075 ( .A(n38494), .B(n38495), .Z(n38470) );
  AND U38076 ( .A(n38496), .B(n38497), .Z(n38495) );
  XOR U38077 ( .A(n38494), .B(n38498), .Z(n38496) );
  XNOR U38078 ( .A(n38431), .B(n38476), .Z(n38478) );
  XNOR U38079 ( .A(n38499), .B(n38500), .Z(n38431) );
  AND U38080 ( .A(n873), .B(n38501), .Z(n38500) );
  XNOR U38081 ( .A(n38502), .B(n38503), .Z(n38501) );
  XOR U38082 ( .A(n38504), .B(n38505), .Z(n38476) );
  AND U38083 ( .A(n38506), .B(n38507), .Z(n38505) );
  XNOR U38084 ( .A(n38504), .B(n38492), .Z(n38507) );
  IV U38085 ( .A(n38442), .Z(n38492) );
  XNOR U38086 ( .A(n38508), .B(n38485), .Z(n38442) );
  XNOR U38087 ( .A(n38509), .B(n38491), .Z(n38485) );
  XOR U38088 ( .A(n38510), .B(n38511), .Z(n38491) );
  NOR U38089 ( .A(n38512), .B(n38513), .Z(n38511) );
  XNOR U38090 ( .A(n38510), .B(n38514), .Z(n38512) );
  XNOR U38091 ( .A(n38490), .B(n38482), .Z(n38509) );
  XOR U38092 ( .A(n38515), .B(n38516), .Z(n38482) );
  AND U38093 ( .A(n38517), .B(n38518), .Z(n38516) );
  XNOR U38094 ( .A(n38515), .B(n38519), .Z(n38517) );
  XNOR U38095 ( .A(n38520), .B(n38487), .Z(n38490) );
  XOR U38096 ( .A(n38521), .B(n38522), .Z(n38487) );
  AND U38097 ( .A(n38523), .B(n38524), .Z(n38522) );
  XOR U38098 ( .A(n38521), .B(n38525), .Z(n38523) );
  XNOR U38099 ( .A(n38526), .B(n38527), .Z(n38520) );
  NOR U38100 ( .A(n38528), .B(n38529), .Z(n38527) );
  XOR U38101 ( .A(n38526), .B(n38530), .Z(n38528) );
  XNOR U38102 ( .A(n38486), .B(n38493), .Z(n38508) );
  NOR U38103 ( .A(n38448), .B(n38531), .Z(n38493) );
  XOR U38104 ( .A(n38498), .B(n38497), .Z(n38486) );
  XNOR U38105 ( .A(n38532), .B(n38494), .Z(n38497) );
  XOR U38106 ( .A(n38533), .B(n38534), .Z(n38494) );
  AND U38107 ( .A(n38535), .B(n38536), .Z(n38534) );
  XOR U38108 ( .A(n38533), .B(n38537), .Z(n38535) );
  XNOR U38109 ( .A(n38538), .B(n38539), .Z(n38532) );
  NOR U38110 ( .A(n38540), .B(n38541), .Z(n38539) );
  XNOR U38111 ( .A(n38538), .B(n38542), .Z(n38540) );
  XOR U38112 ( .A(n38543), .B(n38544), .Z(n38498) );
  NOR U38113 ( .A(n38545), .B(n38546), .Z(n38544) );
  XNOR U38114 ( .A(n38543), .B(n38547), .Z(n38545) );
  XNOR U38115 ( .A(n38439), .B(n38504), .Z(n38506) );
  XNOR U38116 ( .A(n38548), .B(n38549), .Z(n38439) );
  AND U38117 ( .A(n873), .B(n38550), .Z(n38549) );
  XNOR U38118 ( .A(n38551), .B(n38552), .Z(n38550) );
  AND U38119 ( .A(n38445), .B(n38448), .Z(n38504) );
  XOR U38120 ( .A(n38553), .B(n38531), .Z(n38448) );
  XNOR U38121 ( .A(p_input[2048]), .B(p_input[672]), .Z(n38531) );
  XOR U38122 ( .A(n38519), .B(n38518), .Z(n38553) );
  XNOR U38123 ( .A(n38554), .B(n38525), .Z(n38518) );
  XNOR U38124 ( .A(n38514), .B(n38513), .Z(n38525) );
  XOR U38125 ( .A(n38555), .B(n38510), .Z(n38513) );
  XNOR U38126 ( .A(n29266), .B(p_input[682]), .Z(n38510) );
  XNOR U38127 ( .A(p_input[2059]), .B(p_input[683]), .Z(n38555) );
  XOR U38128 ( .A(p_input[2060]), .B(p_input[684]), .Z(n38514) );
  XNOR U38129 ( .A(n38524), .B(n38515), .Z(n38554) );
  XNOR U38130 ( .A(n29494), .B(p_input[673]), .Z(n38515) );
  XOR U38131 ( .A(n38556), .B(n38530), .Z(n38524) );
  XNOR U38132 ( .A(p_input[2063]), .B(p_input[687]), .Z(n38530) );
  XOR U38133 ( .A(n38521), .B(n38529), .Z(n38556) );
  XOR U38134 ( .A(n38557), .B(n38526), .Z(n38529) );
  XOR U38135 ( .A(p_input[2061]), .B(p_input[685]), .Z(n38526) );
  XNOR U38136 ( .A(p_input[2062]), .B(p_input[686]), .Z(n38557) );
  XNOR U38137 ( .A(n29036), .B(p_input[681]), .Z(n38521) );
  XNOR U38138 ( .A(n38537), .B(n38536), .Z(n38519) );
  XNOR U38139 ( .A(n38558), .B(n38542), .Z(n38536) );
  XOR U38140 ( .A(p_input[2056]), .B(p_input[680]), .Z(n38542) );
  XOR U38141 ( .A(n38533), .B(n38541), .Z(n38558) );
  XOR U38142 ( .A(n38559), .B(n38538), .Z(n38541) );
  XOR U38143 ( .A(p_input[2054]), .B(p_input[678]), .Z(n38538) );
  XNOR U38144 ( .A(p_input[2055]), .B(p_input[679]), .Z(n38559) );
  XNOR U38145 ( .A(n29039), .B(p_input[674]), .Z(n38533) );
  XNOR U38146 ( .A(n38547), .B(n38546), .Z(n38537) );
  XOR U38147 ( .A(n38560), .B(n38543), .Z(n38546) );
  XOR U38148 ( .A(p_input[2051]), .B(p_input[675]), .Z(n38543) );
  XNOR U38149 ( .A(p_input[2052]), .B(p_input[676]), .Z(n38560) );
  XOR U38150 ( .A(p_input[2053]), .B(p_input[677]), .Z(n38547) );
  XNOR U38151 ( .A(n38561), .B(n38562), .Z(n38445) );
  AND U38152 ( .A(n873), .B(n38563), .Z(n38562) );
  XNOR U38153 ( .A(n38564), .B(n38565), .Z(n873) );
  AND U38154 ( .A(n38566), .B(n38567), .Z(n38565) );
  XOR U38155 ( .A(n38459), .B(n38564), .Z(n38567) );
  XNOR U38156 ( .A(n38568), .B(n38564), .Z(n38566) );
  XOR U38157 ( .A(n38569), .B(n38570), .Z(n38564) );
  AND U38158 ( .A(n38571), .B(n38572), .Z(n38570) );
  XOR U38159 ( .A(n38474), .B(n38569), .Z(n38572) );
  XOR U38160 ( .A(n38569), .B(n38475), .Z(n38571) );
  XOR U38161 ( .A(n38573), .B(n38574), .Z(n38569) );
  AND U38162 ( .A(n38575), .B(n38576), .Z(n38574) );
  XOR U38163 ( .A(n38502), .B(n38573), .Z(n38576) );
  XOR U38164 ( .A(n38573), .B(n38503), .Z(n38575) );
  XOR U38165 ( .A(n38577), .B(n38578), .Z(n38573) );
  AND U38166 ( .A(n38579), .B(n38580), .Z(n38578) );
  XOR U38167 ( .A(n38577), .B(n38551), .Z(n38580) );
  XNOR U38168 ( .A(n38581), .B(n38582), .Z(n38405) );
  AND U38169 ( .A(n877), .B(n38583), .Z(n38582) );
  XNOR U38170 ( .A(n38584), .B(n38585), .Z(n877) );
  AND U38171 ( .A(n38586), .B(n38587), .Z(n38585) );
  XOR U38172 ( .A(n38584), .B(n38415), .Z(n38587) );
  XNOR U38173 ( .A(n38584), .B(n38375), .Z(n38586) );
  XOR U38174 ( .A(n38588), .B(n38589), .Z(n38584) );
  AND U38175 ( .A(n38590), .B(n38591), .Z(n38589) );
  XOR U38176 ( .A(n38588), .B(n38383), .Z(n38590) );
  XOR U38177 ( .A(n38592), .B(n38593), .Z(n38366) );
  AND U38178 ( .A(n881), .B(n38583), .Z(n38593) );
  XNOR U38179 ( .A(n38581), .B(n38592), .Z(n38583) );
  XNOR U38180 ( .A(n38594), .B(n38595), .Z(n881) );
  AND U38181 ( .A(n38596), .B(n38597), .Z(n38595) );
  XNOR U38182 ( .A(n38598), .B(n38594), .Z(n38597) );
  IV U38183 ( .A(n38415), .Z(n38598) );
  XOR U38184 ( .A(n38568), .B(n38599), .Z(n38415) );
  AND U38185 ( .A(n884), .B(n38600), .Z(n38599) );
  XOR U38186 ( .A(n38458), .B(n38455), .Z(n38600) );
  IV U38187 ( .A(n38568), .Z(n38458) );
  XNOR U38188 ( .A(n38375), .B(n38594), .Z(n38596) );
  XOR U38189 ( .A(n38601), .B(n38602), .Z(n38375) );
  AND U38190 ( .A(n900), .B(n38603), .Z(n38602) );
  XOR U38191 ( .A(n38588), .B(n38604), .Z(n38594) );
  AND U38192 ( .A(n38605), .B(n38591), .Z(n38604) );
  XNOR U38193 ( .A(n38425), .B(n38588), .Z(n38591) );
  XOR U38194 ( .A(n38475), .B(n38606), .Z(n38425) );
  AND U38195 ( .A(n884), .B(n38607), .Z(n38606) );
  XOR U38196 ( .A(n38471), .B(n38475), .Z(n38607) );
  XNOR U38197 ( .A(n38608), .B(n38588), .Z(n38605) );
  IV U38198 ( .A(n38383), .Z(n38608) );
  XOR U38199 ( .A(n38609), .B(n38610), .Z(n38383) );
  AND U38200 ( .A(n900), .B(n38611), .Z(n38610) );
  XOR U38201 ( .A(n38612), .B(n38613), .Z(n38588) );
  AND U38202 ( .A(n38614), .B(n38615), .Z(n38613) );
  XNOR U38203 ( .A(n38435), .B(n38612), .Z(n38615) );
  XOR U38204 ( .A(n38503), .B(n38616), .Z(n38435) );
  AND U38205 ( .A(n884), .B(n38617), .Z(n38616) );
  XOR U38206 ( .A(n38499), .B(n38503), .Z(n38617) );
  XOR U38207 ( .A(n38612), .B(n38392), .Z(n38614) );
  XOR U38208 ( .A(n38618), .B(n38619), .Z(n38392) );
  AND U38209 ( .A(n900), .B(n38620), .Z(n38619) );
  XOR U38210 ( .A(n38621), .B(n38622), .Z(n38612) );
  AND U38211 ( .A(n38623), .B(n38624), .Z(n38622) );
  XNOR U38212 ( .A(n38621), .B(n38443), .Z(n38624) );
  XOR U38213 ( .A(n38552), .B(n38625), .Z(n38443) );
  AND U38214 ( .A(n884), .B(n38626), .Z(n38625) );
  XOR U38215 ( .A(n38548), .B(n38552), .Z(n38626) );
  XNOR U38216 ( .A(n38627), .B(n38621), .Z(n38623) );
  IV U38217 ( .A(n38402), .Z(n38627) );
  XOR U38218 ( .A(n38628), .B(n38629), .Z(n38402) );
  AND U38219 ( .A(n900), .B(n38630), .Z(n38629) );
  AND U38220 ( .A(n38592), .B(n38581), .Z(n38621) );
  XNOR U38221 ( .A(n38631), .B(n38632), .Z(n38581) );
  AND U38222 ( .A(n884), .B(n38563), .Z(n38632) );
  XNOR U38223 ( .A(n38561), .B(n38631), .Z(n38563) );
  XNOR U38224 ( .A(n38633), .B(n38634), .Z(n884) );
  AND U38225 ( .A(n38635), .B(n38636), .Z(n38634) );
  XNOR U38226 ( .A(n38633), .B(n38455), .Z(n38636) );
  IV U38227 ( .A(n38459), .Z(n38455) );
  XOR U38228 ( .A(n38637), .B(n38638), .Z(n38459) );
  AND U38229 ( .A(n888), .B(n38639), .Z(n38638) );
  XOR U38230 ( .A(n38640), .B(n38637), .Z(n38639) );
  XNOR U38231 ( .A(n38633), .B(n38568), .Z(n38635) );
  XOR U38232 ( .A(n38641), .B(n38642), .Z(n38568) );
  AND U38233 ( .A(n896), .B(n38603), .Z(n38642) );
  XOR U38234 ( .A(n38601), .B(n38641), .Z(n38603) );
  XOR U38235 ( .A(n38643), .B(n38644), .Z(n38633) );
  AND U38236 ( .A(n38645), .B(n38646), .Z(n38644) );
  XNOR U38237 ( .A(n38643), .B(n38471), .Z(n38646) );
  IV U38238 ( .A(n38474), .Z(n38471) );
  XOR U38239 ( .A(n38647), .B(n38648), .Z(n38474) );
  AND U38240 ( .A(n888), .B(n38649), .Z(n38648) );
  XOR U38241 ( .A(n38650), .B(n38647), .Z(n38649) );
  XOR U38242 ( .A(n38475), .B(n38643), .Z(n38645) );
  XOR U38243 ( .A(n38651), .B(n38652), .Z(n38475) );
  AND U38244 ( .A(n896), .B(n38611), .Z(n38652) );
  XOR U38245 ( .A(n38651), .B(n38609), .Z(n38611) );
  XOR U38246 ( .A(n38653), .B(n38654), .Z(n38643) );
  AND U38247 ( .A(n38655), .B(n38656), .Z(n38654) );
  XNOR U38248 ( .A(n38653), .B(n38499), .Z(n38656) );
  IV U38249 ( .A(n38502), .Z(n38499) );
  XOR U38250 ( .A(n38657), .B(n38658), .Z(n38502) );
  AND U38251 ( .A(n888), .B(n38659), .Z(n38658) );
  XNOR U38252 ( .A(n38660), .B(n38657), .Z(n38659) );
  XOR U38253 ( .A(n38503), .B(n38653), .Z(n38655) );
  XOR U38254 ( .A(n38661), .B(n38662), .Z(n38503) );
  AND U38255 ( .A(n896), .B(n38620), .Z(n38662) );
  XOR U38256 ( .A(n38661), .B(n38618), .Z(n38620) );
  XOR U38257 ( .A(n38577), .B(n38663), .Z(n38653) );
  AND U38258 ( .A(n38579), .B(n38664), .Z(n38663) );
  XNOR U38259 ( .A(n38577), .B(n38548), .Z(n38664) );
  IV U38260 ( .A(n38551), .Z(n38548) );
  XOR U38261 ( .A(n38665), .B(n38666), .Z(n38551) );
  AND U38262 ( .A(n888), .B(n38667), .Z(n38666) );
  XOR U38263 ( .A(n38668), .B(n38665), .Z(n38667) );
  XOR U38264 ( .A(n38552), .B(n38577), .Z(n38579) );
  XOR U38265 ( .A(n38669), .B(n38670), .Z(n38552) );
  AND U38266 ( .A(n896), .B(n38630), .Z(n38670) );
  XOR U38267 ( .A(n38669), .B(n38628), .Z(n38630) );
  AND U38268 ( .A(n38631), .B(n38561), .Z(n38577) );
  XNOR U38269 ( .A(n38671), .B(n38672), .Z(n38561) );
  AND U38270 ( .A(n888), .B(n38673), .Z(n38672) );
  XNOR U38271 ( .A(n38674), .B(n38671), .Z(n38673) );
  XNOR U38272 ( .A(n38675), .B(n38676), .Z(n888) );
  AND U38273 ( .A(n38677), .B(n38678), .Z(n38676) );
  XOR U38274 ( .A(n38640), .B(n38675), .Z(n38678) );
  AND U38275 ( .A(n38679), .B(n38680), .Z(n38640) );
  XNOR U38276 ( .A(n38637), .B(n38675), .Z(n38677) );
  XNOR U38277 ( .A(n38681), .B(n38682), .Z(n38637) );
  AND U38278 ( .A(n892), .B(n38683), .Z(n38682) );
  XNOR U38279 ( .A(n38684), .B(n38685), .Z(n38683) );
  XOR U38280 ( .A(n38686), .B(n38687), .Z(n38675) );
  AND U38281 ( .A(n38688), .B(n38689), .Z(n38687) );
  XNOR U38282 ( .A(n38686), .B(n38679), .Z(n38689) );
  IV U38283 ( .A(n38650), .Z(n38679) );
  XOR U38284 ( .A(n38690), .B(n38691), .Z(n38650) );
  XOR U38285 ( .A(n38692), .B(n38680), .Z(n38691) );
  AND U38286 ( .A(n38660), .B(n38693), .Z(n38680) );
  AND U38287 ( .A(n38694), .B(n38695), .Z(n38692) );
  XOR U38288 ( .A(n38696), .B(n38690), .Z(n38694) );
  XNOR U38289 ( .A(n38647), .B(n38686), .Z(n38688) );
  XNOR U38290 ( .A(n38697), .B(n38698), .Z(n38647) );
  AND U38291 ( .A(n892), .B(n38699), .Z(n38698) );
  XNOR U38292 ( .A(n38700), .B(n38701), .Z(n38699) );
  XOR U38293 ( .A(n38702), .B(n38703), .Z(n38686) );
  AND U38294 ( .A(n38704), .B(n38705), .Z(n38703) );
  XNOR U38295 ( .A(n38702), .B(n38660), .Z(n38705) );
  XOR U38296 ( .A(n38706), .B(n38695), .Z(n38660) );
  XNOR U38297 ( .A(n38707), .B(n38690), .Z(n38695) );
  XOR U38298 ( .A(n38708), .B(n38709), .Z(n38690) );
  AND U38299 ( .A(n38710), .B(n38711), .Z(n38709) );
  XOR U38300 ( .A(n38712), .B(n38708), .Z(n38710) );
  XNOR U38301 ( .A(n38713), .B(n38714), .Z(n38707) );
  AND U38302 ( .A(n38715), .B(n38716), .Z(n38714) );
  XOR U38303 ( .A(n38713), .B(n38717), .Z(n38715) );
  XNOR U38304 ( .A(n38696), .B(n38693), .Z(n38706) );
  AND U38305 ( .A(n38718), .B(n38719), .Z(n38693) );
  XOR U38306 ( .A(n38720), .B(n38721), .Z(n38696) );
  AND U38307 ( .A(n38722), .B(n38723), .Z(n38721) );
  XOR U38308 ( .A(n38720), .B(n38724), .Z(n38722) );
  XNOR U38309 ( .A(n38657), .B(n38702), .Z(n38704) );
  XNOR U38310 ( .A(n38725), .B(n38726), .Z(n38657) );
  AND U38311 ( .A(n892), .B(n38727), .Z(n38726) );
  XNOR U38312 ( .A(n38728), .B(n38729), .Z(n38727) );
  XOR U38313 ( .A(n38730), .B(n38731), .Z(n38702) );
  AND U38314 ( .A(n38732), .B(n38733), .Z(n38731) );
  XNOR U38315 ( .A(n38730), .B(n38718), .Z(n38733) );
  IV U38316 ( .A(n38668), .Z(n38718) );
  XNOR U38317 ( .A(n38734), .B(n38711), .Z(n38668) );
  XNOR U38318 ( .A(n38735), .B(n38717), .Z(n38711) );
  XOR U38319 ( .A(n38736), .B(n38737), .Z(n38717) );
  NOR U38320 ( .A(n38738), .B(n38739), .Z(n38737) );
  XNOR U38321 ( .A(n38736), .B(n38740), .Z(n38738) );
  XNOR U38322 ( .A(n38716), .B(n38708), .Z(n38735) );
  XOR U38323 ( .A(n38741), .B(n38742), .Z(n38708) );
  AND U38324 ( .A(n38743), .B(n38744), .Z(n38742) );
  XNOR U38325 ( .A(n38741), .B(n38745), .Z(n38743) );
  XNOR U38326 ( .A(n38746), .B(n38713), .Z(n38716) );
  XOR U38327 ( .A(n38747), .B(n38748), .Z(n38713) );
  AND U38328 ( .A(n38749), .B(n38750), .Z(n38748) );
  XOR U38329 ( .A(n38747), .B(n38751), .Z(n38749) );
  XNOR U38330 ( .A(n38752), .B(n38753), .Z(n38746) );
  NOR U38331 ( .A(n38754), .B(n38755), .Z(n38753) );
  XOR U38332 ( .A(n38752), .B(n38756), .Z(n38754) );
  XNOR U38333 ( .A(n38712), .B(n38719), .Z(n38734) );
  NOR U38334 ( .A(n38674), .B(n38757), .Z(n38719) );
  XOR U38335 ( .A(n38724), .B(n38723), .Z(n38712) );
  XNOR U38336 ( .A(n38758), .B(n38720), .Z(n38723) );
  XOR U38337 ( .A(n38759), .B(n38760), .Z(n38720) );
  AND U38338 ( .A(n38761), .B(n38762), .Z(n38760) );
  XOR U38339 ( .A(n38759), .B(n38763), .Z(n38761) );
  XNOR U38340 ( .A(n38764), .B(n38765), .Z(n38758) );
  NOR U38341 ( .A(n38766), .B(n38767), .Z(n38765) );
  XNOR U38342 ( .A(n38764), .B(n38768), .Z(n38766) );
  XOR U38343 ( .A(n38769), .B(n38770), .Z(n38724) );
  NOR U38344 ( .A(n38771), .B(n38772), .Z(n38770) );
  XNOR U38345 ( .A(n38769), .B(n38773), .Z(n38771) );
  XNOR U38346 ( .A(n38665), .B(n38730), .Z(n38732) );
  XNOR U38347 ( .A(n38774), .B(n38775), .Z(n38665) );
  AND U38348 ( .A(n892), .B(n38776), .Z(n38775) );
  XNOR U38349 ( .A(n38777), .B(n38778), .Z(n38776) );
  AND U38350 ( .A(n38671), .B(n38674), .Z(n38730) );
  XOR U38351 ( .A(n38779), .B(n38757), .Z(n38674) );
  XNOR U38352 ( .A(p_input[2048]), .B(p_input[688]), .Z(n38757) );
  XOR U38353 ( .A(n38745), .B(n38744), .Z(n38779) );
  XNOR U38354 ( .A(n38780), .B(n38751), .Z(n38744) );
  XNOR U38355 ( .A(n38740), .B(n38739), .Z(n38751) );
  XOR U38356 ( .A(n38781), .B(n38736), .Z(n38739) );
  XNOR U38357 ( .A(n29266), .B(p_input[698]), .Z(n38736) );
  XNOR U38358 ( .A(p_input[2059]), .B(p_input[699]), .Z(n38781) );
  XOR U38359 ( .A(p_input[2060]), .B(p_input[700]), .Z(n38740) );
  XNOR U38360 ( .A(n38750), .B(n38741), .Z(n38780) );
  XNOR U38361 ( .A(n29494), .B(p_input[689]), .Z(n38741) );
  XOR U38362 ( .A(n38782), .B(n38756), .Z(n38750) );
  XNOR U38363 ( .A(p_input[2063]), .B(p_input[703]), .Z(n38756) );
  XOR U38364 ( .A(n38747), .B(n38755), .Z(n38782) );
  XOR U38365 ( .A(n38783), .B(n38752), .Z(n38755) );
  XOR U38366 ( .A(p_input[2061]), .B(p_input[701]), .Z(n38752) );
  XNOR U38367 ( .A(p_input[2062]), .B(p_input[702]), .Z(n38783) );
  XNOR U38368 ( .A(n29036), .B(p_input[697]), .Z(n38747) );
  XNOR U38369 ( .A(n38763), .B(n38762), .Z(n38745) );
  XNOR U38370 ( .A(n38784), .B(n38768), .Z(n38762) );
  XOR U38371 ( .A(p_input[2056]), .B(p_input[696]), .Z(n38768) );
  XOR U38372 ( .A(n38759), .B(n38767), .Z(n38784) );
  XOR U38373 ( .A(n38785), .B(n38764), .Z(n38767) );
  XOR U38374 ( .A(p_input[2054]), .B(p_input[694]), .Z(n38764) );
  XNOR U38375 ( .A(p_input[2055]), .B(p_input[695]), .Z(n38785) );
  XNOR U38376 ( .A(n29039), .B(p_input[690]), .Z(n38759) );
  XNOR U38377 ( .A(n38773), .B(n38772), .Z(n38763) );
  XOR U38378 ( .A(n38786), .B(n38769), .Z(n38772) );
  XOR U38379 ( .A(p_input[2051]), .B(p_input[691]), .Z(n38769) );
  XNOR U38380 ( .A(p_input[2052]), .B(p_input[692]), .Z(n38786) );
  XOR U38381 ( .A(p_input[2053]), .B(p_input[693]), .Z(n38773) );
  XNOR U38382 ( .A(n38787), .B(n38788), .Z(n38671) );
  AND U38383 ( .A(n892), .B(n38789), .Z(n38788) );
  XNOR U38384 ( .A(n38790), .B(n38791), .Z(n892) );
  AND U38385 ( .A(n38792), .B(n38793), .Z(n38791) );
  XOR U38386 ( .A(n38685), .B(n38790), .Z(n38793) );
  XNOR U38387 ( .A(n38794), .B(n38790), .Z(n38792) );
  XOR U38388 ( .A(n38795), .B(n38796), .Z(n38790) );
  AND U38389 ( .A(n38797), .B(n38798), .Z(n38796) );
  XOR U38390 ( .A(n38700), .B(n38795), .Z(n38798) );
  XOR U38391 ( .A(n38795), .B(n38701), .Z(n38797) );
  XOR U38392 ( .A(n38799), .B(n38800), .Z(n38795) );
  AND U38393 ( .A(n38801), .B(n38802), .Z(n38800) );
  XOR U38394 ( .A(n38728), .B(n38799), .Z(n38802) );
  XOR U38395 ( .A(n38799), .B(n38729), .Z(n38801) );
  XOR U38396 ( .A(n38803), .B(n38804), .Z(n38799) );
  AND U38397 ( .A(n38805), .B(n38806), .Z(n38804) );
  XOR U38398 ( .A(n38803), .B(n38777), .Z(n38806) );
  XNOR U38399 ( .A(n38807), .B(n38808), .Z(n38631) );
  AND U38400 ( .A(n896), .B(n38809), .Z(n38808) );
  XNOR U38401 ( .A(n38810), .B(n38811), .Z(n896) );
  AND U38402 ( .A(n38812), .B(n38813), .Z(n38811) );
  XOR U38403 ( .A(n38810), .B(n38641), .Z(n38813) );
  XNOR U38404 ( .A(n38810), .B(n38601), .Z(n38812) );
  XOR U38405 ( .A(n38814), .B(n38815), .Z(n38810) );
  AND U38406 ( .A(n38816), .B(n38817), .Z(n38815) );
  XOR U38407 ( .A(n38814), .B(n38609), .Z(n38816) );
  XOR U38408 ( .A(n38818), .B(n38819), .Z(n38592) );
  AND U38409 ( .A(n900), .B(n38809), .Z(n38819) );
  XNOR U38410 ( .A(n38807), .B(n38818), .Z(n38809) );
  XNOR U38411 ( .A(n38820), .B(n38821), .Z(n900) );
  AND U38412 ( .A(n38822), .B(n38823), .Z(n38821) );
  XNOR U38413 ( .A(n38824), .B(n38820), .Z(n38823) );
  IV U38414 ( .A(n38641), .Z(n38824) );
  XOR U38415 ( .A(n38794), .B(n38825), .Z(n38641) );
  AND U38416 ( .A(n903), .B(n38826), .Z(n38825) );
  XOR U38417 ( .A(n38684), .B(n38681), .Z(n38826) );
  IV U38418 ( .A(n38794), .Z(n38684) );
  XNOR U38419 ( .A(n38601), .B(n38820), .Z(n38822) );
  XOR U38420 ( .A(n38827), .B(n38828), .Z(n38601) );
  AND U38421 ( .A(n919), .B(n38829), .Z(n38828) );
  XOR U38422 ( .A(n38814), .B(n38830), .Z(n38820) );
  AND U38423 ( .A(n38831), .B(n38817), .Z(n38830) );
  XNOR U38424 ( .A(n38651), .B(n38814), .Z(n38817) );
  XOR U38425 ( .A(n38701), .B(n38832), .Z(n38651) );
  AND U38426 ( .A(n903), .B(n38833), .Z(n38832) );
  XOR U38427 ( .A(n38697), .B(n38701), .Z(n38833) );
  XNOR U38428 ( .A(n38834), .B(n38814), .Z(n38831) );
  IV U38429 ( .A(n38609), .Z(n38834) );
  XOR U38430 ( .A(n38835), .B(n38836), .Z(n38609) );
  AND U38431 ( .A(n919), .B(n38837), .Z(n38836) );
  XOR U38432 ( .A(n38838), .B(n38839), .Z(n38814) );
  AND U38433 ( .A(n38840), .B(n38841), .Z(n38839) );
  XNOR U38434 ( .A(n38661), .B(n38838), .Z(n38841) );
  XOR U38435 ( .A(n38729), .B(n38842), .Z(n38661) );
  AND U38436 ( .A(n903), .B(n38843), .Z(n38842) );
  XOR U38437 ( .A(n38725), .B(n38729), .Z(n38843) );
  XOR U38438 ( .A(n38838), .B(n38618), .Z(n38840) );
  XOR U38439 ( .A(n38844), .B(n38845), .Z(n38618) );
  AND U38440 ( .A(n919), .B(n38846), .Z(n38845) );
  XOR U38441 ( .A(n38847), .B(n38848), .Z(n38838) );
  AND U38442 ( .A(n38849), .B(n38850), .Z(n38848) );
  XNOR U38443 ( .A(n38847), .B(n38669), .Z(n38850) );
  XOR U38444 ( .A(n38778), .B(n38851), .Z(n38669) );
  AND U38445 ( .A(n903), .B(n38852), .Z(n38851) );
  XOR U38446 ( .A(n38774), .B(n38778), .Z(n38852) );
  XNOR U38447 ( .A(n38853), .B(n38847), .Z(n38849) );
  IV U38448 ( .A(n38628), .Z(n38853) );
  XOR U38449 ( .A(n38854), .B(n38855), .Z(n38628) );
  AND U38450 ( .A(n919), .B(n38856), .Z(n38855) );
  AND U38451 ( .A(n38818), .B(n38807), .Z(n38847) );
  XNOR U38452 ( .A(n38857), .B(n38858), .Z(n38807) );
  AND U38453 ( .A(n903), .B(n38789), .Z(n38858) );
  XNOR U38454 ( .A(n38787), .B(n38857), .Z(n38789) );
  XNOR U38455 ( .A(n38859), .B(n38860), .Z(n903) );
  AND U38456 ( .A(n38861), .B(n38862), .Z(n38860) );
  XNOR U38457 ( .A(n38859), .B(n38681), .Z(n38862) );
  IV U38458 ( .A(n38685), .Z(n38681) );
  XOR U38459 ( .A(n38863), .B(n38864), .Z(n38685) );
  AND U38460 ( .A(n907), .B(n38865), .Z(n38864) );
  XOR U38461 ( .A(n38866), .B(n38863), .Z(n38865) );
  XNOR U38462 ( .A(n38859), .B(n38794), .Z(n38861) );
  XOR U38463 ( .A(n38867), .B(n38868), .Z(n38794) );
  AND U38464 ( .A(n915), .B(n38829), .Z(n38868) );
  XOR U38465 ( .A(n38827), .B(n38867), .Z(n38829) );
  XOR U38466 ( .A(n38869), .B(n38870), .Z(n38859) );
  AND U38467 ( .A(n38871), .B(n38872), .Z(n38870) );
  XNOR U38468 ( .A(n38869), .B(n38697), .Z(n38872) );
  IV U38469 ( .A(n38700), .Z(n38697) );
  XOR U38470 ( .A(n38873), .B(n38874), .Z(n38700) );
  AND U38471 ( .A(n907), .B(n38875), .Z(n38874) );
  XOR U38472 ( .A(n38876), .B(n38873), .Z(n38875) );
  XOR U38473 ( .A(n38701), .B(n38869), .Z(n38871) );
  XOR U38474 ( .A(n38877), .B(n38878), .Z(n38701) );
  AND U38475 ( .A(n915), .B(n38837), .Z(n38878) );
  XOR U38476 ( .A(n38877), .B(n38835), .Z(n38837) );
  XOR U38477 ( .A(n38879), .B(n38880), .Z(n38869) );
  AND U38478 ( .A(n38881), .B(n38882), .Z(n38880) );
  XNOR U38479 ( .A(n38879), .B(n38725), .Z(n38882) );
  IV U38480 ( .A(n38728), .Z(n38725) );
  XOR U38481 ( .A(n38883), .B(n38884), .Z(n38728) );
  AND U38482 ( .A(n907), .B(n38885), .Z(n38884) );
  XNOR U38483 ( .A(n38886), .B(n38883), .Z(n38885) );
  XOR U38484 ( .A(n38729), .B(n38879), .Z(n38881) );
  XOR U38485 ( .A(n38887), .B(n38888), .Z(n38729) );
  AND U38486 ( .A(n915), .B(n38846), .Z(n38888) );
  XOR U38487 ( .A(n38887), .B(n38844), .Z(n38846) );
  XOR U38488 ( .A(n38803), .B(n38889), .Z(n38879) );
  AND U38489 ( .A(n38805), .B(n38890), .Z(n38889) );
  XNOR U38490 ( .A(n38803), .B(n38774), .Z(n38890) );
  IV U38491 ( .A(n38777), .Z(n38774) );
  XOR U38492 ( .A(n38891), .B(n38892), .Z(n38777) );
  AND U38493 ( .A(n907), .B(n38893), .Z(n38892) );
  XOR U38494 ( .A(n38894), .B(n38891), .Z(n38893) );
  XOR U38495 ( .A(n38778), .B(n38803), .Z(n38805) );
  XOR U38496 ( .A(n38895), .B(n38896), .Z(n38778) );
  AND U38497 ( .A(n915), .B(n38856), .Z(n38896) );
  XOR U38498 ( .A(n38895), .B(n38854), .Z(n38856) );
  AND U38499 ( .A(n38857), .B(n38787), .Z(n38803) );
  XNOR U38500 ( .A(n38897), .B(n38898), .Z(n38787) );
  AND U38501 ( .A(n907), .B(n38899), .Z(n38898) );
  XNOR U38502 ( .A(n38900), .B(n38897), .Z(n38899) );
  XNOR U38503 ( .A(n38901), .B(n38902), .Z(n907) );
  AND U38504 ( .A(n38903), .B(n38904), .Z(n38902) );
  XOR U38505 ( .A(n38866), .B(n38901), .Z(n38904) );
  AND U38506 ( .A(n38905), .B(n38906), .Z(n38866) );
  XNOR U38507 ( .A(n38863), .B(n38901), .Z(n38903) );
  XNOR U38508 ( .A(n38907), .B(n38908), .Z(n38863) );
  AND U38509 ( .A(n911), .B(n38909), .Z(n38908) );
  XNOR U38510 ( .A(n38910), .B(n38911), .Z(n38909) );
  XOR U38511 ( .A(n38912), .B(n38913), .Z(n38901) );
  AND U38512 ( .A(n38914), .B(n38915), .Z(n38913) );
  XNOR U38513 ( .A(n38912), .B(n38905), .Z(n38915) );
  IV U38514 ( .A(n38876), .Z(n38905) );
  XOR U38515 ( .A(n38916), .B(n38917), .Z(n38876) );
  XOR U38516 ( .A(n38918), .B(n38906), .Z(n38917) );
  AND U38517 ( .A(n38886), .B(n38919), .Z(n38906) );
  AND U38518 ( .A(n38920), .B(n38921), .Z(n38918) );
  XOR U38519 ( .A(n38922), .B(n38916), .Z(n38920) );
  XNOR U38520 ( .A(n38873), .B(n38912), .Z(n38914) );
  XNOR U38521 ( .A(n38923), .B(n38924), .Z(n38873) );
  AND U38522 ( .A(n911), .B(n38925), .Z(n38924) );
  XNOR U38523 ( .A(n38926), .B(n38927), .Z(n38925) );
  XOR U38524 ( .A(n38928), .B(n38929), .Z(n38912) );
  AND U38525 ( .A(n38930), .B(n38931), .Z(n38929) );
  XNOR U38526 ( .A(n38928), .B(n38886), .Z(n38931) );
  XOR U38527 ( .A(n38932), .B(n38921), .Z(n38886) );
  XNOR U38528 ( .A(n38933), .B(n38916), .Z(n38921) );
  XOR U38529 ( .A(n38934), .B(n38935), .Z(n38916) );
  AND U38530 ( .A(n38936), .B(n38937), .Z(n38935) );
  XOR U38531 ( .A(n38938), .B(n38934), .Z(n38936) );
  XNOR U38532 ( .A(n38939), .B(n38940), .Z(n38933) );
  AND U38533 ( .A(n38941), .B(n38942), .Z(n38940) );
  XOR U38534 ( .A(n38939), .B(n38943), .Z(n38941) );
  XNOR U38535 ( .A(n38922), .B(n38919), .Z(n38932) );
  AND U38536 ( .A(n38944), .B(n38945), .Z(n38919) );
  XOR U38537 ( .A(n38946), .B(n38947), .Z(n38922) );
  AND U38538 ( .A(n38948), .B(n38949), .Z(n38947) );
  XOR U38539 ( .A(n38946), .B(n38950), .Z(n38948) );
  XNOR U38540 ( .A(n38883), .B(n38928), .Z(n38930) );
  XNOR U38541 ( .A(n38951), .B(n38952), .Z(n38883) );
  AND U38542 ( .A(n911), .B(n38953), .Z(n38952) );
  XNOR U38543 ( .A(n38954), .B(n38955), .Z(n38953) );
  XOR U38544 ( .A(n38956), .B(n38957), .Z(n38928) );
  AND U38545 ( .A(n38958), .B(n38959), .Z(n38957) );
  XNOR U38546 ( .A(n38956), .B(n38944), .Z(n38959) );
  IV U38547 ( .A(n38894), .Z(n38944) );
  XNOR U38548 ( .A(n38960), .B(n38937), .Z(n38894) );
  XNOR U38549 ( .A(n38961), .B(n38943), .Z(n38937) );
  XOR U38550 ( .A(n38962), .B(n38963), .Z(n38943) );
  NOR U38551 ( .A(n38964), .B(n38965), .Z(n38963) );
  XNOR U38552 ( .A(n38962), .B(n38966), .Z(n38964) );
  XNOR U38553 ( .A(n38942), .B(n38934), .Z(n38961) );
  XOR U38554 ( .A(n38967), .B(n38968), .Z(n38934) );
  AND U38555 ( .A(n38969), .B(n38970), .Z(n38968) );
  XNOR U38556 ( .A(n38967), .B(n38971), .Z(n38969) );
  XNOR U38557 ( .A(n38972), .B(n38939), .Z(n38942) );
  XOR U38558 ( .A(n38973), .B(n38974), .Z(n38939) );
  AND U38559 ( .A(n38975), .B(n38976), .Z(n38974) );
  XOR U38560 ( .A(n38973), .B(n38977), .Z(n38975) );
  XNOR U38561 ( .A(n38978), .B(n38979), .Z(n38972) );
  NOR U38562 ( .A(n38980), .B(n38981), .Z(n38979) );
  XOR U38563 ( .A(n38978), .B(n38982), .Z(n38980) );
  XNOR U38564 ( .A(n38938), .B(n38945), .Z(n38960) );
  NOR U38565 ( .A(n38900), .B(n38983), .Z(n38945) );
  XOR U38566 ( .A(n38950), .B(n38949), .Z(n38938) );
  XNOR U38567 ( .A(n38984), .B(n38946), .Z(n38949) );
  XOR U38568 ( .A(n38985), .B(n38986), .Z(n38946) );
  AND U38569 ( .A(n38987), .B(n38988), .Z(n38986) );
  XOR U38570 ( .A(n38985), .B(n38989), .Z(n38987) );
  XNOR U38571 ( .A(n38990), .B(n38991), .Z(n38984) );
  NOR U38572 ( .A(n38992), .B(n38993), .Z(n38991) );
  XNOR U38573 ( .A(n38990), .B(n38994), .Z(n38992) );
  XOR U38574 ( .A(n38995), .B(n38996), .Z(n38950) );
  NOR U38575 ( .A(n38997), .B(n38998), .Z(n38996) );
  XNOR U38576 ( .A(n38995), .B(n38999), .Z(n38997) );
  XNOR U38577 ( .A(n38891), .B(n38956), .Z(n38958) );
  XNOR U38578 ( .A(n39000), .B(n39001), .Z(n38891) );
  AND U38579 ( .A(n911), .B(n39002), .Z(n39001) );
  XNOR U38580 ( .A(n39003), .B(n39004), .Z(n39002) );
  AND U38581 ( .A(n38897), .B(n38900), .Z(n38956) );
  XOR U38582 ( .A(n39005), .B(n38983), .Z(n38900) );
  XNOR U38583 ( .A(p_input[2048]), .B(p_input[704]), .Z(n38983) );
  XOR U38584 ( .A(n38971), .B(n38970), .Z(n39005) );
  XNOR U38585 ( .A(n39006), .B(n38977), .Z(n38970) );
  XNOR U38586 ( .A(n38966), .B(n38965), .Z(n38977) );
  XOR U38587 ( .A(n39007), .B(n38962), .Z(n38965) );
  XNOR U38588 ( .A(n29266), .B(p_input[714]), .Z(n38962) );
  XNOR U38589 ( .A(p_input[2059]), .B(p_input[715]), .Z(n39007) );
  XOR U38590 ( .A(p_input[2060]), .B(p_input[716]), .Z(n38966) );
  XNOR U38591 ( .A(n38976), .B(n38967), .Z(n39006) );
  XNOR U38592 ( .A(n29494), .B(p_input[705]), .Z(n38967) );
  XOR U38593 ( .A(n39008), .B(n38982), .Z(n38976) );
  XNOR U38594 ( .A(p_input[2063]), .B(p_input[719]), .Z(n38982) );
  XOR U38595 ( .A(n38973), .B(n38981), .Z(n39008) );
  XOR U38596 ( .A(n39009), .B(n38978), .Z(n38981) );
  XOR U38597 ( .A(p_input[2061]), .B(p_input[717]), .Z(n38978) );
  XNOR U38598 ( .A(p_input[2062]), .B(p_input[718]), .Z(n39009) );
  XNOR U38599 ( .A(n29036), .B(p_input[713]), .Z(n38973) );
  XNOR U38600 ( .A(n38989), .B(n38988), .Z(n38971) );
  XNOR U38601 ( .A(n39010), .B(n38994), .Z(n38988) );
  XOR U38602 ( .A(p_input[2056]), .B(p_input[712]), .Z(n38994) );
  XOR U38603 ( .A(n38985), .B(n38993), .Z(n39010) );
  XOR U38604 ( .A(n39011), .B(n38990), .Z(n38993) );
  XOR U38605 ( .A(p_input[2054]), .B(p_input[710]), .Z(n38990) );
  XNOR U38606 ( .A(p_input[2055]), .B(p_input[711]), .Z(n39011) );
  XNOR U38607 ( .A(n29039), .B(p_input[706]), .Z(n38985) );
  XNOR U38608 ( .A(n38999), .B(n38998), .Z(n38989) );
  XOR U38609 ( .A(n39012), .B(n38995), .Z(n38998) );
  XOR U38610 ( .A(p_input[2051]), .B(p_input[707]), .Z(n38995) );
  XNOR U38611 ( .A(p_input[2052]), .B(p_input[708]), .Z(n39012) );
  XOR U38612 ( .A(p_input[2053]), .B(p_input[709]), .Z(n38999) );
  XNOR U38613 ( .A(n39013), .B(n39014), .Z(n38897) );
  AND U38614 ( .A(n911), .B(n39015), .Z(n39014) );
  XNOR U38615 ( .A(n39016), .B(n39017), .Z(n911) );
  AND U38616 ( .A(n39018), .B(n39019), .Z(n39017) );
  XOR U38617 ( .A(n38911), .B(n39016), .Z(n39019) );
  XNOR U38618 ( .A(n39020), .B(n39016), .Z(n39018) );
  XOR U38619 ( .A(n39021), .B(n39022), .Z(n39016) );
  AND U38620 ( .A(n39023), .B(n39024), .Z(n39022) );
  XOR U38621 ( .A(n38926), .B(n39021), .Z(n39024) );
  XOR U38622 ( .A(n39021), .B(n38927), .Z(n39023) );
  XOR U38623 ( .A(n39025), .B(n39026), .Z(n39021) );
  AND U38624 ( .A(n39027), .B(n39028), .Z(n39026) );
  XOR U38625 ( .A(n38954), .B(n39025), .Z(n39028) );
  XOR U38626 ( .A(n39025), .B(n38955), .Z(n39027) );
  XOR U38627 ( .A(n39029), .B(n39030), .Z(n39025) );
  AND U38628 ( .A(n39031), .B(n39032), .Z(n39030) );
  XOR U38629 ( .A(n39029), .B(n39003), .Z(n39032) );
  XNOR U38630 ( .A(n39033), .B(n39034), .Z(n38857) );
  AND U38631 ( .A(n915), .B(n39035), .Z(n39034) );
  XNOR U38632 ( .A(n39036), .B(n39037), .Z(n915) );
  AND U38633 ( .A(n39038), .B(n39039), .Z(n39037) );
  XOR U38634 ( .A(n39036), .B(n38867), .Z(n39039) );
  XNOR U38635 ( .A(n39036), .B(n38827), .Z(n39038) );
  XOR U38636 ( .A(n39040), .B(n39041), .Z(n39036) );
  AND U38637 ( .A(n39042), .B(n39043), .Z(n39041) );
  XOR U38638 ( .A(n39040), .B(n38835), .Z(n39042) );
  XOR U38639 ( .A(n39044), .B(n39045), .Z(n38818) );
  AND U38640 ( .A(n919), .B(n39035), .Z(n39045) );
  XNOR U38641 ( .A(n39033), .B(n39044), .Z(n39035) );
  XNOR U38642 ( .A(n39046), .B(n39047), .Z(n919) );
  AND U38643 ( .A(n39048), .B(n39049), .Z(n39047) );
  XNOR U38644 ( .A(n39050), .B(n39046), .Z(n39049) );
  IV U38645 ( .A(n38867), .Z(n39050) );
  XOR U38646 ( .A(n39020), .B(n39051), .Z(n38867) );
  AND U38647 ( .A(n922), .B(n39052), .Z(n39051) );
  XOR U38648 ( .A(n38910), .B(n38907), .Z(n39052) );
  IV U38649 ( .A(n39020), .Z(n38910) );
  XNOR U38650 ( .A(n38827), .B(n39046), .Z(n39048) );
  XOR U38651 ( .A(n39053), .B(n39054), .Z(n38827) );
  AND U38652 ( .A(n938), .B(n39055), .Z(n39054) );
  XOR U38653 ( .A(n39040), .B(n39056), .Z(n39046) );
  AND U38654 ( .A(n39057), .B(n39043), .Z(n39056) );
  XNOR U38655 ( .A(n38877), .B(n39040), .Z(n39043) );
  XOR U38656 ( .A(n38927), .B(n39058), .Z(n38877) );
  AND U38657 ( .A(n922), .B(n39059), .Z(n39058) );
  XOR U38658 ( .A(n38923), .B(n38927), .Z(n39059) );
  XNOR U38659 ( .A(n39060), .B(n39040), .Z(n39057) );
  IV U38660 ( .A(n38835), .Z(n39060) );
  XOR U38661 ( .A(n39061), .B(n39062), .Z(n38835) );
  AND U38662 ( .A(n938), .B(n39063), .Z(n39062) );
  XOR U38663 ( .A(n39064), .B(n39065), .Z(n39040) );
  AND U38664 ( .A(n39066), .B(n39067), .Z(n39065) );
  XNOR U38665 ( .A(n38887), .B(n39064), .Z(n39067) );
  XOR U38666 ( .A(n38955), .B(n39068), .Z(n38887) );
  AND U38667 ( .A(n922), .B(n39069), .Z(n39068) );
  XOR U38668 ( .A(n38951), .B(n38955), .Z(n39069) );
  XOR U38669 ( .A(n39064), .B(n38844), .Z(n39066) );
  XOR U38670 ( .A(n39070), .B(n39071), .Z(n38844) );
  AND U38671 ( .A(n938), .B(n39072), .Z(n39071) );
  XOR U38672 ( .A(n39073), .B(n39074), .Z(n39064) );
  AND U38673 ( .A(n39075), .B(n39076), .Z(n39074) );
  XNOR U38674 ( .A(n39073), .B(n38895), .Z(n39076) );
  XOR U38675 ( .A(n39004), .B(n39077), .Z(n38895) );
  AND U38676 ( .A(n922), .B(n39078), .Z(n39077) );
  XOR U38677 ( .A(n39000), .B(n39004), .Z(n39078) );
  XNOR U38678 ( .A(n39079), .B(n39073), .Z(n39075) );
  IV U38679 ( .A(n38854), .Z(n39079) );
  XOR U38680 ( .A(n39080), .B(n39081), .Z(n38854) );
  AND U38681 ( .A(n938), .B(n39082), .Z(n39081) );
  AND U38682 ( .A(n39044), .B(n39033), .Z(n39073) );
  XNOR U38683 ( .A(n39083), .B(n39084), .Z(n39033) );
  AND U38684 ( .A(n922), .B(n39015), .Z(n39084) );
  XNOR U38685 ( .A(n39013), .B(n39083), .Z(n39015) );
  XNOR U38686 ( .A(n39085), .B(n39086), .Z(n922) );
  AND U38687 ( .A(n39087), .B(n39088), .Z(n39086) );
  XNOR U38688 ( .A(n39085), .B(n38907), .Z(n39088) );
  IV U38689 ( .A(n38911), .Z(n38907) );
  XOR U38690 ( .A(n39089), .B(n39090), .Z(n38911) );
  AND U38691 ( .A(n926), .B(n39091), .Z(n39090) );
  XOR U38692 ( .A(n39092), .B(n39089), .Z(n39091) );
  XNOR U38693 ( .A(n39085), .B(n39020), .Z(n39087) );
  XOR U38694 ( .A(n39093), .B(n39094), .Z(n39020) );
  AND U38695 ( .A(n934), .B(n39055), .Z(n39094) );
  XOR U38696 ( .A(n39053), .B(n39093), .Z(n39055) );
  XOR U38697 ( .A(n39095), .B(n39096), .Z(n39085) );
  AND U38698 ( .A(n39097), .B(n39098), .Z(n39096) );
  XNOR U38699 ( .A(n39095), .B(n38923), .Z(n39098) );
  IV U38700 ( .A(n38926), .Z(n38923) );
  XOR U38701 ( .A(n39099), .B(n39100), .Z(n38926) );
  AND U38702 ( .A(n926), .B(n39101), .Z(n39100) );
  XOR U38703 ( .A(n39102), .B(n39099), .Z(n39101) );
  XOR U38704 ( .A(n38927), .B(n39095), .Z(n39097) );
  XOR U38705 ( .A(n39103), .B(n39104), .Z(n38927) );
  AND U38706 ( .A(n934), .B(n39063), .Z(n39104) );
  XOR U38707 ( .A(n39103), .B(n39061), .Z(n39063) );
  XOR U38708 ( .A(n39105), .B(n39106), .Z(n39095) );
  AND U38709 ( .A(n39107), .B(n39108), .Z(n39106) );
  XNOR U38710 ( .A(n39105), .B(n38951), .Z(n39108) );
  IV U38711 ( .A(n38954), .Z(n38951) );
  XOR U38712 ( .A(n39109), .B(n39110), .Z(n38954) );
  AND U38713 ( .A(n926), .B(n39111), .Z(n39110) );
  XNOR U38714 ( .A(n39112), .B(n39109), .Z(n39111) );
  XOR U38715 ( .A(n38955), .B(n39105), .Z(n39107) );
  XOR U38716 ( .A(n39113), .B(n39114), .Z(n38955) );
  AND U38717 ( .A(n934), .B(n39072), .Z(n39114) );
  XOR U38718 ( .A(n39113), .B(n39070), .Z(n39072) );
  XOR U38719 ( .A(n39029), .B(n39115), .Z(n39105) );
  AND U38720 ( .A(n39031), .B(n39116), .Z(n39115) );
  XNOR U38721 ( .A(n39029), .B(n39000), .Z(n39116) );
  IV U38722 ( .A(n39003), .Z(n39000) );
  XOR U38723 ( .A(n39117), .B(n39118), .Z(n39003) );
  AND U38724 ( .A(n926), .B(n39119), .Z(n39118) );
  XOR U38725 ( .A(n39120), .B(n39117), .Z(n39119) );
  XOR U38726 ( .A(n39004), .B(n39029), .Z(n39031) );
  XOR U38727 ( .A(n39121), .B(n39122), .Z(n39004) );
  AND U38728 ( .A(n934), .B(n39082), .Z(n39122) );
  XOR U38729 ( .A(n39121), .B(n39080), .Z(n39082) );
  AND U38730 ( .A(n39083), .B(n39013), .Z(n39029) );
  XNOR U38731 ( .A(n39123), .B(n39124), .Z(n39013) );
  AND U38732 ( .A(n926), .B(n39125), .Z(n39124) );
  XNOR U38733 ( .A(n39126), .B(n39123), .Z(n39125) );
  XNOR U38734 ( .A(n39127), .B(n39128), .Z(n926) );
  AND U38735 ( .A(n39129), .B(n39130), .Z(n39128) );
  XOR U38736 ( .A(n39092), .B(n39127), .Z(n39130) );
  AND U38737 ( .A(n39131), .B(n39132), .Z(n39092) );
  XNOR U38738 ( .A(n39089), .B(n39127), .Z(n39129) );
  XNOR U38739 ( .A(n39133), .B(n39134), .Z(n39089) );
  AND U38740 ( .A(n930), .B(n39135), .Z(n39134) );
  XNOR U38741 ( .A(n39136), .B(n39137), .Z(n39135) );
  XOR U38742 ( .A(n39138), .B(n39139), .Z(n39127) );
  AND U38743 ( .A(n39140), .B(n39141), .Z(n39139) );
  XNOR U38744 ( .A(n39138), .B(n39131), .Z(n39141) );
  IV U38745 ( .A(n39102), .Z(n39131) );
  XOR U38746 ( .A(n39142), .B(n39143), .Z(n39102) );
  XOR U38747 ( .A(n39144), .B(n39132), .Z(n39143) );
  AND U38748 ( .A(n39112), .B(n39145), .Z(n39132) );
  AND U38749 ( .A(n39146), .B(n39147), .Z(n39144) );
  XOR U38750 ( .A(n39148), .B(n39142), .Z(n39146) );
  XNOR U38751 ( .A(n39099), .B(n39138), .Z(n39140) );
  XNOR U38752 ( .A(n39149), .B(n39150), .Z(n39099) );
  AND U38753 ( .A(n930), .B(n39151), .Z(n39150) );
  XNOR U38754 ( .A(n39152), .B(n39153), .Z(n39151) );
  XOR U38755 ( .A(n39154), .B(n39155), .Z(n39138) );
  AND U38756 ( .A(n39156), .B(n39157), .Z(n39155) );
  XNOR U38757 ( .A(n39154), .B(n39112), .Z(n39157) );
  XOR U38758 ( .A(n39158), .B(n39147), .Z(n39112) );
  XNOR U38759 ( .A(n39159), .B(n39142), .Z(n39147) );
  XOR U38760 ( .A(n39160), .B(n39161), .Z(n39142) );
  AND U38761 ( .A(n39162), .B(n39163), .Z(n39161) );
  XOR U38762 ( .A(n39164), .B(n39160), .Z(n39162) );
  XNOR U38763 ( .A(n39165), .B(n39166), .Z(n39159) );
  AND U38764 ( .A(n39167), .B(n39168), .Z(n39166) );
  XOR U38765 ( .A(n39165), .B(n39169), .Z(n39167) );
  XNOR U38766 ( .A(n39148), .B(n39145), .Z(n39158) );
  AND U38767 ( .A(n39170), .B(n39171), .Z(n39145) );
  XOR U38768 ( .A(n39172), .B(n39173), .Z(n39148) );
  AND U38769 ( .A(n39174), .B(n39175), .Z(n39173) );
  XOR U38770 ( .A(n39172), .B(n39176), .Z(n39174) );
  XNOR U38771 ( .A(n39109), .B(n39154), .Z(n39156) );
  XNOR U38772 ( .A(n39177), .B(n39178), .Z(n39109) );
  AND U38773 ( .A(n930), .B(n39179), .Z(n39178) );
  XNOR U38774 ( .A(n39180), .B(n39181), .Z(n39179) );
  XOR U38775 ( .A(n39182), .B(n39183), .Z(n39154) );
  AND U38776 ( .A(n39184), .B(n39185), .Z(n39183) );
  XNOR U38777 ( .A(n39182), .B(n39170), .Z(n39185) );
  IV U38778 ( .A(n39120), .Z(n39170) );
  XNOR U38779 ( .A(n39186), .B(n39163), .Z(n39120) );
  XNOR U38780 ( .A(n39187), .B(n39169), .Z(n39163) );
  XOR U38781 ( .A(n39188), .B(n39189), .Z(n39169) );
  NOR U38782 ( .A(n39190), .B(n39191), .Z(n39189) );
  XNOR U38783 ( .A(n39188), .B(n39192), .Z(n39190) );
  XNOR U38784 ( .A(n39168), .B(n39160), .Z(n39187) );
  XOR U38785 ( .A(n39193), .B(n39194), .Z(n39160) );
  AND U38786 ( .A(n39195), .B(n39196), .Z(n39194) );
  XNOR U38787 ( .A(n39193), .B(n39197), .Z(n39195) );
  XNOR U38788 ( .A(n39198), .B(n39165), .Z(n39168) );
  XOR U38789 ( .A(n39199), .B(n39200), .Z(n39165) );
  AND U38790 ( .A(n39201), .B(n39202), .Z(n39200) );
  XOR U38791 ( .A(n39199), .B(n39203), .Z(n39201) );
  XNOR U38792 ( .A(n39204), .B(n39205), .Z(n39198) );
  NOR U38793 ( .A(n39206), .B(n39207), .Z(n39205) );
  XOR U38794 ( .A(n39204), .B(n39208), .Z(n39206) );
  XNOR U38795 ( .A(n39164), .B(n39171), .Z(n39186) );
  NOR U38796 ( .A(n39126), .B(n39209), .Z(n39171) );
  XOR U38797 ( .A(n39176), .B(n39175), .Z(n39164) );
  XNOR U38798 ( .A(n39210), .B(n39172), .Z(n39175) );
  XOR U38799 ( .A(n39211), .B(n39212), .Z(n39172) );
  AND U38800 ( .A(n39213), .B(n39214), .Z(n39212) );
  XOR U38801 ( .A(n39211), .B(n39215), .Z(n39213) );
  XNOR U38802 ( .A(n39216), .B(n39217), .Z(n39210) );
  NOR U38803 ( .A(n39218), .B(n39219), .Z(n39217) );
  XNOR U38804 ( .A(n39216), .B(n39220), .Z(n39218) );
  XOR U38805 ( .A(n39221), .B(n39222), .Z(n39176) );
  NOR U38806 ( .A(n39223), .B(n39224), .Z(n39222) );
  XNOR U38807 ( .A(n39221), .B(n39225), .Z(n39223) );
  XNOR U38808 ( .A(n39117), .B(n39182), .Z(n39184) );
  XNOR U38809 ( .A(n39226), .B(n39227), .Z(n39117) );
  AND U38810 ( .A(n930), .B(n39228), .Z(n39227) );
  XNOR U38811 ( .A(n39229), .B(n39230), .Z(n39228) );
  AND U38812 ( .A(n39123), .B(n39126), .Z(n39182) );
  XOR U38813 ( .A(n39231), .B(n39209), .Z(n39126) );
  XNOR U38814 ( .A(p_input[2048]), .B(p_input[720]), .Z(n39209) );
  XOR U38815 ( .A(n39197), .B(n39196), .Z(n39231) );
  XNOR U38816 ( .A(n39232), .B(n39203), .Z(n39196) );
  XNOR U38817 ( .A(n39192), .B(n39191), .Z(n39203) );
  XOR U38818 ( .A(n39233), .B(n39188), .Z(n39191) );
  XNOR U38819 ( .A(n29266), .B(p_input[730]), .Z(n39188) );
  XNOR U38820 ( .A(p_input[2059]), .B(p_input[731]), .Z(n39233) );
  XOR U38821 ( .A(p_input[2060]), .B(p_input[732]), .Z(n39192) );
  XNOR U38822 ( .A(n39202), .B(n39193), .Z(n39232) );
  XNOR U38823 ( .A(n29494), .B(p_input[721]), .Z(n39193) );
  XOR U38824 ( .A(n39234), .B(n39208), .Z(n39202) );
  XNOR U38825 ( .A(p_input[2063]), .B(p_input[735]), .Z(n39208) );
  XOR U38826 ( .A(n39199), .B(n39207), .Z(n39234) );
  XOR U38827 ( .A(n39235), .B(n39204), .Z(n39207) );
  XOR U38828 ( .A(p_input[2061]), .B(p_input[733]), .Z(n39204) );
  XNOR U38829 ( .A(p_input[2062]), .B(p_input[734]), .Z(n39235) );
  XNOR U38830 ( .A(n29036), .B(p_input[729]), .Z(n39199) );
  XNOR U38831 ( .A(n39215), .B(n39214), .Z(n39197) );
  XNOR U38832 ( .A(n39236), .B(n39220), .Z(n39214) );
  XOR U38833 ( .A(p_input[2056]), .B(p_input[728]), .Z(n39220) );
  XOR U38834 ( .A(n39211), .B(n39219), .Z(n39236) );
  XOR U38835 ( .A(n39237), .B(n39216), .Z(n39219) );
  XOR U38836 ( .A(p_input[2054]), .B(p_input[726]), .Z(n39216) );
  XNOR U38837 ( .A(p_input[2055]), .B(p_input[727]), .Z(n39237) );
  XNOR U38838 ( .A(n29039), .B(p_input[722]), .Z(n39211) );
  XNOR U38839 ( .A(n39225), .B(n39224), .Z(n39215) );
  XOR U38840 ( .A(n39238), .B(n39221), .Z(n39224) );
  XOR U38841 ( .A(p_input[2051]), .B(p_input[723]), .Z(n39221) );
  XNOR U38842 ( .A(p_input[2052]), .B(p_input[724]), .Z(n39238) );
  XOR U38843 ( .A(p_input[2053]), .B(p_input[725]), .Z(n39225) );
  XNOR U38844 ( .A(n39239), .B(n39240), .Z(n39123) );
  AND U38845 ( .A(n930), .B(n39241), .Z(n39240) );
  XNOR U38846 ( .A(n39242), .B(n39243), .Z(n930) );
  AND U38847 ( .A(n39244), .B(n39245), .Z(n39243) );
  XOR U38848 ( .A(n39137), .B(n39242), .Z(n39245) );
  XNOR U38849 ( .A(n39246), .B(n39242), .Z(n39244) );
  XOR U38850 ( .A(n39247), .B(n39248), .Z(n39242) );
  AND U38851 ( .A(n39249), .B(n39250), .Z(n39248) );
  XOR U38852 ( .A(n39152), .B(n39247), .Z(n39250) );
  XOR U38853 ( .A(n39247), .B(n39153), .Z(n39249) );
  XOR U38854 ( .A(n39251), .B(n39252), .Z(n39247) );
  AND U38855 ( .A(n39253), .B(n39254), .Z(n39252) );
  XOR U38856 ( .A(n39180), .B(n39251), .Z(n39254) );
  XOR U38857 ( .A(n39251), .B(n39181), .Z(n39253) );
  XOR U38858 ( .A(n39255), .B(n39256), .Z(n39251) );
  AND U38859 ( .A(n39257), .B(n39258), .Z(n39256) );
  XOR U38860 ( .A(n39255), .B(n39229), .Z(n39258) );
  XNOR U38861 ( .A(n39259), .B(n39260), .Z(n39083) );
  AND U38862 ( .A(n934), .B(n39261), .Z(n39260) );
  XNOR U38863 ( .A(n39262), .B(n39263), .Z(n934) );
  AND U38864 ( .A(n39264), .B(n39265), .Z(n39263) );
  XOR U38865 ( .A(n39262), .B(n39093), .Z(n39265) );
  XNOR U38866 ( .A(n39262), .B(n39053), .Z(n39264) );
  XOR U38867 ( .A(n39266), .B(n39267), .Z(n39262) );
  AND U38868 ( .A(n39268), .B(n39269), .Z(n39267) );
  XOR U38869 ( .A(n39266), .B(n39061), .Z(n39268) );
  XOR U38870 ( .A(n39270), .B(n39271), .Z(n39044) );
  AND U38871 ( .A(n938), .B(n39261), .Z(n39271) );
  XNOR U38872 ( .A(n39259), .B(n39270), .Z(n39261) );
  XNOR U38873 ( .A(n39272), .B(n39273), .Z(n938) );
  AND U38874 ( .A(n39274), .B(n39275), .Z(n39273) );
  XNOR U38875 ( .A(n39276), .B(n39272), .Z(n39275) );
  IV U38876 ( .A(n39093), .Z(n39276) );
  XOR U38877 ( .A(n39246), .B(n39277), .Z(n39093) );
  AND U38878 ( .A(n941), .B(n39278), .Z(n39277) );
  XOR U38879 ( .A(n39136), .B(n39133), .Z(n39278) );
  IV U38880 ( .A(n39246), .Z(n39136) );
  XNOR U38881 ( .A(n39053), .B(n39272), .Z(n39274) );
  XOR U38882 ( .A(n39279), .B(n39280), .Z(n39053) );
  AND U38883 ( .A(n957), .B(n39281), .Z(n39280) );
  XOR U38884 ( .A(n39266), .B(n39282), .Z(n39272) );
  AND U38885 ( .A(n39283), .B(n39269), .Z(n39282) );
  XNOR U38886 ( .A(n39103), .B(n39266), .Z(n39269) );
  XOR U38887 ( .A(n39153), .B(n39284), .Z(n39103) );
  AND U38888 ( .A(n941), .B(n39285), .Z(n39284) );
  XOR U38889 ( .A(n39149), .B(n39153), .Z(n39285) );
  XNOR U38890 ( .A(n39286), .B(n39266), .Z(n39283) );
  IV U38891 ( .A(n39061), .Z(n39286) );
  XOR U38892 ( .A(n39287), .B(n39288), .Z(n39061) );
  AND U38893 ( .A(n957), .B(n39289), .Z(n39288) );
  XOR U38894 ( .A(n39290), .B(n39291), .Z(n39266) );
  AND U38895 ( .A(n39292), .B(n39293), .Z(n39291) );
  XNOR U38896 ( .A(n39113), .B(n39290), .Z(n39293) );
  XOR U38897 ( .A(n39181), .B(n39294), .Z(n39113) );
  AND U38898 ( .A(n941), .B(n39295), .Z(n39294) );
  XOR U38899 ( .A(n39177), .B(n39181), .Z(n39295) );
  XOR U38900 ( .A(n39290), .B(n39070), .Z(n39292) );
  XOR U38901 ( .A(n39296), .B(n39297), .Z(n39070) );
  AND U38902 ( .A(n957), .B(n39298), .Z(n39297) );
  XOR U38903 ( .A(n39299), .B(n39300), .Z(n39290) );
  AND U38904 ( .A(n39301), .B(n39302), .Z(n39300) );
  XNOR U38905 ( .A(n39299), .B(n39121), .Z(n39302) );
  XOR U38906 ( .A(n39230), .B(n39303), .Z(n39121) );
  AND U38907 ( .A(n941), .B(n39304), .Z(n39303) );
  XOR U38908 ( .A(n39226), .B(n39230), .Z(n39304) );
  XNOR U38909 ( .A(n39305), .B(n39299), .Z(n39301) );
  IV U38910 ( .A(n39080), .Z(n39305) );
  XOR U38911 ( .A(n39306), .B(n39307), .Z(n39080) );
  AND U38912 ( .A(n957), .B(n39308), .Z(n39307) );
  AND U38913 ( .A(n39270), .B(n39259), .Z(n39299) );
  XNOR U38914 ( .A(n39309), .B(n39310), .Z(n39259) );
  AND U38915 ( .A(n941), .B(n39241), .Z(n39310) );
  XNOR U38916 ( .A(n39239), .B(n39309), .Z(n39241) );
  XNOR U38917 ( .A(n39311), .B(n39312), .Z(n941) );
  AND U38918 ( .A(n39313), .B(n39314), .Z(n39312) );
  XNOR U38919 ( .A(n39311), .B(n39133), .Z(n39314) );
  IV U38920 ( .A(n39137), .Z(n39133) );
  XOR U38921 ( .A(n39315), .B(n39316), .Z(n39137) );
  AND U38922 ( .A(n945), .B(n39317), .Z(n39316) );
  XOR U38923 ( .A(n39318), .B(n39315), .Z(n39317) );
  XNOR U38924 ( .A(n39311), .B(n39246), .Z(n39313) );
  XOR U38925 ( .A(n39319), .B(n39320), .Z(n39246) );
  AND U38926 ( .A(n953), .B(n39281), .Z(n39320) );
  XOR U38927 ( .A(n39279), .B(n39319), .Z(n39281) );
  XOR U38928 ( .A(n39321), .B(n39322), .Z(n39311) );
  AND U38929 ( .A(n39323), .B(n39324), .Z(n39322) );
  XNOR U38930 ( .A(n39321), .B(n39149), .Z(n39324) );
  IV U38931 ( .A(n39152), .Z(n39149) );
  XOR U38932 ( .A(n39325), .B(n39326), .Z(n39152) );
  AND U38933 ( .A(n945), .B(n39327), .Z(n39326) );
  XOR U38934 ( .A(n39328), .B(n39325), .Z(n39327) );
  XOR U38935 ( .A(n39153), .B(n39321), .Z(n39323) );
  XOR U38936 ( .A(n39329), .B(n39330), .Z(n39153) );
  AND U38937 ( .A(n953), .B(n39289), .Z(n39330) );
  XOR U38938 ( .A(n39329), .B(n39287), .Z(n39289) );
  XOR U38939 ( .A(n39331), .B(n39332), .Z(n39321) );
  AND U38940 ( .A(n39333), .B(n39334), .Z(n39332) );
  XNOR U38941 ( .A(n39331), .B(n39177), .Z(n39334) );
  IV U38942 ( .A(n39180), .Z(n39177) );
  XOR U38943 ( .A(n39335), .B(n39336), .Z(n39180) );
  AND U38944 ( .A(n945), .B(n39337), .Z(n39336) );
  XNOR U38945 ( .A(n39338), .B(n39335), .Z(n39337) );
  XOR U38946 ( .A(n39181), .B(n39331), .Z(n39333) );
  XOR U38947 ( .A(n39339), .B(n39340), .Z(n39181) );
  AND U38948 ( .A(n953), .B(n39298), .Z(n39340) );
  XOR U38949 ( .A(n39339), .B(n39296), .Z(n39298) );
  XOR U38950 ( .A(n39255), .B(n39341), .Z(n39331) );
  AND U38951 ( .A(n39257), .B(n39342), .Z(n39341) );
  XNOR U38952 ( .A(n39255), .B(n39226), .Z(n39342) );
  IV U38953 ( .A(n39229), .Z(n39226) );
  XOR U38954 ( .A(n39343), .B(n39344), .Z(n39229) );
  AND U38955 ( .A(n945), .B(n39345), .Z(n39344) );
  XOR U38956 ( .A(n39346), .B(n39343), .Z(n39345) );
  XOR U38957 ( .A(n39230), .B(n39255), .Z(n39257) );
  XOR U38958 ( .A(n39347), .B(n39348), .Z(n39230) );
  AND U38959 ( .A(n953), .B(n39308), .Z(n39348) );
  XOR U38960 ( .A(n39347), .B(n39306), .Z(n39308) );
  AND U38961 ( .A(n39309), .B(n39239), .Z(n39255) );
  XNOR U38962 ( .A(n39349), .B(n39350), .Z(n39239) );
  AND U38963 ( .A(n945), .B(n39351), .Z(n39350) );
  XNOR U38964 ( .A(n39352), .B(n39349), .Z(n39351) );
  XNOR U38965 ( .A(n39353), .B(n39354), .Z(n945) );
  AND U38966 ( .A(n39355), .B(n39356), .Z(n39354) );
  XOR U38967 ( .A(n39318), .B(n39353), .Z(n39356) );
  AND U38968 ( .A(n39357), .B(n39358), .Z(n39318) );
  XNOR U38969 ( .A(n39315), .B(n39353), .Z(n39355) );
  XNOR U38970 ( .A(n39359), .B(n39360), .Z(n39315) );
  AND U38971 ( .A(n949), .B(n39361), .Z(n39360) );
  XNOR U38972 ( .A(n39362), .B(n39363), .Z(n39361) );
  XOR U38973 ( .A(n39364), .B(n39365), .Z(n39353) );
  AND U38974 ( .A(n39366), .B(n39367), .Z(n39365) );
  XNOR U38975 ( .A(n39364), .B(n39357), .Z(n39367) );
  IV U38976 ( .A(n39328), .Z(n39357) );
  XOR U38977 ( .A(n39368), .B(n39369), .Z(n39328) );
  XOR U38978 ( .A(n39370), .B(n39358), .Z(n39369) );
  AND U38979 ( .A(n39338), .B(n39371), .Z(n39358) );
  AND U38980 ( .A(n39372), .B(n39373), .Z(n39370) );
  XOR U38981 ( .A(n39374), .B(n39368), .Z(n39372) );
  XNOR U38982 ( .A(n39325), .B(n39364), .Z(n39366) );
  XNOR U38983 ( .A(n39375), .B(n39376), .Z(n39325) );
  AND U38984 ( .A(n949), .B(n39377), .Z(n39376) );
  XNOR U38985 ( .A(n39378), .B(n39379), .Z(n39377) );
  XOR U38986 ( .A(n39380), .B(n39381), .Z(n39364) );
  AND U38987 ( .A(n39382), .B(n39383), .Z(n39381) );
  XNOR U38988 ( .A(n39380), .B(n39338), .Z(n39383) );
  XOR U38989 ( .A(n39384), .B(n39373), .Z(n39338) );
  XNOR U38990 ( .A(n39385), .B(n39368), .Z(n39373) );
  XOR U38991 ( .A(n39386), .B(n39387), .Z(n39368) );
  AND U38992 ( .A(n39388), .B(n39389), .Z(n39387) );
  XOR U38993 ( .A(n39390), .B(n39386), .Z(n39388) );
  XNOR U38994 ( .A(n39391), .B(n39392), .Z(n39385) );
  AND U38995 ( .A(n39393), .B(n39394), .Z(n39392) );
  XOR U38996 ( .A(n39391), .B(n39395), .Z(n39393) );
  XNOR U38997 ( .A(n39374), .B(n39371), .Z(n39384) );
  AND U38998 ( .A(n39396), .B(n39397), .Z(n39371) );
  XOR U38999 ( .A(n39398), .B(n39399), .Z(n39374) );
  AND U39000 ( .A(n39400), .B(n39401), .Z(n39399) );
  XOR U39001 ( .A(n39398), .B(n39402), .Z(n39400) );
  XNOR U39002 ( .A(n39335), .B(n39380), .Z(n39382) );
  XNOR U39003 ( .A(n39403), .B(n39404), .Z(n39335) );
  AND U39004 ( .A(n949), .B(n39405), .Z(n39404) );
  XNOR U39005 ( .A(n39406), .B(n39407), .Z(n39405) );
  XOR U39006 ( .A(n39408), .B(n39409), .Z(n39380) );
  AND U39007 ( .A(n39410), .B(n39411), .Z(n39409) );
  XNOR U39008 ( .A(n39408), .B(n39396), .Z(n39411) );
  IV U39009 ( .A(n39346), .Z(n39396) );
  XNOR U39010 ( .A(n39412), .B(n39389), .Z(n39346) );
  XNOR U39011 ( .A(n39413), .B(n39395), .Z(n39389) );
  XOR U39012 ( .A(n39414), .B(n39415), .Z(n39395) );
  NOR U39013 ( .A(n39416), .B(n39417), .Z(n39415) );
  XNOR U39014 ( .A(n39414), .B(n39418), .Z(n39416) );
  XNOR U39015 ( .A(n39394), .B(n39386), .Z(n39413) );
  XOR U39016 ( .A(n39419), .B(n39420), .Z(n39386) );
  AND U39017 ( .A(n39421), .B(n39422), .Z(n39420) );
  XNOR U39018 ( .A(n39419), .B(n39423), .Z(n39421) );
  XNOR U39019 ( .A(n39424), .B(n39391), .Z(n39394) );
  XOR U39020 ( .A(n39425), .B(n39426), .Z(n39391) );
  AND U39021 ( .A(n39427), .B(n39428), .Z(n39426) );
  XOR U39022 ( .A(n39425), .B(n39429), .Z(n39427) );
  XNOR U39023 ( .A(n39430), .B(n39431), .Z(n39424) );
  NOR U39024 ( .A(n39432), .B(n39433), .Z(n39431) );
  XOR U39025 ( .A(n39430), .B(n39434), .Z(n39432) );
  XNOR U39026 ( .A(n39390), .B(n39397), .Z(n39412) );
  NOR U39027 ( .A(n39352), .B(n39435), .Z(n39397) );
  XOR U39028 ( .A(n39402), .B(n39401), .Z(n39390) );
  XNOR U39029 ( .A(n39436), .B(n39398), .Z(n39401) );
  XOR U39030 ( .A(n39437), .B(n39438), .Z(n39398) );
  AND U39031 ( .A(n39439), .B(n39440), .Z(n39438) );
  XOR U39032 ( .A(n39437), .B(n39441), .Z(n39439) );
  XNOR U39033 ( .A(n39442), .B(n39443), .Z(n39436) );
  NOR U39034 ( .A(n39444), .B(n39445), .Z(n39443) );
  XNOR U39035 ( .A(n39442), .B(n39446), .Z(n39444) );
  XOR U39036 ( .A(n39447), .B(n39448), .Z(n39402) );
  NOR U39037 ( .A(n39449), .B(n39450), .Z(n39448) );
  XNOR U39038 ( .A(n39447), .B(n39451), .Z(n39449) );
  XNOR U39039 ( .A(n39343), .B(n39408), .Z(n39410) );
  XNOR U39040 ( .A(n39452), .B(n39453), .Z(n39343) );
  AND U39041 ( .A(n949), .B(n39454), .Z(n39453) );
  XNOR U39042 ( .A(n39455), .B(n39456), .Z(n39454) );
  AND U39043 ( .A(n39349), .B(n39352), .Z(n39408) );
  XOR U39044 ( .A(n39457), .B(n39435), .Z(n39352) );
  XNOR U39045 ( .A(p_input[2048]), .B(p_input[736]), .Z(n39435) );
  XOR U39046 ( .A(n39423), .B(n39422), .Z(n39457) );
  XNOR U39047 ( .A(n39458), .B(n39429), .Z(n39422) );
  XNOR U39048 ( .A(n39418), .B(n39417), .Z(n39429) );
  XOR U39049 ( .A(n39459), .B(n39414), .Z(n39417) );
  XNOR U39050 ( .A(n29266), .B(p_input[746]), .Z(n39414) );
  XNOR U39051 ( .A(p_input[2059]), .B(p_input[747]), .Z(n39459) );
  XOR U39052 ( .A(p_input[2060]), .B(p_input[748]), .Z(n39418) );
  XNOR U39053 ( .A(n39428), .B(n39419), .Z(n39458) );
  XNOR U39054 ( .A(n29494), .B(p_input[737]), .Z(n39419) );
  XOR U39055 ( .A(n39460), .B(n39434), .Z(n39428) );
  XNOR U39056 ( .A(p_input[2063]), .B(p_input[751]), .Z(n39434) );
  XOR U39057 ( .A(n39425), .B(n39433), .Z(n39460) );
  XOR U39058 ( .A(n39461), .B(n39430), .Z(n39433) );
  XOR U39059 ( .A(p_input[2061]), .B(p_input[749]), .Z(n39430) );
  XNOR U39060 ( .A(p_input[2062]), .B(p_input[750]), .Z(n39461) );
  XNOR U39061 ( .A(n29036), .B(p_input[745]), .Z(n39425) );
  XNOR U39062 ( .A(n39441), .B(n39440), .Z(n39423) );
  XNOR U39063 ( .A(n39462), .B(n39446), .Z(n39440) );
  XOR U39064 ( .A(p_input[2056]), .B(p_input[744]), .Z(n39446) );
  XOR U39065 ( .A(n39437), .B(n39445), .Z(n39462) );
  XOR U39066 ( .A(n39463), .B(n39442), .Z(n39445) );
  XOR U39067 ( .A(p_input[2054]), .B(p_input[742]), .Z(n39442) );
  XNOR U39068 ( .A(p_input[2055]), .B(p_input[743]), .Z(n39463) );
  XNOR U39069 ( .A(n29039), .B(p_input[738]), .Z(n39437) );
  XNOR U39070 ( .A(n39451), .B(n39450), .Z(n39441) );
  XOR U39071 ( .A(n39464), .B(n39447), .Z(n39450) );
  XOR U39072 ( .A(p_input[2051]), .B(p_input[739]), .Z(n39447) );
  XNOR U39073 ( .A(p_input[2052]), .B(p_input[740]), .Z(n39464) );
  XOR U39074 ( .A(p_input[2053]), .B(p_input[741]), .Z(n39451) );
  XNOR U39075 ( .A(n39465), .B(n39466), .Z(n39349) );
  AND U39076 ( .A(n949), .B(n39467), .Z(n39466) );
  XNOR U39077 ( .A(n39468), .B(n39469), .Z(n949) );
  AND U39078 ( .A(n39470), .B(n39471), .Z(n39469) );
  XOR U39079 ( .A(n39363), .B(n39468), .Z(n39471) );
  XNOR U39080 ( .A(n39472), .B(n39468), .Z(n39470) );
  XOR U39081 ( .A(n39473), .B(n39474), .Z(n39468) );
  AND U39082 ( .A(n39475), .B(n39476), .Z(n39474) );
  XOR U39083 ( .A(n39378), .B(n39473), .Z(n39476) );
  XOR U39084 ( .A(n39473), .B(n39379), .Z(n39475) );
  XOR U39085 ( .A(n39477), .B(n39478), .Z(n39473) );
  AND U39086 ( .A(n39479), .B(n39480), .Z(n39478) );
  XOR U39087 ( .A(n39406), .B(n39477), .Z(n39480) );
  XOR U39088 ( .A(n39477), .B(n39407), .Z(n39479) );
  XOR U39089 ( .A(n39481), .B(n39482), .Z(n39477) );
  AND U39090 ( .A(n39483), .B(n39484), .Z(n39482) );
  XOR U39091 ( .A(n39481), .B(n39455), .Z(n39484) );
  XNOR U39092 ( .A(n39485), .B(n39486), .Z(n39309) );
  AND U39093 ( .A(n953), .B(n39487), .Z(n39486) );
  XNOR U39094 ( .A(n39488), .B(n39489), .Z(n953) );
  AND U39095 ( .A(n39490), .B(n39491), .Z(n39489) );
  XOR U39096 ( .A(n39488), .B(n39319), .Z(n39491) );
  XNOR U39097 ( .A(n39488), .B(n39279), .Z(n39490) );
  XOR U39098 ( .A(n39492), .B(n39493), .Z(n39488) );
  AND U39099 ( .A(n39494), .B(n39495), .Z(n39493) );
  XOR U39100 ( .A(n39492), .B(n39287), .Z(n39494) );
  XOR U39101 ( .A(n39496), .B(n39497), .Z(n39270) );
  AND U39102 ( .A(n957), .B(n39487), .Z(n39497) );
  XNOR U39103 ( .A(n39485), .B(n39496), .Z(n39487) );
  XNOR U39104 ( .A(n39498), .B(n39499), .Z(n957) );
  AND U39105 ( .A(n39500), .B(n39501), .Z(n39499) );
  XNOR U39106 ( .A(n39502), .B(n39498), .Z(n39501) );
  IV U39107 ( .A(n39319), .Z(n39502) );
  XOR U39108 ( .A(n39472), .B(n39503), .Z(n39319) );
  AND U39109 ( .A(n960), .B(n39504), .Z(n39503) );
  XOR U39110 ( .A(n39362), .B(n39359), .Z(n39504) );
  IV U39111 ( .A(n39472), .Z(n39362) );
  XNOR U39112 ( .A(n39279), .B(n39498), .Z(n39500) );
  XOR U39113 ( .A(n39505), .B(n39506), .Z(n39279) );
  AND U39114 ( .A(n976), .B(n39507), .Z(n39506) );
  XOR U39115 ( .A(n39492), .B(n39508), .Z(n39498) );
  AND U39116 ( .A(n39509), .B(n39495), .Z(n39508) );
  XNOR U39117 ( .A(n39329), .B(n39492), .Z(n39495) );
  XOR U39118 ( .A(n39379), .B(n39510), .Z(n39329) );
  AND U39119 ( .A(n960), .B(n39511), .Z(n39510) );
  XOR U39120 ( .A(n39375), .B(n39379), .Z(n39511) );
  XNOR U39121 ( .A(n39512), .B(n39492), .Z(n39509) );
  IV U39122 ( .A(n39287), .Z(n39512) );
  XOR U39123 ( .A(n39513), .B(n39514), .Z(n39287) );
  AND U39124 ( .A(n976), .B(n39515), .Z(n39514) );
  XOR U39125 ( .A(n39516), .B(n39517), .Z(n39492) );
  AND U39126 ( .A(n39518), .B(n39519), .Z(n39517) );
  XNOR U39127 ( .A(n39339), .B(n39516), .Z(n39519) );
  XOR U39128 ( .A(n39407), .B(n39520), .Z(n39339) );
  AND U39129 ( .A(n960), .B(n39521), .Z(n39520) );
  XOR U39130 ( .A(n39403), .B(n39407), .Z(n39521) );
  XOR U39131 ( .A(n39516), .B(n39296), .Z(n39518) );
  XOR U39132 ( .A(n39522), .B(n39523), .Z(n39296) );
  AND U39133 ( .A(n976), .B(n39524), .Z(n39523) );
  XOR U39134 ( .A(n39525), .B(n39526), .Z(n39516) );
  AND U39135 ( .A(n39527), .B(n39528), .Z(n39526) );
  XNOR U39136 ( .A(n39525), .B(n39347), .Z(n39528) );
  XOR U39137 ( .A(n39456), .B(n39529), .Z(n39347) );
  AND U39138 ( .A(n960), .B(n39530), .Z(n39529) );
  XOR U39139 ( .A(n39452), .B(n39456), .Z(n39530) );
  XNOR U39140 ( .A(n39531), .B(n39525), .Z(n39527) );
  IV U39141 ( .A(n39306), .Z(n39531) );
  XOR U39142 ( .A(n39532), .B(n39533), .Z(n39306) );
  AND U39143 ( .A(n976), .B(n39534), .Z(n39533) );
  AND U39144 ( .A(n39496), .B(n39485), .Z(n39525) );
  XNOR U39145 ( .A(n39535), .B(n39536), .Z(n39485) );
  AND U39146 ( .A(n960), .B(n39467), .Z(n39536) );
  XNOR U39147 ( .A(n39465), .B(n39535), .Z(n39467) );
  XNOR U39148 ( .A(n39537), .B(n39538), .Z(n960) );
  AND U39149 ( .A(n39539), .B(n39540), .Z(n39538) );
  XNOR U39150 ( .A(n39537), .B(n39359), .Z(n39540) );
  IV U39151 ( .A(n39363), .Z(n39359) );
  XOR U39152 ( .A(n39541), .B(n39542), .Z(n39363) );
  AND U39153 ( .A(n964), .B(n39543), .Z(n39542) );
  XOR U39154 ( .A(n39544), .B(n39541), .Z(n39543) );
  XNOR U39155 ( .A(n39537), .B(n39472), .Z(n39539) );
  XOR U39156 ( .A(n39545), .B(n39546), .Z(n39472) );
  AND U39157 ( .A(n972), .B(n39507), .Z(n39546) );
  XOR U39158 ( .A(n39505), .B(n39545), .Z(n39507) );
  XOR U39159 ( .A(n39547), .B(n39548), .Z(n39537) );
  AND U39160 ( .A(n39549), .B(n39550), .Z(n39548) );
  XNOR U39161 ( .A(n39547), .B(n39375), .Z(n39550) );
  IV U39162 ( .A(n39378), .Z(n39375) );
  XOR U39163 ( .A(n39551), .B(n39552), .Z(n39378) );
  AND U39164 ( .A(n964), .B(n39553), .Z(n39552) );
  XOR U39165 ( .A(n39554), .B(n39551), .Z(n39553) );
  XOR U39166 ( .A(n39379), .B(n39547), .Z(n39549) );
  XOR U39167 ( .A(n39555), .B(n39556), .Z(n39379) );
  AND U39168 ( .A(n972), .B(n39515), .Z(n39556) );
  XOR U39169 ( .A(n39555), .B(n39513), .Z(n39515) );
  XOR U39170 ( .A(n39557), .B(n39558), .Z(n39547) );
  AND U39171 ( .A(n39559), .B(n39560), .Z(n39558) );
  XNOR U39172 ( .A(n39557), .B(n39403), .Z(n39560) );
  IV U39173 ( .A(n39406), .Z(n39403) );
  XOR U39174 ( .A(n39561), .B(n39562), .Z(n39406) );
  AND U39175 ( .A(n964), .B(n39563), .Z(n39562) );
  XNOR U39176 ( .A(n39564), .B(n39561), .Z(n39563) );
  XOR U39177 ( .A(n39407), .B(n39557), .Z(n39559) );
  XOR U39178 ( .A(n39565), .B(n39566), .Z(n39407) );
  AND U39179 ( .A(n972), .B(n39524), .Z(n39566) );
  XOR U39180 ( .A(n39565), .B(n39522), .Z(n39524) );
  XOR U39181 ( .A(n39481), .B(n39567), .Z(n39557) );
  AND U39182 ( .A(n39483), .B(n39568), .Z(n39567) );
  XNOR U39183 ( .A(n39481), .B(n39452), .Z(n39568) );
  IV U39184 ( .A(n39455), .Z(n39452) );
  XOR U39185 ( .A(n39569), .B(n39570), .Z(n39455) );
  AND U39186 ( .A(n964), .B(n39571), .Z(n39570) );
  XOR U39187 ( .A(n39572), .B(n39569), .Z(n39571) );
  XOR U39188 ( .A(n39456), .B(n39481), .Z(n39483) );
  XOR U39189 ( .A(n39573), .B(n39574), .Z(n39456) );
  AND U39190 ( .A(n972), .B(n39534), .Z(n39574) );
  XOR U39191 ( .A(n39573), .B(n39532), .Z(n39534) );
  AND U39192 ( .A(n39535), .B(n39465), .Z(n39481) );
  XNOR U39193 ( .A(n39575), .B(n39576), .Z(n39465) );
  AND U39194 ( .A(n964), .B(n39577), .Z(n39576) );
  XNOR U39195 ( .A(n39578), .B(n39575), .Z(n39577) );
  XNOR U39196 ( .A(n39579), .B(n39580), .Z(n964) );
  AND U39197 ( .A(n39581), .B(n39582), .Z(n39580) );
  XOR U39198 ( .A(n39544), .B(n39579), .Z(n39582) );
  AND U39199 ( .A(n39583), .B(n39584), .Z(n39544) );
  XNOR U39200 ( .A(n39541), .B(n39579), .Z(n39581) );
  XNOR U39201 ( .A(n39585), .B(n39586), .Z(n39541) );
  AND U39202 ( .A(n968), .B(n39587), .Z(n39586) );
  XNOR U39203 ( .A(n39588), .B(n39589), .Z(n39587) );
  XOR U39204 ( .A(n39590), .B(n39591), .Z(n39579) );
  AND U39205 ( .A(n39592), .B(n39593), .Z(n39591) );
  XNOR U39206 ( .A(n39590), .B(n39583), .Z(n39593) );
  IV U39207 ( .A(n39554), .Z(n39583) );
  XOR U39208 ( .A(n39594), .B(n39595), .Z(n39554) );
  XOR U39209 ( .A(n39596), .B(n39584), .Z(n39595) );
  AND U39210 ( .A(n39564), .B(n39597), .Z(n39584) );
  AND U39211 ( .A(n39598), .B(n39599), .Z(n39596) );
  XOR U39212 ( .A(n39600), .B(n39594), .Z(n39598) );
  XNOR U39213 ( .A(n39551), .B(n39590), .Z(n39592) );
  XNOR U39214 ( .A(n39601), .B(n39602), .Z(n39551) );
  AND U39215 ( .A(n968), .B(n39603), .Z(n39602) );
  XNOR U39216 ( .A(n39604), .B(n39605), .Z(n39603) );
  XOR U39217 ( .A(n39606), .B(n39607), .Z(n39590) );
  AND U39218 ( .A(n39608), .B(n39609), .Z(n39607) );
  XNOR U39219 ( .A(n39606), .B(n39564), .Z(n39609) );
  XOR U39220 ( .A(n39610), .B(n39599), .Z(n39564) );
  XNOR U39221 ( .A(n39611), .B(n39594), .Z(n39599) );
  XOR U39222 ( .A(n39612), .B(n39613), .Z(n39594) );
  AND U39223 ( .A(n39614), .B(n39615), .Z(n39613) );
  XOR U39224 ( .A(n39616), .B(n39612), .Z(n39614) );
  XNOR U39225 ( .A(n39617), .B(n39618), .Z(n39611) );
  AND U39226 ( .A(n39619), .B(n39620), .Z(n39618) );
  XOR U39227 ( .A(n39617), .B(n39621), .Z(n39619) );
  XNOR U39228 ( .A(n39600), .B(n39597), .Z(n39610) );
  AND U39229 ( .A(n39622), .B(n39623), .Z(n39597) );
  XOR U39230 ( .A(n39624), .B(n39625), .Z(n39600) );
  AND U39231 ( .A(n39626), .B(n39627), .Z(n39625) );
  XOR U39232 ( .A(n39624), .B(n39628), .Z(n39626) );
  XNOR U39233 ( .A(n39561), .B(n39606), .Z(n39608) );
  XNOR U39234 ( .A(n39629), .B(n39630), .Z(n39561) );
  AND U39235 ( .A(n968), .B(n39631), .Z(n39630) );
  XNOR U39236 ( .A(n39632), .B(n39633), .Z(n39631) );
  XOR U39237 ( .A(n39634), .B(n39635), .Z(n39606) );
  AND U39238 ( .A(n39636), .B(n39637), .Z(n39635) );
  XNOR U39239 ( .A(n39634), .B(n39622), .Z(n39637) );
  IV U39240 ( .A(n39572), .Z(n39622) );
  XNOR U39241 ( .A(n39638), .B(n39615), .Z(n39572) );
  XNOR U39242 ( .A(n39639), .B(n39621), .Z(n39615) );
  XOR U39243 ( .A(n39640), .B(n39641), .Z(n39621) );
  NOR U39244 ( .A(n39642), .B(n39643), .Z(n39641) );
  XNOR U39245 ( .A(n39640), .B(n39644), .Z(n39642) );
  XNOR U39246 ( .A(n39620), .B(n39612), .Z(n39639) );
  XOR U39247 ( .A(n39645), .B(n39646), .Z(n39612) );
  AND U39248 ( .A(n39647), .B(n39648), .Z(n39646) );
  XNOR U39249 ( .A(n39645), .B(n39649), .Z(n39647) );
  XNOR U39250 ( .A(n39650), .B(n39617), .Z(n39620) );
  XOR U39251 ( .A(n39651), .B(n39652), .Z(n39617) );
  AND U39252 ( .A(n39653), .B(n39654), .Z(n39652) );
  XOR U39253 ( .A(n39651), .B(n39655), .Z(n39653) );
  XNOR U39254 ( .A(n39656), .B(n39657), .Z(n39650) );
  NOR U39255 ( .A(n39658), .B(n39659), .Z(n39657) );
  XOR U39256 ( .A(n39656), .B(n39660), .Z(n39658) );
  XNOR U39257 ( .A(n39616), .B(n39623), .Z(n39638) );
  NOR U39258 ( .A(n39578), .B(n39661), .Z(n39623) );
  XOR U39259 ( .A(n39628), .B(n39627), .Z(n39616) );
  XNOR U39260 ( .A(n39662), .B(n39624), .Z(n39627) );
  XOR U39261 ( .A(n39663), .B(n39664), .Z(n39624) );
  AND U39262 ( .A(n39665), .B(n39666), .Z(n39664) );
  XOR U39263 ( .A(n39663), .B(n39667), .Z(n39665) );
  XNOR U39264 ( .A(n39668), .B(n39669), .Z(n39662) );
  NOR U39265 ( .A(n39670), .B(n39671), .Z(n39669) );
  XNOR U39266 ( .A(n39668), .B(n39672), .Z(n39670) );
  XOR U39267 ( .A(n39673), .B(n39674), .Z(n39628) );
  NOR U39268 ( .A(n39675), .B(n39676), .Z(n39674) );
  XNOR U39269 ( .A(n39673), .B(n39677), .Z(n39675) );
  XNOR U39270 ( .A(n39569), .B(n39634), .Z(n39636) );
  XNOR U39271 ( .A(n39678), .B(n39679), .Z(n39569) );
  AND U39272 ( .A(n968), .B(n39680), .Z(n39679) );
  XNOR U39273 ( .A(n39681), .B(n39682), .Z(n39680) );
  AND U39274 ( .A(n39575), .B(n39578), .Z(n39634) );
  XOR U39275 ( .A(n39683), .B(n39661), .Z(n39578) );
  XNOR U39276 ( .A(p_input[2048]), .B(p_input[752]), .Z(n39661) );
  XOR U39277 ( .A(n39649), .B(n39648), .Z(n39683) );
  XNOR U39278 ( .A(n39684), .B(n39655), .Z(n39648) );
  XNOR U39279 ( .A(n39644), .B(n39643), .Z(n39655) );
  XOR U39280 ( .A(n39685), .B(n39640), .Z(n39643) );
  XNOR U39281 ( .A(n29266), .B(p_input[762]), .Z(n39640) );
  XNOR U39282 ( .A(p_input[2059]), .B(p_input[763]), .Z(n39685) );
  XOR U39283 ( .A(p_input[2060]), .B(p_input[764]), .Z(n39644) );
  XNOR U39284 ( .A(n39654), .B(n39645), .Z(n39684) );
  XNOR U39285 ( .A(n29494), .B(p_input[753]), .Z(n39645) );
  XOR U39286 ( .A(n39686), .B(n39660), .Z(n39654) );
  XNOR U39287 ( .A(p_input[2063]), .B(p_input[767]), .Z(n39660) );
  XOR U39288 ( .A(n39651), .B(n39659), .Z(n39686) );
  XOR U39289 ( .A(n39687), .B(n39656), .Z(n39659) );
  XOR U39290 ( .A(p_input[2061]), .B(p_input[765]), .Z(n39656) );
  XNOR U39291 ( .A(p_input[2062]), .B(p_input[766]), .Z(n39687) );
  XNOR U39292 ( .A(n29036), .B(p_input[761]), .Z(n39651) );
  XNOR U39293 ( .A(n39667), .B(n39666), .Z(n39649) );
  XNOR U39294 ( .A(n39688), .B(n39672), .Z(n39666) );
  XOR U39295 ( .A(p_input[2056]), .B(p_input[760]), .Z(n39672) );
  XOR U39296 ( .A(n39663), .B(n39671), .Z(n39688) );
  XOR U39297 ( .A(n39689), .B(n39668), .Z(n39671) );
  XOR U39298 ( .A(p_input[2054]), .B(p_input[758]), .Z(n39668) );
  XNOR U39299 ( .A(p_input[2055]), .B(p_input[759]), .Z(n39689) );
  XNOR U39300 ( .A(n29039), .B(p_input[754]), .Z(n39663) );
  XNOR U39301 ( .A(n39677), .B(n39676), .Z(n39667) );
  XOR U39302 ( .A(n39690), .B(n39673), .Z(n39676) );
  XOR U39303 ( .A(p_input[2051]), .B(p_input[755]), .Z(n39673) );
  XNOR U39304 ( .A(p_input[2052]), .B(p_input[756]), .Z(n39690) );
  XOR U39305 ( .A(p_input[2053]), .B(p_input[757]), .Z(n39677) );
  XNOR U39306 ( .A(n39691), .B(n39692), .Z(n39575) );
  AND U39307 ( .A(n968), .B(n39693), .Z(n39692) );
  XNOR U39308 ( .A(n39694), .B(n39695), .Z(n968) );
  AND U39309 ( .A(n39696), .B(n39697), .Z(n39695) );
  XOR U39310 ( .A(n39589), .B(n39694), .Z(n39697) );
  XNOR U39311 ( .A(n39698), .B(n39694), .Z(n39696) );
  XOR U39312 ( .A(n39699), .B(n39700), .Z(n39694) );
  AND U39313 ( .A(n39701), .B(n39702), .Z(n39700) );
  XOR U39314 ( .A(n39604), .B(n39699), .Z(n39702) );
  XOR U39315 ( .A(n39699), .B(n39605), .Z(n39701) );
  XOR U39316 ( .A(n39703), .B(n39704), .Z(n39699) );
  AND U39317 ( .A(n39705), .B(n39706), .Z(n39704) );
  XOR U39318 ( .A(n39632), .B(n39703), .Z(n39706) );
  XOR U39319 ( .A(n39703), .B(n39633), .Z(n39705) );
  XOR U39320 ( .A(n39707), .B(n39708), .Z(n39703) );
  AND U39321 ( .A(n39709), .B(n39710), .Z(n39708) );
  XOR U39322 ( .A(n39707), .B(n39681), .Z(n39710) );
  XNOR U39323 ( .A(n39711), .B(n39712), .Z(n39535) );
  AND U39324 ( .A(n972), .B(n39713), .Z(n39712) );
  XNOR U39325 ( .A(n39714), .B(n39715), .Z(n972) );
  AND U39326 ( .A(n39716), .B(n39717), .Z(n39715) );
  XOR U39327 ( .A(n39714), .B(n39545), .Z(n39717) );
  XNOR U39328 ( .A(n39714), .B(n39505), .Z(n39716) );
  XOR U39329 ( .A(n39718), .B(n39719), .Z(n39714) );
  AND U39330 ( .A(n39720), .B(n39721), .Z(n39719) );
  XOR U39331 ( .A(n39718), .B(n39513), .Z(n39720) );
  XOR U39332 ( .A(n39722), .B(n39723), .Z(n39496) );
  AND U39333 ( .A(n976), .B(n39713), .Z(n39723) );
  XNOR U39334 ( .A(n39711), .B(n39722), .Z(n39713) );
  XNOR U39335 ( .A(n39724), .B(n39725), .Z(n976) );
  AND U39336 ( .A(n39726), .B(n39727), .Z(n39725) );
  XNOR U39337 ( .A(n39728), .B(n39724), .Z(n39727) );
  IV U39338 ( .A(n39545), .Z(n39728) );
  XOR U39339 ( .A(n39698), .B(n39729), .Z(n39545) );
  AND U39340 ( .A(n979), .B(n39730), .Z(n39729) );
  XOR U39341 ( .A(n39588), .B(n39585), .Z(n39730) );
  IV U39342 ( .A(n39698), .Z(n39588) );
  XNOR U39343 ( .A(n39505), .B(n39724), .Z(n39726) );
  XOR U39344 ( .A(n39731), .B(n39732), .Z(n39505) );
  AND U39345 ( .A(n995), .B(n39733), .Z(n39732) );
  XOR U39346 ( .A(n39718), .B(n39734), .Z(n39724) );
  AND U39347 ( .A(n39735), .B(n39721), .Z(n39734) );
  XNOR U39348 ( .A(n39555), .B(n39718), .Z(n39721) );
  XOR U39349 ( .A(n39605), .B(n39736), .Z(n39555) );
  AND U39350 ( .A(n979), .B(n39737), .Z(n39736) );
  XOR U39351 ( .A(n39601), .B(n39605), .Z(n39737) );
  XNOR U39352 ( .A(n39738), .B(n39718), .Z(n39735) );
  IV U39353 ( .A(n39513), .Z(n39738) );
  XOR U39354 ( .A(n39739), .B(n39740), .Z(n39513) );
  AND U39355 ( .A(n995), .B(n39741), .Z(n39740) );
  XOR U39356 ( .A(n39742), .B(n39743), .Z(n39718) );
  AND U39357 ( .A(n39744), .B(n39745), .Z(n39743) );
  XNOR U39358 ( .A(n39565), .B(n39742), .Z(n39745) );
  XOR U39359 ( .A(n39633), .B(n39746), .Z(n39565) );
  AND U39360 ( .A(n979), .B(n39747), .Z(n39746) );
  XOR U39361 ( .A(n39629), .B(n39633), .Z(n39747) );
  XOR U39362 ( .A(n39742), .B(n39522), .Z(n39744) );
  XOR U39363 ( .A(n39748), .B(n39749), .Z(n39522) );
  AND U39364 ( .A(n995), .B(n39750), .Z(n39749) );
  XOR U39365 ( .A(n39751), .B(n39752), .Z(n39742) );
  AND U39366 ( .A(n39753), .B(n39754), .Z(n39752) );
  XNOR U39367 ( .A(n39751), .B(n39573), .Z(n39754) );
  XOR U39368 ( .A(n39682), .B(n39755), .Z(n39573) );
  AND U39369 ( .A(n979), .B(n39756), .Z(n39755) );
  XOR U39370 ( .A(n39678), .B(n39682), .Z(n39756) );
  XNOR U39371 ( .A(n39757), .B(n39751), .Z(n39753) );
  IV U39372 ( .A(n39532), .Z(n39757) );
  XOR U39373 ( .A(n39758), .B(n39759), .Z(n39532) );
  AND U39374 ( .A(n995), .B(n39760), .Z(n39759) );
  AND U39375 ( .A(n39722), .B(n39711), .Z(n39751) );
  XNOR U39376 ( .A(n39761), .B(n39762), .Z(n39711) );
  AND U39377 ( .A(n979), .B(n39693), .Z(n39762) );
  XNOR U39378 ( .A(n39691), .B(n39761), .Z(n39693) );
  XNOR U39379 ( .A(n39763), .B(n39764), .Z(n979) );
  AND U39380 ( .A(n39765), .B(n39766), .Z(n39764) );
  XNOR U39381 ( .A(n39763), .B(n39585), .Z(n39766) );
  IV U39382 ( .A(n39589), .Z(n39585) );
  XOR U39383 ( .A(n39767), .B(n39768), .Z(n39589) );
  AND U39384 ( .A(n983), .B(n39769), .Z(n39768) );
  XOR U39385 ( .A(n39770), .B(n39767), .Z(n39769) );
  XNOR U39386 ( .A(n39763), .B(n39698), .Z(n39765) );
  XOR U39387 ( .A(n39771), .B(n39772), .Z(n39698) );
  AND U39388 ( .A(n991), .B(n39733), .Z(n39772) );
  XOR U39389 ( .A(n39731), .B(n39771), .Z(n39733) );
  XOR U39390 ( .A(n39773), .B(n39774), .Z(n39763) );
  AND U39391 ( .A(n39775), .B(n39776), .Z(n39774) );
  XNOR U39392 ( .A(n39773), .B(n39601), .Z(n39776) );
  IV U39393 ( .A(n39604), .Z(n39601) );
  XOR U39394 ( .A(n39777), .B(n39778), .Z(n39604) );
  AND U39395 ( .A(n983), .B(n39779), .Z(n39778) );
  XOR U39396 ( .A(n39780), .B(n39777), .Z(n39779) );
  XOR U39397 ( .A(n39605), .B(n39773), .Z(n39775) );
  XOR U39398 ( .A(n39781), .B(n39782), .Z(n39605) );
  AND U39399 ( .A(n991), .B(n39741), .Z(n39782) );
  XOR U39400 ( .A(n39781), .B(n39739), .Z(n39741) );
  XOR U39401 ( .A(n39783), .B(n39784), .Z(n39773) );
  AND U39402 ( .A(n39785), .B(n39786), .Z(n39784) );
  XNOR U39403 ( .A(n39783), .B(n39629), .Z(n39786) );
  IV U39404 ( .A(n39632), .Z(n39629) );
  XOR U39405 ( .A(n39787), .B(n39788), .Z(n39632) );
  AND U39406 ( .A(n983), .B(n39789), .Z(n39788) );
  XNOR U39407 ( .A(n39790), .B(n39787), .Z(n39789) );
  XOR U39408 ( .A(n39633), .B(n39783), .Z(n39785) );
  XOR U39409 ( .A(n39791), .B(n39792), .Z(n39633) );
  AND U39410 ( .A(n991), .B(n39750), .Z(n39792) );
  XOR U39411 ( .A(n39791), .B(n39748), .Z(n39750) );
  XOR U39412 ( .A(n39707), .B(n39793), .Z(n39783) );
  AND U39413 ( .A(n39709), .B(n39794), .Z(n39793) );
  XNOR U39414 ( .A(n39707), .B(n39678), .Z(n39794) );
  IV U39415 ( .A(n39681), .Z(n39678) );
  XOR U39416 ( .A(n39795), .B(n39796), .Z(n39681) );
  AND U39417 ( .A(n983), .B(n39797), .Z(n39796) );
  XOR U39418 ( .A(n39798), .B(n39795), .Z(n39797) );
  XOR U39419 ( .A(n39682), .B(n39707), .Z(n39709) );
  XOR U39420 ( .A(n39799), .B(n39800), .Z(n39682) );
  AND U39421 ( .A(n991), .B(n39760), .Z(n39800) );
  XOR U39422 ( .A(n39799), .B(n39758), .Z(n39760) );
  AND U39423 ( .A(n39761), .B(n39691), .Z(n39707) );
  XNOR U39424 ( .A(n39801), .B(n39802), .Z(n39691) );
  AND U39425 ( .A(n983), .B(n39803), .Z(n39802) );
  XNOR U39426 ( .A(n39804), .B(n39801), .Z(n39803) );
  XNOR U39427 ( .A(n39805), .B(n39806), .Z(n983) );
  AND U39428 ( .A(n39807), .B(n39808), .Z(n39806) );
  XOR U39429 ( .A(n39770), .B(n39805), .Z(n39808) );
  AND U39430 ( .A(n39809), .B(n39810), .Z(n39770) );
  XNOR U39431 ( .A(n39767), .B(n39805), .Z(n39807) );
  XNOR U39432 ( .A(n39811), .B(n39812), .Z(n39767) );
  AND U39433 ( .A(n987), .B(n39813), .Z(n39812) );
  XNOR U39434 ( .A(n39814), .B(n39815), .Z(n39813) );
  XOR U39435 ( .A(n39816), .B(n39817), .Z(n39805) );
  AND U39436 ( .A(n39818), .B(n39819), .Z(n39817) );
  XNOR U39437 ( .A(n39816), .B(n39809), .Z(n39819) );
  IV U39438 ( .A(n39780), .Z(n39809) );
  XOR U39439 ( .A(n39820), .B(n39821), .Z(n39780) );
  XOR U39440 ( .A(n39822), .B(n39810), .Z(n39821) );
  AND U39441 ( .A(n39790), .B(n39823), .Z(n39810) );
  AND U39442 ( .A(n39824), .B(n39825), .Z(n39822) );
  XOR U39443 ( .A(n39826), .B(n39820), .Z(n39824) );
  XNOR U39444 ( .A(n39777), .B(n39816), .Z(n39818) );
  XNOR U39445 ( .A(n39827), .B(n39828), .Z(n39777) );
  AND U39446 ( .A(n987), .B(n39829), .Z(n39828) );
  XNOR U39447 ( .A(n39830), .B(n39831), .Z(n39829) );
  XOR U39448 ( .A(n39832), .B(n39833), .Z(n39816) );
  AND U39449 ( .A(n39834), .B(n39835), .Z(n39833) );
  XNOR U39450 ( .A(n39832), .B(n39790), .Z(n39835) );
  XOR U39451 ( .A(n39836), .B(n39825), .Z(n39790) );
  XNOR U39452 ( .A(n39837), .B(n39820), .Z(n39825) );
  XOR U39453 ( .A(n39838), .B(n39839), .Z(n39820) );
  AND U39454 ( .A(n39840), .B(n39841), .Z(n39839) );
  XOR U39455 ( .A(n39842), .B(n39838), .Z(n39840) );
  XNOR U39456 ( .A(n39843), .B(n39844), .Z(n39837) );
  AND U39457 ( .A(n39845), .B(n39846), .Z(n39844) );
  XOR U39458 ( .A(n39843), .B(n39847), .Z(n39845) );
  XNOR U39459 ( .A(n39826), .B(n39823), .Z(n39836) );
  AND U39460 ( .A(n39848), .B(n39849), .Z(n39823) );
  XOR U39461 ( .A(n39850), .B(n39851), .Z(n39826) );
  AND U39462 ( .A(n39852), .B(n39853), .Z(n39851) );
  XOR U39463 ( .A(n39850), .B(n39854), .Z(n39852) );
  XNOR U39464 ( .A(n39787), .B(n39832), .Z(n39834) );
  XNOR U39465 ( .A(n39855), .B(n39856), .Z(n39787) );
  AND U39466 ( .A(n987), .B(n39857), .Z(n39856) );
  XNOR U39467 ( .A(n39858), .B(n39859), .Z(n39857) );
  XOR U39468 ( .A(n39860), .B(n39861), .Z(n39832) );
  AND U39469 ( .A(n39862), .B(n39863), .Z(n39861) );
  XNOR U39470 ( .A(n39860), .B(n39848), .Z(n39863) );
  IV U39471 ( .A(n39798), .Z(n39848) );
  XNOR U39472 ( .A(n39864), .B(n39841), .Z(n39798) );
  XNOR U39473 ( .A(n39865), .B(n39847), .Z(n39841) );
  XOR U39474 ( .A(n39866), .B(n39867), .Z(n39847) );
  NOR U39475 ( .A(n39868), .B(n39869), .Z(n39867) );
  XNOR U39476 ( .A(n39866), .B(n39870), .Z(n39868) );
  XNOR U39477 ( .A(n39846), .B(n39838), .Z(n39865) );
  XOR U39478 ( .A(n39871), .B(n39872), .Z(n39838) );
  AND U39479 ( .A(n39873), .B(n39874), .Z(n39872) );
  XNOR U39480 ( .A(n39871), .B(n39875), .Z(n39873) );
  XNOR U39481 ( .A(n39876), .B(n39843), .Z(n39846) );
  XOR U39482 ( .A(n39877), .B(n39878), .Z(n39843) );
  AND U39483 ( .A(n39879), .B(n39880), .Z(n39878) );
  XOR U39484 ( .A(n39877), .B(n39881), .Z(n39879) );
  XNOR U39485 ( .A(n39882), .B(n39883), .Z(n39876) );
  NOR U39486 ( .A(n39884), .B(n39885), .Z(n39883) );
  XOR U39487 ( .A(n39882), .B(n39886), .Z(n39884) );
  XNOR U39488 ( .A(n39842), .B(n39849), .Z(n39864) );
  NOR U39489 ( .A(n39804), .B(n39887), .Z(n39849) );
  XOR U39490 ( .A(n39854), .B(n39853), .Z(n39842) );
  XNOR U39491 ( .A(n39888), .B(n39850), .Z(n39853) );
  XOR U39492 ( .A(n39889), .B(n39890), .Z(n39850) );
  AND U39493 ( .A(n39891), .B(n39892), .Z(n39890) );
  XOR U39494 ( .A(n39889), .B(n39893), .Z(n39891) );
  XNOR U39495 ( .A(n39894), .B(n39895), .Z(n39888) );
  NOR U39496 ( .A(n39896), .B(n39897), .Z(n39895) );
  XNOR U39497 ( .A(n39894), .B(n39898), .Z(n39896) );
  XOR U39498 ( .A(n39899), .B(n39900), .Z(n39854) );
  NOR U39499 ( .A(n39901), .B(n39902), .Z(n39900) );
  XNOR U39500 ( .A(n39899), .B(n39903), .Z(n39901) );
  XNOR U39501 ( .A(n39795), .B(n39860), .Z(n39862) );
  XNOR U39502 ( .A(n39904), .B(n39905), .Z(n39795) );
  AND U39503 ( .A(n987), .B(n39906), .Z(n39905) );
  XNOR U39504 ( .A(n39907), .B(n39908), .Z(n39906) );
  AND U39505 ( .A(n39801), .B(n39804), .Z(n39860) );
  XOR U39506 ( .A(n39909), .B(n39887), .Z(n39804) );
  XNOR U39507 ( .A(p_input[2048]), .B(p_input[768]), .Z(n39887) );
  XOR U39508 ( .A(n39875), .B(n39874), .Z(n39909) );
  XNOR U39509 ( .A(n39910), .B(n39881), .Z(n39874) );
  XNOR U39510 ( .A(n39870), .B(n39869), .Z(n39881) );
  XOR U39511 ( .A(n39911), .B(n39866), .Z(n39869) );
  XNOR U39512 ( .A(n29266), .B(p_input[778]), .Z(n39866) );
  XNOR U39513 ( .A(p_input[2059]), .B(p_input[779]), .Z(n39911) );
  XOR U39514 ( .A(p_input[2060]), .B(p_input[780]), .Z(n39870) );
  XNOR U39515 ( .A(n39880), .B(n39871), .Z(n39910) );
  XNOR U39516 ( .A(n29494), .B(p_input[769]), .Z(n39871) );
  XOR U39517 ( .A(n39912), .B(n39886), .Z(n39880) );
  XNOR U39518 ( .A(p_input[2063]), .B(p_input[783]), .Z(n39886) );
  XOR U39519 ( .A(n39877), .B(n39885), .Z(n39912) );
  XOR U39520 ( .A(n39913), .B(n39882), .Z(n39885) );
  XOR U39521 ( .A(p_input[2061]), .B(p_input[781]), .Z(n39882) );
  XNOR U39522 ( .A(p_input[2062]), .B(p_input[782]), .Z(n39913) );
  XNOR U39523 ( .A(n29036), .B(p_input[777]), .Z(n39877) );
  XNOR U39524 ( .A(n39893), .B(n39892), .Z(n39875) );
  XNOR U39525 ( .A(n39914), .B(n39898), .Z(n39892) );
  XOR U39526 ( .A(p_input[2056]), .B(p_input[776]), .Z(n39898) );
  XOR U39527 ( .A(n39889), .B(n39897), .Z(n39914) );
  XOR U39528 ( .A(n39915), .B(n39894), .Z(n39897) );
  XOR U39529 ( .A(p_input[2054]), .B(p_input[774]), .Z(n39894) );
  XNOR U39530 ( .A(p_input[2055]), .B(p_input[775]), .Z(n39915) );
  XNOR U39531 ( .A(n29039), .B(p_input[770]), .Z(n39889) );
  XNOR U39532 ( .A(n39903), .B(n39902), .Z(n39893) );
  XOR U39533 ( .A(n39916), .B(n39899), .Z(n39902) );
  XOR U39534 ( .A(p_input[2051]), .B(p_input[771]), .Z(n39899) );
  XNOR U39535 ( .A(p_input[2052]), .B(p_input[772]), .Z(n39916) );
  XOR U39536 ( .A(p_input[2053]), .B(p_input[773]), .Z(n39903) );
  XNOR U39537 ( .A(n39917), .B(n39918), .Z(n39801) );
  AND U39538 ( .A(n987), .B(n39919), .Z(n39918) );
  XNOR U39539 ( .A(n39920), .B(n39921), .Z(n987) );
  AND U39540 ( .A(n39922), .B(n39923), .Z(n39921) );
  XOR U39541 ( .A(n39815), .B(n39920), .Z(n39923) );
  XNOR U39542 ( .A(n39924), .B(n39920), .Z(n39922) );
  XOR U39543 ( .A(n39925), .B(n39926), .Z(n39920) );
  AND U39544 ( .A(n39927), .B(n39928), .Z(n39926) );
  XOR U39545 ( .A(n39830), .B(n39925), .Z(n39928) );
  XOR U39546 ( .A(n39925), .B(n39831), .Z(n39927) );
  XOR U39547 ( .A(n39929), .B(n39930), .Z(n39925) );
  AND U39548 ( .A(n39931), .B(n39932), .Z(n39930) );
  XOR U39549 ( .A(n39858), .B(n39929), .Z(n39932) );
  XOR U39550 ( .A(n39929), .B(n39859), .Z(n39931) );
  XOR U39551 ( .A(n39933), .B(n39934), .Z(n39929) );
  AND U39552 ( .A(n39935), .B(n39936), .Z(n39934) );
  XOR U39553 ( .A(n39933), .B(n39907), .Z(n39936) );
  XNOR U39554 ( .A(n39937), .B(n39938), .Z(n39761) );
  AND U39555 ( .A(n991), .B(n39939), .Z(n39938) );
  XNOR U39556 ( .A(n39940), .B(n39941), .Z(n991) );
  AND U39557 ( .A(n39942), .B(n39943), .Z(n39941) );
  XOR U39558 ( .A(n39940), .B(n39771), .Z(n39943) );
  XNOR U39559 ( .A(n39940), .B(n39731), .Z(n39942) );
  XOR U39560 ( .A(n39944), .B(n39945), .Z(n39940) );
  AND U39561 ( .A(n39946), .B(n39947), .Z(n39945) );
  XOR U39562 ( .A(n39944), .B(n39739), .Z(n39946) );
  XOR U39563 ( .A(n39948), .B(n39949), .Z(n39722) );
  AND U39564 ( .A(n995), .B(n39939), .Z(n39949) );
  XNOR U39565 ( .A(n39937), .B(n39948), .Z(n39939) );
  XNOR U39566 ( .A(n39950), .B(n39951), .Z(n995) );
  AND U39567 ( .A(n39952), .B(n39953), .Z(n39951) );
  XNOR U39568 ( .A(n39954), .B(n39950), .Z(n39953) );
  IV U39569 ( .A(n39771), .Z(n39954) );
  XOR U39570 ( .A(n39924), .B(n39955), .Z(n39771) );
  AND U39571 ( .A(n998), .B(n39956), .Z(n39955) );
  XOR U39572 ( .A(n39814), .B(n39811), .Z(n39956) );
  IV U39573 ( .A(n39924), .Z(n39814) );
  XNOR U39574 ( .A(n39731), .B(n39950), .Z(n39952) );
  XOR U39575 ( .A(n39957), .B(n39958), .Z(n39731) );
  AND U39576 ( .A(n1014), .B(n39959), .Z(n39958) );
  XOR U39577 ( .A(n39944), .B(n39960), .Z(n39950) );
  AND U39578 ( .A(n39961), .B(n39947), .Z(n39960) );
  XNOR U39579 ( .A(n39781), .B(n39944), .Z(n39947) );
  XOR U39580 ( .A(n39831), .B(n39962), .Z(n39781) );
  AND U39581 ( .A(n998), .B(n39963), .Z(n39962) );
  XOR U39582 ( .A(n39827), .B(n39831), .Z(n39963) );
  XNOR U39583 ( .A(n39964), .B(n39944), .Z(n39961) );
  IV U39584 ( .A(n39739), .Z(n39964) );
  XOR U39585 ( .A(n39965), .B(n39966), .Z(n39739) );
  AND U39586 ( .A(n1014), .B(n39967), .Z(n39966) );
  XOR U39587 ( .A(n39968), .B(n39969), .Z(n39944) );
  AND U39588 ( .A(n39970), .B(n39971), .Z(n39969) );
  XNOR U39589 ( .A(n39791), .B(n39968), .Z(n39971) );
  XOR U39590 ( .A(n39859), .B(n39972), .Z(n39791) );
  AND U39591 ( .A(n998), .B(n39973), .Z(n39972) );
  XOR U39592 ( .A(n39855), .B(n39859), .Z(n39973) );
  XOR U39593 ( .A(n39968), .B(n39748), .Z(n39970) );
  XOR U39594 ( .A(n39974), .B(n39975), .Z(n39748) );
  AND U39595 ( .A(n1014), .B(n39976), .Z(n39975) );
  XOR U39596 ( .A(n39977), .B(n39978), .Z(n39968) );
  AND U39597 ( .A(n39979), .B(n39980), .Z(n39978) );
  XNOR U39598 ( .A(n39977), .B(n39799), .Z(n39980) );
  XOR U39599 ( .A(n39908), .B(n39981), .Z(n39799) );
  AND U39600 ( .A(n998), .B(n39982), .Z(n39981) );
  XOR U39601 ( .A(n39904), .B(n39908), .Z(n39982) );
  XNOR U39602 ( .A(n39983), .B(n39977), .Z(n39979) );
  IV U39603 ( .A(n39758), .Z(n39983) );
  XOR U39604 ( .A(n39984), .B(n39985), .Z(n39758) );
  AND U39605 ( .A(n1014), .B(n39986), .Z(n39985) );
  AND U39606 ( .A(n39948), .B(n39937), .Z(n39977) );
  XNOR U39607 ( .A(n39987), .B(n39988), .Z(n39937) );
  AND U39608 ( .A(n998), .B(n39919), .Z(n39988) );
  XNOR U39609 ( .A(n39917), .B(n39987), .Z(n39919) );
  XNOR U39610 ( .A(n39989), .B(n39990), .Z(n998) );
  AND U39611 ( .A(n39991), .B(n39992), .Z(n39990) );
  XNOR U39612 ( .A(n39989), .B(n39811), .Z(n39992) );
  IV U39613 ( .A(n39815), .Z(n39811) );
  XOR U39614 ( .A(n39993), .B(n39994), .Z(n39815) );
  AND U39615 ( .A(n1002), .B(n39995), .Z(n39994) );
  XOR U39616 ( .A(n39996), .B(n39993), .Z(n39995) );
  XNOR U39617 ( .A(n39989), .B(n39924), .Z(n39991) );
  XOR U39618 ( .A(n39997), .B(n39998), .Z(n39924) );
  AND U39619 ( .A(n1010), .B(n39959), .Z(n39998) );
  XOR U39620 ( .A(n39957), .B(n39997), .Z(n39959) );
  XOR U39621 ( .A(n39999), .B(n40000), .Z(n39989) );
  AND U39622 ( .A(n40001), .B(n40002), .Z(n40000) );
  XNOR U39623 ( .A(n39999), .B(n39827), .Z(n40002) );
  IV U39624 ( .A(n39830), .Z(n39827) );
  XOR U39625 ( .A(n40003), .B(n40004), .Z(n39830) );
  AND U39626 ( .A(n1002), .B(n40005), .Z(n40004) );
  XOR U39627 ( .A(n40006), .B(n40003), .Z(n40005) );
  XOR U39628 ( .A(n39831), .B(n39999), .Z(n40001) );
  XOR U39629 ( .A(n40007), .B(n40008), .Z(n39831) );
  AND U39630 ( .A(n1010), .B(n39967), .Z(n40008) );
  XOR U39631 ( .A(n40007), .B(n39965), .Z(n39967) );
  XOR U39632 ( .A(n40009), .B(n40010), .Z(n39999) );
  AND U39633 ( .A(n40011), .B(n40012), .Z(n40010) );
  XNOR U39634 ( .A(n40009), .B(n39855), .Z(n40012) );
  IV U39635 ( .A(n39858), .Z(n39855) );
  XOR U39636 ( .A(n40013), .B(n40014), .Z(n39858) );
  AND U39637 ( .A(n1002), .B(n40015), .Z(n40014) );
  XNOR U39638 ( .A(n40016), .B(n40013), .Z(n40015) );
  XOR U39639 ( .A(n39859), .B(n40009), .Z(n40011) );
  XOR U39640 ( .A(n40017), .B(n40018), .Z(n39859) );
  AND U39641 ( .A(n1010), .B(n39976), .Z(n40018) );
  XOR U39642 ( .A(n40017), .B(n39974), .Z(n39976) );
  XOR U39643 ( .A(n39933), .B(n40019), .Z(n40009) );
  AND U39644 ( .A(n39935), .B(n40020), .Z(n40019) );
  XNOR U39645 ( .A(n39933), .B(n39904), .Z(n40020) );
  IV U39646 ( .A(n39907), .Z(n39904) );
  XOR U39647 ( .A(n40021), .B(n40022), .Z(n39907) );
  AND U39648 ( .A(n1002), .B(n40023), .Z(n40022) );
  XOR U39649 ( .A(n40024), .B(n40021), .Z(n40023) );
  XOR U39650 ( .A(n39908), .B(n39933), .Z(n39935) );
  XOR U39651 ( .A(n40025), .B(n40026), .Z(n39908) );
  AND U39652 ( .A(n1010), .B(n39986), .Z(n40026) );
  XOR U39653 ( .A(n40025), .B(n39984), .Z(n39986) );
  AND U39654 ( .A(n39987), .B(n39917), .Z(n39933) );
  XNOR U39655 ( .A(n40027), .B(n40028), .Z(n39917) );
  AND U39656 ( .A(n1002), .B(n40029), .Z(n40028) );
  XNOR U39657 ( .A(n40030), .B(n40027), .Z(n40029) );
  XNOR U39658 ( .A(n40031), .B(n40032), .Z(n1002) );
  AND U39659 ( .A(n40033), .B(n40034), .Z(n40032) );
  XOR U39660 ( .A(n39996), .B(n40031), .Z(n40034) );
  AND U39661 ( .A(n40035), .B(n40036), .Z(n39996) );
  XNOR U39662 ( .A(n39993), .B(n40031), .Z(n40033) );
  XNOR U39663 ( .A(n40037), .B(n40038), .Z(n39993) );
  AND U39664 ( .A(n1006), .B(n40039), .Z(n40038) );
  XNOR U39665 ( .A(n40040), .B(n40041), .Z(n40039) );
  XOR U39666 ( .A(n40042), .B(n40043), .Z(n40031) );
  AND U39667 ( .A(n40044), .B(n40045), .Z(n40043) );
  XNOR U39668 ( .A(n40042), .B(n40035), .Z(n40045) );
  IV U39669 ( .A(n40006), .Z(n40035) );
  XOR U39670 ( .A(n40046), .B(n40047), .Z(n40006) );
  XOR U39671 ( .A(n40048), .B(n40036), .Z(n40047) );
  AND U39672 ( .A(n40016), .B(n40049), .Z(n40036) );
  AND U39673 ( .A(n40050), .B(n40051), .Z(n40048) );
  XOR U39674 ( .A(n40052), .B(n40046), .Z(n40050) );
  XNOR U39675 ( .A(n40003), .B(n40042), .Z(n40044) );
  XNOR U39676 ( .A(n40053), .B(n40054), .Z(n40003) );
  AND U39677 ( .A(n1006), .B(n40055), .Z(n40054) );
  XNOR U39678 ( .A(n40056), .B(n40057), .Z(n40055) );
  XOR U39679 ( .A(n40058), .B(n40059), .Z(n40042) );
  AND U39680 ( .A(n40060), .B(n40061), .Z(n40059) );
  XNOR U39681 ( .A(n40058), .B(n40016), .Z(n40061) );
  XOR U39682 ( .A(n40062), .B(n40051), .Z(n40016) );
  XNOR U39683 ( .A(n40063), .B(n40046), .Z(n40051) );
  XOR U39684 ( .A(n40064), .B(n40065), .Z(n40046) );
  AND U39685 ( .A(n40066), .B(n40067), .Z(n40065) );
  XOR U39686 ( .A(n40068), .B(n40064), .Z(n40066) );
  XNOR U39687 ( .A(n40069), .B(n40070), .Z(n40063) );
  AND U39688 ( .A(n40071), .B(n40072), .Z(n40070) );
  XOR U39689 ( .A(n40069), .B(n40073), .Z(n40071) );
  XNOR U39690 ( .A(n40052), .B(n40049), .Z(n40062) );
  AND U39691 ( .A(n40074), .B(n40075), .Z(n40049) );
  XOR U39692 ( .A(n40076), .B(n40077), .Z(n40052) );
  AND U39693 ( .A(n40078), .B(n40079), .Z(n40077) );
  XOR U39694 ( .A(n40076), .B(n40080), .Z(n40078) );
  XNOR U39695 ( .A(n40013), .B(n40058), .Z(n40060) );
  XNOR U39696 ( .A(n40081), .B(n40082), .Z(n40013) );
  AND U39697 ( .A(n1006), .B(n40083), .Z(n40082) );
  XNOR U39698 ( .A(n40084), .B(n40085), .Z(n40083) );
  XOR U39699 ( .A(n40086), .B(n40087), .Z(n40058) );
  AND U39700 ( .A(n40088), .B(n40089), .Z(n40087) );
  XNOR U39701 ( .A(n40086), .B(n40074), .Z(n40089) );
  IV U39702 ( .A(n40024), .Z(n40074) );
  XNOR U39703 ( .A(n40090), .B(n40067), .Z(n40024) );
  XNOR U39704 ( .A(n40091), .B(n40073), .Z(n40067) );
  XOR U39705 ( .A(n40092), .B(n40093), .Z(n40073) );
  NOR U39706 ( .A(n40094), .B(n40095), .Z(n40093) );
  XNOR U39707 ( .A(n40092), .B(n40096), .Z(n40094) );
  XNOR U39708 ( .A(n40072), .B(n40064), .Z(n40091) );
  XOR U39709 ( .A(n40097), .B(n40098), .Z(n40064) );
  AND U39710 ( .A(n40099), .B(n40100), .Z(n40098) );
  XNOR U39711 ( .A(n40097), .B(n40101), .Z(n40099) );
  XNOR U39712 ( .A(n40102), .B(n40069), .Z(n40072) );
  XOR U39713 ( .A(n40103), .B(n40104), .Z(n40069) );
  AND U39714 ( .A(n40105), .B(n40106), .Z(n40104) );
  XOR U39715 ( .A(n40103), .B(n40107), .Z(n40105) );
  XNOR U39716 ( .A(n40108), .B(n40109), .Z(n40102) );
  NOR U39717 ( .A(n40110), .B(n40111), .Z(n40109) );
  XOR U39718 ( .A(n40108), .B(n40112), .Z(n40110) );
  XNOR U39719 ( .A(n40068), .B(n40075), .Z(n40090) );
  NOR U39720 ( .A(n40030), .B(n40113), .Z(n40075) );
  XOR U39721 ( .A(n40080), .B(n40079), .Z(n40068) );
  XNOR U39722 ( .A(n40114), .B(n40076), .Z(n40079) );
  XOR U39723 ( .A(n40115), .B(n40116), .Z(n40076) );
  AND U39724 ( .A(n40117), .B(n40118), .Z(n40116) );
  XOR U39725 ( .A(n40115), .B(n40119), .Z(n40117) );
  XNOR U39726 ( .A(n40120), .B(n40121), .Z(n40114) );
  NOR U39727 ( .A(n40122), .B(n40123), .Z(n40121) );
  XNOR U39728 ( .A(n40120), .B(n40124), .Z(n40122) );
  XOR U39729 ( .A(n40125), .B(n40126), .Z(n40080) );
  NOR U39730 ( .A(n40127), .B(n40128), .Z(n40126) );
  XNOR U39731 ( .A(n40125), .B(n40129), .Z(n40127) );
  XNOR U39732 ( .A(n40021), .B(n40086), .Z(n40088) );
  XNOR U39733 ( .A(n40130), .B(n40131), .Z(n40021) );
  AND U39734 ( .A(n1006), .B(n40132), .Z(n40131) );
  XNOR U39735 ( .A(n40133), .B(n40134), .Z(n40132) );
  AND U39736 ( .A(n40027), .B(n40030), .Z(n40086) );
  XOR U39737 ( .A(n40135), .B(n40113), .Z(n40030) );
  XNOR U39738 ( .A(p_input[2048]), .B(p_input[784]), .Z(n40113) );
  XOR U39739 ( .A(n40101), .B(n40100), .Z(n40135) );
  XNOR U39740 ( .A(n40136), .B(n40107), .Z(n40100) );
  XNOR U39741 ( .A(n40096), .B(n40095), .Z(n40107) );
  XOR U39742 ( .A(n40137), .B(n40092), .Z(n40095) );
  XNOR U39743 ( .A(n29266), .B(p_input[794]), .Z(n40092) );
  XNOR U39744 ( .A(p_input[2059]), .B(p_input[795]), .Z(n40137) );
  XOR U39745 ( .A(p_input[2060]), .B(p_input[796]), .Z(n40096) );
  XNOR U39746 ( .A(n40106), .B(n40097), .Z(n40136) );
  XNOR U39747 ( .A(n29494), .B(p_input[785]), .Z(n40097) );
  XOR U39748 ( .A(n40138), .B(n40112), .Z(n40106) );
  XNOR U39749 ( .A(p_input[2063]), .B(p_input[799]), .Z(n40112) );
  XOR U39750 ( .A(n40103), .B(n40111), .Z(n40138) );
  XOR U39751 ( .A(n40139), .B(n40108), .Z(n40111) );
  XOR U39752 ( .A(p_input[2061]), .B(p_input[797]), .Z(n40108) );
  XNOR U39753 ( .A(p_input[2062]), .B(p_input[798]), .Z(n40139) );
  XNOR U39754 ( .A(n29036), .B(p_input[793]), .Z(n40103) );
  XNOR U39755 ( .A(n40119), .B(n40118), .Z(n40101) );
  XNOR U39756 ( .A(n40140), .B(n40124), .Z(n40118) );
  XOR U39757 ( .A(p_input[2056]), .B(p_input[792]), .Z(n40124) );
  XOR U39758 ( .A(n40115), .B(n40123), .Z(n40140) );
  XOR U39759 ( .A(n40141), .B(n40120), .Z(n40123) );
  XOR U39760 ( .A(p_input[2054]), .B(p_input[790]), .Z(n40120) );
  XNOR U39761 ( .A(p_input[2055]), .B(p_input[791]), .Z(n40141) );
  XNOR U39762 ( .A(n29039), .B(p_input[786]), .Z(n40115) );
  XNOR U39763 ( .A(n40129), .B(n40128), .Z(n40119) );
  XOR U39764 ( .A(n40142), .B(n40125), .Z(n40128) );
  XOR U39765 ( .A(p_input[2051]), .B(p_input[787]), .Z(n40125) );
  XNOR U39766 ( .A(p_input[2052]), .B(p_input[788]), .Z(n40142) );
  XOR U39767 ( .A(p_input[2053]), .B(p_input[789]), .Z(n40129) );
  XNOR U39768 ( .A(n40143), .B(n40144), .Z(n40027) );
  AND U39769 ( .A(n1006), .B(n40145), .Z(n40144) );
  XNOR U39770 ( .A(n40146), .B(n40147), .Z(n1006) );
  AND U39771 ( .A(n40148), .B(n40149), .Z(n40147) );
  XOR U39772 ( .A(n40041), .B(n40146), .Z(n40149) );
  XNOR U39773 ( .A(n40150), .B(n40146), .Z(n40148) );
  XOR U39774 ( .A(n40151), .B(n40152), .Z(n40146) );
  AND U39775 ( .A(n40153), .B(n40154), .Z(n40152) );
  XOR U39776 ( .A(n40056), .B(n40151), .Z(n40154) );
  XOR U39777 ( .A(n40151), .B(n40057), .Z(n40153) );
  XOR U39778 ( .A(n40155), .B(n40156), .Z(n40151) );
  AND U39779 ( .A(n40157), .B(n40158), .Z(n40156) );
  XOR U39780 ( .A(n40084), .B(n40155), .Z(n40158) );
  XOR U39781 ( .A(n40155), .B(n40085), .Z(n40157) );
  XOR U39782 ( .A(n40159), .B(n40160), .Z(n40155) );
  AND U39783 ( .A(n40161), .B(n40162), .Z(n40160) );
  XOR U39784 ( .A(n40159), .B(n40133), .Z(n40162) );
  XNOR U39785 ( .A(n40163), .B(n40164), .Z(n39987) );
  AND U39786 ( .A(n1010), .B(n40165), .Z(n40164) );
  XNOR U39787 ( .A(n40166), .B(n40167), .Z(n1010) );
  AND U39788 ( .A(n40168), .B(n40169), .Z(n40167) );
  XOR U39789 ( .A(n40166), .B(n39997), .Z(n40169) );
  XNOR U39790 ( .A(n40166), .B(n39957), .Z(n40168) );
  XOR U39791 ( .A(n40170), .B(n40171), .Z(n40166) );
  AND U39792 ( .A(n40172), .B(n40173), .Z(n40171) );
  XOR U39793 ( .A(n40170), .B(n39965), .Z(n40172) );
  XOR U39794 ( .A(n40174), .B(n40175), .Z(n39948) );
  AND U39795 ( .A(n1014), .B(n40165), .Z(n40175) );
  XNOR U39796 ( .A(n40163), .B(n40174), .Z(n40165) );
  XNOR U39797 ( .A(n40176), .B(n40177), .Z(n1014) );
  AND U39798 ( .A(n40178), .B(n40179), .Z(n40177) );
  XNOR U39799 ( .A(n40180), .B(n40176), .Z(n40179) );
  IV U39800 ( .A(n39997), .Z(n40180) );
  XOR U39801 ( .A(n40150), .B(n40181), .Z(n39997) );
  AND U39802 ( .A(n1017), .B(n40182), .Z(n40181) );
  XOR U39803 ( .A(n40040), .B(n40037), .Z(n40182) );
  IV U39804 ( .A(n40150), .Z(n40040) );
  XNOR U39805 ( .A(n39957), .B(n40176), .Z(n40178) );
  XOR U39806 ( .A(n40183), .B(n40184), .Z(n39957) );
  AND U39807 ( .A(n1033), .B(n40185), .Z(n40184) );
  XOR U39808 ( .A(n40170), .B(n40186), .Z(n40176) );
  AND U39809 ( .A(n40187), .B(n40173), .Z(n40186) );
  XNOR U39810 ( .A(n40007), .B(n40170), .Z(n40173) );
  XOR U39811 ( .A(n40057), .B(n40188), .Z(n40007) );
  AND U39812 ( .A(n1017), .B(n40189), .Z(n40188) );
  XOR U39813 ( .A(n40053), .B(n40057), .Z(n40189) );
  XNOR U39814 ( .A(n40190), .B(n40170), .Z(n40187) );
  IV U39815 ( .A(n39965), .Z(n40190) );
  XOR U39816 ( .A(n40191), .B(n40192), .Z(n39965) );
  AND U39817 ( .A(n1033), .B(n40193), .Z(n40192) );
  XOR U39818 ( .A(n40194), .B(n40195), .Z(n40170) );
  AND U39819 ( .A(n40196), .B(n40197), .Z(n40195) );
  XNOR U39820 ( .A(n40017), .B(n40194), .Z(n40197) );
  XOR U39821 ( .A(n40085), .B(n40198), .Z(n40017) );
  AND U39822 ( .A(n1017), .B(n40199), .Z(n40198) );
  XOR U39823 ( .A(n40081), .B(n40085), .Z(n40199) );
  XOR U39824 ( .A(n40194), .B(n39974), .Z(n40196) );
  XOR U39825 ( .A(n40200), .B(n40201), .Z(n39974) );
  AND U39826 ( .A(n1033), .B(n40202), .Z(n40201) );
  XOR U39827 ( .A(n40203), .B(n40204), .Z(n40194) );
  AND U39828 ( .A(n40205), .B(n40206), .Z(n40204) );
  XNOR U39829 ( .A(n40203), .B(n40025), .Z(n40206) );
  XOR U39830 ( .A(n40134), .B(n40207), .Z(n40025) );
  AND U39831 ( .A(n1017), .B(n40208), .Z(n40207) );
  XOR U39832 ( .A(n40130), .B(n40134), .Z(n40208) );
  XNOR U39833 ( .A(n40209), .B(n40203), .Z(n40205) );
  IV U39834 ( .A(n39984), .Z(n40209) );
  XOR U39835 ( .A(n40210), .B(n40211), .Z(n39984) );
  AND U39836 ( .A(n1033), .B(n40212), .Z(n40211) );
  AND U39837 ( .A(n40174), .B(n40163), .Z(n40203) );
  XNOR U39838 ( .A(n40213), .B(n40214), .Z(n40163) );
  AND U39839 ( .A(n1017), .B(n40145), .Z(n40214) );
  XNOR U39840 ( .A(n40143), .B(n40213), .Z(n40145) );
  XNOR U39841 ( .A(n40215), .B(n40216), .Z(n1017) );
  AND U39842 ( .A(n40217), .B(n40218), .Z(n40216) );
  XNOR U39843 ( .A(n40215), .B(n40037), .Z(n40218) );
  IV U39844 ( .A(n40041), .Z(n40037) );
  XOR U39845 ( .A(n40219), .B(n40220), .Z(n40041) );
  AND U39846 ( .A(n1021), .B(n40221), .Z(n40220) );
  XOR U39847 ( .A(n40222), .B(n40219), .Z(n40221) );
  XNOR U39848 ( .A(n40215), .B(n40150), .Z(n40217) );
  XOR U39849 ( .A(n40223), .B(n40224), .Z(n40150) );
  AND U39850 ( .A(n1029), .B(n40185), .Z(n40224) );
  XOR U39851 ( .A(n40183), .B(n40223), .Z(n40185) );
  XOR U39852 ( .A(n40225), .B(n40226), .Z(n40215) );
  AND U39853 ( .A(n40227), .B(n40228), .Z(n40226) );
  XNOR U39854 ( .A(n40225), .B(n40053), .Z(n40228) );
  IV U39855 ( .A(n40056), .Z(n40053) );
  XOR U39856 ( .A(n40229), .B(n40230), .Z(n40056) );
  AND U39857 ( .A(n1021), .B(n40231), .Z(n40230) );
  XOR U39858 ( .A(n40232), .B(n40229), .Z(n40231) );
  XOR U39859 ( .A(n40057), .B(n40225), .Z(n40227) );
  XOR U39860 ( .A(n40233), .B(n40234), .Z(n40057) );
  AND U39861 ( .A(n1029), .B(n40193), .Z(n40234) );
  XOR U39862 ( .A(n40233), .B(n40191), .Z(n40193) );
  XOR U39863 ( .A(n40235), .B(n40236), .Z(n40225) );
  AND U39864 ( .A(n40237), .B(n40238), .Z(n40236) );
  XNOR U39865 ( .A(n40235), .B(n40081), .Z(n40238) );
  IV U39866 ( .A(n40084), .Z(n40081) );
  XOR U39867 ( .A(n40239), .B(n40240), .Z(n40084) );
  AND U39868 ( .A(n1021), .B(n40241), .Z(n40240) );
  XNOR U39869 ( .A(n40242), .B(n40239), .Z(n40241) );
  XOR U39870 ( .A(n40085), .B(n40235), .Z(n40237) );
  XOR U39871 ( .A(n40243), .B(n40244), .Z(n40085) );
  AND U39872 ( .A(n1029), .B(n40202), .Z(n40244) );
  XOR U39873 ( .A(n40243), .B(n40200), .Z(n40202) );
  XOR U39874 ( .A(n40159), .B(n40245), .Z(n40235) );
  AND U39875 ( .A(n40161), .B(n40246), .Z(n40245) );
  XNOR U39876 ( .A(n40159), .B(n40130), .Z(n40246) );
  IV U39877 ( .A(n40133), .Z(n40130) );
  XOR U39878 ( .A(n40247), .B(n40248), .Z(n40133) );
  AND U39879 ( .A(n1021), .B(n40249), .Z(n40248) );
  XOR U39880 ( .A(n40250), .B(n40247), .Z(n40249) );
  XOR U39881 ( .A(n40134), .B(n40159), .Z(n40161) );
  XOR U39882 ( .A(n40251), .B(n40252), .Z(n40134) );
  AND U39883 ( .A(n1029), .B(n40212), .Z(n40252) );
  XOR U39884 ( .A(n40251), .B(n40210), .Z(n40212) );
  AND U39885 ( .A(n40213), .B(n40143), .Z(n40159) );
  XNOR U39886 ( .A(n40253), .B(n40254), .Z(n40143) );
  AND U39887 ( .A(n1021), .B(n40255), .Z(n40254) );
  XNOR U39888 ( .A(n40256), .B(n40253), .Z(n40255) );
  XNOR U39889 ( .A(n40257), .B(n40258), .Z(n1021) );
  AND U39890 ( .A(n40259), .B(n40260), .Z(n40258) );
  XOR U39891 ( .A(n40222), .B(n40257), .Z(n40260) );
  AND U39892 ( .A(n40261), .B(n40262), .Z(n40222) );
  XNOR U39893 ( .A(n40219), .B(n40257), .Z(n40259) );
  XNOR U39894 ( .A(n40263), .B(n40264), .Z(n40219) );
  AND U39895 ( .A(n1025), .B(n40265), .Z(n40264) );
  XNOR U39896 ( .A(n40266), .B(n40267), .Z(n40265) );
  XOR U39897 ( .A(n40268), .B(n40269), .Z(n40257) );
  AND U39898 ( .A(n40270), .B(n40271), .Z(n40269) );
  XNOR U39899 ( .A(n40268), .B(n40261), .Z(n40271) );
  IV U39900 ( .A(n40232), .Z(n40261) );
  XOR U39901 ( .A(n40272), .B(n40273), .Z(n40232) );
  XOR U39902 ( .A(n40274), .B(n40262), .Z(n40273) );
  AND U39903 ( .A(n40242), .B(n40275), .Z(n40262) );
  AND U39904 ( .A(n40276), .B(n40277), .Z(n40274) );
  XOR U39905 ( .A(n40278), .B(n40272), .Z(n40276) );
  XNOR U39906 ( .A(n40229), .B(n40268), .Z(n40270) );
  XNOR U39907 ( .A(n40279), .B(n40280), .Z(n40229) );
  AND U39908 ( .A(n1025), .B(n40281), .Z(n40280) );
  XNOR U39909 ( .A(n40282), .B(n40283), .Z(n40281) );
  XOR U39910 ( .A(n40284), .B(n40285), .Z(n40268) );
  AND U39911 ( .A(n40286), .B(n40287), .Z(n40285) );
  XNOR U39912 ( .A(n40284), .B(n40242), .Z(n40287) );
  XOR U39913 ( .A(n40288), .B(n40277), .Z(n40242) );
  XNOR U39914 ( .A(n40289), .B(n40272), .Z(n40277) );
  XOR U39915 ( .A(n40290), .B(n40291), .Z(n40272) );
  AND U39916 ( .A(n40292), .B(n40293), .Z(n40291) );
  XOR U39917 ( .A(n40294), .B(n40290), .Z(n40292) );
  XNOR U39918 ( .A(n40295), .B(n40296), .Z(n40289) );
  AND U39919 ( .A(n40297), .B(n40298), .Z(n40296) );
  XOR U39920 ( .A(n40295), .B(n40299), .Z(n40297) );
  XNOR U39921 ( .A(n40278), .B(n40275), .Z(n40288) );
  AND U39922 ( .A(n40300), .B(n40301), .Z(n40275) );
  XOR U39923 ( .A(n40302), .B(n40303), .Z(n40278) );
  AND U39924 ( .A(n40304), .B(n40305), .Z(n40303) );
  XOR U39925 ( .A(n40302), .B(n40306), .Z(n40304) );
  XNOR U39926 ( .A(n40239), .B(n40284), .Z(n40286) );
  XNOR U39927 ( .A(n40307), .B(n40308), .Z(n40239) );
  AND U39928 ( .A(n1025), .B(n40309), .Z(n40308) );
  XNOR U39929 ( .A(n40310), .B(n40311), .Z(n40309) );
  XOR U39930 ( .A(n40312), .B(n40313), .Z(n40284) );
  AND U39931 ( .A(n40314), .B(n40315), .Z(n40313) );
  XNOR U39932 ( .A(n40312), .B(n40300), .Z(n40315) );
  IV U39933 ( .A(n40250), .Z(n40300) );
  XNOR U39934 ( .A(n40316), .B(n40293), .Z(n40250) );
  XNOR U39935 ( .A(n40317), .B(n40299), .Z(n40293) );
  XOR U39936 ( .A(n40318), .B(n40319), .Z(n40299) );
  NOR U39937 ( .A(n40320), .B(n40321), .Z(n40319) );
  XNOR U39938 ( .A(n40318), .B(n40322), .Z(n40320) );
  XNOR U39939 ( .A(n40298), .B(n40290), .Z(n40317) );
  XOR U39940 ( .A(n40323), .B(n40324), .Z(n40290) );
  AND U39941 ( .A(n40325), .B(n40326), .Z(n40324) );
  XNOR U39942 ( .A(n40323), .B(n40327), .Z(n40325) );
  XNOR U39943 ( .A(n40328), .B(n40295), .Z(n40298) );
  XOR U39944 ( .A(n40329), .B(n40330), .Z(n40295) );
  AND U39945 ( .A(n40331), .B(n40332), .Z(n40330) );
  XOR U39946 ( .A(n40329), .B(n40333), .Z(n40331) );
  XNOR U39947 ( .A(n40334), .B(n40335), .Z(n40328) );
  NOR U39948 ( .A(n40336), .B(n40337), .Z(n40335) );
  XOR U39949 ( .A(n40334), .B(n40338), .Z(n40336) );
  XNOR U39950 ( .A(n40294), .B(n40301), .Z(n40316) );
  NOR U39951 ( .A(n40256), .B(n40339), .Z(n40301) );
  XOR U39952 ( .A(n40306), .B(n40305), .Z(n40294) );
  XNOR U39953 ( .A(n40340), .B(n40302), .Z(n40305) );
  XOR U39954 ( .A(n40341), .B(n40342), .Z(n40302) );
  AND U39955 ( .A(n40343), .B(n40344), .Z(n40342) );
  XOR U39956 ( .A(n40341), .B(n40345), .Z(n40343) );
  XNOR U39957 ( .A(n40346), .B(n40347), .Z(n40340) );
  NOR U39958 ( .A(n40348), .B(n40349), .Z(n40347) );
  XNOR U39959 ( .A(n40346), .B(n40350), .Z(n40348) );
  XOR U39960 ( .A(n40351), .B(n40352), .Z(n40306) );
  NOR U39961 ( .A(n40353), .B(n40354), .Z(n40352) );
  XNOR U39962 ( .A(n40351), .B(n40355), .Z(n40353) );
  XNOR U39963 ( .A(n40247), .B(n40312), .Z(n40314) );
  XNOR U39964 ( .A(n40356), .B(n40357), .Z(n40247) );
  AND U39965 ( .A(n1025), .B(n40358), .Z(n40357) );
  XNOR U39966 ( .A(n40359), .B(n40360), .Z(n40358) );
  AND U39967 ( .A(n40253), .B(n40256), .Z(n40312) );
  XOR U39968 ( .A(n40361), .B(n40339), .Z(n40256) );
  XNOR U39969 ( .A(p_input[2048]), .B(p_input[800]), .Z(n40339) );
  XOR U39970 ( .A(n40327), .B(n40326), .Z(n40361) );
  XNOR U39971 ( .A(n40362), .B(n40333), .Z(n40326) );
  XNOR U39972 ( .A(n40322), .B(n40321), .Z(n40333) );
  XOR U39973 ( .A(n40363), .B(n40318), .Z(n40321) );
  XNOR U39974 ( .A(n29266), .B(p_input[810]), .Z(n40318) );
  XNOR U39975 ( .A(p_input[2059]), .B(p_input[811]), .Z(n40363) );
  XOR U39976 ( .A(p_input[2060]), .B(p_input[812]), .Z(n40322) );
  XNOR U39977 ( .A(n40332), .B(n40323), .Z(n40362) );
  XNOR U39978 ( .A(n29494), .B(p_input[801]), .Z(n40323) );
  XOR U39979 ( .A(n40364), .B(n40338), .Z(n40332) );
  XNOR U39980 ( .A(p_input[2063]), .B(p_input[815]), .Z(n40338) );
  XOR U39981 ( .A(n40329), .B(n40337), .Z(n40364) );
  XOR U39982 ( .A(n40365), .B(n40334), .Z(n40337) );
  XOR U39983 ( .A(p_input[2061]), .B(p_input[813]), .Z(n40334) );
  XNOR U39984 ( .A(p_input[2062]), .B(p_input[814]), .Z(n40365) );
  XNOR U39985 ( .A(n29036), .B(p_input[809]), .Z(n40329) );
  XNOR U39986 ( .A(n40345), .B(n40344), .Z(n40327) );
  XNOR U39987 ( .A(n40366), .B(n40350), .Z(n40344) );
  XOR U39988 ( .A(p_input[2056]), .B(p_input[808]), .Z(n40350) );
  XOR U39989 ( .A(n40341), .B(n40349), .Z(n40366) );
  XOR U39990 ( .A(n40367), .B(n40346), .Z(n40349) );
  XOR U39991 ( .A(p_input[2054]), .B(p_input[806]), .Z(n40346) );
  XNOR U39992 ( .A(p_input[2055]), .B(p_input[807]), .Z(n40367) );
  XNOR U39993 ( .A(n29039), .B(p_input[802]), .Z(n40341) );
  XNOR U39994 ( .A(n40355), .B(n40354), .Z(n40345) );
  XOR U39995 ( .A(n40368), .B(n40351), .Z(n40354) );
  XOR U39996 ( .A(p_input[2051]), .B(p_input[803]), .Z(n40351) );
  XNOR U39997 ( .A(p_input[2052]), .B(p_input[804]), .Z(n40368) );
  XOR U39998 ( .A(p_input[2053]), .B(p_input[805]), .Z(n40355) );
  XNOR U39999 ( .A(n40369), .B(n40370), .Z(n40253) );
  AND U40000 ( .A(n1025), .B(n40371), .Z(n40370) );
  XNOR U40001 ( .A(n40372), .B(n40373), .Z(n1025) );
  AND U40002 ( .A(n40374), .B(n40375), .Z(n40373) );
  XOR U40003 ( .A(n40267), .B(n40372), .Z(n40375) );
  XNOR U40004 ( .A(n40376), .B(n40372), .Z(n40374) );
  XOR U40005 ( .A(n40377), .B(n40378), .Z(n40372) );
  AND U40006 ( .A(n40379), .B(n40380), .Z(n40378) );
  XOR U40007 ( .A(n40282), .B(n40377), .Z(n40380) );
  XOR U40008 ( .A(n40377), .B(n40283), .Z(n40379) );
  XOR U40009 ( .A(n40381), .B(n40382), .Z(n40377) );
  AND U40010 ( .A(n40383), .B(n40384), .Z(n40382) );
  XOR U40011 ( .A(n40310), .B(n40381), .Z(n40384) );
  XOR U40012 ( .A(n40381), .B(n40311), .Z(n40383) );
  XOR U40013 ( .A(n40385), .B(n40386), .Z(n40381) );
  AND U40014 ( .A(n40387), .B(n40388), .Z(n40386) );
  XOR U40015 ( .A(n40385), .B(n40359), .Z(n40388) );
  XNOR U40016 ( .A(n40389), .B(n40390), .Z(n40213) );
  AND U40017 ( .A(n1029), .B(n40391), .Z(n40390) );
  XNOR U40018 ( .A(n40392), .B(n40393), .Z(n1029) );
  AND U40019 ( .A(n40394), .B(n40395), .Z(n40393) );
  XOR U40020 ( .A(n40392), .B(n40223), .Z(n40395) );
  XNOR U40021 ( .A(n40392), .B(n40183), .Z(n40394) );
  XOR U40022 ( .A(n40396), .B(n40397), .Z(n40392) );
  AND U40023 ( .A(n40398), .B(n40399), .Z(n40397) );
  XOR U40024 ( .A(n40396), .B(n40191), .Z(n40398) );
  XOR U40025 ( .A(n40400), .B(n40401), .Z(n40174) );
  AND U40026 ( .A(n1033), .B(n40391), .Z(n40401) );
  XNOR U40027 ( .A(n40389), .B(n40400), .Z(n40391) );
  XNOR U40028 ( .A(n40402), .B(n40403), .Z(n1033) );
  AND U40029 ( .A(n40404), .B(n40405), .Z(n40403) );
  XNOR U40030 ( .A(n40406), .B(n40402), .Z(n40405) );
  IV U40031 ( .A(n40223), .Z(n40406) );
  XOR U40032 ( .A(n40376), .B(n40407), .Z(n40223) );
  AND U40033 ( .A(n1036), .B(n40408), .Z(n40407) );
  XOR U40034 ( .A(n40266), .B(n40263), .Z(n40408) );
  IV U40035 ( .A(n40376), .Z(n40266) );
  XNOR U40036 ( .A(n40183), .B(n40402), .Z(n40404) );
  XOR U40037 ( .A(n40409), .B(n40410), .Z(n40183) );
  AND U40038 ( .A(n1052), .B(n40411), .Z(n40410) );
  XOR U40039 ( .A(n40396), .B(n40412), .Z(n40402) );
  AND U40040 ( .A(n40413), .B(n40399), .Z(n40412) );
  XNOR U40041 ( .A(n40233), .B(n40396), .Z(n40399) );
  XOR U40042 ( .A(n40283), .B(n40414), .Z(n40233) );
  AND U40043 ( .A(n1036), .B(n40415), .Z(n40414) );
  XOR U40044 ( .A(n40279), .B(n40283), .Z(n40415) );
  XNOR U40045 ( .A(n40416), .B(n40396), .Z(n40413) );
  IV U40046 ( .A(n40191), .Z(n40416) );
  XOR U40047 ( .A(n40417), .B(n40418), .Z(n40191) );
  AND U40048 ( .A(n1052), .B(n40419), .Z(n40418) );
  XOR U40049 ( .A(n40420), .B(n40421), .Z(n40396) );
  AND U40050 ( .A(n40422), .B(n40423), .Z(n40421) );
  XNOR U40051 ( .A(n40243), .B(n40420), .Z(n40423) );
  XOR U40052 ( .A(n40311), .B(n40424), .Z(n40243) );
  AND U40053 ( .A(n1036), .B(n40425), .Z(n40424) );
  XOR U40054 ( .A(n40307), .B(n40311), .Z(n40425) );
  XOR U40055 ( .A(n40420), .B(n40200), .Z(n40422) );
  XOR U40056 ( .A(n40426), .B(n40427), .Z(n40200) );
  AND U40057 ( .A(n1052), .B(n40428), .Z(n40427) );
  XOR U40058 ( .A(n40429), .B(n40430), .Z(n40420) );
  AND U40059 ( .A(n40431), .B(n40432), .Z(n40430) );
  XNOR U40060 ( .A(n40429), .B(n40251), .Z(n40432) );
  XOR U40061 ( .A(n40360), .B(n40433), .Z(n40251) );
  AND U40062 ( .A(n1036), .B(n40434), .Z(n40433) );
  XOR U40063 ( .A(n40356), .B(n40360), .Z(n40434) );
  XNOR U40064 ( .A(n40435), .B(n40429), .Z(n40431) );
  IV U40065 ( .A(n40210), .Z(n40435) );
  XOR U40066 ( .A(n40436), .B(n40437), .Z(n40210) );
  AND U40067 ( .A(n1052), .B(n40438), .Z(n40437) );
  AND U40068 ( .A(n40400), .B(n40389), .Z(n40429) );
  XNOR U40069 ( .A(n40439), .B(n40440), .Z(n40389) );
  AND U40070 ( .A(n1036), .B(n40371), .Z(n40440) );
  XNOR U40071 ( .A(n40369), .B(n40439), .Z(n40371) );
  XNOR U40072 ( .A(n40441), .B(n40442), .Z(n1036) );
  AND U40073 ( .A(n40443), .B(n40444), .Z(n40442) );
  XNOR U40074 ( .A(n40441), .B(n40263), .Z(n40444) );
  IV U40075 ( .A(n40267), .Z(n40263) );
  XOR U40076 ( .A(n40445), .B(n40446), .Z(n40267) );
  AND U40077 ( .A(n1040), .B(n40447), .Z(n40446) );
  XOR U40078 ( .A(n40448), .B(n40445), .Z(n40447) );
  XNOR U40079 ( .A(n40441), .B(n40376), .Z(n40443) );
  XOR U40080 ( .A(n40449), .B(n40450), .Z(n40376) );
  AND U40081 ( .A(n1048), .B(n40411), .Z(n40450) );
  XOR U40082 ( .A(n40409), .B(n40449), .Z(n40411) );
  XOR U40083 ( .A(n40451), .B(n40452), .Z(n40441) );
  AND U40084 ( .A(n40453), .B(n40454), .Z(n40452) );
  XNOR U40085 ( .A(n40451), .B(n40279), .Z(n40454) );
  IV U40086 ( .A(n40282), .Z(n40279) );
  XOR U40087 ( .A(n40455), .B(n40456), .Z(n40282) );
  AND U40088 ( .A(n1040), .B(n40457), .Z(n40456) );
  XOR U40089 ( .A(n40458), .B(n40455), .Z(n40457) );
  XOR U40090 ( .A(n40283), .B(n40451), .Z(n40453) );
  XOR U40091 ( .A(n40459), .B(n40460), .Z(n40283) );
  AND U40092 ( .A(n1048), .B(n40419), .Z(n40460) );
  XOR U40093 ( .A(n40459), .B(n40417), .Z(n40419) );
  XOR U40094 ( .A(n40461), .B(n40462), .Z(n40451) );
  AND U40095 ( .A(n40463), .B(n40464), .Z(n40462) );
  XNOR U40096 ( .A(n40461), .B(n40307), .Z(n40464) );
  IV U40097 ( .A(n40310), .Z(n40307) );
  XOR U40098 ( .A(n40465), .B(n40466), .Z(n40310) );
  AND U40099 ( .A(n1040), .B(n40467), .Z(n40466) );
  XNOR U40100 ( .A(n40468), .B(n40465), .Z(n40467) );
  XOR U40101 ( .A(n40311), .B(n40461), .Z(n40463) );
  XOR U40102 ( .A(n40469), .B(n40470), .Z(n40311) );
  AND U40103 ( .A(n1048), .B(n40428), .Z(n40470) );
  XOR U40104 ( .A(n40469), .B(n40426), .Z(n40428) );
  XOR U40105 ( .A(n40385), .B(n40471), .Z(n40461) );
  AND U40106 ( .A(n40387), .B(n40472), .Z(n40471) );
  XNOR U40107 ( .A(n40385), .B(n40356), .Z(n40472) );
  IV U40108 ( .A(n40359), .Z(n40356) );
  XOR U40109 ( .A(n40473), .B(n40474), .Z(n40359) );
  AND U40110 ( .A(n1040), .B(n40475), .Z(n40474) );
  XOR U40111 ( .A(n40476), .B(n40473), .Z(n40475) );
  XOR U40112 ( .A(n40360), .B(n40385), .Z(n40387) );
  XOR U40113 ( .A(n40477), .B(n40478), .Z(n40360) );
  AND U40114 ( .A(n1048), .B(n40438), .Z(n40478) );
  XOR U40115 ( .A(n40477), .B(n40436), .Z(n40438) );
  AND U40116 ( .A(n40439), .B(n40369), .Z(n40385) );
  XNOR U40117 ( .A(n40479), .B(n40480), .Z(n40369) );
  AND U40118 ( .A(n1040), .B(n40481), .Z(n40480) );
  XNOR U40119 ( .A(n40482), .B(n40479), .Z(n40481) );
  XNOR U40120 ( .A(n40483), .B(n40484), .Z(n1040) );
  AND U40121 ( .A(n40485), .B(n40486), .Z(n40484) );
  XOR U40122 ( .A(n40448), .B(n40483), .Z(n40486) );
  AND U40123 ( .A(n40487), .B(n40488), .Z(n40448) );
  XNOR U40124 ( .A(n40445), .B(n40483), .Z(n40485) );
  XNOR U40125 ( .A(n40489), .B(n40490), .Z(n40445) );
  AND U40126 ( .A(n1044), .B(n40491), .Z(n40490) );
  XNOR U40127 ( .A(n40492), .B(n40493), .Z(n40491) );
  XOR U40128 ( .A(n40494), .B(n40495), .Z(n40483) );
  AND U40129 ( .A(n40496), .B(n40497), .Z(n40495) );
  XNOR U40130 ( .A(n40494), .B(n40487), .Z(n40497) );
  IV U40131 ( .A(n40458), .Z(n40487) );
  XOR U40132 ( .A(n40498), .B(n40499), .Z(n40458) );
  XOR U40133 ( .A(n40500), .B(n40488), .Z(n40499) );
  AND U40134 ( .A(n40468), .B(n40501), .Z(n40488) );
  AND U40135 ( .A(n40502), .B(n40503), .Z(n40500) );
  XOR U40136 ( .A(n40504), .B(n40498), .Z(n40502) );
  XNOR U40137 ( .A(n40455), .B(n40494), .Z(n40496) );
  XNOR U40138 ( .A(n40505), .B(n40506), .Z(n40455) );
  AND U40139 ( .A(n1044), .B(n40507), .Z(n40506) );
  XNOR U40140 ( .A(n40508), .B(n40509), .Z(n40507) );
  XOR U40141 ( .A(n40510), .B(n40511), .Z(n40494) );
  AND U40142 ( .A(n40512), .B(n40513), .Z(n40511) );
  XNOR U40143 ( .A(n40510), .B(n40468), .Z(n40513) );
  XOR U40144 ( .A(n40514), .B(n40503), .Z(n40468) );
  XNOR U40145 ( .A(n40515), .B(n40498), .Z(n40503) );
  XOR U40146 ( .A(n40516), .B(n40517), .Z(n40498) );
  AND U40147 ( .A(n40518), .B(n40519), .Z(n40517) );
  XOR U40148 ( .A(n40520), .B(n40516), .Z(n40518) );
  XNOR U40149 ( .A(n40521), .B(n40522), .Z(n40515) );
  AND U40150 ( .A(n40523), .B(n40524), .Z(n40522) );
  XOR U40151 ( .A(n40521), .B(n40525), .Z(n40523) );
  XNOR U40152 ( .A(n40504), .B(n40501), .Z(n40514) );
  AND U40153 ( .A(n40526), .B(n40527), .Z(n40501) );
  XOR U40154 ( .A(n40528), .B(n40529), .Z(n40504) );
  AND U40155 ( .A(n40530), .B(n40531), .Z(n40529) );
  XOR U40156 ( .A(n40528), .B(n40532), .Z(n40530) );
  XNOR U40157 ( .A(n40465), .B(n40510), .Z(n40512) );
  XNOR U40158 ( .A(n40533), .B(n40534), .Z(n40465) );
  AND U40159 ( .A(n1044), .B(n40535), .Z(n40534) );
  XNOR U40160 ( .A(n40536), .B(n40537), .Z(n40535) );
  XOR U40161 ( .A(n40538), .B(n40539), .Z(n40510) );
  AND U40162 ( .A(n40540), .B(n40541), .Z(n40539) );
  XNOR U40163 ( .A(n40538), .B(n40526), .Z(n40541) );
  IV U40164 ( .A(n40476), .Z(n40526) );
  XNOR U40165 ( .A(n40542), .B(n40519), .Z(n40476) );
  XNOR U40166 ( .A(n40543), .B(n40525), .Z(n40519) );
  XOR U40167 ( .A(n40544), .B(n40545), .Z(n40525) );
  NOR U40168 ( .A(n40546), .B(n40547), .Z(n40545) );
  XNOR U40169 ( .A(n40544), .B(n40548), .Z(n40546) );
  XNOR U40170 ( .A(n40524), .B(n40516), .Z(n40543) );
  XOR U40171 ( .A(n40549), .B(n40550), .Z(n40516) );
  AND U40172 ( .A(n40551), .B(n40552), .Z(n40550) );
  XNOR U40173 ( .A(n40549), .B(n40553), .Z(n40551) );
  XNOR U40174 ( .A(n40554), .B(n40521), .Z(n40524) );
  XOR U40175 ( .A(n40555), .B(n40556), .Z(n40521) );
  AND U40176 ( .A(n40557), .B(n40558), .Z(n40556) );
  XOR U40177 ( .A(n40555), .B(n40559), .Z(n40557) );
  XNOR U40178 ( .A(n40560), .B(n40561), .Z(n40554) );
  NOR U40179 ( .A(n40562), .B(n40563), .Z(n40561) );
  XOR U40180 ( .A(n40560), .B(n40564), .Z(n40562) );
  XNOR U40181 ( .A(n40520), .B(n40527), .Z(n40542) );
  NOR U40182 ( .A(n40482), .B(n40565), .Z(n40527) );
  XOR U40183 ( .A(n40532), .B(n40531), .Z(n40520) );
  XNOR U40184 ( .A(n40566), .B(n40528), .Z(n40531) );
  XOR U40185 ( .A(n40567), .B(n40568), .Z(n40528) );
  AND U40186 ( .A(n40569), .B(n40570), .Z(n40568) );
  XOR U40187 ( .A(n40567), .B(n40571), .Z(n40569) );
  XNOR U40188 ( .A(n40572), .B(n40573), .Z(n40566) );
  NOR U40189 ( .A(n40574), .B(n40575), .Z(n40573) );
  XNOR U40190 ( .A(n40572), .B(n40576), .Z(n40574) );
  XOR U40191 ( .A(n40577), .B(n40578), .Z(n40532) );
  NOR U40192 ( .A(n40579), .B(n40580), .Z(n40578) );
  XNOR U40193 ( .A(n40577), .B(n40581), .Z(n40579) );
  XNOR U40194 ( .A(n40473), .B(n40538), .Z(n40540) );
  XNOR U40195 ( .A(n40582), .B(n40583), .Z(n40473) );
  AND U40196 ( .A(n1044), .B(n40584), .Z(n40583) );
  XNOR U40197 ( .A(n40585), .B(n40586), .Z(n40584) );
  AND U40198 ( .A(n40479), .B(n40482), .Z(n40538) );
  XOR U40199 ( .A(n40587), .B(n40565), .Z(n40482) );
  XNOR U40200 ( .A(p_input[2048]), .B(p_input[816]), .Z(n40565) );
  XOR U40201 ( .A(n40553), .B(n40552), .Z(n40587) );
  XNOR U40202 ( .A(n40588), .B(n40559), .Z(n40552) );
  XNOR U40203 ( .A(n40548), .B(n40547), .Z(n40559) );
  XOR U40204 ( .A(n40589), .B(n40544), .Z(n40547) );
  XNOR U40205 ( .A(n29266), .B(p_input[826]), .Z(n40544) );
  XNOR U40206 ( .A(p_input[2059]), .B(p_input[827]), .Z(n40589) );
  XOR U40207 ( .A(p_input[2060]), .B(p_input[828]), .Z(n40548) );
  XNOR U40208 ( .A(n40558), .B(n40549), .Z(n40588) );
  XNOR U40209 ( .A(n29494), .B(p_input[817]), .Z(n40549) );
  XOR U40210 ( .A(n40590), .B(n40564), .Z(n40558) );
  XNOR U40211 ( .A(p_input[2063]), .B(p_input[831]), .Z(n40564) );
  XOR U40212 ( .A(n40555), .B(n40563), .Z(n40590) );
  XOR U40213 ( .A(n40591), .B(n40560), .Z(n40563) );
  XOR U40214 ( .A(p_input[2061]), .B(p_input[829]), .Z(n40560) );
  XNOR U40215 ( .A(p_input[2062]), .B(p_input[830]), .Z(n40591) );
  XNOR U40216 ( .A(n29036), .B(p_input[825]), .Z(n40555) );
  XNOR U40217 ( .A(n40571), .B(n40570), .Z(n40553) );
  XNOR U40218 ( .A(n40592), .B(n40576), .Z(n40570) );
  XOR U40219 ( .A(p_input[2056]), .B(p_input[824]), .Z(n40576) );
  XOR U40220 ( .A(n40567), .B(n40575), .Z(n40592) );
  XOR U40221 ( .A(n40593), .B(n40572), .Z(n40575) );
  XOR U40222 ( .A(p_input[2054]), .B(p_input[822]), .Z(n40572) );
  XNOR U40223 ( .A(p_input[2055]), .B(p_input[823]), .Z(n40593) );
  XNOR U40224 ( .A(n29039), .B(p_input[818]), .Z(n40567) );
  XNOR U40225 ( .A(n40581), .B(n40580), .Z(n40571) );
  XOR U40226 ( .A(n40594), .B(n40577), .Z(n40580) );
  XOR U40227 ( .A(p_input[2051]), .B(p_input[819]), .Z(n40577) );
  XNOR U40228 ( .A(p_input[2052]), .B(p_input[820]), .Z(n40594) );
  XOR U40229 ( .A(p_input[2053]), .B(p_input[821]), .Z(n40581) );
  XNOR U40230 ( .A(n40595), .B(n40596), .Z(n40479) );
  AND U40231 ( .A(n1044), .B(n40597), .Z(n40596) );
  XNOR U40232 ( .A(n40598), .B(n40599), .Z(n1044) );
  AND U40233 ( .A(n40600), .B(n40601), .Z(n40599) );
  XOR U40234 ( .A(n40493), .B(n40598), .Z(n40601) );
  XNOR U40235 ( .A(n40602), .B(n40598), .Z(n40600) );
  XOR U40236 ( .A(n40603), .B(n40604), .Z(n40598) );
  AND U40237 ( .A(n40605), .B(n40606), .Z(n40604) );
  XOR U40238 ( .A(n40508), .B(n40603), .Z(n40606) );
  XOR U40239 ( .A(n40603), .B(n40509), .Z(n40605) );
  XOR U40240 ( .A(n40607), .B(n40608), .Z(n40603) );
  AND U40241 ( .A(n40609), .B(n40610), .Z(n40608) );
  XOR U40242 ( .A(n40536), .B(n40607), .Z(n40610) );
  XOR U40243 ( .A(n40607), .B(n40537), .Z(n40609) );
  XOR U40244 ( .A(n40611), .B(n40612), .Z(n40607) );
  AND U40245 ( .A(n40613), .B(n40614), .Z(n40612) );
  XOR U40246 ( .A(n40611), .B(n40585), .Z(n40614) );
  XNOR U40247 ( .A(n40615), .B(n40616), .Z(n40439) );
  AND U40248 ( .A(n1048), .B(n40617), .Z(n40616) );
  XNOR U40249 ( .A(n40618), .B(n40619), .Z(n1048) );
  AND U40250 ( .A(n40620), .B(n40621), .Z(n40619) );
  XOR U40251 ( .A(n40618), .B(n40449), .Z(n40621) );
  XNOR U40252 ( .A(n40618), .B(n40409), .Z(n40620) );
  XOR U40253 ( .A(n40622), .B(n40623), .Z(n40618) );
  AND U40254 ( .A(n40624), .B(n40625), .Z(n40623) );
  XOR U40255 ( .A(n40622), .B(n40417), .Z(n40624) );
  XOR U40256 ( .A(n40626), .B(n40627), .Z(n40400) );
  AND U40257 ( .A(n1052), .B(n40617), .Z(n40627) );
  XNOR U40258 ( .A(n40615), .B(n40626), .Z(n40617) );
  XNOR U40259 ( .A(n40628), .B(n40629), .Z(n1052) );
  AND U40260 ( .A(n40630), .B(n40631), .Z(n40629) );
  XNOR U40261 ( .A(n40632), .B(n40628), .Z(n40631) );
  IV U40262 ( .A(n40449), .Z(n40632) );
  XOR U40263 ( .A(n40602), .B(n40633), .Z(n40449) );
  AND U40264 ( .A(n1055), .B(n40634), .Z(n40633) );
  XOR U40265 ( .A(n40492), .B(n40489), .Z(n40634) );
  IV U40266 ( .A(n40602), .Z(n40492) );
  XNOR U40267 ( .A(n40409), .B(n40628), .Z(n40630) );
  XOR U40268 ( .A(n40635), .B(n40636), .Z(n40409) );
  AND U40269 ( .A(n1071), .B(n40637), .Z(n40636) );
  XOR U40270 ( .A(n40622), .B(n40638), .Z(n40628) );
  AND U40271 ( .A(n40639), .B(n40625), .Z(n40638) );
  XNOR U40272 ( .A(n40459), .B(n40622), .Z(n40625) );
  XOR U40273 ( .A(n40509), .B(n40640), .Z(n40459) );
  AND U40274 ( .A(n1055), .B(n40641), .Z(n40640) );
  XOR U40275 ( .A(n40505), .B(n40509), .Z(n40641) );
  XNOR U40276 ( .A(n40642), .B(n40622), .Z(n40639) );
  IV U40277 ( .A(n40417), .Z(n40642) );
  XOR U40278 ( .A(n40643), .B(n40644), .Z(n40417) );
  AND U40279 ( .A(n1071), .B(n40645), .Z(n40644) );
  XOR U40280 ( .A(n40646), .B(n40647), .Z(n40622) );
  AND U40281 ( .A(n40648), .B(n40649), .Z(n40647) );
  XNOR U40282 ( .A(n40469), .B(n40646), .Z(n40649) );
  XOR U40283 ( .A(n40537), .B(n40650), .Z(n40469) );
  AND U40284 ( .A(n1055), .B(n40651), .Z(n40650) );
  XOR U40285 ( .A(n40533), .B(n40537), .Z(n40651) );
  XOR U40286 ( .A(n40646), .B(n40426), .Z(n40648) );
  XOR U40287 ( .A(n40652), .B(n40653), .Z(n40426) );
  AND U40288 ( .A(n1071), .B(n40654), .Z(n40653) );
  XOR U40289 ( .A(n40655), .B(n40656), .Z(n40646) );
  AND U40290 ( .A(n40657), .B(n40658), .Z(n40656) );
  XNOR U40291 ( .A(n40655), .B(n40477), .Z(n40658) );
  XOR U40292 ( .A(n40586), .B(n40659), .Z(n40477) );
  AND U40293 ( .A(n1055), .B(n40660), .Z(n40659) );
  XOR U40294 ( .A(n40582), .B(n40586), .Z(n40660) );
  XNOR U40295 ( .A(n40661), .B(n40655), .Z(n40657) );
  IV U40296 ( .A(n40436), .Z(n40661) );
  XOR U40297 ( .A(n40662), .B(n40663), .Z(n40436) );
  AND U40298 ( .A(n1071), .B(n40664), .Z(n40663) );
  AND U40299 ( .A(n40626), .B(n40615), .Z(n40655) );
  XNOR U40300 ( .A(n40665), .B(n40666), .Z(n40615) );
  AND U40301 ( .A(n1055), .B(n40597), .Z(n40666) );
  XNOR U40302 ( .A(n40595), .B(n40665), .Z(n40597) );
  XNOR U40303 ( .A(n40667), .B(n40668), .Z(n1055) );
  AND U40304 ( .A(n40669), .B(n40670), .Z(n40668) );
  XNOR U40305 ( .A(n40667), .B(n40489), .Z(n40670) );
  IV U40306 ( .A(n40493), .Z(n40489) );
  XOR U40307 ( .A(n40671), .B(n40672), .Z(n40493) );
  AND U40308 ( .A(n1059), .B(n40673), .Z(n40672) );
  XOR U40309 ( .A(n40674), .B(n40671), .Z(n40673) );
  XNOR U40310 ( .A(n40667), .B(n40602), .Z(n40669) );
  XOR U40311 ( .A(n40675), .B(n40676), .Z(n40602) );
  AND U40312 ( .A(n1067), .B(n40637), .Z(n40676) );
  XOR U40313 ( .A(n40635), .B(n40675), .Z(n40637) );
  XOR U40314 ( .A(n40677), .B(n40678), .Z(n40667) );
  AND U40315 ( .A(n40679), .B(n40680), .Z(n40678) );
  XNOR U40316 ( .A(n40677), .B(n40505), .Z(n40680) );
  IV U40317 ( .A(n40508), .Z(n40505) );
  XOR U40318 ( .A(n40681), .B(n40682), .Z(n40508) );
  AND U40319 ( .A(n1059), .B(n40683), .Z(n40682) );
  XOR U40320 ( .A(n40684), .B(n40681), .Z(n40683) );
  XOR U40321 ( .A(n40509), .B(n40677), .Z(n40679) );
  XOR U40322 ( .A(n40685), .B(n40686), .Z(n40509) );
  AND U40323 ( .A(n1067), .B(n40645), .Z(n40686) );
  XOR U40324 ( .A(n40685), .B(n40643), .Z(n40645) );
  XOR U40325 ( .A(n40687), .B(n40688), .Z(n40677) );
  AND U40326 ( .A(n40689), .B(n40690), .Z(n40688) );
  XNOR U40327 ( .A(n40687), .B(n40533), .Z(n40690) );
  IV U40328 ( .A(n40536), .Z(n40533) );
  XOR U40329 ( .A(n40691), .B(n40692), .Z(n40536) );
  AND U40330 ( .A(n1059), .B(n40693), .Z(n40692) );
  XNOR U40331 ( .A(n40694), .B(n40691), .Z(n40693) );
  XOR U40332 ( .A(n40537), .B(n40687), .Z(n40689) );
  XOR U40333 ( .A(n40695), .B(n40696), .Z(n40537) );
  AND U40334 ( .A(n1067), .B(n40654), .Z(n40696) );
  XOR U40335 ( .A(n40695), .B(n40652), .Z(n40654) );
  XOR U40336 ( .A(n40611), .B(n40697), .Z(n40687) );
  AND U40337 ( .A(n40613), .B(n40698), .Z(n40697) );
  XNOR U40338 ( .A(n40611), .B(n40582), .Z(n40698) );
  IV U40339 ( .A(n40585), .Z(n40582) );
  XOR U40340 ( .A(n40699), .B(n40700), .Z(n40585) );
  AND U40341 ( .A(n1059), .B(n40701), .Z(n40700) );
  XOR U40342 ( .A(n40702), .B(n40699), .Z(n40701) );
  XOR U40343 ( .A(n40586), .B(n40611), .Z(n40613) );
  XOR U40344 ( .A(n40703), .B(n40704), .Z(n40586) );
  AND U40345 ( .A(n1067), .B(n40664), .Z(n40704) );
  XOR U40346 ( .A(n40703), .B(n40662), .Z(n40664) );
  AND U40347 ( .A(n40665), .B(n40595), .Z(n40611) );
  XNOR U40348 ( .A(n40705), .B(n40706), .Z(n40595) );
  AND U40349 ( .A(n1059), .B(n40707), .Z(n40706) );
  XNOR U40350 ( .A(n40708), .B(n40705), .Z(n40707) );
  XNOR U40351 ( .A(n40709), .B(n40710), .Z(n1059) );
  AND U40352 ( .A(n40711), .B(n40712), .Z(n40710) );
  XOR U40353 ( .A(n40674), .B(n40709), .Z(n40712) );
  AND U40354 ( .A(n40713), .B(n40714), .Z(n40674) );
  XNOR U40355 ( .A(n40671), .B(n40709), .Z(n40711) );
  XNOR U40356 ( .A(n40715), .B(n40716), .Z(n40671) );
  AND U40357 ( .A(n1063), .B(n40717), .Z(n40716) );
  XNOR U40358 ( .A(n40718), .B(n40719), .Z(n40717) );
  XOR U40359 ( .A(n40720), .B(n40721), .Z(n40709) );
  AND U40360 ( .A(n40722), .B(n40723), .Z(n40721) );
  XNOR U40361 ( .A(n40720), .B(n40713), .Z(n40723) );
  IV U40362 ( .A(n40684), .Z(n40713) );
  XOR U40363 ( .A(n40724), .B(n40725), .Z(n40684) );
  XOR U40364 ( .A(n40726), .B(n40714), .Z(n40725) );
  AND U40365 ( .A(n40694), .B(n40727), .Z(n40714) );
  AND U40366 ( .A(n40728), .B(n40729), .Z(n40726) );
  XOR U40367 ( .A(n40730), .B(n40724), .Z(n40728) );
  XNOR U40368 ( .A(n40681), .B(n40720), .Z(n40722) );
  XNOR U40369 ( .A(n40731), .B(n40732), .Z(n40681) );
  AND U40370 ( .A(n1063), .B(n40733), .Z(n40732) );
  XNOR U40371 ( .A(n40734), .B(n40735), .Z(n40733) );
  XOR U40372 ( .A(n40736), .B(n40737), .Z(n40720) );
  AND U40373 ( .A(n40738), .B(n40739), .Z(n40737) );
  XNOR U40374 ( .A(n40736), .B(n40694), .Z(n40739) );
  XOR U40375 ( .A(n40740), .B(n40729), .Z(n40694) );
  XNOR U40376 ( .A(n40741), .B(n40724), .Z(n40729) );
  XOR U40377 ( .A(n40742), .B(n40743), .Z(n40724) );
  AND U40378 ( .A(n40744), .B(n40745), .Z(n40743) );
  XOR U40379 ( .A(n40746), .B(n40742), .Z(n40744) );
  XNOR U40380 ( .A(n40747), .B(n40748), .Z(n40741) );
  AND U40381 ( .A(n40749), .B(n40750), .Z(n40748) );
  XOR U40382 ( .A(n40747), .B(n40751), .Z(n40749) );
  XNOR U40383 ( .A(n40730), .B(n40727), .Z(n40740) );
  AND U40384 ( .A(n40752), .B(n40753), .Z(n40727) );
  XOR U40385 ( .A(n40754), .B(n40755), .Z(n40730) );
  AND U40386 ( .A(n40756), .B(n40757), .Z(n40755) );
  XOR U40387 ( .A(n40754), .B(n40758), .Z(n40756) );
  XNOR U40388 ( .A(n40691), .B(n40736), .Z(n40738) );
  XNOR U40389 ( .A(n40759), .B(n40760), .Z(n40691) );
  AND U40390 ( .A(n1063), .B(n40761), .Z(n40760) );
  XNOR U40391 ( .A(n40762), .B(n40763), .Z(n40761) );
  XOR U40392 ( .A(n40764), .B(n40765), .Z(n40736) );
  AND U40393 ( .A(n40766), .B(n40767), .Z(n40765) );
  XNOR U40394 ( .A(n40764), .B(n40752), .Z(n40767) );
  IV U40395 ( .A(n40702), .Z(n40752) );
  XNOR U40396 ( .A(n40768), .B(n40745), .Z(n40702) );
  XNOR U40397 ( .A(n40769), .B(n40751), .Z(n40745) );
  XOR U40398 ( .A(n40770), .B(n40771), .Z(n40751) );
  NOR U40399 ( .A(n40772), .B(n40773), .Z(n40771) );
  XNOR U40400 ( .A(n40770), .B(n40774), .Z(n40772) );
  XNOR U40401 ( .A(n40750), .B(n40742), .Z(n40769) );
  XOR U40402 ( .A(n40775), .B(n40776), .Z(n40742) );
  AND U40403 ( .A(n40777), .B(n40778), .Z(n40776) );
  XNOR U40404 ( .A(n40775), .B(n40779), .Z(n40777) );
  XNOR U40405 ( .A(n40780), .B(n40747), .Z(n40750) );
  XOR U40406 ( .A(n40781), .B(n40782), .Z(n40747) );
  AND U40407 ( .A(n40783), .B(n40784), .Z(n40782) );
  XOR U40408 ( .A(n40781), .B(n40785), .Z(n40783) );
  XNOR U40409 ( .A(n40786), .B(n40787), .Z(n40780) );
  NOR U40410 ( .A(n40788), .B(n40789), .Z(n40787) );
  XOR U40411 ( .A(n40786), .B(n40790), .Z(n40788) );
  XNOR U40412 ( .A(n40746), .B(n40753), .Z(n40768) );
  NOR U40413 ( .A(n40708), .B(n40791), .Z(n40753) );
  XOR U40414 ( .A(n40758), .B(n40757), .Z(n40746) );
  XNOR U40415 ( .A(n40792), .B(n40754), .Z(n40757) );
  XOR U40416 ( .A(n40793), .B(n40794), .Z(n40754) );
  AND U40417 ( .A(n40795), .B(n40796), .Z(n40794) );
  XOR U40418 ( .A(n40793), .B(n40797), .Z(n40795) );
  XNOR U40419 ( .A(n40798), .B(n40799), .Z(n40792) );
  NOR U40420 ( .A(n40800), .B(n40801), .Z(n40799) );
  XNOR U40421 ( .A(n40798), .B(n40802), .Z(n40800) );
  XOR U40422 ( .A(n40803), .B(n40804), .Z(n40758) );
  NOR U40423 ( .A(n40805), .B(n40806), .Z(n40804) );
  XNOR U40424 ( .A(n40803), .B(n40807), .Z(n40805) );
  XNOR U40425 ( .A(n40699), .B(n40764), .Z(n40766) );
  XNOR U40426 ( .A(n40808), .B(n40809), .Z(n40699) );
  AND U40427 ( .A(n1063), .B(n40810), .Z(n40809) );
  XNOR U40428 ( .A(n40811), .B(n40812), .Z(n40810) );
  AND U40429 ( .A(n40705), .B(n40708), .Z(n40764) );
  XOR U40430 ( .A(n40813), .B(n40791), .Z(n40708) );
  XNOR U40431 ( .A(p_input[2048]), .B(p_input[832]), .Z(n40791) );
  XOR U40432 ( .A(n40779), .B(n40778), .Z(n40813) );
  XNOR U40433 ( .A(n40814), .B(n40785), .Z(n40778) );
  XNOR U40434 ( .A(n40774), .B(n40773), .Z(n40785) );
  XOR U40435 ( .A(n40815), .B(n40770), .Z(n40773) );
  XNOR U40436 ( .A(n29266), .B(p_input[842]), .Z(n40770) );
  XNOR U40437 ( .A(p_input[2059]), .B(p_input[843]), .Z(n40815) );
  XOR U40438 ( .A(p_input[2060]), .B(p_input[844]), .Z(n40774) );
  XNOR U40439 ( .A(n40784), .B(n40775), .Z(n40814) );
  XNOR U40440 ( .A(n29494), .B(p_input[833]), .Z(n40775) );
  XOR U40441 ( .A(n40816), .B(n40790), .Z(n40784) );
  XNOR U40442 ( .A(p_input[2063]), .B(p_input[847]), .Z(n40790) );
  XOR U40443 ( .A(n40781), .B(n40789), .Z(n40816) );
  XOR U40444 ( .A(n40817), .B(n40786), .Z(n40789) );
  XOR U40445 ( .A(p_input[2061]), .B(p_input[845]), .Z(n40786) );
  XNOR U40446 ( .A(p_input[2062]), .B(p_input[846]), .Z(n40817) );
  XNOR U40447 ( .A(n29036), .B(p_input[841]), .Z(n40781) );
  XNOR U40448 ( .A(n40797), .B(n40796), .Z(n40779) );
  XNOR U40449 ( .A(n40818), .B(n40802), .Z(n40796) );
  XOR U40450 ( .A(p_input[2056]), .B(p_input[840]), .Z(n40802) );
  XOR U40451 ( .A(n40793), .B(n40801), .Z(n40818) );
  XOR U40452 ( .A(n40819), .B(n40798), .Z(n40801) );
  XOR U40453 ( .A(p_input[2054]), .B(p_input[838]), .Z(n40798) );
  XNOR U40454 ( .A(p_input[2055]), .B(p_input[839]), .Z(n40819) );
  XNOR U40455 ( .A(n29039), .B(p_input[834]), .Z(n40793) );
  XNOR U40456 ( .A(n40807), .B(n40806), .Z(n40797) );
  XOR U40457 ( .A(n40820), .B(n40803), .Z(n40806) );
  XOR U40458 ( .A(p_input[2051]), .B(p_input[835]), .Z(n40803) );
  XNOR U40459 ( .A(p_input[2052]), .B(p_input[836]), .Z(n40820) );
  XOR U40460 ( .A(p_input[2053]), .B(p_input[837]), .Z(n40807) );
  XNOR U40461 ( .A(n40821), .B(n40822), .Z(n40705) );
  AND U40462 ( .A(n1063), .B(n40823), .Z(n40822) );
  XNOR U40463 ( .A(n40824), .B(n40825), .Z(n1063) );
  AND U40464 ( .A(n40826), .B(n40827), .Z(n40825) );
  XOR U40465 ( .A(n40719), .B(n40824), .Z(n40827) );
  XNOR U40466 ( .A(n40828), .B(n40824), .Z(n40826) );
  XOR U40467 ( .A(n40829), .B(n40830), .Z(n40824) );
  AND U40468 ( .A(n40831), .B(n40832), .Z(n40830) );
  XOR U40469 ( .A(n40734), .B(n40829), .Z(n40832) );
  XOR U40470 ( .A(n40829), .B(n40735), .Z(n40831) );
  XOR U40471 ( .A(n40833), .B(n40834), .Z(n40829) );
  AND U40472 ( .A(n40835), .B(n40836), .Z(n40834) );
  XOR U40473 ( .A(n40762), .B(n40833), .Z(n40836) );
  XOR U40474 ( .A(n40833), .B(n40763), .Z(n40835) );
  XOR U40475 ( .A(n40837), .B(n40838), .Z(n40833) );
  AND U40476 ( .A(n40839), .B(n40840), .Z(n40838) );
  XOR U40477 ( .A(n40837), .B(n40811), .Z(n40840) );
  XNOR U40478 ( .A(n40841), .B(n40842), .Z(n40665) );
  AND U40479 ( .A(n1067), .B(n40843), .Z(n40842) );
  XNOR U40480 ( .A(n40844), .B(n40845), .Z(n1067) );
  AND U40481 ( .A(n40846), .B(n40847), .Z(n40845) );
  XOR U40482 ( .A(n40844), .B(n40675), .Z(n40847) );
  XNOR U40483 ( .A(n40844), .B(n40635), .Z(n40846) );
  XOR U40484 ( .A(n40848), .B(n40849), .Z(n40844) );
  AND U40485 ( .A(n40850), .B(n40851), .Z(n40849) );
  XOR U40486 ( .A(n40848), .B(n40643), .Z(n40850) );
  XOR U40487 ( .A(n40852), .B(n40853), .Z(n40626) );
  AND U40488 ( .A(n1071), .B(n40843), .Z(n40853) );
  XNOR U40489 ( .A(n40841), .B(n40852), .Z(n40843) );
  XNOR U40490 ( .A(n40854), .B(n40855), .Z(n1071) );
  AND U40491 ( .A(n40856), .B(n40857), .Z(n40855) );
  XNOR U40492 ( .A(n40858), .B(n40854), .Z(n40857) );
  IV U40493 ( .A(n40675), .Z(n40858) );
  XOR U40494 ( .A(n40828), .B(n40859), .Z(n40675) );
  AND U40495 ( .A(n1074), .B(n40860), .Z(n40859) );
  XOR U40496 ( .A(n40718), .B(n40715), .Z(n40860) );
  IV U40497 ( .A(n40828), .Z(n40718) );
  XNOR U40498 ( .A(n40635), .B(n40854), .Z(n40856) );
  XOR U40499 ( .A(n40861), .B(n40862), .Z(n40635) );
  AND U40500 ( .A(n1090), .B(n40863), .Z(n40862) );
  XOR U40501 ( .A(n40848), .B(n40864), .Z(n40854) );
  AND U40502 ( .A(n40865), .B(n40851), .Z(n40864) );
  XNOR U40503 ( .A(n40685), .B(n40848), .Z(n40851) );
  XOR U40504 ( .A(n40735), .B(n40866), .Z(n40685) );
  AND U40505 ( .A(n1074), .B(n40867), .Z(n40866) );
  XOR U40506 ( .A(n40731), .B(n40735), .Z(n40867) );
  XNOR U40507 ( .A(n40868), .B(n40848), .Z(n40865) );
  IV U40508 ( .A(n40643), .Z(n40868) );
  XOR U40509 ( .A(n40869), .B(n40870), .Z(n40643) );
  AND U40510 ( .A(n1090), .B(n40871), .Z(n40870) );
  XOR U40511 ( .A(n40872), .B(n40873), .Z(n40848) );
  AND U40512 ( .A(n40874), .B(n40875), .Z(n40873) );
  XNOR U40513 ( .A(n40695), .B(n40872), .Z(n40875) );
  XOR U40514 ( .A(n40763), .B(n40876), .Z(n40695) );
  AND U40515 ( .A(n1074), .B(n40877), .Z(n40876) );
  XOR U40516 ( .A(n40759), .B(n40763), .Z(n40877) );
  XOR U40517 ( .A(n40872), .B(n40652), .Z(n40874) );
  XOR U40518 ( .A(n40878), .B(n40879), .Z(n40652) );
  AND U40519 ( .A(n1090), .B(n40880), .Z(n40879) );
  XOR U40520 ( .A(n40881), .B(n40882), .Z(n40872) );
  AND U40521 ( .A(n40883), .B(n40884), .Z(n40882) );
  XNOR U40522 ( .A(n40881), .B(n40703), .Z(n40884) );
  XOR U40523 ( .A(n40812), .B(n40885), .Z(n40703) );
  AND U40524 ( .A(n1074), .B(n40886), .Z(n40885) );
  XOR U40525 ( .A(n40808), .B(n40812), .Z(n40886) );
  XNOR U40526 ( .A(n40887), .B(n40881), .Z(n40883) );
  IV U40527 ( .A(n40662), .Z(n40887) );
  XOR U40528 ( .A(n40888), .B(n40889), .Z(n40662) );
  AND U40529 ( .A(n1090), .B(n40890), .Z(n40889) );
  AND U40530 ( .A(n40852), .B(n40841), .Z(n40881) );
  XNOR U40531 ( .A(n40891), .B(n40892), .Z(n40841) );
  AND U40532 ( .A(n1074), .B(n40823), .Z(n40892) );
  XNOR U40533 ( .A(n40821), .B(n40891), .Z(n40823) );
  XNOR U40534 ( .A(n40893), .B(n40894), .Z(n1074) );
  AND U40535 ( .A(n40895), .B(n40896), .Z(n40894) );
  XNOR U40536 ( .A(n40893), .B(n40715), .Z(n40896) );
  IV U40537 ( .A(n40719), .Z(n40715) );
  XOR U40538 ( .A(n40897), .B(n40898), .Z(n40719) );
  AND U40539 ( .A(n1078), .B(n40899), .Z(n40898) );
  XOR U40540 ( .A(n40900), .B(n40897), .Z(n40899) );
  XNOR U40541 ( .A(n40893), .B(n40828), .Z(n40895) );
  XOR U40542 ( .A(n40901), .B(n40902), .Z(n40828) );
  AND U40543 ( .A(n1086), .B(n40863), .Z(n40902) );
  XOR U40544 ( .A(n40861), .B(n40901), .Z(n40863) );
  XOR U40545 ( .A(n40903), .B(n40904), .Z(n40893) );
  AND U40546 ( .A(n40905), .B(n40906), .Z(n40904) );
  XNOR U40547 ( .A(n40903), .B(n40731), .Z(n40906) );
  IV U40548 ( .A(n40734), .Z(n40731) );
  XOR U40549 ( .A(n40907), .B(n40908), .Z(n40734) );
  AND U40550 ( .A(n1078), .B(n40909), .Z(n40908) );
  XOR U40551 ( .A(n40910), .B(n40907), .Z(n40909) );
  XOR U40552 ( .A(n40735), .B(n40903), .Z(n40905) );
  XOR U40553 ( .A(n40911), .B(n40912), .Z(n40735) );
  AND U40554 ( .A(n1086), .B(n40871), .Z(n40912) );
  XOR U40555 ( .A(n40911), .B(n40869), .Z(n40871) );
  XOR U40556 ( .A(n40913), .B(n40914), .Z(n40903) );
  AND U40557 ( .A(n40915), .B(n40916), .Z(n40914) );
  XNOR U40558 ( .A(n40913), .B(n40759), .Z(n40916) );
  IV U40559 ( .A(n40762), .Z(n40759) );
  XOR U40560 ( .A(n40917), .B(n40918), .Z(n40762) );
  AND U40561 ( .A(n1078), .B(n40919), .Z(n40918) );
  XNOR U40562 ( .A(n40920), .B(n40917), .Z(n40919) );
  XOR U40563 ( .A(n40763), .B(n40913), .Z(n40915) );
  XOR U40564 ( .A(n40921), .B(n40922), .Z(n40763) );
  AND U40565 ( .A(n1086), .B(n40880), .Z(n40922) );
  XOR U40566 ( .A(n40921), .B(n40878), .Z(n40880) );
  XOR U40567 ( .A(n40837), .B(n40923), .Z(n40913) );
  AND U40568 ( .A(n40839), .B(n40924), .Z(n40923) );
  XNOR U40569 ( .A(n40837), .B(n40808), .Z(n40924) );
  IV U40570 ( .A(n40811), .Z(n40808) );
  XOR U40571 ( .A(n40925), .B(n40926), .Z(n40811) );
  AND U40572 ( .A(n1078), .B(n40927), .Z(n40926) );
  XOR U40573 ( .A(n40928), .B(n40925), .Z(n40927) );
  XOR U40574 ( .A(n40812), .B(n40837), .Z(n40839) );
  XOR U40575 ( .A(n40929), .B(n40930), .Z(n40812) );
  AND U40576 ( .A(n1086), .B(n40890), .Z(n40930) );
  XOR U40577 ( .A(n40929), .B(n40888), .Z(n40890) );
  AND U40578 ( .A(n40891), .B(n40821), .Z(n40837) );
  XNOR U40579 ( .A(n40931), .B(n40932), .Z(n40821) );
  AND U40580 ( .A(n1078), .B(n40933), .Z(n40932) );
  XNOR U40581 ( .A(n40934), .B(n40931), .Z(n40933) );
  XNOR U40582 ( .A(n40935), .B(n40936), .Z(n1078) );
  AND U40583 ( .A(n40937), .B(n40938), .Z(n40936) );
  XOR U40584 ( .A(n40900), .B(n40935), .Z(n40938) );
  AND U40585 ( .A(n40939), .B(n40940), .Z(n40900) );
  XNOR U40586 ( .A(n40897), .B(n40935), .Z(n40937) );
  XNOR U40587 ( .A(n40941), .B(n40942), .Z(n40897) );
  AND U40588 ( .A(n1082), .B(n40943), .Z(n40942) );
  XNOR U40589 ( .A(n40944), .B(n40945), .Z(n40943) );
  XOR U40590 ( .A(n40946), .B(n40947), .Z(n40935) );
  AND U40591 ( .A(n40948), .B(n40949), .Z(n40947) );
  XNOR U40592 ( .A(n40946), .B(n40939), .Z(n40949) );
  IV U40593 ( .A(n40910), .Z(n40939) );
  XOR U40594 ( .A(n40950), .B(n40951), .Z(n40910) );
  XOR U40595 ( .A(n40952), .B(n40940), .Z(n40951) );
  AND U40596 ( .A(n40920), .B(n40953), .Z(n40940) );
  AND U40597 ( .A(n40954), .B(n40955), .Z(n40952) );
  XOR U40598 ( .A(n40956), .B(n40950), .Z(n40954) );
  XNOR U40599 ( .A(n40907), .B(n40946), .Z(n40948) );
  XNOR U40600 ( .A(n40957), .B(n40958), .Z(n40907) );
  AND U40601 ( .A(n1082), .B(n40959), .Z(n40958) );
  XNOR U40602 ( .A(n40960), .B(n40961), .Z(n40959) );
  XOR U40603 ( .A(n40962), .B(n40963), .Z(n40946) );
  AND U40604 ( .A(n40964), .B(n40965), .Z(n40963) );
  XNOR U40605 ( .A(n40962), .B(n40920), .Z(n40965) );
  XOR U40606 ( .A(n40966), .B(n40955), .Z(n40920) );
  XNOR U40607 ( .A(n40967), .B(n40950), .Z(n40955) );
  XOR U40608 ( .A(n40968), .B(n40969), .Z(n40950) );
  AND U40609 ( .A(n40970), .B(n40971), .Z(n40969) );
  XOR U40610 ( .A(n40972), .B(n40968), .Z(n40970) );
  XNOR U40611 ( .A(n40973), .B(n40974), .Z(n40967) );
  AND U40612 ( .A(n40975), .B(n40976), .Z(n40974) );
  XOR U40613 ( .A(n40973), .B(n40977), .Z(n40975) );
  XNOR U40614 ( .A(n40956), .B(n40953), .Z(n40966) );
  AND U40615 ( .A(n40978), .B(n40979), .Z(n40953) );
  XOR U40616 ( .A(n40980), .B(n40981), .Z(n40956) );
  AND U40617 ( .A(n40982), .B(n40983), .Z(n40981) );
  XOR U40618 ( .A(n40980), .B(n40984), .Z(n40982) );
  XNOR U40619 ( .A(n40917), .B(n40962), .Z(n40964) );
  XNOR U40620 ( .A(n40985), .B(n40986), .Z(n40917) );
  AND U40621 ( .A(n1082), .B(n40987), .Z(n40986) );
  XNOR U40622 ( .A(n40988), .B(n40989), .Z(n40987) );
  XOR U40623 ( .A(n40990), .B(n40991), .Z(n40962) );
  AND U40624 ( .A(n40992), .B(n40993), .Z(n40991) );
  XNOR U40625 ( .A(n40990), .B(n40978), .Z(n40993) );
  IV U40626 ( .A(n40928), .Z(n40978) );
  XNOR U40627 ( .A(n40994), .B(n40971), .Z(n40928) );
  XNOR U40628 ( .A(n40995), .B(n40977), .Z(n40971) );
  XOR U40629 ( .A(n40996), .B(n40997), .Z(n40977) );
  NOR U40630 ( .A(n40998), .B(n40999), .Z(n40997) );
  XNOR U40631 ( .A(n40996), .B(n41000), .Z(n40998) );
  XNOR U40632 ( .A(n40976), .B(n40968), .Z(n40995) );
  XOR U40633 ( .A(n41001), .B(n41002), .Z(n40968) );
  AND U40634 ( .A(n41003), .B(n41004), .Z(n41002) );
  XNOR U40635 ( .A(n41001), .B(n41005), .Z(n41003) );
  XNOR U40636 ( .A(n41006), .B(n40973), .Z(n40976) );
  XOR U40637 ( .A(n41007), .B(n41008), .Z(n40973) );
  AND U40638 ( .A(n41009), .B(n41010), .Z(n41008) );
  XOR U40639 ( .A(n41007), .B(n41011), .Z(n41009) );
  XNOR U40640 ( .A(n41012), .B(n41013), .Z(n41006) );
  NOR U40641 ( .A(n41014), .B(n41015), .Z(n41013) );
  XOR U40642 ( .A(n41012), .B(n41016), .Z(n41014) );
  XNOR U40643 ( .A(n40972), .B(n40979), .Z(n40994) );
  NOR U40644 ( .A(n40934), .B(n41017), .Z(n40979) );
  XOR U40645 ( .A(n40984), .B(n40983), .Z(n40972) );
  XNOR U40646 ( .A(n41018), .B(n40980), .Z(n40983) );
  XOR U40647 ( .A(n41019), .B(n41020), .Z(n40980) );
  AND U40648 ( .A(n41021), .B(n41022), .Z(n41020) );
  XOR U40649 ( .A(n41019), .B(n41023), .Z(n41021) );
  XNOR U40650 ( .A(n41024), .B(n41025), .Z(n41018) );
  NOR U40651 ( .A(n41026), .B(n41027), .Z(n41025) );
  XNOR U40652 ( .A(n41024), .B(n41028), .Z(n41026) );
  XOR U40653 ( .A(n41029), .B(n41030), .Z(n40984) );
  NOR U40654 ( .A(n41031), .B(n41032), .Z(n41030) );
  XNOR U40655 ( .A(n41029), .B(n41033), .Z(n41031) );
  XNOR U40656 ( .A(n40925), .B(n40990), .Z(n40992) );
  XNOR U40657 ( .A(n41034), .B(n41035), .Z(n40925) );
  AND U40658 ( .A(n1082), .B(n41036), .Z(n41035) );
  XNOR U40659 ( .A(n41037), .B(n41038), .Z(n41036) );
  AND U40660 ( .A(n40931), .B(n40934), .Z(n40990) );
  XOR U40661 ( .A(n41039), .B(n41017), .Z(n40934) );
  XNOR U40662 ( .A(p_input[2048]), .B(p_input[848]), .Z(n41017) );
  XOR U40663 ( .A(n41005), .B(n41004), .Z(n41039) );
  XNOR U40664 ( .A(n41040), .B(n41011), .Z(n41004) );
  XNOR U40665 ( .A(n41000), .B(n40999), .Z(n41011) );
  XOR U40666 ( .A(n41041), .B(n40996), .Z(n40999) );
  XNOR U40667 ( .A(n29266), .B(p_input[858]), .Z(n40996) );
  XNOR U40668 ( .A(p_input[2059]), .B(p_input[859]), .Z(n41041) );
  XOR U40669 ( .A(p_input[2060]), .B(p_input[860]), .Z(n41000) );
  XNOR U40670 ( .A(n41010), .B(n41001), .Z(n41040) );
  XNOR U40671 ( .A(n29494), .B(p_input[849]), .Z(n41001) );
  XOR U40672 ( .A(n41042), .B(n41016), .Z(n41010) );
  XNOR U40673 ( .A(p_input[2063]), .B(p_input[863]), .Z(n41016) );
  XOR U40674 ( .A(n41007), .B(n41015), .Z(n41042) );
  XOR U40675 ( .A(n41043), .B(n41012), .Z(n41015) );
  XOR U40676 ( .A(p_input[2061]), .B(p_input[861]), .Z(n41012) );
  XNOR U40677 ( .A(p_input[2062]), .B(p_input[862]), .Z(n41043) );
  XNOR U40678 ( .A(n29036), .B(p_input[857]), .Z(n41007) );
  XNOR U40679 ( .A(n41023), .B(n41022), .Z(n41005) );
  XNOR U40680 ( .A(n41044), .B(n41028), .Z(n41022) );
  XOR U40681 ( .A(p_input[2056]), .B(p_input[856]), .Z(n41028) );
  XOR U40682 ( .A(n41019), .B(n41027), .Z(n41044) );
  XOR U40683 ( .A(n41045), .B(n41024), .Z(n41027) );
  XOR U40684 ( .A(p_input[2054]), .B(p_input[854]), .Z(n41024) );
  XNOR U40685 ( .A(p_input[2055]), .B(p_input[855]), .Z(n41045) );
  XNOR U40686 ( .A(n29039), .B(p_input[850]), .Z(n41019) );
  XNOR U40687 ( .A(n41033), .B(n41032), .Z(n41023) );
  XOR U40688 ( .A(n41046), .B(n41029), .Z(n41032) );
  XOR U40689 ( .A(p_input[2051]), .B(p_input[851]), .Z(n41029) );
  XNOR U40690 ( .A(p_input[2052]), .B(p_input[852]), .Z(n41046) );
  XOR U40691 ( .A(p_input[2053]), .B(p_input[853]), .Z(n41033) );
  XNOR U40692 ( .A(n41047), .B(n41048), .Z(n40931) );
  AND U40693 ( .A(n1082), .B(n41049), .Z(n41048) );
  XNOR U40694 ( .A(n41050), .B(n41051), .Z(n1082) );
  AND U40695 ( .A(n41052), .B(n41053), .Z(n41051) );
  XOR U40696 ( .A(n40945), .B(n41050), .Z(n41053) );
  XNOR U40697 ( .A(n41054), .B(n41050), .Z(n41052) );
  XOR U40698 ( .A(n41055), .B(n41056), .Z(n41050) );
  AND U40699 ( .A(n41057), .B(n41058), .Z(n41056) );
  XOR U40700 ( .A(n40960), .B(n41055), .Z(n41058) );
  XOR U40701 ( .A(n41055), .B(n40961), .Z(n41057) );
  XOR U40702 ( .A(n41059), .B(n41060), .Z(n41055) );
  AND U40703 ( .A(n41061), .B(n41062), .Z(n41060) );
  XOR U40704 ( .A(n40988), .B(n41059), .Z(n41062) );
  XOR U40705 ( .A(n41059), .B(n40989), .Z(n41061) );
  XOR U40706 ( .A(n41063), .B(n41064), .Z(n41059) );
  AND U40707 ( .A(n41065), .B(n41066), .Z(n41064) );
  XOR U40708 ( .A(n41063), .B(n41037), .Z(n41066) );
  XNOR U40709 ( .A(n41067), .B(n41068), .Z(n40891) );
  AND U40710 ( .A(n1086), .B(n41069), .Z(n41068) );
  XNOR U40711 ( .A(n41070), .B(n41071), .Z(n1086) );
  AND U40712 ( .A(n41072), .B(n41073), .Z(n41071) );
  XOR U40713 ( .A(n41070), .B(n40901), .Z(n41073) );
  XNOR U40714 ( .A(n41070), .B(n40861), .Z(n41072) );
  XOR U40715 ( .A(n41074), .B(n41075), .Z(n41070) );
  AND U40716 ( .A(n41076), .B(n41077), .Z(n41075) );
  XOR U40717 ( .A(n41074), .B(n40869), .Z(n41076) );
  XOR U40718 ( .A(n41078), .B(n41079), .Z(n40852) );
  AND U40719 ( .A(n1090), .B(n41069), .Z(n41079) );
  XNOR U40720 ( .A(n41067), .B(n41078), .Z(n41069) );
  XNOR U40721 ( .A(n41080), .B(n41081), .Z(n1090) );
  AND U40722 ( .A(n41082), .B(n41083), .Z(n41081) );
  XNOR U40723 ( .A(n41084), .B(n41080), .Z(n41083) );
  IV U40724 ( .A(n40901), .Z(n41084) );
  XOR U40725 ( .A(n41054), .B(n41085), .Z(n40901) );
  AND U40726 ( .A(n1093), .B(n41086), .Z(n41085) );
  XOR U40727 ( .A(n40944), .B(n40941), .Z(n41086) );
  IV U40728 ( .A(n41054), .Z(n40944) );
  XNOR U40729 ( .A(n40861), .B(n41080), .Z(n41082) );
  XOR U40730 ( .A(n41087), .B(n41088), .Z(n40861) );
  AND U40731 ( .A(n1109), .B(n41089), .Z(n41088) );
  XOR U40732 ( .A(n41074), .B(n41090), .Z(n41080) );
  AND U40733 ( .A(n41091), .B(n41077), .Z(n41090) );
  XNOR U40734 ( .A(n40911), .B(n41074), .Z(n41077) );
  XOR U40735 ( .A(n40961), .B(n41092), .Z(n40911) );
  AND U40736 ( .A(n1093), .B(n41093), .Z(n41092) );
  XOR U40737 ( .A(n40957), .B(n40961), .Z(n41093) );
  XNOR U40738 ( .A(n41094), .B(n41074), .Z(n41091) );
  IV U40739 ( .A(n40869), .Z(n41094) );
  XOR U40740 ( .A(n41095), .B(n41096), .Z(n40869) );
  AND U40741 ( .A(n1109), .B(n41097), .Z(n41096) );
  XOR U40742 ( .A(n41098), .B(n41099), .Z(n41074) );
  AND U40743 ( .A(n41100), .B(n41101), .Z(n41099) );
  XNOR U40744 ( .A(n40921), .B(n41098), .Z(n41101) );
  XOR U40745 ( .A(n40989), .B(n41102), .Z(n40921) );
  AND U40746 ( .A(n1093), .B(n41103), .Z(n41102) );
  XOR U40747 ( .A(n40985), .B(n40989), .Z(n41103) );
  XOR U40748 ( .A(n41098), .B(n40878), .Z(n41100) );
  XOR U40749 ( .A(n41104), .B(n41105), .Z(n40878) );
  AND U40750 ( .A(n1109), .B(n41106), .Z(n41105) );
  XOR U40751 ( .A(n41107), .B(n41108), .Z(n41098) );
  AND U40752 ( .A(n41109), .B(n41110), .Z(n41108) );
  XNOR U40753 ( .A(n41107), .B(n40929), .Z(n41110) );
  XOR U40754 ( .A(n41038), .B(n41111), .Z(n40929) );
  AND U40755 ( .A(n1093), .B(n41112), .Z(n41111) );
  XOR U40756 ( .A(n41034), .B(n41038), .Z(n41112) );
  XNOR U40757 ( .A(n41113), .B(n41107), .Z(n41109) );
  IV U40758 ( .A(n40888), .Z(n41113) );
  XOR U40759 ( .A(n41114), .B(n41115), .Z(n40888) );
  AND U40760 ( .A(n1109), .B(n41116), .Z(n41115) );
  AND U40761 ( .A(n41078), .B(n41067), .Z(n41107) );
  XNOR U40762 ( .A(n41117), .B(n41118), .Z(n41067) );
  AND U40763 ( .A(n1093), .B(n41049), .Z(n41118) );
  XNOR U40764 ( .A(n41047), .B(n41117), .Z(n41049) );
  XNOR U40765 ( .A(n41119), .B(n41120), .Z(n1093) );
  AND U40766 ( .A(n41121), .B(n41122), .Z(n41120) );
  XNOR U40767 ( .A(n41119), .B(n40941), .Z(n41122) );
  IV U40768 ( .A(n40945), .Z(n40941) );
  XOR U40769 ( .A(n41123), .B(n41124), .Z(n40945) );
  AND U40770 ( .A(n1097), .B(n41125), .Z(n41124) );
  XOR U40771 ( .A(n41126), .B(n41123), .Z(n41125) );
  XNOR U40772 ( .A(n41119), .B(n41054), .Z(n41121) );
  XOR U40773 ( .A(n41127), .B(n41128), .Z(n41054) );
  AND U40774 ( .A(n1105), .B(n41089), .Z(n41128) );
  XOR U40775 ( .A(n41087), .B(n41127), .Z(n41089) );
  XOR U40776 ( .A(n41129), .B(n41130), .Z(n41119) );
  AND U40777 ( .A(n41131), .B(n41132), .Z(n41130) );
  XNOR U40778 ( .A(n41129), .B(n40957), .Z(n41132) );
  IV U40779 ( .A(n40960), .Z(n40957) );
  XOR U40780 ( .A(n41133), .B(n41134), .Z(n40960) );
  AND U40781 ( .A(n1097), .B(n41135), .Z(n41134) );
  XOR U40782 ( .A(n41136), .B(n41133), .Z(n41135) );
  XOR U40783 ( .A(n40961), .B(n41129), .Z(n41131) );
  XOR U40784 ( .A(n41137), .B(n41138), .Z(n40961) );
  AND U40785 ( .A(n1105), .B(n41097), .Z(n41138) );
  XOR U40786 ( .A(n41137), .B(n41095), .Z(n41097) );
  XOR U40787 ( .A(n41139), .B(n41140), .Z(n41129) );
  AND U40788 ( .A(n41141), .B(n41142), .Z(n41140) );
  XNOR U40789 ( .A(n41139), .B(n40985), .Z(n41142) );
  IV U40790 ( .A(n40988), .Z(n40985) );
  XOR U40791 ( .A(n41143), .B(n41144), .Z(n40988) );
  AND U40792 ( .A(n1097), .B(n41145), .Z(n41144) );
  XNOR U40793 ( .A(n41146), .B(n41143), .Z(n41145) );
  XOR U40794 ( .A(n40989), .B(n41139), .Z(n41141) );
  XOR U40795 ( .A(n41147), .B(n41148), .Z(n40989) );
  AND U40796 ( .A(n1105), .B(n41106), .Z(n41148) );
  XOR U40797 ( .A(n41147), .B(n41104), .Z(n41106) );
  XOR U40798 ( .A(n41063), .B(n41149), .Z(n41139) );
  AND U40799 ( .A(n41065), .B(n41150), .Z(n41149) );
  XNOR U40800 ( .A(n41063), .B(n41034), .Z(n41150) );
  IV U40801 ( .A(n41037), .Z(n41034) );
  XOR U40802 ( .A(n41151), .B(n41152), .Z(n41037) );
  AND U40803 ( .A(n1097), .B(n41153), .Z(n41152) );
  XOR U40804 ( .A(n41154), .B(n41151), .Z(n41153) );
  XOR U40805 ( .A(n41038), .B(n41063), .Z(n41065) );
  XOR U40806 ( .A(n41155), .B(n41156), .Z(n41038) );
  AND U40807 ( .A(n1105), .B(n41116), .Z(n41156) );
  XOR U40808 ( .A(n41155), .B(n41114), .Z(n41116) );
  AND U40809 ( .A(n41117), .B(n41047), .Z(n41063) );
  XNOR U40810 ( .A(n41157), .B(n41158), .Z(n41047) );
  AND U40811 ( .A(n1097), .B(n41159), .Z(n41158) );
  XNOR U40812 ( .A(n41160), .B(n41157), .Z(n41159) );
  XNOR U40813 ( .A(n41161), .B(n41162), .Z(n1097) );
  AND U40814 ( .A(n41163), .B(n41164), .Z(n41162) );
  XOR U40815 ( .A(n41126), .B(n41161), .Z(n41164) );
  AND U40816 ( .A(n41165), .B(n41166), .Z(n41126) );
  XNOR U40817 ( .A(n41123), .B(n41161), .Z(n41163) );
  XNOR U40818 ( .A(n41167), .B(n41168), .Z(n41123) );
  AND U40819 ( .A(n1101), .B(n41169), .Z(n41168) );
  XNOR U40820 ( .A(n41170), .B(n41171), .Z(n41169) );
  XOR U40821 ( .A(n41172), .B(n41173), .Z(n41161) );
  AND U40822 ( .A(n41174), .B(n41175), .Z(n41173) );
  XNOR U40823 ( .A(n41172), .B(n41165), .Z(n41175) );
  IV U40824 ( .A(n41136), .Z(n41165) );
  XOR U40825 ( .A(n41176), .B(n41177), .Z(n41136) );
  XOR U40826 ( .A(n41178), .B(n41166), .Z(n41177) );
  AND U40827 ( .A(n41146), .B(n41179), .Z(n41166) );
  AND U40828 ( .A(n41180), .B(n41181), .Z(n41178) );
  XOR U40829 ( .A(n41182), .B(n41176), .Z(n41180) );
  XNOR U40830 ( .A(n41133), .B(n41172), .Z(n41174) );
  XNOR U40831 ( .A(n41183), .B(n41184), .Z(n41133) );
  AND U40832 ( .A(n1101), .B(n41185), .Z(n41184) );
  XNOR U40833 ( .A(n41186), .B(n41187), .Z(n41185) );
  XOR U40834 ( .A(n41188), .B(n41189), .Z(n41172) );
  AND U40835 ( .A(n41190), .B(n41191), .Z(n41189) );
  XNOR U40836 ( .A(n41188), .B(n41146), .Z(n41191) );
  XOR U40837 ( .A(n41192), .B(n41181), .Z(n41146) );
  XNOR U40838 ( .A(n41193), .B(n41176), .Z(n41181) );
  XOR U40839 ( .A(n41194), .B(n41195), .Z(n41176) );
  AND U40840 ( .A(n41196), .B(n41197), .Z(n41195) );
  XOR U40841 ( .A(n41198), .B(n41194), .Z(n41196) );
  XNOR U40842 ( .A(n41199), .B(n41200), .Z(n41193) );
  AND U40843 ( .A(n41201), .B(n41202), .Z(n41200) );
  XOR U40844 ( .A(n41199), .B(n41203), .Z(n41201) );
  XNOR U40845 ( .A(n41182), .B(n41179), .Z(n41192) );
  AND U40846 ( .A(n41204), .B(n41205), .Z(n41179) );
  XOR U40847 ( .A(n41206), .B(n41207), .Z(n41182) );
  AND U40848 ( .A(n41208), .B(n41209), .Z(n41207) );
  XOR U40849 ( .A(n41206), .B(n41210), .Z(n41208) );
  XNOR U40850 ( .A(n41143), .B(n41188), .Z(n41190) );
  XNOR U40851 ( .A(n41211), .B(n41212), .Z(n41143) );
  AND U40852 ( .A(n1101), .B(n41213), .Z(n41212) );
  XNOR U40853 ( .A(n41214), .B(n41215), .Z(n41213) );
  XOR U40854 ( .A(n41216), .B(n41217), .Z(n41188) );
  AND U40855 ( .A(n41218), .B(n41219), .Z(n41217) );
  XNOR U40856 ( .A(n41216), .B(n41204), .Z(n41219) );
  IV U40857 ( .A(n41154), .Z(n41204) );
  XNOR U40858 ( .A(n41220), .B(n41197), .Z(n41154) );
  XNOR U40859 ( .A(n41221), .B(n41203), .Z(n41197) );
  XOR U40860 ( .A(n41222), .B(n41223), .Z(n41203) );
  NOR U40861 ( .A(n41224), .B(n41225), .Z(n41223) );
  XNOR U40862 ( .A(n41222), .B(n41226), .Z(n41224) );
  XNOR U40863 ( .A(n41202), .B(n41194), .Z(n41221) );
  XOR U40864 ( .A(n41227), .B(n41228), .Z(n41194) );
  AND U40865 ( .A(n41229), .B(n41230), .Z(n41228) );
  XNOR U40866 ( .A(n41227), .B(n41231), .Z(n41229) );
  XNOR U40867 ( .A(n41232), .B(n41199), .Z(n41202) );
  XOR U40868 ( .A(n41233), .B(n41234), .Z(n41199) );
  AND U40869 ( .A(n41235), .B(n41236), .Z(n41234) );
  XOR U40870 ( .A(n41233), .B(n41237), .Z(n41235) );
  XNOR U40871 ( .A(n41238), .B(n41239), .Z(n41232) );
  NOR U40872 ( .A(n41240), .B(n41241), .Z(n41239) );
  XOR U40873 ( .A(n41238), .B(n41242), .Z(n41240) );
  XNOR U40874 ( .A(n41198), .B(n41205), .Z(n41220) );
  NOR U40875 ( .A(n41160), .B(n41243), .Z(n41205) );
  XOR U40876 ( .A(n41210), .B(n41209), .Z(n41198) );
  XNOR U40877 ( .A(n41244), .B(n41206), .Z(n41209) );
  XOR U40878 ( .A(n41245), .B(n41246), .Z(n41206) );
  AND U40879 ( .A(n41247), .B(n41248), .Z(n41246) );
  XOR U40880 ( .A(n41245), .B(n41249), .Z(n41247) );
  XNOR U40881 ( .A(n41250), .B(n41251), .Z(n41244) );
  NOR U40882 ( .A(n41252), .B(n41253), .Z(n41251) );
  XNOR U40883 ( .A(n41250), .B(n41254), .Z(n41252) );
  XOR U40884 ( .A(n41255), .B(n41256), .Z(n41210) );
  NOR U40885 ( .A(n41257), .B(n41258), .Z(n41256) );
  XNOR U40886 ( .A(n41255), .B(n41259), .Z(n41257) );
  XNOR U40887 ( .A(n41151), .B(n41216), .Z(n41218) );
  XNOR U40888 ( .A(n41260), .B(n41261), .Z(n41151) );
  AND U40889 ( .A(n1101), .B(n41262), .Z(n41261) );
  XNOR U40890 ( .A(n41263), .B(n41264), .Z(n41262) );
  AND U40891 ( .A(n41157), .B(n41160), .Z(n41216) );
  XOR U40892 ( .A(n41265), .B(n41243), .Z(n41160) );
  XNOR U40893 ( .A(p_input[2048]), .B(p_input[864]), .Z(n41243) );
  XOR U40894 ( .A(n41231), .B(n41230), .Z(n41265) );
  XNOR U40895 ( .A(n41266), .B(n41237), .Z(n41230) );
  XNOR U40896 ( .A(n41226), .B(n41225), .Z(n41237) );
  XOR U40897 ( .A(n41267), .B(n41222), .Z(n41225) );
  XNOR U40898 ( .A(n29266), .B(p_input[874]), .Z(n41222) );
  XNOR U40899 ( .A(p_input[2059]), .B(p_input[875]), .Z(n41267) );
  XOR U40900 ( .A(p_input[2060]), .B(p_input[876]), .Z(n41226) );
  XNOR U40901 ( .A(n41236), .B(n41227), .Z(n41266) );
  XNOR U40902 ( .A(n29494), .B(p_input[865]), .Z(n41227) );
  XOR U40903 ( .A(n41268), .B(n41242), .Z(n41236) );
  XNOR U40904 ( .A(p_input[2063]), .B(p_input[879]), .Z(n41242) );
  XOR U40905 ( .A(n41233), .B(n41241), .Z(n41268) );
  XOR U40906 ( .A(n41269), .B(n41238), .Z(n41241) );
  XOR U40907 ( .A(p_input[2061]), .B(p_input[877]), .Z(n41238) );
  XNOR U40908 ( .A(p_input[2062]), .B(p_input[878]), .Z(n41269) );
  XNOR U40909 ( .A(n29036), .B(p_input[873]), .Z(n41233) );
  XNOR U40910 ( .A(n41249), .B(n41248), .Z(n41231) );
  XNOR U40911 ( .A(n41270), .B(n41254), .Z(n41248) );
  XOR U40912 ( .A(p_input[2056]), .B(p_input[872]), .Z(n41254) );
  XOR U40913 ( .A(n41245), .B(n41253), .Z(n41270) );
  XOR U40914 ( .A(n41271), .B(n41250), .Z(n41253) );
  XOR U40915 ( .A(p_input[2054]), .B(p_input[870]), .Z(n41250) );
  XNOR U40916 ( .A(p_input[2055]), .B(p_input[871]), .Z(n41271) );
  XNOR U40917 ( .A(n29039), .B(p_input[866]), .Z(n41245) );
  XNOR U40918 ( .A(n41259), .B(n41258), .Z(n41249) );
  XOR U40919 ( .A(n41272), .B(n41255), .Z(n41258) );
  XOR U40920 ( .A(p_input[2051]), .B(p_input[867]), .Z(n41255) );
  XNOR U40921 ( .A(p_input[2052]), .B(p_input[868]), .Z(n41272) );
  XOR U40922 ( .A(p_input[2053]), .B(p_input[869]), .Z(n41259) );
  XNOR U40923 ( .A(n41273), .B(n41274), .Z(n41157) );
  AND U40924 ( .A(n1101), .B(n41275), .Z(n41274) );
  XNOR U40925 ( .A(n41276), .B(n41277), .Z(n1101) );
  AND U40926 ( .A(n41278), .B(n41279), .Z(n41277) );
  XOR U40927 ( .A(n41171), .B(n41276), .Z(n41279) );
  XNOR U40928 ( .A(n41280), .B(n41276), .Z(n41278) );
  XOR U40929 ( .A(n41281), .B(n41282), .Z(n41276) );
  AND U40930 ( .A(n41283), .B(n41284), .Z(n41282) );
  XOR U40931 ( .A(n41186), .B(n41281), .Z(n41284) );
  XOR U40932 ( .A(n41281), .B(n41187), .Z(n41283) );
  XOR U40933 ( .A(n41285), .B(n41286), .Z(n41281) );
  AND U40934 ( .A(n41287), .B(n41288), .Z(n41286) );
  XOR U40935 ( .A(n41214), .B(n41285), .Z(n41288) );
  XOR U40936 ( .A(n41285), .B(n41215), .Z(n41287) );
  XOR U40937 ( .A(n41289), .B(n41290), .Z(n41285) );
  AND U40938 ( .A(n41291), .B(n41292), .Z(n41290) );
  XOR U40939 ( .A(n41289), .B(n41263), .Z(n41292) );
  XNOR U40940 ( .A(n41293), .B(n41294), .Z(n41117) );
  AND U40941 ( .A(n1105), .B(n41295), .Z(n41294) );
  XNOR U40942 ( .A(n41296), .B(n41297), .Z(n1105) );
  AND U40943 ( .A(n41298), .B(n41299), .Z(n41297) );
  XOR U40944 ( .A(n41296), .B(n41127), .Z(n41299) );
  XNOR U40945 ( .A(n41296), .B(n41087), .Z(n41298) );
  XOR U40946 ( .A(n41300), .B(n41301), .Z(n41296) );
  AND U40947 ( .A(n41302), .B(n41303), .Z(n41301) );
  XOR U40948 ( .A(n41300), .B(n41095), .Z(n41302) );
  XOR U40949 ( .A(n41304), .B(n41305), .Z(n41078) );
  AND U40950 ( .A(n1109), .B(n41295), .Z(n41305) );
  XNOR U40951 ( .A(n41293), .B(n41304), .Z(n41295) );
  XNOR U40952 ( .A(n41306), .B(n41307), .Z(n1109) );
  AND U40953 ( .A(n41308), .B(n41309), .Z(n41307) );
  XNOR U40954 ( .A(n41310), .B(n41306), .Z(n41309) );
  IV U40955 ( .A(n41127), .Z(n41310) );
  XOR U40956 ( .A(n41280), .B(n41311), .Z(n41127) );
  AND U40957 ( .A(n1112), .B(n41312), .Z(n41311) );
  XOR U40958 ( .A(n41170), .B(n41167), .Z(n41312) );
  IV U40959 ( .A(n41280), .Z(n41170) );
  XNOR U40960 ( .A(n41087), .B(n41306), .Z(n41308) );
  XOR U40961 ( .A(n41313), .B(n41314), .Z(n41087) );
  AND U40962 ( .A(n1128), .B(n41315), .Z(n41314) );
  XOR U40963 ( .A(n41300), .B(n41316), .Z(n41306) );
  AND U40964 ( .A(n41317), .B(n41303), .Z(n41316) );
  XNOR U40965 ( .A(n41137), .B(n41300), .Z(n41303) );
  XOR U40966 ( .A(n41187), .B(n41318), .Z(n41137) );
  AND U40967 ( .A(n1112), .B(n41319), .Z(n41318) );
  XOR U40968 ( .A(n41183), .B(n41187), .Z(n41319) );
  XNOR U40969 ( .A(n41320), .B(n41300), .Z(n41317) );
  IV U40970 ( .A(n41095), .Z(n41320) );
  XOR U40971 ( .A(n41321), .B(n41322), .Z(n41095) );
  AND U40972 ( .A(n1128), .B(n41323), .Z(n41322) );
  XOR U40973 ( .A(n41324), .B(n41325), .Z(n41300) );
  AND U40974 ( .A(n41326), .B(n41327), .Z(n41325) );
  XNOR U40975 ( .A(n41147), .B(n41324), .Z(n41327) );
  XOR U40976 ( .A(n41215), .B(n41328), .Z(n41147) );
  AND U40977 ( .A(n1112), .B(n41329), .Z(n41328) );
  XOR U40978 ( .A(n41211), .B(n41215), .Z(n41329) );
  XOR U40979 ( .A(n41324), .B(n41104), .Z(n41326) );
  XOR U40980 ( .A(n41330), .B(n41331), .Z(n41104) );
  AND U40981 ( .A(n1128), .B(n41332), .Z(n41331) );
  XOR U40982 ( .A(n41333), .B(n41334), .Z(n41324) );
  AND U40983 ( .A(n41335), .B(n41336), .Z(n41334) );
  XNOR U40984 ( .A(n41333), .B(n41155), .Z(n41336) );
  XOR U40985 ( .A(n41264), .B(n41337), .Z(n41155) );
  AND U40986 ( .A(n1112), .B(n41338), .Z(n41337) );
  XOR U40987 ( .A(n41260), .B(n41264), .Z(n41338) );
  XNOR U40988 ( .A(n41339), .B(n41333), .Z(n41335) );
  IV U40989 ( .A(n41114), .Z(n41339) );
  XOR U40990 ( .A(n41340), .B(n41341), .Z(n41114) );
  AND U40991 ( .A(n1128), .B(n41342), .Z(n41341) );
  AND U40992 ( .A(n41304), .B(n41293), .Z(n41333) );
  XNOR U40993 ( .A(n41343), .B(n41344), .Z(n41293) );
  AND U40994 ( .A(n1112), .B(n41275), .Z(n41344) );
  XNOR U40995 ( .A(n41273), .B(n41343), .Z(n41275) );
  XNOR U40996 ( .A(n41345), .B(n41346), .Z(n1112) );
  AND U40997 ( .A(n41347), .B(n41348), .Z(n41346) );
  XNOR U40998 ( .A(n41345), .B(n41167), .Z(n41348) );
  IV U40999 ( .A(n41171), .Z(n41167) );
  XOR U41000 ( .A(n41349), .B(n41350), .Z(n41171) );
  AND U41001 ( .A(n1116), .B(n41351), .Z(n41350) );
  XOR U41002 ( .A(n41352), .B(n41349), .Z(n41351) );
  XNOR U41003 ( .A(n41345), .B(n41280), .Z(n41347) );
  XOR U41004 ( .A(n41353), .B(n41354), .Z(n41280) );
  AND U41005 ( .A(n1124), .B(n41315), .Z(n41354) );
  XOR U41006 ( .A(n41313), .B(n41353), .Z(n41315) );
  XOR U41007 ( .A(n41355), .B(n41356), .Z(n41345) );
  AND U41008 ( .A(n41357), .B(n41358), .Z(n41356) );
  XNOR U41009 ( .A(n41355), .B(n41183), .Z(n41358) );
  IV U41010 ( .A(n41186), .Z(n41183) );
  XOR U41011 ( .A(n41359), .B(n41360), .Z(n41186) );
  AND U41012 ( .A(n1116), .B(n41361), .Z(n41360) );
  XOR U41013 ( .A(n41362), .B(n41359), .Z(n41361) );
  XOR U41014 ( .A(n41187), .B(n41355), .Z(n41357) );
  XOR U41015 ( .A(n41363), .B(n41364), .Z(n41187) );
  AND U41016 ( .A(n1124), .B(n41323), .Z(n41364) );
  XOR U41017 ( .A(n41363), .B(n41321), .Z(n41323) );
  XOR U41018 ( .A(n41365), .B(n41366), .Z(n41355) );
  AND U41019 ( .A(n41367), .B(n41368), .Z(n41366) );
  XNOR U41020 ( .A(n41365), .B(n41211), .Z(n41368) );
  IV U41021 ( .A(n41214), .Z(n41211) );
  XOR U41022 ( .A(n41369), .B(n41370), .Z(n41214) );
  AND U41023 ( .A(n1116), .B(n41371), .Z(n41370) );
  XNOR U41024 ( .A(n41372), .B(n41369), .Z(n41371) );
  XOR U41025 ( .A(n41215), .B(n41365), .Z(n41367) );
  XOR U41026 ( .A(n41373), .B(n41374), .Z(n41215) );
  AND U41027 ( .A(n1124), .B(n41332), .Z(n41374) );
  XOR U41028 ( .A(n41373), .B(n41330), .Z(n41332) );
  XOR U41029 ( .A(n41289), .B(n41375), .Z(n41365) );
  AND U41030 ( .A(n41291), .B(n41376), .Z(n41375) );
  XNOR U41031 ( .A(n41289), .B(n41260), .Z(n41376) );
  IV U41032 ( .A(n41263), .Z(n41260) );
  XOR U41033 ( .A(n41377), .B(n41378), .Z(n41263) );
  AND U41034 ( .A(n1116), .B(n41379), .Z(n41378) );
  XOR U41035 ( .A(n41380), .B(n41377), .Z(n41379) );
  XOR U41036 ( .A(n41264), .B(n41289), .Z(n41291) );
  XOR U41037 ( .A(n41381), .B(n41382), .Z(n41264) );
  AND U41038 ( .A(n1124), .B(n41342), .Z(n41382) );
  XOR U41039 ( .A(n41381), .B(n41340), .Z(n41342) );
  AND U41040 ( .A(n41343), .B(n41273), .Z(n41289) );
  XNOR U41041 ( .A(n41383), .B(n41384), .Z(n41273) );
  AND U41042 ( .A(n1116), .B(n41385), .Z(n41384) );
  XNOR U41043 ( .A(n41386), .B(n41383), .Z(n41385) );
  XNOR U41044 ( .A(n41387), .B(n41388), .Z(n1116) );
  AND U41045 ( .A(n41389), .B(n41390), .Z(n41388) );
  XOR U41046 ( .A(n41352), .B(n41387), .Z(n41390) );
  AND U41047 ( .A(n41391), .B(n41392), .Z(n41352) );
  XNOR U41048 ( .A(n41349), .B(n41387), .Z(n41389) );
  XNOR U41049 ( .A(n41393), .B(n41394), .Z(n41349) );
  AND U41050 ( .A(n1120), .B(n41395), .Z(n41394) );
  XNOR U41051 ( .A(n41396), .B(n41397), .Z(n41395) );
  XOR U41052 ( .A(n41398), .B(n41399), .Z(n41387) );
  AND U41053 ( .A(n41400), .B(n41401), .Z(n41399) );
  XNOR U41054 ( .A(n41398), .B(n41391), .Z(n41401) );
  IV U41055 ( .A(n41362), .Z(n41391) );
  XOR U41056 ( .A(n41402), .B(n41403), .Z(n41362) );
  XOR U41057 ( .A(n41404), .B(n41392), .Z(n41403) );
  AND U41058 ( .A(n41372), .B(n41405), .Z(n41392) );
  AND U41059 ( .A(n41406), .B(n41407), .Z(n41404) );
  XOR U41060 ( .A(n41408), .B(n41402), .Z(n41406) );
  XNOR U41061 ( .A(n41359), .B(n41398), .Z(n41400) );
  XNOR U41062 ( .A(n41409), .B(n41410), .Z(n41359) );
  AND U41063 ( .A(n1120), .B(n41411), .Z(n41410) );
  XNOR U41064 ( .A(n41412), .B(n41413), .Z(n41411) );
  XOR U41065 ( .A(n41414), .B(n41415), .Z(n41398) );
  AND U41066 ( .A(n41416), .B(n41417), .Z(n41415) );
  XNOR U41067 ( .A(n41414), .B(n41372), .Z(n41417) );
  XOR U41068 ( .A(n41418), .B(n41407), .Z(n41372) );
  XNOR U41069 ( .A(n41419), .B(n41402), .Z(n41407) );
  XOR U41070 ( .A(n41420), .B(n41421), .Z(n41402) );
  AND U41071 ( .A(n41422), .B(n41423), .Z(n41421) );
  XOR U41072 ( .A(n41424), .B(n41420), .Z(n41422) );
  XNOR U41073 ( .A(n41425), .B(n41426), .Z(n41419) );
  AND U41074 ( .A(n41427), .B(n41428), .Z(n41426) );
  XOR U41075 ( .A(n41425), .B(n41429), .Z(n41427) );
  XNOR U41076 ( .A(n41408), .B(n41405), .Z(n41418) );
  AND U41077 ( .A(n41430), .B(n41431), .Z(n41405) );
  XOR U41078 ( .A(n41432), .B(n41433), .Z(n41408) );
  AND U41079 ( .A(n41434), .B(n41435), .Z(n41433) );
  XOR U41080 ( .A(n41432), .B(n41436), .Z(n41434) );
  XNOR U41081 ( .A(n41369), .B(n41414), .Z(n41416) );
  XNOR U41082 ( .A(n41437), .B(n41438), .Z(n41369) );
  AND U41083 ( .A(n1120), .B(n41439), .Z(n41438) );
  XNOR U41084 ( .A(n41440), .B(n41441), .Z(n41439) );
  XOR U41085 ( .A(n41442), .B(n41443), .Z(n41414) );
  AND U41086 ( .A(n41444), .B(n41445), .Z(n41443) );
  XNOR U41087 ( .A(n41442), .B(n41430), .Z(n41445) );
  IV U41088 ( .A(n41380), .Z(n41430) );
  XNOR U41089 ( .A(n41446), .B(n41423), .Z(n41380) );
  XNOR U41090 ( .A(n41447), .B(n41429), .Z(n41423) );
  XOR U41091 ( .A(n41448), .B(n41449), .Z(n41429) );
  NOR U41092 ( .A(n41450), .B(n41451), .Z(n41449) );
  XNOR U41093 ( .A(n41448), .B(n41452), .Z(n41450) );
  XNOR U41094 ( .A(n41428), .B(n41420), .Z(n41447) );
  XOR U41095 ( .A(n41453), .B(n41454), .Z(n41420) );
  AND U41096 ( .A(n41455), .B(n41456), .Z(n41454) );
  XNOR U41097 ( .A(n41453), .B(n41457), .Z(n41455) );
  XNOR U41098 ( .A(n41458), .B(n41425), .Z(n41428) );
  XOR U41099 ( .A(n41459), .B(n41460), .Z(n41425) );
  AND U41100 ( .A(n41461), .B(n41462), .Z(n41460) );
  XOR U41101 ( .A(n41459), .B(n41463), .Z(n41461) );
  XNOR U41102 ( .A(n41464), .B(n41465), .Z(n41458) );
  NOR U41103 ( .A(n41466), .B(n41467), .Z(n41465) );
  XOR U41104 ( .A(n41464), .B(n41468), .Z(n41466) );
  XNOR U41105 ( .A(n41424), .B(n41431), .Z(n41446) );
  NOR U41106 ( .A(n41386), .B(n41469), .Z(n41431) );
  XOR U41107 ( .A(n41436), .B(n41435), .Z(n41424) );
  XNOR U41108 ( .A(n41470), .B(n41432), .Z(n41435) );
  XOR U41109 ( .A(n41471), .B(n41472), .Z(n41432) );
  AND U41110 ( .A(n41473), .B(n41474), .Z(n41472) );
  XOR U41111 ( .A(n41471), .B(n41475), .Z(n41473) );
  XNOR U41112 ( .A(n41476), .B(n41477), .Z(n41470) );
  NOR U41113 ( .A(n41478), .B(n41479), .Z(n41477) );
  XNOR U41114 ( .A(n41476), .B(n41480), .Z(n41478) );
  XOR U41115 ( .A(n41481), .B(n41482), .Z(n41436) );
  NOR U41116 ( .A(n41483), .B(n41484), .Z(n41482) );
  XNOR U41117 ( .A(n41481), .B(n41485), .Z(n41483) );
  XNOR U41118 ( .A(n41377), .B(n41442), .Z(n41444) );
  XNOR U41119 ( .A(n41486), .B(n41487), .Z(n41377) );
  AND U41120 ( .A(n1120), .B(n41488), .Z(n41487) );
  XNOR U41121 ( .A(n41489), .B(n41490), .Z(n41488) );
  AND U41122 ( .A(n41383), .B(n41386), .Z(n41442) );
  XOR U41123 ( .A(n41491), .B(n41469), .Z(n41386) );
  XNOR U41124 ( .A(p_input[2048]), .B(p_input[880]), .Z(n41469) );
  XOR U41125 ( .A(n41457), .B(n41456), .Z(n41491) );
  XNOR U41126 ( .A(n41492), .B(n41463), .Z(n41456) );
  XNOR U41127 ( .A(n41452), .B(n41451), .Z(n41463) );
  XOR U41128 ( .A(n41493), .B(n41448), .Z(n41451) );
  XNOR U41129 ( .A(n29266), .B(p_input[890]), .Z(n41448) );
  XNOR U41130 ( .A(p_input[2059]), .B(p_input[891]), .Z(n41493) );
  XOR U41131 ( .A(p_input[2060]), .B(p_input[892]), .Z(n41452) );
  XNOR U41132 ( .A(n41462), .B(n41453), .Z(n41492) );
  XNOR U41133 ( .A(n29494), .B(p_input[881]), .Z(n41453) );
  XOR U41134 ( .A(n41494), .B(n41468), .Z(n41462) );
  XNOR U41135 ( .A(p_input[2063]), .B(p_input[895]), .Z(n41468) );
  XOR U41136 ( .A(n41459), .B(n41467), .Z(n41494) );
  XOR U41137 ( .A(n41495), .B(n41464), .Z(n41467) );
  XOR U41138 ( .A(p_input[2061]), .B(p_input[893]), .Z(n41464) );
  XNOR U41139 ( .A(p_input[2062]), .B(p_input[894]), .Z(n41495) );
  XNOR U41140 ( .A(n29036), .B(p_input[889]), .Z(n41459) );
  XNOR U41141 ( .A(n41475), .B(n41474), .Z(n41457) );
  XNOR U41142 ( .A(n41496), .B(n41480), .Z(n41474) );
  XOR U41143 ( .A(p_input[2056]), .B(p_input[888]), .Z(n41480) );
  XOR U41144 ( .A(n41471), .B(n41479), .Z(n41496) );
  XOR U41145 ( .A(n41497), .B(n41476), .Z(n41479) );
  XOR U41146 ( .A(p_input[2054]), .B(p_input[886]), .Z(n41476) );
  XNOR U41147 ( .A(p_input[2055]), .B(p_input[887]), .Z(n41497) );
  XNOR U41148 ( .A(n29039), .B(p_input[882]), .Z(n41471) );
  XNOR U41149 ( .A(n41485), .B(n41484), .Z(n41475) );
  XOR U41150 ( .A(n41498), .B(n41481), .Z(n41484) );
  XOR U41151 ( .A(p_input[2051]), .B(p_input[883]), .Z(n41481) );
  XNOR U41152 ( .A(p_input[2052]), .B(p_input[884]), .Z(n41498) );
  XOR U41153 ( .A(p_input[2053]), .B(p_input[885]), .Z(n41485) );
  XNOR U41154 ( .A(n41499), .B(n41500), .Z(n41383) );
  AND U41155 ( .A(n1120), .B(n41501), .Z(n41500) );
  XNOR U41156 ( .A(n41502), .B(n41503), .Z(n1120) );
  AND U41157 ( .A(n41504), .B(n41505), .Z(n41503) );
  XOR U41158 ( .A(n41397), .B(n41502), .Z(n41505) );
  XNOR U41159 ( .A(n41506), .B(n41502), .Z(n41504) );
  XOR U41160 ( .A(n41507), .B(n41508), .Z(n41502) );
  AND U41161 ( .A(n41509), .B(n41510), .Z(n41508) );
  XOR U41162 ( .A(n41412), .B(n41507), .Z(n41510) );
  XOR U41163 ( .A(n41507), .B(n41413), .Z(n41509) );
  XOR U41164 ( .A(n41511), .B(n41512), .Z(n41507) );
  AND U41165 ( .A(n41513), .B(n41514), .Z(n41512) );
  XOR U41166 ( .A(n41440), .B(n41511), .Z(n41514) );
  XOR U41167 ( .A(n41511), .B(n41441), .Z(n41513) );
  XOR U41168 ( .A(n41515), .B(n41516), .Z(n41511) );
  AND U41169 ( .A(n41517), .B(n41518), .Z(n41516) );
  XOR U41170 ( .A(n41515), .B(n41489), .Z(n41518) );
  XNOR U41171 ( .A(n41519), .B(n41520), .Z(n41343) );
  AND U41172 ( .A(n1124), .B(n41521), .Z(n41520) );
  XNOR U41173 ( .A(n41522), .B(n41523), .Z(n1124) );
  AND U41174 ( .A(n41524), .B(n41525), .Z(n41523) );
  XOR U41175 ( .A(n41522), .B(n41353), .Z(n41525) );
  XNOR U41176 ( .A(n41522), .B(n41313), .Z(n41524) );
  XOR U41177 ( .A(n41526), .B(n41527), .Z(n41522) );
  AND U41178 ( .A(n41528), .B(n41529), .Z(n41527) );
  XOR U41179 ( .A(n41526), .B(n41321), .Z(n41528) );
  XOR U41180 ( .A(n41530), .B(n41531), .Z(n41304) );
  AND U41181 ( .A(n1128), .B(n41521), .Z(n41531) );
  XNOR U41182 ( .A(n41519), .B(n41530), .Z(n41521) );
  XNOR U41183 ( .A(n41532), .B(n41533), .Z(n1128) );
  AND U41184 ( .A(n41534), .B(n41535), .Z(n41533) );
  XNOR U41185 ( .A(n41536), .B(n41532), .Z(n41535) );
  IV U41186 ( .A(n41353), .Z(n41536) );
  XOR U41187 ( .A(n41506), .B(n41537), .Z(n41353) );
  AND U41188 ( .A(n1131), .B(n41538), .Z(n41537) );
  XOR U41189 ( .A(n41396), .B(n41393), .Z(n41538) );
  IV U41190 ( .A(n41506), .Z(n41396) );
  XNOR U41191 ( .A(n41313), .B(n41532), .Z(n41534) );
  XOR U41192 ( .A(n41539), .B(n41540), .Z(n41313) );
  AND U41193 ( .A(n1147), .B(n41541), .Z(n41540) );
  XOR U41194 ( .A(n41526), .B(n41542), .Z(n41532) );
  AND U41195 ( .A(n41543), .B(n41529), .Z(n41542) );
  XNOR U41196 ( .A(n41363), .B(n41526), .Z(n41529) );
  XOR U41197 ( .A(n41413), .B(n41544), .Z(n41363) );
  AND U41198 ( .A(n1131), .B(n41545), .Z(n41544) );
  XOR U41199 ( .A(n41409), .B(n41413), .Z(n41545) );
  XNOR U41200 ( .A(n41546), .B(n41526), .Z(n41543) );
  IV U41201 ( .A(n41321), .Z(n41546) );
  XOR U41202 ( .A(n41547), .B(n41548), .Z(n41321) );
  AND U41203 ( .A(n1147), .B(n41549), .Z(n41548) );
  XOR U41204 ( .A(n41550), .B(n41551), .Z(n41526) );
  AND U41205 ( .A(n41552), .B(n41553), .Z(n41551) );
  XNOR U41206 ( .A(n41373), .B(n41550), .Z(n41553) );
  XOR U41207 ( .A(n41441), .B(n41554), .Z(n41373) );
  AND U41208 ( .A(n1131), .B(n41555), .Z(n41554) );
  XOR U41209 ( .A(n41437), .B(n41441), .Z(n41555) );
  XOR U41210 ( .A(n41550), .B(n41330), .Z(n41552) );
  XOR U41211 ( .A(n41556), .B(n41557), .Z(n41330) );
  AND U41212 ( .A(n1147), .B(n41558), .Z(n41557) );
  XOR U41213 ( .A(n41559), .B(n41560), .Z(n41550) );
  AND U41214 ( .A(n41561), .B(n41562), .Z(n41560) );
  XNOR U41215 ( .A(n41559), .B(n41381), .Z(n41562) );
  XOR U41216 ( .A(n41490), .B(n41563), .Z(n41381) );
  AND U41217 ( .A(n1131), .B(n41564), .Z(n41563) );
  XOR U41218 ( .A(n41486), .B(n41490), .Z(n41564) );
  XNOR U41219 ( .A(n41565), .B(n41559), .Z(n41561) );
  IV U41220 ( .A(n41340), .Z(n41565) );
  XOR U41221 ( .A(n41566), .B(n41567), .Z(n41340) );
  AND U41222 ( .A(n1147), .B(n41568), .Z(n41567) );
  AND U41223 ( .A(n41530), .B(n41519), .Z(n41559) );
  XNOR U41224 ( .A(n41569), .B(n41570), .Z(n41519) );
  AND U41225 ( .A(n1131), .B(n41501), .Z(n41570) );
  XNOR U41226 ( .A(n41499), .B(n41569), .Z(n41501) );
  XNOR U41227 ( .A(n41571), .B(n41572), .Z(n1131) );
  AND U41228 ( .A(n41573), .B(n41574), .Z(n41572) );
  XNOR U41229 ( .A(n41571), .B(n41393), .Z(n41574) );
  IV U41230 ( .A(n41397), .Z(n41393) );
  XOR U41231 ( .A(n41575), .B(n41576), .Z(n41397) );
  AND U41232 ( .A(n1135), .B(n41577), .Z(n41576) );
  XOR U41233 ( .A(n41578), .B(n41575), .Z(n41577) );
  XNOR U41234 ( .A(n41571), .B(n41506), .Z(n41573) );
  XOR U41235 ( .A(n41579), .B(n41580), .Z(n41506) );
  AND U41236 ( .A(n1143), .B(n41541), .Z(n41580) );
  XOR U41237 ( .A(n41539), .B(n41579), .Z(n41541) );
  XOR U41238 ( .A(n41581), .B(n41582), .Z(n41571) );
  AND U41239 ( .A(n41583), .B(n41584), .Z(n41582) );
  XNOR U41240 ( .A(n41581), .B(n41409), .Z(n41584) );
  IV U41241 ( .A(n41412), .Z(n41409) );
  XOR U41242 ( .A(n41585), .B(n41586), .Z(n41412) );
  AND U41243 ( .A(n1135), .B(n41587), .Z(n41586) );
  XOR U41244 ( .A(n41588), .B(n41585), .Z(n41587) );
  XOR U41245 ( .A(n41413), .B(n41581), .Z(n41583) );
  XOR U41246 ( .A(n41589), .B(n41590), .Z(n41413) );
  AND U41247 ( .A(n1143), .B(n41549), .Z(n41590) );
  XOR U41248 ( .A(n41589), .B(n41547), .Z(n41549) );
  XOR U41249 ( .A(n41591), .B(n41592), .Z(n41581) );
  AND U41250 ( .A(n41593), .B(n41594), .Z(n41592) );
  XNOR U41251 ( .A(n41591), .B(n41437), .Z(n41594) );
  IV U41252 ( .A(n41440), .Z(n41437) );
  XOR U41253 ( .A(n41595), .B(n41596), .Z(n41440) );
  AND U41254 ( .A(n1135), .B(n41597), .Z(n41596) );
  XNOR U41255 ( .A(n41598), .B(n41595), .Z(n41597) );
  XOR U41256 ( .A(n41441), .B(n41591), .Z(n41593) );
  XOR U41257 ( .A(n41599), .B(n41600), .Z(n41441) );
  AND U41258 ( .A(n1143), .B(n41558), .Z(n41600) );
  XOR U41259 ( .A(n41599), .B(n41556), .Z(n41558) );
  XOR U41260 ( .A(n41515), .B(n41601), .Z(n41591) );
  AND U41261 ( .A(n41517), .B(n41602), .Z(n41601) );
  XNOR U41262 ( .A(n41515), .B(n41486), .Z(n41602) );
  IV U41263 ( .A(n41489), .Z(n41486) );
  XOR U41264 ( .A(n41603), .B(n41604), .Z(n41489) );
  AND U41265 ( .A(n1135), .B(n41605), .Z(n41604) );
  XOR U41266 ( .A(n41606), .B(n41603), .Z(n41605) );
  XOR U41267 ( .A(n41490), .B(n41515), .Z(n41517) );
  XOR U41268 ( .A(n41607), .B(n41608), .Z(n41490) );
  AND U41269 ( .A(n1143), .B(n41568), .Z(n41608) );
  XOR U41270 ( .A(n41607), .B(n41566), .Z(n41568) );
  AND U41271 ( .A(n41569), .B(n41499), .Z(n41515) );
  XNOR U41272 ( .A(n41609), .B(n41610), .Z(n41499) );
  AND U41273 ( .A(n1135), .B(n41611), .Z(n41610) );
  XNOR U41274 ( .A(n41612), .B(n41609), .Z(n41611) );
  XNOR U41275 ( .A(n41613), .B(n41614), .Z(n1135) );
  AND U41276 ( .A(n41615), .B(n41616), .Z(n41614) );
  XOR U41277 ( .A(n41578), .B(n41613), .Z(n41616) );
  AND U41278 ( .A(n41617), .B(n41618), .Z(n41578) );
  XNOR U41279 ( .A(n41575), .B(n41613), .Z(n41615) );
  XNOR U41280 ( .A(n41619), .B(n41620), .Z(n41575) );
  AND U41281 ( .A(n1139), .B(n41621), .Z(n41620) );
  XNOR U41282 ( .A(n41622), .B(n41623), .Z(n41621) );
  XOR U41283 ( .A(n41624), .B(n41625), .Z(n41613) );
  AND U41284 ( .A(n41626), .B(n41627), .Z(n41625) );
  XNOR U41285 ( .A(n41624), .B(n41617), .Z(n41627) );
  IV U41286 ( .A(n41588), .Z(n41617) );
  XOR U41287 ( .A(n41628), .B(n41629), .Z(n41588) );
  XOR U41288 ( .A(n41630), .B(n41618), .Z(n41629) );
  AND U41289 ( .A(n41598), .B(n41631), .Z(n41618) );
  AND U41290 ( .A(n41632), .B(n41633), .Z(n41630) );
  XOR U41291 ( .A(n41634), .B(n41628), .Z(n41632) );
  XNOR U41292 ( .A(n41585), .B(n41624), .Z(n41626) );
  XNOR U41293 ( .A(n41635), .B(n41636), .Z(n41585) );
  AND U41294 ( .A(n1139), .B(n41637), .Z(n41636) );
  XNOR U41295 ( .A(n41638), .B(n41639), .Z(n41637) );
  XOR U41296 ( .A(n41640), .B(n41641), .Z(n41624) );
  AND U41297 ( .A(n41642), .B(n41643), .Z(n41641) );
  XNOR U41298 ( .A(n41640), .B(n41598), .Z(n41643) );
  XOR U41299 ( .A(n41644), .B(n41633), .Z(n41598) );
  XNOR U41300 ( .A(n41645), .B(n41628), .Z(n41633) );
  XOR U41301 ( .A(n41646), .B(n41647), .Z(n41628) );
  AND U41302 ( .A(n41648), .B(n41649), .Z(n41647) );
  XOR U41303 ( .A(n41650), .B(n41646), .Z(n41648) );
  XNOR U41304 ( .A(n41651), .B(n41652), .Z(n41645) );
  AND U41305 ( .A(n41653), .B(n41654), .Z(n41652) );
  XOR U41306 ( .A(n41651), .B(n41655), .Z(n41653) );
  XNOR U41307 ( .A(n41634), .B(n41631), .Z(n41644) );
  AND U41308 ( .A(n41656), .B(n41657), .Z(n41631) );
  XOR U41309 ( .A(n41658), .B(n41659), .Z(n41634) );
  AND U41310 ( .A(n41660), .B(n41661), .Z(n41659) );
  XOR U41311 ( .A(n41658), .B(n41662), .Z(n41660) );
  XNOR U41312 ( .A(n41595), .B(n41640), .Z(n41642) );
  XNOR U41313 ( .A(n41663), .B(n41664), .Z(n41595) );
  AND U41314 ( .A(n1139), .B(n41665), .Z(n41664) );
  XNOR U41315 ( .A(n41666), .B(n41667), .Z(n41665) );
  XOR U41316 ( .A(n41668), .B(n41669), .Z(n41640) );
  AND U41317 ( .A(n41670), .B(n41671), .Z(n41669) );
  XNOR U41318 ( .A(n41668), .B(n41656), .Z(n41671) );
  IV U41319 ( .A(n41606), .Z(n41656) );
  XNOR U41320 ( .A(n41672), .B(n41649), .Z(n41606) );
  XNOR U41321 ( .A(n41673), .B(n41655), .Z(n41649) );
  XOR U41322 ( .A(n41674), .B(n41675), .Z(n41655) );
  NOR U41323 ( .A(n41676), .B(n41677), .Z(n41675) );
  XNOR U41324 ( .A(n41674), .B(n41678), .Z(n41676) );
  XNOR U41325 ( .A(n41654), .B(n41646), .Z(n41673) );
  XOR U41326 ( .A(n41679), .B(n41680), .Z(n41646) );
  AND U41327 ( .A(n41681), .B(n41682), .Z(n41680) );
  XNOR U41328 ( .A(n41679), .B(n41683), .Z(n41681) );
  XNOR U41329 ( .A(n41684), .B(n41651), .Z(n41654) );
  XOR U41330 ( .A(n41685), .B(n41686), .Z(n41651) );
  AND U41331 ( .A(n41687), .B(n41688), .Z(n41686) );
  XOR U41332 ( .A(n41685), .B(n41689), .Z(n41687) );
  XNOR U41333 ( .A(n41690), .B(n41691), .Z(n41684) );
  NOR U41334 ( .A(n41692), .B(n41693), .Z(n41691) );
  XOR U41335 ( .A(n41690), .B(n41694), .Z(n41692) );
  XNOR U41336 ( .A(n41650), .B(n41657), .Z(n41672) );
  NOR U41337 ( .A(n41612), .B(n41695), .Z(n41657) );
  XOR U41338 ( .A(n41662), .B(n41661), .Z(n41650) );
  XNOR U41339 ( .A(n41696), .B(n41658), .Z(n41661) );
  XOR U41340 ( .A(n41697), .B(n41698), .Z(n41658) );
  AND U41341 ( .A(n41699), .B(n41700), .Z(n41698) );
  XOR U41342 ( .A(n41697), .B(n41701), .Z(n41699) );
  XNOR U41343 ( .A(n41702), .B(n41703), .Z(n41696) );
  NOR U41344 ( .A(n41704), .B(n41705), .Z(n41703) );
  XNOR U41345 ( .A(n41702), .B(n41706), .Z(n41704) );
  XOR U41346 ( .A(n41707), .B(n41708), .Z(n41662) );
  NOR U41347 ( .A(n41709), .B(n41710), .Z(n41708) );
  XNOR U41348 ( .A(n41707), .B(n41711), .Z(n41709) );
  XNOR U41349 ( .A(n41603), .B(n41668), .Z(n41670) );
  XNOR U41350 ( .A(n41712), .B(n41713), .Z(n41603) );
  AND U41351 ( .A(n1139), .B(n41714), .Z(n41713) );
  XNOR U41352 ( .A(n41715), .B(n41716), .Z(n41714) );
  AND U41353 ( .A(n41609), .B(n41612), .Z(n41668) );
  XOR U41354 ( .A(n41717), .B(n41695), .Z(n41612) );
  XNOR U41355 ( .A(p_input[2048]), .B(p_input[896]), .Z(n41695) );
  XOR U41356 ( .A(n41683), .B(n41682), .Z(n41717) );
  XNOR U41357 ( .A(n41718), .B(n41689), .Z(n41682) );
  XNOR U41358 ( .A(n41678), .B(n41677), .Z(n41689) );
  XOR U41359 ( .A(n41719), .B(n41674), .Z(n41677) );
  XNOR U41360 ( .A(n29266), .B(p_input[906]), .Z(n41674) );
  XNOR U41361 ( .A(p_input[2059]), .B(p_input[907]), .Z(n41719) );
  XOR U41362 ( .A(p_input[2060]), .B(p_input[908]), .Z(n41678) );
  XNOR U41363 ( .A(n41688), .B(n41679), .Z(n41718) );
  XNOR U41364 ( .A(n29494), .B(p_input[897]), .Z(n41679) );
  XOR U41365 ( .A(n41720), .B(n41694), .Z(n41688) );
  XNOR U41366 ( .A(p_input[2063]), .B(p_input[911]), .Z(n41694) );
  XOR U41367 ( .A(n41685), .B(n41693), .Z(n41720) );
  XOR U41368 ( .A(n41721), .B(n41690), .Z(n41693) );
  XOR U41369 ( .A(p_input[2061]), .B(p_input[909]), .Z(n41690) );
  XNOR U41370 ( .A(p_input[2062]), .B(p_input[910]), .Z(n41721) );
  XNOR U41371 ( .A(n29036), .B(p_input[905]), .Z(n41685) );
  XNOR U41372 ( .A(n41701), .B(n41700), .Z(n41683) );
  XNOR U41373 ( .A(n41722), .B(n41706), .Z(n41700) );
  XOR U41374 ( .A(p_input[2056]), .B(p_input[904]), .Z(n41706) );
  XOR U41375 ( .A(n41697), .B(n41705), .Z(n41722) );
  XOR U41376 ( .A(n41723), .B(n41702), .Z(n41705) );
  XOR U41377 ( .A(p_input[2054]), .B(p_input[902]), .Z(n41702) );
  XNOR U41378 ( .A(p_input[2055]), .B(p_input[903]), .Z(n41723) );
  XNOR U41379 ( .A(n29039), .B(p_input[898]), .Z(n41697) );
  XNOR U41380 ( .A(n41711), .B(n41710), .Z(n41701) );
  XOR U41381 ( .A(n41724), .B(n41707), .Z(n41710) );
  XOR U41382 ( .A(p_input[2051]), .B(p_input[899]), .Z(n41707) );
  XNOR U41383 ( .A(p_input[2052]), .B(p_input[900]), .Z(n41724) );
  XOR U41384 ( .A(p_input[2053]), .B(p_input[901]), .Z(n41711) );
  XNOR U41385 ( .A(n41725), .B(n41726), .Z(n41609) );
  AND U41386 ( .A(n1139), .B(n41727), .Z(n41726) );
  XNOR U41387 ( .A(n41728), .B(n41729), .Z(n1139) );
  AND U41388 ( .A(n41730), .B(n41731), .Z(n41729) );
  XOR U41389 ( .A(n41623), .B(n41728), .Z(n41731) );
  XNOR U41390 ( .A(n41732), .B(n41728), .Z(n41730) );
  XOR U41391 ( .A(n41733), .B(n41734), .Z(n41728) );
  AND U41392 ( .A(n41735), .B(n41736), .Z(n41734) );
  XOR U41393 ( .A(n41638), .B(n41733), .Z(n41736) );
  XOR U41394 ( .A(n41733), .B(n41639), .Z(n41735) );
  XOR U41395 ( .A(n41737), .B(n41738), .Z(n41733) );
  AND U41396 ( .A(n41739), .B(n41740), .Z(n41738) );
  XOR U41397 ( .A(n41666), .B(n41737), .Z(n41740) );
  XOR U41398 ( .A(n41737), .B(n41667), .Z(n41739) );
  XOR U41399 ( .A(n41741), .B(n41742), .Z(n41737) );
  AND U41400 ( .A(n41743), .B(n41744), .Z(n41742) );
  XOR U41401 ( .A(n41741), .B(n41715), .Z(n41744) );
  XNOR U41402 ( .A(n41745), .B(n41746), .Z(n41569) );
  AND U41403 ( .A(n1143), .B(n41747), .Z(n41746) );
  XNOR U41404 ( .A(n41748), .B(n41749), .Z(n1143) );
  AND U41405 ( .A(n41750), .B(n41751), .Z(n41749) );
  XOR U41406 ( .A(n41748), .B(n41579), .Z(n41751) );
  XNOR U41407 ( .A(n41748), .B(n41539), .Z(n41750) );
  XOR U41408 ( .A(n41752), .B(n41753), .Z(n41748) );
  AND U41409 ( .A(n41754), .B(n41755), .Z(n41753) );
  XOR U41410 ( .A(n41752), .B(n41547), .Z(n41754) );
  XOR U41411 ( .A(n41756), .B(n41757), .Z(n41530) );
  AND U41412 ( .A(n1147), .B(n41747), .Z(n41757) );
  XNOR U41413 ( .A(n41745), .B(n41756), .Z(n41747) );
  XNOR U41414 ( .A(n41758), .B(n41759), .Z(n1147) );
  AND U41415 ( .A(n41760), .B(n41761), .Z(n41759) );
  XNOR U41416 ( .A(n41762), .B(n41758), .Z(n41761) );
  IV U41417 ( .A(n41579), .Z(n41762) );
  XOR U41418 ( .A(n41732), .B(n41763), .Z(n41579) );
  AND U41419 ( .A(n1150), .B(n41764), .Z(n41763) );
  XOR U41420 ( .A(n41622), .B(n41619), .Z(n41764) );
  IV U41421 ( .A(n41732), .Z(n41622) );
  XNOR U41422 ( .A(n41539), .B(n41758), .Z(n41760) );
  XOR U41423 ( .A(n41765), .B(n41766), .Z(n41539) );
  AND U41424 ( .A(n1166), .B(n41767), .Z(n41766) );
  XOR U41425 ( .A(n41752), .B(n41768), .Z(n41758) );
  AND U41426 ( .A(n41769), .B(n41755), .Z(n41768) );
  XNOR U41427 ( .A(n41589), .B(n41752), .Z(n41755) );
  XOR U41428 ( .A(n41639), .B(n41770), .Z(n41589) );
  AND U41429 ( .A(n1150), .B(n41771), .Z(n41770) );
  XOR U41430 ( .A(n41635), .B(n41639), .Z(n41771) );
  XNOR U41431 ( .A(n41772), .B(n41752), .Z(n41769) );
  IV U41432 ( .A(n41547), .Z(n41772) );
  XOR U41433 ( .A(n41773), .B(n41774), .Z(n41547) );
  AND U41434 ( .A(n1166), .B(n41775), .Z(n41774) );
  XOR U41435 ( .A(n41776), .B(n41777), .Z(n41752) );
  AND U41436 ( .A(n41778), .B(n41779), .Z(n41777) );
  XNOR U41437 ( .A(n41599), .B(n41776), .Z(n41779) );
  XOR U41438 ( .A(n41667), .B(n41780), .Z(n41599) );
  AND U41439 ( .A(n1150), .B(n41781), .Z(n41780) );
  XOR U41440 ( .A(n41663), .B(n41667), .Z(n41781) );
  XOR U41441 ( .A(n41776), .B(n41556), .Z(n41778) );
  XOR U41442 ( .A(n41782), .B(n41783), .Z(n41556) );
  AND U41443 ( .A(n1166), .B(n41784), .Z(n41783) );
  XOR U41444 ( .A(n41785), .B(n41786), .Z(n41776) );
  AND U41445 ( .A(n41787), .B(n41788), .Z(n41786) );
  XNOR U41446 ( .A(n41785), .B(n41607), .Z(n41788) );
  XOR U41447 ( .A(n41716), .B(n41789), .Z(n41607) );
  AND U41448 ( .A(n1150), .B(n41790), .Z(n41789) );
  XOR U41449 ( .A(n41712), .B(n41716), .Z(n41790) );
  XNOR U41450 ( .A(n41791), .B(n41785), .Z(n41787) );
  IV U41451 ( .A(n41566), .Z(n41791) );
  XOR U41452 ( .A(n41792), .B(n41793), .Z(n41566) );
  AND U41453 ( .A(n1166), .B(n41794), .Z(n41793) );
  AND U41454 ( .A(n41756), .B(n41745), .Z(n41785) );
  XNOR U41455 ( .A(n41795), .B(n41796), .Z(n41745) );
  AND U41456 ( .A(n1150), .B(n41727), .Z(n41796) );
  XNOR U41457 ( .A(n41725), .B(n41795), .Z(n41727) );
  XNOR U41458 ( .A(n41797), .B(n41798), .Z(n1150) );
  AND U41459 ( .A(n41799), .B(n41800), .Z(n41798) );
  XNOR U41460 ( .A(n41797), .B(n41619), .Z(n41800) );
  IV U41461 ( .A(n41623), .Z(n41619) );
  XOR U41462 ( .A(n41801), .B(n41802), .Z(n41623) );
  AND U41463 ( .A(n1154), .B(n41803), .Z(n41802) );
  XOR U41464 ( .A(n41804), .B(n41801), .Z(n41803) );
  XNOR U41465 ( .A(n41797), .B(n41732), .Z(n41799) );
  XOR U41466 ( .A(n41805), .B(n41806), .Z(n41732) );
  AND U41467 ( .A(n1162), .B(n41767), .Z(n41806) );
  XOR U41468 ( .A(n41765), .B(n41805), .Z(n41767) );
  XOR U41469 ( .A(n41807), .B(n41808), .Z(n41797) );
  AND U41470 ( .A(n41809), .B(n41810), .Z(n41808) );
  XNOR U41471 ( .A(n41807), .B(n41635), .Z(n41810) );
  IV U41472 ( .A(n41638), .Z(n41635) );
  XOR U41473 ( .A(n41811), .B(n41812), .Z(n41638) );
  AND U41474 ( .A(n1154), .B(n41813), .Z(n41812) );
  XOR U41475 ( .A(n41814), .B(n41811), .Z(n41813) );
  XOR U41476 ( .A(n41639), .B(n41807), .Z(n41809) );
  XOR U41477 ( .A(n41815), .B(n41816), .Z(n41639) );
  AND U41478 ( .A(n1162), .B(n41775), .Z(n41816) );
  XOR U41479 ( .A(n41815), .B(n41773), .Z(n41775) );
  XOR U41480 ( .A(n41817), .B(n41818), .Z(n41807) );
  AND U41481 ( .A(n41819), .B(n41820), .Z(n41818) );
  XNOR U41482 ( .A(n41817), .B(n41663), .Z(n41820) );
  IV U41483 ( .A(n41666), .Z(n41663) );
  XOR U41484 ( .A(n41821), .B(n41822), .Z(n41666) );
  AND U41485 ( .A(n1154), .B(n41823), .Z(n41822) );
  XNOR U41486 ( .A(n41824), .B(n41821), .Z(n41823) );
  XOR U41487 ( .A(n41667), .B(n41817), .Z(n41819) );
  XOR U41488 ( .A(n41825), .B(n41826), .Z(n41667) );
  AND U41489 ( .A(n1162), .B(n41784), .Z(n41826) );
  XOR U41490 ( .A(n41825), .B(n41782), .Z(n41784) );
  XOR U41491 ( .A(n41741), .B(n41827), .Z(n41817) );
  AND U41492 ( .A(n41743), .B(n41828), .Z(n41827) );
  XNOR U41493 ( .A(n41741), .B(n41712), .Z(n41828) );
  IV U41494 ( .A(n41715), .Z(n41712) );
  XOR U41495 ( .A(n41829), .B(n41830), .Z(n41715) );
  AND U41496 ( .A(n1154), .B(n41831), .Z(n41830) );
  XOR U41497 ( .A(n41832), .B(n41829), .Z(n41831) );
  XOR U41498 ( .A(n41716), .B(n41741), .Z(n41743) );
  XOR U41499 ( .A(n41833), .B(n41834), .Z(n41716) );
  AND U41500 ( .A(n1162), .B(n41794), .Z(n41834) );
  XOR U41501 ( .A(n41833), .B(n41792), .Z(n41794) );
  AND U41502 ( .A(n41795), .B(n41725), .Z(n41741) );
  XNOR U41503 ( .A(n41835), .B(n41836), .Z(n41725) );
  AND U41504 ( .A(n1154), .B(n41837), .Z(n41836) );
  XNOR U41505 ( .A(n41838), .B(n41835), .Z(n41837) );
  XNOR U41506 ( .A(n41839), .B(n41840), .Z(n1154) );
  AND U41507 ( .A(n41841), .B(n41842), .Z(n41840) );
  XOR U41508 ( .A(n41804), .B(n41839), .Z(n41842) );
  AND U41509 ( .A(n41843), .B(n41844), .Z(n41804) );
  XNOR U41510 ( .A(n41801), .B(n41839), .Z(n41841) );
  XNOR U41511 ( .A(n41845), .B(n41846), .Z(n41801) );
  AND U41512 ( .A(n1158), .B(n41847), .Z(n41846) );
  XNOR U41513 ( .A(n41848), .B(n41849), .Z(n41847) );
  XOR U41514 ( .A(n41850), .B(n41851), .Z(n41839) );
  AND U41515 ( .A(n41852), .B(n41853), .Z(n41851) );
  XNOR U41516 ( .A(n41850), .B(n41843), .Z(n41853) );
  IV U41517 ( .A(n41814), .Z(n41843) );
  XOR U41518 ( .A(n41854), .B(n41855), .Z(n41814) );
  XOR U41519 ( .A(n41856), .B(n41844), .Z(n41855) );
  AND U41520 ( .A(n41824), .B(n41857), .Z(n41844) );
  AND U41521 ( .A(n41858), .B(n41859), .Z(n41856) );
  XOR U41522 ( .A(n41860), .B(n41854), .Z(n41858) );
  XNOR U41523 ( .A(n41811), .B(n41850), .Z(n41852) );
  XNOR U41524 ( .A(n41861), .B(n41862), .Z(n41811) );
  AND U41525 ( .A(n1158), .B(n41863), .Z(n41862) );
  XNOR U41526 ( .A(n41864), .B(n41865), .Z(n41863) );
  XOR U41527 ( .A(n41866), .B(n41867), .Z(n41850) );
  AND U41528 ( .A(n41868), .B(n41869), .Z(n41867) );
  XNOR U41529 ( .A(n41866), .B(n41824), .Z(n41869) );
  XOR U41530 ( .A(n41870), .B(n41859), .Z(n41824) );
  XNOR U41531 ( .A(n41871), .B(n41854), .Z(n41859) );
  XOR U41532 ( .A(n41872), .B(n41873), .Z(n41854) );
  AND U41533 ( .A(n41874), .B(n41875), .Z(n41873) );
  XOR U41534 ( .A(n41876), .B(n41872), .Z(n41874) );
  XNOR U41535 ( .A(n41877), .B(n41878), .Z(n41871) );
  AND U41536 ( .A(n41879), .B(n41880), .Z(n41878) );
  XOR U41537 ( .A(n41877), .B(n41881), .Z(n41879) );
  XNOR U41538 ( .A(n41860), .B(n41857), .Z(n41870) );
  AND U41539 ( .A(n41882), .B(n41883), .Z(n41857) );
  XOR U41540 ( .A(n41884), .B(n41885), .Z(n41860) );
  AND U41541 ( .A(n41886), .B(n41887), .Z(n41885) );
  XOR U41542 ( .A(n41884), .B(n41888), .Z(n41886) );
  XNOR U41543 ( .A(n41821), .B(n41866), .Z(n41868) );
  XNOR U41544 ( .A(n41889), .B(n41890), .Z(n41821) );
  AND U41545 ( .A(n1158), .B(n41891), .Z(n41890) );
  XNOR U41546 ( .A(n41892), .B(n41893), .Z(n41891) );
  XOR U41547 ( .A(n41894), .B(n41895), .Z(n41866) );
  AND U41548 ( .A(n41896), .B(n41897), .Z(n41895) );
  XNOR U41549 ( .A(n41894), .B(n41882), .Z(n41897) );
  IV U41550 ( .A(n41832), .Z(n41882) );
  XNOR U41551 ( .A(n41898), .B(n41875), .Z(n41832) );
  XNOR U41552 ( .A(n41899), .B(n41881), .Z(n41875) );
  XOR U41553 ( .A(n41900), .B(n41901), .Z(n41881) );
  NOR U41554 ( .A(n41902), .B(n41903), .Z(n41901) );
  XNOR U41555 ( .A(n41900), .B(n41904), .Z(n41902) );
  XNOR U41556 ( .A(n41880), .B(n41872), .Z(n41899) );
  XOR U41557 ( .A(n41905), .B(n41906), .Z(n41872) );
  AND U41558 ( .A(n41907), .B(n41908), .Z(n41906) );
  XNOR U41559 ( .A(n41905), .B(n41909), .Z(n41907) );
  XNOR U41560 ( .A(n41910), .B(n41877), .Z(n41880) );
  XOR U41561 ( .A(n41911), .B(n41912), .Z(n41877) );
  AND U41562 ( .A(n41913), .B(n41914), .Z(n41912) );
  XOR U41563 ( .A(n41911), .B(n41915), .Z(n41913) );
  XNOR U41564 ( .A(n41916), .B(n41917), .Z(n41910) );
  NOR U41565 ( .A(n41918), .B(n41919), .Z(n41917) );
  XOR U41566 ( .A(n41916), .B(n41920), .Z(n41918) );
  XNOR U41567 ( .A(n41876), .B(n41883), .Z(n41898) );
  NOR U41568 ( .A(n41838), .B(n41921), .Z(n41883) );
  XOR U41569 ( .A(n41888), .B(n41887), .Z(n41876) );
  XNOR U41570 ( .A(n41922), .B(n41884), .Z(n41887) );
  XOR U41571 ( .A(n41923), .B(n41924), .Z(n41884) );
  AND U41572 ( .A(n41925), .B(n41926), .Z(n41924) );
  XOR U41573 ( .A(n41923), .B(n41927), .Z(n41925) );
  XNOR U41574 ( .A(n41928), .B(n41929), .Z(n41922) );
  NOR U41575 ( .A(n41930), .B(n41931), .Z(n41929) );
  XNOR U41576 ( .A(n41928), .B(n41932), .Z(n41930) );
  XOR U41577 ( .A(n41933), .B(n41934), .Z(n41888) );
  NOR U41578 ( .A(n41935), .B(n41936), .Z(n41934) );
  XNOR U41579 ( .A(n41933), .B(n41937), .Z(n41935) );
  XNOR U41580 ( .A(n41829), .B(n41894), .Z(n41896) );
  XNOR U41581 ( .A(n41938), .B(n41939), .Z(n41829) );
  AND U41582 ( .A(n1158), .B(n41940), .Z(n41939) );
  XNOR U41583 ( .A(n41941), .B(n41942), .Z(n41940) );
  AND U41584 ( .A(n41835), .B(n41838), .Z(n41894) );
  XOR U41585 ( .A(n41943), .B(n41921), .Z(n41838) );
  XNOR U41586 ( .A(p_input[2048]), .B(p_input[912]), .Z(n41921) );
  XOR U41587 ( .A(n41909), .B(n41908), .Z(n41943) );
  XNOR U41588 ( .A(n41944), .B(n41915), .Z(n41908) );
  XNOR U41589 ( .A(n41904), .B(n41903), .Z(n41915) );
  XOR U41590 ( .A(n41945), .B(n41900), .Z(n41903) );
  XNOR U41591 ( .A(n29266), .B(p_input[922]), .Z(n41900) );
  XNOR U41592 ( .A(p_input[2059]), .B(p_input[923]), .Z(n41945) );
  XOR U41593 ( .A(p_input[2060]), .B(p_input[924]), .Z(n41904) );
  XNOR U41594 ( .A(n41914), .B(n41905), .Z(n41944) );
  XNOR U41595 ( .A(n29494), .B(p_input[913]), .Z(n41905) );
  XOR U41596 ( .A(n41946), .B(n41920), .Z(n41914) );
  XNOR U41597 ( .A(p_input[2063]), .B(p_input[927]), .Z(n41920) );
  XOR U41598 ( .A(n41911), .B(n41919), .Z(n41946) );
  XOR U41599 ( .A(n41947), .B(n41916), .Z(n41919) );
  XOR U41600 ( .A(p_input[2061]), .B(p_input[925]), .Z(n41916) );
  XNOR U41601 ( .A(p_input[2062]), .B(p_input[926]), .Z(n41947) );
  XNOR U41602 ( .A(n29036), .B(p_input[921]), .Z(n41911) );
  XNOR U41603 ( .A(n41927), .B(n41926), .Z(n41909) );
  XNOR U41604 ( .A(n41948), .B(n41932), .Z(n41926) );
  XOR U41605 ( .A(p_input[2056]), .B(p_input[920]), .Z(n41932) );
  XOR U41606 ( .A(n41923), .B(n41931), .Z(n41948) );
  XOR U41607 ( .A(n41949), .B(n41928), .Z(n41931) );
  XOR U41608 ( .A(p_input[2054]), .B(p_input[918]), .Z(n41928) );
  XNOR U41609 ( .A(p_input[2055]), .B(p_input[919]), .Z(n41949) );
  XNOR U41610 ( .A(n29039), .B(p_input[914]), .Z(n41923) );
  XNOR U41611 ( .A(n41937), .B(n41936), .Z(n41927) );
  XOR U41612 ( .A(n41950), .B(n41933), .Z(n41936) );
  XOR U41613 ( .A(p_input[2051]), .B(p_input[915]), .Z(n41933) );
  XNOR U41614 ( .A(p_input[2052]), .B(p_input[916]), .Z(n41950) );
  XOR U41615 ( .A(p_input[2053]), .B(p_input[917]), .Z(n41937) );
  XNOR U41616 ( .A(n41951), .B(n41952), .Z(n41835) );
  AND U41617 ( .A(n1158), .B(n41953), .Z(n41952) );
  XNOR U41618 ( .A(n41954), .B(n41955), .Z(n1158) );
  AND U41619 ( .A(n41956), .B(n41957), .Z(n41955) );
  XOR U41620 ( .A(n41849), .B(n41954), .Z(n41957) );
  XNOR U41621 ( .A(n41958), .B(n41954), .Z(n41956) );
  XOR U41622 ( .A(n41959), .B(n41960), .Z(n41954) );
  AND U41623 ( .A(n41961), .B(n41962), .Z(n41960) );
  XOR U41624 ( .A(n41864), .B(n41959), .Z(n41962) );
  XOR U41625 ( .A(n41959), .B(n41865), .Z(n41961) );
  XOR U41626 ( .A(n41963), .B(n41964), .Z(n41959) );
  AND U41627 ( .A(n41965), .B(n41966), .Z(n41964) );
  XOR U41628 ( .A(n41892), .B(n41963), .Z(n41966) );
  XOR U41629 ( .A(n41963), .B(n41893), .Z(n41965) );
  XOR U41630 ( .A(n41967), .B(n41968), .Z(n41963) );
  AND U41631 ( .A(n41969), .B(n41970), .Z(n41968) );
  XOR U41632 ( .A(n41967), .B(n41941), .Z(n41970) );
  XNOR U41633 ( .A(n41971), .B(n41972), .Z(n41795) );
  AND U41634 ( .A(n1162), .B(n41973), .Z(n41972) );
  XNOR U41635 ( .A(n41974), .B(n41975), .Z(n1162) );
  AND U41636 ( .A(n41976), .B(n41977), .Z(n41975) );
  XOR U41637 ( .A(n41974), .B(n41805), .Z(n41977) );
  XNOR U41638 ( .A(n41974), .B(n41765), .Z(n41976) );
  XOR U41639 ( .A(n41978), .B(n41979), .Z(n41974) );
  AND U41640 ( .A(n41980), .B(n41981), .Z(n41979) );
  XOR U41641 ( .A(n41978), .B(n41773), .Z(n41980) );
  XOR U41642 ( .A(n41982), .B(n41983), .Z(n41756) );
  AND U41643 ( .A(n1166), .B(n41973), .Z(n41983) );
  XNOR U41644 ( .A(n41971), .B(n41982), .Z(n41973) );
  XNOR U41645 ( .A(n41984), .B(n41985), .Z(n1166) );
  AND U41646 ( .A(n41986), .B(n41987), .Z(n41985) );
  XNOR U41647 ( .A(n41988), .B(n41984), .Z(n41987) );
  IV U41648 ( .A(n41805), .Z(n41988) );
  XOR U41649 ( .A(n41958), .B(n41989), .Z(n41805) );
  AND U41650 ( .A(n1169), .B(n41990), .Z(n41989) );
  XOR U41651 ( .A(n41848), .B(n41845), .Z(n41990) );
  IV U41652 ( .A(n41958), .Z(n41848) );
  XNOR U41653 ( .A(n41765), .B(n41984), .Z(n41986) );
  XOR U41654 ( .A(n41991), .B(n41992), .Z(n41765) );
  AND U41655 ( .A(n1185), .B(n41993), .Z(n41992) );
  XOR U41656 ( .A(n41978), .B(n41994), .Z(n41984) );
  AND U41657 ( .A(n41995), .B(n41981), .Z(n41994) );
  XNOR U41658 ( .A(n41815), .B(n41978), .Z(n41981) );
  XOR U41659 ( .A(n41865), .B(n41996), .Z(n41815) );
  AND U41660 ( .A(n1169), .B(n41997), .Z(n41996) );
  XOR U41661 ( .A(n41861), .B(n41865), .Z(n41997) );
  XNOR U41662 ( .A(n41998), .B(n41978), .Z(n41995) );
  IV U41663 ( .A(n41773), .Z(n41998) );
  XOR U41664 ( .A(n41999), .B(n42000), .Z(n41773) );
  AND U41665 ( .A(n1185), .B(n42001), .Z(n42000) );
  XOR U41666 ( .A(n42002), .B(n42003), .Z(n41978) );
  AND U41667 ( .A(n42004), .B(n42005), .Z(n42003) );
  XNOR U41668 ( .A(n41825), .B(n42002), .Z(n42005) );
  XOR U41669 ( .A(n41893), .B(n42006), .Z(n41825) );
  AND U41670 ( .A(n1169), .B(n42007), .Z(n42006) );
  XOR U41671 ( .A(n41889), .B(n41893), .Z(n42007) );
  XOR U41672 ( .A(n42002), .B(n41782), .Z(n42004) );
  XOR U41673 ( .A(n42008), .B(n42009), .Z(n41782) );
  AND U41674 ( .A(n1185), .B(n42010), .Z(n42009) );
  XOR U41675 ( .A(n42011), .B(n42012), .Z(n42002) );
  AND U41676 ( .A(n42013), .B(n42014), .Z(n42012) );
  XNOR U41677 ( .A(n42011), .B(n41833), .Z(n42014) );
  XOR U41678 ( .A(n41942), .B(n42015), .Z(n41833) );
  AND U41679 ( .A(n1169), .B(n42016), .Z(n42015) );
  XOR U41680 ( .A(n41938), .B(n41942), .Z(n42016) );
  XNOR U41681 ( .A(n42017), .B(n42011), .Z(n42013) );
  IV U41682 ( .A(n41792), .Z(n42017) );
  XOR U41683 ( .A(n42018), .B(n42019), .Z(n41792) );
  AND U41684 ( .A(n1185), .B(n42020), .Z(n42019) );
  AND U41685 ( .A(n41982), .B(n41971), .Z(n42011) );
  XNOR U41686 ( .A(n42021), .B(n42022), .Z(n41971) );
  AND U41687 ( .A(n1169), .B(n41953), .Z(n42022) );
  XNOR U41688 ( .A(n41951), .B(n42021), .Z(n41953) );
  XNOR U41689 ( .A(n42023), .B(n42024), .Z(n1169) );
  AND U41690 ( .A(n42025), .B(n42026), .Z(n42024) );
  XNOR U41691 ( .A(n42023), .B(n41845), .Z(n42026) );
  IV U41692 ( .A(n41849), .Z(n41845) );
  XOR U41693 ( .A(n42027), .B(n42028), .Z(n41849) );
  AND U41694 ( .A(n1173), .B(n42029), .Z(n42028) );
  XOR U41695 ( .A(n42030), .B(n42027), .Z(n42029) );
  XNOR U41696 ( .A(n42023), .B(n41958), .Z(n42025) );
  XOR U41697 ( .A(n42031), .B(n42032), .Z(n41958) );
  AND U41698 ( .A(n1181), .B(n41993), .Z(n42032) );
  XOR U41699 ( .A(n41991), .B(n42031), .Z(n41993) );
  XOR U41700 ( .A(n42033), .B(n42034), .Z(n42023) );
  AND U41701 ( .A(n42035), .B(n42036), .Z(n42034) );
  XNOR U41702 ( .A(n42033), .B(n41861), .Z(n42036) );
  IV U41703 ( .A(n41864), .Z(n41861) );
  XOR U41704 ( .A(n42037), .B(n42038), .Z(n41864) );
  AND U41705 ( .A(n1173), .B(n42039), .Z(n42038) );
  XOR U41706 ( .A(n42040), .B(n42037), .Z(n42039) );
  XOR U41707 ( .A(n41865), .B(n42033), .Z(n42035) );
  XOR U41708 ( .A(n42041), .B(n42042), .Z(n41865) );
  AND U41709 ( .A(n1181), .B(n42001), .Z(n42042) );
  XOR U41710 ( .A(n42041), .B(n41999), .Z(n42001) );
  XOR U41711 ( .A(n42043), .B(n42044), .Z(n42033) );
  AND U41712 ( .A(n42045), .B(n42046), .Z(n42044) );
  XNOR U41713 ( .A(n42043), .B(n41889), .Z(n42046) );
  IV U41714 ( .A(n41892), .Z(n41889) );
  XOR U41715 ( .A(n42047), .B(n42048), .Z(n41892) );
  AND U41716 ( .A(n1173), .B(n42049), .Z(n42048) );
  XNOR U41717 ( .A(n42050), .B(n42047), .Z(n42049) );
  XOR U41718 ( .A(n41893), .B(n42043), .Z(n42045) );
  XOR U41719 ( .A(n42051), .B(n42052), .Z(n41893) );
  AND U41720 ( .A(n1181), .B(n42010), .Z(n42052) );
  XOR U41721 ( .A(n42051), .B(n42008), .Z(n42010) );
  XOR U41722 ( .A(n41967), .B(n42053), .Z(n42043) );
  AND U41723 ( .A(n41969), .B(n42054), .Z(n42053) );
  XNOR U41724 ( .A(n41967), .B(n41938), .Z(n42054) );
  IV U41725 ( .A(n41941), .Z(n41938) );
  XOR U41726 ( .A(n42055), .B(n42056), .Z(n41941) );
  AND U41727 ( .A(n1173), .B(n42057), .Z(n42056) );
  XOR U41728 ( .A(n42058), .B(n42055), .Z(n42057) );
  XOR U41729 ( .A(n41942), .B(n41967), .Z(n41969) );
  XOR U41730 ( .A(n42059), .B(n42060), .Z(n41942) );
  AND U41731 ( .A(n1181), .B(n42020), .Z(n42060) );
  XOR U41732 ( .A(n42059), .B(n42018), .Z(n42020) );
  AND U41733 ( .A(n42021), .B(n41951), .Z(n41967) );
  XNOR U41734 ( .A(n42061), .B(n42062), .Z(n41951) );
  AND U41735 ( .A(n1173), .B(n42063), .Z(n42062) );
  XNOR U41736 ( .A(n42064), .B(n42061), .Z(n42063) );
  XNOR U41737 ( .A(n42065), .B(n42066), .Z(n1173) );
  AND U41738 ( .A(n42067), .B(n42068), .Z(n42066) );
  XOR U41739 ( .A(n42030), .B(n42065), .Z(n42068) );
  AND U41740 ( .A(n42069), .B(n42070), .Z(n42030) );
  XNOR U41741 ( .A(n42027), .B(n42065), .Z(n42067) );
  XNOR U41742 ( .A(n42071), .B(n42072), .Z(n42027) );
  AND U41743 ( .A(n1177), .B(n42073), .Z(n42072) );
  XNOR U41744 ( .A(n42074), .B(n42075), .Z(n42073) );
  XOR U41745 ( .A(n42076), .B(n42077), .Z(n42065) );
  AND U41746 ( .A(n42078), .B(n42079), .Z(n42077) );
  XNOR U41747 ( .A(n42076), .B(n42069), .Z(n42079) );
  IV U41748 ( .A(n42040), .Z(n42069) );
  XOR U41749 ( .A(n42080), .B(n42081), .Z(n42040) );
  XOR U41750 ( .A(n42082), .B(n42070), .Z(n42081) );
  AND U41751 ( .A(n42050), .B(n42083), .Z(n42070) );
  AND U41752 ( .A(n42084), .B(n42085), .Z(n42082) );
  XOR U41753 ( .A(n42086), .B(n42080), .Z(n42084) );
  XNOR U41754 ( .A(n42037), .B(n42076), .Z(n42078) );
  XNOR U41755 ( .A(n42087), .B(n42088), .Z(n42037) );
  AND U41756 ( .A(n1177), .B(n42089), .Z(n42088) );
  XNOR U41757 ( .A(n42090), .B(n42091), .Z(n42089) );
  XOR U41758 ( .A(n42092), .B(n42093), .Z(n42076) );
  AND U41759 ( .A(n42094), .B(n42095), .Z(n42093) );
  XNOR U41760 ( .A(n42092), .B(n42050), .Z(n42095) );
  XOR U41761 ( .A(n42096), .B(n42085), .Z(n42050) );
  XNOR U41762 ( .A(n42097), .B(n42080), .Z(n42085) );
  XOR U41763 ( .A(n42098), .B(n42099), .Z(n42080) );
  AND U41764 ( .A(n42100), .B(n42101), .Z(n42099) );
  XOR U41765 ( .A(n42102), .B(n42098), .Z(n42100) );
  XNOR U41766 ( .A(n42103), .B(n42104), .Z(n42097) );
  AND U41767 ( .A(n42105), .B(n42106), .Z(n42104) );
  XOR U41768 ( .A(n42103), .B(n42107), .Z(n42105) );
  XNOR U41769 ( .A(n42086), .B(n42083), .Z(n42096) );
  AND U41770 ( .A(n42108), .B(n42109), .Z(n42083) );
  XOR U41771 ( .A(n42110), .B(n42111), .Z(n42086) );
  AND U41772 ( .A(n42112), .B(n42113), .Z(n42111) );
  XOR U41773 ( .A(n42110), .B(n42114), .Z(n42112) );
  XNOR U41774 ( .A(n42047), .B(n42092), .Z(n42094) );
  XNOR U41775 ( .A(n42115), .B(n42116), .Z(n42047) );
  AND U41776 ( .A(n1177), .B(n42117), .Z(n42116) );
  XNOR U41777 ( .A(n42118), .B(n42119), .Z(n42117) );
  XOR U41778 ( .A(n42120), .B(n42121), .Z(n42092) );
  AND U41779 ( .A(n42122), .B(n42123), .Z(n42121) );
  XNOR U41780 ( .A(n42120), .B(n42108), .Z(n42123) );
  IV U41781 ( .A(n42058), .Z(n42108) );
  XNOR U41782 ( .A(n42124), .B(n42101), .Z(n42058) );
  XNOR U41783 ( .A(n42125), .B(n42107), .Z(n42101) );
  XOR U41784 ( .A(n42126), .B(n42127), .Z(n42107) );
  NOR U41785 ( .A(n42128), .B(n42129), .Z(n42127) );
  XNOR U41786 ( .A(n42126), .B(n42130), .Z(n42128) );
  XNOR U41787 ( .A(n42106), .B(n42098), .Z(n42125) );
  XOR U41788 ( .A(n42131), .B(n42132), .Z(n42098) );
  AND U41789 ( .A(n42133), .B(n42134), .Z(n42132) );
  XNOR U41790 ( .A(n42131), .B(n42135), .Z(n42133) );
  XNOR U41791 ( .A(n42136), .B(n42103), .Z(n42106) );
  XOR U41792 ( .A(n42137), .B(n42138), .Z(n42103) );
  AND U41793 ( .A(n42139), .B(n42140), .Z(n42138) );
  XOR U41794 ( .A(n42137), .B(n42141), .Z(n42139) );
  XNOR U41795 ( .A(n42142), .B(n42143), .Z(n42136) );
  NOR U41796 ( .A(n42144), .B(n42145), .Z(n42143) );
  XOR U41797 ( .A(n42142), .B(n42146), .Z(n42144) );
  XNOR U41798 ( .A(n42102), .B(n42109), .Z(n42124) );
  NOR U41799 ( .A(n42064), .B(n42147), .Z(n42109) );
  XOR U41800 ( .A(n42114), .B(n42113), .Z(n42102) );
  XNOR U41801 ( .A(n42148), .B(n42110), .Z(n42113) );
  XOR U41802 ( .A(n42149), .B(n42150), .Z(n42110) );
  AND U41803 ( .A(n42151), .B(n42152), .Z(n42150) );
  XOR U41804 ( .A(n42149), .B(n42153), .Z(n42151) );
  XNOR U41805 ( .A(n42154), .B(n42155), .Z(n42148) );
  NOR U41806 ( .A(n42156), .B(n42157), .Z(n42155) );
  XNOR U41807 ( .A(n42154), .B(n42158), .Z(n42156) );
  XOR U41808 ( .A(n42159), .B(n42160), .Z(n42114) );
  NOR U41809 ( .A(n42161), .B(n42162), .Z(n42160) );
  XNOR U41810 ( .A(n42159), .B(n42163), .Z(n42161) );
  XNOR U41811 ( .A(n42055), .B(n42120), .Z(n42122) );
  XNOR U41812 ( .A(n42164), .B(n42165), .Z(n42055) );
  AND U41813 ( .A(n1177), .B(n42166), .Z(n42165) );
  XNOR U41814 ( .A(n42167), .B(n42168), .Z(n42166) );
  AND U41815 ( .A(n42061), .B(n42064), .Z(n42120) );
  XOR U41816 ( .A(n42169), .B(n42147), .Z(n42064) );
  XNOR U41817 ( .A(p_input[2048]), .B(p_input[928]), .Z(n42147) );
  XOR U41818 ( .A(n42135), .B(n42134), .Z(n42169) );
  XNOR U41819 ( .A(n42170), .B(n42141), .Z(n42134) );
  XNOR U41820 ( .A(n42130), .B(n42129), .Z(n42141) );
  XOR U41821 ( .A(n42171), .B(n42126), .Z(n42129) );
  XNOR U41822 ( .A(n29266), .B(p_input[938]), .Z(n42126) );
  XNOR U41823 ( .A(p_input[2059]), .B(p_input[939]), .Z(n42171) );
  XOR U41824 ( .A(p_input[2060]), .B(p_input[940]), .Z(n42130) );
  XNOR U41825 ( .A(n42140), .B(n42131), .Z(n42170) );
  XNOR U41826 ( .A(n29494), .B(p_input[929]), .Z(n42131) );
  XOR U41827 ( .A(n42172), .B(n42146), .Z(n42140) );
  XNOR U41828 ( .A(p_input[2063]), .B(p_input[943]), .Z(n42146) );
  XOR U41829 ( .A(n42137), .B(n42145), .Z(n42172) );
  XOR U41830 ( .A(n42173), .B(n42142), .Z(n42145) );
  XOR U41831 ( .A(p_input[2061]), .B(p_input[941]), .Z(n42142) );
  XNOR U41832 ( .A(p_input[2062]), .B(p_input[942]), .Z(n42173) );
  XNOR U41833 ( .A(n29036), .B(p_input[937]), .Z(n42137) );
  XNOR U41834 ( .A(n42153), .B(n42152), .Z(n42135) );
  XNOR U41835 ( .A(n42174), .B(n42158), .Z(n42152) );
  XOR U41836 ( .A(p_input[2056]), .B(p_input[936]), .Z(n42158) );
  XOR U41837 ( .A(n42149), .B(n42157), .Z(n42174) );
  XOR U41838 ( .A(n42175), .B(n42154), .Z(n42157) );
  XOR U41839 ( .A(p_input[2054]), .B(p_input[934]), .Z(n42154) );
  XNOR U41840 ( .A(p_input[2055]), .B(p_input[935]), .Z(n42175) );
  XNOR U41841 ( .A(n29039), .B(p_input[930]), .Z(n42149) );
  XNOR U41842 ( .A(n42163), .B(n42162), .Z(n42153) );
  XOR U41843 ( .A(n42176), .B(n42159), .Z(n42162) );
  XOR U41844 ( .A(p_input[2051]), .B(p_input[931]), .Z(n42159) );
  XNOR U41845 ( .A(p_input[2052]), .B(p_input[932]), .Z(n42176) );
  XOR U41846 ( .A(p_input[2053]), .B(p_input[933]), .Z(n42163) );
  XNOR U41847 ( .A(n42177), .B(n42178), .Z(n42061) );
  AND U41848 ( .A(n1177), .B(n42179), .Z(n42178) );
  XNOR U41849 ( .A(n42180), .B(n42181), .Z(n1177) );
  AND U41850 ( .A(n42182), .B(n42183), .Z(n42181) );
  XOR U41851 ( .A(n42075), .B(n42180), .Z(n42183) );
  XNOR U41852 ( .A(n42184), .B(n42180), .Z(n42182) );
  XOR U41853 ( .A(n42185), .B(n42186), .Z(n42180) );
  AND U41854 ( .A(n42187), .B(n42188), .Z(n42186) );
  XOR U41855 ( .A(n42090), .B(n42185), .Z(n42188) );
  XOR U41856 ( .A(n42185), .B(n42091), .Z(n42187) );
  XOR U41857 ( .A(n42189), .B(n42190), .Z(n42185) );
  AND U41858 ( .A(n42191), .B(n42192), .Z(n42190) );
  XOR U41859 ( .A(n42118), .B(n42189), .Z(n42192) );
  XOR U41860 ( .A(n42189), .B(n42119), .Z(n42191) );
  XOR U41861 ( .A(n42193), .B(n42194), .Z(n42189) );
  AND U41862 ( .A(n42195), .B(n42196), .Z(n42194) );
  XOR U41863 ( .A(n42193), .B(n42167), .Z(n42196) );
  XNOR U41864 ( .A(n42197), .B(n42198), .Z(n42021) );
  AND U41865 ( .A(n1181), .B(n42199), .Z(n42198) );
  XNOR U41866 ( .A(n42200), .B(n42201), .Z(n1181) );
  AND U41867 ( .A(n42202), .B(n42203), .Z(n42201) );
  XOR U41868 ( .A(n42200), .B(n42031), .Z(n42203) );
  XNOR U41869 ( .A(n42200), .B(n41991), .Z(n42202) );
  XOR U41870 ( .A(n42204), .B(n42205), .Z(n42200) );
  AND U41871 ( .A(n42206), .B(n42207), .Z(n42205) );
  XOR U41872 ( .A(n42204), .B(n41999), .Z(n42206) );
  XOR U41873 ( .A(n42208), .B(n42209), .Z(n41982) );
  AND U41874 ( .A(n1185), .B(n42199), .Z(n42209) );
  XNOR U41875 ( .A(n42197), .B(n42208), .Z(n42199) );
  XNOR U41876 ( .A(n42210), .B(n42211), .Z(n1185) );
  AND U41877 ( .A(n42212), .B(n42213), .Z(n42211) );
  XNOR U41878 ( .A(n42214), .B(n42210), .Z(n42213) );
  IV U41879 ( .A(n42031), .Z(n42214) );
  XOR U41880 ( .A(n42184), .B(n42215), .Z(n42031) );
  AND U41881 ( .A(n1188), .B(n42216), .Z(n42215) );
  XOR U41882 ( .A(n42074), .B(n42071), .Z(n42216) );
  IV U41883 ( .A(n42184), .Z(n42074) );
  XNOR U41884 ( .A(n41991), .B(n42210), .Z(n42212) );
  XOR U41885 ( .A(n42217), .B(n42218), .Z(n41991) );
  AND U41886 ( .A(n1204), .B(n42219), .Z(n42218) );
  XOR U41887 ( .A(n42204), .B(n42220), .Z(n42210) );
  AND U41888 ( .A(n42221), .B(n42207), .Z(n42220) );
  XNOR U41889 ( .A(n42041), .B(n42204), .Z(n42207) );
  XOR U41890 ( .A(n42091), .B(n42222), .Z(n42041) );
  AND U41891 ( .A(n1188), .B(n42223), .Z(n42222) );
  XOR U41892 ( .A(n42087), .B(n42091), .Z(n42223) );
  XNOR U41893 ( .A(n42224), .B(n42204), .Z(n42221) );
  IV U41894 ( .A(n41999), .Z(n42224) );
  XOR U41895 ( .A(n42225), .B(n42226), .Z(n41999) );
  AND U41896 ( .A(n1204), .B(n42227), .Z(n42226) );
  XOR U41897 ( .A(n42228), .B(n42229), .Z(n42204) );
  AND U41898 ( .A(n42230), .B(n42231), .Z(n42229) );
  XNOR U41899 ( .A(n42051), .B(n42228), .Z(n42231) );
  XOR U41900 ( .A(n42119), .B(n42232), .Z(n42051) );
  AND U41901 ( .A(n1188), .B(n42233), .Z(n42232) );
  XOR U41902 ( .A(n42115), .B(n42119), .Z(n42233) );
  XOR U41903 ( .A(n42228), .B(n42008), .Z(n42230) );
  XOR U41904 ( .A(n42234), .B(n42235), .Z(n42008) );
  AND U41905 ( .A(n1204), .B(n42236), .Z(n42235) );
  XOR U41906 ( .A(n42237), .B(n42238), .Z(n42228) );
  AND U41907 ( .A(n42239), .B(n42240), .Z(n42238) );
  XNOR U41908 ( .A(n42237), .B(n42059), .Z(n42240) );
  XOR U41909 ( .A(n42168), .B(n42241), .Z(n42059) );
  AND U41910 ( .A(n1188), .B(n42242), .Z(n42241) );
  XOR U41911 ( .A(n42164), .B(n42168), .Z(n42242) );
  XNOR U41912 ( .A(n42243), .B(n42237), .Z(n42239) );
  IV U41913 ( .A(n42018), .Z(n42243) );
  XOR U41914 ( .A(n42244), .B(n42245), .Z(n42018) );
  AND U41915 ( .A(n1204), .B(n42246), .Z(n42245) );
  AND U41916 ( .A(n42208), .B(n42197), .Z(n42237) );
  XNOR U41917 ( .A(n42247), .B(n42248), .Z(n42197) );
  AND U41918 ( .A(n1188), .B(n42179), .Z(n42248) );
  XNOR U41919 ( .A(n42177), .B(n42247), .Z(n42179) );
  XNOR U41920 ( .A(n42249), .B(n42250), .Z(n1188) );
  AND U41921 ( .A(n42251), .B(n42252), .Z(n42250) );
  XNOR U41922 ( .A(n42249), .B(n42071), .Z(n42252) );
  IV U41923 ( .A(n42075), .Z(n42071) );
  XOR U41924 ( .A(n42253), .B(n42254), .Z(n42075) );
  AND U41925 ( .A(n1192), .B(n42255), .Z(n42254) );
  XOR U41926 ( .A(n42256), .B(n42253), .Z(n42255) );
  XNOR U41927 ( .A(n42249), .B(n42184), .Z(n42251) );
  XOR U41928 ( .A(n42257), .B(n42258), .Z(n42184) );
  AND U41929 ( .A(n1200), .B(n42219), .Z(n42258) );
  XOR U41930 ( .A(n42217), .B(n42257), .Z(n42219) );
  XOR U41931 ( .A(n42259), .B(n42260), .Z(n42249) );
  AND U41932 ( .A(n42261), .B(n42262), .Z(n42260) );
  XNOR U41933 ( .A(n42259), .B(n42087), .Z(n42262) );
  IV U41934 ( .A(n42090), .Z(n42087) );
  XOR U41935 ( .A(n42263), .B(n42264), .Z(n42090) );
  AND U41936 ( .A(n1192), .B(n42265), .Z(n42264) );
  XOR U41937 ( .A(n42266), .B(n42263), .Z(n42265) );
  XOR U41938 ( .A(n42091), .B(n42259), .Z(n42261) );
  XOR U41939 ( .A(n42267), .B(n42268), .Z(n42091) );
  AND U41940 ( .A(n1200), .B(n42227), .Z(n42268) );
  XOR U41941 ( .A(n42267), .B(n42225), .Z(n42227) );
  XOR U41942 ( .A(n42269), .B(n42270), .Z(n42259) );
  AND U41943 ( .A(n42271), .B(n42272), .Z(n42270) );
  XNOR U41944 ( .A(n42269), .B(n42115), .Z(n42272) );
  IV U41945 ( .A(n42118), .Z(n42115) );
  XOR U41946 ( .A(n42273), .B(n42274), .Z(n42118) );
  AND U41947 ( .A(n1192), .B(n42275), .Z(n42274) );
  XNOR U41948 ( .A(n42276), .B(n42273), .Z(n42275) );
  XOR U41949 ( .A(n42119), .B(n42269), .Z(n42271) );
  XOR U41950 ( .A(n42277), .B(n42278), .Z(n42119) );
  AND U41951 ( .A(n1200), .B(n42236), .Z(n42278) );
  XOR U41952 ( .A(n42277), .B(n42234), .Z(n42236) );
  XOR U41953 ( .A(n42193), .B(n42279), .Z(n42269) );
  AND U41954 ( .A(n42195), .B(n42280), .Z(n42279) );
  XNOR U41955 ( .A(n42193), .B(n42164), .Z(n42280) );
  IV U41956 ( .A(n42167), .Z(n42164) );
  XOR U41957 ( .A(n42281), .B(n42282), .Z(n42167) );
  AND U41958 ( .A(n1192), .B(n42283), .Z(n42282) );
  XOR U41959 ( .A(n42284), .B(n42281), .Z(n42283) );
  XOR U41960 ( .A(n42168), .B(n42193), .Z(n42195) );
  XOR U41961 ( .A(n42285), .B(n42286), .Z(n42168) );
  AND U41962 ( .A(n1200), .B(n42246), .Z(n42286) );
  XOR U41963 ( .A(n42285), .B(n42244), .Z(n42246) );
  AND U41964 ( .A(n42247), .B(n42177), .Z(n42193) );
  XNOR U41965 ( .A(n42287), .B(n42288), .Z(n42177) );
  AND U41966 ( .A(n1192), .B(n42289), .Z(n42288) );
  XNOR U41967 ( .A(n42290), .B(n42287), .Z(n42289) );
  XNOR U41968 ( .A(n42291), .B(n42292), .Z(n1192) );
  AND U41969 ( .A(n42293), .B(n42294), .Z(n42292) );
  XOR U41970 ( .A(n42256), .B(n42291), .Z(n42294) );
  AND U41971 ( .A(n42295), .B(n42296), .Z(n42256) );
  XNOR U41972 ( .A(n42253), .B(n42291), .Z(n42293) );
  XNOR U41973 ( .A(n42297), .B(n42298), .Z(n42253) );
  AND U41974 ( .A(n1196), .B(n42299), .Z(n42298) );
  XNOR U41975 ( .A(n42300), .B(n42301), .Z(n42299) );
  XOR U41976 ( .A(n42302), .B(n42303), .Z(n42291) );
  AND U41977 ( .A(n42304), .B(n42305), .Z(n42303) );
  XNOR U41978 ( .A(n42302), .B(n42295), .Z(n42305) );
  IV U41979 ( .A(n42266), .Z(n42295) );
  XOR U41980 ( .A(n42306), .B(n42307), .Z(n42266) );
  XOR U41981 ( .A(n42308), .B(n42296), .Z(n42307) );
  AND U41982 ( .A(n42276), .B(n42309), .Z(n42296) );
  AND U41983 ( .A(n42310), .B(n42311), .Z(n42308) );
  XOR U41984 ( .A(n42312), .B(n42306), .Z(n42310) );
  XNOR U41985 ( .A(n42263), .B(n42302), .Z(n42304) );
  XNOR U41986 ( .A(n42313), .B(n42314), .Z(n42263) );
  AND U41987 ( .A(n1196), .B(n42315), .Z(n42314) );
  XNOR U41988 ( .A(n42316), .B(n42317), .Z(n42315) );
  XOR U41989 ( .A(n42318), .B(n42319), .Z(n42302) );
  AND U41990 ( .A(n42320), .B(n42321), .Z(n42319) );
  XNOR U41991 ( .A(n42318), .B(n42276), .Z(n42321) );
  XOR U41992 ( .A(n42322), .B(n42311), .Z(n42276) );
  XNOR U41993 ( .A(n42323), .B(n42306), .Z(n42311) );
  XOR U41994 ( .A(n42324), .B(n42325), .Z(n42306) );
  AND U41995 ( .A(n42326), .B(n42327), .Z(n42325) );
  XOR U41996 ( .A(n42328), .B(n42324), .Z(n42326) );
  XNOR U41997 ( .A(n42329), .B(n42330), .Z(n42323) );
  AND U41998 ( .A(n42331), .B(n42332), .Z(n42330) );
  XOR U41999 ( .A(n42329), .B(n42333), .Z(n42331) );
  XNOR U42000 ( .A(n42312), .B(n42309), .Z(n42322) );
  AND U42001 ( .A(n42334), .B(n42335), .Z(n42309) );
  XOR U42002 ( .A(n42336), .B(n42337), .Z(n42312) );
  AND U42003 ( .A(n42338), .B(n42339), .Z(n42337) );
  XOR U42004 ( .A(n42336), .B(n42340), .Z(n42338) );
  XNOR U42005 ( .A(n42273), .B(n42318), .Z(n42320) );
  XNOR U42006 ( .A(n42341), .B(n42342), .Z(n42273) );
  AND U42007 ( .A(n1196), .B(n42343), .Z(n42342) );
  XNOR U42008 ( .A(n42344), .B(n42345), .Z(n42343) );
  XOR U42009 ( .A(n42346), .B(n42347), .Z(n42318) );
  AND U42010 ( .A(n42348), .B(n42349), .Z(n42347) );
  XNOR U42011 ( .A(n42346), .B(n42334), .Z(n42349) );
  IV U42012 ( .A(n42284), .Z(n42334) );
  XNOR U42013 ( .A(n42350), .B(n42327), .Z(n42284) );
  XNOR U42014 ( .A(n42351), .B(n42333), .Z(n42327) );
  XOR U42015 ( .A(n42352), .B(n42353), .Z(n42333) );
  NOR U42016 ( .A(n42354), .B(n42355), .Z(n42353) );
  XNOR U42017 ( .A(n42352), .B(n42356), .Z(n42354) );
  XNOR U42018 ( .A(n42332), .B(n42324), .Z(n42351) );
  XOR U42019 ( .A(n42357), .B(n42358), .Z(n42324) );
  AND U42020 ( .A(n42359), .B(n42360), .Z(n42358) );
  XNOR U42021 ( .A(n42357), .B(n42361), .Z(n42359) );
  XNOR U42022 ( .A(n42362), .B(n42329), .Z(n42332) );
  XOR U42023 ( .A(n42363), .B(n42364), .Z(n42329) );
  AND U42024 ( .A(n42365), .B(n42366), .Z(n42364) );
  XOR U42025 ( .A(n42363), .B(n42367), .Z(n42365) );
  XNOR U42026 ( .A(n42368), .B(n42369), .Z(n42362) );
  NOR U42027 ( .A(n42370), .B(n42371), .Z(n42369) );
  XOR U42028 ( .A(n42368), .B(n42372), .Z(n42370) );
  XNOR U42029 ( .A(n42328), .B(n42335), .Z(n42350) );
  NOR U42030 ( .A(n42290), .B(n42373), .Z(n42335) );
  XOR U42031 ( .A(n42340), .B(n42339), .Z(n42328) );
  XNOR U42032 ( .A(n42374), .B(n42336), .Z(n42339) );
  XOR U42033 ( .A(n42375), .B(n42376), .Z(n42336) );
  AND U42034 ( .A(n42377), .B(n42378), .Z(n42376) );
  XOR U42035 ( .A(n42375), .B(n42379), .Z(n42377) );
  XNOR U42036 ( .A(n42380), .B(n42381), .Z(n42374) );
  NOR U42037 ( .A(n42382), .B(n42383), .Z(n42381) );
  XNOR U42038 ( .A(n42380), .B(n42384), .Z(n42382) );
  XOR U42039 ( .A(n42385), .B(n42386), .Z(n42340) );
  NOR U42040 ( .A(n42387), .B(n42388), .Z(n42386) );
  XNOR U42041 ( .A(n42385), .B(n42389), .Z(n42387) );
  XNOR U42042 ( .A(n42281), .B(n42346), .Z(n42348) );
  XNOR U42043 ( .A(n42390), .B(n42391), .Z(n42281) );
  AND U42044 ( .A(n1196), .B(n42392), .Z(n42391) );
  XNOR U42045 ( .A(n42393), .B(n42394), .Z(n42392) );
  AND U42046 ( .A(n42287), .B(n42290), .Z(n42346) );
  XOR U42047 ( .A(n42395), .B(n42373), .Z(n42290) );
  XNOR U42048 ( .A(p_input[2048]), .B(p_input[944]), .Z(n42373) );
  XOR U42049 ( .A(n42361), .B(n42360), .Z(n42395) );
  XNOR U42050 ( .A(n42396), .B(n42367), .Z(n42360) );
  XNOR U42051 ( .A(n42356), .B(n42355), .Z(n42367) );
  XOR U42052 ( .A(n42397), .B(n42352), .Z(n42355) );
  XNOR U42053 ( .A(n29266), .B(p_input[954]), .Z(n42352) );
  XNOR U42054 ( .A(p_input[2059]), .B(p_input[955]), .Z(n42397) );
  XOR U42055 ( .A(p_input[2060]), .B(p_input[956]), .Z(n42356) );
  XNOR U42056 ( .A(n42366), .B(n42357), .Z(n42396) );
  XNOR U42057 ( .A(n29494), .B(p_input[945]), .Z(n42357) );
  XOR U42058 ( .A(n42398), .B(n42372), .Z(n42366) );
  XNOR U42059 ( .A(p_input[2063]), .B(p_input[959]), .Z(n42372) );
  XOR U42060 ( .A(n42363), .B(n42371), .Z(n42398) );
  XOR U42061 ( .A(n42399), .B(n42368), .Z(n42371) );
  XOR U42062 ( .A(p_input[2061]), .B(p_input[957]), .Z(n42368) );
  XNOR U42063 ( .A(p_input[2062]), .B(p_input[958]), .Z(n42399) );
  XNOR U42064 ( .A(n29036), .B(p_input[953]), .Z(n42363) );
  XNOR U42065 ( .A(n42379), .B(n42378), .Z(n42361) );
  XNOR U42066 ( .A(n42400), .B(n42384), .Z(n42378) );
  XOR U42067 ( .A(p_input[2056]), .B(p_input[952]), .Z(n42384) );
  XOR U42068 ( .A(n42375), .B(n42383), .Z(n42400) );
  XOR U42069 ( .A(n42401), .B(n42380), .Z(n42383) );
  XOR U42070 ( .A(p_input[2054]), .B(p_input[950]), .Z(n42380) );
  XNOR U42071 ( .A(p_input[2055]), .B(p_input[951]), .Z(n42401) );
  XNOR U42072 ( .A(n29039), .B(p_input[946]), .Z(n42375) );
  XNOR U42073 ( .A(n42389), .B(n42388), .Z(n42379) );
  XOR U42074 ( .A(n42402), .B(n42385), .Z(n42388) );
  XOR U42075 ( .A(p_input[2051]), .B(p_input[947]), .Z(n42385) );
  XNOR U42076 ( .A(p_input[2052]), .B(p_input[948]), .Z(n42402) );
  XOR U42077 ( .A(p_input[2053]), .B(p_input[949]), .Z(n42389) );
  XNOR U42078 ( .A(n42403), .B(n42404), .Z(n42287) );
  AND U42079 ( .A(n1196), .B(n42405), .Z(n42404) );
  XNOR U42080 ( .A(n42406), .B(n42407), .Z(n1196) );
  AND U42081 ( .A(n42408), .B(n42409), .Z(n42407) );
  XOR U42082 ( .A(n42301), .B(n42406), .Z(n42409) );
  XNOR U42083 ( .A(n42410), .B(n42406), .Z(n42408) );
  XOR U42084 ( .A(n42411), .B(n42412), .Z(n42406) );
  AND U42085 ( .A(n42413), .B(n42414), .Z(n42412) );
  XOR U42086 ( .A(n42316), .B(n42411), .Z(n42414) );
  XOR U42087 ( .A(n42411), .B(n42317), .Z(n42413) );
  XOR U42088 ( .A(n42415), .B(n42416), .Z(n42411) );
  AND U42089 ( .A(n42417), .B(n42418), .Z(n42416) );
  XOR U42090 ( .A(n42344), .B(n42415), .Z(n42418) );
  XOR U42091 ( .A(n42415), .B(n42345), .Z(n42417) );
  XOR U42092 ( .A(n42419), .B(n42420), .Z(n42415) );
  AND U42093 ( .A(n42421), .B(n42422), .Z(n42420) );
  XOR U42094 ( .A(n42419), .B(n42393), .Z(n42422) );
  XNOR U42095 ( .A(n42423), .B(n42424), .Z(n42247) );
  AND U42096 ( .A(n1200), .B(n42425), .Z(n42424) );
  XNOR U42097 ( .A(n42426), .B(n42427), .Z(n1200) );
  AND U42098 ( .A(n42428), .B(n42429), .Z(n42427) );
  XOR U42099 ( .A(n42426), .B(n42257), .Z(n42429) );
  XNOR U42100 ( .A(n42426), .B(n42217), .Z(n42428) );
  XOR U42101 ( .A(n42430), .B(n42431), .Z(n42426) );
  AND U42102 ( .A(n42432), .B(n42433), .Z(n42431) );
  XOR U42103 ( .A(n42430), .B(n42225), .Z(n42432) );
  XOR U42104 ( .A(n42434), .B(n42435), .Z(n42208) );
  AND U42105 ( .A(n1204), .B(n42425), .Z(n42435) );
  XNOR U42106 ( .A(n42423), .B(n42434), .Z(n42425) );
  XNOR U42107 ( .A(n42436), .B(n42437), .Z(n1204) );
  AND U42108 ( .A(n42438), .B(n42439), .Z(n42437) );
  XNOR U42109 ( .A(n42440), .B(n42436), .Z(n42439) );
  IV U42110 ( .A(n42257), .Z(n42440) );
  XOR U42111 ( .A(n42410), .B(n42441), .Z(n42257) );
  AND U42112 ( .A(n1207), .B(n42442), .Z(n42441) );
  XOR U42113 ( .A(n42300), .B(n42297), .Z(n42442) );
  IV U42114 ( .A(n42410), .Z(n42300) );
  XNOR U42115 ( .A(n42217), .B(n42436), .Z(n42438) );
  XOR U42116 ( .A(n42443), .B(n42444), .Z(n42217) );
  AND U42117 ( .A(n1223), .B(n42445), .Z(n42444) );
  XOR U42118 ( .A(n42430), .B(n42446), .Z(n42436) );
  AND U42119 ( .A(n42447), .B(n42433), .Z(n42446) );
  XNOR U42120 ( .A(n42267), .B(n42430), .Z(n42433) );
  XOR U42121 ( .A(n42317), .B(n42448), .Z(n42267) );
  AND U42122 ( .A(n1207), .B(n42449), .Z(n42448) );
  XOR U42123 ( .A(n42313), .B(n42317), .Z(n42449) );
  XNOR U42124 ( .A(n42450), .B(n42430), .Z(n42447) );
  IV U42125 ( .A(n42225), .Z(n42450) );
  XOR U42126 ( .A(n42451), .B(n42452), .Z(n42225) );
  AND U42127 ( .A(n1223), .B(n42453), .Z(n42452) );
  XOR U42128 ( .A(n42454), .B(n42455), .Z(n42430) );
  AND U42129 ( .A(n42456), .B(n42457), .Z(n42455) );
  XNOR U42130 ( .A(n42277), .B(n42454), .Z(n42457) );
  XOR U42131 ( .A(n42345), .B(n42458), .Z(n42277) );
  AND U42132 ( .A(n1207), .B(n42459), .Z(n42458) );
  XOR U42133 ( .A(n42341), .B(n42345), .Z(n42459) );
  XOR U42134 ( .A(n42454), .B(n42234), .Z(n42456) );
  XOR U42135 ( .A(n42460), .B(n42461), .Z(n42234) );
  AND U42136 ( .A(n1223), .B(n42462), .Z(n42461) );
  XOR U42137 ( .A(n42463), .B(n42464), .Z(n42454) );
  AND U42138 ( .A(n42465), .B(n42466), .Z(n42464) );
  XNOR U42139 ( .A(n42463), .B(n42285), .Z(n42466) );
  XOR U42140 ( .A(n42394), .B(n42467), .Z(n42285) );
  AND U42141 ( .A(n1207), .B(n42468), .Z(n42467) );
  XOR U42142 ( .A(n42390), .B(n42394), .Z(n42468) );
  XNOR U42143 ( .A(n42469), .B(n42463), .Z(n42465) );
  IV U42144 ( .A(n42244), .Z(n42469) );
  XOR U42145 ( .A(n42470), .B(n42471), .Z(n42244) );
  AND U42146 ( .A(n1223), .B(n42472), .Z(n42471) );
  AND U42147 ( .A(n42434), .B(n42423), .Z(n42463) );
  XNOR U42148 ( .A(n42473), .B(n42474), .Z(n42423) );
  AND U42149 ( .A(n1207), .B(n42405), .Z(n42474) );
  XNOR U42150 ( .A(n42403), .B(n42473), .Z(n42405) );
  XNOR U42151 ( .A(n42475), .B(n42476), .Z(n1207) );
  AND U42152 ( .A(n42477), .B(n42478), .Z(n42476) );
  XNOR U42153 ( .A(n42475), .B(n42297), .Z(n42478) );
  IV U42154 ( .A(n42301), .Z(n42297) );
  XOR U42155 ( .A(n42479), .B(n42480), .Z(n42301) );
  AND U42156 ( .A(n1211), .B(n42481), .Z(n42480) );
  XOR U42157 ( .A(n42482), .B(n42479), .Z(n42481) );
  XNOR U42158 ( .A(n42475), .B(n42410), .Z(n42477) );
  XOR U42159 ( .A(n42483), .B(n42484), .Z(n42410) );
  AND U42160 ( .A(n1219), .B(n42445), .Z(n42484) );
  XOR U42161 ( .A(n42443), .B(n42483), .Z(n42445) );
  XOR U42162 ( .A(n42485), .B(n42486), .Z(n42475) );
  AND U42163 ( .A(n42487), .B(n42488), .Z(n42486) );
  XNOR U42164 ( .A(n42485), .B(n42313), .Z(n42488) );
  IV U42165 ( .A(n42316), .Z(n42313) );
  XOR U42166 ( .A(n42489), .B(n42490), .Z(n42316) );
  AND U42167 ( .A(n1211), .B(n42491), .Z(n42490) );
  XOR U42168 ( .A(n42492), .B(n42489), .Z(n42491) );
  XOR U42169 ( .A(n42317), .B(n42485), .Z(n42487) );
  XOR U42170 ( .A(n42493), .B(n42494), .Z(n42317) );
  AND U42171 ( .A(n1219), .B(n42453), .Z(n42494) );
  XOR U42172 ( .A(n42493), .B(n42451), .Z(n42453) );
  XOR U42173 ( .A(n42495), .B(n42496), .Z(n42485) );
  AND U42174 ( .A(n42497), .B(n42498), .Z(n42496) );
  XNOR U42175 ( .A(n42495), .B(n42341), .Z(n42498) );
  IV U42176 ( .A(n42344), .Z(n42341) );
  XOR U42177 ( .A(n42499), .B(n42500), .Z(n42344) );
  AND U42178 ( .A(n1211), .B(n42501), .Z(n42500) );
  XNOR U42179 ( .A(n42502), .B(n42499), .Z(n42501) );
  XOR U42180 ( .A(n42345), .B(n42495), .Z(n42497) );
  XOR U42181 ( .A(n42503), .B(n42504), .Z(n42345) );
  AND U42182 ( .A(n1219), .B(n42462), .Z(n42504) );
  XOR U42183 ( .A(n42503), .B(n42460), .Z(n42462) );
  XOR U42184 ( .A(n42419), .B(n42505), .Z(n42495) );
  AND U42185 ( .A(n42421), .B(n42506), .Z(n42505) );
  XNOR U42186 ( .A(n42419), .B(n42390), .Z(n42506) );
  IV U42187 ( .A(n42393), .Z(n42390) );
  XOR U42188 ( .A(n42507), .B(n42508), .Z(n42393) );
  AND U42189 ( .A(n1211), .B(n42509), .Z(n42508) );
  XOR U42190 ( .A(n42510), .B(n42507), .Z(n42509) );
  XOR U42191 ( .A(n42394), .B(n42419), .Z(n42421) );
  XOR U42192 ( .A(n42511), .B(n42512), .Z(n42394) );
  AND U42193 ( .A(n1219), .B(n42472), .Z(n42512) );
  XOR U42194 ( .A(n42511), .B(n42470), .Z(n42472) );
  AND U42195 ( .A(n42473), .B(n42403), .Z(n42419) );
  XNOR U42196 ( .A(n42513), .B(n42514), .Z(n42403) );
  AND U42197 ( .A(n1211), .B(n42515), .Z(n42514) );
  XNOR U42198 ( .A(n42516), .B(n42513), .Z(n42515) );
  XNOR U42199 ( .A(n42517), .B(n42518), .Z(n1211) );
  AND U42200 ( .A(n42519), .B(n42520), .Z(n42518) );
  XOR U42201 ( .A(n42482), .B(n42517), .Z(n42520) );
  AND U42202 ( .A(n42521), .B(n42522), .Z(n42482) );
  XNOR U42203 ( .A(n42479), .B(n42517), .Z(n42519) );
  XNOR U42204 ( .A(n42523), .B(n42524), .Z(n42479) );
  AND U42205 ( .A(n1215), .B(n42525), .Z(n42524) );
  XNOR U42206 ( .A(n42526), .B(n42527), .Z(n42525) );
  XOR U42207 ( .A(n42528), .B(n42529), .Z(n42517) );
  AND U42208 ( .A(n42530), .B(n42531), .Z(n42529) );
  XNOR U42209 ( .A(n42528), .B(n42521), .Z(n42531) );
  IV U42210 ( .A(n42492), .Z(n42521) );
  XOR U42211 ( .A(n42532), .B(n42533), .Z(n42492) );
  XOR U42212 ( .A(n42534), .B(n42522), .Z(n42533) );
  AND U42213 ( .A(n42502), .B(n42535), .Z(n42522) );
  AND U42214 ( .A(n42536), .B(n42537), .Z(n42534) );
  XOR U42215 ( .A(n42538), .B(n42532), .Z(n42536) );
  XNOR U42216 ( .A(n42489), .B(n42528), .Z(n42530) );
  XNOR U42217 ( .A(n42539), .B(n42540), .Z(n42489) );
  AND U42218 ( .A(n1215), .B(n42541), .Z(n42540) );
  XNOR U42219 ( .A(n42542), .B(n42543), .Z(n42541) );
  XOR U42220 ( .A(n42544), .B(n42545), .Z(n42528) );
  AND U42221 ( .A(n42546), .B(n42547), .Z(n42545) );
  XNOR U42222 ( .A(n42544), .B(n42502), .Z(n42547) );
  XOR U42223 ( .A(n42548), .B(n42537), .Z(n42502) );
  XNOR U42224 ( .A(n42549), .B(n42532), .Z(n42537) );
  XOR U42225 ( .A(n42550), .B(n42551), .Z(n42532) );
  AND U42226 ( .A(n42552), .B(n42553), .Z(n42551) );
  XOR U42227 ( .A(n42554), .B(n42550), .Z(n42552) );
  XNOR U42228 ( .A(n42555), .B(n42556), .Z(n42549) );
  AND U42229 ( .A(n42557), .B(n42558), .Z(n42556) );
  XOR U42230 ( .A(n42555), .B(n42559), .Z(n42557) );
  XNOR U42231 ( .A(n42538), .B(n42535), .Z(n42548) );
  AND U42232 ( .A(n42560), .B(n42561), .Z(n42535) );
  XOR U42233 ( .A(n42562), .B(n42563), .Z(n42538) );
  AND U42234 ( .A(n42564), .B(n42565), .Z(n42563) );
  XOR U42235 ( .A(n42562), .B(n42566), .Z(n42564) );
  XNOR U42236 ( .A(n42499), .B(n42544), .Z(n42546) );
  XNOR U42237 ( .A(n42567), .B(n42568), .Z(n42499) );
  AND U42238 ( .A(n1215), .B(n42569), .Z(n42568) );
  XNOR U42239 ( .A(n42570), .B(n42571), .Z(n42569) );
  XOR U42240 ( .A(n42572), .B(n42573), .Z(n42544) );
  AND U42241 ( .A(n42574), .B(n42575), .Z(n42573) );
  XNOR U42242 ( .A(n42572), .B(n42560), .Z(n42575) );
  IV U42243 ( .A(n42510), .Z(n42560) );
  XNOR U42244 ( .A(n42576), .B(n42553), .Z(n42510) );
  XNOR U42245 ( .A(n42577), .B(n42559), .Z(n42553) );
  XOR U42246 ( .A(n42578), .B(n42579), .Z(n42559) );
  NOR U42247 ( .A(n42580), .B(n42581), .Z(n42579) );
  XNOR U42248 ( .A(n42578), .B(n42582), .Z(n42580) );
  XNOR U42249 ( .A(n42558), .B(n42550), .Z(n42577) );
  XOR U42250 ( .A(n42583), .B(n42584), .Z(n42550) );
  AND U42251 ( .A(n42585), .B(n42586), .Z(n42584) );
  XNOR U42252 ( .A(n42583), .B(n42587), .Z(n42585) );
  XNOR U42253 ( .A(n42588), .B(n42555), .Z(n42558) );
  XOR U42254 ( .A(n42589), .B(n42590), .Z(n42555) );
  AND U42255 ( .A(n42591), .B(n42592), .Z(n42590) );
  XOR U42256 ( .A(n42589), .B(n42593), .Z(n42591) );
  XNOR U42257 ( .A(n42594), .B(n42595), .Z(n42588) );
  NOR U42258 ( .A(n42596), .B(n42597), .Z(n42595) );
  XOR U42259 ( .A(n42594), .B(n42598), .Z(n42596) );
  XNOR U42260 ( .A(n42554), .B(n42561), .Z(n42576) );
  NOR U42261 ( .A(n42516), .B(n42599), .Z(n42561) );
  XOR U42262 ( .A(n42566), .B(n42565), .Z(n42554) );
  XNOR U42263 ( .A(n42600), .B(n42562), .Z(n42565) );
  XOR U42264 ( .A(n42601), .B(n42602), .Z(n42562) );
  AND U42265 ( .A(n42603), .B(n42604), .Z(n42602) );
  XOR U42266 ( .A(n42601), .B(n42605), .Z(n42603) );
  XNOR U42267 ( .A(n42606), .B(n42607), .Z(n42600) );
  NOR U42268 ( .A(n42608), .B(n42609), .Z(n42607) );
  XNOR U42269 ( .A(n42606), .B(n42610), .Z(n42608) );
  XOR U42270 ( .A(n42611), .B(n42612), .Z(n42566) );
  NOR U42271 ( .A(n42613), .B(n42614), .Z(n42612) );
  XNOR U42272 ( .A(n42611), .B(n42615), .Z(n42613) );
  XNOR U42273 ( .A(n42507), .B(n42572), .Z(n42574) );
  XNOR U42274 ( .A(n42616), .B(n42617), .Z(n42507) );
  AND U42275 ( .A(n1215), .B(n42618), .Z(n42617) );
  XNOR U42276 ( .A(n42619), .B(n42620), .Z(n42618) );
  AND U42277 ( .A(n42513), .B(n42516), .Z(n42572) );
  XOR U42278 ( .A(n42621), .B(n42599), .Z(n42516) );
  XNOR U42279 ( .A(p_input[2048]), .B(p_input[960]), .Z(n42599) );
  XOR U42280 ( .A(n42587), .B(n42586), .Z(n42621) );
  XNOR U42281 ( .A(n42622), .B(n42593), .Z(n42586) );
  XNOR U42282 ( .A(n42582), .B(n42581), .Z(n42593) );
  XOR U42283 ( .A(n42623), .B(n42578), .Z(n42581) );
  XNOR U42284 ( .A(n29266), .B(p_input[970]), .Z(n42578) );
  XNOR U42285 ( .A(p_input[2059]), .B(p_input[971]), .Z(n42623) );
  XOR U42286 ( .A(p_input[2060]), .B(p_input[972]), .Z(n42582) );
  XNOR U42287 ( .A(n42592), .B(n42583), .Z(n42622) );
  XNOR U42288 ( .A(n29494), .B(p_input[961]), .Z(n42583) );
  XOR U42289 ( .A(n42624), .B(n42598), .Z(n42592) );
  XNOR U42290 ( .A(p_input[2063]), .B(p_input[975]), .Z(n42598) );
  XOR U42291 ( .A(n42589), .B(n42597), .Z(n42624) );
  XOR U42292 ( .A(n42625), .B(n42594), .Z(n42597) );
  XOR U42293 ( .A(p_input[2061]), .B(p_input[973]), .Z(n42594) );
  XNOR U42294 ( .A(p_input[2062]), .B(p_input[974]), .Z(n42625) );
  XNOR U42295 ( .A(n29036), .B(p_input[969]), .Z(n42589) );
  XNOR U42296 ( .A(n42605), .B(n42604), .Z(n42587) );
  XNOR U42297 ( .A(n42626), .B(n42610), .Z(n42604) );
  XOR U42298 ( .A(p_input[2056]), .B(p_input[968]), .Z(n42610) );
  XOR U42299 ( .A(n42601), .B(n42609), .Z(n42626) );
  XOR U42300 ( .A(n42627), .B(n42606), .Z(n42609) );
  XOR U42301 ( .A(p_input[2054]), .B(p_input[966]), .Z(n42606) );
  XNOR U42302 ( .A(p_input[2055]), .B(p_input[967]), .Z(n42627) );
  XNOR U42303 ( .A(n29039), .B(p_input[962]), .Z(n42601) );
  XNOR U42304 ( .A(n42615), .B(n42614), .Z(n42605) );
  XOR U42305 ( .A(n42628), .B(n42611), .Z(n42614) );
  XOR U42306 ( .A(p_input[2051]), .B(p_input[963]), .Z(n42611) );
  XNOR U42307 ( .A(p_input[2052]), .B(p_input[964]), .Z(n42628) );
  XOR U42308 ( .A(p_input[2053]), .B(p_input[965]), .Z(n42615) );
  XNOR U42309 ( .A(n42629), .B(n42630), .Z(n42513) );
  AND U42310 ( .A(n1215), .B(n42631), .Z(n42630) );
  XNOR U42311 ( .A(n42632), .B(n42633), .Z(n1215) );
  AND U42312 ( .A(n42634), .B(n42635), .Z(n42633) );
  XOR U42313 ( .A(n42527), .B(n42632), .Z(n42635) );
  XNOR U42314 ( .A(n42636), .B(n42632), .Z(n42634) );
  XOR U42315 ( .A(n42637), .B(n42638), .Z(n42632) );
  AND U42316 ( .A(n42639), .B(n42640), .Z(n42638) );
  XOR U42317 ( .A(n42542), .B(n42637), .Z(n42640) );
  XOR U42318 ( .A(n42637), .B(n42543), .Z(n42639) );
  XOR U42319 ( .A(n42641), .B(n42642), .Z(n42637) );
  AND U42320 ( .A(n42643), .B(n42644), .Z(n42642) );
  XOR U42321 ( .A(n42570), .B(n42641), .Z(n42644) );
  XOR U42322 ( .A(n42641), .B(n42571), .Z(n42643) );
  XOR U42323 ( .A(n42645), .B(n42646), .Z(n42641) );
  AND U42324 ( .A(n42647), .B(n42648), .Z(n42646) );
  XOR U42325 ( .A(n42645), .B(n42619), .Z(n42648) );
  XNOR U42326 ( .A(n42649), .B(n42650), .Z(n42473) );
  AND U42327 ( .A(n1219), .B(n42651), .Z(n42650) );
  XNOR U42328 ( .A(n42652), .B(n42653), .Z(n1219) );
  AND U42329 ( .A(n42654), .B(n42655), .Z(n42653) );
  XOR U42330 ( .A(n42652), .B(n42483), .Z(n42655) );
  XNOR U42331 ( .A(n42652), .B(n42443), .Z(n42654) );
  XOR U42332 ( .A(n42656), .B(n42657), .Z(n42652) );
  AND U42333 ( .A(n42658), .B(n42659), .Z(n42657) );
  XOR U42334 ( .A(n42656), .B(n42451), .Z(n42658) );
  XOR U42335 ( .A(n42660), .B(n42661), .Z(n42434) );
  AND U42336 ( .A(n1223), .B(n42651), .Z(n42661) );
  XNOR U42337 ( .A(n42649), .B(n42660), .Z(n42651) );
  XNOR U42338 ( .A(n42662), .B(n42663), .Z(n1223) );
  AND U42339 ( .A(n42664), .B(n42665), .Z(n42663) );
  XNOR U42340 ( .A(n42666), .B(n42662), .Z(n42665) );
  IV U42341 ( .A(n42483), .Z(n42666) );
  XOR U42342 ( .A(n42636), .B(n42667), .Z(n42483) );
  AND U42343 ( .A(n1226), .B(n42668), .Z(n42667) );
  XOR U42344 ( .A(n42526), .B(n42523), .Z(n42668) );
  IV U42345 ( .A(n42636), .Z(n42526) );
  XNOR U42346 ( .A(n42443), .B(n42662), .Z(n42664) );
  XOR U42347 ( .A(n42669), .B(n42670), .Z(n42443) );
  AND U42348 ( .A(n1242), .B(n42671), .Z(n42670) );
  XOR U42349 ( .A(n42656), .B(n42672), .Z(n42662) );
  AND U42350 ( .A(n42673), .B(n42659), .Z(n42672) );
  XNOR U42351 ( .A(n42493), .B(n42656), .Z(n42659) );
  XOR U42352 ( .A(n42543), .B(n42674), .Z(n42493) );
  AND U42353 ( .A(n1226), .B(n42675), .Z(n42674) );
  XOR U42354 ( .A(n42539), .B(n42543), .Z(n42675) );
  XNOR U42355 ( .A(n42676), .B(n42656), .Z(n42673) );
  IV U42356 ( .A(n42451), .Z(n42676) );
  XOR U42357 ( .A(n42677), .B(n42678), .Z(n42451) );
  AND U42358 ( .A(n1242), .B(n42679), .Z(n42678) );
  XOR U42359 ( .A(n42680), .B(n42681), .Z(n42656) );
  AND U42360 ( .A(n42682), .B(n42683), .Z(n42681) );
  XNOR U42361 ( .A(n42503), .B(n42680), .Z(n42683) );
  XOR U42362 ( .A(n42571), .B(n42684), .Z(n42503) );
  AND U42363 ( .A(n1226), .B(n42685), .Z(n42684) );
  XOR U42364 ( .A(n42567), .B(n42571), .Z(n42685) );
  XOR U42365 ( .A(n42680), .B(n42460), .Z(n42682) );
  XOR U42366 ( .A(n42686), .B(n42687), .Z(n42460) );
  AND U42367 ( .A(n1242), .B(n42688), .Z(n42687) );
  XOR U42368 ( .A(n42689), .B(n42690), .Z(n42680) );
  AND U42369 ( .A(n42691), .B(n42692), .Z(n42690) );
  XNOR U42370 ( .A(n42689), .B(n42511), .Z(n42692) );
  XOR U42371 ( .A(n42620), .B(n42693), .Z(n42511) );
  AND U42372 ( .A(n1226), .B(n42694), .Z(n42693) );
  XOR U42373 ( .A(n42616), .B(n42620), .Z(n42694) );
  XNOR U42374 ( .A(n42695), .B(n42689), .Z(n42691) );
  IV U42375 ( .A(n42470), .Z(n42695) );
  XOR U42376 ( .A(n42696), .B(n42697), .Z(n42470) );
  AND U42377 ( .A(n1242), .B(n42698), .Z(n42697) );
  AND U42378 ( .A(n42660), .B(n42649), .Z(n42689) );
  XNOR U42379 ( .A(n42699), .B(n42700), .Z(n42649) );
  AND U42380 ( .A(n1226), .B(n42631), .Z(n42700) );
  XNOR U42381 ( .A(n42629), .B(n42699), .Z(n42631) );
  XNOR U42382 ( .A(n42701), .B(n42702), .Z(n1226) );
  AND U42383 ( .A(n42703), .B(n42704), .Z(n42702) );
  XNOR U42384 ( .A(n42701), .B(n42523), .Z(n42704) );
  IV U42385 ( .A(n42527), .Z(n42523) );
  XOR U42386 ( .A(n42705), .B(n42706), .Z(n42527) );
  AND U42387 ( .A(n1230), .B(n42707), .Z(n42706) );
  XOR U42388 ( .A(n42708), .B(n42705), .Z(n42707) );
  XNOR U42389 ( .A(n42701), .B(n42636), .Z(n42703) );
  XOR U42390 ( .A(n42709), .B(n42710), .Z(n42636) );
  AND U42391 ( .A(n1238), .B(n42671), .Z(n42710) );
  XOR U42392 ( .A(n42669), .B(n42709), .Z(n42671) );
  XOR U42393 ( .A(n42711), .B(n42712), .Z(n42701) );
  AND U42394 ( .A(n42713), .B(n42714), .Z(n42712) );
  XNOR U42395 ( .A(n42711), .B(n42539), .Z(n42714) );
  IV U42396 ( .A(n42542), .Z(n42539) );
  XOR U42397 ( .A(n42715), .B(n42716), .Z(n42542) );
  AND U42398 ( .A(n1230), .B(n42717), .Z(n42716) );
  XOR U42399 ( .A(n42718), .B(n42715), .Z(n42717) );
  XOR U42400 ( .A(n42543), .B(n42711), .Z(n42713) );
  XOR U42401 ( .A(n42719), .B(n42720), .Z(n42543) );
  AND U42402 ( .A(n1238), .B(n42679), .Z(n42720) );
  XOR U42403 ( .A(n42719), .B(n42677), .Z(n42679) );
  XOR U42404 ( .A(n42721), .B(n42722), .Z(n42711) );
  AND U42405 ( .A(n42723), .B(n42724), .Z(n42722) );
  XNOR U42406 ( .A(n42721), .B(n42567), .Z(n42724) );
  IV U42407 ( .A(n42570), .Z(n42567) );
  XOR U42408 ( .A(n42725), .B(n42726), .Z(n42570) );
  AND U42409 ( .A(n1230), .B(n42727), .Z(n42726) );
  XNOR U42410 ( .A(n42728), .B(n42725), .Z(n42727) );
  XOR U42411 ( .A(n42571), .B(n42721), .Z(n42723) );
  XOR U42412 ( .A(n42729), .B(n42730), .Z(n42571) );
  AND U42413 ( .A(n1238), .B(n42688), .Z(n42730) );
  XOR U42414 ( .A(n42729), .B(n42686), .Z(n42688) );
  XOR U42415 ( .A(n42645), .B(n42731), .Z(n42721) );
  AND U42416 ( .A(n42647), .B(n42732), .Z(n42731) );
  XNOR U42417 ( .A(n42645), .B(n42616), .Z(n42732) );
  IV U42418 ( .A(n42619), .Z(n42616) );
  XOR U42419 ( .A(n42733), .B(n42734), .Z(n42619) );
  AND U42420 ( .A(n1230), .B(n42735), .Z(n42734) );
  XOR U42421 ( .A(n42736), .B(n42733), .Z(n42735) );
  XOR U42422 ( .A(n42620), .B(n42645), .Z(n42647) );
  XOR U42423 ( .A(n42737), .B(n42738), .Z(n42620) );
  AND U42424 ( .A(n1238), .B(n42698), .Z(n42738) );
  XOR U42425 ( .A(n42737), .B(n42696), .Z(n42698) );
  AND U42426 ( .A(n42699), .B(n42629), .Z(n42645) );
  XNOR U42427 ( .A(n42739), .B(n42740), .Z(n42629) );
  AND U42428 ( .A(n1230), .B(n42741), .Z(n42740) );
  XNOR U42429 ( .A(n42742), .B(n42739), .Z(n42741) );
  XNOR U42430 ( .A(n42743), .B(n42744), .Z(n1230) );
  AND U42431 ( .A(n42745), .B(n42746), .Z(n42744) );
  XOR U42432 ( .A(n42708), .B(n42743), .Z(n42746) );
  AND U42433 ( .A(n42747), .B(n42748), .Z(n42708) );
  XNOR U42434 ( .A(n42705), .B(n42743), .Z(n42745) );
  XNOR U42435 ( .A(n42749), .B(n42750), .Z(n42705) );
  AND U42436 ( .A(n1234), .B(n42751), .Z(n42750) );
  XNOR U42437 ( .A(n42752), .B(n42753), .Z(n42751) );
  XOR U42438 ( .A(n42754), .B(n42755), .Z(n42743) );
  AND U42439 ( .A(n42756), .B(n42757), .Z(n42755) );
  XNOR U42440 ( .A(n42754), .B(n42747), .Z(n42757) );
  IV U42441 ( .A(n42718), .Z(n42747) );
  XOR U42442 ( .A(n42758), .B(n42759), .Z(n42718) );
  XOR U42443 ( .A(n42760), .B(n42748), .Z(n42759) );
  AND U42444 ( .A(n42728), .B(n42761), .Z(n42748) );
  AND U42445 ( .A(n42762), .B(n42763), .Z(n42760) );
  XOR U42446 ( .A(n42764), .B(n42758), .Z(n42762) );
  XNOR U42447 ( .A(n42715), .B(n42754), .Z(n42756) );
  XNOR U42448 ( .A(n42765), .B(n42766), .Z(n42715) );
  AND U42449 ( .A(n1234), .B(n42767), .Z(n42766) );
  XNOR U42450 ( .A(n42768), .B(n42769), .Z(n42767) );
  XOR U42451 ( .A(n42770), .B(n42771), .Z(n42754) );
  AND U42452 ( .A(n42772), .B(n42773), .Z(n42771) );
  XNOR U42453 ( .A(n42770), .B(n42728), .Z(n42773) );
  XOR U42454 ( .A(n42774), .B(n42763), .Z(n42728) );
  XNOR U42455 ( .A(n42775), .B(n42758), .Z(n42763) );
  XOR U42456 ( .A(n42776), .B(n42777), .Z(n42758) );
  AND U42457 ( .A(n42778), .B(n42779), .Z(n42777) );
  XOR U42458 ( .A(n42780), .B(n42776), .Z(n42778) );
  XNOR U42459 ( .A(n42781), .B(n42782), .Z(n42775) );
  AND U42460 ( .A(n42783), .B(n42784), .Z(n42782) );
  XOR U42461 ( .A(n42781), .B(n42785), .Z(n42783) );
  XNOR U42462 ( .A(n42764), .B(n42761), .Z(n42774) );
  AND U42463 ( .A(n42786), .B(n42787), .Z(n42761) );
  XOR U42464 ( .A(n42788), .B(n42789), .Z(n42764) );
  AND U42465 ( .A(n42790), .B(n42791), .Z(n42789) );
  XOR U42466 ( .A(n42788), .B(n42792), .Z(n42790) );
  XNOR U42467 ( .A(n42725), .B(n42770), .Z(n42772) );
  XNOR U42468 ( .A(n42793), .B(n42794), .Z(n42725) );
  AND U42469 ( .A(n1234), .B(n42795), .Z(n42794) );
  XNOR U42470 ( .A(n42796), .B(n42797), .Z(n42795) );
  XOR U42471 ( .A(n42798), .B(n42799), .Z(n42770) );
  AND U42472 ( .A(n42800), .B(n42801), .Z(n42799) );
  XNOR U42473 ( .A(n42798), .B(n42786), .Z(n42801) );
  IV U42474 ( .A(n42736), .Z(n42786) );
  XNOR U42475 ( .A(n42802), .B(n42779), .Z(n42736) );
  XNOR U42476 ( .A(n42803), .B(n42785), .Z(n42779) );
  XOR U42477 ( .A(n42804), .B(n42805), .Z(n42785) );
  NOR U42478 ( .A(n42806), .B(n42807), .Z(n42805) );
  XNOR U42479 ( .A(n42804), .B(n42808), .Z(n42806) );
  XNOR U42480 ( .A(n42784), .B(n42776), .Z(n42803) );
  XOR U42481 ( .A(n42809), .B(n42810), .Z(n42776) );
  AND U42482 ( .A(n42811), .B(n42812), .Z(n42810) );
  XNOR U42483 ( .A(n42809), .B(n42813), .Z(n42811) );
  XNOR U42484 ( .A(n42814), .B(n42781), .Z(n42784) );
  XOR U42485 ( .A(n42815), .B(n42816), .Z(n42781) );
  AND U42486 ( .A(n42817), .B(n42818), .Z(n42816) );
  XOR U42487 ( .A(n42815), .B(n42819), .Z(n42817) );
  XNOR U42488 ( .A(n42820), .B(n42821), .Z(n42814) );
  NOR U42489 ( .A(n42822), .B(n42823), .Z(n42821) );
  XOR U42490 ( .A(n42820), .B(n42824), .Z(n42822) );
  XNOR U42491 ( .A(n42780), .B(n42787), .Z(n42802) );
  NOR U42492 ( .A(n42742), .B(n42825), .Z(n42787) );
  XOR U42493 ( .A(n42792), .B(n42791), .Z(n42780) );
  XNOR U42494 ( .A(n42826), .B(n42788), .Z(n42791) );
  XOR U42495 ( .A(n42827), .B(n42828), .Z(n42788) );
  AND U42496 ( .A(n42829), .B(n42830), .Z(n42828) );
  XOR U42497 ( .A(n42827), .B(n42831), .Z(n42829) );
  XNOR U42498 ( .A(n42832), .B(n42833), .Z(n42826) );
  NOR U42499 ( .A(n42834), .B(n42835), .Z(n42833) );
  XNOR U42500 ( .A(n42832), .B(n42836), .Z(n42834) );
  XOR U42501 ( .A(n42837), .B(n42838), .Z(n42792) );
  NOR U42502 ( .A(n42839), .B(n42840), .Z(n42838) );
  XNOR U42503 ( .A(n42837), .B(n42841), .Z(n42839) );
  XNOR U42504 ( .A(n42733), .B(n42798), .Z(n42800) );
  XNOR U42505 ( .A(n42842), .B(n42843), .Z(n42733) );
  AND U42506 ( .A(n1234), .B(n42844), .Z(n42843) );
  XNOR U42507 ( .A(n42845), .B(n42846), .Z(n42844) );
  AND U42508 ( .A(n42739), .B(n42742), .Z(n42798) );
  XOR U42509 ( .A(n42847), .B(n42825), .Z(n42742) );
  XNOR U42510 ( .A(p_input[2048]), .B(p_input[976]), .Z(n42825) );
  XOR U42511 ( .A(n42813), .B(n42812), .Z(n42847) );
  XNOR U42512 ( .A(n42848), .B(n42819), .Z(n42812) );
  XNOR U42513 ( .A(n42808), .B(n42807), .Z(n42819) );
  XOR U42514 ( .A(n42849), .B(n42804), .Z(n42807) );
  XNOR U42515 ( .A(n29266), .B(p_input[986]), .Z(n42804) );
  XNOR U42516 ( .A(p_input[2059]), .B(p_input[987]), .Z(n42849) );
  XOR U42517 ( .A(p_input[2060]), .B(p_input[988]), .Z(n42808) );
  XNOR U42518 ( .A(n42818), .B(n42809), .Z(n42848) );
  XNOR U42519 ( .A(n29494), .B(p_input[977]), .Z(n42809) );
  XOR U42520 ( .A(n42850), .B(n42824), .Z(n42818) );
  XNOR U42521 ( .A(p_input[2063]), .B(p_input[991]), .Z(n42824) );
  XOR U42522 ( .A(n42815), .B(n42823), .Z(n42850) );
  XOR U42523 ( .A(n42851), .B(n42820), .Z(n42823) );
  XOR U42524 ( .A(p_input[2061]), .B(p_input[989]), .Z(n42820) );
  XNOR U42525 ( .A(p_input[2062]), .B(p_input[990]), .Z(n42851) );
  XNOR U42526 ( .A(n29036), .B(p_input[985]), .Z(n42815) );
  XNOR U42527 ( .A(n42831), .B(n42830), .Z(n42813) );
  XNOR U42528 ( .A(n42852), .B(n42836), .Z(n42830) );
  XOR U42529 ( .A(p_input[2056]), .B(p_input[984]), .Z(n42836) );
  XOR U42530 ( .A(n42827), .B(n42835), .Z(n42852) );
  XOR U42531 ( .A(n42853), .B(n42832), .Z(n42835) );
  XOR U42532 ( .A(p_input[2054]), .B(p_input[982]), .Z(n42832) );
  XNOR U42533 ( .A(p_input[2055]), .B(p_input[983]), .Z(n42853) );
  XNOR U42534 ( .A(n29039), .B(p_input[978]), .Z(n42827) );
  XNOR U42535 ( .A(n42841), .B(n42840), .Z(n42831) );
  XOR U42536 ( .A(n42854), .B(n42837), .Z(n42840) );
  XOR U42537 ( .A(p_input[2051]), .B(p_input[979]), .Z(n42837) );
  XNOR U42538 ( .A(p_input[2052]), .B(p_input[980]), .Z(n42854) );
  XOR U42539 ( .A(p_input[2053]), .B(p_input[981]), .Z(n42841) );
  XNOR U42540 ( .A(n42855), .B(n42856), .Z(n42739) );
  AND U42541 ( .A(n1234), .B(n42857), .Z(n42856) );
  XNOR U42542 ( .A(n42858), .B(n42859), .Z(n1234) );
  AND U42543 ( .A(n42860), .B(n42861), .Z(n42859) );
  XOR U42544 ( .A(n42753), .B(n42858), .Z(n42861) );
  XNOR U42545 ( .A(n42862), .B(n42858), .Z(n42860) );
  XOR U42546 ( .A(n42863), .B(n42864), .Z(n42858) );
  AND U42547 ( .A(n42865), .B(n42866), .Z(n42864) );
  XOR U42548 ( .A(n42768), .B(n42863), .Z(n42866) );
  XOR U42549 ( .A(n42863), .B(n42769), .Z(n42865) );
  XOR U42550 ( .A(n42867), .B(n42868), .Z(n42863) );
  AND U42551 ( .A(n42869), .B(n42870), .Z(n42868) );
  XOR U42552 ( .A(n42796), .B(n42867), .Z(n42870) );
  XOR U42553 ( .A(n42867), .B(n42797), .Z(n42869) );
  XOR U42554 ( .A(n42871), .B(n42872), .Z(n42867) );
  AND U42555 ( .A(n42873), .B(n42874), .Z(n42872) );
  XOR U42556 ( .A(n42871), .B(n42845), .Z(n42874) );
  XNOR U42557 ( .A(n42875), .B(n42876), .Z(n42699) );
  AND U42558 ( .A(n1238), .B(n42877), .Z(n42876) );
  XNOR U42559 ( .A(n42878), .B(n42879), .Z(n1238) );
  AND U42560 ( .A(n42880), .B(n42881), .Z(n42879) );
  XOR U42561 ( .A(n42878), .B(n42709), .Z(n42881) );
  XNOR U42562 ( .A(n42878), .B(n42669), .Z(n42880) );
  XOR U42563 ( .A(n42882), .B(n42883), .Z(n42878) );
  AND U42564 ( .A(n42884), .B(n42885), .Z(n42883) );
  XOR U42565 ( .A(n42882), .B(n42677), .Z(n42884) );
  XOR U42566 ( .A(n42886), .B(n42887), .Z(n42660) );
  AND U42567 ( .A(n1242), .B(n42877), .Z(n42887) );
  XNOR U42568 ( .A(n42875), .B(n42886), .Z(n42877) );
  XNOR U42569 ( .A(n42888), .B(n42889), .Z(n1242) );
  AND U42570 ( .A(n42890), .B(n42891), .Z(n42889) );
  XNOR U42571 ( .A(n42892), .B(n42888), .Z(n42891) );
  IV U42572 ( .A(n42709), .Z(n42892) );
  XOR U42573 ( .A(n42862), .B(n42893), .Z(n42709) );
  AND U42574 ( .A(n1245), .B(n42894), .Z(n42893) );
  XOR U42575 ( .A(n42752), .B(n42749), .Z(n42894) );
  IV U42576 ( .A(n42862), .Z(n42752) );
  XNOR U42577 ( .A(n42669), .B(n42888), .Z(n42890) );
  XOR U42578 ( .A(n42895), .B(n42896), .Z(n42669) );
  AND U42579 ( .A(n1261), .B(n42897), .Z(n42896) );
  XOR U42580 ( .A(n42882), .B(n42898), .Z(n42888) );
  AND U42581 ( .A(n42899), .B(n42885), .Z(n42898) );
  XNOR U42582 ( .A(n42719), .B(n42882), .Z(n42885) );
  XOR U42583 ( .A(n42769), .B(n42900), .Z(n42719) );
  AND U42584 ( .A(n1245), .B(n42901), .Z(n42900) );
  XOR U42585 ( .A(n42765), .B(n42769), .Z(n42901) );
  XNOR U42586 ( .A(n42902), .B(n42882), .Z(n42899) );
  IV U42587 ( .A(n42677), .Z(n42902) );
  XOR U42588 ( .A(n42903), .B(n42904), .Z(n42677) );
  AND U42589 ( .A(n1261), .B(n42905), .Z(n42904) );
  XOR U42590 ( .A(n42906), .B(n42907), .Z(n42882) );
  AND U42591 ( .A(n42908), .B(n42909), .Z(n42907) );
  XNOR U42592 ( .A(n42729), .B(n42906), .Z(n42909) );
  XOR U42593 ( .A(n42797), .B(n42910), .Z(n42729) );
  AND U42594 ( .A(n1245), .B(n42911), .Z(n42910) );
  XOR U42595 ( .A(n42793), .B(n42797), .Z(n42911) );
  XOR U42596 ( .A(n42906), .B(n42686), .Z(n42908) );
  XOR U42597 ( .A(n42912), .B(n42913), .Z(n42686) );
  AND U42598 ( .A(n1261), .B(n42914), .Z(n42913) );
  XOR U42599 ( .A(n42915), .B(n42916), .Z(n42906) );
  AND U42600 ( .A(n42917), .B(n42918), .Z(n42916) );
  XNOR U42601 ( .A(n42915), .B(n42737), .Z(n42918) );
  XOR U42602 ( .A(n42846), .B(n42919), .Z(n42737) );
  AND U42603 ( .A(n1245), .B(n42920), .Z(n42919) );
  XOR U42604 ( .A(n42842), .B(n42846), .Z(n42920) );
  XNOR U42605 ( .A(n42921), .B(n42915), .Z(n42917) );
  IV U42606 ( .A(n42696), .Z(n42921) );
  XOR U42607 ( .A(n42922), .B(n42923), .Z(n42696) );
  AND U42608 ( .A(n1261), .B(n42924), .Z(n42923) );
  AND U42609 ( .A(n42886), .B(n42875), .Z(n42915) );
  XNOR U42610 ( .A(n42925), .B(n42926), .Z(n42875) );
  AND U42611 ( .A(n1245), .B(n42857), .Z(n42926) );
  XNOR U42612 ( .A(n42855), .B(n42925), .Z(n42857) );
  XNOR U42613 ( .A(n42927), .B(n42928), .Z(n1245) );
  AND U42614 ( .A(n42929), .B(n42930), .Z(n42928) );
  XNOR U42615 ( .A(n42927), .B(n42749), .Z(n42930) );
  IV U42616 ( .A(n42753), .Z(n42749) );
  XOR U42617 ( .A(n42931), .B(n42932), .Z(n42753) );
  AND U42618 ( .A(n1249), .B(n42933), .Z(n42932) );
  XOR U42619 ( .A(n42934), .B(n42931), .Z(n42933) );
  XNOR U42620 ( .A(n42927), .B(n42862), .Z(n42929) );
  XOR U42621 ( .A(n42935), .B(n42936), .Z(n42862) );
  AND U42622 ( .A(n1257), .B(n42897), .Z(n42936) );
  XOR U42623 ( .A(n42895), .B(n42935), .Z(n42897) );
  XOR U42624 ( .A(n42937), .B(n42938), .Z(n42927) );
  AND U42625 ( .A(n42939), .B(n42940), .Z(n42938) );
  XNOR U42626 ( .A(n42937), .B(n42765), .Z(n42940) );
  IV U42627 ( .A(n42768), .Z(n42765) );
  XOR U42628 ( .A(n42941), .B(n42942), .Z(n42768) );
  AND U42629 ( .A(n1249), .B(n42943), .Z(n42942) );
  XOR U42630 ( .A(n42944), .B(n42941), .Z(n42943) );
  XOR U42631 ( .A(n42769), .B(n42937), .Z(n42939) );
  XOR U42632 ( .A(n42945), .B(n42946), .Z(n42769) );
  AND U42633 ( .A(n1257), .B(n42905), .Z(n42946) );
  XOR U42634 ( .A(n42945), .B(n42903), .Z(n42905) );
  XOR U42635 ( .A(n42947), .B(n42948), .Z(n42937) );
  AND U42636 ( .A(n42949), .B(n42950), .Z(n42948) );
  XNOR U42637 ( .A(n42947), .B(n42793), .Z(n42950) );
  IV U42638 ( .A(n42796), .Z(n42793) );
  XOR U42639 ( .A(n42951), .B(n42952), .Z(n42796) );
  AND U42640 ( .A(n1249), .B(n42953), .Z(n42952) );
  XNOR U42641 ( .A(n42954), .B(n42951), .Z(n42953) );
  XOR U42642 ( .A(n42797), .B(n42947), .Z(n42949) );
  XOR U42643 ( .A(n42955), .B(n42956), .Z(n42797) );
  AND U42644 ( .A(n1257), .B(n42914), .Z(n42956) );
  XOR U42645 ( .A(n42955), .B(n42912), .Z(n42914) );
  XOR U42646 ( .A(n42871), .B(n42957), .Z(n42947) );
  AND U42647 ( .A(n42873), .B(n42958), .Z(n42957) );
  XNOR U42648 ( .A(n42871), .B(n42842), .Z(n42958) );
  IV U42649 ( .A(n42845), .Z(n42842) );
  XOR U42650 ( .A(n42959), .B(n42960), .Z(n42845) );
  AND U42651 ( .A(n1249), .B(n42961), .Z(n42960) );
  XOR U42652 ( .A(n42962), .B(n42959), .Z(n42961) );
  XOR U42653 ( .A(n42846), .B(n42871), .Z(n42873) );
  XOR U42654 ( .A(n42963), .B(n42964), .Z(n42846) );
  AND U42655 ( .A(n1257), .B(n42924), .Z(n42964) );
  XOR U42656 ( .A(n42963), .B(n42922), .Z(n42924) );
  AND U42657 ( .A(n42925), .B(n42855), .Z(n42871) );
  XNOR U42658 ( .A(n42965), .B(n42966), .Z(n42855) );
  AND U42659 ( .A(n1249), .B(n42967), .Z(n42966) );
  XNOR U42660 ( .A(n42968), .B(n42965), .Z(n42967) );
  XNOR U42661 ( .A(n42969), .B(n42970), .Z(n1249) );
  AND U42662 ( .A(n42971), .B(n42972), .Z(n42970) );
  XOR U42663 ( .A(n42934), .B(n42969), .Z(n42972) );
  AND U42664 ( .A(n42973), .B(n42974), .Z(n42934) );
  XNOR U42665 ( .A(n42931), .B(n42969), .Z(n42971) );
  XNOR U42666 ( .A(n42975), .B(n42976), .Z(n42931) );
  AND U42667 ( .A(n1253), .B(n42977), .Z(n42976) );
  XNOR U42668 ( .A(n42978), .B(n42979), .Z(n42977) );
  XOR U42669 ( .A(n42980), .B(n42981), .Z(n42969) );
  AND U42670 ( .A(n42982), .B(n42983), .Z(n42981) );
  XNOR U42671 ( .A(n42980), .B(n42973), .Z(n42983) );
  IV U42672 ( .A(n42944), .Z(n42973) );
  XOR U42673 ( .A(n42984), .B(n42985), .Z(n42944) );
  XOR U42674 ( .A(n42986), .B(n42974), .Z(n42985) );
  AND U42675 ( .A(n42954), .B(n42987), .Z(n42974) );
  AND U42676 ( .A(n42988), .B(n42989), .Z(n42986) );
  XOR U42677 ( .A(n42990), .B(n42984), .Z(n42988) );
  XNOR U42678 ( .A(n42941), .B(n42980), .Z(n42982) );
  XNOR U42679 ( .A(n42991), .B(n42992), .Z(n42941) );
  AND U42680 ( .A(n1253), .B(n42993), .Z(n42992) );
  XNOR U42681 ( .A(n42994), .B(n42995), .Z(n42993) );
  XOR U42682 ( .A(n42996), .B(n42997), .Z(n42980) );
  AND U42683 ( .A(n42998), .B(n42999), .Z(n42997) );
  XNOR U42684 ( .A(n42996), .B(n42954), .Z(n42999) );
  XOR U42685 ( .A(n43000), .B(n42989), .Z(n42954) );
  XNOR U42686 ( .A(n43001), .B(n42984), .Z(n42989) );
  XOR U42687 ( .A(n43002), .B(n43003), .Z(n42984) );
  AND U42688 ( .A(n43004), .B(n43005), .Z(n43003) );
  XOR U42689 ( .A(n43006), .B(n43002), .Z(n43004) );
  XNOR U42690 ( .A(n43007), .B(n43008), .Z(n43001) );
  AND U42691 ( .A(n43009), .B(n43010), .Z(n43008) );
  XOR U42692 ( .A(n43007), .B(n43011), .Z(n43009) );
  XNOR U42693 ( .A(n42990), .B(n42987), .Z(n43000) );
  AND U42694 ( .A(n43012), .B(n43013), .Z(n42987) );
  XOR U42695 ( .A(n43014), .B(n43015), .Z(n42990) );
  AND U42696 ( .A(n43016), .B(n43017), .Z(n43015) );
  XOR U42697 ( .A(n43014), .B(n43018), .Z(n43016) );
  XNOR U42698 ( .A(n42951), .B(n42996), .Z(n42998) );
  XNOR U42699 ( .A(n43019), .B(n43020), .Z(n42951) );
  AND U42700 ( .A(n1253), .B(n43021), .Z(n43020) );
  XNOR U42701 ( .A(n43022), .B(n43023), .Z(n43021) );
  XOR U42702 ( .A(n43024), .B(n43025), .Z(n42996) );
  AND U42703 ( .A(n43026), .B(n43027), .Z(n43025) );
  XNOR U42704 ( .A(n43024), .B(n43012), .Z(n43027) );
  IV U42705 ( .A(n42962), .Z(n43012) );
  XNOR U42706 ( .A(n43028), .B(n43005), .Z(n42962) );
  XNOR U42707 ( .A(n43029), .B(n43011), .Z(n43005) );
  XNOR U42708 ( .A(n43030), .B(n43031), .Z(n43011) );
  NOR U42709 ( .A(n43032), .B(n43033), .Z(n43031) );
  XOR U42710 ( .A(n43030), .B(n43034), .Z(n43032) );
  XNOR U42711 ( .A(n43010), .B(n43002), .Z(n43029) );
  XOR U42712 ( .A(n43035), .B(n43036), .Z(n43002) );
  AND U42713 ( .A(n43037), .B(n43038), .Z(n43036) );
  XOR U42714 ( .A(n43035), .B(n43039), .Z(n43037) );
  XNOR U42715 ( .A(n43040), .B(n43007), .Z(n43010) );
  XOR U42716 ( .A(n43041), .B(n43042), .Z(n43007) );
  AND U42717 ( .A(n43043), .B(n43044), .Z(n43042) );
  XNOR U42718 ( .A(n43045), .B(n43046), .Z(n43043) );
  IV U42719 ( .A(n43041), .Z(n43045) );
  XNOR U42720 ( .A(n43047), .B(n43048), .Z(n43040) );
  NOR U42721 ( .A(n43049), .B(n43050), .Z(n43048) );
  XNOR U42722 ( .A(n43047), .B(n43051), .Z(n43049) );
  XNOR U42723 ( .A(n43006), .B(n43013), .Z(n43028) );
  NOR U42724 ( .A(n42968), .B(n43052), .Z(n43013) );
  XOR U42725 ( .A(n43018), .B(n43017), .Z(n43006) );
  XNOR U42726 ( .A(n43053), .B(n43014), .Z(n43017) );
  XOR U42727 ( .A(n43054), .B(n43055), .Z(n43014) );
  AND U42728 ( .A(n43056), .B(n43057), .Z(n43055) );
  XOR U42729 ( .A(n43054), .B(n43058), .Z(n43056) );
  XNOR U42730 ( .A(n43059), .B(n43060), .Z(n43053) );
  NOR U42731 ( .A(n43061), .B(n43062), .Z(n43060) );
  XNOR U42732 ( .A(n43059), .B(n43063), .Z(n43061) );
  XOR U42733 ( .A(n43064), .B(n43065), .Z(n43018) );
  NOR U42734 ( .A(n43066), .B(n43067), .Z(n43065) );
  XNOR U42735 ( .A(n43064), .B(n43068), .Z(n43066) );
  XNOR U42736 ( .A(n42959), .B(n43024), .Z(n43026) );
  XNOR U42737 ( .A(n43069), .B(n43070), .Z(n42959) );
  AND U42738 ( .A(n1253), .B(n43071), .Z(n43070) );
  XNOR U42739 ( .A(n43072), .B(n43073), .Z(n43071) );
  AND U42740 ( .A(n42965), .B(n42968), .Z(n43024) );
  XOR U42741 ( .A(n43074), .B(n43052), .Z(n42968) );
  XNOR U42742 ( .A(p_input[2048]), .B(p_input[992]), .Z(n43052) );
  XNOR U42743 ( .A(n43039), .B(n43038), .Z(n43074) );
  XNOR U42744 ( .A(n43075), .B(n43046), .Z(n43038) );
  XNOR U42745 ( .A(n43034), .B(n43033), .Z(n43046) );
  XNOR U42746 ( .A(n43076), .B(n43030), .Z(n43033) );
  XNOR U42747 ( .A(p_input[1002]), .B(p_input[2058]), .Z(n43030) );
  XOR U42748 ( .A(p_input[1003]), .B(n29030), .Z(n43076) );
  XOR U42749 ( .A(p_input[1004]), .B(p_input[2060]), .Z(n43034) );
  XNOR U42750 ( .A(n43044), .B(n43035), .Z(n43075) );
  XNOR U42751 ( .A(n29494), .B(p_input[993]), .Z(n43035) );
  XNOR U42752 ( .A(n43077), .B(n43051), .Z(n43044) );
  XNOR U42753 ( .A(p_input[1007]), .B(n29033), .Z(n43051) );
  XOR U42754 ( .A(n43041), .B(n43050), .Z(n43077) );
  XOR U42755 ( .A(n43078), .B(n43047), .Z(n43050) );
  XOR U42756 ( .A(p_input[1005]), .B(p_input[2061]), .Z(n43047) );
  XOR U42757 ( .A(p_input[1006]), .B(n29035), .Z(n43078) );
  XOR U42758 ( .A(p_input[1001]), .B(p_input[2057]), .Z(n43041) );
  XOR U42759 ( .A(n43058), .B(n43057), .Z(n43039) );
  XNOR U42760 ( .A(n43079), .B(n43063), .Z(n43057) );
  XOR U42761 ( .A(p_input[1000]), .B(p_input[2056]), .Z(n43063) );
  XOR U42762 ( .A(n43054), .B(n43062), .Z(n43079) );
  XOR U42763 ( .A(n43080), .B(n43059), .Z(n43062) );
  XOR U42764 ( .A(p_input[2054]), .B(p_input[998]), .Z(n43059) );
  XNOR U42765 ( .A(p_input[2055]), .B(p_input[999]), .Z(n43080) );
  XNOR U42766 ( .A(n29039), .B(p_input[994]), .Z(n43054) );
  XNOR U42767 ( .A(n43068), .B(n43067), .Z(n43058) );
  XOR U42768 ( .A(n43081), .B(n43064), .Z(n43067) );
  XOR U42769 ( .A(p_input[2051]), .B(p_input[995]), .Z(n43064) );
  XNOR U42770 ( .A(p_input[2052]), .B(p_input[996]), .Z(n43081) );
  XOR U42771 ( .A(p_input[2053]), .B(p_input[997]), .Z(n43068) );
  XNOR U42772 ( .A(n43082), .B(n43083), .Z(n42965) );
  AND U42773 ( .A(n1253), .B(n43084), .Z(n43083) );
  XNOR U42774 ( .A(n43085), .B(n43086), .Z(n1253) );
  AND U42775 ( .A(n43087), .B(n43088), .Z(n43086) );
  XOR U42776 ( .A(n42979), .B(n43085), .Z(n43088) );
  XNOR U42777 ( .A(n43089), .B(n43085), .Z(n43087) );
  XOR U42778 ( .A(n43090), .B(n43091), .Z(n43085) );
  AND U42779 ( .A(n43092), .B(n43093), .Z(n43091) );
  XOR U42780 ( .A(n42994), .B(n43090), .Z(n43093) );
  XOR U42781 ( .A(n43090), .B(n42995), .Z(n43092) );
  XOR U42782 ( .A(n43094), .B(n43095), .Z(n43090) );
  AND U42783 ( .A(n43096), .B(n43097), .Z(n43095) );
  XOR U42784 ( .A(n43022), .B(n43094), .Z(n43097) );
  XOR U42785 ( .A(n43094), .B(n43023), .Z(n43096) );
  XOR U42786 ( .A(n43098), .B(n43099), .Z(n43094) );
  AND U42787 ( .A(n43100), .B(n43101), .Z(n43099) );
  XOR U42788 ( .A(n43098), .B(n43072), .Z(n43101) );
  XNOR U42789 ( .A(n43102), .B(n43103), .Z(n42925) );
  AND U42790 ( .A(n1257), .B(n43104), .Z(n43103) );
  XNOR U42791 ( .A(n43105), .B(n43106), .Z(n1257) );
  AND U42792 ( .A(n43107), .B(n43108), .Z(n43106) );
  XOR U42793 ( .A(n43105), .B(n42935), .Z(n43108) );
  XNOR U42794 ( .A(n43105), .B(n42895), .Z(n43107) );
  XOR U42795 ( .A(n43109), .B(n43110), .Z(n43105) );
  AND U42796 ( .A(n43111), .B(n43112), .Z(n43110) );
  XOR U42797 ( .A(n43109), .B(n42903), .Z(n43111) );
  XOR U42798 ( .A(n43113), .B(n43114), .Z(n42886) );
  AND U42799 ( .A(n1261), .B(n43104), .Z(n43114) );
  XNOR U42800 ( .A(n43102), .B(n43113), .Z(n43104) );
  XNOR U42801 ( .A(n43115), .B(n43116), .Z(n1261) );
  AND U42802 ( .A(n43117), .B(n43118), .Z(n43116) );
  XNOR U42803 ( .A(n43119), .B(n43115), .Z(n43118) );
  IV U42804 ( .A(n42935), .Z(n43119) );
  XOR U42805 ( .A(n43089), .B(n43120), .Z(n42935) );
  AND U42806 ( .A(n1264), .B(n43121), .Z(n43120) );
  XOR U42807 ( .A(n42978), .B(n42975), .Z(n43121) );
  IV U42808 ( .A(n43089), .Z(n42978) );
  XNOR U42809 ( .A(n42895), .B(n43115), .Z(n43117) );
  XOR U42810 ( .A(n43122), .B(n43123), .Z(n42895) );
  AND U42811 ( .A(n1280), .B(n43124), .Z(n43123) );
  XOR U42812 ( .A(n43109), .B(n43125), .Z(n43115) );
  AND U42813 ( .A(n43126), .B(n43112), .Z(n43125) );
  XNOR U42814 ( .A(n42945), .B(n43109), .Z(n43112) );
  XOR U42815 ( .A(n42995), .B(n43127), .Z(n42945) );
  AND U42816 ( .A(n1264), .B(n43128), .Z(n43127) );
  XOR U42817 ( .A(n42991), .B(n42995), .Z(n43128) );
  XNOR U42818 ( .A(n43129), .B(n43109), .Z(n43126) );
  IV U42819 ( .A(n42903), .Z(n43129) );
  XOR U42820 ( .A(n43130), .B(n43131), .Z(n42903) );
  AND U42821 ( .A(n1280), .B(n43132), .Z(n43131) );
  XOR U42822 ( .A(n43133), .B(n43134), .Z(n43109) );
  AND U42823 ( .A(n43135), .B(n43136), .Z(n43134) );
  XNOR U42824 ( .A(n42955), .B(n43133), .Z(n43136) );
  XOR U42825 ( .A(n43023), .B(n43137), .Z(n42955) );
  AND U42826 ( .A(n1264), .B(n43138), .Z(n43137) );
  XOR U42827 ( .A(n43019), .B(n43023), .Z(n43138) );
  XOR U42828 ( .A(n43133), .B(n42912), .Z(n43135) );
  XOR U42829 ( .A(n43139), .B(n43140), .Z(n42912) );
  AND U42830 ( .A(n1280), .B(n43141), .Z(n43140) );
  XOR U42831 ( .A(n43142), .B(n43143), .Z(n43133) );
  AND U42832 ( .A(n43144), .B(n43145), .Z(n43143) );
  XNOR U42833 ( .A(n43142), .B(n42963), .Z(n43145) );
  XOR U42834 ( .A(n43073), .B(n43146), .Z(n42963) );
  AND U42835 ( .A(n1264), .B(n43147), .Z(n43146) );
  XOR U42836 ( .A(n43069), .B(n43073), .Z(n43147) );
  XNOR U42837 ( .A(n43148), .B(n43142), .Z(n43144) );
  IV U42838 ( .A(n42922), .Z(n43148) );
  XOR U42839 ( .A(n43149), .B(n43150), .Z(n42922) );
  AND U42840 ( .A(n1280), .B(n43151), .Z(n43150) );
  AND U42841 ( .A(n43113), .B(n43102), .Z(n43142) );
  XNOR U42842 ( .A(n43152), .B(n43153), .Z(n43102) );
  AND U42843 ( .A(n1264), .B(n43084), .Z(n43153) );
  XNOR U42844 ( .A(n43082), .B(n43152), .Z(n43084) );
  XNOR U42845 ( .A(n43154), .B(n43155), .Z(n1264) );
  AND U42846 ( .A(n43156), .B(n43157), .Z(n43155) );
  XNOR U42847 ( .A(n43154), .B(n42975), .Z(n43157) );
  IV U42848 ( .A(n42979), .Z(n42975) );
  XOR U42849 ( .A(n43158), .B(n43159), .Z(n42979) );
  AND U42850 ( .A(n1268), .B(n43160), .Z(n43159) );
  XOR U42851 ( .A(n43161), .B(n43158), .Z(n43160) );
  XNOR U42852 ( .A(n43154), .B(n43089), .Z(n43156) );
  XOR U42853 ( .A(n43162), .B(n43163), .Z(n43089) );
  AND U42854 ( .A(n1276), .B(n43124), .Z(n43163) );
  XOR U42855 ( .A(n43122), .B(n43162), .Z(n43124) );
  XOR U42856 ( .A(n43164), .B(n43165), .Z(n43154) );
  AND U42857 ( .A(n43166), .B(n43167), .Z(n43165) );
  XNOR U42858 ( .A(n43164), .B(n42991), .Z(n43167) );
  IV U42859 ( .A(n42994), .Z(n42991) );
  XOR U42860 ( .A(n43168), .B(n43169), .Z(n42994) );
  AND U42861 ( .A(n1268), .B(n43170), .Z(n43169) );
  XOR U42862 ( .A(n43171), .B(n43168), .Z(n43170) );
  XOR U42863 ( .A(n42995), .B(n43164), .Z(n43166) );
  XOR U42864 ( .A(n43172), .B(n43173), .Z(n42995) );
  AND U42865 ( .A(n1276), .B(n43132), .Z(n43173) );
  XOR U42866 ( .A(n43172), .B(n43130), .Z(n43132) );
  XOR U42867 ( .A(n43174), .B(n43175), .Z(n43164) );
  AND U42868 ( .A(n43176), .B(n43177), .Z(n43175) );
  XNOR U42869 ( .A(n43174), .B(n43019), .Z(n43177) );
  IV U42870 ( .A(n43022), .Z(n43019) );
  XOR U42871 ( .A(n43178), .B(n43179), .Z(n43022) );
  AND U42872 ( .A(n1268), .B(n43180), .Z(n43179) );
  XNOR U42873 ( .A(n43181), .B(n43178), .Z(n43180) );
  XOR U42874 ( .A(n43023), .B(n43174), .Z(n43176) );
  XOR U42875 ( .A(n43182), .B(n43183), .Z(n43023) );
  AND U42876 ( .A(n1276), .B(n43141), .Z(n43183) );
  XOR U42877 ( .A(n43182), .B(n43139), .Z(n43141) );
  XOR U42878 ( .A(n43098), .B(n43184), .Z(n43174) );
  AND U42879 ( .A(n43100), .B(n43185), .Z(n43184) );
  XNOR U42880 ( .A(n43098), .B(n43069), .Z(n43185) );
  IV U42881 ( .A(n43072), .Z(n43069) );
  XOR U42882 ( .A(n43186), .B(n43187), .Z(n43072) );
  AND U42883 ( .A(n1268), .B(n43188), .Z(n43187) );
  XOR U42884 ( .A(n43189), .B(n43186), .Z(n43188) );
  XOR U42885 ( .A(n43073), .B(n43098), .Z(n43100) );
  XOR U42886 ( .A(n43190), .B(n43191), .Z(n43073) );
  AND U42887 ( .A(n1276), .B(n43151), .Z(n43191) );
  XOR U42888 ( .A(n43190), .B(n43149), .Z(n43151) );
  AND U42889 ( .A(n43152), .B(n43082), .Z(n43098) );
  XNOR U42890 ( .A(n43192), .B(n43193), .Z(n43082) );
  AND U42891 ( .A(n1268), .B(n43194), .Z(n43193) );
  XNOR U42892 ( .A(n43195), .B(n43192), .Z(n43194) );
  XNOR U42893 ( .A(n43196), .B(n43197), .Z(n1268) );
  AND U42894 ( .A(n43198), .B(n43199), .Z(n43197) );
  XOR U42895 ( .A(n43161), .B(n43196), .Z(n43199) );
  AND U42896 ( .A(n43200), .B(n43201), .Z(n43161) );
  XNOR U42897 ( .A(n43158), .B(n43196), .Z(n43198) );
  XNOR U42898 ( .A(n43202), .B(n43203), .Z(n43158) );
  AND U42899 ( .A(n1272), .B(n43204), .Z(n43203) );
  XNOR U42900 ( .A(n43205), .B(n43206), .Z(n43204) );
  XOR U42901 ( .A(n43207), .B(n43208), .Z(n43196) );
  AND U42902 ( .A(n43209), .B(n43210), .Z(n43208) );
  XNOR U42903 ( .A(n43207), .B(n43200), .Z(n43210) );
  IV U42904 ( .A(n43171), .Z(n43200) );
  XOR U42905 ( .A(n43211), .B(n43212), .Z(n43171) );
  XOR U42906 ( .A(n43213), .B(n43201), .Z(n43212) );
  AND U42907 ( .A(n43181), .B(n43214), .Z(n43201) );
  AND U42908 ( .A(n43215), .B(n43216), .Z(n43213) );
  XOR U42909 ( .A(n43217), .B(n43211), .Z(n43215) );
  XNOR U42910 ( .A(n43168), .B(n43207), .Z(n43209) );
  XNOR U42911 ( .A(n43218), .B(n43219), .Z(n43168) );
  AND U42912 ( .A(n1272), .B(n43220), .Z(n43219) );
  XNOR U42913 ( .A(n43221), .B(n43222), .Z(n43220) );
  XOR U42914 ( .A(n43223), .B(n43224), .Z(n43207) );
  AND U42915 ( .A(n43225), .B(n43226), .Z(n43224) );
  XNOR U42916 ( .A(n43223), .B(n43181), .Z(n43226) );
  XOR U42917 ( .A(n43227), .B(n43216), .Z(n43181) );
  XNOR U42918 ( .A(n43228), .B(n43211), .Z(n43216) );
  XOR U42919 ( .A(n43229), .B(n43230), .Z(n43211) );
  AND U42920 ( .A(n43231), .B(n43232), .Z(n43230) );
  XOR U42921 ( .A(n43233), .B(n43229), .Z(n43231) );
  XNOR U42922 ( .A(n43234), .B(n43235), .Z(n43228) );
  AND U42923 ( .A(n43236), .B(n43237), .Z(n43235) );
  XOR U42924 ( .A(n43234), .B(n43238), .Z(n43236) );
  XNOR U42925 ( .A(n43217), .B(n43214), .Z(n43227) );
  AND U42926 ( .A(n43239), .B(n43240), .Z(n43214) );
  XOR U42927 ( .A(n43241), .B(n43242), .Z(n43217) );
  AND U42928 ( .A(n43243), .B(n43244), .Z(n43242) );
  XOR U42929 ( .A(n43241), .B(n43245), .Z(n43243) );
  XNOR U42930 ( .A(n43178), .B(n43223), .Z(n43225) );
  XNOR U42931 ( .A(n43246), .B(n43247), .Z(n43178) );
  AND U42932 ( .A(n1272), .B(n43248), .Z(n43247) );
  XNOR U42933 ( .A(n43249), .B(n43250), .Z(n43248) );
  XOR U42934 ( .A(n43251), .B(n43252), .Z(n43223) );
  AND U42935 ( .A(n43253), .B(n43254), .Z(n43252) );
  XNOR U42936 ( .A(n43251), .B(n43239), .Z(n43254) );
  IV U42937 ( .A(n43189), .Z(n43239) );
  XNOR U42938 ( .A(n43255), .B(n43232), .Z(n43189) );
  XNOR U42939 ( .A(n43256), .B(n43238), .Z(n43232) );
  XNOR U42940 ( .A(n43257), .B(n43258), .Z(n43238) );
  NOR U42941 ( .A(n43259), .B(n43260), .Z(n43258) );
  XOR U42942 ( .A(n43257), .B(n43261), .Z(n43259) );
  XNOR U42943 ( .A(n43237), .B(n43229), .Z(n43256) );
  XOR U42944 ( .A(n43262), .B(n43263), .Z(n43229) );
  AND U42945 ( .A(n43264), .B(n43265), .Z(n43263) );
  XOR U42946 ( .A(n43262), .B(n43266), .Z(n43264) );
  XNOR U42947 ( .A(n43267), .B(n43234), .Z(n43237) );
  XOR U42948 ( .A(n43268), .B(n43269), .Z(n43234) );
  AND U42949 ( .A(n43270), .B(n43271), .Z(n43269) );
  XNOR U42950 ( .A(n43272), .B(n43273), .Z(n43270) );
  IV U42951 ( .A(n43268), .Z(n43272) );
  XNOR U42952 ( .A(n43274), .B(n43275), .Z(n43267) );
  NOR U42953 ( .A(n43276), .B(n43277), .Z(n43275) );
  XNOR U42954 ( .A(n43274), .B(n43278), .Z(n43276) );
  XNOR U42955 ( .A(n43233), .B(n43240), .Z(n43255) );
  NOR U42956 ( .A(n43195), .B(n43279), .Z(n43240) );
  XOR U42957 ( .A(n43245), .B(n43244), .Z(n43233) );
  XNOR U42958 ( .A(n43280), .B(n43241), .Z(n43244) );
  XOR U42959 ( .A(n43281), .B(n43282), .Z(n43241) );
  AND U42960 ( .A(n43283), .B(n43284), .Z(n43282) );
  XNOR U42961 ( .A(n43285), .B(n43286), .Z(n43283) );
  IV U42962 ( .A(n43281), .Z(n43285) );
  XNOR U42963 ( .A(n43287), .B(n43288), .Z(n43280) );
  NOR U42964 ( .A(n43289), .B(n43290), .Z(n43288) );
  XNOR U42965 ( .A(n43287), .B(n43291), .Z(n43289) );
  XOR U42966 ( .A(n43292), .B(n43293), .Z(n43245) );
  NOR U42967 ( .A(n43294), .B(n43295), .Z(n43293) );
  XNOR U42968 ( .A(n43292), .B(n43296), .Z(n43294) );
  XNOR U42969 ( .A(n43186), .B(n43251), .Z(n43253) );
  XNOR U42970 ( .A(n43297), .B(n43298), .Z(n43186) );
  AND U42971 ( .A(n1272), .B(n43299), .Z(n43298) );
  XNOR U42972 ( .A(n43300), .B(n43301), .Z(n43299) );
  AND U42973 ( .A(n43192), .B(n43195), .Z(n43251) );
  XOR U42974 ( .A(n43302), .B(n43279), .Z(n43195) );
  XNOR U42975 ( .A(p_input[1008]), .B(p_input[2048]), .Z(n43279) );
  XNOR U42976 ( .A(n43266), .B(n43265), .Z(n43302) );
  XNOR U42977 ( .A(n43303), .B(n43273), .Z(n43265) );
  XNOR U42978 ( .A(n43261), .B(n43260), .Z(n43273) );
  XNOR U42979 ( .A(n43304), .B(n43257), .Z(n43260) );
  XNOR U42980 ( .A(p_input[1018]), .B(p_input[2058]), .Z(n43257) );
  XOR U42981 ( .A(p_input[1019]), .B(n29030), .Z(n43304) );
  XOR U42982 ( .A(p_input[1020]), .B(p_input[2060]), .Z(n43261) );
  XOR U42983 ( .A(n43271), .B(n43305), .Z(n43303) );
  IV U42984 ( .A(n43262), .Z(n43305) );
  XOR U42985 ( .A(p_input[1009]), .B(p_input[2049]), .Z(n43262) );
  XNOR U42986 ( .A(n43306), .B(n43278), .Z(n43271) );
  XNOR U42987 ( .A(p_input[1023]), .B(n29033), .Z(n43278) );
  XOR U42988 ( .A(n43268), .B(n43277), .Z(n43306) );
  XOR U42989 ( .A(n43307), .B(n43274), .Z(n43277) );
  XOR U42990 ( .A(p_input[1021]), .B(p_input[2061]), .Z(n43274) );
  XOR U42991 ( .A(p_input[1022]), .B(n29035), .Z(n43307) );
  XOR U42992 ( .A(p_input[1017]), .B(p_input[2057]), .Z(n43268) );
  XOR U42993 ( .A(n43286), .B(n43284), .Z(n43266) );
  XNOR U42994 ( .A(n43308), .B(n43291), .Z(n43284) );
  XOR U42995 ( .A(p_input[1016]), .B(p_input[2056]), .Z(n43291) );
  XOR U42996 ( .A(n43281), .B(n43290), .Z(n43308) );
  XOR U42997 ( .A(n43309), .B(n43287), .Z(n43290) );
  XOR U42998 ( .A(p_input[1014]), .B(p_input[2054]), .Z(n43287) );
  XOR U42999 ( .A(p_input[1015]), .B(n30404), .Z(n43309) );
  XOR U43000 ( .A(p_input[1010]), .B(p_input[2050]), .Z(n43281) );
  XNOR U43001 ( .A(n43296), .B(n43295), .Z(n43286) );
  XOR U43002 ( .A(n43310), .B(n43292), .Z(n43295) );
  XOR U43003 ( .A(p_input[1011]), .B(p_input[2051]), .Z(n43292) );
  XOR U43004 ( .A(p_input[1012]), .B(n30406), .Z(n43310) );
  XOR U43005 ( .A(p_input[1013]), .B(p_input[2053]), .Z(n43296) );
  XNOR U43006 ( .A(n43311), .B(n43312), .Z(n43192) );
  AND U43007 ( .A(n1272), .B(n43313), .Z(n43312) );
  XNOR U43008 ( .A(n43314), .B(n43315), .Z(n1272) );
  AND U43009 ( .A(n43316), .B(n43317), .Z(n43315) );
  XOR U43010 ( .A(n43206), .B(n43314), .Z(n43317) );
  XNOR U43011 ( .A(n43318), .B(n43314), .Z(n43316) );
  XOR U43012 ( .A(n43319), .B(n43320), .Z(n43314) );
  AND U43013 ( .A(n43321), .B(n43322), .Z(n43320) );
  XOR U43014 ( .A(n43221), .B(n43319), .Z(n43322) );
  XOR U43015 ( .A(n43319), .B(n43222), .Z(n43321) );
  XOR U43016 ( .A(n43323), .B(n43324), .Z(n43319) );
  AND U43017 ( .A(n43325), .B(n43326), .Z(n43324) );
  XOR U43018 ( .A(n43249), .B(n43323), .Z(n43326) );
  XOR U43019 ( .A(n43323), .B(n43250), .Z(n43325) );
  XOR U43020 ( .A(n43327), .B(n43328), .Z(n43323) );
  AND U43021 ( .A(n43329), .B(n43330), .Z(n43328) );
  XOR U43022 ( .A(n43327), .B(n43300), .Z(n43330) );
  XNOR U43023 ( .A(n43331), .B(n43332), .Z(n43152) );
  AND U43024 ( .A(n1276), .B(n43333), .Z(n43332) );
  XNOR U43025 ( .A(n43334), .B(n43335), .Z(n1276) );
  AND U43026 ( .A(n43336), .B(n43337), .Z(n43335) );
  XOR U43027 ( .A(n43334), .B(n43162), .Z(n43337) );
  XNOR U43028 ( .A(n43334), .B(n43122), .Z(n43336) );
  XOR U43029 ( .A(n43338), .B(n43339), .Z(n43334) );
  AND U43030 ( .A(n43340), .B(n43341), .Z(n43339) );
  XOR U43031 ( .A(n43338), .B(n43130), .Z(n43340) );
  XOR U43032 ( .A(n43342), .B(n43343), .Z(n43113) );
  AND U43033 ( .A(n1280), .B(n43333), .Z(n43343) );
  XNOR U43034 ( .A(n43331), .B(n43342), .Z(n43333) );
  XNOR U43035 ( .A(n43344), .B(n43345), .Z(n1280) );
  AND U43036 ( .A(n43346), .B(n43347), .Z(n43345) );
  XNOR U43037 ( .A(n43348), .B(n43344), .Z(n43347) );
  IV U43038 ( .A(n43162), .Z(n43348) );
  XOR U43039 ( .A(n43318), .B(n43349), .Z(n43162) );
  AND U43040 ( .A(n1283), .B(n43350), .Z(n43349) );
  XOR U43041 ( .A(n43205), .B(n43202), .Z(n43350) );
  IV U43042 ( .A(n43318), .Z(n43205) );
  XNOR U43043 ( .A(n43122), .B(n43344), .Z(n43346) );
  XOR U43044 ( .A(n43351), .B(n43352), .Z(n43122) );
  AND U43045 ( .A(n1299), .B(n43353), .Z(n43352) );
  XOR U43046 ( .A(n43338), .B(n43354), .Z(n43344) );
  AND U43047 ( .A(n43355), .B(n43341), .Z(n43354) );
  XNOR U43048 ( .A(n43172), .B(n43338), .Z(n43341) );
  XOR U43049 ( .A(n43222), .B(n43356), .Z(n43172) );
  AND U43050 ( .A(n1283), .B(n43357), .Z(n43356) );
  XOR U43051 ( .A(n43218), .B(n43222), .Z(n43357) );
  XNOR U43052 ( .A(n43358), .B(n43338), .Z(n43355) );
  IV U43053 ( .A(n43130), .Z(n43358) );
  XOR U43054 ( .A(n43359), .B(n43360), .Z(n43130) );
  AND U43055 ( .A(n1299), .B(n43361), .Z(n43360) );
  XOR U43056 ( .A(n43362), .B(n43363), .Z(n43338) );
  AND U43057 ( .A(n43364), .B(n43365), .Z(n43363) );
  XNOR U43058 ( .A(n43182), .B(n43362), .Z(n43365) );
  XOR U43059 ( .A(n43250), .B(n43366), .Z(n43182) );
  AND U43060 ( .A(n1283), .B(n43367), .Z(n43366) );
  XOR U43061 ( .A(n43246), .B(n43250), .Z(n43367) );
  XOR U43062 ( .A(n43362), .B(n43139), .Z(n43364) );
  XOR U43063 ( .A(n43368), .B(n43369), .Z(n43139) );
  AND U43064 ( .A(n1299), .B(n43370), .Z(n43369) );
  XOR U43065 ( .A(n43371), .B(n43372), .Z(n43362) );
  AND U43066 ( .A(n43373), .B(n43374), .Z(n43372) );
  XNOR U43067 ( .A(n43371), .B(n43190), .Z(n43374) );
  XOR U43068 ( .A(n43301), .B(n43375), .Z(n43190) );
  AND U43069 ( .A(n1283), .B(n43376), .Z(n43375) );
  XOR U43070 ( .A(n43297), .B(n43301), .Z(n43376) );
  XNOR U43071 ( .A(n43377), .B(n43371), .Z(n43373) );
  IV U43072 ( .A(n43149), .Z(n43377) );
  XOR U43073 ( .A(n43378), .B(n43379), .Z(n43149) );
  AND U43074 ( .A(n1299), .B(n43380), .Z(n43379) );
  AND U43075 ( .A(n43342), .B(n43331), .Z(n43371) );
  XNOR U43076 ( .A(n43381), .B(n43382), .Z(n43331) );
  AND U43077 ( .A(n1283), .B(n43313), .Z(n43382) );
  XNOR U43078 ( .A(n43311), .B(n43381), .Z(n43313) );
  XNOR U43079 ( .A(n43383), .B(n43384), .Z(n1283) );
  AND U43080 ( .A(n43385), .B(n43386), .Z(n43384) );
  XNOR U43081 ( .A(n43383), .B(n43202), .Z(n43386) );
  IV U43082 ( .A(n43206), .Z(n43202) );
  XOR U43083 ( .A(n43387), .B(n43388), .Z(n43206) );
  AND U43084 ( .A(n1287), .B(n43389), .Z(n43388) );
  XOR U43085 ( .A(n43390), .B(n43387), .Z(n43389) );
  XNOR U43086 ( .A(n43383), .B(n43318), .Z(n43385) );
  XOR U43087 ( .A(n43391), .B(n43392), .Z(n43318) );
  AND U43088 ( .A(n1295), .B(n43353), .Z(n43392) );
  XOR U43089 ( .A(n43351), .B(n43391), .Z(n43353) );
  XOR U43090 ( .A(n43393), .B(n43394), .Z(n43383) );
  AND U43091 ( .A(n43395), .B(n43396), .Z(n43394) );
  XNOR U43092 ( .A(n43393), .B(n43218), .Z(n43396) );
  IV U43093 ( .A(n43221), .Z(n43218) );
  XOR U43094 ( .A(n43397), .B(n43398), .Z(n43221) );
  AND U43095 ( .A(n1287), .B(n43399), .Z(n43398) );
  XOR U43096 ( .A(n43400), .B(n43397), .Z(n43399) );
  XOR U43097 ( .A(n43222), .B(n43393), .Z(n43395) );
  XOR U43098 ( .A(n43401), .B(n43402), .Z(n43222) );
  AND U43099 ( .A(n1295), .B(n43361), .Z(n43402) );
  XOR U43100 ( .A(n43401), .B(n43359), .Z(n43361) );
  XOR U43101 ( .A(n43403), .B(n43404), .Z(n43393) );
  AND U43102 ( .A(n43405), .B(n43406), .Z(n43404) );
  XNOR U43103 ( .A(n43403), .B(n43246), .Z(n43406) );
  IV U43104 ( .A(n43249), .Z(n43246) );
  XOR U43105 ( .A(n43407), .B(n43408), .Z(n43249) );
  AND U43106 ( .A(n1287), .B(n43409), .Z(n43408) );
  XNOR U43107 ( .A(n43410), .B(n43407), .Z(n43409) );
  XOR U43108 ( .A(n43250), .B(n43403), .Z(n43405) );
  XOR U43109 ( .A(n43411), .B(n43412), .Z(n43250) );
  AND U43110 ( .A(n1295), .B(n43370), .Z(n43412) );
  XOR U43111 ( .A(n43411), .B(n43368), .Z(n43370) );
  XOR U43112 ( .A(n43327), .B(n43413), .Z(n43403) );
  AND U43113 ( .A(n43329), .B(n43414), .Z(n43413) );
  XNOR U43114 ( .A(n43327), .B(n43297), .Z(n43414) );
  IV U43115 ( .A(n43300), .Z(n43297) );
  XOR U43116 ( .A(n43415), .B(n43416), .Z(n43300) );
  AND U43117 ( .A(n1287), .B(n43417), .Z(n43416) );
  XOR U43118 ( .A(n43418), .B(n43415), .Z(n43417) );
  XOR U43119 ( .A(n43301), .B(n43327), .Z(n43329) );
  XOR U43120 ( .A(n43419), .B(n43420), .Z(n43301) );
  AND U43121 ( .A(n1295), .B(n43380), .Z(n43420) );
  XOR U43122 ( .A(n43419), .B(n43378), .Z(n43380) );
  AND U43123 ( .A(n43381), .B(n43311), .Z(n43327) );
  XNOR U43124 ( .A(n43421), .B(n43422), .Z(n43311) );
  AND U43125 ( .A(n1287), .B(n43423), .Z(n43422) );
  XNOR U43126 ( .A(n43424), .B(n43421), .Z(n43423) );
  XNOR U43127 ( .A(n43425), .B(n43426), .Z(n1287) );
  AND U43128 ( .A(n43427), .B(n43428), .Z(n43426) );
  XOR U43129 ( .A(n43390), .B(n43425), .Z(n43428) );
  AND U43130 ( .A(n43429), .B(n43430), .Z(n43390) );
  XNOR U43131 ( .A(n43387), .B(n43425), .Z(n43427) );
  XNOR U43132 ( .A(n43431), .B(n43432), .Z(n43387) );
  AND U43133 ( .A(n1291), .B(n43433), .Z(n43432) );
  XNOR U43134 ( .A(n43434), .B(n43435), .Z(n43433) );
  XOR U43135 ( .A(n43436), .B(n43437), .Z(n43425) );
  AND U43136 ( .A(n43438), .B(n43439), .Z(n43437) );
  XNOR U43137 ( .A(n43436), .B(n43429), .Z(n43439) );
  IV U43138 ( .A(n43400), .Z(n43429) );
  XOR U43139 ( .A(n43440), .B(n43441), .Z(n43400) );
  XOR U43140 ( .A(n43442), .B(n43430), .Z(n43441) );
  AND U43141 ( .A(n43410), .B(n43443), .Z(n43430) );
  AND U43142 ( .A(n43444), .B(n43445), .Z(n43442) );
  XOR U43143 ( .A(n43446), .B(n43440), .Z(n43444) );
  XNOR U43144 ( .A(n43397), .B(n43436), .Z(n43438) );
  XNOR U43145 ( .A(n43447), .B(n43448), .Z(n43397) );
  AND U43146 ( .A(n1291), .B(n43449), .Z(n43448) );
  XNOR U43147 ( .A(n43450), .B(n43451), .Z(n43449) );
  XOR U43148 ( .A(n43452), .B(n43453), .Z(n43436) );
  AND U43149 ( .A(n43454), .B(n43455), .Z(n43453) );
  XNOR U43150 ( .A(n43452), .B(n43410), .Z(n43455) );
  XOR U43151 ( .A(n43456), .B(n43445), .Z(n43410) );
  XNOR U43152 ( .A(n43457), .B(n43440), .Z(n43445) );
  XOR U43153 ( .A(n43458), .B(n43459), .Z(n43440) );
  AND U43154 ( .A(n43460), .B(n43461), .Z(n43459) );
  XOR U43155 ( .A(n43462), .B(n43458), .Z(n43460) );
  XNOR U43156 ( .A(n43463), .B(n43464), .Z(n43457) );
  AND U43157 ( .A(n43465), .B(n43466), .Z(n43464) );
  XOR U43158 ( .A(n43463), .B(n43467), .Z(n43465) );
  XNOR U43159 ( .A(n43446), .B(n43443), .Z(n43456) );
  AND U43160 ( .A(n43468), .B(n43469), .Z(n43443) );
  XOR U43161 ( .A(n43470), .B(n43471), .Z(n43446) );
  AND U43162 ( .A(n43472), .B(n43473), .Z(n43471) );
  XOR U43163 ( .A(n43470), .B(n43474), .Z(n43472) );
  XNOR U43164 ( .A(n43407), .B(n43452), .Z(n43454) );
  XNOR U43165 ( .A(n43475), .B(n43476), .Z(n43407) );
  AND U43166 ( .A(n1291), .B(n43477), .Z(n43476) );
  XNOR U43167 ( .A(n43478), .B(n43479), .Z(n43477) );
  XOR U43168 ( .A(n43480), .B(n43481), .Z(n43452) );
  AND U43169 ( .A(n43482), .B(n43483), .Z(n43481) );
  XNOR U43170 ( .A(n43480), .B(n43468), .Z(n43483) );
  IV U43171 ( .A(n43418), .Z(n43468) );
  XNOR U43172 ( .A(n43484), .B(n43461), .Z(n43418) );
  XNOR U43173 ( .A(n43485), .B(n43467), .Z(n43461) );
  XNOR U43174 ( .A(n43486), .B(n43487), .Z(n43467) );
  NOR U43175 ( .A(n43488), .B(n43489), .Z(n43487) );
  XOR U43176 ( .A(n43486), .B(n43490), .Z(n43488) );
  XNOR U43177 ( .A(n43466), .B(n43458), .Z(n43485) );
  XOR U43178 ( .A(n43491), .B(n43492), .Z(n43458) );
  AND U43179 ( .A(n43493), .B(n43494), .Z(n43492) );
  XOR U43180 ( .A(n43491), .B(n43495), .Z(n43493) );
  XNOR U43181 ( .A(n43496), .B(n43463), .Z(n43466) );
  XOR U43182 ( .A(n43497), .B(n43498), .Z(n43463) );
  AND U43183 ( .A(n43499), .B(n43500), .Z(n43498) );
  XNOR U43184 ( .A(n43501), .B(n43502), .Z(n43499) );
  IV U43185 ( .A(n43497), .Z(n43501) );
  XNOR U43186 ( .A(n43503), .B(n43504), .Z(n43496) );
  NOR U43187 ( .A(n43505), .B(n43506), .Z(n43504) );
  XNOR U43188 ( .A(n43503), .B(n43507), .Z(n43505) );
  XNOR U43189 ( .A(n43462), .B(n43469), .Z(n43484) );
  NOR U43190 ( .A(n43424), .B(n43508), .Z(n43469) );
  XOR U43191 ( .A(n43474), .B(n43473), .Z(n43462) );
  XNOR U43192 ( .A(n43509), .B(n43470), .Z(n43473) );
  XOR U43193 ( .A(n43510), .B(n43511), .Z(n43470) );
  AND U43194 ( .A(n43512), .B(n43513), .Z(n43511) );
  XNOR U43195 ( .A(n43514), .B(n43515), .Z(n43512) );
  IV U43196 ( .A(n43510), .Z(n43514) );
  XNOR U43197 ( .A(n43516), .B(n43517), .Z(n43509) );
  NOR U43198 ( .A(n43518), .B(n43519), .Z(n43517) );
  XNOR U43199 ( .A(n43516), .B(n43520), .Z(n43518) );
  XOR U43200 ( .A(n43521), .B(n43522), .Z(n43474) );
  NOR U43201 ( .A(n43523), .B(n43524), .Z(n43522) );
  XNOR U43202 ( .A(n43521), .B(n43525), .Z(n43523) );
  XNOR U43203 ( .A(n43415), .B(n43480), .Z(n43482) );
  XNOR U43204 ( .A(n43526), .B(n43527), .Z(n43415) );
  AND U43205 ( .A(n1291), .B(n43528), .Z(n43527) );
  XNOR U43206 ( .A(n43529), .B(n43530), .Z(n43528) );
  AND U43207 ( .A(n43421), .B(n43424), .Z(n43480) );
  XOR U43208 ( .A(n43531), .B(n43508), .Z(n43424) );
  XNOR U43209 ( .A(p_input[1024]), .B(p_input[2048]), .Z(n43508) );
  XNOR U43210 ( .A(n43495), .B(n43494), .Z(n43531) );
  XNOR U43211 ( .A(n43532), .B(n43502), .Z(n43494) );
  XNOR U43212 ( .A(n43490), .B(n43489), .Z(n43502) );
  XNOR U43213 ( .A(n43533), .B(n43486), .Z(n43489) );
  XNOR U43214 ( .A(p_input[1034]), .B(p_input[2058]), .Z(n43486) );
  XOR U43215 ( .A(p_input[1035]), .B(n29030), .Z(n43533) );
  XOR U43216 ( .A(p_input[1036]), .B(p_input[2060]), .Z(n43490) );
  XOR U43217 ( .A(n43500), .B(n43534), .Z(n43532) );
  IV U43218 ( .A(n43491), .Z(n43534) );
  XOR U43219 ( .A(p_input[1025]), .B(p_input[2049]), .Z(n43491) );
  XNOR U43220 ( .A(n43535), .B(n43507), .Z(n43500) );
  XNOR U43221 ( .A(p_input[1039]), .B(n29033), .Z(n43507) );
  XOR U43222 ( .A(n43497), .B(n43506), .Z(n43535) );
  XOR U43223 ( .A(n43536), .B(n43503), .Z(n43506) );
  XOR U43224 ( .A(p_input[1037]), .B(p_input[2061]), .Z(n43503) );
  XOR U43225 ( .A(p_input[1038]), .B(n29035), .Z(n43536) );
  XOR U43226 ( .A(p_input[1033]), .B(p_input[2057]), .Z(n43497) );
  XOR U43227 ( .A(n43515), .B(n43513), .Z(n43495) );
  XNOR U43228 ( .A(n43537), .B(n43520), .Z(n43513) );
  XOR U43229 ( .A(p_input[1032]), .B(p_input[2056]), .Z(n43520) );
  XOR U43230 ( .A(n43510), .B(n43519), .Z(n43537) );
  XOR U43231 ( .A(n43538), .B(n43516), .Z(n43519) );
  XOR U43232 ( .A(p_input[1030]), .B(p_input[2054]), .Z(n43516) );
  XOR U43233 ( .A(p_input[1031]), .B(n30404), .Z(n43538) );
  XOR U43234 ( .A(p_input[1026]), .B(p_input[2050]), .Z(n43510) );
  XNOR U43235 ( .A(n43525), .B(n43524), .Z(n43515) );
  XOR U43236 ( .A(n43539), .B(n43521), .Z(n43524) );
  XOR U43237 ( .A(p_input[1027]), .B(p_input[2051]), .Z(n43521) );
  XOR U43238 ( .A(p_input[1028]), .B(n30406), .Z(n43539) );
  XOR U43239 ( .A(p_input[1029]), .B(p_input[2053]), .Z(n43525) );
  XNOR U43240 ( .A(n43540), .B(n43541), .Z(n43421) );
  AND U43241 ( .A(n1291), .B(n43542), .Z(n43541) );
  XNOR U43242 ( .A(n43543), .B(n43544), .Z(n1291) );
  AND U43243 ( .A(n43545), .B(n43546), .Z(n43544) );
  XOR U43244 ( .A(n43435), .B(n43543), .Z(n43546) );
  XNOR U43245 ( .A(n43547), .B(n43543), .Z(n43545) );
  XOR U43246 ( .A(n43548), .B(n43549), .Z(n43543) );
  AND U43247 ( .A(n43550), .B(n43551), .Z(n43549) );
  XOR U43248 ( .A(n43450), .B(n43548), .Z(n43551) );
  XOR U43249 ( .A(n43548), .B(n43451), .Z(n43550) );
  XOR U43250 ( .A(n43552), .B(n43553), .Z(n43548) );
  AND U43251 ( .A(n43554), .B(n43555), .Z(n43553) );
  XOR U43252 ( .A(n43478), .B(n43552), .Z(n43555) );
  XOR U43253 ( .A(n43552), .B(n43479), .Z(n43554) );
  XOR U43254 ( .A(n43556), .B(n43557), .Z(n43552) );
  AND U43255 ( .A(n43558), .B(n43559), .Z(n43557) );
  XOR U43256 ( .A(n43556), .B(n43529), .Z(n43559) );
  XNOR U43257 ( .A(n43560), .B(n43561), .Z(n43381) );
  AND U43258 ( .A(n1295), .B(n43562), .Z(n43561) );
  XNOR U43259 ( .A(n43563), .B(n43564), .Z(n1295) );
  AND U43260 ( .A(n43565), .B(n43566), .Z(n43564) );
  XOR U43261 ( .A(n43563), .B(n43391), .Z(n43566) );
  XNOR U43262 ( .A(n43563), .B(n43351), .Z(n43565) );
  XOR U43263 ( .A(n43567), .B(n43568), .Z(n43563) );
  AND U43264 ( .A(n43569), .B(n43570), .Z(n43568) );
  XOR U43265 ( .A(n43567), .B(n43359), .Z(n43569) );
  XOR U43266 ( .A(n43571), .B(n43572), .Z(n43342) );
  AND U43267 ( .A(n1299), .B(n43562), .Z(n43572) );
  XNOR U43268 ( .A(n43560), .B(n43571), .Z(n43562) );
  XNOR U43269 ( .A(n43573), .B(n43574), .Z(n1299) );
  AND U43270 ( .A(n43575), .B(n43576), .Z(n43574) );
  XNOR U43271 ( .A(n43577), .B(n43573), .Z(n43576) );
  IV U43272 ( .A(n43391), .Z(n43577) );
  XOR U43273 ( .A(n43547), .B(n43578), .Z(n43391) );
  AND U43274 ( .A(n1302), .B(n43579), .Z(n43578) );
  XOR U43275 ( .A(n43434), .B(n43431), .Z(n43579) );
  IV U43276 ( .A(n43547), .Z(n43434) );
  XNOR U43277 ( .A(n43351), .B(n43573), .Z(n43575) );
  XOR U43278 ( .A(n43580), .B(n43581), .Z(n43351) );
  AND U43279 ( .A(n1318), .B(n43582), .Z(n43581) );
  XOR U43280 ( .A(n43567), .B(n43583), .Z(n43573) );
  AND U43281 ( .A(n43584), .B(n43570), .Z(n43583) );
  XNOR U43282 ( .A(n43401), .B(n43567), .Z(n43570) );
  XOR U43283 ( .A(n43451), .B(n43585), .Z(n43401) );
  AND U43284 ( .A(n1302), .B(n43586), .Z(n43585) );
  XOR U43285 ( .A(n43447), .B(n43451), .Z(n43586) );
  XNOR U43286 ( .A(n43587), .B(n43567), .Z(n43584) );
  IV U43287 ( .A(n43359), .Z(n43587) );
  XOR U43288 ( .A(n43588), .B(n43589), .Z(n43359) );
  AND U43289 ( .A(n1318), .B(n43590), .Z(n43589) );
  XOR U43290 ( .A(n43591), .B(n43592), .Z(n43567) );
  AND U43291 ( .A(n43593), .B(n43594), .Z(n43592) );
  XNOR U43292 ( .A(n43411), .B(n43591), .Z(n43594) );
  XOR U43293 ( .A(n43479), .B(n43595), .Z(n43411) );
  AND U43294 ( .A(n1302), .B(n43596), .Z(n43595) );
  XOR U43295 ( .A(n43475), .B(n43479), .Z(n43596) );
  XOR U43296 ( .A(n43591), .B(n43368), .Z(n43593) );
  XOR U43297 ( .A(n43597), .B(n43598), .Z(n43368) );
  AND U43298 ( .A(n1318), .B(n43599), .Z(n43598) );
  XOR U43299 ( .A(n43600), .B(n43601), .Z(n43591) );
  AND U43300 ( .A(n43602), .B(n43603), .Z(n43601) );
  XNOR U43301 ( .A(n43600), .B(n43419), .Z(n43603) );
  XOR U43302 ( .A(n43530), .B(n43604), .Z(n43419) );
  AND U43303 ( .A(n1302), .B(n43605), .Z(n43604) );
  XOR U43304 ( .A(n43526), .B(n43530), .Z(n43605) );
  XNOR U43305 ( .A(n43606), .B(n43600), .Z(n43602) );
  IV U43306 ( .A(n43378), .Z(n43606) );
  XOR U43307 ( .A(n43607), .B(n43608), .Z(n43378) );
  AND U43308 ( .A(n1318), .B(n43609), .Z(n43608) );
  AND U43309 ( .A(n43571), .B(n43560), .Z(n43600) );
  XNOR U43310 ( .A(n43610), .B(n43611), .Z(n43560) );
  AND U43311 ( .A(n1302), .B(n43542), .Z(n43611) );
  XNOR U43312 ( .A(n43540), .B(n43610), .Z(n43542) );
  XNOR U43313 ( .A(n43612), .B(n43613), .Z(n1302) );
  AND U43314 ( .A(n43614), .B(n43615), .Z(n43613) );
  XNOR U43315 ( .A(n43612), .B(n43431), .Z(n43615) );
  IV U43316 ( .A(n43435), .Z(n43431) );
  XOR U43317 ( .A(n43616), .B(n43617), .Z(n43435) );
  AND U43318 ( .A(n1306), .B(n43618), .Z(n43617) );
  XOR U43319 ( .A(n43619), .B(n43616), .Z(n43618) );
  XNOR U43320 ( .A(n43612), .B(n43547), .Z(n43614) );
  XOR U43321 ( .A(n43620), .B(n43621), .Z(n43547) );
  AND U43322 ( .A(n1314), .B(n43582), .Z(n43621) );
  XOR U43323 ( .A(n43580), .B(n43620), .Z(n43582) );
  XOR U43324 ( .A(n43622), .B(n43623), .Z(n43612) );
  AND U43325 ( .A(n43624), .B(n43625), .Z(n43623) );
  XNOR U43326 ( .A(n43622), .B(n43447), .Z(n43625) );
  IV U43327 ( .A(n43450), .Z(n43447) );
  XOR U43328 ( .A(n43626), .B(n43627), .Z(n43450) );
  AND U43329 ( .A(n1306), .B(n43628), .Z(n43627) );
  XOR U43330 ( .A(n43629), .B(n43626), .Z(n43628) );
  XOR U43331 ( .A(n43451), .B(n43622), .Z(n43624) );
  XOR U43332 ( .A(n43630), .B(n43631), .Z(n43451) );
  AND U43333 ( .A(n1314), .B(n43590), .Z(n43631) );
  XOR U43334 ( .A(n43630), .B(n43588), .Z(n43590) );
  XOR U43335 ( .A(n43632), .B(n43633), .Z(n43622) );
  AND U43336 ( .A(n43634), .B(n43635), .Z(n43633) );
  XNOR U43337 ( .A(n43632), .B(n43475), .Z(n43635) );
  IV U43338 ( .A(n43478), .Z(n43475) );
  XOR U43339 ( .A(n43636), .B(n43637), .Z(n43478) );
  AND U43340 ( .A(n1306), .B(n43638), .Z(n43637) );
  XNOR U43341 ( .A(n43639), .B(n43636), .Z(n43638) );
  XOR U43342 ( .A(n43479), .B(n43632), .Z(n43634) );
  XOR U43343 ( .A(n43640), .B(n43641), .Z(n43479) );
  AND U43344 ( .A(n1314), .B(n43599), .Z(n43641) );
  XOR U43345 ( .A(n43640), .B(n43597), .Z(n43599) );
  XOR U43346 ( .A(n43556), .B(n43642), .Z(n43632) );
  AND U43347 ( .A(n43558), .B(n43643), .Z(n43642) );
  XNOR U43348 ( .A(n43556), .B(n43526), .Z(n43643) );
  IV U43349 ( .A(n43529), .Z(n43526) );
  XOR U43350 ( .A(n43644), .B(n43645), .Z(n43529) );
  AND U43351 ( .A(n1306), .B(n43646), .Z(n43645) );
  XOR U43352 ( .A(n43647), .B(n43644), .Z(n43646) );
  XOR U43353 ( .A(n43530), .B(n43556), .Z(n43558) );
  XOR U43354 ( .A(n43648), .B(n43649), .Z(n43530) );
  AND U43355 ( .A(n1314), .B(n43609), .Z(n43649) );
  XOR U43356 ( .A(n43648), .B(n43607), .Z(n43609) );
  AND U43357 ( .A(n43610), .B(n43540), .Z(n43556) );
  XNOR U43358 ( .A(n43650), .B(n43651), .Z(n43540) );
  AND U43359 ( .A(n1306), .B(n43652), .Z(n43651) );
  XNOR U43360 ( .A(n43653), .B(n43650), .Z(n43652) );
  XNOR U43361 ( .A(n43654), .B(n43655), .Z(n1306) );
  AND U43362 ( .A(n43656), .B(n43657), .Z(n43655) );
  XOR U43363 ( .A(n43619), .B(n43654), .Z(n43657) );
  AND U43364 ( .A(n43658), .B(n43659), .Z(n43619) );
  XNOR U43365 ( .A(n43616), .B(n43654), .Z(n43656) );
  XNOR U43366 ( .A(n43660), .B(n43661), .Z(n43616) );
  AND U43367 ( .A(n1310), .B(n43662), .Z(n43661) );
  XNOR U43368 ( .A(n43663), .B(n43664), .Z(n43662) );
  XOR U43369 ( .A(n43665), .B(n43666), .Z(n43654) );
  AND U43370 ( .A(n43667), .B(n43668), .Z(n43666) );
  XNOR U43371 ( .A(n43665), .B(n43658), .Z(n43668) );
  IV U43372 ( .A(n43629), .Z(n43658) );
  XOR U43373 ( .A(n43669), .B(n43670), .Z(n43629) );
  XOR U43374 ( .A(n43671), .B(n43659), .Z(n43670) );
  AND U43375 ( .A(n43639), .B(n43672), .Z(n43659) );
  AND U43376 ( .A(n43673), .B(n43674), .Z(n43671) );
  XOR U43377 ( .A(n43675), .B(n43669), .Z(n43673) );
  XNOR U43378 ( .A(n43626), .B(n43665), .Z(n43667) );
  XNOR U43379 ( .A(n43676), .B(n43677), .Z(n43626) );
  AND U43380 ( .A(n1310), .B(n43678), .Z(n43677) );
  XNOR U43381 ( .A(n43679), .B(n43680), .Z(n43678) );
  XOR U43382 ( .A(n43681), .B(n43682), .Z(n43665) );
  AND U43383 ( .A(n43683), .B(n43684), .Z(n43682) );
  XNOR U43384 ( .A(n43681), .B(n43639), .Z(n43684) );
  XOR U43385 ( .A(n43685), .B(n43674), .Z(n43639) );
  XNOR U43386 ( .A(n43686), .B(n43669), .Z(n43674) );
  XOR U43387 ( .A(n43687), .B(n43688), .Z(n43669) );
  AND U43388 ( .A(n43689), .B(n43690), .Z(n43688) );
  XOR U43389 ( .A(n43691), .B(n43687), .Z(n43689) );
  XNOR U43390 ( .A(n43692), .B(n43693), .Z(n43686) );
  AND U43391 ( .A(n43694), .B(n43695), .Z(n43693) );
  XOR U43392 ( .A(n43692), .B(n43696), .Z(n43694) );
  XNOR U43393 ( .A(n43675), .B(n43672), .Z(n43685) );
  AND U43394 ( .A(n43697), .B(n43698), .Z(n43672) );
  XOR U43395 ( .A(n43699), .B(n43700), .Z(n43675) );
  AND U43396 ( .A(n43701), .B(n43702), .Z(n43700) );
  XOR U43397 ( .A(n43699), .B(n43703), .Z(n43701) );
  XNOR U43398 ( .A(n43636), .B(n43681), .Z(n43683) );
  XNOR U43399 ( .A(n43704), .B(n43705), .Z(n43636) );
  AND U43400 ( .A(n1310), .B(n43706), .Z(n43705) );
  XNOR U43401 ( .A(n43707), .B(n43708), .Z(n43706) );
  XOR U43402 ( .A(n43709), .B(n43710), .Z(n43681) );
  AND U43403 ( .A(n43711), .B(n43712), .Z(n43710) );
  XNOR U43404 ( .A(n43709), .B(n43697), .Z(n43712) );
  IV U43405 ( .A(n43647), .Z(n43697) );
  XNOR U43406 ( .A(n43713), .B(n43690), .Z(n43647) );
  XNOR U43407 ( .A(n43714), .B(n43696), .Z(n43690) );
  XNOR U43408 ( .A(n43715), .B(n43716), .Z(n43696) );
  NOR U43409 ( .A(n43717), .B(n43718), .Z(n43716) );
  XOR U43410 ( .A(n43715), .B(n43719), .Z(n43717) );
  XNOR U43411 ( .A(n43695), .B(n43687), .Z(n43714) );
  XOR U43412 ( .A(n43720), .B(n43721), .Z(n43687) );
  AND U43413 ( .A(n43722), .B(n43723), .Z(n43721) );
  XOR U43414 ( .A(n43720), .B(n43724), .Z(n43722) );
  XNOR U43415 ( .A(n43725), .B(n43692), .Z(n43695) );
  XOR U43416 ( .A(n43726), .B(n43727), .Z(n43692) );
  AND U43417 ( .A(n43728), .B(n43729), .Z(n43727) );
  XNOR U43418 ( .A(n43730), .B(n43731), .Z(n43728) );
  IV U43419 ( .A(n43726), .Z(n43730) );
  XNOR U43420 ( .A(n43732), .B(n43733), .Z(n43725) );
  NOR U43421 ( .A(n43734), .B(n43735), .Z(n43733) );
  XNOR U43422 ( .A(n43732), .B(n43736), .Z(n43734) );
  XNOR U43423 ( .A(n43691), .B(n43698), .Z(n43713) );
  NOR U43424 ( .A(n43653), .B(n43737), .Z(n43698) );
  XOR U43425 ( .A(n43703), .B(n43702), .Z(n43691) );
  XNOR U43426 ( .A(n43738), .B(n43699), .Z(n43702) );
  XOR U43427 ( .A(n43739), .B(n43740), .Z(n43699) );
  AND U43428 ( .A(n43741), .B(n43742), .Z(n43740) );
  XNOR U43429 ( .A(n43743), .B(n43744), .Z(n43741) );
  IV U43430 ( .A(n43739), .Z(n43743) );
  XNOR U43431 ( .A(n43745), .B(n43746), .Z(n43738) );
  NOR U43432 ( .A(n43747), .B(n43748), .Z(n43746) );
  XNOR U43433 ( .A(n43745), .B(n43749), .Z(n43747) );
  XOR U43434 ( .A(n43750), .B(n43751), .Z(n43703) );
  NOR U43435 ( .A(n43752), .B(n43753), .Z(n43751) );
  XNOR U43436 ( .A(n43750), .B(n43754), .Z(n43752) );
  XNOR U43437 ( .A(n43644), .B(n43709), .Z(n43711) );
  XNOR U43438 ( .A(n43755), .B(n43756), .Z(n43644) );
  AND U43439 ( .A(n1310), .B(n43757), .Z(n43756) );
  XNOR U43440 ( .A(n43758), .B(n43759), .Z(n43757) );
  AND U43441 ( .A(n43650), .B(n43653), .Z(n43709) );
  XOR U43442 ( .A(n43760), .B(n43737), .Z(n43653) );
  XNOR U43443 ( .A(p_input[1040]), .B(p_input[2048]), .Z(n43737) );
  XNOR U43444 ( .A(n43724), .B(n43723), .Z(n43760) );
  XNOR U43445 ( .A(n43761), .B(n43731), .Z(n43723) );
  XNOR U43446 ( .A(n43719), .B(n43718), .Z(n43731) );
  XNOR U43447 ( .A(n43762), .B(n43715), .Z(n43718) );
  XNOR U43448 ( .A(p_input[1050]), .B(p_input[2058]), .Z(n43715) );
  XOR U43449 ( .A(p_input[1051]), .B(n29030), .Z(n43762) );
  XOR U43450 ( .A(p_input[1052]), .B(p_input[2060]), .Z(n43719) );
  XOR U43451 ( .A(n43729), .B(n43763), .Z(n43761) );
  IV U43452 ( .A(n43720), .Z(n43763) );
  XOR U43453 ( .A(p_input[1041]), .B(p_input[2049]), .Z(n43720) );
  XNOR U43454 ( .A(n43764), .B(n43736), .Z(n43729) );
  XNOR U43455 ( .A(p_input[1055]), .B(n29033), .Z(n43736) );
  XOR U43456 ( .A(n43726), .B(n43735), .Z(n43764) );
  XOR U43457 ( .A(n43765), .B(n43732), .Z(n43735) );
  XOR U43458 ( .A(p_input[1053]), .B(p_input[2061]), .Z(n43732) );
  XOR U43459 ( .A(p_input[1054]), .B(n29035), .Z(n43765) );
  XOR U43460 ( .A(p_input[1049]), .B(p_input[2057]), .Z(n43726) );
  XOR U43461 ( .A(n43744), .B(n43742), .Z(n43724) );
  XNOR U43462 ( .A(n43766), .B(n43749), .Z(n43742) );
  XOR U43463 ( .A(p_input[1048]), .B(p_input[2056]), .Z(n43749) );
  XOR U43464 ( .A(n43739), .B(n43748), .Z(n43766) );
  XOR U43465 ( .A(n43767), .B(n43745), .Z(n43748) );
  XOR U43466 ( .A(p_input[1046]), .B(p_input[2054]), .Z(n43745) );
  XOR U43467 ( .A(p_input[1047]), .B(n30404), .Z(n43767) );
  XOR U43468 ( .A(p_input[1042]), .B(p_input[2050]), .Z(n43739) );
  XNOR U43469 ( .A(n43754), .B(n43753), .Z(n43744) );
  XOR U43470 ( .A(n43768), .B(n43750), .Z(n43753) );
  XOR U43471 ( .A(p_input[1043]), .B(p_input[2051]), .Z(n43750) );
  XOR U43472 ( .A(p_input[1044]), .B(n30406), .Z(n43768) );
  XOR U43473 ( .A(p_input[1045]), .B(p_input[2053]), .Z(n43754) );
  XNOR U43474 ( .A(n43769), .B(n43770), .Z(n43650) );
  AND U43475 ( .A(n1310), .B(n43771), .Z(n43770) );
  XNOR U43476 ( .A(n43772), .B(n43773), .Z(n1310) );
  AND U43477 ( .A(n43774), .B(n43775), .Z(n43773) );
  XOR U43478 ( .A(n43664), .B(n43772), .Z(n43775) );
  XNOR U43479 ( .A(n43776), .B(n43772), .Z(n43774) );
  XOR U43480 ( .A(n43777), .B(n43778), .Z(n43772) );
  AND U43481 ( .A(n43779), .B(n43780), .Z(n43778) );
  XOR U43482 ( .A(n43679), .B(n43777), .Z(n43780) );
  XOR U43483 ( .A(n43777), .B(n43680), .Z(n43779) );
  XOR U43484 ( .A(n43781), .B(n43782), .Z(n43777) );
  AND U43485 ( .A(n43783), .B(n43784), .Z(n43782) );
  XOR U43486 ( .A(n43707), .B(n43781), .Z(n43784) );
  XOR U43487 ( .A(n43781), .B(n43708), .Z(n43783) );
  XOR U43488 ( .A(n43785), .B(n43786), .Z(n43781) );
  AND U43489 ( .A(n43787), .B(n43788), .Z(n43786) );
  XOR U43490 ( .A(n43785), .B(n43758), .Z(n43788) );
  XNOR U43491 ( .A(n43789), .B(n43790), .Z(n43610) );
  AND U43492 ( .A(n1314), .B(n43791), .Z(n43790) );
  XNOR U43493 ( .A(n43792), .B(n43793), .Z(n1314) );
  AND U43494 ( .A(n43794), .B(n43795), .Z(n43793) );
  XOR U43495 ( .A(n43792), .B(n43620), .Z(n43795) );
  XNOR U43496 ( .A(n43792), .B(n43580), .Z(n43794) );
  XOR U43497 ( .A(n43796), .B(n43797), .Z(n43792) );
  AND U43498 ( .A(n43798), .B(n43799), .Z(n43797) );
  XOR U43499 ( .A(n43796), .B(n43588), .Z(n43798) );
  XOR U43500 ( .A(n43800), .B(n43801), .Z(n43571) );
  AND U43501 ( .A(n1318), .B(n43791), .Z(n43801) );
  XNOR U43502 ( .A(n43789), .B(n43800), .Z(n43791) );
  XNOR U43503 ( .A(n43802), .B(n43803), .Z(n1318) );
  AND U43504 ( .A(n43804), .B(n43805), .Z(n43803) );
  XNOR U43505 ( .A(n43806), .B(n43802), .Z(n43805) );
  IV U43506 ( .A(n43620), .Z(n43806) );
  XOR U43507 ( .A(n43776), .B(n43807), .Z(n43620) );
  AND U43508 ( .A(n1321), .B(n43808), .Z(n43807) );
  XOR U43509 ( .A(n43663), .B(n43660), .Z(n43808) );
  IV U43510 ( .A(n43776), .Z(n43663) );
  XNOR U43511 ( .A(n43580), .B(n43802), .Z(n43804) );
  XOR U43512 ( .A(n43809), .B(n43810), .Z(n43580) );
  AND U43513 ( .A(n1337), .B(n43811), .Z(n43810) );
  XOR U43514 ( .A(n43796), .B(n43812), .Z(n43802) );
  AND U43515 ( .A(n43813), .B(n43799), .Z(n43812) );
  XNOR U43516 ( .A(n43630), .B(n43796), .Z(n43799) );
  XOR U43517 ( .A(n43680), .B(n43814), .Z(n43630) );
  AND U43518 ( .A(n1321), .B(n43815), .Z(n43814) );
  XOR U43519 ( .A(n43676), .B(n43680), .Z(n43815) );
  XNOR U43520 ( .A(n43816), .B(n43796), .Z(n43813) );
  IV U43521 ( .A(n43588), .Z(n43816) );
  XOR U43522 ( .A(n43817), .B(n43818), .Z(n43588) );
  AND U43523 ( .A(n1337), .B(n43819), .Z(n43818) );
  XOR U43524 ( .A(n43820), .B(n43821), .Z(n43796) );
  AND U43525 ( .A(n43822), .B(n43823), .Z(n43821) );
  XNOR U43526 ( .A(n43640), .B(n43820), .Z(n43823) );
  XOR U43527 ( .A(n43708), .B(n43824), .Z(n43640) );
  AND U43528 ( .A(n1321), .B(n43825), .Z(n43824) );
  XOR U43529 ( .A(n43704), .B(n43708), .Z(n43825) );
  XOR U43530 ( .A(n43820), .B(n43597), .Z(n43822) );
  XOR U43531 ( .A(n43826), .B(n43827), .Z(n43597) );
  AND U43532 ( .A(n1337), .B(n43828), .Z(n43827) );
  XOR U43533 ( .A(n43829), .B(n43830), .Z(n43820) );
  AND U43534 ( .A(n43831), .B(n43832), .Z(n43830) );
  XNOR U43535 ( .A(n43829), .B(n43648), .Z(n43832) );
  XOR U43536 ( .A(n43759), .B(n43833), .Z(n43648) );
  AND U43537 ( .A(n1321), .B(n43834), .Z(n43833) );
  XOR U43538 ( .A(n43755), .B(n43759), .Z(n43834) );
  XNOR U43539 ( .A(n43835), .B(n43829), .Z(n43831) );
  IV U43540 ( .A(n43607), .Z(n43835) );
  XOR U43541 ( .A(n43836), .B(n43837), .Z(n43607) );
  AND U43542 ( .A(n1337), .B(n43838), .Z(n43837) );
  AND U43543 ( .A(n43800), .B(n43789), .Z(n43829) );
  XNOR U43544 ( .A(n43839), .B(n43840), .Z(n43789) );
  AND U43545 ( .A(n1321), .B(n43771), .Z(n43840) );
  XNOR U43546 ( .A(n43769), .B(n43839), .Z(n43771) );
  XNOR U43547 ( .A(n43841), .B(n43842), .Z(n1321) );
  AND U43548 ( .A(n43843), .B(n43844), .Z(n43842) );
  XNOR U43549 ( .A(n43841), .B(n43660), .Z(n43844) );
  IV U43550 ( .A(n43664), .Z(n43660) );
  XOR U43551 ( .A(n43845), .B(n43846), .Z(n43664) );
  AND U43552 ( .A(n1325), .B(n43847), .Z(n43846) );
  XOR U43553 ( .A(n43848), .B(n43845), .Z(n43847) );
  XNOR U43554 ( .A(n43841), .B(n43776), .Z(n43843) );
  XOR U43555 ( .A(n43849), .B(n43850), .Z(n43776) );
  AND U43556 ( .A(n1333), .B(n43811), .Z(n43850) );
  XOR U43557 ( .A(n43809), .B(n43849), .Z(n43811) );
  XOR U43558 ( .A(n43851), .B(n43852), .Z(n43841) );
  AND U43559 ( .A(n43853), .B(n43854), .Z(n43852) );
  XNOR U43560 ( .A(n43851), .B(n43676), .Z(n43854) );
  IV U43561 ( .A(n43679), .Z(n43676) );
  XOR U43562 ( .A(n43855), .B(n43856), .Z(n43679) );
  AND U43563 ( .A(n1325), .B(n43857), .Z(n43856) );
  XOR U43564 ( .A(n43858), .B(n43855), .Z(n43857) );
  XOR U43565 ( .A(n43680), .B(n43851), .Z(n43853) );
  XOR U43566 ( .A(n43859), .B(n43860), .Z(n43680) );
  AND U43567 ( .A(n1333), .B(n43819), .Z(n43860) );
  XOR U43568 ( .A(n43859), .B(n43817), .Z(n43819) );
  XOR U43569 ( .A(n43861), .B(n43862), .Z(n43851) );
  AND U43570 ( .A(n43863), .B(n43864), .Z(n43862) );
  XNOR U43571 ( .A(n43861), .B(n43704), .Z(n43864) );
  IV U43572 ( .A(n43707), .Z(n43704) );
  XOR U43573 ( .A(n43865), .B(n43866), .Z(n43707) );
  AND U43574 ( .A(n1325), .B(n43867), .Z(n43866) );
  XNOR U43575 ( .A(n43868), .B(n43865), .Z(n43867) );
  XOR U43576 ( .A(n43708), .B(n43861), .Z(n43863) );
  XOR U43577 ( .A(n43869), .B(n43870), .Z(n43708) );
  AND U43578 ( .A(n1333), .B(n43828), .Z(n43870) );
  XOR U43579 ( .A(n43869), .B(n43826), .Z(n43828) );
  XOR U43580 ( .A(n43785), .B(n43871), .Z(n43861) );
  AND U43581 ( .A(n43787), .B(n43872), .Z(n43871) );
  XNOR U43582 ( .A(n43785), .B(n43755), .Z(n43872) );
  IV U43583 ( .A(n43758), .Z(n43755) );
  XOR U43584 ( .A(n43873), .B(n43874), .Z(n43758) );
  AND U43585 ( .A(n1325), .B(n43875), .Z(n43874) );
  XOR U43586 ( .A(n43876), .B(n43873), .Z(n43875) );
  XOR U43587 ( .A(n43759), .B(n43785), .Z(n43787) );
  XOR U43588 ( .A(n43877), .B(n43878), .Z(n43759) );
  AND U43589 ( .A(n1333), .B(n43838), .Z(n43878) );
  XOR U43590 ( .A(n43877), .B(n43836), .Z(n43838) );
  AND U43591 ( .A(n43839), .B(n43769), .Z(n43785) );
  XNOR U43592 ( .A(n43879), .B(n43880), .Z(n43769) );
  AND U43593 ( .A(n1325), .B(n43881), .Z(n43880) );
  XNOR U43594 ( .A(n43882), .B(n43879), .Z(n43881) );
  XNOR U43595 ( .A(n43883), .B(n43884), .Z(n1325) );
  AND U43596 ( .A(n43885), .B(n43886), .Z(n43884) );
  XOR U43597 ( .A(n43848), .B(n43883), .Z(n43886) );
  AND U43598 ( .A(n43887), .B(n43888), .Z(n43848) );
  XNOR U43599 ( .A(n43845), .B(n43883), .Z(n43885) );
  XNOR U43600 ( .A(n43889), .B(n43890), .Z(n43845) );
  AND U43601 ( .A(n1329), .B(n43891), .Z(n43890) );
  XNOR U43602 ( .A(n43892), .B(n43893), .Z(n43891) );
  XOR U43603 ( .A(n43894), .B(n43895), .Z(n43883) );
  AND U43604 ( .A(n43896), .B(n43897), .Z(n43895) );
  XNOR U43605 ( .A(n43894), .B(n43887), .Z(n43897) );
  IV U43606 ( .A(n43858), .Z(n43887) );
  XOR U43607 ( .A(n43898), .B(n43899), .Z(n43858) );
  XOR U43608 ( .A(n43900), .B(n43888), .Z(n43899) );
  AND U43609 ( .A(n43868), .B(n43901), .Z(n43888) );
  AND U43610 ( .A(n43902), .B(n43903), .Z(n43900) );
  XOR U43611 ( .A(n43904), .B(n43898), .Z(n43902) );
  XNOR U43612 ( .A(n43855), .B(n43894), .Z(n43896) );
  XNOR U43613 ( .A(n43905), .B(n43906), .Z(n43855) );
  AND U43614 ( .A(n1329), .B(n43907), .Z(n43906) );
  XNOR U43615 ( .A(n43908), .B(n43909), .Z(n43907) );
  XOR U43616 ( .A(n43910), .B(n43911), .Z(n43894) );
  AND U43617 ( .A(n43912), .B(n43913), .Z(n43911) );
  XNOR U43618 ( .A(n43910), .B(n43868), .Z(n43913) );
  XOR U43619 ( .A(n43914), .B(n43903), .Z(n43868) );
  XNOR U43620 ( .A(n43915), .B(n43898), .Z(n43903) );
  XOR U43621 ( .A(n43916), .B(n43917), .Z(n43898) );
  AND U43622 ( .A(n43918), .B(n43919), .Z(n43917) );
  XOR U43623 ( .A(n43920), .B(n43916), .Z(n43918) );
  XNOR U43624 ( .A(n43921), .B(n43922), .Z(n43915) );
  AND U43625 ( .A(n43923), .B(n43924), .Z(n43922) );
  XOR U43626 ( .A(n43921), .B(n43925), .Z(n43923) );
  XNOR U43627 ( .A(n43904), .B(n43901), .Z(n43914) );
  AND U43628 ( .A(n43926), .B(n43927), .Z(n43901) );
  XOR U43629 ( .A(n43928), .B(n43929), .Z(n43904) );
  AND U43630 ( .A(n43930), .B(n43931), .Z(n43929) );
  XOR U43631 ( .A(n43928), .B(n43932), .Z(n43930) );
  XNOR U43632 ( .A(n43865), .B(n43910), .Z(n43912) );
  XNOR U43633 ( .A(n43933), .B(n43934), .Z(n43865) );
  AND U43634 ( .A(n1329), .B(n43935), .Z(n43934) );
  XNOR U43635 ( .A(n43936), .B(n43937), .Z(n43935) );
  XOR U43636 ( .A(n43938), .B(n43939), .Z(n43910) );
  AND U43637 ( .A(n43940), .B(n43941), .Z(n43939) );
  XNOR U43638 ( .A(n43938), .B(n43926), .Z(n43941) );
  IV U43639 ( .A(n43876), .Z(n43926) );
  XNOR U43640 ( .A(n43942), .B(n43919), .Z(n43876) );
  XNOR U43641 ( .A(n43943), .B(n43925), .Z(n43919) );
  XNOR U43642 ( .A(n43944), .B(n43945), .Z(n43925) );
  NOR U43643 ( .A(n43946), .B(n43947), .Z(n43945) );
  XOR U43644 ( .A(n43944), .B(n43948), .Z(n43946) );
  XNOR U43645 ( .A(n43924), .B(n43916), .Z(n43943) );
  XOR U43646 ( .A(n43949), .B(n43950), .Z(n43916) );
  AND U43647 ( .A(n43951), .B(n43952), .Z(n43950) );
  XOR U43648 ( .A(n43949), .B(n43953), .Z(n43951) );
  XNOR U43649 ( .A(n43954), .B(n43921), .Z(n43924) );
  XOR U43650 ( .A(n43955), .B(n43956), .Z(n43921) );
  AND U43651 ( .A(n43957), .B(n43958), .Z(n43956) );
  XNOR U43652 ( .A(n43959), .B(n43960), .Z(n43957) );
  IV U43653 ( .A(n43955), .Z(n43959) );
  XNOR U43654 ( .A(n43961), .B(n43962), .Z(n43954) );
  NOR U43655 ( .A(n43963), .B(n43964), .Z(n43962) );
  XNOR U43656 ( .A(n43961), .B(n43965), .Z(n43963) );
  XNOR U43657 ( .A(n43920), .B(n43927), .Z(n43942) );
  NOR U43658 ( .A(n43882), .B(n43966), .Z(n43927) );
  XOR U43659 ( .A(n43932), .B(n43931), .Z(n43920) );
  XNOR U43660 ( .A(n43967), .B(n43928), .Z(n43931) );
  XOR U43661 ( .A(n43968), .B(n43969), .Z(n43928) );
  AND U43662 ( .A(n43970), .B(n43971), .Z(n43969) );
  XNOR U43663 ( .A(n43972), .B(n43973), .Z(n43970) );
  IV U43664 ( .A(n43968), .Z(n43972) );
  XNOR U43665 ( .A(n43974), .B(n43975), .Z(n43967) );
  NOR U43666 ( .A(n43976), .B(n43977), .Z(n43975) );
  XNOR U43667 ( .A(n43974), .B(n43978), .Z(n43976) );
  XOR U43668 ( .A(n43979), .B(n43980), .Z(n43932) );
  NOR U43669 ( .A(n43981), .B(n43982), .Z(n43980) );
  XNOR U43670 ( .A(n43979), .B(n43983), .Z(n43981) );
  XNOR U43671 ( .A(n43873), .B(n43938), .Z(n43940) );
  XNOR U43672 ( .A(n43984), .B(n43985), .Z(n43873) );
  AND U43673 ( .A(n1329), .B(n43986), .Z(n43985) );
  XNOR U43674 ( .A(n43987), .B(n43988), .Z(n43986) );
  AND U43675 ( .A(n43879), .B(n43882), .Z(n43938) );
  XOR U43676 ( .A(n43989), .B(n43966), .Z(n43882) );
  XNOR U43677 ( .A(p_input[1056]), .B(p_input[2048]), .Z(n43966) );
  XNOR U43678 ( .A(n43953), .B(n43952), .Z(n43989) );
  XNOR U43679 ( .A(n43990), .B(n43960), .Z(n43952) );
  XNOR U43680 ( .A(n43948), .B(n43947), .Z(n43960) );
  XNOR U43681 ( .A(n43991), .B(n43944), .Z(n43947) );
  XNOR U43682 ( .A(p_input[1066]), .B(p_input[2058]), .Z(n43944) );
  XOR U43683 ( .A(p_input[1067]), .B(n29030), .Z(n43991) );
  XOR U43684 ( .A(p_input[1068]), .B(p_input[2060]), .Z(n43948) );
  XOR U43685 ( .A(n43958), .B(n43992), .Z(n43990) );
  IV U43686 ( .A(n43949), .Z(n43992) );
  XOR U43687 ( .A(p_input[1057]), .B(p_input[2049]), .Z(n43949) );
  XNOR U43688 ( .A(n43993), .B(n43965), .Z(n43958) );
  XNOR U43689 ( .A(p_input[1071]), .B(n29033), .Z(n43965) );
  XOR U43690 ( .A(n43955), .B(n43964), .Z(n43993) );
  XOR U43691 ( .A(n43994), .B(n43961), .Z(n43964) );
  XOR U43692 ( .A(p_input[1069]), .B(p_input[2061]), .Z(n43961) );
  XOR U43693 ( .A(p_input[1070]), .B(n29035), .Z(n43994) );
  XOR U43694 ( .A(p_input[1065]), .B(p_input[2057]), .Z(n43955) );
  XOR U43695 ( .A(n43973), .B(n43971), .Z(n43953) );
  XNOR U43696 ( .A(n43995), .B(n43978), .Z(n43971) );
  XOR U43697 ( .A(p_input[1064]), .B(p_input[2056]), .Z(n43978) );
  XOR U43698 ( .A(n43968), .B(n43977), .Z(n43995) );
  XOR U43699 ( .A(n43996), .B(n43974), .Z(n43977) );
  XOR U43700 ( .A(p_input[1062]), .B(p_input[2054]), .Z(n43974) );
  XOR U43701 ( .A(p_input[1063]), .B(n30404), .Z(n43996) );
  XOR U43702 ( .A(p_input[1058]), .B(p_input[2050]), .Z(n43968) );
  XNOR U43703 ( .A(n43983), .B(n43982), .Z(n43973) );
  XOR U43704 ( .A(n43997), .B(n43979), .Z(n43982) );
  XOR U43705 ( .A(p_input[1059]), .B(p_input[2051]), .Z(n43979) );
  XOR U43706 ( .A(p_input[1060]), .B(n30406), .Z(n43997) );
  XOR U43707 ( .A(p_input[1061]), .B(p_input[2053]), .Z(n43983) );
  XNOR U43708 ( .A(n43998), .B(n43999), .Z(n43879) );
  AND U43709 ( .A(n1329), .B(n44000), .Z(n43999) );
  XNOR U43710 ( .A(n44001), .B(n44002), .Z(n1329) );
  AND U43711 ( .A(n44003), .B(n44004), .Z(n44002) );
  XOR U43712 ( .A(n43893), .B(n44001), .Z(n44004) );
  XNOR U43713 ( .A(n44005), .B(n44001), .Z(n44003) );
  XOR U43714 ( .A(n44006), .B(n44007), .Z(n44001) );
  AND U43715 ( .A(n44008), .B(n44009), .Z(n44007) );
  XOR U43716 ( .A(n43908), .B(n44006), .Z(n44009) );
  XOR U43717 ( .A(n44006), .B(n43909), .Z(n44008) );
  XOR U43718 ( .A(n44010), .B(n44011), .Z(n44006) );
  AND U43719 ( .A(n44012), .B(n44013), .Z(n44011) );
  XOR U43720 ( .A(n43936), .B(n44010), .Z(n44013) );
  XOR U43721 ( .A(n44010), .B(n43937), .Z(n44012) );
  XOR U43722 ( .A(n44014), .B(n44015), .Z(n44010) );
  AND U43723 ( .A(n44016), .B(n44017), .Z(n44015) );
  XOR U43724 ( .A(n44014), .B(n43987), .Z(n44017) );
  XNOR U43725 ( .A(n44018), .B(n44019), .Z(n43839) );
  AND U43726 ( .A(n1333), .B(n44020), .Z(n44019) );
  XNOR U43727 ( .A(n44021), .B(n44022), .Z(n1333) );
  AND U43728 ( .A(n44023), .B(n44024), .Z(n44022) );
  XOR U43729 ( .A(n44021), .B(n43849), .Z(n44024) );
  XNOR U43730 ( .A(n44021), .B(n43809), .Z(n44023) );
  XOR U43731 ( .A(n44025), .B(n44026), .Z(n44021) );
  AND U43732 ( .A(n44027), .B(n44028), .Z(n44026) );
  XOR U43733 ( .A(n44025), .B(n43817), .Z(n44027) );
  XOR U43734 ( .A(n44029), .B(n44030), .Z(n43800) );
  AND U43735 ( .A(n1337), .B(n44020), .Z(n44030) );
  XNOR U43736 ( .A(n44018), .B(n44029), .Z(n44020) );
  XNOR U43737 ( .A(n44031), .B(n44032), .Z(n1337) );
  AND U43738 ( .A(n44033), .B(n44034), .Z(n44032) );
  XNOR U43739 ( .A(n44035), .B(n44031), .Z(n44034) );
  IV U43740 ( .A(n43849), .Z(n44035) );
  XOR U43741 ( .A(n44005), .B(n44036), .Z(n43849) );
  AND U43742 ( .A(n1340), .B(n44037), .Z(n44036) );
  XOR U43743 ( .A(n43892), .B(n43889), .Z(n44037) );
  IV U43744 ( .A(n44005), .Z(n43892) );
  XNOR U43745 ( .A(n43809), .B(n44031), .Z(n44033) );
  XOR U43746 ( .A(n44038), .B(n44039), .Z(n43809) );
  AND U43747 ( .A(n1356), .B(n44040), .Z(n44039) );
  XOR U43748 ( .A(n44025), .B(n44041), .Z(n44031) );
  AND U43749 ( .A(n44042), .B(n44028), .Z(n44041) );
  XNOR U43750 ( .A(n43859), .B(n44025), .Z(n44028) );
  XOR U43751 ( .A(n43909), .B(n44043), .Z(n43859) );
  AND U43752 ( .A(n1340), .B(n44044), .Z(n44043) );
  XOR U43753 ( .A(n43905), .B(n43909), .Z(n44044) );
  XNOR U43754 ( .A(n44045), .B(n44025), .Z(n44042) );
  IV U43755 ( .A(n43817), .Z(n44045) );
  XOR U43756 ( .A(n44046), .B(n44047), .Z(n43817) );
  AND U43757 ( .A(n1356), .B(n44048), .Z(n44047) );
  XOR U43758 ( .A(n44049), .B(n44050), .Z(n44025) );
  AND U43759 ( .A(n44051), .B(n44052), .Z(n44050) );
  XNOR U43760 ( .A(n43869), .B(n44049), .Z(n44052) );
  XOR U43761 ( .A(n43937), .B(n44053), .Z(n43869) );
  AND U43762 ( .A(n1340), .B(n44054), .Z(n44053) );
  XOR U43763 ( .A(n43933), .B(n43937), .Z(n44054) );
  XOR U43764 ( .A(n44049), .B(n43826), .Z(n44051) );
  XOR U43765 ( .A(n44055), .B(n44056), .Z(n43826) );
  AND U43766 ( .A(n1356), .B(n44057), .Z(n44056) );
  XOR U43767 ( .A(n44058), .B(n44059), .Z(n44049) );
  AND U43768 ( .A(n44060), .B(n44061), .Z(n44059) );
  XNOR U43769 ( .A(n44058), .B(n43877), .Z(n44061) );
  XOR U43770 ( .A(n43988), .B(n44062), .Z(n43877) );
  AND U43771 ( .A(n1340), .B(n44063), .Z(n44062) );
  XOR U43772 ( .A(n43984), .B(n43988), .Z(n44063) );
  XNOR U43773 ( .A(n44064), .B(n44058), .Z(n44060) );
  IV U43774 ( .A(n43836), .Z(n44064) );
  XOR U43775 ( .A(n44065), .B(n44066), .Z(n43836) );
  AND U43776 ( .A(n1356), .B(n44067), .Z(n44066) );
  AND U43777 ( .A(n44029), .B(n44018), .Z(n44058) );
  XNOR U43778 ( .A(n44068), .B(n44069), .Z(n44018) );
  AND U43779 ( .A(n1340), .B(n44000), .Z(n44069) );
  XNOR U43780 ( .A(n43998), .B(n44068), .Z(n44000) );
  XNOR U43781 ( .A(n44070), .B(n44071), .Z(n1340) );
  AND U43782 ( .A(n44072), .B(n44073), .Z(n44071) );
  XNOR U43783 ( .A(n44070), .B(n43889), .Z(n44073) );
  IV U43784 ( .A(n43893), .Z(n43889) );
  XOR U43785 ( .A(n44074), .B(n44075), .Z(n43893) );
  AND U43786 ( .A(n1344), .B(n44076), .Z(n44075) );
  XOR U43787 ( .A(n44077), .B(n44074), .Z(n44076) );
  XNOR U43788 ( .A(n44070), .B(n44005), .Z(n44072) );
  XOR U43789 ( .A(n44078), .B(n44079), .Z(n44005) );
  AND U43790 ( .A(n1352), .B(n44040), .Z(n44079) );
  XOR U43791 ( .A(n44038), .B(n44078), .Z(n44040) );
  XOR U43792 ( .A(n44080), .B(n44081), .Z(n44070) );
  AND U43793 ( .A(n44082), .B(n44083), .Z(n44081) );
  XNOR U43794 ( .A(n44080), .B(n43905), .Z(n44083) );
  IV U43795 ( .A(n43908), .Z(n43905) );
  XOR U43796 ( .A(n44084), .B(n44085), .Z(n43908) );
  AND U43797 ( .A(n1344), .B(n44086), .Z(n44085) );
  XOR U43798 ( .A(n44087), .B(n44084), .Z(n44086) );
  XOR U43799 ( .A(n43909), .B(n44080), .Z(n44082) );
  XOR U43800 ( .A(n44088), .B(n44089), .Z(n43909) );
  AND U43801 ( .A(n1352), .B(n44048), .Z(n44089) );
  XOR U43802 ( .A(n44088), .B(n44046), .Z(n44048) );
  XOR U43803 ( .A(n44090), .B(n44091), .Z(n44080) );
  AND U43804 ( .A(n44092), .B(n44093), .Z(n44091) );
  XNOR U43805 ( .A(n44090), .B(n43933), .Z(n44093) );
  IV U43806 ( .A(n43936), .Z(n43933) );
  XOR U43807 ( .A(n44094), .B(n44095), .Z(n43936) );
  AND U43808 ( .A(n1344), .B(n44096), .Z(n44095) );
  XNOR U43809 ( .A(n44097), .B(n44094), .Z(n44096) );
  XOR U43810 ( .A(n43937), .B(n44090), .Z(n44092) );
  XOR U43811 ( .A(n44098), .B(n44099), .Z(n43937) );
  AND U43812 ( .A(n1352), .B(n44057), .Z(n44099) );
  XOR U43813 ( .A(n44098), .B(n44055), .Z(n44057) );
  XOR U43814 ( .A(n44014), .B(n44100), .Z(n44090) );
  AND U43815 ( .A(n44016), .B(n44101), .Z(n44100) );
  XNOR U43816 ( .A(n44014), .B(n43984), .Z(n44101) );
  IV U43817 ( .A(n43987), .Z(n43984) );
  XOR U43818 ( .A(n44102), .B(n44103), .Z(n43987) );
  AND U43819 ( .A(n1344), .B(n44104), .Z(n44103) );
  XOR U43820 ( .A(n44105), .B(n44102), .Z(n44104) );
  XOR U43821 ( .A(n43988), .B(n44014), .Z(n44016) );
  XOR U43822 ( .A(n44106), .B(n44107), .Z(n43988) );
  AND U43823 ( .A(n1352), .B(n44067), .Z(n44107) );
  XOR U43824 ( .A(n44106), .B(n44065), .Z(n44067) );
  AND U43825 ( .A(n44068), .B(n43998), .Z(n44014) );
  XNOR U43826 ( .A(n44108), .B(n44109), .Z(n43998) );
  AND U43827 ( .A(n1344), .B(n44110), .Z(n44109) );
  XNOR U43828 ( .A(n44111), .B(n44108), .Z(n44110) );
  XNOR U43829 ( .A(n44112), .B(n44113), .Z(n1344) );
  AND U43830 ( .A(n44114), .B(n44115), .Z(n44113) );
  XOR U43831 ( .A(n44077), .B(n44112), .Z(n44115) );
  AND U43832 ( .A(n44116), .B(n44117), .Z(n44077) );
  XNOR U43833 ( .A(n44074), .B(n44112), .Z(n44114) );
  XNOR U43834 ( .A(n44118), .B(n44119), .Z(n44074) );
  AND U43835 ( .A(n1348), .B(n44120), .Z(n44119) );
  XNOR U43836 ( .A(n44121), .B(n44122), .Z(n44120) );
  XOR U43837 ( .A(n44123), .B(n44124), .Z(n44112) );
  AND U43838 ( .A(n44125), .B(n44126), .Z(n44124) );
  XNOR U43839 ( .A(n44123), .B(n44116), .Z(n44126) );
  IV U43840 ( .A(n44087), .Z(n44116) );
  XOR U43841 ( .A(n44127), .B(n44128), .Z(n44087) );
  XOR U43842 ( .A(n44129), .B(n44117), .Z(n44128) );
  AND U43843 ( .A(n44097), .B(n44130), .Z(n44117) );
  AND U43844 ( .A(n44131), .B(n44132), .Z(n44129) );
  XOR U43845 ( .A(n44133), .B(n44127), .Z(n44131) );
  XNOR U43846 ( .A(n44084), .B(n44123), .Z(n44125) );
  XNOR U43847 ( .A(n44134), .B(n44135), .Z(n44084) );
  AND U43848 ( .A(n1348), .B(n44136), .Z(n44135) );
  XNOR U43849 ( .A(n44137), .B(n44138), .Z(n44136) );
  XOR U43850 ( .A(n44139), .B(n44140), .Z(n44123) );
  AND U43851 ( .A(n44141), .B(n44142), .Z(n44140) );
  XNOR U43852 ( .A(n44139), .B(n44097), .Z(n44142) );
  XOR U43853 ( .A(n44143), .B(n44132), .Z(n44097) );
  XNOR U43854 ( .A(n44144), .B(n44127), .Z(n44132) );
  XOR U43855 ( .A(n44145), .B(n44146), .Z(n44127) );
  AND U43856 ( .A(n44147), .B(n44148), .Z(n44146) );
  XOR U43857 ( .A(n44149), .B(n44145), .Z(n44147) );
  XNOR U43858 ( .A(n44150), .B(n44151), .Z(n44144) );
  AND U43859 ( .A(n44152), .B(n44153), .Z(n44151) );
  XOR U43860 ( .A(n44150), .B(n44154), .Z(n44152) );
  XNOR U43861 ( .A(n44133), .B(n44130), .Z(n44143) );
  AND U43862 ( .A(n44155), .B(n44156), .Z(n44130) );
  XOR U43863 ( .A(n44157), .B(n44158), .Z(n44133) );
  AND U43864 ( .A(n44159), .B(n44160), .Z(n44158) );
  XOR U43865 ( .A(n44157), .B(n44161), .Z(n44159) );
  XNOR U43866 ( .A(n44094), .B(n44139), .Z(n44141) );
  XNOR U43867 ( .A(n44162), .B(n44163), .Z(n44094) );
  AND U43868 ( .A(n1348), .B(n44164), .Z(n44163) );
  XNOR U43869 ( .A(n44165), .B(n44166), .Z(n44164) );
  XOR U43870 ( .A(n44167), .B(n44168), .Z(n44139) );
  AND U43871 ( .A(n44169), .B(n44170), .Z(n44168) );
  XNOR U43872 ( .A(n44167), .B(n44155), .Z(n44170) );
  IV U43873 ( .A(n44105), .Z(n44155) );
  XNOR U43874 ( .A(n44171), .B(n44148), .Z(n44105) );
  XNOR U43875 ( .A(n44172), .B(n44154), .Z(n44148) );
  XNOR U43876 ( .A(n44173), .B(n44174), .Z(n44154) );
  NOR U43877 ( .A(n44175), .B(n44176), .Z(n44174) );
  XOR U43878 ( .A(n44173), .B(n44177), .Z(n44175) );
  XNOR U43879 ( .A(n44153), .B(n44145), .Z(n44172) );
  XOR U43880 ( .A(n44178), .B(n44179), .Z(n44145) );
  AND U43881 ( .A(n44180), .B(n44181), .Z(n44179) );
  XOR U43882 ( .A(n44178), .B(n44182), .Z(n44180) );
  XNOR U43883 ( .A(n44183), .B(n44150), .Z(n44153) );
  XOR U43884 ( .A(n44184), .B(n44185), .Z(n44150) );
  AND U43885 ( .A(n44186), .B(n44187), .Z(n44185) );
  XNOR U43886 ( .A(n44188), .B(n44189), .Z(n44186) );
  IV U43887 ( .A(n44184), .Z(n44188) );
  XNOR U43888 ( .A(n44190), .B(n44191), .Z(n44183) );
  NOR U43889 ( .A(n44192), .B(n44193), .Z(n44191) );
  XNOR U43890 ( .A(n44190), .B(n44194), .Z(n44192) );
  XNOR U43891 ( .A(n44149), .B(n44156), .Z(n44171) );
  NOR U43892 ( .A(n44111), .B(n44195), .Z(n44156) );
  XOR U43893 ( .A(n44161), .B(n44160), .Z(n44149) );
  XNOR U43894 ( .A(n44196), .B(n44157), .Z(n44160) );
  XOR U43895 ( .A(n44197), .B(n44198), .Z(n44157) );
  AND U43896 ( .A(n44199), .B(n44200), .Z(n44198) );
  XNOR U43897 ( .A(n44201), .B(n44202), .Z(n44199) );
  IV U43898 ( .A(n44197), .Z(n44201) );
  XNOR U43899 ( .A(n44203), .B(n44204), .Z(n44196) );
  NOR U43900 ( .A(n44205), .B(n44206), .Z(n44204) );
  XNOR U43901 ( .A(n44203), .B(n44207), .Z(n44205) );
  XOR U43902 ( .A(n44208), .B(n44209), .Z(n44161) );
  NOR U43903 ( .A(n44210), .B(n44211), .Z(n44209) );
  XNOR U43904 ( .A(n44208), .B(n44212), .Z(n44210) );
  XNOR U43905 ( .A(n44102), .B(n44167), .Z(n44169) );
  XNOR U43906 ( .A(n44213), .B(n44214), .Z(n44102) );
  AND U43907 ( .A(n1348), .B(n44215), .Z(n44214) );
  XNOR U43908 ( .A(n44216), .B(n44217), .Z(n44215) );
  AND U43909 ( .A(n44108), .B(n44111), .Z(n44167) );
  XOR U43910 ( .A(n44218), .B(n44195), .Z(n44111) );
  XNOR U43911 ( .A(p_input[1072]), .B(p_input[2048]), .Z(n44195) );
  XNOR U43912 ( .A(n44182), .B(n44181), .Z(n44218) );
  XNOR U43913 ( .A(n44219), .B(n44189), .Z(n44181) );
  XNOR U43914 ( .A(n44177), .B(n44176), .Z(n44189) );
  XNOR U43915 ( .A(n44220), .B(n44173), .Z(n44176) );
  XNOR U43916 ( .A(p_input[1082]), .B(p_input[2058]), .Z(n44173) );
  XOR U43917 ( .A(p_input[1083]), .B(n29030), .Z(n44220) );
  XOR U43918 ( .A(p_input[1084]), .B(p_input[2060]), .Z(n44177) );
  XOR U43919 ( .A(n44187), .B(n44221), .Z(n44219) );
  IV U43920 ( .A(n44178), .Z(n44221) );
  XOR U43921 ( .A(p_input[1073]), .B(p_input[2049]), .Z(n44178) );
  XNOR U43922 ( .A(n44222), .B(n44194), .Z(n44187) );
  XNOR U43923 ( .A(p_input[1087]), .B(n29033), .Z(n44194) );
  XOR U43924 ( .A(n44184), .B(n44193), .Z(n44222) );
  XOR U43925 ( .A(n44223), .B(n44190), .Z(n44193) );
  XOR U43926 ( .A(p_input[1085]), .B(p_input[2061]), .Z(n44190) );
  XOR U43927 ( .A(p_input[1086]), .B(n29035), .Z(n44223) );
  XOR U43928 ( .A(p_input[1081]), .B(p_input[2057]), .Z(n44184) );
  XOR U43929 ( .A(n44202), .B(n44200), .Z(n44182) );
  XNOR U43930 ( .A(n44224), .B(n44207), .Z(n44200) );
  XOR U43931 ( .A(p_input[1080]), .B(p_input[2056]), .Z(n44207) );
  XOR U43932 ( .A(n44197), .B(n44206), .Z(n44224) );
  XOR U43933 ( .A(n44225), .B(n44203), .Z(n44206) );
  XOR U43934 ( .A(p_input[1078]), .B(p_input[2054]), .Z(n44203) );
  XOR U43935 ( .A(p_input[1079]), .B(n30404), .Z(n44225) );
  XOR U43936 ( .A(p_input[1074]), .B(p_input[2050]), .Z(n44197) );
  XNOR U43937 ( .A(n44212), .B(n44211), .Z(n44202) );
  XOR U43938 ( .A(n44226), .B(n44208), .Z(n44211) );
  XOR U43939 ( .A(p_input[1075]), .B(p_input[2051]), .Z(n44208) );
  XOR U43940 ( .A(p_input[1076]), .B(n30406), .Z(n44226) );
  XOR U43941 ( .A(p_input[1077]), .B(p_input[2053]), .Z(n44212) );
  XNOR U43942 ( .A(n44227), .B(n44228), .Z(n44108) );
  AND U43943 ( .A(n1348), .B(n44229), .Z(n44228) );
  XNOR U43944 ( .A(n44230), .B(n44231), .Z(n1348) );
  AND U43945 ( .A(n44232), .B(n44233), .Z(n44231) );
  XOR U43946 ( .A(n44122), .B(n44230), .Z(n44233) );
  XNOR U43947 ( .A(n44234), .B(n44230), .Z(n44232) );
  XOR U43948 ( .A(n44235), .B(n44236), .Z(n44230) );
  AND U43949 ( .A(n44237), .B(n44238), .Z(n44236) );
  XOR U43950 ( .A(n44137), .B(n44235), .Z(n44238) );
  XOR U43951 ( .A(n44235), .B(n44138), .Z(n44237) );
  XOR U43952 ( .A(n44239), .B(n44240), .Z(n44235) );
  AND U43953 ( .A(n44241), .B(n44242), .Z(n44240) );
  XOR U43954 ( .A(n44165), .B(n44239), .Z(n44242) );
  XOR U43955 ( .A(n44239), .B(n44166), .Z(n44241) );
  XOR U43956 ( .A(n44243), .B(n44244), .Z(n44239) );
  AND U43957 ( .A(n44245), .B(n44246), .Z(n44244) );
  XOR U43958 ( .A(n44243), .B(n44216), .Z(n44246) );
  XNOR U43959 ( .A(n44247), .B(n44248), .Z(n44068) );
  AND U43960 ( .A(n1352), .B(n44249), .Z(n44248) );
  XNOR U43961 ( .A(n44250), .B(n44251), .Z(n1352) );
  AND U43962 ( .A(n44252), .B(n44253), .Z(n44251) );
  XOR U43963 ( .A(n44250), .B(n44078), .Z(n44253) );
  XNOR U43964 ( .A(n44250), .B(n44038), .Z(n44252) );
  XOR U43965 ( .A(n44254), .B(n44255), .Z(n44250) );
  AND U43966 ( .A(n44256), .B(n44257), .Z(n44255) );
  XOR U43967 ( .A(n44254), .B(n44046), .Z(n44256) );
  XOR U43968 ( .A(n44258), .B(n44259), .Z(n44029) );
  AND U43969 ( .A(n1356), .B(n44249), .Z(n44259) );
  XNOR U43970 ( .A(n44247), .B(n44258), .Z(n44249) );
  XNOR U43971 ( .A(n44260), .B(n44261), .Z(n1356) );
  AND U43972 ( .A(n44262), .B(n44263), .Z(n44261) );
  XNOR U43973 ( .A(n44264), .B(n44260), .Z(n44263) );
  IV U43974 ( .A(n44078), .Z(n44264) );
  XOR U43975 ( .A(n44234), .B(n44265), .Z(n44078) );
  AND U43976 ( .A(n1359), .B(n44266), .Z(n44265) );
  XOR U43977 ( .A(n44121), .B(n44118), .Z(n44266) );
  IV U43978 ( .A(n44234), .Z(n44121) );
  XNOR U43979 ( .A(n44038), .B(n44260), .Z(n44262) );
  XOR U43980 ( .A(n44267), .B(n44268), .Z(n44038) );
  AND U43981 ( .A(n1375), .B(n44269), .Z(n44268) );
  XOR U43982 ( .A(n44254), .B(n44270), .Z(n44260) );
  AND U43983 ( .A(n44271), .B(n44257), .Z(n44270) );
  XNOR U43984 ( .A(n44088), .B(n44254), .Z(n44257) );
  XOR U43985 ( .A(n44138), .B(n44272), .Z(n44088) );
  AND U43986 ( .A(n1359), .B(n44273), .Z(n44272) );
  XOR U43987 ( .A(n44134), .B(n44138), .Z(n44273) );
  XNOR U43988 ( .A(n44274), .B(n44254), .Z(n44271) );
  IV U43989 ( .A(n44046), .Z(n44274) );
  XOR U43990 ( .A(n44275), .B(n44276), .Z(n44046) );
  AND U43991 ( .A(n1375), .B(n44277), .Z(n44276) );
  XOR U43992 ( .A(n44278), .B(n44279), .Z(n44254) );
  AND U43993 ( .A(n44280), .B(n44281), .Z(n44279) );
  XNOR U43994 ( .A(n44098), .B(n44278), .Z(n44281) );
  XOR U43995 ( .A(n44166), .B(n44282), .Z(n44098) );
  AND U43996 ( .A(n1359), .B(n44283), .Z(n44282) );
  XOR U43997 ( .A(n44162), .B(n44166), .Z(n44283) );
  XOR U43998 ( .A(n44278), .B(n44055), .Z(n44280) );
  XOR U43999 ( .A(n44284), .B(n44285), .Z(n44055) );
  AND U44000 ( .A(n1375), .B(n44286), .Z(n44285) );
  XOR U44001 ( .A(n44287), .B(n44288), .Z(n44278) );
  AND U44002 ( .A(n44289), .B(n44290), .Z(n44288) );
  XNOR U44003 ( .A(n44287), .B(n44106), .Z(n44290) );
  XOR U44004 ( .A(n44217), .B(n44291), .Z(n44106) );
  AND U44005 ( .A(n1359), .B(n44292), .Z(n44291) );
  XOR U44006 ( .A(n44213), .B(n44217), .Z(n44292) );
  XNOR U44007 ( .A(n44293), .B(n44287), .Z(n44289) );
  IV U44008 ( .A(n44065), .Z(n44293) );
  XOR U44009 ( .A(n44294), .B(n44295), .Z(n44065) );
  AND U44010 ( .A(n1375), .B(n44296), .Z(n44295) );
  AND U44011 ( .A(n44258), .B(n44247), .Z(n44287) );
  XNOR U44012 ( .A(n44297), .B(n44298), .Z(n44247) );
  AND U44013 ( .A(n1359), .B(n44229), .Z(n44298) );
  XNOR U44014 ( .A(n44227), .B(n44297), .Z(n44229) );
  XNOR U44015 ( .A(n44299), .B(n44300), .Z(n1359) );
  AND U44016 ( .A(n44301), .B(n44302), .Z(n44300) );
  XNOR U44017 ( .A(n44299), .B(n44118), .Z(n44302) );
  IV U44018 ( .A(n44122), .Z(n44118) );
  XOR U44019 ( .A(n44303), .B(n44304), .Z(n44122) );
  AND U44020 ( .A(n1363), .B(n44305), .Z(n44304) );
  XOR U44021 ( .A(n44306), .B(n44303), .Z(n44305) );
  XNOR U44022 ( .A(n44299), .B(n44234), .Z(n44301) );
  XOR U44023 ( .A(n44307), .B(n44308), .Z(n44234) );
  AND U44024 ( .A(n1371), .B(n44269), .Z(n44308) );
  XOR U44025 ( .A(n44267), .B(n44307), .Z(n44269) );
  XOR U44026 ( .A(n44309), .B(n44310), .Z(n44299) );
  AND U44027 ( .A(n44311), .B(n44312), .Z(n44310) );
  XNOR U44028 ( .A(n44309), .B(n44134), .Z(n44312) );
  IV U44029 ( .A(n44137), .Z(n44134) );
  XOR U44030 ( .A(n44313), .B(n44314), .Z(n44137) );
  AND U44031 ( .A(n1363), .B(n44315), .Z(n44314) );
  XOR U44032 ( .A(n44316), .B(n44313), .Z(n44315) );
  XOR U44033 ( .A(n44138), .B(n44309), .Z(n44311) );
  XOR U44034 ( .A(n44317), .B(n44318), .Z(n44138) );
  AND U44035 ( .A(n1371), .B(n44277), .Z(n44318) );
  XOR U44036 ( .A(n44317), .B(n44275), .Z(n44277) );
  XOR U44037 ( .A(n44319), .B(n44320), .Z(n44309) );
  AND U44038 ( .A(n44321), .B(n44322), .Z(n44320) );
  XNOR U44039 ( .A(n44319), .B(n44162), .Z(n44322) );
  IV U44040 ( .A(n44165), .Z(n44162) );
  XOR U44041 ( .A(n44323), .B(n44324), .Z(n44165) );
  AND U44042 ( .A(n1363), .B(n44325), .Z(n44324) );
  XNOR U44043 ( .A(n44326), .B(n44323), .Z(n44325) );
  XOR U44044 ( .A(n44166), .B(n44319), .Z(n44321) );
  XOR U44045 ( .A(n44327), .B(n44328), .Z(n44166) );
  AND U44046 ( .A(n1371), .B(n44286), .Z(n44328) );
  XOR U44047 ( .A(n44327), .B(n44284), .Z(n44286) );
  XOR U44048 ( .A(n44243), .B(n44329), .Z(n44319) );
  AND U44049 ( .A(n44245), .B(n44330), .Z(n44329) );
  XNOR U44050 ( .A(n44243), .B(n44213), .Z(n44330) );
  IV U44051 ( .A(n44216), .Z(n44213) );
  XOR U44052 ( .A(n44331), .B(n44332), .Z(n44216) );
  AND U44053 ( .A(n1363), .B(n44333), .Z(n44332) );
  XOR U44054 ( .A(n44334), .B(n44331), .Z(n44333) );
  XOR U44055 ( .A(n44217), .B(n44243), .Z(n44245) );
  XOR U44056 ( .A(n44335), .B(n44336), .Z(n44217) );
  AND U44057 ( .A(n1371), .B(n44296), .Z(n44336) );
  XOR U44058 ( .A(n44335), .B(n44294), .Z(n44296) );
  AND U44059 ( .A(n44297), .B(n44227), .Z(n44243) );
  XNOR U44060 ( .A(n44337), .B(n44338), .Z(n44227) );
  AND U44061 ( .A(n1363), .B(n44339), .Z(n44338) );
  XNOR U44062 ( .A(n44340), .B(n44337), .Z(n44339) );
  XNOR U44063 ( .A(n44341), .B(n44342), .Z(n1363) );
  AND U44064 ( .A(n44343), .B(n44344), .Z(n44342) );
  XOR U44065 ( .A(n44306), .B(n44341), .Z(n44344) );
  AND U44066 ( .A(n44345), .B(n44346), .Z(n44306) );
  XNOR U44067 ( .A(n44303), .B(n44341), .Z(n44343) );
  XNOR U44068 ( .A(n44347), .B(n44348), .Z(n44303) );
  AND U44069 ( .A(n1367), .B(n44349), .Z(n44348) );
  XNOR U44070 ( .A(n44350), .B(n44351), .Z(n44349) );
  XOR U44071 ( .A(n44352), .B(n44353), .Z(n44341) );
  AND U44072 ( .A(n44354), .B(n44355), .Z(n44353) );
  XNOR U44073 ( .A(n44352), .B(n44345), .Z(n44355) );
  IV U44074 ( .A(n44316), .Z(n44345) );
  XOR U44075 ( .A(n44356), .B(n44357), .Z(n44316) );
  XOR U44076 ( .A(n44358), .B(n44346), .Z(n44357) );
  AND U44077 ( .A(n44326), .B(n44359), .Z(n44346) );
  AND U44078 ( .A(n44360), .B(n44361), .Z(n44358) );
  XOR U44079 ( .A(n44362), .B(n44356), .Z(n44360) );
  XNOR U44080 ( .A(n44313), .B(n44352), .Z(n44354) );
  XNOR U44081 ( .A(n44363), .B(n44364), .Z(n44313) );
  AND U44082 ( .A(n1367), .B(n44365), .Z(n44364) );
  XNOR U44083 ( .A(n44366), .B(n44367), .Z(n44365) );
  XOR U44084 ( .A(n44368), .B(n44369), .Z(n44352) );
  AND U44085 ( .A(n44370), .B(n44371), .Z(n44369) );
  XNOR U44086 ( .A(n44368), .B(n44326), .Z(n44371) );
  XOR U44087 ( .A(n44372), .B(n44361), .Z(n44326) );
  XNOR U44088 ( .A(n44373), .B(n44356), .Z(n44361) );
  XOR U44089 ( .A(n44374), .B(n44375), .Z(n44356) );
  AND U44090 ( .A(n44376), .B(n44377), .Z(n44375) );
  XOR U44091 ( .A(n44378), .B(n44374), .Z(n44376) );
  XNOR U44092 ( .A(n44379), .B(n44380), .Z(n44373) );
  AND U44093 ( .A(n44381), .B(n44382), .Z(n44380) );
  XOR U44094 ( .A(n44379), .B(n44383), .Z(n44381) );
  XNOR U44095 ( .A(n44362), .B(n44359), .Z(n44372) );
  AND U44096 ( .A(n44384), .B(n44385), .Z(n44359) );
  XOR U44097 ( .A(n44386), .B(n44387), .Z(n44362) );
  AND U44098 ( .A(n44388), .B(n44389), .Z(n44387) );
  XOR U44099 ( .A(n44386), .B(n44390), .Z(n44388) );
  XNOR U44100 ( .A(n44323), .B(n44368), .Z(n44370) );
  XNOR U44101 ( .A(n44391), .B(n44392), .Z(n44323) );
  AND U44102 ( .A(n1367), .B(n44393), .Z(n44392) );
  XNOR U44103 ( .A(n44394), .B(n44395), .Z(n44393) );
  XOR U44104 ( .A(n44396), .B(n44397), .Z(n44368) );
  AND U44105 ( .A(n44398), .B(n44399), .Z(n44397) );
  XNOR U44106 ( .A(n44396), .B(n44384), .Z(n44399) );
  IV U44107 ( .A(n44334), .Z(n44384) );
  XNOR U44108 ( .A(n44400), .B(n44377), .Z(n44334) );
  XNOR U44109 ( .A(n44401), .B(n44383), .Z(n44377) );
  XNOR U44110 ( .A(n44402), .B(n44403), .Z(n44383) );
  NOR U44111 ( .A(n44404), .B(n44405), .Z(n44403) );
  XOR U44112 ( .A(n44402), .B(n44406), .Z(n44404) );
  XNOR U44113 ( .A(n44382), .B(n44374), .Z(n44401) );
  XOR U44114 ( .A(n44407), .B(n44408), .Z(n44374) );
  AND U44115 ( .A(n44409), .B(n44410), .Z(n44408) );
  XOR U44116 ( .A(n44407), .B(n44411), .Z(n44409) );
  XNOR U44117 ( .A(n44412), .B(n44379), .Z(n44382) );
  XOR U44118 ( .A(n44413), .B(n44414), .Z(n44379) );
  AND U44119 ( .A(n44415), .B(n44416), .Z(n44414) );
  XNOR U44120 ( .A(n44417), .B(n44418), .Z(n44415) );
  IV U44121 ( .A(n44413), .Z(n44417) );
  XNOR U44122 ( .A(n44419), .B(n44420), .Z(n44412) );
  NOR U44123 ( .A(n44421), .B(n44422), .Z(n44420) );
  XNOR U44124 ( .A(n44419), .B(n44423), .Z(n44421) );
  XNOR U44125 ( .A(n44378), .B(n44385), .Z(n44400) );
  NOR U44126 ( .A(n44340), .B(n44424), .Z(n44385) );
  XOR U44127 ( .A(n44390), .B(n44389), .Z(n44378) );
  XNOR U44128 ( .A(n44425), .B(n44386), .Z(n44389) );
  XOR U44129 ( .A(n44426), .B(n44427), .Z(n44386) );
  AND U44130 ( .A(n44428), .B(n44429), .Z(n44427) );
  XNOR U44131 ( .A(n44430), .B(n44431), .Z(n44428) );
  IV U44132 ( .A(n44426), .Z(n44430) );
  XNOR U44133 ( .A(n44432), .B(n44433), .Z(n44425) );
  NOR U44134 ( .A(n44434), .B(n44435), .Z(n44433) );
  XNOR U44135 ( .A(n44432), .B(n44436), .Z(n44434) );
  XOR U44136 ( .A(n44437), .B(n44438), .Z(n44390) );
  NOR U44137 ( .A(n44439), .B(n44440), .Z(n44438) );
  XNOR U44138 ( .A(n44437), .B(n44441), .Z(n44439) );
  XNOR U44139 ( .A(n44331), .B(n44396), .Z(n44398) );
  XNOR U44140 ( .A(n44442), .B(n44443), .Z(n44331) );
  AND U44141 ( .A(n1367), .B(n44444), .Z(n44443) );
  XNOR U44142 ( .A(n44445), .B(n44446), .Z(n44444) );
  AND U44143 ( .A(n44337), .B(n44340), .Z(n44396) );
  XOR U44144 ( .A(n44447), .B(n44424), .Z(n44340) );
  XNOR U44145 ( .A(p_input[1088]), .B(p_input[2048]), .Z(n44424) );
  XNOR U44146 ( .A(n44411), .B(n44410), .Z(n44447) );
  XNOR U44147 ( .A(n44448), .B(n44418), .Z(n44410) );
  XNOR U44148 ( .A(n44406), .B(n44405), .Z(n44418) );
  XNOR U44149 ( .A(n44449), .B(n44402), .Z(n44405) );
  XNOR U44150 ( .A(p_input[1098]), .B(p_input[2058]), .Z(n44402) );
  XOR U44151 ( .A(p_input[1099]), .B(n29030), .Z(n44449) );
  XOR U44152 ( .A(p_input[1100]), .B(p_input[2060]), .Z(n44406) );
  XOR U44153 ( .A(n44416), .B(n44450), .Z(n44448) );
  IV U44154 ( .A(n44407), .Z(n44450) );
  XOR U44155 ( .A(p_input[1089]), .B(p_input[2049]), .Z(n44407) );
  XNOR U44156 ( .A(n44451), .B(n44423), .Z(n44416) );
  XNOR U44157 ( .A(p_input[1103]), .B(n29033), .Z(n44423) );
  XOR U44158 ( .A(n44413), .B(n44422), .Z(n44451) );
  XOR U44159 ( .A(n44452), .B(n44419), .Z(n44422) );
  XOR U44160 ( .A(p_input[1101]), .B(p_input[2061]), .Z(n44419) );
  XOR U44161 ( .A(p_input[1102]), .B(n29035), .Z(n44452) );
  XOR U44162 ( .A(p_input[1097]), .B(p_input[2057]), .Z(n44413) );
  XOR U44163 ( .A(n44431), .B(n44429), .Z(n44411) );
  XNOR U44164 ( .A(n44453), .B(n44436), .Z(n44429) );
  XOR U44165 ( .A(p_input[1096]), .B(p_input[2056]), .Z(n44436) );
  XOR U44166 ( .A(n44426), .B(n44435), .Z(n44453) );
  XOR U44167 ( .A(n44454), .B(n44432), .Z(n44435) );
  XOR U44168 ( .A(p_input[1094]), .B(p_input[2054]), .Z(n44432) );
  XOR U44169 ( .A(p_input[1095]), .B(n30404), .Z(n44454) );
  XOR U44170 ( .A(p_input[1090]), .B(p_input[2050]), .Z(n44426) );
  XNOR U44171 ( .A(n44441), .B(n44440), .Z(n44431) );
  XOR U44172 ( .A(n44455), .B(n44437), .Z(n44440) );
  XOR U44173 ( .A(p_input[1091]), .B(p_input[2051]), .Z(n44437) );
  XOR U44174 ( .A(p_input[1092]), .B(n30406), .Z(n44455) );
  XOR U44175 ( .A(p_input[1093]), .B(p_input[2053]), .Z(n44441) );
  XNOR U44176 ( .A(n44456), .B(n44457), .Z(n44337) );
  AND U44177 ( .A(n1367), .B(n44458), .Z(n44457) );
  XNOR U44178 ( .A(n44459), .B(n44460), .Z(n1367) );
  AND U44179 ( .A(n44461), .B(n44462), .Z(n44460) );
  XOR U44180 ( .A(n44351), .B(n44459), .Z(n44462) );
  XNOR U44181 ( .A(n44463), .B(n44459), .Z(n44461) );
  XOR U44182 ( .A(n44464), .B(n44465), .Z(n44459) );
  AND U44183 ( .A(n44466), .B(n44467), .Z(n44465) );
  XOR U44184 ( .A(n44366), .B(n44464), .Z(n44467) );
  XOR U44185 ( .A(n44464), .B(n44367), .Z(n44466) );
  XOR U44186 ( .A(n44468), .B(n44469), .Z(n44464) );
  AND U44187 ( .A(n44470), .B(n44471), .Z(n44469) );
  XOR U44188 ( .A(n44394), .B(n44468), .Z(n44471) );
  XOR U44189 ( .A(n44468), .B(n44395), .Z(n44470) );
  XOR U44190 ( .A(n44472), .B(n44473), .Z(n44468) );
  AND U44191 ( .A(n44474), .B(n44475), .Z(n44473) );
  XOR U44192 ( .A(n44472), .B(n44445), .Z(n44475) );
  XNOR U44193 ( .A(n44476), .B(n44477), .Z(n44297) );
  AND U44194 ( .A(n1371), .B(n44478), .Z(n44477) );
  XNOR U44195 ( .A(n44479), .B(n44480), .Z(n1371) );
  AND U44196 ( .A(n44481), .B(n44482), .Z(n44480) );
  XOR U44197 ( .A(n44479), .B(n44307), .Z(n44482) );
  XNOR U44198 ( .A(n44479), .B(n44267), .Z(n44481) );
  XOR U44199 ( .A(n44483), .B(n44484), .Z(n44479) );
  AND U44200 ( .A(n44485), .B(n44486), .Z(n44484) );
  XOR U44201 ( .A(n44483), .B(n44275), .Z(n44485) );
  XOR U44202 ( .A(n44487), .B(n44488), .Z(n44258) );
  AND U44203 ( .A(n1375), .B(n44478), .Z(n44488) );
  XNOR U44204 ( .A(n44476), .B(n44487), .Z(n44478) );
  XNOR U44205 ( .A(n44489), .B(n44490), .Z(n1375) );
  AND U44206 ( .A(n44491), .B(n44492), .Z(n44490) );
  XNOR U44207 ( .A(n44493), .B(n44489), .Z(n44492) );
  IV U44208 ( .A(n44307), .Z(n44493) );
  XOR U44209 ( .A(n44463), .B(n44494), .Z(n44307) );
  AND U44210 ( .A(n1378), .B(n44495), .Z(n44494) );
  XOR U44211 ( .A(n44350), .B(n44347), .Z(n44495) );
  IV U44212 ( .A(n44463), .Z(n44350) );
  XNOR U44213 ( .A(n44267), .B(n44489), .Z(n44491) );
  XOR U44214 ( .A(n44496), .B(n44497), .Z(n44267) );
  AND U44215 ( .A(n1394), .B(n44498), .Z(n44497) );
  XOR U44216 ( .A(n44483), .B(n44499), .Z(n44489) );
  AND U44217 ( .A(n44500), .B(n44486), .Z(n44499) );
  XNOR U44218 ( .A(n44317), .B(n44483), .Z(n44486) );
  XOR U44219 ( .A(n44367), .B(n44501), .Z(n44317) );
  AND U44220 ( .A(n1378), .B(n44502), .Z(n44501) );
  XOR U44221 ( .A(n44363), .B(n44367), .Z(n44502) );
  XNOR U44222 ( .A(n44503), .B(n44483), .Z(n44500) );
  IV U44223 ( .A(n44275), .Z(n44503) );
  XOR U44224 ( .A(n44504), .B(n44505), .Z(n44275) );
  AND U44225 ( .A(n1394), .B(n44506), .Z(n44505) );
  XOR U44226 ( .A(n44507), .B(n44508), .Z(n44483) );
  AND U44227 ( .A(n44509), .B(n44510), .Z(n44508) );
  XNOR U44228 ( .A(n44327), .B(n44507), .Z(n44510) );
  XOR U44229 ( .A(n44395), .B(n44511), .Z(n44327) );
  AND U44230 ( .A(n1378), .B(n44512), .Z(n44511) );
  XOR U44231 ( .A(n44391), .B(n44395), .Z(n44512) );
  XOR U44232 ( .A(n44507), .B(n44284), .Z(n44509) );
  XOR U44233 ( .A(n44513), .B(n44514), .Z(n44284) );
  AND U44234 ( .A(n1394), .B(n44515), .Z(n44514) );
  XOR U44235 ( .A(n44516), .B(n44517), .Z(n44507) );
  AND U44236 ( .A(n44518), .B(n44519), .Z(n44517) );
  XNOR U44237 ( .A(n44516), .B(n44335), .Z(n44519) );
  XOR U44238 ( .A(n44446), .B(n44520), .Z(n44335) );
  AND U44239 ( .A(n1378), .B(n44521), .Z(n44520) );
  XOR U44240 ( .A(n44442), .B(n44446), .Z(n44521) );
  XNOR U44241 ( .A(n44522), .B(n44516), .Z(n44518) );
  IV U44242 ( .A(n44294), .Z(n44522) );
  XOR U44243 ( .A(n44523), .B(n44524), .Z(n44294) );
  AND U44244 ( .A(n1394), .B(n44525), .Z(n44524) );
  AND U44245 ( .A(n44487), .B(n44476), .Z(n44516) );
  XNOR U44246 ( .A(n44526), .B(n44527), .Z(n44476) );
  AND U44247 ( .A(n1378), .B(n44458), .Z(n44527) );
  XNOR U44248 ( .A(n44456), .B(n44526), .Z(n44458) );
  XNOR U44249 ( .A(n44528), .B(n44529), .Z(n1378) );
  AND U44250 ( .A(n44530), .B(n44531), .Z(n44529) );
  XNOR U44251 ( .A(n44528), .B(n44347), .Z(n44531) );
  IV U44252 ( .A(n44351), .Z(n44347) );
  XOR U44253 ( .A(n44532), .B(n44533), .Z(n44351) );
  AND U44254 ( .A(n1382), .B(n44534), .Z(n44533) );
  XOR U44255 ( .A(n44535), .B(n44532), .Z(n44534) );
  XNOR U44256 ( .A(n44528), .B(n44463), .Z(n44530) );
  XOR U44257 ( .A(n44536), .B(n44537), .Z(n44463) );
  AND U44258 ( .A(n1390), .B(n44498), .Z(n44537) );
  XOR U44259 ( .A(n44496), .B(n44536), .Z(n44498) );
  XOR U44260 ( .A(n44538), .B(n44539), .Z(n44528) );
  AND U44261 ( .A(n44540), .B(n44541), .Z(n44539) );
  XNOR U44262 ( .A(n44538), .B(n44363), .Z(n44541) );
  IV U44263 ( .A(n44366), .Z(n44363) );
  XOR U44264 ( .A(n44542), .B(n44543), .Z(n44366) );
  AND U44265 ( .A(n1382), .B(n44544), .Z(n44543) );
  XOR U44266 ( .A(n44545), .B(n44542), .Z(n44544) );
  XOR U44267 ( .A(n44367), .B(n44538), .Z(n44540) );
  XOR U44268 ( .A(n44546), .B(n44547), .Z(n44367) );
  AND U44269 ( .A(n1390), .B(n44506), .Z(n44547) );
  XOR U44270 ( .A(n44546), .B(n44504), .Z(n44506) );
  XOR U44271 ( .A(n44548), .B(n44549), .Z(n44538) );
  AND U44272 ( .A(n44550), .B(n44551), .Z(n44549) );
  XNOR U44273 ( .A(n44548), .B(n44391), .Z(n44551) );
  IV U44274 ( .A(n44394), .Z(n44391) );
  XOR U44275 ( .A(n44552), .B(n44553), .Z(n44394) );
  AND U44276 ( .A(n1382), .B(n44554), .Z(n44553) );
  XNOR U44277 ( .A(n44555), .B(n44552), .Z(n44554) );
  XOR U44278 ( .A(n44395), .B(n44548), .Z(n44550) );
  XOR U44279 ( .A(n44556), .B(n44557), .Z(n44395) );
  AND U44280 ( .A(n1390), .B(n44515), .Z(n44557) );
  XOR U44281 ( .A(n44556), .B(n44513), .Z(n44515) );
  XOR U44282 ( .A(n44472), .B(n44558), .Z(n44548) );
  AND U44283 ( .A(n44474), .B(n44559), .Z(n44558) );
  XNOR U44284 ( .A(n44472), .B(n44442), .Z(n44559) );
  IV U44285 ( .A(n44445), .Z(n44442) );
  XOR U44286 ( .A(n44560), .B(n44561), .Z(n44445) );
  AND U44287 ( .A(n1382), .B(n44562), .Z(n44561) );
  XOR U44288 ( .A(n44563), .B(n44560), .Z(n44562) );
  XOR U44289 ( .A(n44446), .B(n44472), .Z(n44474) );
  XOR U44290 ( .A(n44564), .B(n44565), .Z(n44446) );
  AND U44291 ( .A(n1390), .B(n44525), .Z(n44565) );
  XOR U44292 ( .A(n44564), .B(n44523), .Z(n44525) );
  AND U44293 ( .A(n44526), .B(n44456), .Z(n44472) );
  XNOR U44294 ( .A(n44566), .B(n44567), .Z(n44456) );
  AND U44295 ( .A(n1382), .B(n44568), .Z(n44567) );
  XNOR U44296 ( .A(n44569), .B(n44566), .Z(n44568) );
  XNOR U44297 ( .A(n44570), .B(n44571), .Z(n1382) );
  AND U44298 ( .A(n44572), .B(n44573), .Z(n44571) );
  XOR U44299 ( .A(n44535), .B(n44570), .Z(n44573) );
  AND U44300 ( .A(n44574), .B(n44575), .Z(n44535) );
  XNOR U44301 ( .A(n44532), .B(n44570), .Z(n44572) );
  XNOR U44302 ( .A(n44576), .B(n44577), .Z(n44532) );
  AND U44303 ( .A(n1386), .B(n44578), .Z(n44577) );
  XNOR U44304 ( .A(n44579), .B(n44580), .Z(n44578) );
  XOR U44305 ( .A(n44581), .B(n44582), .Z(n44570) );
  AND U44306 ( .A(n44583), .B(n44584), .Z(n44582) );
  XNOR U44307 ( .A(n44581), .B(n44574), .Z(n44584) );
  IV U44308 ( .A(n44545), .Z(n44574) );
  XOR U44309 ( .A(n44585), .B(n44586), .Z(n44545) );
  XOR U44310 ( .A(n44587), .B(n44575), .Z(n44586) );
  AND U44311 ( .A(n44555), .B(n44588), .Z(n44575) );
  AND U44312 ( .A(n44589), .B(n44590), .Z(n44587) );
  XOR U44313 ( .A(n44591), .B(n44585), .Z(n44589) );
  XNOR U44314 ( .A(n44542), .B(n44581), .Z(n44583) );
  XNOR U44315 ( .A(n44592), .B(n44593), .Z(n44542) );
  AND U44316 ( .A(n1386), .B(n44594), .Z(n44593) );
  XNOR U44317 ( .A(n44595), .B(n44596), .Z(n44594) );
  XOR U44318 ( .A(n44597), .B(n44598), .Z(n44581) );
  AND U44319 ( .A(n44599), .B(n44600), .Z(n44598) );
  XNOR U44320 ( .A(n44597), .B(n44555), .Z(n44600) );
  XOR U44321 ( .A(n44601), .B(n44590), .Z(n44555) );
  XNOR U44322 ( .A(n44602), .B(n44585), .Z(n44590) );
  XOR U44323 ( .A(n44603), .B(n44604), .Z(n44585) );
  AND U44324 ( .A(n44605), .B(n44606), .Z(n44604) );
  XOR U44325 ( .A(n44607), .B(n44603), .Z(n44605) );
  XNOR U44326 ( .A(n44608), .B(n44609), .Z(n44602) );
  AND U44327 ( .A(n44610), .B(n44611), .Z(n44609) );
  XOR U44328 ( .A(n44608), .B(n44612), .Z(n44610) );
  XNOR U44329 ( .A(n44591), .B(n44588), .Z(n44601) );
  AND U44330 ( .A(n44613), .B(n44614), .Z(n44588) );
  XOR U44331 ( .A(n44615), .B(n44616), .Z(n44591) );
  AND U44332 ( .A(n44617), .B(n44618), .Z(n44616) );
  XOR U44333 ( .A(n44615), .B(n44619), .Z(n44617) );
  XNOR U44334 ( .A(n44552), .B(n44597), .Z(n44599) );
  XNOR U44335 ( .A(n44620), .B(n44621), .Z(n44552) );
  AND U44336 ( .A(n1386), .B(n44622), .Z(n44621) );
  XNOR U44337 ( .A(n44623), .B(n44624), .Z(n44622) );
  XOR U44338 ( .A(n44625), .B(n44626), .Z(n44597) );
  AND U44339 ( .A(n44627), .B(n44628), .Z(n44626) );
  XNOR U44340 ( .A(n44625), .B(n44613), .Z(n44628) );
  IV U44341 ( .A(n44563), .Z(n44613) );
  XNOR U44342 ( .A(n44629), .B(n44606), .Z(n44563) );
  XNOR U44343 ( .A(n44630), .B(n44612), .Z(n44606) );
  XNOR U44344 ( .A(n44631), .B(n44632), .Z(n44612) );
  NOR U44345 ( .A(n44633), .B(n44634), .Z(n44632) );
  XOR U44346 ( .A(n44631), .B(n44635), .Z(n44633) );
  XNOR U44347 ( .A(n44611), .B(n44603), .Z(n44630) );
  XOR U44348 ( .A(n44636), .B(n44637), .Z(n44603) );
  AND U44349 ( .A(n44638), .B(n44639), .Z(n44637) );
  XOR U44350 ( .A(n44636), .B(n44640), .Z(n44638) );
  XNOR U44351 ( .A(n44641), .B(n44608), .Z(n44611) );
  XOR U44352 ( .A(n44642), .B(n44643), .Z(n44608) );
  AND U44353 ( .A(n44644), .B(n44645), .Z(n44643) );
  XNOR U44354 ( .A(n44646), .B(n44647), .Z(n44644) );
  IV U44355 ( .A(n44642), .Z(n44646) );
  XNOR U44356 ( .A(n44648), .B(n44649), .Z(n44641) );
  NOR U44357 ( .A(n44650), .B(n44651), .Z(n44649) );
  XNOR U44358 ( .A(n44648), .B(n44652), .Z(n44650) );
  XNOR U44359 ( .A(n44607), .B(n44614), .Z(n44629) );
  NOR U44360 ( .A(n44569), .B(n44653), .Z(n44614) );
  XOR U44361 ( .A(n44619), .B(n44618), .Z(n44607) );
  XNOR U44362 ( .A(n44654), .B(n44615), .Z(n44618) );
  XOR U44363 ( .A(n44655), .B(n44656), .Z(n44615) );
  AND U44364 ( .A(n44657), .B(n44658), .Z(n44656) );
  XNOR U44365 ( .A(n44659), .B(n44660), .Z(n44657) );
  IV U44366 ( .A(n44655), .Z(n44659) );
  XNOR U44367 ( .A(n44661), .B(n44662), .Z(n44654) );
  NOR U44368 ( .A(n44663), .B(n44664), .Z(n44662) );
  XNOR U44369 ( .A(n44661), .B(n44665), .Z(n44663) );
  XOR U44370 ( .A(n44666), .B(n44667), .Z(n44619) );
  NOR U44371 ( .A(n44668), .B(n44669), .Z(n44667) );
  XNOR U44372 ( .A(n44666), .B(n44670), .Z(n44668) );
  XNOR U44373 ( .A(n44560), .B(n44625), .Z(n44627) );
  XNOR U44374 ( .A(n44671), .B(n44672), .Z(n44560) );
  AND U44375 ( .A(n1386), .B(n44673), .Z(n44672) );
  XNOR U44376 ( .A(n44674), .B(n44675), .Z(n44673) );
  AND U44377 ( .A(n44566), .B(n44569), .Z(n44625) );
  XOR U44378 ( .A(n44676), .B(n44653), .Z(n44569) );
  XNOR U44379 ( .A(p_input[1104]), .B(p_input[2048]), .Z(n44653) );
  XNOR U44380 ( .A(n44640), .B(n44639), .Z(n44676) );
  XNOR U44381 ( .A(n44677), .B(n44647), .Z(n44639) );
  XNOR U44382 ( .A(n44635), .B(n44634), .Z(n44647) );
  XNOR U44383 ( .A(n44678), .B(n44631), .Z(n44634) );
  XNOR U44384 ( .A(p_input[1114]), .B(p_input[2058]), .Z(n44631) );
  XOR U44385 ( .A(p_input[1115]), .B(n29030), .Z(n44678) );
  XOR U44386 ( .A(p_input[1116]), .B(p_input[2060]), .Z(n44635) );
  XOR U44387 ( .A(n44645), .B(n44679), .Z(n44677) );
  IV U44388 ( .A(n44636), .Z(n44679) );
  XOR U44389 ( .A(p_input[1105]), .B(p_input[2049]), .Z(n44636) );
  XNOR U44390 ( .A(n44680), .B(n44652), .Z(n44645) );
  XNOR U44391 ( .A(p_input[1119]), .B(n29033), .Z(n44652) );
  XOR U44392 ( .A(n44642), .B(n44651), .Z(n44680) );
  XOR U44393 ( .A(n44681), .B(n44648), .Z(n44651) );
  XOR U44394 ( .A(p_input[1117]), .B(p_input[2061]), .Z(n44648) );
  XOR U44395 ( .A(p_input[1118]), .B(n29035), .Z(n44681) );
  XOR U44396 ( .A(p_input[1113]), .B(p_input[2057]), .Z(n44642) );
  XOR U44397 ( .A(n44660), .B(n44658), .Z(n44640) );
  XNOR U44398 ( .A(n44682), .B(n44665), .Z(n44658) );
  XOR U44399 ( .A(p_input[1112]), .B(p_input[2056]), .Z(n44665) );
  XOR U44400 ( .A(n44655), .B(n44664), .Z(n44682) );
  XOR U44401 ( .A(n44683), .B(n44661), .Z(n44664) );
  XOR U44402 ( .A(p_input[1110]), .B(p_input[2054]), .Z(n44661) );
  XOR U44403 ( .A(p_input[1111]), .B(n30404), .Z(n44683) );
  XOR U44404 ( .A(p_input[1106]), .B(p_input[2050]), .Z(n44655) );
  XNOR U44405 ( .A(n44670), .B(n44669), .Z(n44660) );
  XOR U44406 ( .A(n44684), .B(n44666), .Z(n44669) );
  XOR U44407 ( .A(p_input[1107]), .B(p_input[2051]), .Z(n44666) );
  XOR U44408 ( .A(p_input[1108]), .B(n30406), .Z(n44684) );
  XOR U44409 ( .A(p_input[1109]), .B(p_input[2053]), .Z(n44670) );
  XNOR U44410 ( .A(n44685), .B(n44686), .Z(n44566) );
  AND U44411 ( .A(n1386), .B(n44687), .Z(n44686) );
  XNOR U44412 ( .A(n44688), .B(n44689), .Z(n1386) );
  AND U44413 ( .A(n44690), .B(n44691), .Z(n44689) );
  XOR U44414 ( .A(n44580), .B(n44688), .Z(n44691) );
  XNOR U44415 ( .A(n44692), .B(n44688), .Z(n44690) );
  XOR U44416 ( .A(n44693), .B(n44694), .Z(n44688) );
  AND U44417 ( .A(n44695), .B(n44696), .Z(n44694) );
  XOR U44418 ( .A(n44595), .B(n44693), .Z(n44696) );
  XOR U44419 ( .A(n44693), .B(n44596), .Z(n44695) );
  XOR U44420 ( .A(n44697), .B(n44698), .Z(n44693) );
  AND U44421 ( .A(n44699), .B(n44700), .Z(n44698) );
  XOR U44422 ( .A(n44623), .B(n44697), .Z(n44700) );
  XOR U44423 ( .A(n44697), .B(n44624), .Z(n44699) );
  XOR U44424 ( .A(n44701), .B(n44702), .Z(n44697) );
  AND U44425 ( .A(n44703), .B(n44704), .Z(n44702) );
  XOR U44426 ( .A(n44701), .B(n44674), .Z(n44704) );
  XNOR U44427 ( .A(n44705), .B(n44706), .Z(n44526) );
  AND U44428 ( .A(n1390), .B(n44707), .Z(n44706) );
  XNOR U44429 ( .A(n44708), .B(n44709), .Z(n1390) );
  AND U44430 ( .A(n44710), .B(n44711), .Z(n44709) );
  XOR U44431 ( .A(n44708), .B(n44536), .Z(n44711) );
  XNOR U44432 ( .A(n44708), .B(n44496), .Z(n44710) );
  XOR U44433 ( .A(n44712), .B(n44713), .Z(n44708) );
  AND U44434 ( .A(n44714), .B(n44715), .Z(n44713) );
  XOR U44435 ( .A(n44712), .B(n44504), .Z(n44714) );
  XOR U44436 ( .A(n44716), .B(n44717), .Z(n44487) );
  AND U44437 ( .A(n1394), .B(n44707), .Z(n44717) );
  XNOR U44438 ( .A(n44705), .B(n44716), .Z(n44707) );
  XNOR U44439 ( .A(n44718), .B(n44719), .Z(n1394) );
  AND U44440 ( .A(n44720), .B(n44721), .Z(n44719) );
  XNOR U44441 ( .A(n44722), .B(n44718), .Z(n44721) );
  IV U44442 ( .A(n44536), .Z(n44722) );
  XOR U44443 ( .A(n44692), .B(n44723), .Z(n44536) );
  AND U44444 ( .A(n1397), .B(n44724), .Z(n44723) );
  XOR U44445 ( .A(n44579), .B(n44576), .Z(n44724) );
  IV U44446 ( .A(n44692), .Z(n44579) );
  XNOR U44447 ( .A(n44496), .B(n44718), .Z(n44720) );
  XOR U44448 ( .A(n44725), .B(n44726), .Z(n44496) );
  AND U44449 ( .A(n1413), .B(n44727), .Z(n44726) );
  XOR U44450 ( .A(n44712), .B(n44728), .Z(n44718) );
  AND U44451 ( .A(n44729), .B(n44715), .Z(n44728) );
  XNOR U44452 ( .A(n44546), .B(n44712), .Z(n44715) );
  XOR U44453 ( .A(n44596), .B(n44730), .Z(n44546) );
  AND U44454 ( .A(n1397), .B(n44731), .Z(n44730) );
  XOR U44455 ( .A(n44592), .B(n44596), .Z(n44731) );
  XNOR U44456 ( .A(n44732), .B(n44712), .Z(n44729) );
  IV U44457 ( .A(n44504), .Z(n44732) );
  XOR U44458 ( .A(n44733), .B(n44734), .Z(n44504) );
  AND U44459 ( .A(n1413), .B(n44735), .Z(n44734) );
  XOR U44460 ( .A(n44736), .B(n44737), .Z(n44712) );
  AND U44461 ( .A(n44738), .B(n44739), .Z(n44737) );
  XNOR U44462 ( .A(n44556), .B(n44736), .Z(n44739) );
  XOR U44463 ( .A(n44624), .B(n44740), .Z(n44556) );
  AND U44464 ( .A(n1397), .B(n44741), .Z(n44740) );
  XOR U44465 ( .A(n44620), .B(n44624), .Z(n44741) );
  XOR U44466 ( .A(n44736), .B(n44513), .Z(n44738) );
  XOR U44467 ( .A(n44742), .B(n44743), .Z(n44513) );
  AND U44468 ( .A(n1413), .B(n44744), .Z(n44743) );
  XOR U44469 ( .A(n44745), .B(n44746), .Z(n44736) );
  AND U44470 ( .A(n44747), .B(n44748), .Z(n44746) );
  XNOR U44471 ( .A(n44745), .B(n44564), .Z(n44748) );
  XOR U44472 ( .A(n44675), .B(n44749), .Z(n44564) );
  AND U44473 ( .A(n1397), .B(n44750), .Z(n44749) );
  XOR U44474 ( .A(n44671), .B(n44675), .Z(n44750) );
  XNOR U44475 ( .A(n44751), .B(n44745), .Z(n44747) );
  IV U44476 ( .A(n44523), .Z(n44751) );
  XOR U44477 ( .A(n44752), .B(n44753), .Z(n44523) );
  AND U44478 ( .A(n1413), .B(n44754), .Z(n44753) );
  AND U44479 ( .A(n44716), .B(n44705), .Z(n44745) );
  XNOR U44480 ( .A(n44755), .B(n44756), .Z(n44705) );
  AND U44481 ( .A(n1397), .B(n44687), .Z(n44756) );
  XNOR U44482 ( .A(n44685), .B(n44755), .Z(n44687) );
  XNOR U44483 ( .A(n44757), .B(n44758), .Z(n1397) );
  AND U44484 ( .A(n44759), .B(n44760), .Z(n44758) );
  XNOR U44485 ( .A(n44757), .B(n44576), .Z(n44760) );
  IV U44486 ( .A(n44580), .Z(n44576) );
  XOR U44487 ( .A(n44761), .B(n44762), .Z(n44580) );
  AND U44488 ( .A(n1401), .B(n44763), .Z(n44762) );
  XOR U44489 ( .A(n44764), .B(n44761), .Z(n44763) );
  XNOR U44490 ( .A(n44757), .B(n44692), .Z(n44759) );
  XOR U44491 ( .A(n44765), .B(n44766), .Z(n44692) );
  AND U44492 ( .A(n1409), .B(n44727), .Z(n44766) );
  XOR U44493 ( .A(n44725), .B(n44765), .Z(n44727) );
  XOR U44494 ( .A(n44767), .B(n44768), .Z(n44757) );
  AND U44495 ( .A(n44769), .B(n44770), .Z(n44768) );
  XNOR U44496 ( .A(n44767), .B(n44592), .Z(n44770) );
  IV U44497 ( .A(n44595), .Z(n44592) );
  XOR U44498 ( .A(n44771), .B(n44772), .Z(n44595) );
  AND U44499 ( .A(n1401), .B(n44773), .Z(n44772) );
  XOR U44500 ( .A(n44774), .B(n44771), .Z(n44773) );
  XOR U44501 ( .A(n44596), .B(n44767), .Z(n44769) );
  XOR U44502 ( .A(n44775), .B(n44776), .Z(n44596) );
  AND U44503 ( .A(n1409), .B(n44735), .Z(n44776) );
  XOR U44504 ( .A(n44775), .B(n44733), .Z(n44735) );
  XOR U44505 ( .A(n44777), .B(n44778), .Z(n44767) );
  AND U44506 ( .A(n44779), .B(n44780), .Z(n44778) );
  XNOR U44507 ( .A(n44777), .B(n44620), .Z(n44780) );
  IV U44508 ( .A(n44623), .Z(n44620) );
  XOR U44509 ( .A(n44781), .B(n44782), .Z(n44623) );
  AND U44510 ( .A(n1401), .B(n44783), .Z(n44782) );
  XNOR U44511 ( .A(n44784), .B(n44781), .Z(n44783) );
  XOR U44512 ( .A(n44624), .B(n44777), .Z(n44779) );
  XOR U44513 ( .A(n44785), .B(n44786), .Z(n44624) );
  AND U44514 ( .A(n1409), .B(n44744), .Z(n44786) );
  XOR U44515 ( .A(n44785), .B(n44742), .Z(n44744) );
  XOR U44516 ( .A(n44701), .B(n44787), .Z(n44777) );
  AND U44517 ( .A(n44703), .B(n44788), .Z(n44787) );
  XNOR U44518 ( .A(n44701), .B(n44671), .Z(n44788) );
  IV U44519 ( .A(n44674), .Z(n44671) );
  XOR U44520 ( .A(n44789), .B(n44790), .Z(n44674) );
  AND U44521 ( .A(n1401), .B(n44791), .Z(n44790) );
  XOR U44522 ( .A(n44792), .B(n44789), .Z(n44791) );
  XOR U44523 ( .A(n44675), .B(n44701), .Z(n44703) );
  XOR U44524 ( .A(n44793), .B(n44794), .Z(n44675) );
  AND U44525 ( .A(n1409), .B(n44754), .Z(n44794) );
  XOR U44526 ( .A(n44793), .B(n44752), .Z(n44754) );
  AND U44527 ( .A(n44755), .B(n44685), .Z(n44701) );
  XNOR U44528 ( .A(n44795), .B(n44796), .Z(n44685) );
  AND U44529 ( .A(n1401), .B(n44797), .Z(n44796) );
  XNOR U44530 ( .A(n44798), .B(n44795), .Z(n44797) );
  XNOR U44531 ( .A(n44799), .B(n44800), .Z(n1401) );
  AND U44532 ( .A(n44801), .B(n44802), .Z(n44800) );
  XOR U44533 ( .A(n44764), .B(n44799), .Z(n44802) );
  AND U44534 ( .A(n44803), .B(n44804), .Z(n44764) );
  XNOR U44535 ( .A(n44761), .B(n44799), .Z(n44801) );
  XNOR U44536 ( .A(n44805), .B(n44806), .Z(n44761) );
  AND U44537 ( .A(n1405), .B(n44807), .Z(n44806) );
  XNOR U44538 ( .A(n44808), .B(n44809), .Z(n44807) );
  XOR U44539 ( .A(n44810), .B(n44811), .Z(n44799) );
  AND U44540 ( .A(n44812), .B(n44813), .Z(n44811) );
  XNOR U44541 ( .A(n44810), .B(n44803), .Z(n44813) );
  IV U44542 ( .A(n44774), .Z(n44803) );
  XOR U44543 ( .A(n44814), .B(n44815), .Z(n44774) );
  XOR U44544 ( .A(n44816), .B(n44804), .Z(n44815) );
  AND U44545 ( .A(n44784), .B(n44817), .Z(n44804) );
  AND U44546 ( .A(n44818), .B(n44819), .Z(n44816) );
  XOR U44547 ( .A(n44820), .B(n44814), .Z(n44818) );
  XNOR U44548 ( .A(n44771), .B(n44810), .Z(n44812) );
  XNOR U44549 ( .A(n44821), .B(n44822), .Z(n44771) );
  AND U44550 ( .A(n1405), .B(n44823), .Z(n44822) );
  XNOR U44551 ( .A(n44824), .B(n44825), .Z(n44823) );
  XOR U44552 ( .A(n44826), .B(n44827), .Z(n44810) );
  AND U44553 ( .A(n44828), .B(n44829), .Z(n44827) );
  XNOR U44554 ( .A(n44826), .B(n44784), .Z(n44829) );
  XOR U44555 ( .A(n44830), .B(n44819), .Z(n44784) );
  XNOR U44556 ( .A(n44831), .B(n44814), .Z(n44819) );
  XOR U44557 ( .A(n44832), .B(n44833), .Z(n44814) );
  AND U44558 ( .A(n44834), .B(n44835), .Z(n44833) );
  XOR U44559 ( .A(n44836), .B(n44832), .Z(n44834) );
  XNOR U44560 ( .A(n44837), .B(n44838), .Z(n44831) );
  AND U44561 ( .A(n44839), .B(n44840), .Z(n44838) );
  XOR U44562 ( .A(n44837), .B(n44841), .Z(n44839) );
  XNOR U44563 ( .A(n44820), .B(n44817), .Z(n44830) );
  AND U44564 ( .A(n44842), .B(n44843), .Z(n44817) );
  XOR U44565 ( .A(n44844), .B(n44845), .Z(n44820) );
  AND U44566 ( .A(n44846), .B(n44847), .Z(n44845) );
  XOR U44567 ( .A(n44844), .B(n44848), .Z(n44846) );
  XNOR U44568 ( .A(n44781), .B(n44826), .Z(n44828) );
  XNOR U44569 ( .A(n44849), .B(n44850), .Z(n44781) );
  AND U44570 ( .A(n1405), .B(n44851), .Z(n44850) );
  XNOR U44571 ( .A(n44852), .B(n44853), .Z(n44851) );
  XOR U44572 ( .A(n44854), .B(n44855), .Z(n44826) );
  AND U44573 ( .A(n44856), .B(n44857), .Z(n44855) );
  XNOR U44574 ( .A(n44854), .B(n44842), .Z(n44857) );
  IV U44575 ( .A(n44792), .Z(n44842) );
  XNOR U44576 ( .A(n44858), .B(n44835), .Z(n44792) );
  XNOR U44577 ( .A(n44859), .B(n44841), .Z(n44835) );
  XNOR U44578 ( .A(n44860), .B(n44861), .Z(n44841) );
  NOR U44579 ( .A(n44862), .B(n44863), .Z(n44861) );
  XOR U44580 ( .A(n44860), .B(n44864), .Z(n44862) );
  XNOR U44581 ( .A(n44840), .B(n44832), .Z(n44859) );
  XOR U44582 ( .A(n44865), .B(n44866), .Z(n44832) );
  AND U44583 ( .A(n44867), .B(n44868), .Z(n44866) );
  XOR U44584 ( .A(n44865), .B(n44869), .Z(n44867) );
  XNOR U44585 ( .A(n44870), .B(n44837), .Z(n44840) );
  XOR U44586 ( .A(n44871), .B(n44872), .Z(n44837) );
  AND U44587 ( .A(n44873), .B(n44874), .Z(n44872) );
  XNOR U44588 ( .A(n44875), .B(n44876), .Z(n44873) );
  IV U44589 ( .A(n44871), .Z(n44875) );
  XNOR U44590 ( .A(n44877), .B(n44878), .Z(n44870) );
  NOR U44591 ( .A(n44879), .B(n44880), .Z(n44878) );
  XNOR U44592 ( .A(n44877), .B(n44881), .Z(n44879) );
  XNOR U44593 ( .A(n44836), .B(n44843), .Z(n44858) );
  NOR U44594 ( .A(n44798), .B(n44882), .Z(n44843) );
  XOR U44595 ( .A(n44848), .B(n44847), .Z(n44836) );
  XNOR U44596 ( .A(n44883), .B(n44844), .Z(n44847) );
  XOR U44597 ( .A(n44884), .B(n44885), .Z(n44844) );
  AND U44598 ( .A(n44886), .B(n44887), .Z(n44885) );
  XNOR U44599 ( .A(n44888), .B(n44889), .Z(n44886) );
  IV U44600 ( .A(n44884), .Z(n44888) );
  XNOR U44601 ( .A(n44890), .B(n44891), .Z(n44883) );
  NOR U44602 ( .A(n44892), .B(n44893), .Z(n44891) );
  XNOR U44603 ( .A(n44890), .B(n44894), .Z(n44892) );
  XOR U44604 ( .A(n44895), .B(n44896), .Z(n44848) );
  NOR U44605 ( .A(n44897), .B(n44898), .Z(n44896) );
  XNOR U44606 ( .A(n44895), .B(n44899), .Z(n44897) );
  XNOR U44607 ( .A(n44789), .B(n44854), .Z(n44856) );
  XNOR U44608 ( .A(n44900), .B(n44901), .Z(n44789) );
  AND U44609 ( .A(n1405), .B(n44902), .Z(n44901) );
  XNOR U44610 ( .A(n44903), .B(n44904), .Z(n44902) );
  AND U44611 ( .A(n44795), .B(n44798), .Z(n44854) );
  XOR U44612 ( .A(n44905), .B(n44882), .Z(n44798) );
  XNOR U44613 ( .A(p_input[1120]), .B(p_input[2048]), .Z(n44882) );
  XNOR U44614 ( .A(n44869), .B(n44868), .Z(n44905) );
  XNOR U44615 ( .A(n44906), .B(n44876), .Z(n44868) );
  XNOR U44616 ( .A(n44864), .B(n44863), .Z(n44876) );
  XNOR U44617 ( .A(n44907), .B(n44860), .Z(n44863) );
  XNOR U44618 ( .A(p_input[1130]), .B(p_input[2058]), .Z(n44860) );
  XOR U44619 ( .A(p_input[1131]), .B(n29030), .Z(n44907) );
  XOR U44620 ( .A(p_input[1132]), .B(p_input[2060]), .Z(n44864) );
  XOR U44621 ( .A(n44874), .B(n44908), .Z(n44906) );
  IV U44622 ( .A(n44865), .Z(n44908) );
  XOR U44623 ( .A(p_input[1121]), .B(p_input[2049]), .Z(n44865) );
  XNOR U44624 ( .A(n44909), .B(n44881), .Z(n44874) );
  XNOR U44625 ( .A(p_input[1135]), .B(n29033), .Z(n44881) );
  XOR U44626 ( .A(n44871), .B(n44880), .Z(n44909) );
  XOR U44627 ( .A(n44910), .B(n44877), .Z(n44880) );
  XOR U44628 ( .A(p_input[1133]), .B(p_input[2061]), .Z(n44877) );
  XOR U44629 ( .A(p_input[1134]), .B(n29035), .Z(n44910) );
  XOR U44630 ( .A(p_input[1129]), .B(p_input[2057]), .Z(n44871) );
  XOR U44631 ( .A(n44889), .B(n44887), .Z(n44869) );
  XNOR U44632 ( .A(n44911), .B(n44894), .Z(n44887) );
  XOR U44633 ( .A(p_input[1128]), .B(p_input[2056]), .Z(n44894) );
  XOR U44634 ( .A(n44884), .B(n44893), .Z(n44911) );
  XOR U44635 ( .A(n44912), .B(n44890), .Z(n44893) );
  XOR U44636 ( .A(p_input[1126]), .B(p_input[2054]), .Z(n44890) );
  XOR U44637 ( .A(p_input[1127]), .B(n30404), .Z(n44912) );
  XOR U44638 ( .A(p_input[1122]), .B(p_input[2050]), .Z(n44884) );
  XNOR U44639 ( .A(n44899), .B(n44898), .Z(n44889) );
  XOR U44640 ( .A(n44913), .B(n44895), .Z(n44898) );
  XOR U44641 ( .A(p_input[1123]), .B(p_input[2051]), .Z(n44895) );
  XOR U44642 ( .A(p_input[1124]), .B(n30406), .Z(n44913) );
  XOR U44643 ( .A(p_input[1125]), .B(p_input[2053]), .Z(n44899) );
  XNOR U44644 ( .A(n44914), .B(n44915), .Z(n44795) );
  AND U44645 ( .A(n1405), .B(n44916), .Z(n44915) );
  XNOR U44646 ( .A(n44917), .B(n44918), .Z(n1405) );
  AND U44647 ( .A(n44919), .B(n44920), .Z(n44918) );
  XOR U44648 ( .A(n44809), .B(n44917), .Z(n44920) );
  XNOR U44649 ( .A(n44921), .B(n44917), .Z(n44919) );
  XOR U44650 ( .A(n44922), .B(n44923), .Z(n44917) );
  AND U44651 ( .A(n44924), .B(n44925), .Z(n44923) );
  XOR U44652 ( .A(n44824), .B(n44922), .Z(n44925) );
  XOR U44653 ( .A(n44922), .B(n44825), .Z(n44924) );
  XOR U44654 ( .A(n44926), .B(n44927), .Z(n44922) );
  AND U44655 ( .A(n44928), .B(n44929), .Z(n44927) );
  XOR U44656 ( .A(n44852), .B(n44926), .Z(n44929) );
  XOR U44657 ( .A(n44926), .B(n44853), .Z(n44928) );
  XOR U44658 ( .A(n44930), .B(n44931), .Z(n44926) );
  AND U44659 ( .A(n44932), .B(n44933), .Z(n44931) );
  XOR U44660 ( .A(n44930), .B(n44903), .Z(n44933) );
  XNOR U44661 ( .A(n44934), .B(n44935), .Z(n44755) );
  AND U44662 ( .A(n1409), .B(n44936), .Z(n44935) );
  XNOR U44663 ( .A(n44937), .B(n44938), .Z(n1409) );
  AND U44664 ( .A(n44939), .B(n44940), .Z(n44938) );
  XOR U44665 ( .A(n44937), .B(n44765), .Z(n44940) );
  XNOR U44666 ( .A(n44937), .B(n44725), .Z(n44939) );
  XOR U44667 ( .A(n44941), .B(n44942), .Z(n44937) );
  AND U44668 ( .A(n44943), .B(n44944), .Z(n44942) );
  XOR U44669 ( .A(n44941), .B(n44733), .Z(n44943) );
  XOR U44670 ( .A(n44945), .B(n44946), .Z(n44716) );
  AND U44671 ( .A(n1413), .B(n44936), .Z(n44946) );
  XNOR U44672 ( .A(n44934), .B(n44945), .Z(n44936) );
  XNOR U44673 ( .A(n44947), .B(n44948), .Z(n1413) );
  AND U44674 ( .A(n44949), .B(n44950), .Z(n44948) );
  XNOR U44675 ( .A(n44951), .B(n44947), .Z(n44950) );
  IV U44676 ( .A(n44765), .Z(n44951) );
  XOR U44677 ( .A(n44921), .B(n44952), .Z(n44765) );
  AND U44678 ( .A(n1416), .B(n44953), .Z(n44952) );
  XOR U44679 ( .A(n44808), .B(n44805), .Z(n44953) );
  IV U44680 ( .A(n44921), .Z(n44808) );
  XNOR U44681 ( .A(n44725), .B(n44947), .Z(n44949) );
  XOR U44682 ( .A(n44954), .B(n44955), .Z(n44725) );
  AND U44683 ( .A(n1432), .B(n44956), .Z(n44955) );
  XOR U44684 ( .A(n44941), .B(n44957), .Z(n44947) );
  AND U44685 ( .A(n44958), .B(n44944), .Z(n44957) );
  XNOR U44686 ( .A(n44775), .B(n44941), .Z(n44944) );
  XOR U44687 ( .A(n44825), .B(n44959), .Z(n44775) );
  AND U44688 ( .A(n1416), .B(n44960), .Z(n44959) );
  XOR U44689 ( .A(n44821), .B(n44825), .Z(n44960) );
  XNOR U44690 ( .A(n44961), .B(n44941), .Z(n44958) );
  IV U44691 ( .A(n44733), .Z(n44961) );
  XOR U44692 ( .A(n44962), .B(n44963), .Z(n44733) );
  AND U44693 ( .A(n1432), .B(n44964), .Z(n44963) );
  XOR U44694 ( .A(n44965), .B(n44966), .Z(n44941) );
  AND U44695 ( .A(n44967), .B(n44968), .Z(n44966) );
  XNOR U44696 ( .A(n44785), .B(n44965), .Z(n44968) );
  XOR U44697 ( .A(n44853), .B(n44969), .Z(n44785) );
  AND U44698 ( .A(n1416), .B(n44970), .Z(n44969) );
  XOR U44699 ( .A(n44849), .B(n44853), .Z(n44970) );
  XOR U44700 ( .A(n44965), .B(n44742), .Z(n44967) );
  XOR U44701 ( .A(n44971), .B(n44972), .Z(n44742) );
  AND U44702 ( .A(n1432), .B(n44973), .Z(n44972) );
  XOR U44703 ( .A(n44974), .B(n44975), .Z(n44965) );
  AND U44704 ( .A(n44976), .B(n44977), .Z(n44975) );
  XNOR U44705 ( .A(n44974), .B(n44793), .Z(n44977) );
  XOR U44706 ( .A(n44904), .B(n44978), .Z(n44793) );
  AND U44707 ( .A(n1416), .B(n44979), .Z(n44978) );
  XOR U44708 ( .A(n44900), .B(n44904), .Z(n44979) );
  XNOR U44709 ( .A(n44980), .B(n44974), .Z(n44976) );
  IV U44710 ( .A(n44752), .Z(n44980) );
  XOR U44711 ( .A(n44981), .B(n44982), .Z(n44752) );
  AND U44712 ( .A(n1432), .B(n44983), .Z(n44982) );
  AND U44713 ( .A(n44945), .B(n44934), .Z(n44974) );
  XNOR U44714 ( .A(n44984), .B(n44985), .Z(n44934) );
  AND U44715 ( .A(n1416), .B(n44916), .Z(n44985) );
  XNOR U44716 ( .A(n44914), .B(n44984), .Z(n44916) );
  XNOR U44717 ( .A(n44986), .B(n44987), .Z(n1416) );
  AND U44718 ( .A(n44988), .B(n44989), .Z(n44987) );
  XNOR U44719 ( .A(n44986), .B(n44805), .Z(n44989) );
  IV U44720 ( .A(n44809), .Z(n44805) );
  XOR U44721 ( .A(n44990), .B(n44991), .Z(n44809) );
  AND U44722 ( .A(n1420), .B(n44992), .Z(n44991) );
  XOR U44723 ( .A(n44993), .B(n44990), .Z(n44992) );
  XNOR U44724 ( .A(n44986), .B(n44921), .Z(n44988) );
  XOR U44725 ( .A(n44994), .B(n44995), .Z(n44921) );
  AND U44726 ( .A(n1428), .B(n44956), .Z(n44995) );
  XOR U44727 ( .A(n44954), .B(n44994), .Z(n44956) );
  XOR U44728 ( .A(n44996), .B(n44997), .Z(n44986) );
  AND U44729 ( .A(n44998), .B(n44999), .Z(n44997) );
  XNOR U44730 ( .A(n44996), .B(n44821), .Z(n44999) );
  IV U44731 ( .A(n44824), .Z(n44821) );
  XOR U44732 ( .A(n45000), .B(n45001), .Z(n44824) );
  AND U44733 ( .A(n1420), .B(n45002), .Z(n45001) );
  XOR U44734 ( .A(n45003), .B(n45000), .Z(n45002) );
  XOR U44735 ( .A(n44825), .B(n44996), .Z(n44998) );
  XOR U44736 ( .A(n45004), .B(n45005), .Z(n44825) );
  AND U44737 ( .A(n1428), .B(n44964), .Z(n45005) );
  XOR U44738 ( .A(n45004), .B(n44962), .Z(n44964) );
  XOR U44739 ( .A(n45006), .B(n45007), .Z(n44996) );
  AND U44740 ( .A(n45008), .B(n45009), .Z(n45007) );
  XNOR U44741 ( .A(n45006), .B(n44849), .Z(n45009) );
  IV U44742 ( .A(n44852), .Z(n44849) );
  XOR U44743 ( .A(n45010), .B(n45011), .Z(n44852) );
  AND U44744 ( .A(n1420), .B(n45012), .Z(n45011) );
  XNOR U44745 ( .A(n45013), .B(n45010), .Z(n45012) );
  XOR U44746 ( .A(n44853), .B(n45006), .Z(n45008) );
  XOR U44747 ( .A(n45014), .B(n45015), .Z(n44853) );
  AND U44748 ( .A(n1428), .B(n44973), .Z(n45015) );
  XOR U44749 ( .A(n45014), .B(n44971), .Z(n44973) );
  XOR U44750 ( .A(n44930), .B(n45016), .Z(n45006) );
  AND U44751 ( .A(n44932), .B(n45017), .Z(n45016) );
  XNOR U44752 ( .A(n44930), .B(n44900), .Z(n45017) );
  IV U44753 ( .A(n44903), .Z(n44900) );
  XOR U44754 ( .A(n45018), .B(n45019), .Z(n44903) );
  AND U44755 ( .A(n1420), .B(n45020), .Z(n45019) );
  XOR U44756 ( .A(n45021), .B(n45018), .Z(n45020) );
  XOR U44757 ( .A(n44904), .B(n44930), .Z(n44932) );
  XOR U44758 ( .A(n45022), .B(n45023), .Z(n44904) );
  AND U44759 ( .A(n1428), .B(n44983), .Z(n45023) );
  XOR U44760 ( .A(n45022), .B(n44981), .Z(n44983) );
  AND U44761 ( .A(n44984), .B(n44914), .Z(n44930) );
  XNOR U44762 ( .A(n45024), .B(n45025), .Z(n44914) );
  AND U44763 ( .A(n1420), .B(n45026), .Z(n45025) );
  XNOR U44764 ( .A(n45027), .B(n45024), .Z(n45026) );
  XNOR U44765 ( .A(n45028), .B(n45029), .Z(n1420) );
  AND U44766 ( .A(n45030), .B(n45031), .Z(n45029) );
  XOR U44767 ( .A(n44993), .B(n45028), .Z(n45031) );
  AND U44768 ( .A(n45032), .B(n45033), .Z(n44993) );
  XNOR U44769 ( .A(n44990), .B(n45028), .Z(n45030) );
  XNOR U44770 ( .A(n45034), .B(n45035), .Z(n44990) );
  AND U44771 ( .A(n1424), .B(n45036), .Z(n45035) );
  XNOR U44772 ( .A(n45037), .B(n45038), .Z(n45036) );
  XOR U44773 ( .A(n45039), .B(n45040), .Z(n45028) );
  AND U44774 ( .A(n45041), .B(n45042), .Z(n45040) );
  XNOR U44775 ( .A(n45039), .B(n45032), .Z(n45042) );
  IV U44776 ( .A(n45003), .Z(n45032) );
  XOR U44777 ( .A(n45043), .B(n45044), .Z(n45003) );
  XOR U44778 ( .A(n45045), .B(n45033), .Z(n45044) );
  AND U44779 ( .A(n45013), .B(n45046), .Z(n45033) );
  AND U44780 ( .A(n45047), .B(n45048), .Z(n45045) );
  XOR U44781 ( .A(n45049), .B(n45043), .Z(n45047) );
  XNOR U44782 ( .A(n45000), .B(n45039), .Z(n45041) );
  XNOR U44783 ( .A(n45050), .B(n45051), .Z(n45000) );
  AND U44784 ( .A(n1424), .B(n45052), .Z(n45051) );
  XNOR U44785 ( .A(n45053), .B(n45054), .Z(n45052) );
  XOR U44786 ( .A(n45055), .B(n45056), .Z(n45039) );
  AND U44787 ( .A(n45057), .B(n45058), .Z(n45056) );
  XNOR U44788 ( .A(n45055), .B(n45013), .Z(n45058) );
  XOR U44789 ( .A(n45059), .B(n45048), .Z(n45013) );
  XNOR U44790 ( .A(n45060), .B(n45043), .Z(n45048) );
  XOR U44791 ( .A(n45061), .B(n45062), .Z(n45043) );
  AND U44792 ( .A(n45063), .B(n45064), .Z(n45062) );
  XOR U44793 ( .A(n45065), .B(n45061), .Z(n45063) );
  XNOR U44794 ( .A(n45066), .B(n45067), .Z(n45060) );
  AND U44795 ( .A(n45068), .B(n45069), .Z(n45067) );
  XOR U44796 ( .A(n45066), .B(n45070), .Z(n45068) );
  XNOR U44797 ( .A(n45049), .B(n45046), .Z(n45059) );
  AND U44798 ( .A(n45071), .B(n45072), .Z(n45046) );
  XOR U44799 ( .A(n45073), .B(n45074), .Z(n45049) );
  AND U44800 ( .A(n45075), .B(n45076), .Z(n45074) );
  XOR U44801 ( .A(n45073), .B(n45077), .Z(n45075) );
  XNOR U44802 ( .A(n45010), .B(n45055), .Z(n45057) );
  XNOR U44803 ( .A(n45078), .B(n45079), .Z(n45010) );
  AND U44804 ( .A(n1424), .B(n45080), .Z(n45079) );
  XNOR U44805 ( .A(n45081), .B(n45082), .Z(n45080) );
  XOR U44806 ( .A(n45083), .B(n45084), .Z(n45055) );
  AND U44807 ( .A(n45085), .B(n45086), .Z(n45084) );
  XNOR U44808 ( .A(n45083), .B(n45071), .Z(n45086) );
  IV U44809 ( .A(n45021), .Z(n45071) );
  XNOR U44810 ( .A(n45087), .B(n45064), .Z(n45021) );
  XNOR U44811 ( .A(n45088), .B(n45070), .Z(n45064) );
  XNOR U44812 ( .A(n45089), .B(n45090), .Z(n45070) );
  NOR U44813 ( .A(n45091), .B(n45092), .Z(n45090) );
  XOR U44814 ( .A(n45089), .B(n45093), .Z(n45091) );
  XNOR U44815 ( .A(n45069), .B(n45061), .Z(n45088) );
  XOR U44816 ( .A(n45094), .B(n45095), .Z(n45061) );
  AND U44817 ( .A(n45096), .B(n45097), .Z(n45095) );
  XOR U44818 ( .A(n45094), .B(n45098), .Z(n45096) );
  XNOR U44819 ( .A(n45099), .B(n45066), .Z(n45069) );
  XOR U44820 ( .A(n45100), .B(n45101), .Z(n45066) );
  AND U44821 ( .A(n45102), .B(n45103), .Z(n45101) );
  XNOR U44822 ( .A(n45104), .B(n45105), .Z(n45102) );
  IV U44823 ( .A(n45100), .Z(n45104) );
  XNOR U44824 ( .A(n45106), .B(n45107), .Z(n45099) );
  NOR U44825 ( .A(n45108), .B(n45109), .Z(n45107) );
  XNOR U44826 ( .A(n45106), .B(n45110), .Z(n45108) );
  XNOR U44827 ( .A(n45065), .B(n45072), .Z(n45087) );
  NOR U44828 ( .A(n45027), .B(n45111), .Z(n45072) );
  XOR U44829 ( .A(n45077), .B(n45076), .Z(n45065) );
  XNOR U44830 ( .A(n45112), .B(n45073), .Z(n45076) );
  XOR U44831 ( .A(n45113), .B(n45114), .Z(n45073) );
  AND U44832 ( .A(n45115), .B(n45116), .Z(n45114) );
  XNOR U44833 ( .A(n45117), .B(n45118), .Z(n45115) );
  IV U44834 ( .A(n45113), .Z(n45117) );
  XNOR U44835 ( .A(n45119), .B(n45120), .Z(n45112) );
  NOR U44836 ( .A(n45121), .B(n45122), .Z(n45120) );
  XNOR U44837 ( .A(n45119), .B(n45123), .Z(n45121) );
  XOR U44838 ( .A(n45124), .B(n45125), .Z(n45077) );
  NOR U44839 ( .A(n45126), .B(n45127), .Z(n45125) );
  XNOR U44840 ( .A(n45124), .B(n45128), .Z(n45126) );
  XNOR U44841 ( .A(n45018), .B(n45083), .Z(n45085) );
  XNOR U44842 ( .A(n45129), .B(n45130), .Z(n45018) );
  AND U44843 ( .A(n1424), .B(n45131), .Z(n45130) );
  XNOR U44844 ( .A(n45132), .B(n45133), .Z(n45131) );
  AND U44845 ( .A(n45024), .B(n45027), .Z(n45083) );
  XOR U44846 ( .A(n45134), .B(n45111), .Z(n45027) );
  XNOR U44847 ( .A(p_input[1136]), .B(p_input[2048]), .Z(n45111) );
  XNOR U44848 ( .A(n45098), .B(n45097), .Z(n45134) );
  XNOR U44849 ( .A(n45135), .B(n45105), .Z(n45097) );
  XNOR U44850 ( .A(n45093), .B(n45092), .Z(n45105) );
  XNOR U44851 ( .A(n45136), .B(n45089), .Z(n45092) );
  XNOR U44852 ( .A(p_input[1146]), .B(p_input[2058]), .Z(n45089) );
  XOR U44853 ( .A(p_input[1147]), .B(n29030), .Z(n45136) );
  XOR U44854 ( .A(p_input[1148]), .B(p_input[2060]), .Z(n45093) );
  XOR U44855 ( .A(n45103), .B(n45137), .Z(n45135) );
  IV U44856 ( .A(n45094), .Z(n45137) );
  XOR U44857 ( .A(p_input[1137]), .B(p_input[2049]), .Z(n45094) );
  XNOR U44858 ( .A(n45138), .B(n45110), .Z(n45103) );
  XNOR U44859 ( .A(p_input[1151]), .B(n29033), .Z(n45110) );
  XOR U44860 ( .A(n45100), .B(n45109), .Z(n45138) );
  XOR U44861 ( .A(n45139), .B(n45106), .Z(n45109) );
  XOR U44862 ( .A(p_input[1149]), .B(p_input[2061]), .Z(n45106) );
  XOR U44863 ( .A(p_input[1150]), .B(n29035), .Z(n45139) );
  XOR U44864 ( .A(p_input[1145]), .B(p_input[2057]), .Z(n45100) );
  XOR U44865 ( .A(n45118), .B(n45116), .Z(n45098) );
  XNOR U44866 ( .A(n45140), .B(n45123), .Z(n45116) );
  XOR U44867 ( .A(p_input[1144]), .B(p_input[2056]), .Z(n45123) );
  XOR U44868 ( .A(n45113), .B(n45122), .Z(n45140) );
  XOR U44869 ( .A(n45141), .B(n45119), .Z(n45122) );
  XOR U44870 ( .A(p_input[1142]), .B(p_input[2054]), .Z(n45119) );
  XOR U44871 ( .A(p_input[1143]), .B(n30404), .Z(n45141) );
  XOR U44872 ( .A(p_input[1138]), .B(p_input[2050]), .Z(n45113) );
  XNOR U44873 ( .A(n45128), .B(n45127), .Z(n45118) );
  XOR U44874 ( .A(n45142), .B(n45124), .Z(n45127) );
  XOR U44875 ( .A(p_input[1139]), .B(p_input[2051]), .Z(n45124) );
  XOR U44876 ( .A(p_input[1140]), .B(n30406), .Z(n45142) );
  XOR U44877 ( .A(p_input[1141]), .B(p_input[2053]), .Z(n45128) );
  XNOR U44878 ( .A(n45143), .B(n45144), .Z(n45024) );
  AND U44879 ( .A(n1424), .B(n45145), .Z(n45144) );
  XNOR U44880 ( .A(n45146), .B(n45147), .Z(n1424) );
  AND U44881 ( .A(n45148), .B(n45149), .Z(n45147) );
  XOR U44882 ( .A(n45038), .B(n45146), .Z(n45149) );
  XNOR U44883 ( .A(n45150), .B(n45146), .Z(n45148) );
  XOR U44884 ( .A(n45151), .B(n45152), .Z(n45146) );
  AND U44885 ( .A(n45153), .B(n45154), .Z(n45152) );
  XOR U44886 ( .A(n45053), .B(n45151), .Z(n45154) );
  XOR U44887 ( .A(n45151), .B(n45054), .Z(n45153) );
  XOR U44888 ( .A(n45155), .B(n45156), .Z(n45151) );
  AND U44889 ( .A(n45157), .B(n45158), .Z(n45156) );
  XOR U44890 ( .A(n45081), .B(n45155), .Z(n45158) );
  XOR U44891 ( .A(n45155), .B(n45082), .Z(n45157) );
  XOR U44892 ( .A(n45159), .B(n45160), .Z(n45155) );
  AND U44893 ( .A(n45161), .B(n45162), .Z(n45160) );
  XOR U44894 ( .A(n45159), .B(n45132), .Z(n45162) );
  XNOR U44895 ( .A(n45163), .B(n45164), .Z(n44984) );
  AND U44896 ( .A(n1428), .B(n45165), .Z(n45164) );
  XNOR U44897 ( .A(n45166), .B(n45167), .Z(n1428) );
  AND U44898 ( .A(n45168), .B(n45169), .Z(n45167) );
  XOR U44899 ( .A(n45166), .B(n44994), .Z(n45169) );
  XNOR U44900 ( .A(n45166), .B(n44954), .Z(n45168) );
  XOR U44901 ( .A(n45170), .B(n45171), .Z(n45166) );
  AND U44902 ( .A(n45172), .B(n45173), .Z(n45171) );
  XOR U44903 ( .A(n45170), .B(n44962), .Z(n45172) );
  XOR U44904 ( .A(n45174), .B(n45175), .Z(n44945) );
  AND U44905 ( .A(n1432), .B(n45165), .Z(n45175) );
  XNOR U44906 ( .A(n45163), .B(n45174), .Z(n45165) );
  XNOR U44907 ( .A(n45176), .B(n45177), .Z(n1432) );
  AND U44908 ( .A(n45178), .B(n45179), .Z(n45177) );
  XNOR U44909 ( .A(n45180), .B(n45176), .Z(n45179) );
  IV U44910 ( .A(n44994), .Z(n45180) );
  XOR U44911 ( .A(n45150), .B(n45181), .Z(n44994) );
  AND U44912 ( .A(n1435), .B(n45182), .Z(n45181) );
  XOR U44913 ( .A(n45037), .B(n45034), .Z(n45182) );
  IV U44914 ( .A(n45150), .Z(n45037) );
  XNOR U44915 ( .A(n44954), .B(n45176), .Z(n45178) );
  XOR U44916 ( .A(n45183), .B(n45184), .Z(n44954) );
  AND U44917 ( .A(n1451), .B(n45185), .Z(n45184) );
  XOR U44918 ( .A(n45170), .B(n45186), .Z(n45176) );
  AND U44919 ( .A(n45187), .B(n45173), .Z(n45186) );
  XNOR U44920 ( .A(n45004), .B(n45170), .Z(n45173) );
  XOR U44921 ( .A(n45054), .B(n45188), .Z(n45004) );
  AND U44922 ( .A(n1435), .B(n45189), .Z(n45188) );
  XOR U44923 ( .A(n45050), .B(n45054), .Z(n45189) );
  XNOR U44924 ( .A(n45190), .B(n45170), .Z(n45187) );
  IV U44925 ( .A(n44962), .Z(n45190) );
  XOR U44926 ( .A(n45191), .B(n45192), .Z(n44962) );
  AND U44927 ( .A(n1451), .B(n45193), .Z(n45192) );
  XOR U44928 ( .A(n45194), .B(n45195), .Z(n45170) );
  AND U44929 ( .A(n45196), .B(n45197), .Z(n45195) );
  XNOR U44930 ( .A(n45014), .B(n45194), .Z(n45197) );
  XOR U44931 ( .A(n45082), .B(n45198), .Z(n45014) );
  AND U44932 ( .A(n1435), .B(n45199), .Z(n45198) );
  XOR U44933 ( .A(n45078), .B(n45082), .Z(n45199) );
  XOR U44934 ( .A(n45194), .B(n44971), .Z(n45196) );
  XOR U44935 ( .A(n45200), .B(n45201), .Z(n44971) );
  AND U44936 ( .A(n1451), .B(n45202), .Z(n45201) );
  XOR U44937 ( .A(n45203), .B(n45204), .Z(n45194) );
  AND U44938 ( .A(n45205), .B(n45206), .Z(n45204) );
  XNOR U44939 ( .A(n45203), .B(n45022), .Z(n45206) );
  XOR U44940 ( .A(n45133), .B(n45207), .Z(n45022) );
  AND U44941 ( .A(n1435), .B(n45208), .Z(n45207) );
  XOR U44942 ( .A(n45129), .B(n45133), .Z(n45208) );
  XNOR U44943 ( .A(n45209), .B(n45203), .Z(n45205) );
  IV U44944 ( .A(n44981), .Z(n45209) );
  XOR U44945 ( .A(n45210), .B(n45211), .Z(n44981) );
  AND U44946 ( .A(n1451), .B(n45212), .Z(n45211) );
  AND U44947 ( .A(n45174), .B(n45163), .Z(n45203) );
  XNOR U44948 ( .A(n45213), .B(n45214), .Z(n45163) );
  AND U44949 ( .A(n1435), .B(n45145), .Z(n45214) );
  XNOR U44950 ( .A(n45143), .B(n45213), .Z(n45145) );
  XNOR U44951 ( .A(n45215), .B(n45216), .Z(n1435) );
  AND U44952 ( .A(n45217), .B(n45218), .Z(n45216) );
  XNOR U44953 ( .A(n45215), .B(n45034), .Z(n45218) );
  IV U44954 ( .A(n45038), .Z(n45034) );
  XOR U44955 ( .A(n45219), .B(n45220), .Z(n45038) );
  AND U44956 ( .A(n1439), .B(n45221), .Z(n45220) );
  XOR U44957 ( .A(n45222), .B(n45219), .Z(n45221) );
  XNOR U44958 ( .A(n45215), .B(n45150), .Z(n45217) );
  XOR U44959 ( .A(n45223), .B(n45224), .Z(n45150) );
  AND U44960 ( .A(n1447), .B(n45185), .Z(n45224) );
  XOR U44961 ( .A(n45183), .B(n45223), .Z(n45185) );
  XOR U44962 ( .A(n45225), .B(n45226), .Z(n45215) );
  AND U44963 ( .A(n45227), .B(n45228), .Z(n45226) );
  XNOR U44964 ( .A(n45225), .B(n45050), .Z(n45228) );
  IV U44965 ( .A(n45053), .Z(n45050) );
  XOR U44966 ( .A(n45229), .B(n45230), .Z(n45053) );
  AND U44967 ( .A(n1439), .B(n45231), .Z(n45230) );
  XOR U44968 ( .A(n45232), .B(n45229), .Z(n45231) );
  XOR U44969 ( .A(n45054), .B(n45225), .Z(n45227) );
  XOR U44970 ( .A(n45233), .B(n45234), .Z(n45054) );
  AND U44971 ( .A(n1447), .B(n45193), .Z(n45234) );
  XOR U44972 ( .A(n45233), .B(n45191), .Z(n45193) );
  XOR U44973 ( .A(n45235), .B(n45236), .Z(n45225) );
  AND U44974 ( .A(n45237), .B(n45238), .Z(n45236) );
  XNOR U44975 ( .A(n45235), .B(n45078), .Z(n45238) );
  IV U44976 ( .A(n45081), .Z(n45078) );
  XOR U44977 ( .A(n45239), .B(n45240), .Z(n45081) );
  AND U44978 ( .A(n1439), .B(n45241), .Z(n45240) );
  XNOR U44979 ( .A(n45242), .B(n45239), .Z(n45241) );
  XOR U44980 ( .A(n45082), .B(n45235), .Z(n45237) );
  XOR U44981 ( .A(n45243), .B(n45244), .Z(n45082) );
  AND U44982 ( .A(n1447), .B(n45202), .Z(n45244) );
  XOR U44983 ( .A(n45243), .B(n45200), .Z(n45202) );
  XOR U44984 ( .A(n45159), .B(n45245), .Z(n45235) );
  AND U44985 ( .A(n45161), .B(n45246), .Z(n45245) );
  XNOR U44986 ( .A(n45159), .B(n45129), .Z(n45246) );
  IV U44987 ( .A(n45132), .Z(n45129) );
  XOR U44988 ( .A(n45247), .B(n45248), .Z(n45132) );
  AND U44989 ( .A(n1439), .B(n45249), .Z(n45248) );
  XOR U44990 ( .A(n45250), .B(n45247), .Z(n45249) );
  XOR U44991 ( .A(n45133), .B(n45159), .Z(n45161) );
  XOR U44992 ( .A(n45251), .B(n45252), .Z(n45133) );
  AND U44993 ( .A(n1447), .B(n45212), .Z(n45252) );
  XOR U44994 ( .A(n45251), .B(n45210), .Z(n45212) );
  AND U44995 ( .A(n45213), .B(n45143), .Z(n45159) );
  XNOR U44996 ( .A(n45253), .B(n45254), .Z(n45143) );
  AND U44997 ( .A(n1439), .B(n45255), .Z(n45254) );
  XNOR U44998 ( .A(n45256), .B(n45253), .Z(n45255) );
  XNOR U44999 ( .A(n45257), .B(n45258), .Z(n1439) );
  AND U45000 ( .A(n45259), .B(n45260), .Z(n45258) );
  XOR U45001 ( .A(n45222), .B(n45257), .Z(n45260) );
  AND U45002 ( .A(n45261), .B(n45262), .Z(n45222) );
  XNOR U45003 ( .A(n45219), .B(n45257), .Z(n45259) );
  XNOR U45004 ( .A(n45263), .B(n45264), .Z(n45219) );
  AND U45005 ( .A(n1443), .B(n45265), .Z(n45264) );
  XNOR U45006 ( .A(n45266), .B(n45267), .Z(n45265) );
  XOR U45007 ( .A(n45268), .B(n45269), .Z(n45257) );
  AND U45008 ( .A(n45270), .B(n45271), .Z(n45269) );
  XNOR U45009 ( .A(n45268), .B(n45261), .Z(n45271) );
  IV U45010 ( .A(n45232), .Z(n45261) );
  XOR U45011 ( .A(n45272), .B(n45273), .Z(n45232) );
  XOR U45012 ( .A(n45274), .B(n45262), .Z(n45273) );
  AND U45013 ( .A(n45242), .B(n45275), .Z(n45262) );
  AND U45014 ( .A(n45276), .B(n45277), .Z(n45274) );
  XOR U45015 ( .A(n45278), .B(n45272), .Z(n45276) );
  XNOR U45016 ( .A(n45229), .B(n45268), .Z(n45270) );
  XNOR U45017 ( .A(n45279), .B(n45280), .Z(n45229) );
  AND U45018 ( .A(n1443), .B(n45281), .Z(n45280) );
  XNOR U45019 ( .A(n45282), .B(n45283), .Z(n45281) );
  XOR U45020 ( .A(n45284), .B(n45285), .Z(n45268) );
  AND U45021 ( .A(n45286), .B(n45287), .Z(n45285) );
  XNOR U45022 ( .A(n45284), .B(n45242), .Z(n45287) );
  XOR U45023 ( .A(n45288), .B(n45277), .Z(n45242) );
  XNOR U45024 ( .A(n45289), .B(n45272), .Z(n45277) );
  XOR U45025 ( .A(n45290), .B(n45291), .Z(n45272) );
  AND U45026 ( .A(n45292), .B(n45293), .Z(n45291) );
  XOR U45027 ( .A(n45294), .B(n45290), .Z(n45292) );
  XNOR U45028 ( .A(n45295), .B(n45296), .Z(n45289) );
  AND U45029 ( .A(n45297), .B(n45298), .Z(n45296) );
  XOR U45030 ( .A(n45295), .B(n45299), .Z(n45297) );
  XNOR U45031 ( .A(n45278), .B(n45275), .Z(n45288) );
  AND U45032 ( .A(n45300), .B(n45301), .Z(n45275) );
  XOR U45033 ( .A(n45302), .B(n45303), .Z(n45278) );
  AND U45034 ( .A(n45304), .B(n45305), .Z(n45303) );
  XOR U45035 ( .A(n45302), .B(n45306), .Z(n45304) );
  XNOR U45036 ( .A(n45239), .B(n45284), .Z(n45286) );
  XNOR U45037 ( .A(n45307), .B(n45308), .Z(n45239) );
  AND U45038 ( .A(n1443), .B(n45309), .Z(n45308) );
  XNOR U45039 ( .A(n45310), .B(n45311), .Z(n45309) );
  XOR U45040 ( .A(n45312), .B(n45313), .Z(n45284) );
  AND U45041 ( .A(n45314), .B(n45315), .Z(n45313) );
  XNOR U45042 ( .A(n45312), .B(n45300), .Z(n45315) );
  IV U45043 ( .A(n45250), .Z(n45300) );
  XNOR U45044 ( .A(n45316), .B(n45293), .Z(n45250) );
  XNOR U45045 ( .A(n45317), .B(n45299), .Z(n45293) );
  XNOR U45046 ( .A(n45318), .B(n45319), .Z(n45299) );
  NOR U45047 ( .A(n45320), .B(n45321), .Z(n45319) );
  XOR U45048 ( .A(n45318), .B(n45322), .Z(n45320) );
  XNOR U45049 ( .A(n45298), .B(n45290), .Z(n45317) );
  XOR U45050 ( .A(n45323), .B(n45324), .Z(n45290) );
  AND U45051 ( .A(n45325), .B(n45326), .Z(n45324) );
  XOR U45052 ( .A(n45323), .B(n45327), .Z(n45325) );
  XNOR U45053 ( .A(n45328), .B(n45295), .Z(n45298) );
  XOR U45054 ( .A(n45329), .B(n45330), .Z(n45295) );
  AND U45055 ( .A(n45331), .B(n45332), .Z(n45330) );
  XNOR U45056 ( .A(n45333), .B(n45334), .Z(n45331) );
  IV U45057 ( .A(n45329), .Z(n45333) );
  XNOR U45058 ( .A(n45335), .B(n45336), .Z(n45328) );
  NOR U45059 ( .A(n45337), .B(n45338), .Z(n45336) );
  XNOR U45060 ( .A(n45335), .B(n45339), .Z(n45337) );
  XNOR U45061 ( .A(n45294), .B(n45301), .Z(n45316) );
  NOR U45062 ( .A(n45256), .B(n45340), .Z(n45301) );
  XOR U45063 ( .A(n45306), .B(n45305), .Z(n45294) );
  XNOR U45064 ( .A(n45341), .B(n45302), .Z(n45305) );
  XOR U45065 ( .A(n45342), .B(n45343), .Z(n45302) );
  AND U45066 ( .A(n45344), .B(n45345), .Z(n45343) );
  XNOR U45067 ( .A(n45346), .B(n45347), .Z(n45344) );
  IV U45068 ( .A(n45342), .Z(n45346) );
  XNOR U45069 ( .A(n45348), .B(n45349), .Z(n45341) );
  NOR U45070 ( .A(n45350), .B(n45351), .Z(n45349) );
  XNOR U45071 ( .A(n45348), .B(n45352), .Z(n45350) );
  XOR U45072 ( .A(n45353), .B(n45354), .Z(n45306) );
  NOR U45073 ( .A(n45355), .B(n45356), .Z(n45354) );
  XNOR U45074 ( .A(n45353), .B(n45357), .Z(n45355) );
  XNOR U45075 ( .A(n45247), .B(n45312), .Z(n45314) );
  XNOR U45076 ( .A(n45358), .B(n45359), .Z(n45247) );
  AND U45077 ( .A(n1443), .B(n45360), .Z(n45359) );
  XNOR U45078 ( .A(n45361), .B(n45362), .Z(n45360) );
  AND U45079 ( .A(n45253), .B(n45256), .Z(n45312) );
  XOR U45080 ( .A(n45363), .B(n45340), .Z(n45256) );
  XNOR U45081 ( .A(p_input[1152]), .B(p_input[2048]), .Z(n45340) );
  XNOR U45082 ( .A(n45327), .B(n45326), .Z(n45363) );
  XNOR U45083 ( .A(n45364), .B(n45334), .Z(n45326) );
  XNOR U45084 ( .A(n45322), .B(n45321), .Z(n45334) );
  XNOR U45085 ( .A(n45365), .B(n45318), .Z(n45321) );
  XNOR U45086 ( .A(p_input[1162]), .B(p_input[2058]), .Z(n45318) );
  XOR U45087 ( .A(p_input[1163]), .B(n29030), .Z(n45365) );
  XOR U45088 ( .A(p_input[1164]), .B(p_input[2060]), .Z(n45322) );
  XOR U45089 ( .A(n45332), .B(n45366), .Z(n45364) );
  IV U45090 ( .A(n45323), .Z(n45366) );
  XOR U45091 ( .A(p_input[1153]), .B(p_input[2049]), .Z(n45323) );
  XNOR U45092 ( .A(n45367), .B(n45339), .Z(n45332) );
  XNOR U45093 ( .A(p_input[1167]), .B(n29033), .Z(n45339) );
  XOR U45094 ( .A(n45329), .B(n45338), .Z(n45367) );
  XOR U45095 ( .A(n45368), .B(n45335), .Z(n45338) );
  XOR U45096 ( .A(p_input[1165]), .B(p_input[2061]), .Z(n45335) );
  XOR U45097 ( .A(p_input[1166]), .B(n29035), .Z(n45368) );
  XOR U45098 ( .A(p_input[1161]), .B(p_input[2057]), .Z(n45329) );
  XOR U45099 ( .A(n45347), .B(n45345), .Z(n45327) );
  XNOR U45100 ( .A(n45369), .B(n45352), .Z(n45345) );
  XOR U45101 ( .A(p_input[1160]), .B(p_input[2056]), .Z(n45352) );
  XOR U45102 ( .A(n45342), .B(n45351), .Z(n45369) );
  XOR U45103 ( .A(n45370), .B(n45348), .Z(n45351) );
  XOR U45104 ( .A(p_input[1158]), .B(p_input[2054]), .Z(n45348) );
  XOR U45105 ( .A(p_input[1159]), .B(n30404), .Z(n45370) );
  XOR U45106 ( .A(p_input[1154]), .B(p_input[2050]), .Z(n45342) );
  XNOR U45107 ( .A(n45357), .B(n45356), .Z(n45347) );
  XOR U45108 ( .A(n45371), .B(n45353), .Z(n45356) );
  XOR U45109 ( .A(p_input[1155]), .B(p_input[2051]), .Z(n45353) );
  XOR U45110 ( .A(p_input[1156]), .B(n30406), .Z(n45371) );
  XOR U45111 ( .A(p_input[1157]), .B(p_input[2053]), .Z(n45357) );
  XNOR U45112 ( .A(n45372), .B(n45373), .Z(n45253) );
  AND U45113 ( .A(n1443), .B(n45374), .Z(n45373) );
  XNOR U45114 ( .A(n45375), .B(n45376), .Z(n1443) );
  AND U45115 ( .A(n45377), .B(n45378), .Z(n45376) );
  XOR U45116 ( .A(n45267), .B(n45375), .Z(n45378) );
  XNOR U45117 ( .A(n45379), .B(n45375), .Z(n45377) );
  XOR U45118 ( .A(n45380), .B(n45381), .Z(n45375) );
  AND U45119 ( .A(n45382), .B(n45383), .Z(n45381) );
  XOR U45120 ( .A(n45282), .B(n45380), .Z(n45383) );
  XOR U45121 ( .A(n45380), .B(n45283), .Z(n45382) );
  XOR U45122 ( .A(n45384), .B(n45385), .Z(n45380) );
  AND U45123 ( .A(n45386), .B(n45387), .Z(n45385) );
  XOR U45124 ( .A(n45310), .B(n45384), .Z(n45387) );
  XOR U45125 ( .A(n45384), .B(n45311), .Z(n45386) );
  XOR U45126 ( .A(n45388), .B(n45389), .Z(n45384) );
  AND U45127 ( .A(n45390), .B(n45391), .Z(n45389) );
  XOR U45128 ( .A(n45388), .B(n45361), .Z(n45391) );
  XNOR U45129 ( .A(n45392), .B(n45393), .Z(n45213) );
  AND U45130 ( .A(n1447), .B(n45394), .Z(n45393) );
  XNOR U45131 ( .A(n45395), .B(n45396), .Z(n1447) );
  AND U45132 ( .A(n45397), .B(n45398), .Z(n45396) );
  XOR U45133 ( .A(n45395), .B(n45223), .Z(n45398) );
  XNOR U45134 ( .A(n45395), .B(n45183), .Z(n45397) );
  XOR U45135 ( .A(n45399), .B(n45400), .Z(n45395) );
  AND U45136 ( .A(n45401), .B(n45402), .Z(n45400) );
  XOR U45137 ( .A(n45399), .B(n45191), .Z(n45401) );
  XOR U45138 ( .A(n45403), .B(n45404), .Z(n45174) );
  AND U45139 ( .A(n1451), .B(n45394), .Z(n45404) );
  XNOR U45140 ( .A(n45392), .B(n45403), .Z(n45394) );
  XNOR U45141 ( .A(n45405), .B(n45406), .Z(n1451) );
  AND U45142 ( .A(n45407), .B(n45408), .Z(n45406) );
  XNOR U45143 ( .A(n45409), .B(n45405), .Z(n45408) );
  IV U45144 ( .A(n45223), .Z(n45409) );
  XOR U45145 ( .A(n45379), .B(n45410), .Z(n45223) );
  AND U45146 ( .A(n1454), .B(n45411), .Z(n45410) );
  XOR U45147 ( .A(n45266), .B(n45263), .Z(n45411) );
  IV U45148 ( .A(n45379), .Z(n45266) );
  XNOR U45149 ( .A(n45183), .B(n45405), .Z(n45407) );
  XOR U45150 ( .A(n45412), .B(n45413), .Z(n45183) );
  AND U45151 ( .A(n1470), .B(n45414), .Z(n45413) );
  XOR U45152 ( .A(n45399), .B(n45415), .Z(n45405) );
  AND U45153 ( .A(n45416), .B(n45402), .Z(n45415) );
  XNOR U45154 ( .A(n45233), .B(n45399), .Z(n45402) );
  XOR U45155 ( .A(n45283), .B(n45417), .Z(n45233) );
  AND U45156 ( .A(n1454), .B(n45418), .Z(n45417) );
  XOR U45157 ( .A(n45279), .B(n45283), .Z(n45418) );
  XNOR U45158 ( .A(n45419), .B(n45399), .Z(n45416) );
  IV U45159 ( .A(n45191), .Z(n45419) );
  XOR U45160 ( .A(n45420), .B(n45421), .Z(n45191) );
  AND U45161 ( .A(n1470), .B(n45422), .Z(n45421) );
  XOR U45162 ( .A(n45423), .B(n45424), .Z(n45399) );
  AND U45163 ( .A(n45425), .B(n45426), .Z(n45424) );
  XNOR U45164 ( .A(n45243), .B(n45423), .Z(n45426) );
  XOR U45165 ( .A(n45311), .B(n45427), .Z(n45243) );
  AND U45166 ( .A(n1454), .B(n45428), .Z(n45427) );
  XOR U45167 ( .A(n45307), .B(n45311), .Z(n45428) );
  XOR U45168 ( .A(n45423), .B(n45200), .Z(n45425) );
  XOR U45169 ( .A(n45429), .B(n45430), .Z(n45200) );
  AND U45170 ( .A(n1470), .B(n45431), .Z(n45430) );
  XOR U45171 ( .A(n45432), .B(n45433), .Z(n45423) );
  AND U45172 ( .A(n45434), .B(n45435), .Z(n45433) );
  XNOR U45173 ( .A(n45432), .B(n45251), .Z(n45435) );
  XOR U45174 ( .A(n45362), .B(n45436), .Z(n45251) );
  AND U45175 ( .A(n1454), .B(n45437), .Z(n45436) );
  XOR U45176 ( .A(n45358), .B(n45362), .Z(n45437) );
  XNOR U45177 ( .A(n45438), .B(n45432), .Z(n45434) );
  IV U45178 ( .A(n45210), .Z(n45438) );
  XOR U45179 ( .A(n45439), .B(n45440), .Z(n45210) );
  AND U45180 ( .A(n1470), .B(n45441), .Z(n45440) );
  AND U45181 ( .A(n45403), .B(n45392), .Z(n45432) );
  XNOR U45182 ( .A(n45442), .B(n45443), .Z(n45392) );
  AND U45183 ( .A(n1454), .B(n45374), .Z(n45443) );
  XNOR U45184 ( .A(n45372), .B(n45442), .Z(n45374) );
  XNOR U45185 ( .A(n45444), .B(n45445), .Z(n1454) );
  AND U45186 ( .A(n45446), .B(n45447), .Z(n45445) );
  XNOR U45187 ( .A(n45444), .B(n45263), .Z(n45447) );
  IV U45188 ( .A(n45267), .Z(n45263) );
  XOR U45189 ( .A(n45448), .B(n45449), .Z(n45267) );
  AND U45190 ( .A(n1458), .B(n45450), .Z(n45449) );
  XOR U45191 ( .A(n45451), .B(n45448), .Z(n45450) );
  XNOR U45192 ( .A(n45444), .B(n45379), .Z(n45446) );
  XOR U45193 ( .A(n45452), .B(n45453), .Z(n45379) );
  AND U45194 ( .A(n1466), .B(n45414), .Z(n45453) );
  XOR U45195 ( .A(n45412), .B(n45452), .Z(n45414) );
  XOR U45196 ( .A(n45454), .B(n45455), .Z(n45444) );
  AND U45197 ( .A(n45456), .B(n45457), .Z(n45455) );
  XNOR U45198 ( .A(n45454), .B(n45279), .Z(n45457) );
  IV U45199 ( .A(n45282), .Z(n45279) );
  XOR U45200 ( .A(n45458), .B(n45459), .Z(n45282) );
  AND U45201 ( .A(n1458), .B(n45460), .Z(n45459) );
  XOR U45202 ( .A(n45461), .B(n45458), .Z(n45460) );
  XOR U45203 ( .A(n45283), .B(n45454), .Z(n45456) );
  XOR U45204 ( .A(n45462), .B(n45463), .Z(n45283) );
  AND U45205 ( .A(n1466), .B(n45422), .Z(n45463) );
  XOR U45206 ( .A(n45462), .B(n45420), .Z(n45422) );
  XOR U45207 ( .A(n45464), .B(n45465), .Z(n45454) );
  AND U45208 ( .A(n45466), .B(n45467), .Z(n45465) );
  XNOR U45209 ( .A(n45464), .B(n45307), .Z(n45467) );
  IV U45210 ( .A(n45310), .Z(n45307) );
  XOR U45211 ( .A(n45468), .B(n45469), .Z(n45310) );
  AND U45212 ( .A(n1458), .B(n45470), .Z(n45469) );
  XNOR U45213 ( .A(n45471), .B(n45468), .Z(n45470) );
  XOR U45214 ( .A(n45311), .B(n45464), .Z(n45466) );
  XOR U45215 ( .A(n45472), .B(n45473), .Z(n45311) );
  AND U45216 ( .A(n1466), .B(n45431), .Z(n45473) );
  XOR U45217 ( .A(n45472), .B(n45429), .Z(n45431) );
  XOR U45218 ( .A(n45388), .B(n45474), .Z(n45464) );
  AND U45219 ( .A(n45390), .B(n45475), .Z(n45474) );
  XNOR U45220 ( .A(n45388), .B(n45358), .Z(n45475) );
  IV U45221 ( .A(n45361), .Z(n45358) );
  XOR U45222 ( .A(n45476), .B(n45477), .Z(n45361) );
  AND U45223 ( .A(n1458), .B(n45478), .Z(n45477) );
  XOR U45224 ( .A(n45479), .B(n45476), .Z(n45478) );
  XOR U45225 ( .A(n45362), .B(n45388), .Z(n45390) );
  XOR U45226 ( .A(n45480), .B(n45481), .Z(n45362) );
  AND U45227 ( .A(n1466), .B(n45441), .Z(n45481) );
  XOR U45228 ( .A(n45480), .B(n45439), .Z(n45441) );
  AND U45229 ( .A(n45442), .B(n45372), .Z(n45388) );
  XNOR U45230 ( .A(n45482), .B(n45483), .Z(n45372) );
  AND U45231 ( .A(n1458), .B(n45484), .Z(n45483) );
  XNOR U45232 ( .A(n45485), .B(n45482), .Z(n45484) );
  XNOR U45233 ( .A(n45486), .B(n45487), .Z(n1458) );
  AND U45234 ( .A(n45488), .B(n45489), .Z(n45487) );
  XOR U45235 ( .A(n45451), .B(n45486), .Z(n45489) );
  AND U45236 ( .A(n45490), .B(n45491), .Z(n45451) );
  XNOR U45237 ( .A(n45448), .B(n45486), .Z(n45488) );
  XNOR U45238 ( .A(n45492), .B(n45493), .Z(n45448) );
  AND U45239 ( .A(n1462), .B(n45494), .Z(n45493) );
  XNOR U45240 ( .A(n45495), .B(n45496), .Z(n45494) );
  XOR U45241 ( .A(n45497), .B(n45498), .Z(n45486) );
  AND U45242 ( .A(n45499), .B(n45500), .Z(n45498) );
  XNOR U45243 ( .A(n45497), .B(n45490), .Z(n45500) );
  IV U45244 ( .A(n45461), .Z(n45490) );
  XOR U45245 ( .A(n45501), .B(n45502), .Z(n45461) );
  XOR U45246 ( .A(n45503), .B(n45491), .Z(n45502) );
  AND U45247 ( .A(n45471), .B(n45504), .Z(n45491) );
  AND U45248 ( .A(n45505), .B(n45506), .Z(n45503) );
  XOR U45249 ( .A(n45507), .B(n45501), .Z(n45505) );
  XNOR U45250 ( .A(n45458), .B(n45497), .Z(n45499) );
  XNOR U45251 ( .A(n45508), .B(n45509), .Z(n45458) );
  AND U45252 ( .A(n1462), .B(n45510), .Z(n45509) );
  XNOR U45253 ( .A(n45511), .B(n45512), .Z(n45510) );
  XOR U45254 ( .A(n45513), .B(n45514), .Z(n45497) );
  AND U45255 ( .A(n45515), .B(n45516), .Z(n45514) );
  XNOR U45256 ( .A(n45513), .B(n45471), .Z(n45516) );
  XOR U45257 ( .A(n45517), .B(n45506), .Z(n45471) );
  XNOR U45258 ( .A(n45518), .B(n45501), .Z(n45506) );
  XOR U45259 ( .A(n45519), .B(n45520), .Z(n45501) );
  AND U45260 ( .A(n45521), .B(n45522), .Z(n45520) );
  XOR U45261 ( .A(n45523), .B(n45519), .Z(n45521) );
  XNOR U45262 ( .A(n45524), .B(n45525), .Z(n45518) );
  AND U45263 ( .A(n45526), .B(n45527), .Z(n45525) );
  XOR U45264 ( .A(n45524), .B(n45528), .Z(n45526) );
  XNOR U45265 ( .A(n45507), .B(n45504), .Z(n45517) );
  AND U45266 ( .A(n45529), .B(n45530), .Z(n45504) );
  XOR U45267 ( .A(n45531), .B(n45532), .Z(n45507) );
  AND U45268 ( .A(n45533), .B(n45534), .Z(n45532) );
  XOR U45269 ( .A(n45531), .B(n45535), .Z(n45533) );
  XNOR U45270 ( .A(n45468), .B(n45513), .Z(n45515) );
  XNOR U45271 ( .A(n45536), .B(n45537), .Z(n45468) );
  AND U45272 ( .A(n1462), .B(n45538), .Z(n45537) );
  XNOR U45273 ( .A(n45539), .B(n45540), .Z(n45538) );
  XOR U45274 ( .A(n45541), .B(n45542), .Z(n45513) );
  AND U45275 ( .A(n45543), .B(n45544), .Z(n45542) );
  XNOR U45276 ( .A(n45541), .B(n45529), .Z(n45544) );
  IV U45277 ( .A(n45479), .Z(n45529) );
  XNOR U45278 ( .A(n45545), .B(n45522), .Z(n45479) );
  XNOR U45279 ( .A(n45546), .B(n45528), .Z(n45522) );
  XNOR U45280 ( .A(n45547), .B(n45548), .Z(n45528) );
  NOR U45281 ( .A(n45549), .B(n45550), .Z(n45548) );
  XOR U45282 ( .A(n45547), .B(n45551), .Z(n45549) );
  XNOR U45283 ( .A(n45527), .B(n45519), .Z(n45546) );
  XOR U45284 ( .A(n45552), .B(n45553), .Z(n45519) );
  AND U45285 ( .A(n45554), .B(n45555), .Z(n45553) );
  XOR U45286 ( .A(n45552), .B(n45556), .Z(n45554) );
  XNOR U45287 ( .A(n45557), .B(n45524), .Z(n45527) );
  XOR U45288 ( .A(n45558), .B(n45559), .Z(n45524) );
  AND U45289 ( .A(n45560), .B(n45561), .Z(n45559) );
  XNOR U45290 ( .A(n45562), .B(n45563), .Z(n45560) );
  IV U45291 ( .A(n45558), .Z(n45562) );
  XNOR U45292 ( .A(n45564), .B(n45565), .Z(n45557) );
  NOR U45293 ( .A(n45566), .B(n45567), .Z(n45565) );
  XNOR U45294 ( .A(n45564), .B(n45568), .Z(n45566) );
  XNOR U45295 ( .A(n45523), .B(n45530), .Z(n45545) );
  NOR U45296 ( .A(n45485), .B(n45569), .Z(n45530) );
  XOR U45297 ( .A(n45535), .B(n45534), .Z(n45523) );
  XNOR U45298 ( .A(n45570), .B(n45531), .Z(n45534) );
  XOR U45299 ( .A(n45571), .B(n45572), .Z(n45531) );
  AND U45300 ( .A(n45573), .B(n45574), .Z(n45572) );
  XNOR U45301 ( .A(n45575), .B(n45576), .Z(n45573) );
  IV U45302 ( .A(n45571), .Z(n45575) );
  XNOR U45303 ( .A(n45577), .B(n45578), .Z(n45570) );
  NOR U45304 ( .A(n45579), .B(n45580), .Z(n45578) );
  XNOR U45305 ( .A(n45577), .B(n45581), .Z(n45579) );
  XOR U45306 ( .A(n45582), .B(n45583), .Z(n45535) );
  NOR U45307 ( .A(n45584), .B(n45585), .Z(n45583) );
  XNOR U45308 ( .A(n45582), .B(n45586), .Z(n45584) );
  XNOR U45309 ( .A(n45476), .B(n45541), .Z(n45543) );
  XNOR U45310 ( .A(n45587), .B(n45588), .Z(n45476) );
  AND U45311 ( .A(n1462), .B(n45589), .Z(n45588) );
  XNOR U45312 ( .A(n45590), .B(n45591), .Z(n45589) );
  AND U45313 ( .A(n45482), .B(n45485), .Z(n45541) );
  XOR U45314 ( .A(n45592), .B(n45569), .Z(n45485) );
  XNOR U45315 ( .A(p_input[1168]), .B(p_input[2048]), .Z(n45569) );
  XNOR U45316 ( .A(n45556), .B(n45555), .Z(n45592) );
  XNOR U45317 ( .A(n45593), .B(n45563), .Z(n45555) );
  XNOR U45318 ( .A(n45551), .B(n45550), .Z(n45563) );
  XNOR U45319 ( .A(n45594), .B(n45547), .Z(n45550) );
  XNOR U45320 ( .A(p_input[1178]), .B(p_input[2058]), .Z(n45547) );
  XOR U45321 ( .A(p_input[1179]), .B(n29030), .Z(n45594) );
  XOR U45322 ( .A(p_input[1180]), .B(p_input[2060]), .Z(n45551) );
  XOR U45323 ( .A(n45561), .B(n45595), .Z(n45593) );
  IV U45324 ( .A(n45552), .Z(n45595) );
  XOR U45325 ( .A(p_input[1169]), .B(p_input[2049]), .Z(n45552) );
  XNOR U45326 ( .A(n45596), .B(n45568), .Z(n45561) );
  XNOR U45327 ( .A(p_input[1183]), .B(n29033), .Z(n45568) );
  XOR U45328 ( .A(n45558), .B(n45567), .Z(n45596) );
  XOR U45329 ( .A(n45597), .B(n45564), .Z(n45567) );
  XOR U45330 ( .A(p_input[1181]), .B(p_input[2061]), .Z(n45564) );
  XOR U45331 ( .A(p_input[1182]), .B(n29035), .Z(n45597) );
  XOR U45332 ( .A(p_input[1177]), .B(p_input[2057]), .Z(n45558) );
  XOR U45333 ( .A(n45576), .B(n45574), .Z(n45556) );
  XNOR U45334 ( .A(n45598), .B(n45581), .Z(n45574) );
  XOR U45335 ( .A(p_input[1176]), .B(p_input[2056]), .Z(n45581) );
  XOR U45336 ( .A(n45571), .B(n45580), .Z(n45598) );
  XOR U45337 ( .A(n45599), .B(n45577), .Z(n45580) );
  XOR U45338 ( .A(p_input[1174]), .B(p_input[2054]), .Z(n45577) );
  XOR U45339 ( .A(p_input[1175]), .B(n30404), .Z(n45599) );
  XOR U45340 ( .A(p_input[1170]), .B(p_input[2050]), .Z(n45571) );
  XNOR U45341 ( .A(n45586), .B(n45585), .Z(n45576) );
  XOR U45342 ( .A(n45600), .B(n45582), .Z(n45585) );
  XOR U45343 ( .A(p_input[1171]), .B(p_input[2051]), .Z(n45582) );
  XOR U45344 ( .A(p_input[1172]), .B(n30406), .Z(n45600) );
  XOR U45345 ( .A(p_input[1173]), .B(p_input[2053]), .Z(n45586) );
  XNOR U45346 ( .A(n45601), .B(n45602), .Z(n45482) );
  AND U45347 ( .A(n1462), .B(n45603), .Z(n45602) );
  XNOR U45348 ( .A(n45604), .B(n45605), .Z(n1462) );
  AND U45349 ( .A(n45606), .B(n45607), .Z(n45605) );
  XOR U45350 ( .A(n45496), .B(n45604), .Z(n45607) );
  XNOR U45351 ( .A(n45608), .B(n45604), .Z(n45606) );
  XOR U45352 ( .A(n45609), .B(n45610), .Z(n45604) );
  AND U45353 ( .A(n45611), .B(n45612), .Z(n45610) );
  XOR U45354 ( .A(n45511), .B(n45609), .Z(n45612) );
  XOR U45355 ( .A(n45609), .B(n45512), .Z(n45611) );
  XOR U45356 ( .A(n45613), .B(n45614), .Z(n45609) );
  AND U45357 ( .A(n45615), .B(n45616), .Z(n45614) );
  XOR U45358 ( .A(n45539), .B(n45613), .Z(n45616) );
  XOR U45359 ( .A(n45613), .B(n45540), .Z(n45615) );
  XOR U45360 ( .A(n45617), .B(n45618), .Z(n45613) );
  AND U45361 ( .A(n45619), .B(n45620), .Z(n45618) );
  XOR U45362 ( .A(n45617), .B(n45590), .Z(n45620) );
  XNOR U45363 ( .A(n45621), .B(n45622), .Z(n45442) );
  AND U45364 ( .A(n1466), .B(n45623), .Z(n45622) );
  XNOR U45365 ( .A(n45624), .B(n45625), .Z(n1466) );
  AND U45366 ( .A(n45626), .B(n45627), .Z(n45625) );
  XOR U45367 ( .A(n45624), .B(n45452), .Z(n45627) );
  XNOR U45368 ( .A(n45624), .B(n45412), .Z(n45626) );
  XOR U45369 ( .A(n45628), .B(n45629), .Z(n45624) );
  AND U45370 ( .A(n45630), .B(n45631), .Z(n45629) );
  XOR U45371 ( .A(n45628), .B(n45420), .Z(n45630) );
  XOR U45372 ( .A(n45632), .B(n45633), .Z(n45403) );
  AND U45373 ( .A(n1470), .B(n45623), .Z(n45633) );
  XNOR U45374 ( .A(n45621), .B(n45632), .Z(n45623) );
  XNOR U45375 ( .A(n45634), .B(n45635), .Z(n1470) );
  AND U45376 ( .A(n45636), .B(n45637), .Z(n45635) );
  XNOR U45377 ( .A(n45638), .B(n45634), .Z(n45637) );
  IV U45378 ( .A(n45452), .Z(n45638) );
  XOR U45379 ( .A(n45608), .B(n45639), .Z(n45452) );
  AND U45380 ( .A(n1473), .B(n45640), .Z(n45639) );
  XOR U45381 ( .A(n45495), .B(n45492), .Z(n45640) );
  IV U45382 ( .A(n45608), .Z(n45495) );
  XNOR U45383 ( .A(n45412), .B(n45634), .Z(n45636) );
  XOR U45384 ( .A(n45641), .B(n45642), .Z(n45412) );
  AND U45385 ( .A(n1489), .B(n45643), .Z(n45642) );
  XOR U45386 ( .A(n45628), .B(n45644), .Z(n45634) );
  AND U45387 ( .A(n45645), .B(n45631), .Z(n45644) );
  XNOR U45388 ( .A(n45462), .B(n45628), .Z(n45631) );
  XOR U45389 ( .A(n45512), .B(n45646), .Z(n45462) );
  AND U45390 ( .A(n1473), .B(n45647), .Z(n45646) );
  XOR U45391 ( .A(n45508), .B(n45512), .Z(n45647) );
  XNOR U45392 ( .A(n45648), .B(n45628), .Z(n45645) );
  IV U45393 ( .A(n45420), .Z(n45648) );
  XOR U45394 ( .A(n45649), .B(n45650), .Z(n45420) );
  AND U45395 ( .A(n1489), .B(n45651), .Z(n45650) );
  XOR U45396 ( .A(n45652), .B(n45653), .Z(n45628) );
  AND U45397 ( .A(n45654), .B(n45655), .Z(n45653) );
  XNOR U45398 ( .A(n45472), .B(n45652), .Z(n45655) );
  XOR U45399 ( .A(n45540), .B(n45656), .Z(n45472) );
  AND U45400 ( .A(n1473), .B(n45657), .Z(n45656) );
  XOR U45401 ( .A(n45536), .B(n45540), .Z(n45657) );
  XOR U45402 ( .A(n45652), .B(n45429), .Z(n45654) );
  XOR U45403 ( .A(n45658), .B(n45659), .Z(n45429) );
  AND U45404 ( .A(n1489), .B(n45660), .Z(n45659) );
  XOR U45405 ( .A(n45661), .B(n45662), .Z(n45652) );
  AND U45406 ( .A(n45663), .B(n45664), .Z(n45662) );
  XNOR U45407 ( .A(n45661), .B(n45480), .Z(n45664) );
  XOR U45408 ( .A(n45591), .B(n45665), .Z(n45480) );
  AND U45409 ( .A(n1473), .B(n45666), .Z(n45665) );
  XOR U45410 ( .A(n45587), .B(n45591), .Z(n45666) );
  XNOR U45411 ( .A(n45667), .B(n45661), .Z(n45663) );
  IV U45412 ( .A(n45439), .Z(n45667) );
  XOR U45413 ( .A(n45668), .B(n45669), .Z(n45439) );
  AND U45414 ( .A(n1489), .B(n45670), .Z(n45669) );
  AND U45415 ( .A(n45632), .B(n45621), .Z(n45661) );
  XNOR U45416 ( .A(n45671), .B(n45672), .Z(n45621) );
  AND U45417 ( .A(n1473), .B(n45603), .Z(n45672) );
  XNOR U45418 ( .A(n45601), .B(n45671), .Z(n45603) );
  XNOR U45419 ( .A(n45673), .B(n45674), .Z(n1473) );
  AND U45420 ( .A(n45675), .B(n45676), .Z(n45674) );
  XNOR U45421 ( .A(n45673), .B(n45492), .Z(n45676) );
  IV U45422 ( .A(n45496), .Z(n45492) );
  XOR U45423 ( .A(n45677), .B(n45678), .Z(n45496) );
  AND U45424 ( .A(n1477), .B(n45679), .Z(n45678) );
  XOR U45425 ( .A(n45680), .B(n45677), .Z(n45679) );
  XNOR U45426 ( .A(n45673), .B(n45608), .Z(n45675) );
  XOR U45427 ( .A(n45681), .B(n45682), .Z(n45608) );
  AND U45428 ( .A(n1485), .B(n45643), .Z(n45682) );
  XOR U45429 ( .A(n45641), .B(n45681), .Z(n45643) );
  XOR U45430 ( .A(n45683), .B(n45684), .Z(n45673) );
  AND U45431 ( .A(n45685), .B(n45686), .Z(n45684) );
  XNOR U45432 ( .A(n45683), .B(n45508), .Z(n45686) );
  IV U45433 ( .A(n45511), .Z(n45508) );
  XOR U45434 ( .A(n45687), .B(n45688), .Z(n45511) );
  AND U45435 ( .A(n1477), .B(n45689), .Z(n45688) );
  XOR U45436 ( .A(n45690), .B(n45687), .Z(n45689) );
  XOR U45437 ( .A(n45512), .B(n45683), .Z(n45685) );
  XOR U45438 ( .A(n45691), .B(n45692), .Z(n45512) );
  AND U45439 ( .A(n1485), .B(n45651), .Z(n45692) );
  XOR U45440 ( .A(n45691), .B(n45649), .Z(n45651) );
  XOR U45441 ( .A(n45693), .B(n45694), .Z(n45683) );
  AND U45442 ( .A(n45695), .B(n45696), .Z(n45694) );
  XNOR U45443 ( .A(n45693), .B(n45536), .Z(n45696) );
  IV U45444 ( .A(n45539), .Z(n45536) );
  XOR U45445 ( .A(n45697), .B(n45698), .Z(n45539) );
  AND U45446 ( .A(n1477), .B(n45699), .Z(n45698) );
  XNOR U45447 ( .A(n45700), .B(n45697), .Z(n45699) );
  XOR U45448 ( .A(n45540), .B(n45693), .Z(n45695) );
  XOR U45449 ( .A(n45701), .B(n45702), .Z(n45540) );
  AND U45450 ( .A(n1485), .B(n45660), .Z(n45702) );
  XOR U45451 ( .A(n45701), .B(n45658), .Z(n45660) );
  XOR U45452 ( .A(n45617), .B(n45703), .Z(n45693) );
  AND U45453 ( .A(n45619), .B(n45704), .Z(n45703) );
  XNOR U45454 ( .A(n45617), .B(n45587), .Z(n45704) );
  IV U45455 ( .A(n45590), .Z(n45587) );
  XOR U45456 ( .A(n45705), .B(n45706), .Z(n45590) );
  AND U45457 ( .A(n1477), .B(n45707), .Z(n45706) );
  XOR U45458 ( .A(n45708), .B(n45705), .Z(n45707) );
  XOR U45459 ( .A(n45591), .B(n45617), .Z(n45619) );
  XOR U45460 ( .A(n45709), .B(n45710), .Z(n45591) );
  AND U45461 ( .A(n1485), .B(n45670), .Z(n45710) );
  XOR U45462 ( .A(n45709), .B(n45668), .Z(n45670) );
  AND U45463 ( .A(n45671), .B(n45601), .Z(n45617) );
  XNOR U45464 ( .A(n45711), .B(n45712), .Z(n45601) );
  AND U45465 ( .A(n1477), .B(n45713), .Z(n45712) );
  XNOR U45466 ( .A(n45714), .B(n45711), .Z(n45713) );
  XNOR U45467 ( .A(n45715), .B(n45716), .Z(n1477) );
  AND U45468 ( .A(n45717), .B(n45718), .Z(n45716) );
  XOR U45469 ( .A(n45680), .B(n45715), .Z(n45718) );
  AND U45470 ( .A(n45719), .B(n45720), .Z(n45680) );
  XNOR U45471 ( .A(n45677), .B(n45715), .Z(n45717) );
  XNOR U45472 ( .A(n45721), .B(n45722), .Z(n45677) );
  AND U45473 ( .A(n1481), .B(n45723), .Z(n45722) );
  XNOR U45474 ( .A(n45724), .B(n45725), .Z(n45723) );
  XOR U45475 ( .A(n45726), .B(n45727), .Z(n45715) );
  AND U45476 ( .A(n45728), .B(n45729), .Z(n45727) );
  XNOR U45477 ( .A(n45726), .B(n45719), .Z(n45729) );
  IV U45478 ( .A(n45690), .Z(n45719) );
  XOR U45479 ( .A(n45730), .B(n45731), .Z(n45690) );
  XOR U45480 ( .A(n45732), .B(n45720), .Z(n45731) );
  AND U45481 ( .A(n45700), .B(n45733), .Z(n45720) );
  AND U45482 ( .A(n45734), .B(n45735), .Z(n45732) );
  XOR U45483 ( .A(n45736), .B(n45730), .Z(n45734) );
  XNOR U45484 ( .A(n45687), .B(n45726), .Z(n45728) );
  XNOR U45485 ( .A(n45737), .B(n45738), .Z(n45687) );
  AND U45486 ( .A(n1481), .B(n45739), .Z(n45738) );
  XNOR U45487 ( .A(n45740), .B(n45741), .Z(n45739) );
  XOR U45488 ( .A(n45742), .B(n45743), .Z(n45726) );
  AND U45489 ( .A(n45744), .B(n45745), .Z(n45743) );
  XNOR U45490 ( .A(n45742), .B(n45700), .Z(n45745) );
  XOR U45491 ( .A(n45746), .B(n45735), .Z(n45700) );
  XNOR U45492 ( .A(n45747), .B(n45730), .Z(n45735) );
  XOR U45493 ( .A(n45748), .B(n45749), .Z(n45730) );
  AND U45494 ( .A(n45750), .B(n45751), .Z(n45749) );
  XOR U45495 ( .A(n45752), .B(n45748), .Z(n45750) );
  XNOR U45496 ( .A(n45753), .B(n45754), .Z(n45747) );
  AND U45497 ( .A(n45755), .B(n45756), .Z(n45754) );
  XOR U45498 ( .A(n45753), .B(n45757), .Z(n45755) );
  XNOR U45499 ( .A(n45736), .B(n45733), .Z(n45746) );
  AND U45500 ( .A(n45758), .B(n45759), .Z(n45733) );
  XOR U45501 ( .A(n45760), .B(n45761), .Z(n45736) );
  AND U45502 ( .A(n45762), .B(n45763), .Z(n45761) );
  XOR U45503 ( .A(n45760), .B(n45764), .Z(n45762) );
  XNOR U45504 ( .A(n45697), .B(n45742), .Z(n45744) );
  XNOR U45505 ( .A(n45765), .B(n45766), .Z(n45697) );
  AND U45506 ( .A(n1481), .B(n45767), .Z(n45766) );
  XNOR U45507 ( .A(n45768), .B(n45769), .Z(n45767) );
  XOR U45508 ( .A(n45770), .B(n45771), .Z(n45742) );
  AND U45509 ( .A(n45772), .B(n45773), .Z(n45771) );
  XNOR U45510 ( .A(n45770), .B(n45758), .Z(n45773) );
  IV U45511 ( .A(n45708), .Z(n45758) );
  XNOR U45512 ( .A(n45774), .B(n45751), .Z(n45708) );
  XNOR U45513 ( .A(n45775), .B(n45757), .Z(n45751) );
  XNOR U45514 ( .A(n45776), .B(n45777), .Z(n45757) );
  NOR U45515 ( .A(n45778), .B(n45779), .Z(n45777) );
  XOR U45516 ( .A(n45776), .B(n45780), .Z(n45778) );
  XNOR U45517 ( .A(n45756), .B(n45748), .Z(n45775) );
  XOR U45518 ( .A(n45781), .B(n45782), .Z(n45748) );
  AND U45519 ( .A(n45783), .B(n45784), .Z(n45782) );
  XOR U45520 ( .A(n45781), .B(n45785), .Z(n45783) );
  XNOR U45521 ( .A(n45786), .B(n45753), .Z(n45756) );
  XOR U45522 ( .A(n45787), .B(n45788), .Z(n45753) );
  AND U45523 ( .A(n45789), .B(n45790), .Z(n45788) );
  XNOR U45524 ( .A(n45791), .B(n45792), .Z(n45789) );
  IV U45525 ( .A(n45787), .Z(n45791) );
  XNOR U45526 ( .A(n45793), .B(n45794), .Z(n45786) );
  NOR U45527 ( .A(n45795), .B(n45796), .Z(n45794) );
  XNOR U45528 ( .A(n45793), .B(n45797), .Z(n45795) );
  XNOR U45529 ( .A(n45752), .B(n45759), .Z(n45774) );
  NOR U45530 ( .A(n45714), .B(n45798), .Z(n45759) );
  XOR U45531 ( .A(n45764), .B(n45763), .Z(n45752) );
  XNOR U45532 ( .A(n45799), .B(n45760), .Z(n45763) );
  XOR U45533 ( .A(n45800), .B(n45801), .Z(n45760) );
  AND U45534 ( .A(n45802), .B(n45803), .Z(n45801) );
  XNOR U45535 ( .A(n45804), .B(n45805), .Z(n45802) );
  IV U45536 ( .A(n45800), .Z(n45804) );
  XNOR U45537 ( .A(n45806), .B(n45807), .Z(n45799) );
  NOR U45538 ( .A(n45808), .B(n45809), .Z(n45807) );
  XNOR U45539 ( .A(n45806), .B(n45810), .Z(n45808) );
  XOR U45540 ( .A(n45811), .B(n45812), .Z(n45764) );
  NOR U45541 ( .A(n45813), .B(n45814), .Z(n45812) );
  XNOR U45542 ( .A(n45811), .B(n45815), .Z(n45813) );
  XNOR U45543 ( .A(n45705), .B(n45770), .Z(n45772) );
  XNOR U45544 ( .A(n45816), .B(n45817), .Z(n45705) );
  AND U45545 ( .A(n1481), .B(n45818), .Z(n45817) );
  XNOR U45546 ( .A(n45819), .B(n45820), .Z(n45818) );
  AND U45547 ( .A(n45711), .B(n45714), .Z(n45770) );
  XOR U45548 ( .A(n45821), .B(n45798), .Z(n45714) );
  XNOR U45549 ( .A(p_input[1184]), .B(p_input[2048]), .Z(n45798) );
  XNOR U45550 ( .A(n45785), .B(n45784), .Z(n45821) );
  XNOR U45551 ( .A(n45822), .B(n45792), .Z(n45784) );
  XNOR U45552 ( .A(n45780), .B(n45779), .Z(n45792) );
  XNOR U45553 ( .A(n45823), .B(n45776), .Z(n45779) );
  XNOR U45554 ( .A(p_input[1194]), .B(p_input[2058]), .Z(n45776) );
  XOR U45555 ( .A(p_input[1195]), .B(n29030), .Z(n45823) );
  XOR U45556 ( .A(p_input[1196]), .B(p_input[2060]), .Z(n45780) );
  XOR U45557 ( .A(n45790), .B(n45824), .Z(n45822) );
  IV U45558 ( .A(n45781), .Z(n45824) );
  XOR U45559 ( .A(p_input[1185]), .B(p_input[2049]), .Z(n45781) );
  XNOR U45560 ( .A(n45825), .B(n45797), .Z(n45790) );
  XNOR U45561 ( .A(p_input[1199]), .B(n29033), .Z(n45797) );
  XOR U45562 ( .A(n45787), .B(n45796), .Z(n45825) );
  XOR U45563 ( .A(n45826), .B(n45793), .Z(n45796) );
  XOR U45564 ( .A(p_input[1197]), .B(p_input[2061]), .Z(n45793) );
  XOR U45565 ( .A(p_input[1198]), .B(n29035), .Z(n45826) );
  XOR U45566 ( .A(p_input[1193]), .B(p_input[2057]), .Z(n45787) );
  XOR U45567 ( .A(n45805), .B(n45803), .Z(n45785) );
  XNOR U45568 ( .A(n45827), .B(n45810), .Z(n45803) );
  XOR U45569 ( .A(p_input[1192]), .B(p_input[2056]), .Z(n45810) );
  XOR U45570 ( .A(n45800), .B(n45809), .Z(n45827) );
  XOR U45571 ( .A(n45828), .B(n45806), .Z(n45809) );
  XOR U45572 ( .A(p_input[1190]), .B(p_input[2054]), .Z(n45806) );
  XOR U45573 ( .A(p_input[1191]), .B(n30404), .Z(n45828) );
  XOR U45574 ( .A(p_input[1186]), .B(p_input[2050]), .Z(n45800) );
  XNOR U45575 ( .A(n45815), .B(n45814), .Z(n45805) );
  XOR U45576 ( .A(n45829), .B(n45811), .Z(n45814) );
  XOR U45577 ( .A(p_input[1187]), .B(p_input[2051]), .Z(n45811) );
  XOR U45578 ( .A(p_input[1188]), .B(n30406), .Z(n45829) );
  XOR U45579 ( .A(p_input[1189]), .B(p_input[2053]), .Z(n45815) );
  XNOR U45580 ( .A(n45830), .B(n45831), .Z(n45711) );
  AND U45581 ( .A(n1481), .B(n45832), .Z(n45831) );
  XNOR U45582 ( .A(n45833), .B(n45834), .Z(n1481) );
  AND U45583 ( .A(n45835), .B(n45836), .Z(n45834) );
  XOR U45584 ( .A(n45725), .B(n45833), .Z(n45836) );
  XNOR U45585 ( .A(n45837), .B(n45833), .Z(n45835) );
  XOR U45586 ( .A(n45838), .B(n45839), .Z(n45833) );
  AND U45587 ( .A(n45840), .B(n45841), .Z(n45839) );
  XOR U45588 ( .A(n45740), .B(n45838), .Z(n45841) );
  XOR U45589 ( .A(n45838), .B(n45741), .Z(n45840) );
  XOR U45590 ( .A(n45842), .B(n45843), .Z(n45838) );
  AND U45591 ( .A(n45844), .B(n45845), .Z(n45843) );
  XOR U45592 ( .A(n45768), .B(n45842), .Z(n45845) );
  XOR U45593 ( .A(n45842), .B(n45769), .Z(n45844) );
  XOR U45594 ( .A(n45846), .B(n45847), .Z(n45842) );
  AND U45595 ( .A(n45848), .B(n45849), .Z(n45847) );
  XOR U45596 ( .A(n45846), .B(n45819), .Z(n45849) );
  XNOR U45597 ( .A(n45850), .B(n45851), .Z(n45671) );
  AND U45598 ( .A(n1485), .B(n45852), .Z(n45851) );
  XNOR U45599 ( .A(n45853), .B(n45854), .Z(n1485) );
  AND U45600 ( .A(n45855), .B(n45856), .Z(n45854) );
  XOR U45601 ( .A(n45853), .B(n45681), .Z(n45856) );
  XNOR U45602 ( .A(n45853), .B(n45641), .Z(n45855) );
  XOR U45603 ( .A(n45857), .B(n45858), .Z(n45853) );
  AND U45604 ( .A(n45859), .B(n45860), .Z(n45858) );
  XOR U45605 ( .A(n45857), .B(n45649), .Z(n45859) );
  XOR U45606 ( .A(n45861), .B(n45862), .Z(n45632) );
  AND U45607 ( .A(n1489), .B(n45852), .Z(n45862) );
  XNOR U45608 ( .A(n45850), .B(n45861), .Z(n45852) );
  XNOR U45609 ( .A(n45863), .B(n45864), .Z(n1489) );
  AND U45610 ( .A(n45865), .B(n45866), .Z(n45864) );
  XNOR U45611 ( .A(n45867), .B(n45863), .Z(n45866) );
  IV U45612 ( .A(n45681), .Z(n45867) );
  XOR U45613 ( .A(n45837), .B(n45868), .Z(n45681) );
  AND U45614 ( .A(n1492), .B(n45869), .Z(n45868) );
  XOR U45615 ( .A(n45724), .B(n45721), .Z(n45869) );
  IV U45616 ( .A(n45837), .Z(n45724) );
  XNOR U45617 ( .A(n45641), .B(n45863), .Z(n45865) );
  XOR U45618 ( .A(n45870), .B(n45871), .Z(n45641) );
  AND U45619 ( .A(n1508), .B(n45872), .Z(n45871) );
  XOR U45620 ( .A(n45857), .B(n45873), .Z(n45863) );
  AND U45621 ( .A(n45874), .B(n45860), .Z(n45873) );
  XNOR U45622 ( .A(n45691), .B(n45857), .Z(n45860) );
  XOR U45623 ( .A(n45741), .B(n45875), .Z(n45691) );
  AND U45624 ( .A(n1492), .B(n45876), .Z(n45875) );
  XOR U45625 ( .A(n45737), .B(n45741), .Z(n45876) );
  XNOR U45626 ( .A(n45877), .B(n45857), .Z(n45874) );
  IV U45627 ( .A(n45649), .Z(n45877) );
  XOR U45628 ( .A(n45878), .B(n45879), .Z(n45649) );
  AND U45629 ( .A(n1508), .B(n45880), .Z(n45879) );
  XOR U45630 ( .A(n45881), .B(n45882), .Z(n45857) );
  AND U45631 ( .A(n45883), .B(n45884), .Z(n45882) );
  XNOR U45632 ( .A(n45701), .B(n45881), .Z(n45884) );
  XOR U45633 ( .A(n45769), .B(n45885), .Z(n45701) );
  AND U45634 ( .A(n1492), .B(n45886), .Z(n45885) );
  XOR U45635 ( .A(n45765), .B(n45769), .Z(n45886) );
  XOR U45636 ( .A(n45881), .B(n45658), .Z(n45883) );
  XOR U45637 ( .A(n45887), .B(n45888), .Z(n45658) );
  AND U45638 ( .A(n1508), .B(n45889), .Z(n45888) );
  XOR U45639 ( .A(n45890), .B(n45891), .Z(n45881) );
  AND U45640 ( .A(n45892), .B(n45893), .Z(n45891) );
  XNOR U45641 ( .A(n45890), .B(n45709), .Z(n45893) );
  XOR U45642 ( .A(n45820), .B(n45894), .Z(n45709) );
  AND U45643 ( .A(n1492), .B(n45895), .Z(n45894) );
  XOR U45644 ( .A(n45816), .B(n45820), .Z(n45895) );
  XNOR U45645 ( .A(n45896), .B(n45890), .Z(n45892) );
  IV U45646 ( .A(n45668), .Z(n45896) );
  XOR U45647 ( .A(n45897), .B(n45898), .Z(n45668) );
  AND U45648 ( .A(n1508), .B(n45899), .Z(n45898) );
  AND U45649 ( .A(n45861), .B(n45850), .Z(n45890) );
  XNOR U45650 ( .A(n45900), .B(n45901), .Z(n45850) );
  AND U45651 ( .A(n1492), .B(n45832), .Z(n45901) );
  XNOR U45652 ( .A(n45830), .B(n45900), .Z(n45832) );
  XNOR U45653 ( .A(n45902), .B(n45903), .Z(n1492) );
  AND U45654 ( .A(n45904), .B(n45905), .Z(n45903) );
  XNOR U45655 ( .A(n45902), .B(n45721), .Z(n45905) );
  IV U45656 ( .A(n45725), .Z(n45721) );
  XOR U45657 ( .A(n45906), .B(n45907), .Z(n45725) );
  AND U45658 ( .A(n1496), .B(n45908), .Z(n45907) );
  XOR U45659 ( .A(n45909), .B(n45906), .Z(n45908) );
  XNOR U45660 ( .A(n45902), .B(n45837), .Z(n45904) );
  XOR U45661 ( .A(n45910), .B(n45911), .Z(n45837) );
  AND U45662 ( .A(n1504), .B(n45872), .Z(n45911) );
  XOR U45663 ( .A(n45870), .B(n45910), .Z(n45872) );
  XOR U45664 ( .A(n45912), .B(n45913), .Z(n45902) );
  AND U45665 ( .A(n45914), .B(n45915), .Z(n45913) );
  XNOR U45666 ( .A(n45912), .B(n45737), .Z(n45915) );
  IV U45667 ( .A(n45740), .Z(n45737) );
  XOR U45668 ( .A(n45916), .B(n45917), .Z(n45740) );
  AND U45669 ( .A(n1496), .B(n45918), .Z(n45917) );
  XOR U45670 ( .A(n45919), .B(n45916), .Z(n45918) );
  XOR U45671 ( .A(n45741), .B(n45912), .Z(n45914) );
  XOR U45672 ( .A(n45920), .B(n45921), .Z(n45741) );
  AND U45673 ( .A(n1504), .B(n45880), .Z(n45921) );
  XOR U45674 ( .A(n45920), .B(n45878), .Z(n45880) );
  XOR U45675 ( .A(n45922), .B(n45923), .Z(n45912) );
  AND U45676 ( .A(n45924), .B(n45925), .Z(n45923) );
  XNOR U45677 ( .A(n45922), .B(n45765), .Z(n45925) );
  IV U45678 ( .A(n45768), .Z(n45765) );
  XOR U45679 ( .A(n45926), .B(n45927), .Z(n45768) );
  AND U45680 ( .A(n1496), .B(n45928), .Z(n45927) );
  XNOR U45681 ( .A(n45929), .B(n45926), .Z(n45928) );
  XOR U45682 ( .A(n45769), .B(n45922), .Z(n45924) );
  XOR U45683 ( .A(n45930), .B(n45931), .Z(n45769) );
  AND U45684 ( .A(n1504), .B(n45889), .Z(n45931) );
  XOR U45685 ( .A(n45930), .B(n45887), .Z(n45889) );
  XOR U45686 ( .A(n45846), .B(n45932), .Z(n45922) );
  AND U45687 ( .A(n45848), .B(n45933), .Z(n45932) );
  XNOR U45688 ( .A(n45846), .B(n45816), .Z(n45933) );
  IV U45689 ( .A(n45819), .Z(n45816) );
  XOR U45690 ( .A(n45934), .B(n45935), .Z(n45819) );
  AND U45691 ( .A(n1496), .B(n45936), .Z(n45935) );
  XOR U45692 ( .A(n45937), .B(n45934), .Z(n45936) );
  XOR U45693 ( .A(n45820), .B(n45846), .Z(n45848) );
  XOR U45694 ( .A(n45938), .B(n45939), .Z(n45820) );
  AND U45695 ( .A(n1504), .B(n45899), .Z(n45939) );
  XOR U45696 ( .A(n45938), .B(n45897), .Z(n45899) );
  AND U45697 ( .A(n45900), .B(n45830), .Z(n45846) );
  XNOR U45698 ( .A(n45940), .B(n45941), .Z(n45830) );
  AND U45699 ( .A(n1496), .B(n45942), .Z(n45941) );
  XNOR U45700 ( .A(n45943), .B(n45940), .Z(n45942) );
  XNOR U45701 ( .A(n45944), .B(n45945), .Z(n1496) );
  AND U45702 ( .A(n45946), .B(n45947), .Z(n45945) );
  XOR U45703 ( .A(n45909), .B(n45944), .Z(n45947) );
  AND U45704 ( .A(n45948), .B(n45949), .Z(n45909) );
  XNOR U45705 ( .A(n45906), .B(n45944), .Z(n45946) );
  XNOR U45706 ( .A(n45950), .B(n45951), .Z(n45906) );
  AND U45707 ( .A(n1500), .B(n45952), .Z(n45951) );
  XNOR U45708 ( .A(n45953), .B(n45954), .Z(n45952) );
  XOR U45709 ( .A(n45955), .B(n45956), .Z(n45944) );
  AND U45710 ( .A(n45957), .B(n45958), .Z(n45956) );
  XNOR U45711 ( .A(n45955), .B(n45948), .Z(n45958) );
  IV U45712 ( .A(n45919), .Z(n45948) );
  XOR U45713 ( .A(n45959), .B(n45960), .Z(n45919) );
  XOR U45714 ( .A(n45961), .B(n45949), .Z(n45960) );
  AND U45715 ( .A(n45929), .B(n45962), .Z(n45949) );
  AND U45716 ( .A(n45963), .B(n45964), .Z(n45961) );
  XOR U45717 ( .A(n45965), .B(n45959), .Z(n45963) );
  XNOR U45718 ( .A(n45916), .B(n45955), .Z(n45957) );
  XNOR U45719 ( .A(n45966), .B(n45967), .Z(n45916) );
  AND U45720 ( .A(n1500), .B(n45968), .Z(n45967) );
  XNOR U45721 ( .A(n45969), .B(n45970), .Z(n45968) );
  XOR U45722 ( .A(n45971), .B(n45972), .Z(n45955) );
  AND U45723 ( .A(n45973), .B(n45974), .Z(n45972) );
  XNOR U45724 ( .A(n45971), .B(n45929), .Z(n45974) );
  XOR U45725 ( .A(n45975), .B(n45964), .Z(n45929) );
  XNOR U45726 ( .A(n45976), .B(n45959), .Z(n45964) );
  XOR U45727 ( .A(n45977), .B(n45978), .Z(n45959) );
  AND U45728 ( .A(n45979), .B(n45980), .Z(n45978) );
  XOR U45729 ( .A(n45981), .B(n45977), .Z(n45979) );
  XNOR U45730 ( .A(n45982), .B(n45983), .Z(n45976) );
  AND U45731 ( .A(n45984), .B(n45985), .Z(n45983) );
  XOR U45732 ( .A(n45982), .B(n45986), .Z(n45984) );
  XNOR U45733 ( .A(n45965), .B(n45962), .Z(n45975) );
  AND U45734 ( .A(n45987), .B(n45988), .Z(n45962) );
  XOR U45735 ( .A(n45989), .B(n45990), .Z(n45965) );
  AND U45736 ( .A(n45991), .B(n45992), .Z(n45990) );
  XOR U45737 ( .A(n45989), .B(n45993), .Z(n45991) );
  XNOR U45738 ( .A(n45926), .B(n45971), .Z(n45973) );
  XNOR U45739 ( .A(n45994), .B(n45995), .Z(n45926) );
  AND U45740 ( .A(n1500), .B(n45996), .Z(n45995) );
  XNOR U45741 ( .A(n45997), .B(n45998), .Z(n45996) );
  XOR U45742 ( .A(n45999), .B(n46000), .Z(n45971) );
  AND U45743 ( .A(n46001), .B(n46002), .Z(n46000) );
  XNOR U45744 ( .A(n45999), .B(n45987), .Z(n46002) );
  IV U45745 ( .A(n45937), .Z(n45987) );
  XNOR U45746 ( .A(n46003), .B(n45980), .Z(n45937) );
  XNOR U45747 ( .A(n46004), .B(n45986), .Z(n45980) );
  XNOR U45748 ( .A(n46005), .B(n46006), .Z(n45986) );
  NOR U45749 ( .A(n46007), .B(n46008), .Z(n46006) );
  XOR U45750 ( .A(n46005), .B(n46009), .Z(n46007) );
  XNOR U45751 ( .A(n45985), .B(n45977), .Z(n46004) );
  XOR U45752 ( .A(n46010), .B(n46011), .Z(n45977) );
  AND U45753 ( .A(n46012), .B(n46013), .Z(n46011) );
  XOR U45754 ( .A(n46010), .B(n46014), .Z(n46012) );
  XNOR U45755 ( .A(n46015), .B(n45982), .Z(n45985) );
  XOR U45756 ( .A(n46016), .B(n46017), .Z(n45982) );
  AND U45757 ( .A(n46018), .B(n46019), .Z(n46017) );
  XNOR U45758 ( .A(n46020), .B(n46021), .Z(n46018) );
  IV U45759 ( .A(n46016), .Z(n46020) );
  XNOR U45760 ( .A(n46022), .B(n46023), .Z(n46015) );
  NOR U45761 ( .A(n46024), .B(n46025), .Z(n46023) );
  XNOR U45762 ( .A(n46022), .B(n46026), .Z(n46024) );
  XNOR U45763 ( .A(n45981), .B(n45988), .Z(n46003) );
  NOR U45764 ( .A(n45943), .B(n46027), .Z(n45988) );
  XOR U45765 ( .A(n45993), .B(n45992), .Z(n45981) );
  XNOR U45766 ( .A(n46028), .B(n45989), .Z(n45992) );
  XOR U45767 ( .A(n46029), .B(n46030), .Z(n45989) );
  AND U45768 ( .A(n46031), .B(n46032), .Z(n46030) );
  XNOR U45769 ( .A(n46033), .B(n46034), .Z(n46031) );
  IV U45770 ( .A(n46029), .Z(n46033) );
  XNOR U45771 ( .A(n46035), .B(n46036), .Z(n46028) );
  NOR U45772 ( .A(n46037), .B(n46038), .Z(n46036) );
  XNOR U45773 ( .A(n46035), .B(n46039), .Z(n46037) );
  XOR U45774 ( .A(n46040), .B(n46041), .Z(n45993) );
  NOR U45775 ( .A(n46042), .B(n46043), .Z(n46041) );
  XNOR U45776 ( .A(n46040), .B(n46044), .Z(n46042) );
  XNOR U45777 ( .A(n45934), .B(n45999), .Z(n46001) );
  XNOR U45778 ( .A(n46045), .B(n46046), .Z(n45934) );
  AND U45779 ( .A(n1500), .B(n46047), .Z(n46046) );
  XNOR U45780 ( .A(n46048), .B(n46049), .Z(n46047) );
  AND U45781 ( .A(n45940), .B(n45943), .Z(n45999) );
  XOR U45782 ( .A(n46050), .B(n46027), .Z(n45943) );
  XNOR U45783 ( .A(p_input[1200]), .B(p_input[2048]), .Z(n46027) );
  XNOR U45784 ( .A(n46014), .B(n46013), .Z(n46050) );
  XNOR U45785 ( .A(n46051), .B(n46021), .Z(n46013) );
  XNOR U45786 ( .A(n46009), .B(n46008), .Z(n46021) );
  XNOR U45787 ( .A(n46052), .B(n46005), .Z(n46008) );
  XNOR U45788 ( .A(p_input[1210]), .B(p_input[2058]), .Z(n46005) );
  XOR U45789 ( .A(p_input[1211]), .B(n29030), .Z(n46052) );
  XOR U45790 ( .A(p_input[1212]), .B(p_input[2060]), .Z(n46009) );
  XOR U45791 ( .A(n46019), .B(n46053), .Z(n46051) );
  IV U45792 ( .A(n46010), .Z(n46053) );
  XOR U45793 ( .A(p_input[1201]), .B(p_input[2049]), .Z(n46010) );
  XNOR U45794 ( .A(n46054), .B(n46026), .Z(n46019) );
  XNOR U45795 ( .A(p_input[1215]), .B(n29033), .Z(n46026) );
  XOR U45796 ( .A(n46016), .B(n46025), .Z(n46054) );
  XOR U45797 ( .A(n46055), .B(n46022), .Z(n46025) );
  XOR U45798 ( .A(p_input[1213]), .B(p_input[2061]), .Z(n46022) );
  XOR U45799 ( .A(p_input[1214]), .B(n29035), .Z(n46055) );
  XOR U45800 ( .A(p_input[1209]), .B(p_input[2057]), .Z(n46016) );
  XOR U45801 ( .A(n46034), .B(n46032), .Z(n46014) );
  XNOR U45802 ( .A(n46056), .B(n46039), .Z(n46032) );
  XOR U45803 ( .A(p_input[1208]), .B(p_input[2056]), .Z(n46039) );
  XOR U45804 ( .A(n46029), .B(n46038), .Z(n46056) );
  XOR U45805 ( .A(n46057), .B(n46035), .Z(n46038) );
  XOR U45806 ( .A(p_input[1206]), .B(p_input[2054]), .Z(n46035) );
  XOR U45807 ( .A(p_input[1207]), .B(n30404), .Z(n46057) );
  XOR U45808 ( .A(p_input[1202]), .B(p_input[2050]), .Z(n46029) );
  XNOR U45809 ( .A(n46044), .B(n46043), .Z(n46034) );
  XOR U45810 ( .A(n46058), .B(n46040), .Z(n46043) );
  XOR U45811 ( .A(p_input[1203]), .B(p_input[2051]), .Z(n46040) );
  XOR U45812 ( .A(p_input[1204]), .B(n30406), .Z(n46058) );
  XOR U45813 ( .A(p_input[1205]), .B(p_input[2053]), .Z(n46044) );
  XNOR U45814 ( .A(n46059), .B(n46060), .Z(n45940) );
  AND U45815 ( .A(n1500), .B(n46061), .Z(n46060) );
  XNOR U45816 ( .A(n46062), .B(n46063), .Z(n1500) );
  AND U45817 ( .A(n46064), .B(n46065), .Z(n46063) );
  XOR U45818 ( .A(n45954), .B(n46062), .Z(n46065) );
  XNOR U45819 ( .A(n46066), .B(n46062), .Z(n46064) );
  XOR U45820 ( .A(n46067), .B(n46068), .Z(n46062) );
  AND U45821 ( .A(n46069), .B(n46070), .Z(n46068) );
  XOR U45822 ( .A(n45969), .B(n46067), .Z(n46070) );
  XOR U45823 ( .A(n46067), .B(n45970), .Z(n46069) );
  XOR U45824 ( .A(n46071), .B(n46072), .Z(n46067) );
  AND U45825 ( .A(n46073), .B(n46074), .Z(n46072) );
  XOR U45826 ( .A(n45997), .B(n46071), .Z(n46074) );
  XOR U45827 ( .A(n46071), .B(n45998), .Z(n46073) );
  XOR U45828 ( .A(n46075), .B(n46076), .Z(n46071) );
  AND U45829 ( .A(n46077), .B(n46078), .Z(n46076) );
  XOR U45830 ( .A(n46075), .B(n46048), .Z(n46078) );
  XNOR U45831 ( .A(n46079), .B(n46080), .Z(n45900) );
  AND U45832 ( .A(n1504), .B(n46081), .Z(n46080) );
  XNOR U45833 ( .A(n46082), .B(n46083), .Z(n1504) );
  AND U45834 ( .A(n46084), .B(n46085), .Z(n46083) );
  XOR U45835 ( .A(n46082), .B(n45910), .Z(n46085) );
  XNOR U45836 ( .A(n46082), .B(n45870), .Z(n46084) );
  XOR U45837 ( .A(n46086), .B(n46087), .Z(n46082) );
  AND U45838 ( .A(n46088), .B(n46089), .Z(n46087) );
  XOR U45839 ( .A(n46086), .B(n45878), .Z(n46088) );
  XOR U45840 ( .A(n46090), .B(n46091), .Z(n45861) );
  AND U45841 ( .A(n1508), .B(n46081), .Z(n46091) );
  XNOR U45842 ( .A(n46079), .B(n46090), .Z(n46081) );
  XNOR U45843 ( .A(n46092), .B(n46093), .Z(n1508) );
  AND U45844 ( .A(n46094), .B(n46095), .Z(n46093) );
  XNOR U45845 ( .A(n46096), .B(n46092), .Z(n46095) );
  IV U45846 ( .A(n45910), .Z(n46096) );
  XOR U45847 ( .A(n46066), .B(n46097), .Z(n45910) );
  AND U45848 ( .A(n1511), .B(n46098), .Z(n46097) );
  XOR U45849 ( .A(n45953), .B(n45950), .Z(n46098) );
  IV U45850 ( .A(n46066), .Z(n45953) );
  XNOR U45851 ( .A(n45870), .B(n46092), .Z(n46094) );
  XOR U45852 ( .A(n46099), .B(n46100), .Z(n45870) );
  AND U45853 ( .A(n1527), .B(n46101), .Z(n46100) );
  XOR U45854 ( .A(n46086), .B(n46102), .Z(n46092) );
  AND U45855 ( .A(n46103), .B(n46089), .Z(n46102) );
  XNOR U45856 ( .A(n45920), .B(n46086), .Z(n46089) );
  XOR U45857 ( .A(n45970), .B(n46104), .Z(n45920) );
  AND U45858 ( .A(n1511), .B(n46105), .Z(n46104) );
  XOR U45859 ( .A(n45966), .B(n45970), .Z(n46105) );
  XNOR U45860 ( .A(n46106), .B(n46086), .Z(n46103) );
  IV U45861 ( .A(n45878), .Z(n46106) );
  XOR U45862 ( .A(n46107), .B(n46108), .Z(n45878) );
  AND U45863 ( .A(n1527), .B(n46109), .Z(n46108) );
  XOR U45864 ( .A(n46110), .B(n46111), .Z(n46086) );
  AND U45865 ( .A(n46112), .B(n46113), .Z(n46111) );
  XNOR U45866 ( .A(n45930), .B(n46110), .Z(n46113) );
  XOR U45867 ( .A(n45998), .B(n46114), .Z(n45930) );
  AND U45868 ( .A(n1511), .B(n46115), .Z(n46114) );
  XOR U45869 ( .A(n45994), .B(n45998), .Z(n46115) );
  XOR U45870 ( .A(n46110), .B(n45887), .Z(n46112) );
  XOR U45871 ( .A(n46116), .B(n46117), .Z(n45887) );
  AND U45872 ( .A(n1527), .B(n46118), .Z(n46117) );
  XOR U45873 ( .A(n46119), .B(n46120), .Z(n46110) );
  AND U45874 ( .A(n46121), .B(n46122), .Z(n46120) );
  XNOR U45875 ( .A(n46119), .B(n45938), .Z(n46122) );
  XOR U45876 ( .A(n46049), .B(n46123), .Z(n45938) );
  AND U45877 ( .A(n1511), .B(n46124), .Z(n46123) );
  XOR U45878 ( .A(n46045), .B(n46049), .Z(n46124) );
  XNOR U45879 ( .A(n46125), .B(n46119), .Z(n46121) );
  IV U45880 ( .A(n45897), .Z(n46125) );
  XOR U45881 ( .A(n46126), .B(n46127), .Z(n45897) );
  AND U45882 ( .A(n1527), .B(n46128), .Z(n46127) );
  AND U45883 ( .A(n46090), .B(n46079), .Z(n46119) );
  XNOR U45884 ( .A(n46129), .B(n46130), .Z(n46079) );
  AND U45885 ( .A(n1511), .B(n46061), .Z(n46130) );
  XNOR U45886 ( .A(n46059), .B(n46129), .Z(n46061) );
  XNOR U45887 ( .A(n46131), .B(n46132), .Z(n1511) );
  AND U45888 ( .A(n46133), .B(n46134), .Z(n46132) );
  XNOR U45889 ( .A(n46131), .B(n45950), .Z(n46134) );
  IV U45890 ( .A(n45954), .Z(n45950) );
  XOR U45891 ( .A(n46135), .B(n46136), .Z(n45954) );
  AND U45892 ( .A(n1515), .B(n46137), .Z(n46136) );
  XOR U45893 ( .A(n46138), .B(n46135), .Z(n46137) );
  XNOR U45894 ( .A(n46131), .B(n46066), .Z(n46133) );
  XOR U45895 ( .A(n46139), .B(n46140), .Z(n46066) );
  AND U45896 ( .A(n1523), .B(n46101), .Z(n46140) );
  XOR U45897 ( .A(n46099), .B(n46139), .Z(n46101) );
  XOR U45898 ( .A(n46141), .B(n46142), .Z(n46131) );
  AND U45899 ( .A(n46143), .B(n46144), .Z(n46142) );
  XNOR U45900 ( .A(n46141), .B(n45966), .Z(n46144) );
  IV U45901 ( .A(n45969), .Z(n45966) );
  XOR U45902 ( .A(n46145), .B(n46146), .Z(n45969) );
  AND U45903 ( .A(n1515), .B(n46147), .Z(n46146) );
  XOR U45904 ( .A(n46148), .B(n46145), .Z(n46147) );
  XOR U45905 ( .A(n45970), .B(n46141), .Z(n46143) );
  XOR U45906 ( .A(n46149), .B(n46150), .Z(n45970) );
  AND U45907 ( .A(n1523), .B(n46109), .Z(n46150) );
  XOR U45908 ( .A(n46149), .B(n46107), .Z(n46109) );
  XOR U45909 ( .A(n46151), .B(n46152), .Z(n46141) );
  AND U45910 ( .A(n46153), .B(n46154), .Z(n46152) );
  XNOR U45911 ( .A(n46151), .B(n45994), .Z(n46154) );
  IV U45912 ( .A(n45997), .Z(n45994) );
  XOR U45913 ( .A(n46155), .B(n46156), .Z(n45997) );
  AND U45914 ( .A(n1515), .B(n46157), .Z(n46156) );
  XNOR U45915 ( .A(n46158), .B(n46155), .Z(n46157) );
  XOR U45916 ( .A(n45998), .B(n46151), .Z(n46153) );
  XOR U45917 ( .A(n46159), .B(n46160), .Z(n45998) );
  AND U45918 ( .A(n1523), .B(n46118), .Z(n46160) );
  XOR U45919 ( .A(n46159), .B(n46116), .Z(n46118) );
  XOR U45920 ( .A(n46075), .B(n46161), .Z(n46151) );
  AND U45921 ( .A(n46077), .B(n46162), .Z(n46161) );
  XNOR U45922 ( .A(n46075), .B(n46045), .Z(n46162) );
  IV U45923 ( .A(n46048), .Z(n46045) );
  XOR U45924 ( .A(n46163), .B(n46164), .Z(n46048) );
  AND U45925 ( .A(n1515), .B(n46165), .Z(n46164) );
  XOR U45926 ( .A(n46166), .B(n46163), .Z(n46165) );
  XOR U45927 ( .A(n46049), .B(n46075), .Z(n46077) );
  XOR U45928 ( .A(n46167), .B(n46168), .Z(n46049) );
  AND U45929 ( .A(n1523), .B(n46128), .Z(n46168) );
  XOR U45930 ( .A(n46167), .B(n46126), .Z(n46128) );
  AND U45931 ( .A(n46129), .B(n46059), .Z(n46075) );
  XNOR U45932 ( .A(n46169), .B(n46170), .Z(n46059) );
  AND U45933 ( .A(n1515), .B(n46171), .Z(n46170) );
  XNOR U45934 ( .A(n46172), .B(n46169), .Z(n46171) );
  XNOR U45935 ( .A(n46173), .B(n46174), .Z(n1515) );
  AND U45936 ( .A(n46175), .B(n46176), .Z(n46174) );
  XOR U45937 ( .A(n46138), .B(n46173), .Z(n46176) );
  AND U45938 ( .A(n46177), .B(n46178), .Z(n46138) );
  XNOR U45939 ( .A(n46135), .B(n46173), .Z(n46175) );
  XNOR U45940 ( .A(n46179), .B(n46180), .Z(n46135) );
  AND U45941 ( .A(n1519), .B(n46181), .Z(n46180) );
  XNOR U45942 ( .A(n46182), .B(n46183), .Z(n46181) );
  XOR U45943 ( .A(n46184), .B(n46185), .Z(n46173) );
  AND U45944 ( .A(n46186), .B(n46187), .Z(n46185) );
  XNOR U45945 ( .A(n46184), .B(n46177), .Z(n46187) );
  IV U45946 ( .A(n46148), .Z(n46177) );
  XOR U45947 ( .A(n46188), .B(n46189), .Z(n46148) );
  XOR U45948 ( .A(n46190), .B(n46178), .Z(n46189) );
  AND U45949 ( .A(n46158), .B(n46191), .Z(n46178) );
  AND U45950 ( .A(n46192), .B(n46193), .Z(n46190) );
  XOR U45951 ( .A(n46194), .B(n46188), .Z(n46192) );
  XNOR U45952 ( .A(n46145), .B(n46184), .Z(n46186) );
  XNOR U45953 ( .A(n46195), .B(n46196), .Z(n46145) );
  AND U45954 ( .A(n1519), .B(n46197), .Z(n46196) );
  XNOR U45955 ( .A(n46198), .B(n46199), .Z(n46197) );
  XOR U45956 ( .A(n46200), .B(n46201), .Z(n46184) );
  AND U45957 ( .A(n46202), .B(n46203), .Z(n46201) );
  XNOR U45958 ( .A(n46200), .B(n46158), .Z(n46203) );
  XOR U45959 ( .A(n46204), .B(n46193), .Z(n46158) );
  XNOR U45960 ( .A(n46205), .B(n46188), .Z(n46193) );
  XOR U45961 ( .A(n46206), .B(n46207), .Z(n46188) );
  AND U45962 ( .A(n46208), .B(n46209), .Z(n46207) );
  XOR U45963 ( .A(n46210), .B(n46206), .Z(n46208) );
  XNOR U45964 ( .A(n46211), .B(n46212), .Z(n46205) );
  AND U45965 ( .A(n46213), .B(n46214), .Z(n46212) );
  XOR U45966 ( .A(n46211), .B(n46215), .Z(n46213) );
  XNOR U45967 ( .A(n46194), .B(n46191), .Z(n46204) );
  AND U45968 ( .A(n46216), .B(n46217), .Z(n46191) );
  XOR U45969 ( .A(n46218), .B(n46219), .Z(n46194) );
  AND U45970 ( .A(n46220), .B(n46221), .Z(n46219) );
  XOR U45971 ( .A(n46218), .B(n46222), .Z(n46220) );
  XNOR U45972 ( .A(n46155), .B(n46200), .Z(n46202) );
  XNOR U45973 ( .A(n46223), .B(n46224), .Z(n46155) );
  AND U45974 ( .A(n1519), .B(n46225), .Z(n46224) );
  XNOR U45975 ( .A(n46226), .B(n46227), .Z(n46225) );
  XOR U45976 ( .A(n46228), .B(n46229), .Z(n46200) );
  AND U45977 ( .A(n46230), .B(n46231), .Z(n46229) );
  XNOR U45978 ( .A(n46228), .B(n46216), .Z(n46231) );
  IV U45979 ( .A(n46166), .Z(n46216) );
  XNOR U45980 ( .A(n46232), .B(n46209), .Z(n46166) );
  XNOR U45981 ( .A(n46233), .B(n46215), .Z(n46209) );
  XNOR U45982 ( .A(n46234), .B(n46235), .Z(n46215) );
  NOR U45983 ( .A(n46236), .B(n46237), .Z(n46235) );
  XOR U45984 ( .A(n46234), .B(n46238), .Z(n46236) );
  XNOR U45985 ( .A(n46214), .B(n46206), .Z(n46233) );
  XOR U45986 ( .A(n46239), .B(n46240), .Z(n46206) );
  AND U45987 ( .A(n46241), .B(n46242), .Z(n46240) );
  XOR U45988 ( .A(n46239), .B(n46243), .Z(n46241) );
  XNOR U45989 ( .A(n46244), .B(n46211), .Z(n46214) );
  XOR U45990 ( .A(n46245), .B(n46246), .Z(n46211) );
  AND U45991 ( .A(n46247), .B(n46248), .Z(n46246) );
  XNOR U45992 ( .A(n46249), .B(n46250), .Z(n46247) );
  IV U45993 ( .A(n46245), .Z(n46249) );
  XNOR U45994 ( .A(n46251), .B(n46252), .Z(n46244) );
  NOR U45995 ( .A(n46253), .B(n46254), .Z(n46252) );
  XNOR U45996 ( .A(n46251), .B(n46255), .Z(n46253) );
  XNOR U45997 ( .A(n46210), .B(n46217), .Z(n46232) );
  NOR U45998 ( .A(n46172), .B(n46256), .Z(n46217) );
  XOR U45999 ( .A(n46222), .B(n46221), .Z(n46210) );
  XNOR U46000 ( .A(n46257), .B(n46218), .Z(n46221) );
  XOR U46001 ( .A(n46258), .B(n46259), .Z(n46218) );
  AND U46002 ( .A(n46260), .B(n46261), .Z(n46259) );
  XNOR U46003 ( .A(n46262), .B(n46263), .Z(n46260) );
  IV U46004 ( .A(n46258), .Z(n46262) );
  XNOR U46005 ( .A(n46264), .B(n46265), .Z(n46257) );
  NOR U46006 ( .A(n46266), .B(n46267), .Z(n46265) );
  XNOR U46007 ( .A(n46264), .B(n46268), .Z(n46266) );
  XOR U46008 ( .A(n46269), .B(n46270), .Z(n46222) );
  NOR U46009 ( .A(n46271), .B(n46272), .Z(n46270) );
  XNOR U46010 ( .A(n46269), .B(n46273), .Z(n46271) );
  XNOR U46011 ( .A(n46163), .B(n46228), .Z(n46230) );
  XNOR U46012 ( .A(n46274), .B(n46275), .Z(n46163) );
  AND U46013 ( .A(n1519), .B(n46276), .Z(n46275) );
  XNOR U46014 ( .A(n46277), .B(n46278), .Z(n46276) );
  AND U46015 ( .A(n46169), .B(n46172), .Z(n46228) );
  XOR U46016 ( .A(n46279), .B(n46256), .Z(n46172) );
  XNOR U46017 ( .A(p_input[1216]), .B(p_input[2048]), .Z(n46256) );
  XNOR U46018 ( .A(n46243), .B(n46242), .Z(n46279) );
  XNOR U46019 ( .A(n46280), .B(n46250), .Z(n46242) );
  XNOR U46020 ( .A(n46238), .B(n46237), .Z(n46250) );
  XNOR U46021 ( .A(n46281), .B(n46234), .Z(n46237) );
  XNOR U46022 ( .A(p_input[1226]), .B(p_input[2058]), .Z(n46234) );
  XOR U46023 ( .A(p_input[1227]), .B(n29030), .Z(n46281) );
  XOR U46024 ( .A(p_input[1228]), .B(p_input[2060]), .Z(n46238) );
  XOR U46025 ( .A(n46248), .B(n46282), .Z(n46280) );
  IV U46026 ( .A(n46239), .Z(n46282) );
  XOR U46027 ( .A(p_input[1217]), .B(p_input[2049]), .Z(n46239) );
  XNOR U46028 ( .A(n46283), .B(n46255), .Z(n46248) );
  XNOR U46029 ( .A(p_input[1231]), .B(n29033), .Z(n46255) );
  XOR U46030 ( .A(n46245), .B(n46254), .Z(n46283) );
  XOR U46031 ( .A(n46284), .B(n46251), .Z(n46254) );
  XOR U46032 ( .A(p_input[1229]), .B(p_input[2061]), .Z(n46251) );
  XOR U46033 ( .A(p_input[1230]), .B(n29035), .Z(n46284) );
  XOR U46034 ( .A(p_input[1225]), .B(p_input[2057]), .Z(n46245) );
  XOR U46035 ( .A(n46263), .B(n46261), .Z(n46243) );
  XNOR U46036 ( .A(n46285), .B(n46268), .Z(n46261) );
  XOR U46037 ( .A(p_input[1224]), .B(p_input[2056]), .Z(n46268) );
  XOR U46038 ( .A(n46258), .B(n46267), .Z(n46285) );
  XOR U46039 ( .A(n46286), .B(n46264), .Z(n46267) );
  XOR U46040 ( .A(p_input[1222]), .B(p_input[2054]), .Z(n46264) );
  XOR U46041 ( .A(p_input[1223]), .B(n30404), .Z(n46286) );
  XOR U46042 ( .A(p_input[1218]), .B(p_input[2050]), .Z(n46258) );
  XNOR U46043 ( .A(n46273), .B(n46272), .Z(n46263) );
  XOR U46044 ( .A(n46287), .B(n46269), .Z(n46272) );
  XOR U46045 ( .A(p_input[1219]), .B(p_input[2051]), .Z(n46269) );
  XOR U46046 ( .A(p_input[1220]), .B(n30406), .Z(n46287) );
  XOR U46047 ( .A(p_input[1221]), .B(p_input[2053]), .Z(n46273) );
  XNOR U46048 ( .A(n46288), .B(n46289), .Z(n46169) );
  AND U46049 ( .A(n1519), .B(n46290), .Z(n46289) );
  XNOR U46050 ( .A(n46291), .B(n46292), .Z(n1519) );
  AND U46051 ( .A(n46293), .B(n46294), .Z(n46292) );
  XOR U46052 ( .A(n46183), .B(n46291), .Z(n46294) );
  XNOR U46053 ( .A(n46295), .B(n46291), .Z(n46293) );
  XOR U46054 ( .A(n46296), .B(n46297), .Z(n46291) );
  AND U46055 ( .A(n46298), .B(n46299), .Z(n46297) );
  XOR U46056 ( .A(n46198), .B(n46296), .Z(n46299) );
  XOR U46057 ( .A(n46296), .B(n46199), .Z(n46298) );
  XOR U46058 ( .A(n46300), .B(n46301), .Z(n46296) );
  AND U46059 ( .A(n46302), .B(n46303), .Z(n46301) );
  XOR U46060 ( .A(n46226), .B(n46300), .Z(n46303) );
  XOR U46061 ( .A(n46300), .B(n46227), .Z(n46302) );
  XOR U46062 ( .A(n46304), .B(n46305), .Z(n46300) );
  AND U46063 ( .A(n46306), .B(n46307), .Z(n46305) );
  XOR U46064 ( .A(n46304), .B(n46277), .Z(n46307) );
  XNOR U46065 ( .A(n46308), .B(n46309), .Z(n46129) );
  AND U46066 ( .A(n1523), .B(n46310), .Z(n46309) );
  XNOR U46067 ( .A(n46311), .B(n46312), .Z(n1523) );
  AND U46068 ( .A(n46313), .B(n46314), .Z(n46312) );
  XOR U46069 ( .A(n46311), .B(n46139), .Z(n46314) );
  XNOR U46070 ( .A(n46311), .B(n46099), .Z(n46313) );
  XOR U46071 ( .A(n46315), .B(n46316), .Z(n46311) );
  AND U46072 ( .A(n46317), .B(n46318), .Z(n46316) );
  XOR U46073 ( .A(n46315), .B(n46107), .Z(n46317) );
  XOR U46074 ( .A(n46319), .B(n46320), .Z(n46090) );
  AND U46075 ( .A(n1527), .B(n46310), .Z(n46320) );
  XNOR U46076 ( .A(n46308), .B(n46319), .Z(n46310) );
  XNOR U46077 ( .A(n46321), .B(n46322), .Z(n1527) );
  AND U46078 ( .A(n46323), .B(n46324), .Z(n46322) );
  XNOR U46079 ( .A(n46325), .B(n46321), .Z(n46324) );
  IV U46080 ( .A(n46139), .Z(n46325) );
  XOR U46081 ( .A(n46295), .B(n46326), .Z(n46139) );
  AND U46082 ( .A(n1530), .B(n46327), .Z(n46326) );
  XOR U46083 ( .A(n46182), .B(n46179), .Z(n46327) );
  IV U46084 ( .A(n46295), .Z(n46182) );
  XNOR U46085 ( .A(n46099), .B(n46321), .Z(n46323) );
  XOR U46086 ( .A(n46328), .B(n46329), .Z(n46099) );
  AND U46087 ( .A(n1546), .B(n46330), .Z(n46329) );
  XOR U46088 ( .A(n46315), .B(n46331), .Z(n46321) );
  AND U46089 ( .A(n46332), .B(n46318), .Z(n46331) );
  XNOR U46090 ( .A(n46149), .B(n46315), .Z(n46318) );
  XOR U46091 ( .A(n46199), .B(n46333), .Z(n46149) );
  AND U46092 ( .A(n1530), .B(n46334), .Z(n46333) );
  XOR U46093 ( .A(n46195), .B(n46199), .Z(n46334) );
  XNOR U46094 ( .A(n46335), .B(n46315), .Z(n46332) );
  IV U46095 ( .A(n46107), .Z(n46335) );
  XOR U46096 ( .A(n46336), .B(n46337), .Z(n46107) );
  AND U46097 ( .A(n1546), .B(n46338), .Z(n46337) );
  XOR U46098 ( .A(n46339), .B(n46340), .Z(n46315) );
  AND U46099 ( .A(n46341), .B(n46342), .Z(n46340) );
  XNOR U46100 ( .A(n46159), .B(n46339), .Z(n46342) );
  XOR U46101 ( .A(n46227), .B(n46343), .Z(n46159) );
  AND U46102 ( .A(n1530), .B(n46344), .Z(n46343) );
  XOR U46103 ( .A(n46223), .B(n46227), .Z(n46344) );
  XOR U46104 ( .A(n46339), .B(n46116), .Z(n46341) );
  XOR U46105 ( .A(n46345), .B(n46346), .Z(n46116) );
  AND U46106 ( .A(n1546), .B(n46347), .Z(n46346) );
  XOR U46107 ( .A(n46348), .B(n46349), .Z(n46339) );
  AND U46108 ( .A(n46350), .B(n46351), .Z(n46349) );
  XNOR U46109 ( .A(n46348), .B(n46167), .Z(n46351) );
  XOR U46110 ( .A(n46278), .B(n46352), .Z(n46167) );
  AND U46111 ( .A(n1530), .B(n46353), .Z(n46352) );
  XOR U46112 ( .A(n46274), .B(n46278), .Z(n46353) );
  XNOR U46113 ( .A(n46354), .B(n46348), .Z(n46350) );
  IV U46114 ( .A(n46126), .Z(n46354) );
  XOR U46115 ( .A(n46355), .B(n46356), .Z(n46126) );
  AND U46116 ( .A(n1546), .B(n46357), .Z(n46356) );
  AND U46117 ( .A(n46319), .B(n46308), .Z(n46348) );
  XNOR U46118 ( .A(n46358), .B(n46359), .Z(n46308) );
  AND U46119 ( .A(n1530), .B(n46290), .Z(n46359) );
  XNOR U46120 ( .A(n46288), .B(n46358), .Z(n46290) );
  XNOR U46121 ( .A(n46360), .B(n46361), .Z(n1530) );
  AND U46122 ( .A(n46362), .B(n46363), .Z(n46361) );
  XNOR U46123 ( .A(n46360), .B(n46179), .Z(n46363) );
  IV U46124 ( .A(n46183), .Z(n46179) );
  XOR U46125 ( .A(n46364), .B(n46365), .Z(n46183) );
  AND U46126 ( .A(n1534), .B(n46366), .Z(n46365) );
  XOR U46127 ( .A(n46367), .B(n46364), .Z(n46366) );
  XNOR U46128 ( .A(n46360), .B(n46295), .Z(n46362) );
  XOR U46129 ( .A(n46368), .B(n46369), .Z(n46295) );
  AND U46130 ( .A(n1542), .B(n46330), .Z(n46369) );
  XOR U46131 ( .A(n46328), .B(n46368), .Z(n46330) );
  XOR U46132 ( .A(n46370), .B(n46371), .Z(n46360) );
  AND U46133 ( .A(n46372), .B(n46373), .Z(n46371) );
  XNOR U46134 ( .A(n46370), .B(n46195), .Z(n46373) );
  IV U46135 ( .A(n46198), .Z(n46195) );
  XOR U46136 ( .A(n46374), .B(n46375), .Z(n46198) );
  AND U46137 ( .A(n1534), .B(n46376), .Z(n46375) );
  XOR U46138 ( .A(n46377), .B(n46374), .Z(n46376) );
  XOR U46139 ( .A(n46199), .B(n46370), .Z(n46372) );
  XOR U46140 ( .A(n46378), .B(n46379), .Z(n46199) );
  AND U46141 ( .A(n1542), .B(n46338), .Z(n46379) );
  XOR U46142 ( .A(n46378), .B(n46336), .Z(n46338) );
  XOR U46143 ( .A(n46380), .B(n46381), .Z(n46370) );
  AND U46144 ( .A(n46382), .B(n46383), .Z(n46381) );
  XNOR U46145 ( .A(n46380), .B(n46223), .Z(n46383) );
  IV U46146 ( .A(n46226), .Z(n46223) );
  XOR U46147 ( .A(n46384), .B(n46385), .Z(n46226) );
  AND U46148 ( .A(n1534), .B(n46386), .Z(n46385) );
  XNOR U46149 ( .A(n46387), .B(n46384), .Z(n46386) );
  XOR U46150 ( .A(n46227), .B(n46380), .Z(n46382) );
  XOR U46151 ( .A(n46388), .B(n46389), .Z(n46227) );
  AND U46152 ( .A(n1542), .B(n46347), .Z(n46389) );
  XOR U46153 ( .A(n46388), .B(n46345), .Z(n46347) );
  XOR U46154 ( .A(n46304), .B(n46390), .Z(n46380) );
  AND U46155 ( .A(n46306), .B(n46391), .Z(n46390) );
  XNOR U46156 ( .A(n46304), .B(n46274), .Z(n46391) );
  IV U46157 ( .A(n46277), .Z(n46274) );
  XOR U46158 ( .A(n46392), .B(n46393), .Z(n46277) );
  AND U46159 ( .A(n1534), .B(n46394), .Z(n46393) );
  XOR U46160 ( .A(n46395), .B(n46392), .Z(n46394) );
  XOR U46161 ( .A(n46278), .B(n46304), .Z(n46306) );
  XOR U46162 ( .A(n46396), .B(n46397), .Z(n46278) );
  AND U46163 ( .A(n1542), .B(n46357), .Z(n46397) );
  XOR U46164 ( .A(n46396), .B(n46355), .Z(n46357) );
  AND U46165 ( .A(n46358), .B(n46288), .Z(n46304) );
  XNOR U46166 ( .A(n46398), .B(n46399), .Z(n46288) );
  AND U46167 ( .A(n1534), .B(n46400), .Z(n46399) );
  XNOR U46168 ( .A(n46401), .B(n46398), .Z(n46400) );
  XNOR U46169 ( .A(n46402), .B(n46403), .Z(n1534) );
  AND U46170 ( .A(n46404), .B(n46405), .Z(n46403) );
  XOR U46171 ( .A(n46367), .B(n46402), .Z(n46405) );
  AND U46172 ( .A(n46406), .B(n46407), .Z(n46367) );
  XNOR U46173 ( .A(n46364), .B(n46402), .Z(n46404) );
  XNOR U46174 ( .A(n46408), .B(n46409), .Z(n46364) );
  AND U46175 ( .A(n1538), .B(n46410), .Z(n46409) );
  XNOR U46176 ( .A(n46411), .B(n46412), .Z(n46410) );
  XOR U46177 ( .A(n46413), .B(n46414), .Z(n46402) );
  AND U46178 ( .A(n46415), .B(n46416), .Z(n46414) );
  XNOR U46179 ( .A(n46413), .B(n46406), .Z(n46416) );
  IV U46180 ( .A(n46377), .Z(n46406) );
  XOR U46181 ( .A(n46417), .B(n46418), .Z(n46377) );
  XOR U46182 ( .A(n46419), .B(n46407), .Z(n46418) );
  AND U46183 ( .A(n46387), .B(n46420), .Z(n46407) );
  AND U46184 ( .A(n46421), .B(n46422), .Z(n46419) );
  XOR U46185 ( .A(n46423), .B(n46417), .Z(n46421) );
  XNOR U46186 ( .A(n46374), .B(n46413), .Z(n46415) );
  XNOR U46187 ( .A(n46424), .B(n46425), .Z(n46374) );
  AND U46188 ( .A(n1538), .B(n46426), .Z(n46425) );
  XNOR U46189 ( .A(n46427), .B(n46428), .Z(n46426) );
  XOR U46190 ( .A(n46429), .B(n46430), .Z(n46413) );
  AND U46191 ( .A(n46431), .B(n46432), .Z(n46430) );
  XNOR U46192 ( .A(n46429), .B(n46387), .Z(n46432) );
  XOR U46193 ( .A(n46433), .B(n46422), .Z(n46387) );
  XNOR U46194 ( .A(n46434), .B(n46417), .Z(n46422) );
  XOR U46195 ( .A(n46435), .B(n46436), .Z(n46417) );
  AND U46196 ( .A(n46437), .B(n46438), .Z(n46436) );
  XOR U46197 ( .A(n46439), .B(n46435), .Z(n46437) );
  XNOR U46198 ( .A(n46440), .B(n46441), .Z(n46434) );
  AND U46199 ( .A(n46442), .B(n46443), .Z(n46441) );
  XOR U46200 ( .A(n46440), .B(n46444), .Z(n46442) );
  XNOR U46201 ( .A(n46423), .B(n46420), .Z(n46433) );
  AND U46202 ( .A(n46445), .B(n46446), .Z(n46420) );
  XOR U46203 ( .A(n46447), .B(n46448), .Z(n46423) );
  AND U46204 ( .A(n46449), .B(n46450), .Z(n46448) );
  XOR U46205 ( .A(n46447), .B(n46451), .Z(n46449) );
  XNOR U46206 ( .A(n46384), .B(n46429), .Z(n46431) );
  XNOR U46207 ( .A(n46452), .B(n46453), .Z(n46384) );
  AND U46208 ( .A(n1538), .B(n46454), .Z(n46453) );
  XNOR U46209 ( .A(n46455), .B(n46456), .Z(n46454) );
  XOR U46210 ( .A(n46457), .B(n46458), .Z(n46429) );
  AND U46211 ( .A(n46459), .B(n46460), .Z(n46458) );
  XNOR U46212 ( .A(n46457), .B(n46445), .Z(n46460) );
  IV U46213 ( .A(n46395), .Z(n46445) );
  XNOR U46214 ( .A(n46461), .B(n46438), .Z(n46395) );
  XNOR U46215 ( .A(n46462), .B(n46444), .Z(n46438) );
  XNOR U46216 ( .A(n46463), .B(n46464), .Z(n46444) );
  NOR U46217 ( .A(n46465), .B(n46466), .Z(n46464) );
  XOR U46218 ( .A(n46463), .B(n46467), .Z(n46465) );
  XNOR U46219 ( .A(n46443), .B(n46435), .Z(n46462) );
  XOR U46220 ( .A(n46468), .B(n46469), .Z(n46435) );
  AND U46221 ( .A(n46470), .B(n46471), .Z(n46469) );
  XOR U46222 ( .A(n46468), .B(n46472), .Z(n46470) );
  XNOR U46223 ( .A(n46473), .B(n46440), .Z(n46443) );
  XOR U46224 ( .A(n46474), .B(n46475), .Z(n46440) );
  AND U46225 ( .A(n46476), .B(n46477), .Z(n46475) );
  XNOR U46226 ( .A(n46478), .B(n46479), .Z(n46476) );
  IV U46227 ( .A(n46474), .Z(n46478) );
  XNOR U46228 ( .A(n46480), .B(n46481), .Z(n46473) );
  NOR U46229 ( .A(n46482), .B(n46483), .Z(n46481) );
  XNOR U46230 ( .A(n46480), .B(n46484), .Z(n46482) );
  XNOR U46231 ( .A(n46439), .B(n46446), .Z(n46461) );
  NOR U46232 ( .A(n46401), .B(n46485), .Z(n46446) );
  XOR U46233 ( .A(n46451), .B(n46450), .Z(n46439) );
  XNOR U46234 ( .A(n46486), .B(n46447), .Z(n46450) );
  XOR U46235 ( .A(n46487), .B(n46488), .Z(n46447) );
  AND U46236 ( .A(n46489), .B(n46490), .Z(n46488) );
  XNOR U46237 ( .A(n46491), .B(n46492), .Z(n46489) );
  IV U46238 ( .A(n46487), .Z(n46491) );
  XNOR U46239 ( .A(n46493), .B(n46494), .Z(n46486) );
  NOR U46240 ( .A(n46495), .B(n46496), .Z(n46494) );
  XNOR U46241 ( .A(n46493), .B(n46497), .Z(n46495) );
  XOR U46242 ( .A(n46498), .B(n46499), .Z(n46451) );
  NOR U46243 ( .A(n46500), .B(n46501), .Z(n46499) );
  XNOR U46244 ( .A(n46498), .B(n46502), .Z(n46500) );
  XNOR U46245 ( .A(n46392), .B(n46457), .Z(n46459) );
  XNOR U46246 ( .A(n46503), .B(n46504), .Z(n46392) );
  AND U46247 ( .A(n1538), .B(n46505), .Z(n46504) );
  XNOR U46248 ( .A(n46506), .B(n46507), .Z(n46505) );
  AND U46249 ( .A(n46398), .B(n46401), .Z(n46457) );
  XOR U46250 ( .A(n46508), .B(n46485), .Z(n46401) );
  XNOR U46251 ( .A(p_input[1232]), .B(p_input[2048]), .Z(n46485) );
  XNOR U46252 ( .A(n46472), .B(n46471), .Z(n46508) );
  XNOR U46253 ( .A(n46509), .B(n46479), .Z(n46471) );
  XNOR U46254 ( .A(n46467), .B(n46466), .Z(n46479) );
  XNOR U46255 ( .A(n46510), .B(n46463), .Z(n46466) );
  XNOR U46256 ( .A(p_input[1242]), .B(p_input[2058]), .Z(n46463) );
  XOR U46257 ( .A(p_input[1243]), .B(n29030), .Z(n46510) );
  XOR U46258 ( .A(p_input[1244]), .B(p_input[2060]), .Z(n46467) );
  XOR U46259 ( .A(n46477), .B(n46511), .Z(n46509) );
  IV U46260 ( .A(n46468), .Z(n46511) );
  XOR U46261 ( .A(p_input[1233]), .B(p_input[2049]), .Z(n46468) );
  XNOR U46262 ( .A(n46512), .B(n46484), .Z(n46477) );
  XNOR U46263 ( .A(p_input[1247]), .B(n29033), .Z(n46484) );
  XOR U46264 ( .A(n46474), .B(n46483), .Z(n46512) );
  XOR U46265 ( .A(n46513), .B(n46480), .Z(n46483) );
  XOR U46266 ( .A(p_input[1245]), .B(p_input[2061]), .Z(n46480) );
  XOR U46267 ( .A(p_input[1246]), .B(n29035), .Z(n46513) );
  XOR U46268 ( .A(p_input[1241]), .B(p_input[2057]), .Z(n46474) );
  XOR U46269 ( .A(n46492), .B(n46490), .Z(n46472) );
  XNOR U46270 ( .A(n46514), .B(n46497), .Z(n46490) );
  XOR U46271 ( .A(p_input[1240]), .B(p_input[2056]), .Z(n46497) );
  XOR U46272 ( .A(n46487), .B(n46496), .Z(n46514) );
  XOR U46273 ( .A(n46515), .B(n46493), .Z(n46496) );
  XOR U46274 ( .A(p_input[1238]), .B(p_input[2054]), .Z(n46493) );
  XOR U46275 ( .A(p_input[1239]), .B(n30404), .Z(n46515) );
  XOR U46276 ( .A(p_input[1234]), .B(p_input[2050]), .Z(n46487) );
  XNOR U46277 ( .A(n46502), .B(n46501), .Z(n46492) );
  XOR U46278 ( .A(n46516), .B(n46498), .Z(n46501) );
  XOR U46279 ( .A(p_input[1235]), .B(p_input[2051]), .Z(n46498) );
  XOR U46280 ( .A(p_input[1236]), .B(n30406), .Z(n46516) );
  XOR U46281 ( .A(p_input[1237]), .B(p_input[2053]), .Z(n46502) );
  XNOR U46282 ( .A(n46517), .B(n46518), .Z(n46398) );
  AND U46283 ( .A(n1538), .B(n46519), .Z(n46518) );
  XNOR U46284 ( .A(n46520), .B(n46521), .Z(n1538) );
  AND U46285 ( .A(n46522), .B(n46523), .Z(n46521) );
  XOR U46286 ( .A(n46412), .B(n46520), .Z(n46523) );
  XNOR U46287 ( .A(n46524), .B(n46520), .Z(n46522) );
  XOR U46288 ( .A(n46525), .B(n46526), .Z(n46520) );
  AND U46289 ( .A(n46527), .B(n46528), .Z(n46526) );
  XOR U46290 ( .A(n46427), .B(n46525), .Z(n46528) );
  XOR U46291 ( .A(n46525), .B(n46428), .Z(n46527) );
  XOR U46292 ( .A(n46529), .B(n46530), .Z(n46525) );
  AND U46293 ( .A(n46531), .B(n46532), .Z(n46530) );
  XOR U46294 ( .A(n46455), .B(n46529), .Z(n46532) );
  XOR U46295 ( .A(n46529), .B(n46456), .Z(n46531) );
  XOR U46296 ( .A(n46533), .B(n46534), .Z(n46529) );
  AND U46297 ( .A(n46535), .B(n46536), .Z(n46534) );
  XOR U46298 ( .A(n46533), .B(n46506), .Z(n46536) );
  XNOR U46299 ( .A(n46537), .B(n46538), .Z(n46358) );
  AND U46300 ( .A(n1542), .B(n46539), .Z(n46538) );
  XNOR U46301 ( .A(n46540), .B(n46541), .Z(n1542) );
  AND U46302 ( .A(n46542), .B(n46543), .Z(n46541) );
  XOR U46303 ( .A(n46540), .B(n46368), .Z(n46543) );
  XNOR U46304 ( .A(n46540), .B(n46328), .Z(n46542) );
  XOR U46305 ( .A(n46544), .B(n46545), .Z(n46540) );
  AND U46306 ( .A(n46546), .B(n46547), .Z(n46545) );
  XOR U46307 ( .A(n46544), .B(n46336), .Z(n46546) );
  XOR U46308 ( .A(n46548), .B(n46549), .Z(n46319) );
  AND U46309 ( .A(n1546), .B(n46539), .Z(n46549) );
  XNOR U46310 ( .A(n46537), .B(n46548), .Z(n46539) );
  XNOR U46311 ( .A(n46550), .B(n46551), .Z(n1546) );
  AND U46312 ( .A(n46552), .B(n46553), .Z(n46551) );
  XNOR U46313 ( .A(n46554), .B(n46550), .Z(n46553) );
  IV U46314 ( .A(n46368), .Z(n46554) );
  XOR U46315 ( .A(n46524), .B(n46555), .Z(n46368) );
  AND U46316 ( .A(n1549), .B(n46556), .Z(n46555) );
  XOR U46317 ( .A(n46411), .B(n46408), .Z(n46556) );
  IV U46318 ( .A(n46524), .Z(n46411) );
  XNOR U46319 ( .A(n46328), .B(n46550), .Z(n46552) );
  XOR U46320 ( .A(n46557), .B(n46558), .Z(n46328) );
  AND U46321 ( .A(n1565), .B(n46559), .Z(n46558) );
  XOR U46322 ( .A(n46544), .B(n46560), .Z(n46550) );
  AND U46323 ( .A(n46561), .B(n46547), .Z(n46560) );
  XNOR U46324 ( .A(n46378), .B(n46544), .Z(n46547) );
  XOR U46325 ( .A(n46428), .B(n46562), .Z(n46378) );
  AND U46326 ( .A(n1549), .B(n46563), .Z(n46562) );
  XOR U46327 ( .A(n46424), .B(n46428), .Z(n46563) );
  XNOR U46328 ( .A(n46564), .B(n46544), .Z(n46561) );
  IV U46329 ( .A(n46336), .Z(n46564) );
  XOR U46330 ( .A(n46565), .B(n46566), .Z(n46336) );
  AND U46331 ( .A(n1565), .B(n46567), .Z(n46566) );
  XOR U46332 ( .A(n46568), .B(n46569), .Z(n46544) );
  AND U46333 ( .A(n46570), .B(n46571), .Z(n46569) );
  XNOR U46334 ( .A(n46388), .B(n46568), .Z(n46571) );
  XOR U46335 ( .A(n46456), .B(n46572), .Z(n46388) );
  AND U46336 ( .A(n1549), .B(n46573), .Z(n46572) );
  XOR U46337 ( .A(n46452), .B(n46456), .Z(n46573) );
  XOR U46338 ( .A(n46568), .B(n46345), .Z(n46570) );
  XOR U46339 ( .A(n46574), .B(n46575), .Z(n46345) );
  AND U46340 ( .A(n1565), .B(n46576), .Z(n46575) );
  XOR U46341 ( .A(n46577), .B(n46578), .Z(n46568) );
  AND U46342 ( .A(n46579), .B(n46580), .Z(n46578) );
  XNOR U46343 ( .A(n46577), .B(n46396), .Z(n46580) );
  XOR U46344 ( .A(n46507), .B(n46581), .Z(n46396) );
  AND U46345 ( .A(n1549), .B(n46582), .Z(n46581) );
  XOR U46346 ( .A(n46503), .B(n46507), .Z(n46582) );
  XNOR U46347 ( .A(n46583), .B(n46577), .Z(n46579) );
  IV U46348 ( .A(n46355), .Z(n46583) );
  XOR U46349 ( .A(n46584), .B(n46585), .Z(n46355) );
  AND U46350 ( .A(n1565), .B(n46586), .Z(n46585) );
  AND U46351 ( .A(n46548), .B(n46537), .Z(n46577) );
  XNOR U46352 ( .A(n46587), .B(n46588), .Z(n46537) );
  AND U46353 ( .A(n1549), .B(n46519), .Z(n46588) );
  XNOR U46354 ( .A(n46517), .B(n46587), .Z(n46519) );
  XNOR U46355 ( .A(n46589), .B(n46590), .Z(n1549) );
  AND U46356 ( .A(n46591), .B(n46592), .Z(n46590) );
  XNOR U46357 ( .A(n46589), .B(n46408), .Z(n46592) );
  IV U46358 ( .A(n46412), .Z(n46408) );
  XOR U46359 ( .A(n46593), .B(n46594), .Z(n46412) );
  AND U46360 ( .A(n1553), .B(n46595), .Z(n46594) );
  XOR U46361 ( .A(n46596), .B(n46593), .Z(n46595) );
  XNOR U46362 ( .A(n46589), .B(n46524), .Z(n46591) );
  XOR U46363 ( .A(n46597), .B(n46598), .Z(n46524) );
  AND U46364 ( .A(n1561), .B(n46559), .Z(n46598) );
  XOR U46365 ( .A(n46557), .B(n46597), .Z(n46559) );
  XOR U46366 ( .A(n46599), .B(n46600), .Z(n46589) );
  AND U46367 ( .A(n46601), .B(n46602), .Z(n46600) );
  XNOR U46368 ( .A(n46599), .B(n46424), .Z(n46602) );
  IV U46369 ( .A(n46427), .Z(n46424) );
  XOR U46370 ( .A(n46603), .B(n46604), .Z(n46427) );
  AND U46371 ( .A(n1553), .B(n46605), .Z(n46604) );
  XOR U46372 ( .A(n46606), .B(n46603), .Z(n46605) );
  XOR U46373 ( .A(n46428), .B(n46599), .Z(n46601) );
  XOR U46374 ( .A(n46607), .B(n46608), .Z(n46428) );
  AND U46375 ( .A(n1561), .B(n46567), .Z(n46608) );
  XOR U46376 ( .A(n46607), .B(n46565), .Z(n46567) );
  XOR U46377 ( .A(n46609), .B(n46610), .Z(n46599) );
  AND U46378 ( .A(n46611), .B(n46612), .Z(n46610) );
  XNOR U46379 ( .A(n46609), .B(n46452), .Z(n46612) );
  IV U46380 ( .A(n46455), .Z(n46452) );
  XOR U46381 ( .A(n46613), .B(n46614), .Z(n46455) );
  AND U46382 ( .A(n1553), .B(n46615), .Z(n46614) );
  XNOR U46383 ( .A(n46616), .B(n46613), .Z(n46615) );
  XOR U46384 ( .A(n46456), .B(n46609), .Z(n46611) );
  XOR U46385 ( .A(n46617), .B(n46618), .Z(n46456) );
  AND U46386 ( .A(n1561), .B(n46576), .Z(n46618) );
  XOR U46387 ( .A(n46617), .B(n46574), .Z(n46576) );
  XOR U46388 ( .A(n46533), .B(n46619), .Z(n46609) );
  AND U46389 ( .A(n46535), .B(n46620), .Z(n46619) );
  XNOR U46390 ( .A(n46533), .B(n46503), .Z(n46620) );
  IV U46391 ( .A(n46506), .Z(n46503) );
  XOR U46392 ( .A(n46621), .B(n46622), .Z(n46506) );
  AND U46393 ( .A(n1553), .B(n46623), .Z(n46622) );
  XOR U46394 ( .A(n46624), .B(n46621), .Z(n46623) );
  XOR U46395 ( .A(n46507), .B(n46533), .Z(n46535) );
  XOR U46396 ( .A(n46625), .B(n46626), .Z(n46507) );
  AND U46397 ( .A(n1561), .B(n46586), .Z(n46626) );
  XOR U46398 ( .A(n46625), .B(n46584), .Z(n46586) );
  AND U46399 ( .A(n46587), .B(n46517), .Z(n46533) );
  XNOR U46400 ( .A(n46627), .B(n46628), .Z(n46517) );
  AND U46401 ( .A(n1553), .B(n46629), .Z(n46628) );
  XNOR U46402 ( .A(n46630), .B(n46627), .Z(n46629) );
  XNOR U46403 ( .A(n46631), .B(n46632), .Z(n1553) );
  AND U46404 ( .A(n46633), .B(n46634), .Z(n46632) );
  XOR U46405 ( .A(n46596), .B(n46631), .Z(n46634) );
  AND U46406 ( .A(n46635), .B(n46636), .Z(n46596) );
  XNOR U46407 ( .A(n46593), .B(n46631), .Z(n46633) );
  XNOR U46408 ( .A(n46637), .B(n46638), .Z(n46593) );
  AND U46409 ( .A(n1557), .B(n46639), .Z(n46638) );
  XNOR U46410 ( .A(n46640), .B(n46641), .Z(n46639) );
  XOR U46411 ( .A(n46642), .B(n46643), .Z(n46631) );
  AND U46412 ( .A(n46644), .B(n46645), .Z(n46643) );
  XNOR U46413 ( .A(n46642), .B(n46635), .Z(n46645) );
  IV U46414 ( .A(n46606), .Z(n46635) );
  XOR U46415 ( .A(n46646), .B(n46647), .Z(n46606) );
  XOR U46416 ( .A(n46648), .B(n46636), .Z(n46647) );
  AND U46417 ( .A(n46616), .B(n46649), .Z(n46636) );
  AND U46418 ( .A(n46650), .B(n46651), .Z(n46648) );
  XOR U46419 ( .A(n46652), .B(n46646), .Z(n46650) );
  XNOR U46420 ( .A(n46603), .B(n46642), .Z(n46644) );
  XNOR U46421 ( .A(n46653), .B(n46654), .Z(n46603) );
  AND U46422 ( .A(n1557), .B(n46655), .Z(n46654) );
  XNOR U46423 ( .A(n46656), .B(n46657), .Z(n46655) );
  XOR U46424 ( .A(n46658), .B(n46659), .Z(n46642) );
  AND U46425 ( .A(n46660), .B(n46661), .Z(n46659) );
  XNOR U46426 ( .A(n46658), .B(n46616), .Z(n46661) );
  XOR U46427 ( .A(n46662), .B(n46651), .Z(n46616) );
  XNOR U46428 ( .A(n46663), .B(n46646), .Z(n46651) );
  XOR U46429 ( .A(n46664), .B(n46665), .Z(n46646) );
  AND U46430 ( .A(n46666), .B(n46667), .Z(n46665) );
  XOR U46431 ( .A(n46668), .B(n46664), .Z(n46666) );
  XNOR U46432 ( .A(n46669), .B(n46670), .Z(n46663) );
  AND U46433 ( .A(n46671), .B(n46672), .Z(n46670) );
  XOR U46434 ( .A(n46669), .B(n46673), .Z(n46671) );
  XNOR U46435 ( .A(n46652), .B(n46649), .Z(n46662) );
  AND U46436 ( .A(n46674), .B(n46675), .Z(n46649) );
  XOR U46437 ( .A(n46676), .B(n46677), .Z(n46652) );
  AND U46438 ( .A(n46678), .B(n46679), .Z(n46677) );
  XOR U46439 ( .A(n46676), .B(n46680), .Z(n46678) );
  XNOR U46440 ( .A(n46613), .B(n46658), .Z(n46660) );
  XNOR U46441 ( .A(n46681), .B(n46682), .Z(n46613) );
  AND U46442 ( .A(n1557), .B(n46683), .Z(n46682) );
  XNOR U46443 ( .A(n46684), .B(n46685), .Z(n46683) );
  XOR U46444 ( .A(n46686), .B(n46687), .Z(n46658) );
  AND U46445 ( .A(n46688), .B(n46689), .Z(n46687) );
  XNOR U46446 ( .A(n46686), .B(n46674), .Z(n46689) );
  IV U46447 ( .A(n46624), .Z(n46674) );
  XNOR U46448 ( .A(n46690), .B(n46667), .Z(n46624) );
  XNOR U46449 ( .A(n46691), .B(n46673), .Z(n46667) );
  XNOR U46450 ( .A(n46692), .B(n46693), .Z(n46673) );
  NOR U46451 ( .A(n46694), .B(n46695), .Z(n46693) );
  XOR U46452 ( .A(n46692), .B(n46696), .Z(n46694) );
  XNOR U46453 ( .A(n46672), .B(n46664), .Z(n46691) );
  XOR U46454 ( .A(n46697), .B(n46698), .Z(n46664) );
  AND U46455 ( .A(n46699), .B(n46700), .Z(n46698) );
  XOR U46456 ( .A(n46697), .B(n46701), .Z(n46699) );
  XNOR U46457 ( .A(n46702), .B(n46669), .Z(n46672) );
  XOR U46458 ( .A(n46703), .B(n46704), .Z(n46669) );
  AND U46459 ( .A(n46705), .B(n46706), .Z(n46704) );
  XNOR U46460 ( .A(n46707), .B(n46708), .Z(n46705) );
  IV U46461 ( .A(n46703), .Z(n46707) );
  XNOR U46462 ( .A(n46709), .B(n46710), .Z(n46702) );
  NOR U46463 ( .A(n46711), .B(n46712), .Z(n46710) );
  XNOR U46464 ( .A(n46709), .B(n46713), .Z(n46711) );
  XNOR U46465 ( .A(n46668), .B(n46675), .Z(n46690) );
  NOR U46466 ( .A(n46630), .B(n46714), .Z(n46675) );
  XOR U46467 ( .A(n46680), .B(n46679), .Z(n46668) );
  XNOR U46468 ( .A(n46715), .B(n46676), .Z(n46679) );
  XOR U46469 ( .A(n46716), .B(n46717), .Z(n46676) );
  AND U46470 ( .A(n46718), .B(n46719), .Z(n46717) );
  XNOR U46471 ( .A(n46720), .B(n46721), .Z(n46718) );
  IV U46472 ( .A(n46716), .Z(n46720) );
  XNOR U46473 ( .A(n46722), .B(n46723), .Z(n46715) );
  NOR U46474 ( .A(n46724), .B(n46725), .Z(n46723) );
  XNOR U46475 ( .A(n46722), .B(n46726), .Z(n46724) );
  XOR U46476 ( .A(n46727), .B(n46728), .Z(n46680) );
  NOR U46477 ( .A(n46729), .B(n46730), .Z(n46728) );
  XNOR U46478 ( .A(n46727), .B(n46731), .Z(n46729) );
  XNOR U46479 ( .A(n46621), .B(n46686), .Z(n46688) );
  XNOR U46480 ( .A(n46732), .B(n46733), .Z(n46621) );
  AND U46481 ( .A(n1557), .B(n46734), .Z(n46733) );
  XNOR U46482 ( .A(n46735), .B(n46736), .Z(n46734) );
  AND U46483 ( .A(n46627), .B(n46630), .Z(n46686) );
  XOR U46484 ( .A(n46737), .B(n46714), .Z(n46630) );
  XNOR U46485 ( .A(p_input[1248]), .B(p_input[2048]), .Z(n46714) );
  XNOR U46486 ( .A(n46701), .B(n46700), .Z(n46737) );
  XNOR U46487 ( .A(n46738), .B(n46708), .Z(n46700) );
  XNOR U46488 ( .A(n46696), .B(n46695), .Z(n46708) );
  XNOR U46489 ( .A(n46739), .B(n46692), .Z(n46695) );
  XNOR U46490 ( .A(p_input[1258]), .B(p_input[2058]), .Z(n46692) );
  XOR U46491 ( .A(p_input[1259]), .B(n29030), .Z(n46739) );
  XOR U46492 ( .A(p_input[1260]), .B(p_input[2060]), .Z(n46696) );
  XOR U46493 ( .A(n46706), .B(n46740), .Z(n46738) );
  IV U46494 ( .A(n46697), .Z(n46740) );
  XOR U46495 ( .A(p_input[1249]), .B(p_input[2049]), .Z(n46697) );
  XNOR U46496 ( .A(n46741), .B(n46713), .Z(n46706) );
  XNOR U46497 ( .A(p_input[1263]), .B(n29033), .Z(n46713) );
  XOR U46498 ( .A(n46703), .B(n46712), .Z(n46741) );
  XOR U46499 ( .A(n46742), .B(n46709), .Z(n46712) );
  XOR U46500 ( .A(p_input[1261]), .B(p_input[2061]), .Z(n46709) );
  XOR U46501 ( .A(p_input[1262]), .B(n29035), .Z(n46742) );
  XOR U46502 ( .A(p_input[1257]), .B(p_input[2057]), .Z(n46703) );
  XOR U46503 ( .A(n46721), .B(n46719), .Z(n46701) );
  XNOR U46504 ( .A(n46743), .B(n46726), .Z(n46719) );
  XOR U46505 ( .A(p_input[1256]), .B(p_input[2056]), .Z(n46726) );
  XOR U46506 ( .A(n46716), .B(n46725), .Z(n46743) );
  XOR U46507 ( .A(n46744), .B(n46722), .Z(n46725) );
  XOR U46508 ( .A(p_input[1254]), .B(p_input[2054]), .Z(n46722) );
  XOR U46509 ( .A(p_input[1255]), .B(n30404), .Z(n46744) );
  XOR U46510 ( .A(p_input[1250]), .B(p_input[2050]), .Z(n46716) );
  XNOR U46511 ( .A(n46731), .B(n46730), .Z(n46721) );
  XOR U46512 ( .A(n46745), .B(n46727), .Z(n46730) );
  XOR U46513 ( .A(p_input[1251]), .B(p_input[2051]), .Z(n46727) );
  XOR U46514 ( .A(p_input[1252]), .B(n30406), .Z(n46745) );
  XOR U46515 ( .A(p_input[1253]), .B(p_input[2053]), .Z(n46731) );
  XNOR U46516 ( .A(n46746), .B(n46747), .Z(n46627) );
  AND U46517 ( .A(n1557), .B(n46748), .Z(n46747) );
  XNOR U46518 ( .A(n46749), .B(n46750), .Z(n1557) );
  AND U46519 ( .A(n46751), .B(n46752), .Z(n46750) );
  XOR U46520 ( .A(n46641), .B(n46749), .Z(n46752) );
  XNOR U46521 ( .A(n46753), .B(n46749), .Z(n46751) );
  XOR U46522 ( .A(n46754), .B(n46755), .Z(n46749) );
  AND U46523 ( .A(n46756), .B(n46757), .Z(n46755) );
  XOR U46524 ( .A(n46656), .B(n46754), .Z(n46757) );
  XOR U46525 ( .A(n46754), .B(n46657), .Z(n46756) );
  XOR U46526 ( .A(n46758), .B(n46759), .Z(n46754) );
  AND U46527 ( .A(n46760), .B(n46761), .Z(n46759) );
  XOR U46528 ( .A(n46684), .B(n46758), .Z(n46761) );
  XOR U46529 ( .A(n46758), .B(n46685), .Z(n46760) );
  XOR U46530 ( .A(n46762), .B(n46763), .Z(n46758) );
  AND U46531 ( .A(n46764), .B(n46765), .Z(n46763) );
  XOR U46532 ( .A(n46762), .B(n46735), .Z(n46765) );
  XNOR U46533 ( .A(n46766), .B(n46767), .Z(n46587) );
  AND U46534 ( .A(n1561), .B(n46768), .Z(n46767) );
  XNOR U46535 ( .A(n46769), .B(n46770), .Z(n1561) );
  AND U46536 ( .A(n46771), .B(n46772), .Z(n46770) );
  XOR U46537 ( .A(n46769), .B(n46597), .Z(n46772) );
  XNOR U46538 ( .A(n46769), .B(n46557), .Z(n46771) );
  XOR U46539 ( .A(n46773), .B(n46774), .Z(n46769) );
  AND U46540 ( .A(n46775), .B(n46776), .Z(n46774) );
  XOR U46541 ( .A(n46773), .B(n46565), .Z(n46775) );
  XOR U46542 ( .A(n46777), .B(n46778), .Z(n46548) );
  AND U46543 ( .A(n1565), .B(n46768), .Z(n46778) );
  XNOR U46544 ( .A(n46766), .B(n46777), .Z(n46768) );
  XNOR U46545 ( .A(n46779), .B(n46780), .Z(n1565) );
  AND U46546 ( .A(n46781), .B(n46782), .Z(n46780) );
  XNOR U46547 ( .A(n46783), .B(n46779), .Z(n46782) );
  IV U46548 ( .A(n46597), .Z(n46783) );
  XOR U46549 ( .A(n46753), .B(n46784), .Z(n46597) );
  AND U46550 ( .A(n1568), .B(n46785), .Z(n46784) );
  XOR U46551 ( .A(n46640), .B(n46637), .Z(n46785) );
  IV U46552 ( .A(n46753), .Z(n46640) );
  XNOR U46553 ( .A(n46557), .B(n46779), .Z(n46781) );
  XOR U46554 ( .A(n46786), .B(n46787), .Z(n46557) );
  AND U46555 ( .A(n1584), .B(n46788), .Z(n46787) );
  XOR U46556 ( .A(n46773), .B(n46789), .Z(n46779) );
  AND U46557 ( .A(n46790), .B(n46776), .Z(n46789) );
  XNOR U46558 ( .A(n46607), .B(n46773), .Z(n46776) );
  XOR U46559 ( .A(n46657), .B(n46791), .Z(n46607) );
  AND U46560 ( .A(n1568), .B(n46792), .Z(n46791) );
  XOR U46561 ( .A(n46653), .B(n46657), .Z(n46792) );
  XNOR U46562 ( .A(n46793), .B(n46773), .Z(n46790) );
  IV U46563 ( .A(n46565), .Z(n46793) );
  XOR U46564 ( .A(n46794), .B(n46795), .Z(n46565) );
  AND U46565 ( .A(n1584), .B(n46796), .Z(n46795) );
  XOR U46566 ( .A(n46797), .B(n46798), .Z(n46773) );
  AND U46567 ( .A(n46799), .B(n46800), .Z(n46798) );
  XNOR U46568 ( .A(n46617), .B(n46797), .Z(n46800) );
  XOR U46569 ( .A(n46685), .B(n46801), .Z(n46617) );
  AND U46570 ( .A(n1568), .B(n46802), .Z(n46801) );
  XOR U46571 ( .A(n46681), .B(n46685), .Z(n46802) );
  XOR U46572 ( .A(n46797), .B(n46574), .Z(n46799) );
  XOR U46573 ( .A(n46803), .B(n46804), .Z(n46574) );
  AND U46574 ( .A(n1584), .B(n46805), .Z(n46804) );
  XOR U46575 ( .A(n46806), .B(n46807), .Z(n46797) );
  AND U46576 ( .A(n46808), .B(n46809), .Z(n46807) );
  XNOR U46577 ( .A(n46806), .B(n46625), .Z(n46809) );
  XOR U46578 ( .A(n46736), .B(n46810), .Z(n46625) );
  AND U46579 ( .A(n1568), .B(n46811), .Z(n46810) );
  XOR U46580 ( .A(n46732), .B(n46736), .Z(n46811) );
  XNOR U46581 ( .A(n46812), .B(n46806), .Z(n46808) );
  IV U46582 ( .A(n46584), .Z(n46812) );
  XOR U46583 ( .A(n46813), .B(n46814), .Z(n46584) );
  AND U46584 ( .A(n1584), .B(n46815), .Z(n46814) );
  AND U46585 ( .A(n46777), .B(n46766), .Z(n46806) );
  XNOR U46586 ( .A(n46816), .B(n46817), .Z(n46766) );
  AND U46587 ( .A(n1568), .B(n46748), .Z(n46817) );
  XNOR U46588 ( .A(n46746), .B(n46816), .Z(n46748) );
  XNOR U46589 ( .A(n46818), .B(n46819), .Z(n1568) );
  AND U46590 ( .A(n46820), .B(n46821), .Z(n46819) );
  XNOR U46591 ( .A(n46818), .B(n46637), .Z(n46821) );
  IV U46592 ( .A(n46641), .Z(n46637) );
  XOR U46593 ( .A(n46822), .B(n46823), .Z(n46641) );
  AND U46594 ( .A(n1572), .B(n46824), .Z(n46823) );
  XOR U46595 ( .A(n46825), .B(n46822), .Z(n46824) );
  XNOR U46596 ( .A(n46818), .B(n46753), .Z(n46820) );
  XOR U46597 ( .A(n46826), .B(n46827), .Z(n46753) );
  AND U46598 ( .A(n1580), .B(n46788), .Z(n46827) );
  XOR U46599 ( .A(n46786), .B(n46826), .Z(n46788) );
  XOR U46600 ( .A(n46828), .B(n46829), .Z(n46818) );
  AND U46601 ( .A(n46830), .B(n46831), .Z(n46829) );
  XNOR U46602 ( .A(n46828), .B(n46653), .Z(n46831) );
  IV U46603 ( .A(n46656), .Z(n46653) );
  XOR U46604 ( .A(n46832), .B(n46833), .Z(n46656) );
  AND U46605 ( .A(n1572), .B(n46834), .Z(n46833) );
  XOR U46606 ( .A(n46835), .B(n46832), .Z(n46834) );
  XOR U46607 ( .A(n46657), .B(n46828), .Z(n46830) );
  XOR U46608 ( .A(n46836), .B(n46837), .Z(n46657) );
  AND U46609 ( .A(n1580), .B(n46796), .Z(n46837) );
  XOR U46610 ( .A(n46836), .B(n46794), .Z(n46796) );
  XOR U46611 ( .A(n46838), .B(n46839), .Z(n46828) );
  AND U46612 ( .A(n46840), .B(n46841), .Z(n46839) );
  XNOR U46613 ( .A(n46838), .B(n46681), .Z(n46841) );
  IV U46614 ( .A(n46684), .Z(n46681) );
  XOR U46615 ( .A(n46842), .B(n46843), .Z(n46684) );
  AND U46616 ( .A(n1572), .B(n46844), .Z(n46843) );
  XNOR U46617 ( .A(n46845), .B(n46842), .Z(n46844) );
  XOR U46618 ( .A(n46685), .B(n46838), .Z(n46840) );
  XOR U46619 ( .A(n46846), .B(n46847), .Z(n46685) );
  AND U46620 ( .A(n1580), .B(n46805), .Z(n46847) );
  XOR U46621 ( .A(n46846), .B(n46803), .Z(n46805) );
  XOR U46622 ( .A(n46762), .B(n46848), .Z(n46838) );
  AND U46623 ( .A(n46764), .B(n46849), .Z(n46848) );
  XNOR U46624 ( .A(n46762), .B(n46732), .Z(n46849) );
  IV U46625 ( .A(n46735), .Z(n46732) );
  XOR U46626 ( .A(n46850), .B(n46851), .Z(n46735) );
  AND U46627 ( .A(n1572), .B(n46852), .Z(n46851) );
  XOR U46628 ( .A(n46853), .B(n46850), .Z(n46852) );
  XOR U46629 ( .A(n46736), .B(n46762), .Z(n46764) );
  XOR U46630 ( .A(n46854), .B(n46855), .Z(n46736) );
  AND U46631 ( .A(n1580), .B(n46815), .Z(n46855) );
  XOR U46632 ( .A(n46854), .B(n46813), .Z(n46815) );
  AND U46633 ( .A(n46816), .B(n46746), .Z(n46762) );
  XNOR U46634 ( .A(n46856), .B(n46857), .Z(n46746) );
  AND U46635 ( .A(n1572), .B(n46858), .Z(n46857) );
  XNOR U46636 ( .A(n46859), .B(n46856), .Z(n46858) );
  XNOR U46637 ( .A(n46860), .B(n46861), .Z(n1572) );
  AND U46638 ( .A(n46862), .B(n46863), .Z(n46861) );
  XOR U46639 ( .A(n46825), .B(n46860), .Z(n46863) );
  AND U46640 ( .A(n46864), .B(n46865), .Z(n46825) );
  XNOR U46641 ( .A(n46822), .B(n46860), .Z(n46862) );
  XNOR U46642 ( .A(n46866), .B(n46867), .Z(n46822) );
  AND U46643 ( .A(n1576), .B(n46868), .Z(n46867) );
  XNOR U46644 ( .A(n46869), .B(n46870), .Z(n46868) );
  XOR U46645 ( .A(n46871), .B(n46872), .Z(n46860) );
  AND U46646 ( .A(n46873), .B(n46874), .Z(n46872) );
  XNOR U46647 ( .A(n46871), .B(n46864), .Z(n46874) );
  IV U46648 ( .A(n46835), .Z(n46864) );
  XOR U46649 ( .A(n46875), .B(n46876), .Z(n46835) );
  XOR U46650 ( .A(n46877), .B(n46865), .Z(n46876) );
  AND U46651 ( .A(n46845), .B(n46878), .Z(n46865) );
  AND U46652 ( .A(n46879), .B(n46880), .Z(n46877) );
  XOR U46653 ( .A(n46881), .B(n46875), .Z(n46879) );
  XNOR U46654 ( .A(n46832), .B(n46871), .Z(n46873) );
  XNOR U46655 ( .A(n46882), .B(n46883), .Z(n46832) );
  AND U46656 ( .A(n1576), .B(n46884), .Z(n46883) );
  XNOR U46657 ( .A(n46885), .B(n46886), .Z(n46884) );
  XOR U46658 ( .A(n46887), .B(n46888), .Z(n46871) );
  AND U46659 ( .A(n46889), .B(n46890), .Z(n46888) );
  XNOR U46660 ( .A(n46887), .B(n46845), .Z(n46890) );
  XOR U46661 ( .A(n46891), .B(n46880), .Z(n46845) );
  XNOR U46662 ( .A(n46892), .B(n46875), .Z(n46880) );
  XOR U46663 ( .A(n46893), .B(n46894), .Z(n46875) );
  AND U46664 ( .A(n46895), .B(n46896), .Z(n46894) );
  XOR U46665 ( .A(n46897), .B(n46893), .Z(n46895) );
  XNOR U46666 ( .A(n46898), .B(n46899), .Z(n46892) );
  AND U46667 ( .A(n46900), .B(n46901), .Z(n46899) );
  XOR U46668 ( .A(n46898), .B(n46902), .Z(n46900) );
  XNOR U46669 ( .A(n46881), .B(n46878), .Z(n46891) );
  AND U46670 ( .A(n46903), .B(n46904), .Z(n46878) );
  XOR U46671 ( .A(n46905), .B(n46906), .Z(n46881) );
  AND U46672 ( .A(n46907), .B(n46908), .Z(n46906) );
  XOR U46673 ( .A(n46905), .B(n46909), .Z(n46907) );
  XNOR U46674 ( .A(n46842), .B(n46887), .Z(n46889) );
  XNOR U46675 ( .A(n46910), .B(n46911), .Z(n46842) );
  AND U46676 ( .A(n1576), .B(n46912), .Z(n46911) );
  XNOR U46677 ( .A(n46913), .B(n46914), .Z(n46912) );
  XOR U46678 ( .A(n46915), .B(n46916), .Z(n46887) );
  AND U46679 ( .A(n46917), .B(n46918), .Z(n46916) );
  XNOR U46680 ( .A(n46915), .B(n46903), .Z(n46918) );
  IV U46681 ( .A(n46853), .Z(n46903) );
  XNOR U46682 ( .A(n46919), .B(n46896), .Z(n46853) );
  XNOR U46683 ( .A(n46920), .B(n46902), .Z(n46896) );
  XNOR U46684 ( .A(n46921), .B(n46922), .Z(n46902) );
  NOR U46685 ( .A(n46923), .B(n46924), .Z(n46922) );
  XOR U46686 ( .A(n46921), .B(n46925), .Z(n46923) );
  XNOR U46687 ( .A(n46901), .B(n46893), .Z(n46920) );
  XOR U46688 ( .A(n46926), .B(n46927), .Z(n46893) );
  AND U46689 ( .A(n46928), .B(n46929), .Z(n46927) );
  XOR U46690 ( .A(n46926), .B(n46930), .Z(n46928) );
  XNOR U46691 ( .A(n46931), .B(n46898), .Z(n46901) );
  XOR U46692 ( .A(n46932), .B(n46933), .Z(n46898) );
  AND U46693 ( .A(n46934), .B(n46935), .Z(n46933) );
  XNOR U46694 ( .A(n46936), .B(n46937), .Z(n46934) );
  IV U46695 ( .A(n46932), .Z(n46936) );
  XNOR U46696 ( .A(n46938), .B(n46939), .Z(n46931) );
  NOR U46697 ( .A(n46940), .B(n46941), .Z(n46939) );
  XNOR U46698 ( .A(n46938), .B(n46942), .Z(n46940) );
  XNOR U46699 ( .A(n46897), .B(n46904), .Z(n46919) );
  NOR U46700 ( .A(n46859), .B(n46943), .Z(n46904) );
  XOR U46701 ( .A(n46909), .B(n46908), .Z(n46897) );
  XNOR U46702 ( .A(n46944), .B(n46905), .Z(n46908) );
  XOR U46703 ( .A(n46945), .B(n46946), .Z(n46905) );
  AND U46704 ( .A(n46947), .B(n46948), .Z(n46946) );
  XNOR U46705 ( .A(n46949), .B(n46950), .Z(n46947) );
  IV U46706 ( .A(n46945), .Z(n46949) );
  XNOR U46707 ( .A(n46951), .B(n46952), .Z(n46944) );
  NOR U46708 ( .A(n46953), .B(n46954), .Z(n46952) );
  XNOR U46709 ( .A(n46951), .B(n46955), .Z(n46953) );
  XOR U46710 ( .A(n46956), .B(n46957), .Z(n46909) );
  NOR U46711 ( .A(n46958), .B(n46959), .Z(n46957) );
  XNOR U46712 ( .A(n46956), .B(n46960), .Z(n46958) );
  XNOR U46713 ( .A(n46850), .B(n46915), .Z(n46917) );
  XNOR U46714 ( .A(n46961), .B(n46962), .Z(n46850) );
  AND U46715 ( .A(n1576), .B(n46963), .Z(n46962) );
  XNOR U46716 ( .A(n46964), .B(n46965), .Z(n46963) );
  AND U46717 ( .A(n46856), .B(n46859), .Z(n46915) );
  XOR U46718 ( .A(n46966), .B(n46943), .Z(n46859) );
  XNOR U46719 ( .A(p_input[1264]), .B(p_input[2048]), .Z(n46943) );
  XNOR U46720 ( .A(n46930), .B(n46929), .Z(n46966) );
  XNOR U46721 ( .A(n46967), .B(n46937), .Z(n46929) );
  XNOR U46722 ( .A(n46925), .B(n46924), .Z(n46937) );
  XNOR U46723 ( .A(n46968), .B(n46921), .Z(n46924) );
  XNOR U46724 ( .A(p_input[1274]), .B(p_input[2058]), .Z(n46921) );
  XOR U46725 ( .A(p_input[1275]), .B(n29030), .Z(n46968) );
  XOR U46726 ( .A(p_input[1276]), .B(p_input[2060]), .Z(n46925) );
  XOR U46727 ( .A(n46935), .B(n46969), .Z(n46967) );
  IV U46728 ( .A(n46926), .Z(n46969) );
  XOR U46729 ( .A(p_input[1265]), .B(p_input[2049]), .Z(n46926) );
  XNOR U46730 ( .A(n46970), .B(n46942), .Z(n46935) );
  XNOR U46731 ( .A(p_input[1279]), .B(n29033), .Z(n46942) );
  XOR U46732 ( .A(n46932), .B(n46941), .Z(n46970) );
  XOR U46733 ( .A(n46971), .B(n46938), .Z(n46941) );
  XOR U46734 ( .A(p_input[1277]), .B(p_input[2061]), .Z(n46938) );
  XOR U46735 ( .A(p_input[1278]), .B(n29035), .Z(n46971) );
  XOR U46736 ( .A(p_input[1273]), .B(p_input[2057]), .Z(n46932) );
  XOR U46737 ( .A(n46950), .B(n46948), .Z(n46930) );
  XNOR U46738 ( .A(n46972), .B(n46955), .Z(n46948) );
  XOR U46739 ( .A(p_input[1272]), .B(p_input[2056]), .Z(n46955) );
  XOR U46740 ( .A(n46945), .B(n46954), .Z(n46972) );
  XOR U46741 ( .A(n46973), .B(n46951), .Z(n46954) );
  XOR U46742 ( .A(p_input[1270]), .B(p_input[2054]), .Z(n46951) );
  XOR U46743 ( .A(p_input[1271]), .B(n30404), .Z(n46973) );
  XOR U46744 ( .A(p_input[1266]), .B(p_input[2050]), .Z(n46945) );
  XNOR U46745 ( .A(n46960), .B(n46959), .Z(n46950) );
  XOR U46746 ( .A(n46974), .B(n46956), .Z(n46959) );
  XOR U46747 ( .A(p_input[1267]), .B(p_input[2051]), .Z(n46956) );
  XOR U46748 ( .A(p_input[1268]), .B(n30406), .Z(n46974) );
  XOR U46749 ( .A(p_input[1269]), .B(p_input[2053]), .Z(n46960) );
  XNOR U46750 ( .A(n46975), .B(n46976), .Z(n46856) );
  AND U46751 ( .A(n1576), .B(n46977), .Z(n46976) );
  XNOR U46752 ( .A(n46978), .B(n46979), .Z(n1576) );
  AND U46753 ( .A(n46980), .B(n46981), .Z(n46979) );
  XOR U46754 ( .A(n46870), .B(n46978), .Z(n46981) );
  XNOR U46755 ( .A(n46982), .B(n46978), .Z(n46980) );
  XOR U46756 ( .A(n46983), .B(n46984), .Z(n46978) );
  AND U46757 ( .A(n46985), .B(n46986), .Z(n46984) );
  XOR U46758 ( .A(n46885), .B(n46983), .Z(n46986) );
  XOR U46759 ( .A(n46983), .B(n46886), .Z(n46985) );
  XOR U46760 ( .A(n46987), .B(n46988), .Z(n46983) );
  AND U46761 ( .A(n46989), .B(n46990), .Z(n46988) );
  XOR U46762 ( .A(n46913), .B(n46987), .Z(n46990) );
  XOR U46763 ( .A(n46987), .B(n46914), .Z(n46989) );
  XOR U46764 ( .A(n46991), .B(n46992), .Z(n46987) );
  AND U46765 ( .A(n46993), .B(n46994), .Z(n46992) );
  XOR U46766 ( .A(n46991), .B(n46964), .Z(n46994) );
  XNOR U46767 ( .A(n46995), .B(n46996), .Z(n46816) );
  AND U46768 ( .A(n1580), .B(n46997), .Z(n46996) );
  XNOR U46769 ( .A(n46998), .B(n46999), .Z(n1580) );
  AND U46770 ( .A(n47000), .B(n47001), .Z(n46999) );
  XOR U46771 ( .A(n46998), .B(n46826), .Z(n47001) );
  XNOR U46772 ( .A(n46998), .B(n46786), .Z(n47000) );
  XOR U46773 ( .A(n47002), .B(n47003), .Z(n46998) );
  AND U46774 ( .A(n47004), .B(n47005), .Z(n47003) );
  XOR U46775 ( .A(n47002), .B(n46794), .Z(n47004) );
  XOR U46776 ( .A(n47006), .B(n47007), .Z(n46777) );
  AND U46777 ( .A(n1584), .B(n46997), .Z(n47007) );
  XNOR U46778 ( .A(n46995), .B(n47006), .Z(n46997) );
  XNOR U46779 ( .A(n47008), .B(n47009), .Z(n1584) );
  AND U46780 ( .A(n47010), .B(n47011), .Z(n47009) );
  XNOR U46781 ( .A(n47012), .B(n47008), .Z(n47011) );
  IV U46782 ( .A(n46826), .Z(n47012) );
  XOR U46783 ( .A(n46982), .B(n47013), .Z(n46826) );
  AND U46784 ( .A(n1587), .B(n47014), .Z(n47013) );
  XOR U46785 ( .A(n46869), .B(n46866), .Z(n47014) );
  IV U46786 ( .A(n46982), .Z(n46869) );
  XNOR U46787 ( .A(n46786), .B(n47008), .Z(n47010) );
  XOR U46788 ( .A(n47015), .B(n47016), .Z(n46786) );
  AND U46789 ( .A(n1603), .B(n47017), .Z(n47016) );
  XOR U46790 ( .A(n47002), .B(n47018), .Z(n47008) );
  AND U46791 ( .A(n47019), .B(n47005), .Z(n47018) );
  XNOR U46792 ( .A(n46836), .B(n47002), .Z(n47005) );
  XOR U46793 ( .A(n46886), .B(n47020), .Z(n46836) );
  AND U46794 ( .A(n1587), .B(n47021), .Z(n47020) );
  XOR U46795 ( .A(n46882), .B(n46886), .Z(n47021) );
  XNOR U46796 ( .A(n47022), .B(n47002), .Z(n47019) );
  IV U46797 ( .A(n46794), .Z(n47022) );
  XOR U46798 ( .A(n47023), .B(n47024), .Z(n46794) );
  AND U46799 ( .A(n1603), .B(n47025), .Z(n47024) );
  XOR U46800 ( .A(n47026), .B(n47027), .Z(n47002) );
  AND U46801 ( .A(n47028), .B(n47029), .Z(n47027) );
  XNOR U46802 ( .A(n46846), .B(n47026), .Z(n47029) );
  XOR U46803 ( .A(n46914), .B(n47030), .Z(n46846) );
  AND U46804 ( .A(n1587), .B(n47031), .Z(n47030) );
  XOR U46805 ( .A(n46910), .B(n46914), .Z(n47031) );
  XOR U46806 ( .A(n47026), .B(n46803), .Z(n47028) );
  XOR U46807 ( .A(n47032), .B(n47033), .Z(n46803) );
  AND U46808 ( .A(n1603), .B(n47034), .Z(n47033) );
  XOR U46809 ( .A(n47035), .B(n47036), .Z(n47026) );
  AND U46810 ( .A(n47037), .B(n47038), .Z(n47036) );
  XNOR U46811 ( .A(n47035), .B(n46854), .Z(n47038) );
  XOR U46812 ( .A(n46965), .B(n47039), .Z(n46854) );
  AND U46813 ( .A(n1587), .B(n47040), .Z(n47039) );
  XOR U46814 ( .A(n46961), .B(n46965), .Z(n47040) );
  XNOR U46815 ( .A(n47041), .B(n47035), .Z(n47037) );
  IV U46816 ( .A(n46813), .Z(n47041) );
  XOR U46817 ( .A(n47042), .B(n47043), .Z(n46813) );
  AND U46818 ( .A(n1603), .B(n47044), .Z(n47043) );
  AND U46819 ( .A(n47006), .B(n46995), .Z(n47035) );
  XNOR U46820 ( .A(n47045), .B(n47046), .Z(n46995) );
  AND U46821 ( .A(n1587), .B(n46977), .Z(n47046) );
  XNOR U46822 ( .A(n46975), .B(n47045), .Z(n46977) );
  XNOR U46823 ( .A(n47047), .B(n47048), .Z(n1587) );
  AND U46824 ( .A(n47049), .B(n47050), .Z(n47048) );
  XNOR U46825 ( .A(n47047), .B(n46866), .Z(n47050) );
  IV U46826 ( .A(n46870), .Z(n46866) );
  XOR U46827 ( .A(n47051), .B(n47052), .Z(n46870) );
  AND U46828 ( .A(n1591), .B(n47053), .Z(n47052) );
  XOR U46829 ( .A(n47054), .B(n47051), .Z(n47053) );
  XNOR U46830 ( .A(n47047), .B(n46982), .Z(n47049) );
  XOR U46831 ( .A(n47055), .B(n47056), .Z(n46982) );
  AND U46832 ( .A(n1599), .B(n47017), .Z(n47056) );
  XOR U46833 ( .A(n47015), .B(n47055), .Z(n47017) );
  XOR U46834 ( .A(n47057), .B(n47058), .Z(n47047) );
  AND U46835 ( .A(n47059), .B(n47060), .Z(n47058) );
  XNOR U46836 ( .A(n47057), .B(n46882), .Z(n47060) );
  IV U46837 ( .A(n46885), .Z(n46882) );
  XOR U46838 ( .A(n47061), .B(n47062), .Z(n46885) );
  AND U46839 ( .A(n1591), .B(n47063), .Z(n47062) );
  XOR U46840 ( .A(n47064), .B(n47061), .Z(n47063) );
  XOR U46841 ( .A(n46886), .B(n47057), .Z(n47059) );
  XOR U46842 ( .A(n47065), .B(n47066), .Z(n46886) );
  AND U46843 ( .A(n1599), .B(n47025), .Z(n47066) );
  XOR U46844 ( .A(n47065), .B(n47023), .Z(n47025) );
  XOR U46845 ( .A(n47067), .B(n47068), .Z(n47057) );
  AND U46846 ( .A(n47069), .B(n47070), .Z(n47068) );
  XNOR U46847 ( .A(n47067), .B(n46910), .Z(n47070) );
  IV U46848 ( .A(n46913), .Z(n46910) );
  XOR U46849 ( .A(n47071), .B(n47072), .Z(n46913) );
  AND U46850 ( .A(n1591), .B(n47073), .Z(n47072) );
  XNOR U46851 ( .A(n47074), .B(n47071), .Z(n47073) );
  XOR U46852 ( .A(n46914), .B(n47067), .Z(n47069) );
  XOR U46853 ( .A(n47075), .B(n47076), .Z(n46914) );
  AND U46854 ( .A(n1599), .B(n47034), .Z(n47076) );
  XOR U46855 ( .A(n47075), .B(n47032), .Z(n47034) );
  XOR U46856 ( .A(n46991), .B(n47077), .Z(n47067) );
  AND U46857 ( .A(n46993), .B(n47078), .Z(n47077) );
  XNOR U46858 ( .A(n46991), .B(n46961), .Z(n47078) );
  IV U46859 ( .A(n46964), .Z(n46961) );
  XOR U46860 ( .A(n47079), .B(n47080), .Z(n46964) );
  AND U46861 ( .A(n1591), .B(n47081), .Z(n47080) );
  XOR U46862 ( .A(n47082), .B(n47079), .Z(n47081) );
  XOR U46863 ( .A(n46965), .B(n46991), .Z(n46993) );
  XOR U46864 ( .A(n47083), .B(n47084), .Z(n46965) );
  AND U46865 ( .A(n1599), .B(n47044), .Z(n47084) );
  XOR U46866 ( .A(n47083), .B(n47042), .Z(n47044) );
  AND U46867 ( .A(n47045), .B(n46975), .Z(n46991) );
  XNOR U46868 ( .A(n47085), .B(n47086), .Z(n46975) );
  AND U46869 ( .A(n1591), .B(n47087), .Z(n47086) );
  XNOR U46870 ( .A(n47088), .B(n47085), .Z(n47087) );
  XNOR U46871 ( .A(n47089), .B(n47090), .Z(n1591) );
  AND U46872 ( .A(n47091), .B(n47092), .Z(n47090) );
  XOR U46873 ( .A(n47054), .B(n47089), .Z(n47092) );
  AND U46874 ( .A(n47093), .B(n47094), .Z(n47054) );
  XNOR U46875 ( .A(n47051), .B(n47089), .Z(n47091) );
  XNOR U46876 ( .A(n47095), .B(n47096), .Z(n47051) );
  AND U46877 ( .A(n1595), .B(n47097), .Z(n47096) );
  XNOR U46878 ( .A(n47098), .B(n47099), .Z(n47097) );
  XOR U46879 ( .A(n47100), .B(n47101), .Z(n47089) );
  AND U46880 ( .A(n47102), .B(n47103), .Z(n47101) );
  XNOR U46881 ( .A(n47100), .B(n47093), .Z(n47103) );
  IV U46882 ( .A(n47064), .Z(n47093) );
  XOR U46883 ( .A(n47104), .B(n47105), .Z(n47064) );
  XOR U46884 ( .A(n47106), .B(n47094), .Z(n47105) );
  AND U46885 ( .A(n47074), .B(n47107), .Z(n47094) );
  AND U46886 ( .A(n47108), .B(n47109), .Z(n47106) );
  XOR U46887 ( .A(n47110), .B(n47104), .Z(n47108) );
  XNOR U46888 ( .A(n47061), .B(n47100), .Z(n47102) );
  XNOR U46889 ( .A(n47111), .B(n47112), .Z(n47061) );
  AND U46890 ( .A(n1595), .B(n47113), .Z(n47112) );
  XNOR U46891 ( .A(n47114), .B(n47115), .Z(n47113) );
  XOR U46892 ( .A(n47116), .B(n47117), .Z(n47100) );
  AND U46893 ( .A(n47118), .B(n47119), .Z(n47117) );
  XNOR U46894 ( .A(n47116), .B(n47074), .Z(n47119) );
  XOR U46895 ( .A(n47120), .B(n47109), .Z(n47074) );
  XNOR U46896 ( .A(n47121), .B(n47104), .Z(n47109) );
  XOR U46897 ( .A(n47122), .B(n47123), .Z(n47104) );
  AND U46898 ( .A(n47124), .B(n47125), .Z(n47123) );
  XOR U46899 ( .A(n47126), .B(n47122), .Z(n47124) );
  XNOR U46900 ( .A(n47127), .B(n47128), .Z(n47121) );
  AND U46901 ( .A(n47129), .B(n47130), .Z(n47128) );
  XOR U46902 ( .A(n47127), .B(n47131), .Z(n47129) );
  XNOR U46903 ( .A(n47110), .B(n47107), .Z(n47120) );
  AND U46904 ( .A(n47132), .B(n47133), .Z(n47107) );
  XOR U46905 ( .A(n47134), .B(n47135), .Z(n47110) );
  AND U46906 ( .A(n47136), .B(n47137), .Z(n47135) );
  XOR U46907 ( .A(n47134), .B(n47138), .Z(n47136) );
  XNOR U46908 ( .A(n47071), .B(n47116), .Z(n47118) );
  XNOR U46909 ( .A(n47139), .B(n47140), .Z(n47071) );
  AND U46910 ( .A(n1595), .B(n47141), .Z(n47140) );
  XNOR U46911 ( .A(n47142), .B(n47143), .Z(n47141) );
  XOR U46912 ( .A(n47144), .B(n47145), .Z(n47116) );
  AND U46913 ( .A(n47146), .B(n47147), .Z(n47145) );
  XNOR U46914 ( .A(n47144), .B(n47132), .Z(n47147) );
  IV U46915 ( .A(n47082), .Z(n47132) );
  XNOR U46916 ( .A(n47148), .B(n47125), .Z(n47082) );
  XNOR U46917 ( .A(n47149), .B(n47131), .Z(n47125) );
  XNOR U46918 ( .A(n47150), .B(n47151), .Z(n47131) );
  NOR U46919 ( .A(n47152), .B(n47153), .Z(n47151) );
  XOR U46920 ( .A(n47150), .B(n47154), .Z(n47152) );
  XNOR U46921 ( .A(n47130), .B(n47122), .Z(n47149) );
  XOR U46922 ( .A(n47155), .B(n47156), .Z(n47122) );
  AND U46923 ( .A(n47157), .B(n47158), .Z(n47156) );
  XOR U46924 ( .A(n47155), .B(n47159), .Z(n47157) );
  XNOR U46925 ( .A(n47160), .B(n47127), .Z(n47130) );
  XOR U46926 ( .A(n47161), .B(n47162), .Z(n47127) );
  AND U46927 ( .A(n47163), .B(n47164), .Z(n47162) );
  XNOR U46928 ( .A(n47165), .B(n47166), .Z(n47163) );
  IV U46929 ( .A(n47161), .Z(n47165) );
  XNOR U46930 ( .A(n47167), .B(n47168), .Z(n47160) );
  NOR U46931 ( .A(n47169), .B(n47170), .Z(n47168) );
  XNOR U46932 ( .A(n47167), .B(n47171), .Z(n47169) );
  XNOR U46933 ( .A(n47126), .B(n47133), .Z(n47148) );
  NOR U46934 ( .A(n47088), .B(n47172), .Z(n47133) );
  XOR U46935 ( .A(n47138), .B(n47137), .Z(n47126) );
  XNOR U46936 ( .A(n47173), .B(n47134), .Z(n47137) );
  XOR U46937 ( .A(n47174), .B(n47175), .Z(n47134) );
  AND U46938 ( .A(n47176), .B(n47177), .Z(n47175) );
  XNOR U46939 ( .A(n47178), .B(n47179), .Z(n47176) );
  IV U46940 ( .A(n47174), .Z(n47178) );
  XNOR U46941 ( .A(n47180), .B(n47181), .Z(n47173) );
  NOR U46942 ( .A(n47182), .B(n47183), .Z(n47181) );
  XNOR U46943 ( .A(n47180), .B(n47184), .Z(n47182) );
  XOR U46944 ( .A(n47185), .B(n47186), .Z(n47138) );
  NOR U46945 ( .A(n47187), .B(n47188), .Z(n47186) );
  XNOR U46946 ( .A(n47185), .B(n47189), .Z(n47187) );
  XNOR U46947 ( .A(n47079), .B(n47144), .Z(n47146) );
  XNOR U46948 ( .A(n47190), .B(n47191), .Z(n47079) );
  AND U46949 ( .A(n1595), .B(n47192), .Z(n47191) );
  XNOR U46950 ( .A(n47193), .B(n47194), .Z(n47192) );
  AND U46951 ( .A(n47085), .B(n47088), .Z(n47144) );
  XOR U46952 ( .A(n47195), .B(n47172), .Z(n47088) );
  XNOR U46953 ( .A(p_input[1280]), .B(p_input[2048]), .Z(n47172) );
  XNOR U46954 ( .A(n47159), .B(n47158), .Z(n47195) );
  XNOR U46955 ( .A(n47196), .B(n47166), .Z(n47158) );
  XNOR U46956 ( .A(n47154), .B(n47153), .Z(n47166) );
  XNOR U46957 ( .A(n47197), .B(n47150), .Z(n47153) );
  XNOR U46958 ( .A(p_input[1290]), .B(p_input[2058]), .Z(n47150) );
  XOR U46959 ( .A(p_input[1291]), .B(n29030), .Z(n47197) );
  XOR U46960 ( .A(p_input[1292]), .B(p_input[2060]), .Z(n47154) );
  XOR U46961 ( .A(n47164), .B(n47198), .Z(n47196) );
  IV U46962 ( .A(n47155), .Z(n47198) );
  XOR U46963 ( .A(p_input[1281]), .B(p_input[2049]), .Z(n47155) );
  XNOR U46964 ( .A(n47199), .B(n47171), .Z(n47164) );
  XNOR U46965 ( .A(p_input[1295]), .B(n29033), .Z(n47171) );
  XOR U46966 ( .A(n47161), .B(n47170), .Z(n47199) );
  XOR U46967 ( .A(n47200), .B(n47167), .Z(n47170) );
  XOR U46968 ( .A(p_input[1293]), .B(p_input[2061]), .Z(n47167) );
  XOR U46969 ( .A(p_input[1294]), .B(n29035), .Z(n47200) );
  XOR U46970 ( .A(p_input[1289]), .B(p_input[2057]), .Z(n47161) );
  XOR U46971 ( .A(n47179), .B(n47177), .Z(n47159) );
  XNOR U46972 ( .A(n47201), .B(n47184), .Z(n47177) );
  XOR U46973 ( .A(p_input[1288]), .B(p_input[2056]), .Z(n47184) );
  XOR U46974 ( .A(n47174), .B(n47183), .Z(n47201) );
  XOR U46975 ( .A(n47202), .B(n47180), .Z(n47183) );
  XOR U46976 ( .A(p_input[1286]), .B(p_input[2054]), .Z(n47180) );
  XOR U46977 ( .A(p_input[1287]), .B(n30404), .Z(n47202) );
  XOR U46978 ( .A(p_input[1282]), .B(p_input[2050]), .Z(n47174) );
  XNOR U46979 ( .A(n47189), .B(n47188), .Z(n47179) );
  XOR U46980 ( .A(n47203), .B(n47185), .Z(n47188) );
  XOR U46981 ( .A(p_input[1283]), .B(p_input[2051]), .Z(n47185) );
  XOR U46982 ( .A(p_input[1284]), .B(n30406), .Z(n47203) );
  XOR U46983 ( .A(p_input[1285]), .B(p_input[2053]), .Z(n47189) );
  XNOR U46984 ( .A(n47204), .B(n47205), .Z(n47085) );
  AND U46985 ( .A(n1595), .B(n47206), .Z(n47205) );
  XNOR U46986 ( .A(n47207), .B(n47208), .Z(n1595) );
  AND U46987 ( .A(n47209), .B(n47210), .Z(n47208) );
  XOR U46988 ( .A(n47099), .B(n47207), .Z(n47210) );
  XNOR U46989 ( .A(n47211), .B(n47207), .Z(n47209) );
  XOR U46990 ( .A(n47212), .B(n47213), .Z(n47207) );
  AND U46991 ( .A(n47214), .B(n47215), .Z(n47213) );
  XOR U46992 ( .A(n47114), .B(n47212), .Z(n47215) );
  XOR U46993 ( .A(n47212), .B(n47115), .Z(n47214) );
  XOR U46994 ( .A(n47216), .B(n47217), .Z(n47212) );
  AND U46995 ( .A(n47218), .B(n47219), .Z(n47217) );
  XOR U46996 ( .A(n47142), .B(n47216), .Z(n47219) );
  XOR U46997 ( .A(n47216), .B(n47143), .Z(n47218) );
  XOR U46998 ( .A(n47220), .B(n47221), .Z(n47216) );
  AND U46999 ( .A(n47222), .B(n47223), .Z(n47221) );
  XOR U47000 ( .A(n47220), .B(n47193), .Z(n47223) );
  XNOR U47001 ( .A(n47224), .B(n47225), .Z(n47045) );
  AND U47002 ( .A(n1599), .B(n47226), .Z(n47225) );
  XNOR U47003 ( .A(n47227), .B(n47228), .Z(n1599) );
  AND U47004 ( .A(n47229), .B(n47230), .Z(n47228) );
  XOR U47005 ( .A(n47227), .B(n47055), .Z(n47230) );
  XNOR U47006 ( .A(n47227), .B(n47015), .Z(n47229) );
  XOR U47007 ( .A(n47231), .B(n47232), .Z(n47227) );
  AND U47008 ( .A(n47233), .B(n47234), .Z(n47232) );
  XOR U47009 ( .A(n47231), .B(n47023), .Z(n47233) );
  XOR U47010 ( .A(n47235), .B(n47236), .Z(n47006) );
  AND U47011 ( .A(n1603), .B(n47226), .Z(n47236) );
  XNOR U47012 ( .A(n47224), .B(n47235), .Z(n47226) );
  XNOR U47013 ( .A(n47237), .B(n47238), .Z(n1603) );
  AND U47014 ( .A(n47239), .B(n47240), .Z(n47238) );
  XNOR U47015 ( .A(n47241), .B(n47237), .Z(n47240) );
  IV U47016 ( .A(n47055), .Z(n47241) );
  XOR U47017 ( .A(n47211), .B(n47242), .Z(n47055) );
  AND U47018 ( .A(n1606), .B(n47243), .Z(n47242) );
  XOR U47019 ( .A(n47098), .B(n47095), .Z(n47243) );
  IV U47020 ( .A(n47211), .Z(n47098) );
  XNOR U47021 ( .A(n47015), .B(n47237), .Z(n47239) );
  XOR U47022 ( .A(n47244), .B(n47245), .Z(n47015) );
  AND U47023 ( .A(n1622), .B(n47246), .Z(n47245) );
  XOR U47024 ( .A(n47231), .B(n47247), .Z(n47237) );
  AND U47025 ( .A(n47248), .B(n47234), .Z(n47247) );
  XNOR U47026 ( .A(n47065), .B(n47231), .Z(n47234) );
  XOR U47027 ( .A(n47115), .B(n47249), .Z(n47065) );
  AND U47028 ( .A(n1606), .B(n47250), .Z(n47249) );
  XOR U47029 ( .A(n47111), .B(n47115), .Z(n47250) );
  XNOR U47030 ( .A(n47251), .B(n47231), .Z(n47248) );
  IV U47031 ( .A(n47023), .Z(n47251) );
  XOR U47032 ( .A(n47252), .B(n47253), .Z(n47023) );
  AND U47033 ( .A(n1622), .B(n47254), .Z(n47253) );
  XOR U47034 ( .A(n47255), .B(n47256), .Z(n47231) );
  AND U47035 ( .A(n47257), .B(n47258), .Z(n47256) );
  XNOR U47036 ( .A(n47075), .B(n47255), .Z(n47258) );
  XOR U47037 ( .A(n47143), .B(n47259), .Z(n47075) );
  AND U47038 ( .A(n1606), .B(n47260), .Z(n47259) );
  XOR U47039 ( .A(n47139), .B(n47143), .Z(n47260) );
  XOR U47040 ( .A(n47255), .B(n47032), .Z(n47257) );
  XOR U47041 ( .A(n47261), .B(n47262), .Z(n47032) );
  AND U47042 ( .A(n1622), .B(n47263), .Z(n47262) );
  XOR U47043 ( .A(n47264), .B(n47265), .Z(n47255) );
  AND U47044 ( .A(n47266), .B(n47267), .Z(n47265) );
  XNOR U47045 ( .A(n47264), .B(n47083), .Z(n47267) );
  XOR U47046 ( .A(n47194), .B(n47268), .Z(n47083) );
  AND U47047 ( .A(n1606), .B(n47269), .Z(n47268) );
  XOR U47048 ( .A(n47190), .B(n47194), .Z(n47269) );
  XNOR U47049 ( .A(n47270), .B(n47264), .Z(n47266) );
  IV U47050 ( .A(n47042), .Z(n47270) );
  XOR U47051 ( .A(n47271), .B(n47272), .Z(n47042) );
  AND U47052 ( .A(n1622), .B(n47273), .Z(n47272) );
  AND U47053 ( .A(n47235), .B(n47224), .Z(n47264) );
  XNOR U47054 ( .A(n47274), .B(n47275), .Z(n47224) );
  AND U47055 ( .A(n1606), .B(n47206), .Z(n47275) );
  XNOR U47056 ( .A(n47204), .B(n47274), .Z(n47206) );
  XNOR U47057 ( .A(n47276), .B(n47277), .Z(n1606) );
  AND U47058 ( .A(n47278), .B(n47279), .Z(n47277) );
  XNOR U47059 ( .A(n47276), .B(n47095), .Z(n47279) );
  IV U47060 ( .A(n47099), .Z(n47095) );
  XOR U47061 ( .A(n47280), .B(n47281), .Z(n47099) );
  AND U47062 ( .A(n1610), .B(n47282), .Z(n47281) );
  XOR U47063 ( .A(n47283), .B(n47280), .Z(n47282) );
  XNOR U47064 ( .A(n47276), .B(n47211), .Z(n47278) );
  XOR U47065 ( .A(n47284), .B(n47285), .Z(n47211) );
  AND U47066 ( .A(n1618), .B(n47246), .Z(n47285) );
  XOR U47067 ( .A(n47244), .B(n47284), .Z(n47246) );
  XOR U47068 ( .A(n47286), .B(n47287), .Z(n47276) );
  AND U47069 ( .A(n47288), .B(n47289), .Z(n47287) );
  XNOR U47070 ( .A(n47286), .B(n47111), .Z(n47289) );
  IV U47071 ( .A(n47114), .Z(n47111) );
  XOR U47072 ( .A(n47290), .B(n47291), .Z(n47114) );
  AND U47073 ( .A(n1610), .B(n47292), .Z(n47291) );
  XOR U47074 ( .A(n47293), .B(n47290), .Z(n47292) );
  XOR U47075 ( .A(n47115), .B(n47286), .Z(n47288) );
  XOR U47076 ( .A(n47294), .B(n47295), .Z(n47115) );
  AND U47077 ( .A(n1618), .B(n47254), .Z(n47295) );
  XOR U47078 ( .A(n47294), .B(n47252), .Z(n47254) );
  XOR U47079 ( .A(n47296), .B(n47297), .Z(n47286) );
  AND U47080 ( .A(n47298), .B(n47299), .Z(n47297) );
  XNOR U47081 ( .A(n47296), .B(n47139), .Z(n47299) );
  IV U47082 ( .A(n47142), .Z(n47139) );
  XOR U47083 ( .A(n47300), .B(n47301), .Z(n47142) );
  AND U47084 ( .A(n1610), .B(n47302), .Z(n47301) );
  XNOR U47085 ( .A(n47303), .B(n47300), .Z(n47302) );
  XOR U47086 ( .A(n47143), .B(n47296), .Z(n47298) );
  XOR U47087 ( .A(n47304), .B(n47305), .Z(n47143) );
  AND U47088 ( .A(n1618), .B(n47263), .Z(n47305) );
  XOR U47089 ( .A(n47304), .B(n47261), .Z(n47263) );
  XOR U47090 ( .A(n47220), .B(n47306), .Z(n47296) );
  AND U47091 ( .A(n47222), .B(n47307), .Z(n47306) );
  XNOR U47092 ( .A(n47220), .B(n47190), .Z(n47307) );
  IV U47093 ( .A(n47193), .Z(n47190) );
  XOR U47094 ( .A(n47308), .B(n47309), .Z(n47193) );
  AND U47095 ( .A(n1610), .B(n47310), .Z(n47309) );
  XOR U47096 ( .A(n47311), .B(n47308), .Z(n47310) );
  XOR U47097 ( .A(n47194), .B(n47220), .Z(n47222) );
  XOR U47098 ( .A(n47312), .B(n47313), .Z(n47194) );
  AND U47099 ( .A(n1618), .B(n47273), .Z(n47313) );
  XOR U47100 ( .A(n47312), .B(n47271), .Z(n47273) );
  AND U47101 ( .A(n47274), .B(n47204), .Z(n47220) );
  XNOR U47102 ( .A(n47314), .B(n47315), .Z(n47204) );
  AND U47103 ( .A(n1610), .B(n47316), .Z(n47315) );
  XNOR U47104 ( .A(n47317), .B(n47314), .Z(n47316) );
  XNOR U47105 ( .A(n47318), .B(n47319), .Z(n1610) );
  AND U47106 ( .A(n47320), .B(n47321), .Z(n47319) );
  XOR U47107 ( .A(n47283), .B(n47318), .Z(n47321) );
  AND U47108 ( .A(n47322), .B(n47323), .Z(n47283) );
  XNOR U47109 ( .A(n47280), .B(n47318), .Z(n47320) );
  XNOR U47110 ( .A(n47324), .B(n47325), .Z(n47280) );
  AND U47111 ( .A(n1614), .B(n47326), .Z(n47325) );
  XNOR U47112 ( .A(n47327), .B(n47328), .Z(n47326) );
  XOR U47113 ( .A(n47329), .B(n47330), .Z(n47318) );
  AND U47114 ( .A(n47331), .B(n47332), .Z(n47330) );
  XNOR U47115 ( .A(n47329), .B(n47322), .Z(n47332) );
  IV U47116 ( .A(n47293), .Z(n47322) );
  XOR U47117 ( .A(n47333), .B(n47334), .Z(n47293) );
  XOR U47118 ( .A(n47335), .B(n47323), .Z(n47334) );
  AND U47119 ( .A(n47303), .B(n47336), .Z(n47323) );
  AND U47120 ( .A(n47337), .B(n47338), .Z(n47335) );
  XOR U47121 ( .A(n47339), .B(n47333), .Z(n47337) );
  XNOR U47122 ( .A(n47290), .B(n47329), .Z(n47331) );
  XNOR U47123 ( .A(n47340), .B(n47341), .Z(n47290) );
  AND U47124 ( .A(n1614), .B(n47342), .Z(n47341) );
  XNOR U47125 ( .A(n47343), .B(n47344), .Z(n47342) );
  XOR U47126 ( .A(n47345), .B(n47346), .Z(n47329) );
  AND U47127 ( .A(n47347), .B(n47348), .Z(n47346) );
  XNOR U47128 ( .A(n47345), .B(n47303), .Z(n47348) );
  XOR U47129 ( .A(n47349), .B(n47338), .Z(n47303) );
  XNOR U47130 ( .A(n47350), .B(n47333), .Z(n47338) );
  XOR U47131 ( .A(n47351), .B(n47352), .Z(n47333) );
  AND U47132 ( .A(n47353), .B(n47354), .Z(n47352) );
  XOR U47133 ( .A(n47355), .B(n47351), .Z(n47353) );
  XNOR U47134 ( .A(n47356), .B(n47357), .Z(n47350) );
  AND U47135 ( .A(n47358), .B(n47359), .Z(n47357) );
  XOR U47136 ( .A(n47356), .B(n47360), .Z(n47358) );
  XNOR U47137 ( .A(n47339), .B(n47336), .Z(n47349) );
  AND U47138 ( .A(n47361), .B(n47362), .Z(n47336) );
  XOR U47139 ( .A(n47363), .B(n47364), .Z(n47339) );
  AND U47140 ( .A(n47365), .B(n47366), .Z(n47364) );
  XOR U47141 ( .A(n47363), .B(n47367), .Z(n47365) );
  XNOR U47142 ( .A(n47300), .B(n47345), .Z(n47347) );
  XNOR U47143 ( .A(n47368), .B(n47369), .Z(n47300) );
  AND U47144 ( .A(n1614), .B(n47370), .Z(n47369) );
  XNOR U47145 ( .A(n47371), .B(n47372), .Z(n47370) );
  XOR U47146 ( .A(n47373), .B(n47374), .Z(n47345) );
  AND U47147 ( .A(n47375), .B(n47376), .Z(n47374) );
  XNOR U47148 ( .A(n47373), .B(n47361), .Z(n47376) );
  IV U47149 ( .A(n47311), .Z(n47361) );
  XNOR U47150 ( .A(n47377), .B(n47354), .Z(n47311) );
  XNOR U47151 ( .A(n47378), .B(n47360), .Z(n47354) );
  XNOR U47152 ( .A(n47379), .B(n47380), .Z(n47360) );
  NOR U47153 ( .A(n47381), .B(n47382), .Z(n47380) );
  XOR U47154 ( .A(n47379), .B(n47383), .Z(n47381) );
  XNOR U47155 ( .A(n47359), .B(n47351), .Z(n47378) );
  XOR U47156 ( .A(n47384), .B(n47385), .Z(n47351) );
  AND U47157 ( .A(n47386), .B(n47387), .Z(n47385) );
  XOR U47158 ( .A(n47384), .B(n47388), .Z(n47386) );
  XNOR U47159 ( .A(n47389), .B(n47356), .Z(n47359) );
  XOR U47160 ( .A(n47390), .B(n47391), .Z(n47356) );
  AND U47161 ( .A(n47392), .B(n47393), .Z(n47391) );
  XNOR U47162 ( .A(n47394), .B(n47395), .Z(n47392) );
  IV U47163 ( .A(n47390), .Z(n47394) );
  XNOR U47164 ( .A(n47396), .B(n47397), .Z(n47389) );
  NOR U47165 ( .A(n47398), .B(n47399), .Z(n47397) );
  XNOR U47166 ( .A(n47396), .B(n47400), .Z(n47398) );
  XNOR U47167 ( .A(n47355), .B(n47362), .Z(n47377) );
  NOR U47168 ( .A(n47317), .B(n47401), .Z(n47362) );
  XOR U47169 ( .A(n47367), .B(n47366), .Z(n47355) );
  XNOR U47170 ( .A(n47402), .B(n47363), .Z(n47366) );
  XOR U47171 ( .A(n47403), .B(n47404), .Z(n47363) );
  AND U47172 ( .A(n47405), .B(n47406), .Z(n47404) );
  XNOR U47173 ( .A(n47407), .B(n47408), .Z(n47405) );
  IV U47174 ( .A(n47403), .Z(n47407) );
  XNOR U47175 ( .A(n47409), .B(n47410), .Z(n47402) );
  NOR U47176 ( .A(n47411), .B(n47412), .Z(n47410) );
  XNOR U47177 ( .A(n47409), .B(n47413), .Z(n47411) );
  XOR U47178 ( .A(n47414), .B(n47415), .Z(n47367) );
  NOR U47179 ( .A(n47416), .B(n47417), .Z(n47415) );
  XNOR U47180 ( .A(n47414), .B(n47418), .Z(n47416) );
  XNOR U47181 ( .A(n47308), .B(n47373), .Z(n47375) );
  XNOR U47182 ( .A(n47419), .B(n47420), .Z(n47308) );
  AND U47183 ( .A(n1614), .B(n47421), .Z(n47420) );
  XNOR U47184 ( .A(n47422), .B(n47423), .Z(n47421) );
  AND U47185 ( .A(n47314), .B(n47317), .Z(n47373) );
  XOR U47186 ( .A(n47424), .B(n47401), .Z(n47317) );
  XNOR U47187 ( .A(p_input[1296]), .B(p_input[2048]), .Z(n47401) );
  XNOR U47188 ( .A(n47388), .B(n47387), .Z(n47424) );
  XNOR U47189 ( .A(n47425), .B(n47395), .Z(n47387) );
  XNOR U47190 ( .A(n47383), .B(n47382), .Z(n47395) );
  XNOR U47191 ( .A(n47426), .B(n47379), .Z(n47382) );
  XNOR U47192 ( .A(p_input[1306]), .B(p_input[2058]), .Z(n47379) );
  XOR U47193 ( .A(p_input[1307]), .B(n29030), .Z(n47426) );
  XOR U47194 ( .A(p_input[1308]), .B(p_input[2060]), .Z(n47383) );
  XOR U47195 ( .A(n47393), .B(n47427), .Z(n47425) );
  IV U47196 ( .A(n47384), .Z(n47427) );
  XOR U47197 ( .A(p_input[1297]), .B(p_input[2049]), .Z(n47384) );
  XNOR U47198 ( .A(n47428), .B(n47400), .Z(n47393) );
  XNOR U47199 ( .A(p_input[1311]), .B(n29033), .Z(n47400) );
  XOR U47200 ( .A(n47390), .B(n47399), .Z(n47428) );
  XOR U47201 ( .A(n47429), .B(n47396), .Z(n47399) );
  XOR U47202 ( .A(p_input[1309]), .B(p_input[2061]), .Z(n47396) );
  XOR U47203 ( .A(p_input[1310]), .B(n29035), .Z(n47429) );
  XOR U47204 ( .A(p_input[1305]), .B(p_input[2057]), .Z(n47390) );
  XOR U47205 ( .A(n47408), .B(n47406), .Z(n47388) );
  XNOR U47206 ( .A(n47430), .B(n47413), .Z(n47406) );
  XOR U47207 ( .A(p_input[1304]), .B(p_input[2056]), .Z(n47413) );
  XOR U47208 ( .A(n47403), .B(n47412), .Z(n47430) );
  XOR U47209 ( .A(n47431), .B(n47409), .Z(n47412) );
  XOR U47210 ( .A(p_input[1302]), .B(p_input[2054]), .Z(n47409) );
  XOR U47211 ( .A(p_input[1303]), .B(n30404), .Z(n47431) );
  XOR U47212 ( .A(p_input[1298]), .B(p_input[2050]), .Z(n47403) );
  XNOR U47213 ( .A(n47418), .B(n47417), .Z(n47408) );
  XOR U47214 ( .A(n47432), .B(n47414), .Z(n47417) );
  XOR U47215 ( .A(p_input[1299]), .B(p_input[2051]), .Z(n47414) );
  XOR U47216 ( .A(p_input[1300]), .B(n30406), .Z(n47432) );
  XOR U47217 ( .A(p_input[1301]), .B(p_input[2053]), .Z(n47418) );
  XNOR U47218 ( .A(n47433), .B(n47434), .Z(n47314) );
  AND U47219 ( .A(n1614), .B(n47435), .Z(n47434) );
  XNOR U47220 ( .A(n47436), .B(n47437), .Z(n1614) );
  AND U47221 ( .A(n47438), .B(n47439), .Z(n47437) );
  XOR U47222 ( .A(n47328), .B(n47436), .Z(n47439) );
  XNOR U47223 ( .A(n47440), .B(n47436), .Z(n47438) );
  XOR U47224 ( .A(n47441), .B(n47442), .Z(n47436) );
  AND U47225 ( .A(n47443), .B(n47444), .Z(n47442) );
  XOR U47226 ( .A(n47343), .B(n47441), .Z(n47444) );
  XOR U47227 ( .A(n47441), .B(n47344), .Z(n47443) );
  XOR U47228 ( .A(n47445), .B(n47446), .Z(n47441) );
  AND U47229 ( .A(n47447), .B(n47448), .Z(n47446) );
  XOR U47230 ( .A(n47371), .B(n47445), .Z(n47448) );
  XOR U47231 ( .A(n47445), .B(n47372), .Z(n47447) );
  XOR U47232 ( .A(n47449), .B(n47450), .Z(n47445) );
  AND U47233 ( .A(n47451), .B(n47452), .Z(n47450) );
  XOR U47234 ( .A(n47449), .B(n47422), .Z(n47452) );
  XNOR U47235 ( .A(n47453), .B(n47454), .Z(n47274) );
  AND U47236 ( .A(n1618), .B(n47455), .Z(n47454) );
  XNOR U47237 ( .A(n47456), .B(n47457), .Z(n1618) );
  AND U47238 ( .A(n47458), .B(n47459), .Z(n47457) );
  XOR U47239 ( .A(n47456), .B(n47284), .Z(n47459) );
  XNOR U47240 ( .A(n47456), .B(n47244), .Z(n47458) );
  XOR U47241 ( .A(n47460), .B(n47461), .Z(n47456) );
  AND U47242 ( .A(n47462), .B(n47463), .Z(n47461) );
  XOR U47243 ( .A(n47460), .B(n47252), .Z(n47462) );
  XOR U47244 ( .A(n47464), .B(n47465), .Z(n47235) );
  AND U47245 ( .A(n1622), .B(n47455), .Z(n47465) );
  XNOR U47246 ( .A(n47453), .B(n47464), .Z(n47455) );
  XNOR U47247 ( .A(n47466), .B(n47467), .Z(n1622) );
  AND U47248 ( .A(n47468), .B(n47469), .Z(n47467) );
  XNOR U47249 ( .A(n47470), .B(n47466), .Z(n47469) );
  IV U47250 ( .A(n47284), .Z(n47470) );
  XOR U47251 ( .A(n47440), .B(n47471), .Z(n47284) );
  AND U47252 ( .A(n1625), .B(n47472), .Z(n47471) );
  XOR U47253 ( .A(n47327), .B(n47324), .Z(n47472) );
  IV U47254 ( .A(n47440), .Z(n47327) );
  XNOR U47255 ( .A(n47244), .B(n47466), .Z(n47468) );
  XOR U47256 ( .A(n47473), .B(n47474), .Z(n47244) );
  AND U47257 ( .A(n1641), .B(n47475), .Z(n47474) );
  XOR U47258 ( .A(n47460), .B(n47476), .Z(n47466) );
  AND U47259 ( .A(n47477), .B(n47463), .Z(n47476) );
  XNOR U47260 ( .A(n47294), .B(n47460), .Z(n47463) );
  XOR U47261 ( .A(n47344), .B(n47478), .Z(n47294) );
  AND U47262 ( .A(n1625), .B(n47479), .Z(n47478) );
  XOR U47263 ( .A(n47340), .B(n47344), .Z(n47479) );
  XNOR U47264 ( .A(n47480), .B(n47460), .Z(n47477) );
  IV U47265 ( .A(n47252), .Z(n47480) );
  XOR U47266 ( .A(n47481), .B(n47482), .Z(n47252) );
  AND U47267 ( .A(n1641), .B(n47483), .Z(n47482) );
  XOR U47268 ( .A(n47484), .B(n47485), .Z(n47460) );
  AND U47269 ( .A(n47486), .B(n47487), .Z(n47485) );
  XNOR U47270 ( .A(n47304), .B(n47484), .Z(n47487) );
  XOR U47271 ( .A(n47372), .B(n47488), .Z(n47304) );
  AND U47272 ( .A(n1625), .B(n47489), .Z(n47488) );
  XOR U47273 ( .A(n47368), .B(n47372), .Z(n47489) );
  XOR U47274 ( .A(n47484), .B(n47261), .Z(n47486) );
  XOR U47275 ( .A(n47490), .B(n47491), .Z(n47261) );
  AND U47276 ( .A(n1641), .B(n47492), .Z(n47491) );
  XOR U47277 ( .A(n47493), .B(n47494), .Z(n47484) );
  AND U47278 ( .A(n47495), .B(n47496), .Z(n47494) );
  XNOR U47279 ( .A(n47493), .B(n47312), .Z(n47496) );
  XOR U47280 ( .A(n47423), .B(n47497), .Z(n47312) );
  AND U47281 ( .A(n1625), .B(n47498), .Z(n47497) );
  XOR U47282 ( .A(n47419), .B(n47423), .Z(n47498) );
  XNOR U47283 ( .A(n47499), .B(n47493), .Z(n47495) );
  IV U47284 ( .A(n47271), .Z(n47499) );
  XOR U47285 ( .A(n47500), .B(n47501), .Z(n47271) );
  AND U47286 ( .A(n1641), .B(n47502), .Z(n47501) );
  AND U47287 ( .A(n47464), .B(n47453), .Z(n47493) );
  XNOR U47288 ( .A(n47503), .B(n47504), .Z(n47453) );
  AND U47289 ( .A(n1625), .B(n47435), .Z(n47504) );
  XNOR U47290 ( .A(n47433), .B(n47503), .Z(n47435) );
  XNOR U47291 ( .A(n47505), .B(n47506), .Z(n1625) );
  AND U47292 ( .A(n47507), .B(n47508), .Z(n47506) );
  XNOR U47293 ( .A(n47505), .B(n47324), .Z(n47508) );
  IV U47294 ( .A(n47328), .Z(n47324) );
  XOR U47295 ( .A(n47509), .B(n47510), .Z(n47328) );
  AND U47296 ( .A(n1629), .B(n47511), .Z(n47510) );
  XOR U47297 ( .A(n47512), .B(n47509), .Z(n47511) );
  XNOR U47298 ( .A(n47505), .B(n47440), .Z(n47507) );
  XOR U47299 ( .A(n47513), .B(n47514), .Z(n47440) );
  AND U47300 ( .A(n1637), .B(n47475), .Z(n47514) );
  XOR U47301 ( .A(n47473), .B(n47513), .Z(n47475) );
  XOR U47302 ( .A(n47515), .B(n47516), .Z(n47505) );
  AND U47303 ( .A(n47517), .B(n47518), .Z(n47516) );
  XNOR U47304 ( .A(n47515), .B(n47340), .Z(n47518) );
  IV U47305 ( .A(n47343), .Z(n47340) );
  XOR U47306 ( .A(n47519), .B(n47520), .Z(n47343) );
  AND U47307 ( .A(n1629), .B(n47521), .Z(n47520) );
  XOR U47308 ( .A(n47522), .B(n47519), .Z(n47521) );
  XOR U47309 ( .A(n47344), .B(n47515), .Z(n47517) );
  XOR U47310 ( .A(n47523), .B(n47524), .Z(n47344) );
  AND U47311 ( .A(n1637), .B(n47483), .Z(n47524) );
  XOR U47312 ( .A(n47523), .B(n47481), .Z(n47483) );
  XOR U47313 ( .A(n47525), .B(n47526), .Z(n47515) );
  AND U47314 ( .A(n47527), .B(n47528), .Z(n47526) );
  XNOR U47315 ( .A(n47525), .B(n47368), .Z(n47528) );
  IV U47316 ( .A(n47371), .Z(n47368) );
  XOR U47317 ( .A(n47529), .B(n47530), .Z(n47371) );
  AND U47318 ( .A(n1629), .B(n47531), .Z(n47530) );
  XNOR U47319 ( .A(n47532), .B(n47529), .Z(n47531) );
  XOR U47320 ( .A(n47372), .B(n47525), .Z(n47527) );
  XOR U47321 ( .A(n47533), .B(n47534), .Z(n47372) );
  AND U47322 ( .A(n1637), .B(n47492), .Z(n47534) );
  XOR U47323 ( .A(n47533), .B(n47490), .Z(n47492) );
  XOR U47324 ( .A(n47449), .B(n47535), .Z(n47525) );
  AND U47325 ( .A(n47451), .B(n47536), .Z(n47535) );
  XNOR U47326 ( .A(n47449), .B(n47419), .Z(n47536) );
  IV U47327 ( .A(n47422), .Z(n47419) );
  XOR U47328 ( .A(n47537), .B(n47538), .Z(n47422) );
  AND U47329 ( .A(n1629), .B(n47539), .Z(n47538) );
  XOR U47330 ( .A(n47540), .B(n47537), .Z(n47539) );
  XOR U47331 ( .A(n47423), .B(n47449), .Z(n47451) );
  XOR U47332 ( .A(n47541), .B(n47542), .Z(n47423) );
  AND U47333 ( .A(n1637), .B(n47502), .Z(n47542) );
  XOR U47334 ( .A(n47541), .B(n47500), .Z(n47502) );
  AND U47335 ( .A(n47503), .B(n47433), .Z(n47449) );
  XNOR U47336 ( .A(n47543), .B(n47544), .Z(n47433) );
  AND U47337 ( .A(n1629), .B(n47545), .Z(n47544) );
  XNOR U47338 ( .A(n47546), .B(n47543), .Z(n47545) );
  XNOR U47339 ( .A(n47547), .B(n47548), .Z(n1629) );
  AND U47340 ( .A(n47549), .B(n47550), .Z(n47548) );
  XOR U47341 ( .A(n47512), .B(n47547), .Z(n47550) );
  AND U47342 ( .A(n47551), .B(n47552), .Z(n47512) );
  XNOR U47343 ( .A(n47509), .B(n47547), .Z(n47549) );
  XNOR U47344 ( .A(n47553), .B(n47554), .Z(n47509) );
  AND U47345 ( .A(n1633), .B(n47555), .Z(n47554) );
  XNOR U47346 ( .A(n47556), .B(n47557), .Z(n47555) );
  XOR U47347 ( .A(n47558), .B(n47559), .Z(n47547) );
  AND U47348 ( .A(n47560), .B(n47561), .Z(n47559) );
  XNOR U47349 ( .A(n47558), .B(n47551), .Z(n47561) );
  IV U47350 ( .A(n47522), .Z(n47551) );
  XOR U47351 ( .A(n47562), .B(n47563), .Z(n47522) );
  XOR U47352 ( .A(n47564), .B(n47552), .Z(n47563) );
  AND U47353 ( .A(n47532), .B(n47565), .Z(n47552) );
  AND U47354 ( .A(n47566), .B(n47567), .Z(n47564) );
  XOR U47355 ( .A(n47568), .B(n47562), .Z(n47566) );
  XNOR U47356 ( .A(n47519), .B(n47558), .Z(n47560) );
  XNOR U47357 ( .A(n47569), .B(n47570), .Z(n47519) );
  AND U47358 ( .A(n1633), .B(n47571), .Z(n47570) );
  XNOR U47359 ( .A(n47572), .B(n47573), .Z(n47571) );
  XOR U47360 ( .A(n47574), .B(n47575), .Z(n47558) );
  AND U47361 ( .A(n47576), .B(n47577), .Z(n47575) );
  XNOR U47362 ( .A(n47574), .B(n47532), .Z(n47577) );
  XOR U47363 ( .A(n47578), .B(n47567), .Z(n47532) );
  XNOR U47364 ( .A(n47579), .B(n47562), .Z(n47567) );
  XOR U47365 ( .A(n47580), .B(n47581), .Z(n47562) );
  AND U47366 ( .A(n47582), .B(n47583), .Z(n47581) );
  XOR U47367 ( .A(n47584), .B(n47580), .Z(n47582) );
  XNOR U47368 ( .A(n47585), .B(n47586), .Z(n47579) );
  AND U47369 ( .A(n47587), .B(n47588), .Z(n47586) );
  XOR U47370 ( .A(n47585), .B(n47589), .Z(n47587) );
  XNOR U47371 ( .A(n47568), .B(n47565), .Z(n47578) );
  AND U47372 ( .A(n47590), .B(n47591), .Z(n47565) );
  XOR U47373 ( .A(n47592), .B(n47593), .Z(n47568) );
  AND U47374 ( .A(n47594), .B(n47595), .Z(n47593) );
  XOR U47375 ( .A(n47592), .B(n47596), .Z(n47594) );
  XNOR U47376 ( .A(n47529), .B(n47574), .Z(n47576) );
  XNOR U47377 ( .A(n47597), .B(n47598), .Z(n47529) );
  AND U47378 ( .A(n1633), .B(n47599), .Z(n47598) );
  XNOR U47379 ( .A(n47600), .B(n47601), .Z(n47599) );
  XOR U47380 ( .A(n47602), .B(n47603), .Z(n47574) );
  AND U47381 ( .A(n47604), .B(n47605), .Z(n47603) );
  XNOR U47382 ( .A(n47602), .B(n47590), .Z(n47605) );
  IV U47383 ( .A(n47540), .Z(n47590) );
  XNOR U47384 ( .A(n47606), .B(n47583), .Z(n47540) );
  XNOR U47385 ( .A(n47607), .B(n47589), .Z(n47583) );
  XNOR U47386 ( .A(n47608), .B(n47609), .Z(n47589) );
  NOR U47387 ( .A(n47610), .B(n47611), .Z(n47609) );
  XOR U47388 ( .A(n47608), .B(n47612), .Z(n47610) );
  XNOR U47389 ( .A(n47588), .B(n47580), .Z(n47607) );
  XOR U47390 ( .A(n47613), .B(n47614), .Z(n47580) );
  AND U47391 ( .A(n47615), .B(n47616), .Z(n47614) );
  XOR U47392 ( .A(n47613), .B(n47617), .Z(n47615) );
  XNOR U47393 ( .A(n47618), .B(n47585), .Z(n47588) );
  XOR U47394 ( .A(n47619), .B(n47620), .Z(n47585) );
  AND U47395 ( .A(n47621), .B(n47622), .Z(n47620) );
  XNOR U47396 ( .A(n47623), .B(n47624), .Z(n47621) );
  IV U47397 ( .A(n47619), .Z(n47623) );
  XNOR U47398 ( .A(n47625), .B(n47626), .Z(n47618) );
  NOR U47399 ( .A(n47627), .B(n47628), .Z(n47626) );
  XNOR U47400 ( .A(n47625), .B(n47629), .Z(n47627) );
  XNOR U47401 ( .A(n47584), .B(n47591), .Z(n47606) );
  NOR U47402 ( .A(n47546), .B(n47630), .Z(n47591) );
  XOR U47403 ( .A(n47596), .B(n47595), .Z(n47584) );
  XNOR U47404 ( .A(n47631), .B(n47592), .Z(n47595) );
  XOR U47405 ( .A(n47632), .B(n47633), .Z(n47592) );
  AND U47406 ( .A(n47634), .B(n47635), .Z(n47633) );
  XNOR U47407 ( .A(n47636), .B(n47637), .Z(n47634) );
  IV U47408 ( .A(n47632), .Z(n47636) );
  XNOR U47409 ( .A(n47638), .B(n47639), .Z(n47631) );
  NOR U47410 ( .A(n47640), .B(n47641), .Z(n47639) );
  XNOR U47411 ( .A(n47638), .B(n47642), .Z(n47640) );
  XOR U47412 ( .A(n47643), .B(n47644), .Z(n47596) );
  NOR U47413 ( .A(n47645), .B(n47646), .Z(n47644) );
  XNOR U47414 ( .A(n47643), .B(n47647), .Z(n47645) );
  XNOR U47415 ( .A(n47537), .B(n47602), .Z(n47604) );
  XNOR U47416 ( .A(n47648), .B(n47649), .Z(n47537) );
  AND U47417 ( .A(n1633), .B(n47650), .Z(n47649) );
  XNOR U47418 ( .A(n47651), .B(n47652), .Z(n47650) );
  AND U47419 ( .A(n47543), .B(n47546), .Z(n47602) );
  XOR U47420 ( .A(n47653), .B(n47630), .Z(n47546) );
  XNOR U47421 ( .A(p_input[1312]), .B(p_input[2048]), .Z(n47630) );
  XNOR U47422 ( .A(n47617), .B(n47616), .Z(n47653) );
  XNOR U47423 ( .A(n47654), .B(n47624), .Z(n47616) );
  XNOR U47424 ( .A(n47612), .B(n47611), .Z(n47624) );
  XNOR U47425 ( .A(n47655), .B(n47608), .Z(n47611) );
  XNOR U47426 ( .A(p_input[1322]), .B(p_input[2058]), .Z(n47608) );
  XOR U47427 ( .A(p_input[1323]), .B(n29030), .Z(n47655) );
  XOR U47428 ( .A(p_input[1324]), .B(p_input[2060]), .Z(n47612) );
  XOR U47429 ( .A(n47622), .B(n47656), .Z(n47654) );
  IV U47430 ( .A(n47613), .Z(n47656) );
  XOR U47431 ( .A(p_input[1313]), .B(p_input[2049]), .Z(n47613) );
  XNOR U47432 ( .A(n47657), .B(n47629), .Z(n47622) );
  XNOR U47433 ( .A(p_input[1327]), .B(n29033), .Z(n47629) );
  XOR U47434 ( .A(n47619), .B(n47628), .Z(n47657) );
  XOR U47435 ( .A(n47658), .B(n47625), .Z(n47628) );
  XOR U47436 ( .A(p_input[1325]), .B(p_input[2061]), .Z(n47625) );
  XOR U47437 ( .A(p_input[1326]), .B(n29035), .Z(n47658) );
  XOR U47438 ( .A(p_input[1321]), .B(p_input[2057]), .Z(n47619) );
  XOR U47439 ( .A(n47637), .B(n47635), .Z(n47617) );
  XNOR U47440 ( .A(n47659), .B(n47642), .Z(n47635) );
  XOR U47441 ( .A(p_input[1320]), .B(p_input[2056]), .Z(n47642) );
  XOR U47442 ( .A(n47632), .B(n47641), .Z(n47659) );
  XOR U47443 ( .A(n47660), .B(n47638), .Z(n47641) );
  XOR U47444 ( .A(p_input[1318]), .B(p_input[2054]), .Z(n47638) );
  XOR U47445 ( .A(p_input[1319]), .B(n30404), .Z(n47660) );
  XOR U47446 ( .A(p_input[1314]), .B(p_input[2050]), .Z(n47632) );
  XNOR U47447 ( .A(n47647), .B(n47646), .Z(n47637) );
  XOR U47448 ( .A(n47661), .B(n47643), .Z(n47646) );
  XOR U47449 ( .A(p_input[1315]), .B(p_input[2051]), .Z(n47643) );
  XOR U47450 ( .A(p_input[1316]), .B(n30406), .Z(n47661) );
  XOR U47451 ( .A(p_input[1317]), .B(p_input[2053]), .Z(n47647) );
  XNOR U47452 ( .A(n47662), .B(n47663), .Z(n47543) );
  AND U47453 ( .A(n1633), .B(n47664), .Z(n47663) );
  XNOR U47454 ( .A(n47665), .B(n47666), .Z(n1633) );
  AND U47455 ( .A(n47667), .B(n47668), .Z(n47666) );
  XOR U47456 ( .A(n47557), .B(n47665), .Z(n47668) );
  XNOR U47457 ( .A(n47669), .B(n47665), .Z(n47667) );
  XOR U47458 ( .A(n47670), .B(n47671), .Z(n47665) );
  AND U47459 ( .A(n47672), .B(n47673), .Z(n47671) );
  XOR U47460 ( .A(n47572), .B(n47670), .Z(n47673) );
  XOR U47461 ( .A(n47670), .B(n47573), .Z(n47672) );
  XOR U47462 ( .A(n47674), .B(n47675), .Z(n47670) );
  AND U47463 ( .A(n47676), .B(n47677), .Z(n47675) );
  XOR U47464 ( .A(n47600), .B(n47674), .Z(n47677) );
  XOR U47465 ( .A(n47674), .B(n47601), .Z(n47676) );
  XOR U47466 ( .A(n47678), .B(n47679), .Z(n47674) );
  AND U47467 ( .A(n47680), .B(n47681), .Z(n47679) );
  XOR U47468 ( .A(n47678), .B(n47651), .Z(n47681) );
  XNOR U47469 ( .A(n47682), .B(n47683), .Z(n47503) );
  AND U47470 ( .A(n1637), .B(n47684), .Z(n47683) );
  XNOR U47471 ( .A(n47685), .B(n47686), .Z(n1637) );
  AND U47472 ( .A(n47687), .B(n47688), .Z(n47686) );
  XOR U47473 ( .A(n47685), .B(n47513), .Z(n47688) );
  XNOR U47474 ( .A(n47685), .B(n47473), .Z(n47687) );
  XOR U47475 ( .A(n47689), .B(n47690), .Z(n47685) );
  AND U47476 ( .A(n47691), .B(n47692), .Z(n47690) );
  XOR U47477 ( .A(n47689), .B(n47481), .Z(n47691) );
  XOR U47478 ( .A(n47693), .B(n47694), .Z(n47464) );
  AND U47479 ( .A(n1641), .B(n47684), .Z(n47694) );
  XNOR U47480 ( .A(n47682), .B(n47693), .Z(n47684) );
  XNOR U47481 ( .A(n47695), .B(n47696), .Z(n1641) );
  AND U47482 ( .A(n47697), .B(n47698), .Z(n47696) );
  XNOR U47483 ( .A(n47699), .B(n47695), .Z(n47698) );
  IV U47484 ( .A(n47513), .Z(n47699) );
  XOR U47485 ( .A(n47669), .B(n47700), .Z(n47513) );
  AND U47486 ( .A(n1644), .B(n47701), .Z(n47700) );
  XOR U47487 ( .A(n47556), .B(n47553), .Z(n47701) );
  IV U47488 ( .A(n47669), .Z(n47556) );
  XNOR U47489 ( .A(n47473), .B(n47695), .Z(n47697) );
  XOR U47490 ( .A(n47702), .B(n47703), .Z(n47473) );
  AND U47491 ( .A(n1660), .B(n47704), .Z(n47703) );
  XOR U47492 ( .A(n47689), .B(n47705), .Z(n47695) );
  AND U47493 ( .A(n47706), .B(n47692), .Z(n47705) );
  XNOR U47494 ( .A(n47523), .B(n47689), .Z(n47692) );
  XOR U47495 ( .A(n47573), .B(n47707), .Z(n47523) );
  AND U47496 ( .A(n1644), .B(n47708), .Z(n47707) );
  XOR U47497 ( .A(n47569), .B(n47573), .Z(n47708) );
  XNOR U47498 ( .A(n47709), .B(n47689), .Z(n47706) );
  IV U47499 ( .A(n47481), .Z(n47709) );
  XOR U47500 ( .A(n47710), .B(n47711), .Z(n47481) );
  AND U47501 ( .A(n1660), .B(n47712), .Z(n47711) );
  XOR U47502 ( .A(n47713), .B(n47714), .Z(n47689) );
  AND U47503 ( .A(n47715), .B(n47716), .Z(n47714) );
  XNOR U47504 ( .A(n47533), .B(n47713), .Z(n47716) );
  XOR U47505 ( .A(n47601), .B(n47717), .Z(n47533) );
  AND U47506 ( .A(n1644), .B(n47718), .Z(n47717) );
  XOR U47507 ( .A(n47597), .B(n47601), .Z(n47718) );
  XOR U47508 ( .A(n47713), .B(n47490), .Z(n47715) );
  XOR U47509 ( .A(n47719), .B(n47720), .Z(n47490) );
  AND U47510 ( .A(n1660), .B(n47721), .Z(n47720) );
  XOR U47511 ( .A(n47722), .B(n47723), .Z(n47713) );
  AND U47512 ( .A(n47724), .B(n47725), .Z(n47723) );
  XNOR U47513 ( .A(n47722), .B(n47541), .Z(n47725) );
  XOR U47514 ( .A(n47652), .B(n47726), .Z(n47541) );
  AND U47515 ( .A(n1644), .B(n47727), .Z(n47726) );
  XOR U47516 ( .A(n47648), .B(n47652), .Z(n47727) );
  XNOR U47517 ( .A(n47728), .B(n47722), .Z(n47724) );
  IV U47518 ( .A(n47500), .Z(n47728) );
  XOR U47519 ( .A(n47729), .B(n47730), .Z(n47500) );
  AND U47520 ( .A(n1660), .B(n47731), .Z(n47730) );
  AND U47521 ( .A(n47693), .B(n47682), .Z(n47722) );
  XNOR U47522 ( .A(n47732), .B(n47733), .Z(n47682) );
  AND U47523 ( .A(n1644), .B(n47664), .Z(n47733) );
  XNOR U47524 ( .A(n47662), .B(n47732), .Z(n47664) );
  XNOR U47525 ( .A(n47734), .B(n47735), .Z(n1644) );
  AND U47526 ( .A(n47736), .B(n47737), .Z(n47735) );
  XNOR U47527 ( .A(n47734), .B(n47553), .Z(n47737) );
  IV U47528 ( .A(n47557), .Z(n47553) );
  XOR U47529 ( .A(n47738), .B(n47739), .Z(n47557) );
  AND U47530 ( .A(n1648), .B(n47740), .Z(n47739) );
  XOR U47531 ( .A(n47741), .B(n47738), .Z(n47740) );
  XNOR U47532 ( .A(n47734), .B(n47669), .Z(n47736) );
  XOR U47533 ( .A(n47742), .B(n47743), .Z(n47669) );
  AND U47534 ( .A(n1656), .B(n47704), .Z(n47743) );
  XOR U47535 ( .A(n47702), .B(n47742), .Z(n47704) );
  XOR U47536 ( .A(n47744), .B(n47745), .Z(n47734) );
  AND U47537 ( .A(n47746), .B(n47747), .Z(n47745) );
  XNOR U47538 ( .A(n47744), .B(n47569), .Z(n47747) );
  IV U47539 ( .A(n47572), .Z(n47569) );
  XOR U47540 ( .A(n47748), .B(n47749), .Z(n47572) );
  AND U47541 ( .A(n1648), .B(n47750), .Z(n47749) );
  XOR U47542 ( .A(n47751), .B(n47748), .Z(n47750) );
  XOR U47543 ( .A(n47573), .B(n47744), .Z(n47746) );
  XOR U47544 ( .A(n47752), .B(n47753), .Z(n47573) );
  AND U47545 ( .A(n1656), .B(n47712), .Z(n47753) );
  XOR U47546 ( .A(n47752), .B(n47710), .Z(n47712) );
  XOR U47547 ( .A(n47754), .B(n47755), .Z(n47744) );
  AND U47548 ( .A(n47756), .B(n47757), .Z(n47755) );
  XNOR U47549 ( .A(n47754), .B(n47597), .Z(n47757) );
  IV U47550 ( .A(n47600), .Z(n47597) );
  XOR U47551 ( .A(n47758), .B(n47759), .Z(n47600) );
  AND U47552 ( .A(n1648), .B(n47760), .Z(n47759) );
  XNOR U47553 ( .A(n47761), .B(n47758), .Z(n47760) );
  XOR U47554 ( .A(n47601), .B(n47754), .Z(n47756) );
  XOR U47555 ( .A(n47762), .B(n47763), .Z(n47601) );
  AND U47556 ( .A(n1656), .B(n47721), .Z(n47763) );
  XOR U47557 ( .A(n47762), .B(n47719), .Z(n47721) );
  XOR U47558 ( .A(n47678), .B(n47764), .Z(n47754) );
  AND U47559 ( .A(n47680), .B(n47765), .Z(n47764) );
  XNOR U47560 ( .A(n47678), .B(n47648), .Z(n47765) );
  IV U47561 ( .A(n47651), .Z(n47648) );
  XOR U47562 ( .A(n47766), .B(n47767), .Z(n47651) );
  AND U47563 ( .A(n1648), .B(n47768), .Z(n47767) );
  XOR U47564 ( .A(n47769), .B(n47766), .Z(n47768) );
  XOR U47565 ( .A(n47652), .B(n47678), .Z(n47680) );
  XOR U47566 ( .A(n47770), .B(n47771), .Z(n47652) );
  AND U47567 ( .A(n1656), .B(n47731), .Z(n47771) );
  XOR U47568 ( .A(n47770), .B(n47729), .Z(n47731) );
  AND U47569 ( .A(n47732), .B(n47662), .Z(n47678) );
  XNOR U47570 ( .A(n47772), .B(n47773), .Z(n47662) );
  AND U47571 ( .A(n1648), .B(n47774), .Z(n47773) );
  XNOR U47572 ( .A(n47775), .B(n47772), .Z(n47774) );
  XNOR U47573 ( .A(n47776), .B(n47777), .Z(n1648) );
  AND U47574 ( .A(n47778), .B(n47779), .Z(n47777) );
  XOR U47575 ( .A(n47741), .B(n47776), .Z(n47779) );
  AND U47576 ( .A(n47780), .B(n47781), .Z(n47741) );
  XNOR U47577 ( .A(n47738), .B(n47776), .Z(n47778) );
  XNOR U47578 ( .A(n47782), .B(n47783), .Z(n47738) );
  AND U47579 ( .A(n1652), .B(n47784), .Z(n47783) );
  XNOR U47580 ( .A(n47785), .B(n47786), .Z(n47784) );
  XOR U47581 ( .A(n47787), .B(n47788), .Z(n47776) );
  AND U47582 ( .A(n47789), .B(n47790), .Z(n47788) );
  XNOR U47583 ( .A(n47787), .B(n47780), .Z(n47790) );
  IV U47584 ( .A(n47751), .Z(n47780) );
  XOR U47585 ( .A(n47791), .B(n47792), .Z(n47751) );
  XOR U47586 ( .A(n47793), .B(n47781), .Z(n47792) );
  AND U47587 ( .A(n47761), .B(n47794), .Z(n47781) );
  AND U47588 ( .A(n47795), .B(n47796), .Z(n47793) );
  XOR U47589 ( .A(n47797), .B(n47791), .Z(n47795) );
  XNOR U47590 ( .A(n47748), .B(n47787), .Z(n47789) );
  XNOR U47591 ( .A(n47798), .B(n47799), .Z(n47748) );
  AND U47592 ( .A(n1652), .B(n47800), .Z(n47799) );
  XNOR U47593 ( .A(n47801), .B(n47802), .Z(n47800) );
  XOR U47594 ( .A(n47803), .B(n47804), .Z(n47787) );
  AND U47595 ( .A(n47805), .B(n47806), .Z(n47804) );
  XNOR U47596 ( .A(n47803), .B(n47761), .Z(n47806) );
  XOR U47597 ( .A(n47807), .B(n47796), .Z(n47761) );
  XNOR U47598 ( .A(n47808), .B(n47791), .Z(n47796) );
  XOR U47599 ( .A(n47809), .B(n47810), .Z(n47791) );
  AND U47600 ( .A(n47811), .B(n47812), .Z(n47810) );
  XOR U47601 ( .A(n47813), .B(n47809), .Z(n47811) );
  XNOR U47602 ( .A(n47814), .B(n47815), .Z(n47808) );
  AND U47603 ( .A(n47816), .B(n47817), .Z(n47815) );
  XOR U47604 ( .A(n47814), .B(n47818), .Z(n47816) );
  XNOR U47605 ( .A(n47797), .B(n47794), .Z(n47807) );
  AND U47606 ( .A(n47819), .B(n47820), .Z(n47794) );
  XOR U47607 ( .A(n47821), .B(n47822), .Z(n47797) );
  AND U47608 ( .A(n47823), .B(n47824), .Z(n47822) );
  XOR U47609 ( .A(n47821), .B(n47825), .Z(n47823) );
  XNOR U47610 ( .A(n47758), .B(n47803), .Z(n47805) );
  XNOR U47611 ( .A(n47826), .B(n47827), .Z(n47758) );
  AND U47612 ( .A(n1652), .B(n47828), .Z(n47827) );
  XNOR U47613 ( .A(n47829), .B(n47830), .Z(n47828) );
  XOR U47614 ( .A(n47831), .B(n47832), .Z(n47803) );
  AND U47615 ( .A(n47833), .B(n47834), .Z(n47832) );
  XNOR U47616 ( .A(n47831), .B(n47819), .Z(n47834) );
  IV U47617 ( .A(n47769), .Z(n47819) );
  XNOR U47618 ( .A(n47835), .B(n47812), .Z(n47769) );
  XNOR U47619 ( .A(n47836), .B(n47818), .Z(n47812) );
  XNOR U47620 ( .A(n47837), .B(n47838), .Z(n47818) );
  NOR U47621 ( .A(n47839), .B(n47840), .Z(n47838) );
  XOR U47622 ( .A(n47837), .B(n47841), .Z(n47839) );
  XNOR U47623 ( .A(n47817), .B(n47809), .Z(n47836) );
  XOR U47624 ( .A(n47842), .B(n47843), .Z(n47809) );
  AND U47625 ( .A(n47844), .B(n47845), .Z(n47843) );
  XOR U47626 ( .A(n47842), .B(n47846), .Z(n47844) );
  XNOR U47627 ( .A(n47847), .B(n47814), .Z(n47817) );
  XOR U47628 ( .A(n47848), .B(n47849), .Z(n47814) );
  AND U47629 ( .A(n47850), .B(n47851), .Z(n47849) );
  XNOR U47630 ( .A(n47852), .B(n47853), .Z(n47850) );
  IV U47631 ( .A(n47848), .Z(n47852) );
  XNOR U47632 ( .A(n47854), .B(n47855), .Z(n47847) );
  NOR U47633 ( .A(n47856), .B(n47857), .Z(n47855) );
  XNOR U47634 ( .A(n47854), .B(n47858), .Z(n47856) );
  XNOR U47635 ( .A(n47813), .B(n47820), .Z(n47835) );
  NOR U47636 ( .A(n47775), .B(n47859), .Z(n47820) );
  XOR U47637 ( .A(n47825), .B(n47824), .Z(n47813) );
  XNOR U47638 ( .A(n47860), .B(n47821), .Z(n47824) );
  XOR U47639 ( .A(n47861), .B(n47862), .Z(n47821) );
  AND U47640 ( .A(n47863), .B(n47864), .Z(n47862) );
  XNOR U47641 ( .A(n47865), .B(n47866), .Z(n47863) );
  IV U47642 ( .A(n47861), .Z(n47865) );
  XNOR U47643 ( .A(n47867), .B(n47868), .Z(n47860) );
  NOR U47644 ( .A(n47869), .B(n47870), .Z(n47868) );
  XNOR U47645 ( .A(n47867), .B(n47871), .Z(n47869) );
  XOR U47646 ( .A(n47872), .B(n47873), .Z(n47825) );
  NOR U47647 ( .A(n47874), .B(n47875), .Z(n47873) );
  XNOR U47648 ( .A(n47872), .B(n47876), .Z(n47874) );
  XNOR U47649 ( .A(n47766), .B(n47831), .Z(n47833) );
  XNOR U47650 ( .A(n47877), .B(n47878), .Z(n47766) );
  AND U47651 ( .A(n1652), .B(n47879), .Z(n47878) );
  XNOR U47652 ( .A(n47880), .B(n47881), .Z(n47879) );
  AND U47653 ( .A(n47772), .B(n47775), .Z(n47831) );
  XOR U47654 ( .A(n47882), .B(n47859), .Z(n47775) );
  XNOR U47655 ( .A(p_input[1328]), .B(p_input[2048]), .Z(n47859) );
  XNOR U47656 ( .A(n47846), .B(n47845), .Z(n47882) );
  XNOR U47657 ( .A(n47883), .B(n47853), .Z(n47845) );
  XNOR U47658 ( .A(n47841), .B(n47840), .Z(n47853) );
  XNOR U47659 ( .A(n47884), .B(n47837), .Z(n47840) );
  XNOR U47660 ( .A(p_input[1338]), .B(p_input[2058]), .Z(n47837) );
  XOR U47661 ( .A(p_input[1339]), .B(n29030), .Z(n47884) );
  XOR U47662 ( .A(p_input[1340]), .B(p_input[2060]), .Z(n47841) );
  XOR U47663 ( .A(n47851), .B(n47885), .Z(n47883) );
  IV U47664 ( .A(n47842), .Z(n47885) );
  XOR U47665 ( .A(p_input[1329]), .B(p_input[2049]), .Z(n47842) );
  XNOR U47666 ( .A(n47886), .B(n47858), .Z(n47851) );
  XNOR U47667 ( .A(p_input[1343]), .B(n29033), .Z(n47858) );
  XOR U47668 ( .A(n47848), .B(n47857), .Z(n47886) );
  XOR U47669 ( .A(n47887), .B(n47854), .Z(n47857) );
  XOR U47670 ( .A(p_input[1341]), .B(p_input[2061]), .Z(n47854) );
  XOR U47671 ( .A(p_input[1342]), .B(n29035), .Z(n47887) );
  XOR U47672 ( .A(p_input[1337]), .B(p_input[2057]), .Z(n47848) );
  XOR U47673 ( .A(n47866), .B(n47864), .Z(n47846) );
  XNOR U47674 ( .A(n47888), .B(n47871), .Z(n47864) );
  XOR U47675 ( .A(p_input[1336]), .B(p_input[2056]), .Z(n47871) );
  XOR U47676 ( .A(n47861), .B(n47870), .Z(n47888) );
  XOR U47677 ( .A(n47889), .B(n47867), .Z(n47870) );
  XOR U47678 ( .A(p_input[1334]), .B(p_input[2054]), .Z(n47867) );
  XOR U47679 ( .A(p_input[1335]), .B(n30404), .Z(n47889) );
  XOR U47680 ( .A(p_input[1330]), .B(p_input[2050]), .Z(n47861) );
  XNOR U47681 ( .A(n47876), .B(n47875), .Z(n47866) );
  XOR U47682 ( .A(n47890), .B(n47872), .Z(n47875) );
  XOR U47683 ( .A(p_input[1331]), .B(p_input[2051]), .Z(n47872) );
  XOR U47684 ( .A(p_input[1332]), .B(n30406), .Z(n47890) );
  XOR U47685 ( .A(p_input[1333]), .B(p_input[2053]), .Z(n47876) );
  XNOR U47686 ( .A(n47891), .B(n47892), .Z(n47772) );
  AND U47687 ( .A(n1652), .B(n47893), .Z(n47892) );
  XNOR U47688 ( .A(n47894), .B(n47895), .Z(n1652) );
  AND U47689 ( .A(n47896), .B(n47897), .Z(n47895) );
  XOR U47690 ( .A(n47786), .B(n47894), .Z(n47897) );
  XNOR U47691 ( .A(n47898), .B(n47894), .Z(n47896) );
  XOR U47692 ( .A(n47899), .B(n47900), .Z(n47894) );
  AND U47693 ( .A(n47901), .B(n47902), .Z(n47900) );
  XOR U47694 ( .A(n47801), .B(n47899), .Z(n47902) );
  XOR U47695 ( .A(n47899), .B(n47802), .Z(n47901) );
  XOR U47696 ( .A(n47903), .B(n47904), .Z(n47899) );
  AND U47697 ( .A(n47905), .B(n47906), .Z(n47904) );
  XOR U47698 ( .A(n47829), .B(n47903), .Z(n47906) );
  XOR U47699 ( .A(n47903), .B(n47830), .Z(n47905) );
  XOR U47700 ( .A(n47907), .B(n47908), .Z(n47903) );
  AND U47701 ( .A(n47909), .B(n47910), .Z(n47908) );
  XOR U47702 ( .A(n47907), .B(n47880), .Z(n47910) );
  XNOR U47703 ( .A(n47911), .B(n47912), .Z(n47732) );
  AND U47704 ( .A(n1656), .B(n47913), .Z(n47912) );
  XNOR U47705 ( .A(n47914), .B(n47915), .Z(n1656) );
  AND U47706 ( .A(n47916), .B(n47917), .Z(n47915) );
  XOR U47707 ( .A(n47914), .B(n47742), .Z(n47917) );
  XNOR U47708 ( .A(n47914), .B(n47702), .Z(n47916) );
  XOR U47709 ( .A(n47918), .B(n47919), .Z(n47914) );
  AND U47710 ( .A(n47920), .B(n47921), .Z(n47919) );
  XOR U47711 ( .A(n47918), .B(n47710), .Z(n47920) );
  XOR U47712 ( .A(n47922), .B(n47923), .Z(n47693) );
  AND U47713 ( .A(n1660), .B(n47913), .Z(n47923) );
  XNOR U47714 ( .A(n47911), .B(n47922), .Z(n47913) );
  XNOR U47715 ( .A(n47924), .B(n47925), .Z(n1660) );
  AND U47716 ( .A(n47926), .B(n47927), .Z(n47925) );
  XNOR U47717 ( .A(n47928), .B(n47924), .Z(n47927) );
  IV U47718 ( .A(n47742), .Z(n47928) );
  XOR U47719 ( .A(n47898), .B(n47929), .Z(n47742) );
  AND U47720 ( .A(n1663), .B(n47930), .Z(n47929) );
  XOR U47721 ( .A(n47785), .B(n47782), .Z(n47930) );
  IV U47722 ( .A(n47898), .Z(n47785) );
  XNOR U47723 ( .A(n47702), .B(n47924), .Z(n47926) );
  XOR U47724 ( .A(n47931), .B(n47932), .Z(n47702) );
  AND U47725 ( .A(n1679), .B(n47933), .Z(n47932) );
  XOR U47726 ( .A(n47918), .B(n47934), .Z(n47924) );
  AND U47727 ( .A(n47935), .B(n47921), .Z(n47934) );
  XNOR U47728 ( .A(n47752), .B(n47918), .Z(n47921) );
  XOR U47729 ( .A(n47802), .B(n47936), .Z(n47752) );
  AND U47730 ( .A(n1663), .B(n47937), .Z(n47936) );
  XOR U47731 ( .A(n47798), .B(n47802), .Z(n47937) );
  XNOR U47732 ( .A(n47938), .B(n47918), .Z(n47935) );
  IV U47733 ( .A(n47710), .Z(n47938) );
  XOR U47734 ( .A(n47939), .B(n47940), .Z(n47710) );
  AND U47735 ( .A(n1679), .B(n47941), .Z(n47940) );
  XOR U47736 ( .A(n47942), .B(n47943), .Z(n47918) );
  AND U47737 ( .A(n47944), .B(n47945), .Z(n47943) );
  XNOR U47738 ( .A(n47762), .B(n47942), .Z(n47945) );
  XOR U47739 ( .A(n47830), .B(n47946), .Z(n47762) );
  AND U47740 ( .A(n1663), .B(n47947), .Z(n47946) );
  XOR U47741 ( .A(n47826), .B(n47830), .Z(n47947) );
  XOR U47742 ( .A(n47942), .B(n47719), .Z(n47944) );
  XOR U47743 ( .A(n47948), .B(n47949), .Z(n47719) );
  AND U47744 ( .A(n1679), .B(n47950), .Z(n47949) );
  XOR U47745 ( .A(n47951), .B(n47952), .Z(n47942) );
  AND U47746 ( .A(n47953), .B(n47954), .Z(n47952) );
  XNOR U47747 ( .A(n47951), .B(n47770), .Z(n47954) );
  XOR U47748 ( .A(n47881), .B(n47955), .Z(n47770) );
  AND U47749 ( .A(n1663), .B(n47956), .Z(n47955) );
  XOR U47750 ( .A(n47877), .B(n47881), .Z(n47956) );
  XNOR U47751 ( .A(n47957), .B(n47951), .Z(n47953) );
  IV U47752 ( .A(n47729), .Z(n47957) );
  XOR U47753 ( .A(n47958), .B(n47959), .Z(n47729) );
  AND U47754 ( .A(n1679), .B(n47960), .Z(n47959) );
  AND U47755 ( .A(n47922), .B(n47911), .Z(n47951) );
  XNOR U47756 ( .A(n47961), .B(n47962), .Z(n47911) );
  AND U47757 ( .A(n1663), .B(n47893), .Z(n47962) );
  XNOR U47758 ( .A(n47891), .B(n47961), .Z(n47893) );
  XNOR U47759 ( .A(n47963), .B(n47964), .Z(n1663) );
  AND U47760 ( .A(n47965), .B(n47966), .Z(n47964) );
  XNOR U47761 ( .A(n47963), .B(n47782), .Z(n47966) );
  IV U47762 ( .A(n47786), .Z(n47782) );
  XOR U47763 ( .A(n47967), .B(n47968), .Z(n47786) );
  AND U47764 ( .A(n1667), .B(n47969), .Z(n47968) );
  XOR U47765 ( .A(n47970), .B(n47967), .Z(n47969) );
  XNOR U47766 ( .A(n47963), .B(n47898), .Z(n47965) );
  XOR U47767 ( .A(n47971), .B(n47972), .Z(n47898) );
  AND U47768 ( .A(n1675), .B(n47933), .Z(n47972) );
  XOR U47769 ( .A(n47931), .B(n47971), .Z(n47933) );
  XOR U47770 ( .A(n47973), .B(n47974), .Z(n47963) );
  AND U47771 ( .A(n47975), .B(n47976), .Z(n47974) );
  XNOR U47772 ( .A(n47973), .B(n47798), .Z(n47976) );
  IV U47773 ( .A(n47801), .Z(n47798) );
  XOR U47774 ( .A(n47977), .B(n47978), .Z(n47801) );
  AND U47775 ( .A(n1667), .B(n47979), .Z(n47978) );
  XOR U47776 ( .A(n47980), .B(n47977), .Z(n47979) );
  XOR U47777 ( .A(n47802), .B(n47973), .Z(n47975) );
  XOR U47778 ( .A(n47981), .B(n47982), .Z(n47802) );
  AND U47779 ( .A(n1675), .B(n47941), .Z(n47982) );
  XOR U47780 ( .A(n47981), .B(n47939), .Z(n47941) );
  XOR U47781 ( .A(n47983), .B(n47984), .Z(n47973) );
  AND U47782 ( .A(n47985), .B(n47986), .Z(n47984) );
  XNOR U47783 ( .A(n47983), .B(n47826), .Z(n47986) );
  IV U47784 ( .A(n47829), .Z(n47826) );
  XOR U47785 ( .A(n47987), .B(n47988), .Z(n47829) );
  AND U47786 ( .A(n1667), .B(n47989), .Z(n47988) );
  XNOR U47787 ( .A(n47990), .B(n47987), .Z(n47989) );
  XOR U47788 ( .A(n47830), .B(n47983), .Z(n47985) );
  XOR U47789 ( .A(n47991), .B(n47992), .Z(n47830) );
  AND U47790 ( .A(n1675), .B(n47950), .Z(n47992) );
  XOR U47791 ( .A(n47991), .B(n47948), .Z(n47950) );
  XOR U47792 ( .A(n47907), .B(n47993), .Z(n47983) );
  AND U47793 ( .A(n47909), .B(n47994), .Z(n47993) );
  XNOR U47794 ( .A(n47907), .B(n47877), .Z(n47994) );
  IV U47795 ( .A(n47880), .Z(n47877) );
  XOR U47796 ( .A(n47995), .B(n47996), .Z(n47880) );
  AND U47797 ( .A(n1667), .B(n47997), .Z(n47996) );
  XOR U47798 ( .A(n47998), .B(n47995), .Z(n47997) );
  XOR U47799 ( .A(n47881), .B(n47907), .Z(n47909) );
  XOR U47800 ( .A(n47999), .B(n48000), .Z(n47881) );
  AND U47801 ( .A(n1675), .B(n47960), .Z(n48000) );
  XOR U47802 ( .A(n47999), .B(n47958), .Z(n47960) );
  AND U47803 ( .A(n47961), .B(n47891), .Z(n47907) );
  XNOR U47804 ( .A(n48001), .B(n48002), .Z(n47891) );
  AND U47805 ( .A(n1667), .B(n48003), .Z(n48002) );
  XNOR U47806 ( .A(n48004), .B(n48001), .Z(n48003) );
  XNOR U47807 ( .A(n48005), .B(n48006), .Z(n1667) );
  AND U47808 ( .A(n48007), .B(n48008), .Z(n48006) );
  XOR U47809 ( .A(n47970), .B(n48005), .Z(n48008) );
  AND U47810 ( .A(n48009), .B(n48010), .Z(n47970) );
  XNOR U47811 ( .A(n47967), .B(n48005), .Z(n48007) );
  XNOR U47812 ( .A(n48011), .B(n48012), .Z(n47967) );
  AND U47813 ( .A(n1671), .B(n48013), .Z(n48012) );
  XNOR U47814 ( .A(n48014), .B(n48015), .Z(n48013) );
  XOR U47815 ( .A(n48016), .B(n48017), .Z(n48005) );
  AND U47816 ( .A(n48018), .B(n48019), .Z(n48017) );
  XNOR U47817 ( .A(n48016), .B(n48009), .Z(n48019) );
  IV U47818 ( .A(n47980), .Z(n48009) );
  XOR U47819 ( .A(n48020), .B(n48021), .Z(n47980) );
  XOR U47820 ( .A(n48022), .B(n48010), .Z(n48021) );
  AND U47821 ( .A(n47990), .B(n48023), .Z(n48010) );
  AND U47822 ( .A(n48024), .B(n48025), .Z(n48022) );
  XOR U47823 ( .A(n48026), .B(n48020), .Z(n48024) );
  XNOR U47824 ( .A(n47977), .B(n48016), .Z(n48018) );
  XNOR U47825 ( .A(n48027), .B(n48028), .Z(n47977) );
  AND U47826 ( .A(n1671), .B(n48029), .Z(n48028) );
  XNOR U47827 ( .A(n48030), .B(n48031), .Z(n48029) );
  XOR U47828 ( .A(n48032), .B(n48033), .Z(n48016) );
  AND U47829 ( .A(n48034), .B(n48035), .Z(n48033) );
  XNOR U47830 ( .A(n48032), .B(n47990), .Z(n48035) );
  XOR U47831 ( .A(n48036), .B(n48025), .Z(n47990) );
  XNOR U47832 ( .A(n48037), .B(n48020), .Z(n48025) );
  XOR U47833 ( .A(n48038), .B(n48039), .Z(n48020) );
  AND U47834 ( .A(n48040), .B(n48041), .Z(n48039) );
  XOR U47835 ( .A(n48042), .B(n48038), .Z(n48040) );
  XNOR U47836 ( .A(n48043), .B(n48044), .Z(n48037) );
  AND U47837 ( .A(n48045), .B(n48046), .Z(n48044) );
  XOR U47838 ( .A(n48043), .B(n48047), .Z(n48045) );
  XNOR U47839 ( .A(n48026), .B(n48023), .Z(n48036) );
  AND U47840 ( .A(n48048), .B(n48049), .Z(n48023) );
  XOR U47841 ( .A(n48050), .B(n48051), .Z(n48026) );
  AND U47842 ( .A(n48052), .B(n48053), .Z(n48051) );
  XOR U47843 ( .A(n48050), .B(n48054), .Z(n48052) );
  XNOR U47844 ( .A(n47987), .B(n48032), .Z(n48034) );
  XNOR U47845 ( .A(n48055), .B(n48056), .Z(n47987) );
  AND U47846 ( .A(n1671), .B(n48057), .Z(n48056) );
  XNOR U47847 ( .A(n48058), .B(n48059), .Z(n48057) );
  XOR U47848 ( .A(n48060), .B(n48061), .Z(n48032) );
  AND U47849 ( .A(n48062), .B(n48063), .Z(n48061) );
  XNOR U47850 ( .A(n48060), .B(n48048), .Z(n48063) );
  IV U47851 ( .A(n47998), .Z(n48048) );
  XNOR U47852 ( .A(n48064), .B(n48041), .Z(n47998) );
  XNOR U47853 ( .A(n48065), .B(n48047), .Z(n48041) );
  XNOR U47854 ( .A(n48066), .B(n48067), .Z(n48047) );
  NOR U47855 ( .A(n48068), .B(n48069), .Z(n48067) );
  XOR U47856 ( .A(n48066), .B(n48070), .Z(n48068) );
  XNOR U47857 ( .A(n48046), .B(n48038), .Z(n48065) );
  XOR U47858 ( .A(n48071), .B(n48072), .Z(n48038) );
  AND U47859 ( .A(n48073), .B(n48074), .Z(n48072) );
  XOR U47860 ( .A(n48071), .B(n48075), .Z(n48073) );
  XNOR U47861 ( .A(n48076), .B(n48043), .Z(n48046) );
  XOR U47862 ( .A(n48077), .B(n48078), .Z(n48043) );
  AND U47863 ( .A(n48079), .B(n48080), .Z(n48078) );
  XNOR U47864 ( .A(n48081), .B(n48082), .Z(n48079) );
  IV U47865 ( .A(n48077), .Z(n48081) );
  XNOR U47866 ( .A(n48083), .B(n48084), .Z(n48076) );
  NOR U47867 ( .A(n48085), .B(n48086), .Z(n48084) );
  XNOR U47868 ( .A(n48083), .B(n48087), .Z(n48085) );
  XNOR U47869 ( .A(n48042), .B(n48049), .Z(n48064) );
  NOR U47870 ( .A(n48004), .B(n48088), .Z(n48049) );
  XOR U47871 ( .A(n48054), .B(n48053), .Z(n48042) );
  XNOR U47872 ( .A(n48089), .B(n48050), .Z(n48053) );
  XOR U47873 ( .A(n48090), .B(n48091), .Z(n48050) );
  AND U47874 ( .A(n48092), .B(n48093), .Z(n48091) );
  XNOR U47875 ( .A(n48094), .B(n48095), .Z(n48092) );
  IV U47876 ( .A(n48090), .Z(n48094) );
  XNOR U47877 ( .A(n48096), .B(n48097), .Z(n48089) );
  NOR U47878 ( .A(n48098), .B(n48099), .Z(n48097) );
  XNOR U47879 ( .A(n48096), .B(n48100), .Z(n48098) );
  XOR U47880 ( .A(n48101), .B(n48102), .Z(n48054) );
  NOR U47881 ( .A(n48103), .B(n48104), .Z(n48102) );
  XNOR U47882 ( .A(n48101), .B(n48105), .Z(n48103) );
  XNOR U47883 ( .A(n47995), .B(n48060), .Z(n48062) );
  XNOR U47884 ( .A(n48106), .B(n48107), .Z(n47995) );
  AND U47885 ( .A(n1671), .B(n48108), .Z(n48107) );
  XNOR U47886 ( .A(n48109), .B(n48110), .Z(n48108) );
  AND U47887 ( .A(n48001), .B(n48004), .Z(n48060) );
  XOR U47888 ( .A(n48111), .B(n48088), .Z(n48004) );
  XNOR U47889 ( .A(p_input[1344]), .B(p_input[2048]), .Z(n48088) );
  XNOR U47890 ( .A(n48075), .B(n48074), .Z(n48111) );
  XNOR U47891 ( .A(n48112), .B(n48082), .Z(n48074) );
  XNOR U47892 ( .A(n48070), .B(n48069), .Z(n48082) );
  XNOR U47893 ( .A(n48113), .B(n48066), .Z(n48069) );
  XNOR U47894 ( .A(p_input[1354]), .B(p_input[2058]), .Z(n48066) );
  XOR U47895 ( .A(p_input[1355]), .B(n29030), .Z(n48113) );
  XOR U47896 ( .A(p_input[1356]), .B(p_input[2060]), .Z(n48070) );
  XOR U47897 ( .A(n48080), .B(n48114), .Z(n48112) );
  IV U47898 ( .A(n48071), .Z(n48114) );
  XOR U47899 ( .A(p_input[1345]), .B(p_input[2049]), .Z(n48071) );
  XNOR U47900 ( .A(n48115), .B(n48087), .Z(n48080) );
  XNOR U47901 ( .A(p_input[1359]), .B(n29033), .Z(n48087) );
  XOR U47902 ( .A(n48077), .B(n48086), .Z(n48115) );
  XOR U47903 ( .A(n48116), .B(n48083), .Z(n48086) );
  XOR U47904 ( .A(p_input[1357]), .B(p_input[2061]), .Z(n48083) );
  XOR U47905 ( .A(p_input[1358]), .B(n29035), .Z(n48116) );
  XOR U47906 ( .A(p_input[1353]), .B(p_input[2057]), .Z(n48077) );
  XOR U47907 ( .A(n48095), .B(n48093), .Z(n48075) );
  XNOR U47908 ( .A(n48117), .B(n48100), .Z(n48093) );
  XOR U47909 ( .A(p_input[1352]), .B(p_input[2056]), .Z(n48100) );
  XOR U47910 ( .A(n48090), .B(n48099), .Z(n48117) );
  XOR U47911 ( .A(n48118), .B(n48096), .Z(n48099) );
  XOR U47912 ( .A(p_input[1350]), .B(p_input[2054]), .Z(n48096) );
  XOR U47913 ( .A(p_input[1351]), .B(n30404), .Z(n48118) );
  XOR U47914 ( .A(p_input[1346]), .B(p_input[2050]), .Z(n48090) );
  XNOR U47915 ( .A(n48105), .B(n48104), .Z(n48095) );
  XOR U47916 ( .A(n48119), .B(n48101), .Z(n48104) );
  XOR U47917 ( .A(p_input[1347]), .B(p_input[2051]), .Z(n48101) );
  XOR U47918 ( .A(p_input[1348]), .B(n30406), .Z(n48119) );
  XOR U47919 ( .A(p_input[1349]), .B(p_input[2053]), .Z(n48105) );
  XNOR U47920 ( .A(n48120), .B(n48121), .Z(n48001) );
  AND U47921 ( .A(n1671), .B(n48122), .Z(n48121) );
  XNOR U47922 ( .A(n48123), .B(n48124), .Z(n1671) );
  AND U47923 ( .A(n48125), .B(n48126), .Z(n48124) );
  XOR U47924 ( .A(n48015), .B(n48123), .Z(n48126) );
  XNOR U47925 ( .A(n48127), .B(n48123), .Z(n48125) );
  XOR U47926 ( .A(n48128), .B(n48129), .Z(n48123) );
  AND U47927 ( .A(n48130), .B(n48131), .Z(n48129) );
  XOR U47928 ( .A(n48030), .B(n48128), .Z(n48131) );
  XOR U47929 ( .A(n48128), .B(n48031), .Z(n48130) );
  XOR U47930 ( .A(n48132), .B(n48133), .Z(n48128) );
  AND U47931 ( .A(n48134), .B(n48135), .Z(n48133) );
  XOR U47932 ( .A(n48058), .B(n48132), .Z(n48135) );
  XOR U47933 ( .A(n48132), .B(n48059), .Z(n48134) );
  XOR U47934 ( .A(n48136), .B(n48137), .Z(n48132) );
  AND U47935 ( .A(n48138), .B(n48139), .Z(n48137) );
  XOR U47936 ( .A(n48136), .B(n48109), .Z(n48139) );
  XNOR U47937 ( .A(n48140), .B(n48141), .Z(n47961) );
  AND U47938 ( .A(n1675), .B(n48142), .Z(n48141) );
  XNOR U47939 ( .A(n48143), .B(n48144), .Z(n1675) );
  AND U47940 ( .A(n48145), .B(n48146), .Z(n48144) );
  XOR U47941 ( .A(n48143), .B(n47971), .Z(n48146) );
  XNOR U47942 ( .A(n48143), .B(n47931), .Z(n48145) );
  XOR U47943 ( .A(n48147), .B(n48148), .Z(n48143) );
  AND U47944 ( .A(n48149), .B(n48150), .Z(n48148) );
  XOR U47945 ( .A(n48147), .B(n47939), .Z(n48149) );
  XOR U47946 ( .A(n48151), .B(n48152), .Z(n47922) );
  AND U47947 ( .A(n1679), .B(n48142), .Z(n48152) );
  XNOR U47948 ( .A(n48140), .B(n48151), .Z(n48142) );
  XNOR U47949 ( .A(n48153), .B(n48154), .Z(n1679) );
  AND U47950 ( .A(n48155), .B(n48156), .Z(n48154) );
  XNOR U47951 ( .A(n48157), .B(n48153), .Z(n48156) );
  IV U47952 ( .A(n47971), .Z(n48157) );
  XOR U47953 ( .A(n48127), .B(n48158), .Z(n47971) );
  AND U47954 ( .A(n1682), .B(n48159), .Z(n48158) );
  XOR U47955 ( .A(n48014), .B(n48011), .Z(n48159) );
  IV U47956 ( .A(n48127), .Z(n48014) );
  XNOR U47957 ( .A(n47931), .B(n48153), .Z(n48155) );
  XOR U47958 ( .A(n48160), .B(n48161), .Z(n47931) );
  AND U47959 ( .A(n1698), .B(n48162), .Z(n48161) );
  XOR U47960 ( .A(n48147), .B(n48163), .Z(n48153) );
  AND U47961 ( .A(n48164), .B(n48150), .Z(n48163) );
  XNOR U47962 ( .A(n47981), .B(n48147), .Z(n48150) );
  XOR U47963 ( .A(n48031), .B(n48165), .Z(n47981) );
  AND U47964 ( .A(n1682), .B(n48166), .Z(n48165) );
  XOR U47965 ( .A(n48027), .B(n48031), .Z(n48166) );
  XNOR U47966 ( .A(n48167), .B(n48147), .Z(n48164) );
  IV U47967 ( .A(n47939), .Z(n48167) );
  XOR U47968 ( .A(n48168), .B(n48169), .Z(n47939) );
  AND U47969 ( .A(n1698), .B(n48170), .Z(n48169) );
  XOR U47970 ( .A(n48171), .B(n48172), .Z(n48147) );
  AND U47971 ( .A(n48173), .B(n48174), .Z(n48172) );
  XNOR U47972 ( .A(n47991), .B(n48171), .Z(n48174) );
  XOR U47973 ( .A(n48059), .B(n48175), .Z(n47991) );
  AND U47974 ( .A(n1682), .B(n48176), .Z(n48175) );
  XOR U47975 ( .A(n48055), .B(n48059), .Z(n48176) );
  XOR U47976 ( .A(n48171), .B(n47948), .Z(n48173) );
  XOR U47977 ( .A(n48177), .B(n48178), .Z(n47948) );
  AND U47978 ( .A(n1698), .B(n48179), .Z(n48178) );
  XOR U47979 ( .A(n48180), .B(n48181), .Z(n48171) );
  AND U47980 ( .A(n48182), .B(n48183), .Z(n48181) );
  XNOR U47981 ( .A(n48180), .B(n47999), .Z(n48183) );
  XOR U47982 ( .A(n48110), .B(n48184), .Z(n47999) );
  AND U47983 ( .A(n1682), .B(n48185), .Z(n48184) );
  XOR U47984 ( .A(n48106), .B(n48110), .Z(n48185) );
  XNOR U47985 ( .A(n48186), .B(n48180), .Z(n48182) );
  IV U47986 ( .A(n47958), .Z(n48186) );
  XOR U47987 ( .A(n48187), .B(n48188), .Z(n47958) );
  AND U47988 ( .A(n1698), .B(n48189), .Z(n48188) );
  AND U47989 ( .A(n48151), .B(n48140), .Z(n48180) );
  XNOR U47990 ( .A(n48190), .B(n48191), .Z(n48140) );
  AND U47991 ( .A(n1682), .B(n48122), .Z(n48191) );
  XNOR U47992 ( .A(n48120), .B(n48190), .Z(n48122) );
  XNOR U47993 ( .A(n48192), .B(n48193), .Z(n1682) );
  AND U47994 ( .A(n48194), .B(n48195), .Z(n48193) );
  XNOR U47995 ( .A(n48192), .B(n48011), .Z(n48195) );
  IV U47996 ( .A(n48015), .Z(n48011) );
  XOR U47997 ( .A(n48196), .B(n48197), .Z(n48015) );
  AND U47998 ( .A(n1686), .B(n48198), .Z(n48197) );
  XOR U47999 ( .A(n48199), .B(n48196), .Z(n48198) );
  XNOR U48000 ( .A(n48192), .B(n48127), .Z(n48194) );
  XOR U48001 ( .A(n48200), .B(n48201), .Z(n48127) );
  AND U48002 ( .A(n1694), .B(n48162), .Z(n48201) );
  XOR U48003 ( .A(n48160), .B(n48200), .Z(n48162) );
  XOR U48004 ( .A(n48202), .B(n48203), .Z(n48192) );
  AND U48005 ( .A(n48204), .B(n48205), .Z(n48203) );
  XNOR U48006 ( .A(n48202), .B(n48027), .Z(n48205) );
  IV U48007 ( .A(n48030), .Z(n48027) );
  XOR U48008 ( .A(n48206), .B(n48207), .Z(n48030) );
  AND U48009 ( .A(n1686), .B(n48208), .Z(n48207) );
  XOR U48010 ( .A(n48209), .B(n48206), .Z(n48208) );
  XOR U48011 ( .A(n48031), .B(n48202), .Z(n48204) );
  XOR U48012 ( .A(n48210), .B(n48211), .Z(n48031) );
  AND U48013 ( .A(n1694), .B(n48170), .Z(n48211) );
  XOR U48014 ( .A(n48210), .B(n48168), .Z(n48170) );
  XOR U48015 ( .A(n48212), .B(n48213), .Z(n48202) );
  AND U48016 ( .A(n48214), .B(n48215), .Z(n48213) );
  XNOR U48017 ( .A(n48212), .B(n48055), .Z(n48215) );
  IV U48018 ( .A(n48058), .Z(n48055) );
  XOR U48019 ( .A(n48216), .B(n48217), .Z(n48058) );
  AND U48020 ( .A(n1686), .B(n48218), .Z(n48217) );
  XNOR U48021 ( .A(n48219), .B(n48216), .Z(n48218) );
  XOR U48022 ( .A(n48059), .B(n48212), .Z(n48214) );
  XOR U48023 ( .A(n48220), .B(n48221), .Z(n48059) );
  AND U48024 ( .A(n1694), .B(n48179), .Z(n48221) );
  XOR U48025 ( .A(n48220), .B(n48177), .Z(n48179) );
  XOR U48026 ( .A(n48136), .B(n48222), .Z(n48212) );
  AND U48027 ( .A(n48138), .B(n48223), .Z(n48222) );
  XNOR U48028 ( .A(n48136), .B(n48106), .Z(n48223) );
  IV U48029 ( .A(n48109), .Z(n48106) );
  XOR U48030 ( .A(n48224), .B(n48225), .Z(n48109) );
  AND U48031 ( .A(n1686), .B(n48226), .Z(n48225) );
  XOR U48032 ( .A(n48227), .B(n48224), .Z(n48226) );
  XOR U48033 ( .A(n48110), .B(n48136), .Z(n48138) );
  XOR U48034 ( .A(n48228), .B(n48229), .Z(n48110) );
  AND U48035 ( .A(n1694), .B(n48189), .Z(n48229) );
  XOR U48036 ( .A(n48228), .B(n48187), .Z(n48189) );
  AND U48037 ( .A(n48190), .B(n48120), .Z(n48136) );
  XNOR U48038 ( .A(n48230), .B(n48231), .Z(n48120) );
  AND U48039 ( .A(n1686), .B(n48232), .Z(n48231) );
  XNOR U48040 ( .A(n48233), .B(n48230), .Z(n48232) );
  XNOR U48041 ( .A(n48234), .B(n48235), .Z(n1686) );
  AND U48042 ( .A(n48236), .B(n48237), .Z(n48235) );
  XOR U48043 ( .A(n48199), .B(n48234), .Z(n48237) );
  AND U48044 ( .A(n48238), .B(n48239), .Z(n48199) );
  XNOR U48045 ( .A(n48196), .B(n48234), .Z(n48236) );
  XNOR U48046 ( .A(n48240), .B(n48241), .Z(n48196) );
  AND U48047 ( .A(n1690), .B(n48242), .Z(n48241) );
  XNOR U48048 ( .A(n48243), .B(n48244), .Z(n48242) );
  XOR U48049 ( .A(n48245), .B(n48246), .Z(n48234) );
  AND U48050 ( .A(n48247), .B(n48248), .Z(n48246) );
  XNOR U48051 ( .A(n48245), .B(n48238), .Z(n48248) );
  IV U48052 ( .A(n48209), .Z(n48238) );
  XOR U48053 ( .A(n48249), .B(n48250), .Z(n48209) );
  XOR U48054 ( .A(n48251), .B(n48239), .Z(n48250) );
  AND U48055 ( .A(n48219), .B(n48252), .Z(n48239) );
  AND U48056 ( .A(n48253), .B(n48254), .Z(n48251) );
  XOR U48057 ( .A(n48255), .B(n48249), .Z(n48253) );
  XNOR U48058 ( .A(n48206), .B(n48245), .Z(n48247) );
  XNOR U48059 ( .A(n48256), .B(n48257), .Z(n48206) );
  AND U48060 ( .A(n1690), .B(n48258), .Z(n48257) );
  XNOR U48061 ( .A(n48259), .B(n48260), .Z(n48258) );
  XOR U48062 ( .A(n48261), .B(n48262), .Z(n48245) );
  AND U48063 ( .A(n48263), .B(n48264), .Z(n48262) );
  XNOR U48064 ( .A(n48261), .B(n48219), .Z(n48264) );
  XOR U48065 ( .A(n48265), .B(n48254), .Z(n48219) );
  XNOR U48066 ( .A(n48266), .B(n48249), .Z(n48254) );
  XOR U48067 ( .A(n48267), .B(n48268), .Z(n48249) );
  AND U48068 ( .A(n48269), .B(n48270), .Z(n48268) );
  XOR U48069 ( .A(n48271), .B(n48267), .Z(n48269) );
  XNOR U48070 ( .A(n48272), .B(n48273), .Z(n48266) );
  AND U48071 ( .A(n48274), .B(n48275), .Z(n48273) );
  XOR U48072 ( .A(n48272), .B(n48276), .Z(n48274) );
  XNOR U48073 ( .A(n48255), .B(n48252), .Z(n48265) );
  AND U48074 ( .A(n48277), .B(n48278), .Z(n48252) );
  XOR U48075 ( .A(n48279), .B(n48280), .Z(n48255) );
  AND U48076 ( .A(n48281), .B(n48282), .Z(n48280) );
  XOR U48077 ( .A(n48279), .B(n48283), .Z(n48281) );
  XNOR U48078 ( .A(n48216), .B(n48261), .Z(n48263) );
  XNOR U48079 ( .A(n48284), .B(n48285), .Z(n48216) );
  AND U48080 ( .A(n1690), .B(n48286), .Z(n48285) );
  XNOR U48081 ( .A(n48287), .B(n48288), .Z(n48286) );
  XOR U48082 ( .A(n48289), .B(n48290), .Z(n48261) );
  AND U48083 ( .A(n48291), .B(n48292), .Z(n48290) );
  XNOR U48084 ( .A(n48289), .B(n48277), .Z(n48292) );
  IV U48085 ( .A(n48227), .Z(n48277) );
  XNOR U48086 ( .A(n48293), .B(n48270), .Z(n48227) );
  XNOR U48087 ( .A(n48294), .B(n48276), .Z(n48270) );
  XNOR U48088 ( .A(n48295), .B(n48296), .Z(n48276) );
  NOR U48089 ( .A(n48297), .B(n48298), .Z(n48296) );
  XOR U48090 ( .A(n48295), .B(n48299), .Z(n48297) );
  XNOR U48091 ( .A(n48275), .B(n48267), .Z(n48294) );
  XOR U48092 ( .A(n48300), .B(n48301), .Z(n48267) );
  AND U48093 ( .A(n48302), .B(n48303), .Z(n48301) );
  XOR U48094 ( .A(n48300), .B(n48304), .Z(n48302) );
  XNOR U48095 ( .A(n48305), .B(n48272), .Z(n48275) );
  XOR U48096 ( .A(n48306), .B(n48307), .Z(n48272) );
  AND U48097 ( .A(n48308), .B(n48309), .Z(n48307) );
  XNOR U48098 ( .A(n48310), .B(n48311), .Z(n48308) );
  IV U48099 ( .A(n48306), .Z(n48310) );
  XNOR U48100 ( .A(n48312), .B(n48313), .Z(n48305) );
  NOR U48101 ( .A(n48314), .B(n48315), .Z(n48313) );
  XNOR U48102 ( .A(n48312), .B(n48316), .Z(n48314) );
  XNOR U48103 ( .A(n48271), .B(n48278), .Z(n48293) );
  NOR U48104 ( .A(n48233), .B(n48317), .Z(n48278) );
  XOR U48105 ( .A(n48283), .B(n48282), .Z(n48271) );
  XNOR U48106 ( .A(n48318), .B(n48279), .Z(n48282) );
  XOR U48107 ( .A(n48319), .B(n48320), .Z(n48279) );
  AND U48108 ( .A(n48321), .B(n48322), .Z(n48320) );
  XNOR U48109 ( .A(n48323), .B(n48324), .Z(n48321) );
  IV U48110 ( .A(n48319), .Z(n48323) );
  XNOR U48111 ( .A(n48325), .B(n48326), .Z(n48318) );
  NOR U48112 ( .A(n48327), .B(n48328), .Z(n48326) );
  XNOR U48113 ( .A(n48325), .B(n48329), .Z(n48327) );
  XOR U48114 ( .A(n48330), .B(n48331), .Z(n48283) );
  NOR U48115 ( .A(n48332), .B(n48333), .Z(n48331) );
  XNOR U48116 ( .A(n48330), .B(n48334), .Z(n48332) );
  XNOR U48117 ( .A(n48224), .B(n48289), .Z(n48291) );
  XNOR U48118 ( .A(n48335), .B(n48336), .Z(n48224) );
  AND U48119 ( .A(n1690), .B(n48337), .Z(n48336) );
  XNOR U48120 ( .A(n48338), .B(n48339), .Z(n48337) );
  AND U48121 ( .A(n48230), .B(n48233), .Z(n48289) );
  XOR U48122 ( .A(n48340), .B(n48317), .Z(n48233) );
  XNOR U48123 ( .A(p_input[1360]), .B(p_input[2048]), .Z(n48317) );
  XNOR U48124 ( .A(n48304), .B(n48303), .Z(n48340) );
  XNOR U48125 ( .A(n48341), .B(n48311), .Z(n48303) );
  XNOR U48126 ( .A(n48299), .B(n48298), .Z(n48311) );
  XNOR U48127 ( .A(n48342), .B(n48295), .Z(n48298) );
  XNOR U48128 ( .A(p_input[1370]), .B(p_input[2058]), .Z(n48295) );
  XOR U48129 ( .A(p_input[1371]), .B(n29030), .Z(n48342) );
  XOR U48130 ( .A(p_input[1372]), .B(p_input[2060]), .Z(n48299) );
  XOR U48131 ( .A(n48309), .B(n48343), .Z(n48341) );
  IV U48132 ( .A(n48300), .Z(n48343) );
  XOR U48133 ( .A(p_input[1361]), .B(p_input[2049]), .Z(n48300) );
  XNOR U48134 ( .A(n48344), .B(n48316), .Z(n48309) );
  XNOR U48135 ( .A(p_input[1375]), .B(n29033), .Z(n48316) );
  XOR U48136 ( .A(n48306), .B(n48315), .Z(n48344) );
  XOR U48137 ( .A(n48345), .B(n48312), .Z(n48315) );
  XOR U48138 ( .A(p_input[1373]), .B(p_input[2061]), .Z(n48312) );
  XOR U48139 ( .A(p_input[1374]), .B(n29035), .Z(n48345) );
  XOR U48140 ( .A(p_input[1369]), .B(p_input[2057]), .Z(n48306) );
  XOR U48141 ( .A(n48324), .B(n48322), .Z(n48304) );
  XNOR U48142 ( .A(n48346), .B(n48329), .Z(n48322) );
  XOR U48143 ( .A(p_input[1368]), .B(p_input[2056]), .Z(n48329) );
  XOR U48144 ( .A(n48319), .B(n48328), .Z(n48346) );
  XOR U48145 ( .A(n48347), .B(n48325), .Z(n48328) );
  XOR U48146 ( .A(p_input[1366]), .B(p_input[2054]), .Z(n48325) );
  XOR U48147 ( .A(p_input[1367]), .B(n30404), .Z(n48347) );
  XOR U48148 ( .A(p_input[1362]), .B(p_input[2050]), .Z(n48319) );
  XNOR U48149 ( .A(n48334), .B(n48333), .Z(n48324) );
  XOR U48150 ( .A(n48348), .B(n48330), .Z(n48333) );
  XOR U48151 ( .A(p_input[1363]), .B(p_input[2051]), .Z(n48330) );
  XOR U48152 ( .A(p_input[1364]), .B(n30406), .Z(n48348) );
  XOR U48153 ( .A(p_input[1365]), .B(p_input[2053]), .Z(n48334) );
  XNOR U48154 ( .A(n48349), .B(n48350), .Z(n48230) );
  AND U48155 ( .A(n1690), .B(n48351), .Z(n48350) );
  XNOR U48156 ( .A(n48352), .B(n48353), .Z(n1690) );
  AND U48157 ( .A(n48354), .B(n48355), .Z(n48353) );
  XOR U48158 ( .A(n48244), .B(n48352), .Z(n48355) );
  XNOR U48159 ( .A(n48356), .B(n48352), .Z(n48354) );
  XOR U48160 ( .A(n48357), .B(n48358), .Z(n48352) );
  AND U48161 ( .A(n48359), .B(n48360), .Z(n48358) );
  XOR U48162 ( .A(n48259), .B(n48357), .Z(n48360) );
  XOR U48163 ( .A(n48357), .B(n48260), .Z(n48359) );
  XOR U48164 ( .A(n48361), .B(n48362), .Z(n48357) );
  AND U48165 ( .A(n48363), .B(n48364), .Z(n48362) );
  XOR U48166 ( .A(n48287), .B(n48361), .Z(n48364) );
  XOR U48167 ( .A(n48361), .B(n48288), .Z(n48363) );
  XOR U48168 ( .A(n48365), .B(n48366), .Z(n48361) );
  AND U48169 ( .A(n48367), .B(n48368), .Z(n48366) );
  XOR U48170 ( .A(n48365), .B(n48338), .Z(n48368) );
  XNOR U48171 ( .A(n48369), .B(n48370), .Z(n48190) );
  AND U48172 ( .A(n1694), .B(n48371), .Z(n48370) );
  XNOR U48173 ( .A(n48372), .B(n48373), .Z(n1694) );
  AND U48174 ( .A(n48374), .B(n48375), .Z(n48373) );
  XOR U48175 ( .A(n48372), .B(n48200), .Z(n48375) );
  XNOR U48176 ( .A(n48372), .B(n48160), .Z(n48374) );
  XOR U48177 ( .A(n48376), .B(n48377), .Z(n48372) );
  AND U48178 ( .A(n48378), .B(n48379), .Z(n48377) );
  XOR U48179 ( .A(n48376), .B(n48168), .Z(n48378) );
  XOR U48180 ( .A(n48380), .B(n48381), .Z(n48151) );
  AND U48181 ( .A(n1698), .B(n48371), .Z(n48381) );
  XNOR U48182 ( .A(n48369), .B(n48380), .Z(n48371) );
  XNOR U48183 ( .A(n48382), .B(n48383), .Z(n1698) );
  AND U48184 ( .A(n48384), .B(n48385), .Z(n48383) );
  XNOR U48185 ( .A(n48386), .B(n48382), .Z(n48385) );
  IV U48186 ( .A(n48200), .Z(n48386) );
  XOR U48187 ( .A(n48356), .B(n48387), .Z(n48200) );
  AND U48188 ( .A(n1701), .B(n48388), .Z(n48387) );
  XOR U48189 ( .A(n48243), .B(n48240), .Z(n48388) );
  IV U48190 ( .A(n48356), .Z(n48243) );
  XNOR U48191 ( .A(n48160), .B(n48382), .Z(n48384) );
  XOR U48192 ( .A(n48389), .B(n48390), .Z(n48160) );
  AND U48193 ( .A(n1717), .B(n48391), .Z(n48390) );
  XOR U48194 ( .A(n48376), .B(n48392), .Z(n48382) );
  AND U48195 ( .A(n48393), .B(n48379), .Z(n48392) );
  XNOR U48196 ( .A(n48210), .B(n48376), .Z(n48379) );
  XOR U48197 ( .A(n48260), .B(n48394), .Z(n48210) );
  AND U48198 ( .A(n1701), .B(n48395), .Z(n48394) );
  XOR U48199 ( .A(n48256), .B(n48260), .Z(n48395) );
  XNOR U48200 ( .A(n48396), .B(n48376), .Z(n48393) );
  IV U48201 ( .A(n48168), .Z(n48396) );
  XOR U48202 ( .A(n48397), .B(n48398), .Z(n48168) );
  AND U48203 ( .A(n1717), .B(n48399), .Z(n48398) );
  XOR U48204 ( .A(n48400), .B(n48401), .Z(n48376) );
  AND U48205 ( .A(n48402), .B(n48403), .Z(n48401) );
  XNOR U48206 ( .A(n48220), .B(n48400), .Z(n48403) );
  XOR U48207 ( .A(n48288), .B(n48404), .Z(n48220) );
  AND U48208 ( .A(n1701), .B(n48405), .Z(n48404) );
  XOR U48209 ( .A(n48284), .B(n48288), .Z(n48405) );
  XOR U48210 ( .A(n48400), .B(n48177), .Z(n48402) );
  XOR U48211 ( .A(n48406), .B(n48407), .Z(n48177) );
  AND U48212 ( .A(n1717), .B(n48408), .Z(n48407) );
  XOR U48213 ( .A(n48409), .B(n48410), .Z(n48400) );
  AND U48214 ( .A(n48411), .B(n48412), .Z(n48410) );
  XNOR U48215 ( .A(n48409), .B(n48228), .Z(n48412) );
  XOR U48216 ( .A(n48339), .B(n48413), .Z(n48228) );
  AND U48217 ( .A(n1701), .B(n48414), .Z(n48413) );
  XOR U48218 ( .A(n48335), .B(n48339), .Z(n48414) );
  XNOR U48219 ( .A(n48415), .B(n48409), .Z(n48411) );
  IV U48220 ( .A(n48187), .Z(n48415) );
  XOR U48221 ( .A(n48416), .B(n48417), .Z(n48187) );
  AND U48222 ( .A(n1717), .B(n48418), .Z(n48417) );
  AND U48223 ( .A(n48380), .B(n48369), .Z(n48409) );
  XNOR U48224 ( .A(n48419), .B(n48420), .Z(n48369) );
  AND U48225 ( .A(n1701), .B(n48351), .Z(n48420) );
  XNOR U48226 ( .A(n48349), .B(n48419), .Z(n48351) );
  XNOR U48227 ( .A(n48421), .B(n48422), .Z(n1701) );
  AND U48228 ( .A(n48423), .B(n48424), .Z(n48422) );
  XNOR U48229 ( .A(n48421), .B(n48240), .Z(n48424) );
  IV U48230 ( .A(n48244), .Z(n48240) );
  XOR U48231 ( .A(n48425), .B(n48426), .Z(n48244) );
  AND U48232 ( .A(n1705), .B(n48427), .Z(n48426) );
  XOR U48233 ( .A(n48428), .B(n48425), .Z(n48427) );
  XNOR U48234 ( .A(n48421), .B(n48356), .Z(n48423) );
  XOR U48235 ( .A(n48429), .B(n48430), .Z(n48356) );
  AND U48236 ( .A(n1713), .B(n48391), .Z(n48430) );
  XOR U48237 ( .A(n48389), .B(n48429), .Z(n48391) );
  XOR U48238 ( .A(n48431), .B(n48432), .Z(n48421) );
  AND U48239 ( .A(n48433), .B(n48434), .Z(n48432) );
  XNOR U48240 ( .A(n48431), .B(n48256), .Z(n48434) );
  IV U48241 ( .A(n48259), .Z(n48256) );
  XOR U48242 ( .A(n48435), .B(n48436), .Z(n48259) );
  AND U48243 ( .A(n1705), .B(n48437), .Z(n48436) );
  XOR U48244 ( .A(n48438), .B(n48435), .Z(n48437) );
  XOR U48245 ( .A(n48260), .B(n48431), .Z(n48433) );
  XOR U48246 ( .A(n48439), .B(n48440), .Z(n48260) );
  AND U48247 ( .A(n1713), .B(n48399), .Z(n48440) );
  XOR U48248 ( .A(n48439), .B(n48397), .Z(n48399) );
  XOR U48249 ( .A(n48441), .B(n48442), .Z(n48431) );
  AND U48250 ( .A(n48443), .B(n48444), .Z(n48442) );
  XNOR U48251 ( .A(n48441), .B(n48284), .Z(n48444) );
  IV U48252 ( .A(n48287), .Z(n48284) );
  XOR U48253 ( .A(n48445), .B(n48446), .Z(n48287) );
  AND U48254 ( .A(n1705), .B(n48447), .Z(n48446) );
  XNOR U48255 ( .A(n48448), .B(n48445), .Z(n48447) );
  XOR U48256 ( .A(n48288), .B(n48441), .Z(n48443) );
  XOR U48257 ( .A(n48449), .B(n48450), .Z(n48288) );
  AND U48258 ( .A(n1713), .B(n48408), .Z(n48450) );
  XOR U48259 ( .A(n48449), .B(n48406), .Z(n48408) );
  XOR U48260 ( .A(n48365), .B(n48451), .Z(n48441) );
  AND U48261 ( .A(n48367), .B(n48452), .Z(n48451) );
  XNOR U48262 ( .A(n48365), .B(n48335), .Z(n48452) );
  IV U48263 ( .A(n48338), .Z(n48335) );
  XOR U48264 ( .A(n48453), .B(n48454), .Z(n48338) );
  AND U48265 ( .A(n1705), .B(n48455), .Z(n48454) );
  XOR U48266 ( .A(n48456), .B(n48453), .Z(n48455) );
  XOR U48267 ( .A(n48339), .B(n48365), .Z(n48367) );
  XOR U48268 ( .A(n48457), .B(n48458), .Z(n48339) );
  AND U48269 ( .A(n1713), .B(n48418), .Z(n48458) );
  XOR U48270 ( .A(n48457), .B(n48416), .Z(n48418) );
  AND U48271 ( .A(n48419), .B(n48349), .Z(n48365) );
  XNOR U48272 ( .A(n48459), .B(n48460), .Z(n48349) );
  AND U48273 ( .A(n1705), .B(n48461), .Z(n48460) );
  XNOR U48274 ( .A(n48462), .B(n48459), .Z(n48461) );
  XNOR U48275 ( .A(n48463), .B(n48464), .Z(n1705) );
  AND U48276 ( .A(n48465), .B(n48466), .Z(n48464) );
  XOR U48277 ( .A(n48428), .B(n48463), .Z(n48466) );
  AND U48278 ( .A(n48467), .B(n48468), .Z(n48428) );
  XNOR U48279 ( .A(n48425), .B(n48463), .Z(n48465) );
  XNOR U48280 ( .A(n48469), .B(n48470), .Z(n48425) );
  AND U48281 ( .A(n1709), .B(n48471), .Z(n48470) );
  XNOR U48282 ( .A(n48472), .B(n48473), .Z(n48471) );
  XOR U48283 ( .A(n48474), .B(n48475), .Z(n48463) );
  AND U48284 ( .A(n48476), .B(n48477), .Z(n48475) );
  XNOR U48285 ( .A(n48474), .B(n48467), .Z(n48477) );
  IV U48286 ( .A(n48438), .Z(n48467) );
  XOR U48287 ( .A(n48478), .B(n48479), .Z(n48438) );
  XOR U48288 ( .A(n48480), .B(n48468), .Z(n48479) );
  AND U48289 ( .A(n48448), .B(n48481), .Z(n48468) );
  AND U48290 ( .A(n48482), .B(n48483), .Z(n48480) );
  XOR U48291 ( .A(n48484), .B(n48478), .Z(n48482) );
  XNOR U48292 ( .A(n48435), .B(n48474), .Z(n48476) );
  XNOR U48293 ( .A(n48485), .B(n48486), .Z(n48435) );
  AND U48294 ( .A(n1709), .B(n48487), .Z(n48486) );
  XNOR U48295 ( .A(n48488), .B(n48489), .Z(n48487) );
  XOR U48296 ( .A(n48490), .B(n48491), .Z(n48474) );
  AND U48297 ( .A(n48492), .B(n48493), .Z(n48491) );
  XNOR U48298 ( .A(n48490), .B(n48448), .Z(n48493) );
  XOR U48299 ( .A(n48494), .B(n48483), .Z(n48448) );
  XNOR U48300 ( .A(n48495), .B(n48478), .Z(n48483) );
  XOR U48301 ( .A(n48496), .B(n48497), .Z(n48478) );
  AND U48302 ( .A(n48498), .B(n48499), .Z(n48497) );
  XOR U48303 ( .A(n48500), .B(n48496), .Z(n48498) );
  XNOR U48304 ( .A(n48501), .B(n48502), .Z(n48495) );
  AND U48305 ( .A(n48503), .B(n48504), .Z(n48502) );
  XOR U48306 ( .A(n48501), .B(n48505), .Z(n48503) );
  XNOR U48307 ( .A(n48484), .B(n48481), .Z(n48494) );
  AND U48308 ( .A(n48506), .B(n48507), .Z(n48481) );
  XOR U48309 ( .A(n48508), .B(n48509), .Z(n48484) );
  AND U48310 ( .A(n48510), .B(n48511), .Z(n48509) );
  XOR U48311 ( .A(n48508), .B(n48512), .Z(n48510) );
  XNOR U48312 ( .A(n48445), .B(n48490), .Z(n48492) );
  XNOR U48313 ( .A(n48513), .B(n48514), .Z(n48445) );
  AND U48314 ( .A(n1709), .B(n48515), .Z(n48514) );
  XNOR U48315 ( .A(n48516), .B(n48517), .Z(n48515) );
  XOR U48316 ( .A(n48518), .B(n48519), .Z(n48490) );
  AND U48317 ( .A(n48520), .B(n48521), .Z(n48519) );
  XNOR U48318 ( .A(n48518), .B(n48506), .Z(n48521) );
  IV U48319 ( .A(n48456), .Z(n48506) );
  XNOR U48320 ( .A(n48522), .B(n48499), .Z(n48456) );
  XNOR U48321 ( .A(n48523), .B(n48505), .Z(n48499) );
  XNOR U48322 ( .A(n48524), .B(n48525), .Z(n48505) );
  NOR U48323 ( .A(n48526), .B(n48527), .Z(n48525) );
  XOR U48324 ( .A(n48524), .B(n48528), .Z(n48526) );
  XNOR U48325 ( .A(n48504), .B(n48496), .Z(n48523) );
  XOR U48326 ( .A(n48529), .B(n48530), .Z(n48496) );
  AND U48327 ( .A(n48531), .B(n48532), .Z(n48530) );
  XOR U48328 ( .A(n48529), .B(n48533), .Z(n48531) );
  XNOR U48329 ( .A(n48534), .B(n48501), .Z(n48504) );
  XOR U48330 ( .A(n48535), .B(n48536), .Z(n48501) );
  AND U48331 ( .A(n48537), .B(n48538), .Z(n48536) );
  XNOR U48332 ( .A(n48539), .B(n48540), .Z(n48537) );
  IV U48333 ( .A(n48535), .Z(n48539) );
  XNOR U48334 ( .A(n48541), .B(n48542), .Z(n48534) );
  NOR U48335 ( .A(n48543), .B(n48544), .Z(n48542) );
  XNOR U48336 ( .A(n48541), .B(n48545), .Z(n48543) );
  XNOR U48337 ( .A(n48500), .B(n48507), .Z(n48522) );
  NOR U48338 ( .A(n48462), .B(n48546), .Z(n48507) );
  XOR U48339 ( .A(n48512), .B(n48511), .Z(n48500) );
  XNOR U48340 ( .A(n48547), .B(n48508), .Z(n48511) );
  XOR U48341 ( .A(n48548), .B(n48549), .Z(n48508) );
  AND U48342 ( .A(n48550), .B(n48551), .Z(n48549) );
  XNOR U48343 ( .A(n48552), .B(n48553), .Z(n48550) );
  IV U48344 ( .A(n48548), .Z(n48552) );
  XNOR U48345 ( .A(n48554), .B(n48555), .Z(n48547) );
  NOR U48346 ( .A(n48556), .B(n48557), .Z(n48555) );
  XNOR U48347 ( .A(n48554), .B(n48558), .Z(n48556) );
  XOR U48348 ( .A(n48559), .B(n48560), .Z(n48512) );
  NOR U48349 ( .A(n48561), .B(n48562), .Z(n48560) );
  XNOR U48350 ( .A(n48559), .B(n48563), .Z(n48561) );
  XNOR U48351 ( .A(n48453), .B(n48518), .Z(n48520) );
  XNOR U48352 ( .A(n48564), .B(n48565), .Z(n48453) );
  AND U48353 ( .A(n1709), .B(n48566), .Z(n48565) );
  XNOR U48354 ( .A(n48567), .B(n48568), .Z(n48566) );
  AND U48355 ( .A(n48459), .B(n48462), .Z(n48518) );
  XOR U48356 ( .A(n48569), .B(n48546), .Z(n48462) );
  XNOR U48357 ( .A(p_input[1376]), .B(p_input[2048]), .Z(n48546) );
  XNOR U48358 ( .A(n48533), .B(n48532), .Z(n48569) );
  XNOR U48359 ( .A(n48570), .B(n48540), .Z(n48532) );
  XNOR U48360 ( .A(n48528), .B(n48527), .Z(n48540) );
  XNOR U48361 ( .A(n48571), .B(n48524), .Z(n48527) );
  XNOR U48362 ( .A(p_input[1386]), .B(p_input[2058]), .Z(n48524) );
  XOR U48363 ( .A(p_input[1387]), .B(n29030), .Z(n48571) );
  XOR U48364 ( .A(p_input[1388]), .B(p_input[2060]), .Z(n48528) );
  XOR U48365 ( .A(n48538), .B(n48572), .Z(n48570) );
  IV U48366 ( .A(n48529), .Z(n48572) );
  XOR U48367 ( .A(p_input[1377]), .B(p_input[2049]), .Z(n48529) );
  XNOR U48368 ( .A(n48573), .B(n48545), .Z(n48538) );
  XNOR U48369 ( .A(p_input[1391]), .B(n29033), .Z(n48545) );
  XOR U48370 ( .A(n48535), .B(n48544), .Z(n48573) );
  XOR U48371 ( .A(n48574), .B(n48541), .Z(n48544) );
  XOR U48372 ( .A(p_input[1389]), .B(p_input[2061]), .Z(n48541) );
  XOR U48373 ( .A(p_input[1390]), .B(n29035), .Z(n48574) );
  XOR U48374 ( .A(p_input[1385]), .B(p_input[2057]), .Z(n48535) );
  XOR U48375 ( .A(n48553), .B(n48551), .Z(n48533) );
  XNOR U48376 ( .A(n48575), .B(n48558), .Z(n48551) );
  XOR U48377 ( .A(p_input[1384]), .B(p_input[2056]), .Z(n48558) );
  XOR U48378 ( .A(n48548), .B(n48557), .Z(n48575) );
  XOR U48379 ( .A(n48576), .B(n48554), .Z(n48557) );
  XOR U48380 ( .A(p_input[1382]), .B(p_input[2054]), .Z(n48554) );
  XOR U48381 ( .A(p_input[1383]), .B(n30404), .Z(n48576) );
  XOR U48382 ( .A(p_input[1378]), .B(p_input[2050]), .Z(n48548) );
  XNOR U48383 ( .A(n48563), .B(n48562), .Z(n48553) );
  XOR U48384 ( .A(n48577), .B(n48559), .Z(n48562) );
  XOR U48385 ( .A(p_input[1379]), .B(p_input[2051]), .Z(n48559) );
  XOR U48386 ( .A(p_input[1380]), .B(n30406), .Z(n48577) );
  XOR U48387 ( .A(p_input[1381]), .B(p_input[2053]), .Z(n48563) );
  XNOR U48388 ( .A(n48578), .B(n48579), .Z(n48459) );
  AND U48389 ( .A(n1709), .B(n48580), .Z(n48579) );
  XNOR U48390 ( .A(n48581), .B(n48582), .Z(n1709) );
  AND U48391 ( .A(n48583), .B(n48584), .Z(n48582) );
  XOR U48392 ( .A(n48473), .B(n48581), .Z(n48584) );
  XNOR U48393 ( .A(n48585), .B(n48581), .Z(n48583) );
  XOR U48394 ( .A(n48586), .B(n48587), .Z(n48581) );
  AND U48395 ( .A(n48588), .B(n48589), .Z(n48587) );
  XOR U48396 ( .A(n48488), .B(n48586), .Z(n48589) );
  XOR U48397 ( .A(n48586), .B(n48489), .Z(n48588) );
  XOR U48398 ( .A(n48590), .B(n48591), .Z(n48586) );
  AND U48399 ( .A(n48592), .B(n48593), .Z(n48591) );
  XOR U48400 ( .A(n48516), .B(n48590), .Z(n48593) );
  XOR U48401 ( .A(n48590), .B(n48517), .Z(n48592) );
  XOR U48402 ( .A(n48594), .B(n48595), .Z(n48590) );
  AND U48403 ( .A(n48596), .B(n48597), .Z(n48595) );
  XOR U48404 ( .A(n48594), .B(n48567), .Z(n48597) );
  XNOR U48405 ( .A(n48598), .B(n48599), .Z(n48419) );
  AND U48406 ( .A(n1713), .B(n48600), .Z(n48599) );
  XNOR U48407 ( .A(n48601), .B(n48602), .Z(n1713) );
  AND U48408 ( .A(n48603), .B(n48604), .Z(n48602) );
  XOR U48409 ( .A(n48601), .B(n48429), .Z(n48604) );
  XNOR U48410 ( .A(n48601), .B(n48389), .Z(n48603) );
  XOR U48411 ( .A(n48605), .B(n48606), .Z(n48601) );
  AND U48412 ( .A(n48607), .B(n48608), .Z(n48606) );
  XOR U48413 ( .A(n48605), .B(n48397), .Z(n48607) );
  XOR U48414 ( .A(n48609), .B(n48610), .Z(n48380) );
  AND U48415 ( .A(n1717), .B(n48600), .Z(n48610) );
  XNOR U48416 ( .A(n48598), .B(n48609), .Z(n48600) );
  XNOR U48417 ( .A(n48611), .B(n48612), .Z(n1717) );
  AND U48418 ( .A(n48613), .B(n48614), .Z(n48612) );
  XNOR U48419 ( .A(n48615), .B(n48611), .Z(n48614) );
  IV U48420 ( .A(n48429), .Z(n48615) );
  XOR U48421 ( .A(n48585), .B(n48616), .Z(n48429) );
  AND U48422 ( .A(n1720), .B(n48617), .Z(n48616) );
  XOR U48423 ( .A(n48472), .B(n48469), .Z(n48617) );
  IV U48424 ( .A(n48585), .Z(n48472) );
  XNOR U48425 ( .A(n48389), .B(n48611), .Z(n48613) );
  XOR U48426 ( .A(n48618), .B(n48619), .Z(n48389) );
  AND U48427 ( .A(n1736), .B(n48620), .Z(n48619) );
  XOR U48428 ( .A(n48605), .B(n48621), .Z(n48611) );
  AND U48429 ( .A(n48622), .B(n48608), .Z(n48621) );
  XNOR U48430 ( .A(n48439), .B(n48605), .Z(n48608) );
  XOR U48431 ( .A(n48489), .B(n48623), .Z(n48439) );
  AND U48432 ( .A(n1720), .B(n48624), .Z(n48623) );
  XOR U48433 ( .A(n48485), .B(n48489), .Z(n48624) );
  XNOR U48434 ( .A(n48625), .B(n48605), .Z(n48622) );
  IV U48435 ( .A(n48397), .Z(n48625) );
  XOR U48436 ( .A(n48626), .B(n48627), .Z(n48397) );
  AND U48437 ( .A(n1736), .B(n48628), .Z(n48627) );
  XOR U48438 ( .A(n48629), .B(n48630), .Z(n48605) );
  AND U48439 ( .A(n48631), .B(n48632), .Z(n48630) );
  XNOR U48440 ( .A(n48449), .B(n48629), .Z(n48632) );
  XOR U48441 ( .A(n48517), .B(n48633), .Z(n48449) );
  AND U48442 ( .A(n1720), .B(n48634), .Z(n48633) );
  XOR U48443 ( .A(n48513), .B(n48517), .Z(n48634) );
  XOR U48444 ( .A(n48629), .B(n48406), .Z(n48631) );
  XOR U48445 ( .A(n48635), .B(n48636), .Z(n48406) );
  AND U48446 ( .A(n1736), .B(n48637), .Z(n48636) );
  XOR U48447 ( .A(n48638), .B(n48639), .Z(n48629) );
  AND U48448 ( .A(n48640), .B(n48641), .Z(n48639) );
  XNOR U48449 ( .A(n48638), .B(n48457), .Z(n48641) );
  XOR U48450 ( .A(n48568), .B(n48642), .Z(n48457) );
  AND U48451 ( .A(n1720), .B(n48643), .Z(n48642) );
  XOR U48452 ( .A(n48564), .B(n48568), .Z(n48643) );
  XNOR U48453 ( .A(n48644), .B(n48638), .Z(n48640) );
  IV U48454 ( .A(n48416), .Z(n48644) );
  XOR U48455 ( .A(n48645), .B(n48646), .Z(n48416) );
  AND U48456 ( .A(n1736), .B(n48647), .Z(n48646) );
  AND U48457 ( .A(n48609), .B(n48598), .Z(n48638) );
  XNOR U48458 ( .A(n48648), .B(n48649), .Z(n48598) );
  AND U48459 ( .A(n1720), .B(n48580), .Z(n48649) );
  XNOR U48460 ( .A(n48578), .B(n48648), .Z(n48580) );
  XNOR U48461 ( .A(n48650), .B(n48651), .Z(n1720) );
  AND U48462 ( .A(n48652), .B(n48653), .Z(n48651) );
  XNOR U48463 ( .A(n48650), .B(n48469), .Z(n48653) );
  IV U48464 ( .A(n48473), .Z(n48469) );
  XOR U48465 ( .A(n48654), .B(n48655), .Z(n48473) );
  AND U48466 ( .A(n1724), .B(n48656), .Z(n48655) );
  XOR U48467 ( .A(n48657), .B(n48654), .Z(n48656) );
  XNOR U48468 ( .A(n48650), .B(n48585), .Z(n48652) );
  XOR U48469 ( .A(n48658), .B(n48659), .Z(n48585) );
  AND U48470 ( .A(n1732), .B(n48620), .Z(n48659) );
  XOR U48471 ( .A(n48618), .B(n48658), .Z(n48620) );
  XOR U48472 ( .A(n48660), .B(n48661), .Z(n48650) );
  AND U48473 ( .A(n48662), .B(n48663), .Z(n48661) );
  XNOR U48474 ( .A(n48660), .B(n48485), .Z(n48663) );
  IV U48475 ( .A(n48488), .Z(n48485) );
  XOR U48476 ( .A(n48664), .B(n48665), .Z(n48488) );
  AND U48477 ( .A(n1724), .B(n48666), .Z(n48665) );
  XOR U48478 ( .A(n48667), .B(n48664), .Z(n48666) );
  XOR U48479 ( .A(n48489), .B(n48660), .Z(n48662) );
  XOR U48480 ( .A(n48668), .B(n48669), .Z(n48489) );
  AND U48481 ( .A(n1732), .B(n48628), .Z(n48669) );
  XOR U48482 ( .A(n48668), .B(n48626), .Z(n48628) );
  XOR U48483 ( .A(n48670), .B(n48671), .Z(n48660) );
  AND U48484 ( .A(n48672), .B(n48673), .Z(n48671) );
  XNOR U48485 ( .A(n48670), .B(n48513), .Z(n48673) );
  IV U48486 ( .A(n48516), .Z(n48513) );
  XOR U48487 ( .A(n48674), .B(n48675), .Z(n48516) );
  AND U48488 ( .A(n1724), .B(n48676), .Z(n48675) );
  XNOR U48489 ( .A(n48677), .B(n48674), .Z(n48676) );
  XOR U48490 ( .A(n48517), .B(n48670), .Z(n48672) );
  XOR U48491 ( .A(n48678), .B(n48679), .Z(n48517) );
  AND U48492 ( .A(n1732), .B(n48637), .Z(n48679) );
  XOR U48493 ( .A(n48678), .B(n48635), .Z(n48637) );
  XOR U48494 ( .A(n48594), .B(n48680), .Z(n48670) );
  AND U48495 ( .A(n48596), .B(n48681), .Z(n48680) );
  XNOR U48496 ( .A(n48594), .B(n48564), .Z(n48681) );
  IV U48497 ( .A(n48567), .Z(n48564) );
  XOR U48498 ( .A(n48682), .B(n48683), .Z(n48567) );
  AND U48499 ( .A(n1724), .B(n48684), .Z(n48683) );
  XOR U48500 ( .A(n48685), .B(n48682), .Z(n48684) );
  XOR U48501 ( .A(n48568), .B(n48594), .Z(n48596) );
  XOR U48502 ( .A(n48686), .B(n48687), .Z(n48568) );
  AND U48503 ( .A(n1732), .B(n48647), .Z(n48687) );
  XOR U48504 ( .A(n48686), .B(n48645), .Z(n48647) );
  AND U48505 ( .A(n48648), .B(n48578), .Z(n48594) );
  XNOR U48506 ( .A(n48688), .B(n48689), .Z(n48578) );
  AND U48507 ( .A(n1724), .B(n48690), .Z(n48689) );
  XNOR U48508 ( .A(n48691), .B(n48688), .Z(n48690) );
  XNOR U48509 ( .A(n48692), .B(n48693), .Z(n1724) );
  AND U48510 ( .A(n48694), .B(n48695), .Z(n48693) );
  XOR U48511 ( .A(n48657), .B(n48692), .Z(n48695) );
  AND U48512 ( .A(n48696), .B(n48697), .Z(n48657) );
  XNOR U48513 ( .A(n48654), .B(n48692), .Z(n48694) );
  XNOR U48514 ( .A(n48698), .B(n48699), .Z(n48654) );
  AND U48515 ( .A(n1728), .B(n48700), .Z(n48699) );
  XNOR U48516 ( .A(n48701), .B(n48702), .Z(n48700) );
  XOR U48517 ( .A(n48703), .B(n48704), .Z(n48692) );
  AND U48518 ( .A(n48705), .B(n48706), .Z(n48704) );
  XNOR U48519 ( .A(n48703), .B(n48696), .Z(n48706) );
  IV U48520 ( .A(n48667), .Z(n48696) );
  XOR U48521 ( .A(n48707), .B(n48708), .Z(n48667) );
  XOR U48522 ( .A(n48709), .B(n48697), .Z(n48708) );
  AND U48523 ( .A(n48677), .B(n48710), .Z(n48697) );
  AND U48524 ( .A(n48711), .B(n48712), .Z(n48709) );
  XOR U48525 ( .A(n48713), .B(n48707), .Z(n48711) );
  XNOR U48526 ( .A(n48664), .B(n48703), .Z(n48705) );
  XNOR U48527 ( .A(n48714), .B(n48715), .Z(n48664) );
  AND U48528 ( .A(n1728), .B(n48716), .Z(n48715) );
  XNOR U48529 ( .A(n48717), .B(n48718), .Z(n48716) );
  XOR U48530 ( .A(n48719), .B(n48720), .Z(n48703) );
  AND U48531 ( .A(n48721), .B(n48722), .Z(n48720) );
  XNOR U48532 ( .A(n48719), .B(n48677), .Z(n48722) );
  XOR U48533 ( .A(n48723), .B(n48712), .Z(n48677) );
  XNOR U48534 ( .A(n48724), .B(n48707), .Z(n48712) );
  XOR U48535 ( .A(n48725), .B(n48726), .Z(n48707) );
  AND U48536 ( .A(n48727), .B(n48728), .Z(n48726) );
  XOR U48537 ( .A(n48729), .B(n48725), .Z(n48727) );
  XNOR U48538 ( .A(n48730), .B(n48731), .Z(n48724) );
  AND U48539 ( .A(n48732), .B(n48733), .Z(n48731) );
  XOR U48540 ( .A(n48730), .B(n48734), .Z(n48732) );
  XNOR U48541 ( .A(n48713), .B(n48710), .Z(n48723) );
  AND U48542 ( .A(n48735), .B(n48736), .Z(n48710) );
  XOR U48543 ( .A(n48737), .B(n48738), .Z(n48713) );
  AND U48544 ( .A(n48739), .B(n48740), .Z(n48738) );
  XOR U48545 ( .A(n48737), .B(n48741), .Z(n48739) );
  XNOR U48546 ( .A(n48674), .B(n48719), .Z(n48721) );
  XNOR U48547 ( .A(n48742), .B(n48743), .Z(n48674) );
  AND U48548 ( .A(n1728), .B(n48744), .Z(n48743) );
  XNOR U48549 ( .A(n48745), .B(n48746), .Z(n48744) );
  XOR U48550 ( .A(n48747), .B(n48748), .Z(n48719) );
  AND U48551 ( .A(n48749), .B(n48750), .Z(n48748) );
  XNOR U48552 ( .A(n48747), .B(n48735), .Z(n48750) );
  IV U48553 ( .A(n48685), .Z(n48735) );
  XNOR U48554 ( .A(n48751), .B(n48728), .Z(n48685) );
  XNOR U48555 ( .A(n48752), .B(n48734), .Z(n48728) );
  XNOR U48556 ( .A(n48753), .B(n48754), .Z(n48734) );
  NOR U48557 ( .A(n48755), .B(n48756), .Z(n48754) );
  XOR U48558 ( .A(n48753), .B(n48757), .Z(n48755) );
  XNOR U48559 ( .A(n48733), .B(n48725), .Z(n48752) );
  XOR U48560 ( .A(n48758), .B(n48759), .Z(n48725) );
  AND U48561 ( .A(n48760), .B(n48761), .Z(n48759) );
  XOR U48562 ( .A(n48758), .B(n48762), .Z(n48760) );
  XNOR U48563 ( .A(n48763), .B(n48730), .Z(n48733) );
  XOR U48564 ( .A(n48764), .B(n48765), .Z(n48730) );
  AND U48565 ( .A(n48766), .B(n48767), .Z(n48765) );
  XNOR U48566 ( .A(n48768), .B(n48769), .Z(n48766) );
  IV U48567 ( .A(n48764), .Z(n48768) );
  XNOR U48568 ( .A(n48770), .B(n48771), .Z(n48763) );
  NOR U48569 ( .A(n48772), .B(n48773), .Z(n48771) );
  XNOR U48570 ( .A(n48770), .B(n48774), .Z(n48772) );
  XNOR U48571 ( .A(n48729), .B(n48736), .Z(n48751) );
  NOR U48572 ( .A(n48691), .B(n48775), .Z(n48736) );
  XOR U48573 ( .A(n48741), .B(n48740), .Z(n48729) );
  XNOR U48574 ( .A(n48776), .B(n48737), .Z(n48740) );
  XOR U48575 ( .A(n48777), .B(n48778), .Z(n48737) );
  AND U48576 ( .A(n48779), .B(n48780), .Z(n48778) );
  XNOR U48577 ( .A(n48781), .B(n48782), .Z(n48779) );
  IV U48578 ( .A(n48777), .Z(n48781) );
  XNOR U48579 ( .A(n48783), .B(n48784), .Z(n48776) );
  NOR U48580 ( .A(n48785), .B(n48786), .Z(n48784) );
  XNOR U48581 ( .A(n48783), .B(n48787), .Z(n48785) );
  XOR U48582 ( .A(n48788), .B(n48789), .Z(n48741) );
  NOR U48583 ( .A(n48790), .B(n48791), .Z(n48789) );
  XNOR U48584 ( .A(n48788), .B(n48792), .Z(n48790) );
  XNOR U48585 ( .A(n48682), .B(n48747), .Z(n48749) );
  XNOR U48586 ( .A(n48793), .B(n48794), .Z(n48682) );
  AND U48587 ( .A(n1728), .B(n48795), .Z(n48794) );
  XNOR U48588 ( .A(n48796), .B(n48797), .Z(n48795) );
  AND U48589 ( .A(n48688), .B(n48691), .Z(n48747) );
  XOR U48590 ( .A(n48798), .B(n48775), .Z(n48691) );
  XNOR U48591 ( .A(p_input[1392]), .B(p_input[2048]), .Z(n48775) );
  XNOR U48592 ( .A(n48762), .B(n48761), .Z(n48798) );
  XNOR U48593 ( .A(n48799), .B(n48769), .Z(n48761) );
  XNOR U48594 ( .A(n48757), .B(n48756), .Z(n48769) );
  XNOR U48595 ( .A(n48800), .B(n48753), .Z(n48756) );
  XNOR U48596 ( .A(p_input[1402]), .B(p_input[2058]), .Z(n48753) );
  XOR U48597 ( .A(p_input[1403]), .B(n29030), .Z(n48800) );
  XOR U48598 ( .A(p_input[1404]), .B(p_input[2060]), .Z(n48757) );
  XOR U48599 ( .A(n48767), .B(n48801), .Z(n48799) );
  IV U48600 ( .A(n48758), .Z(n48801) );
  XOR U48601 ( .A(p_input[1393]), .B(p_input[2049]), .Z(n48758) );
  XNOR U48602 ( .A(n48802), .B(n48774), .Z(n48767) );
  XNOR U48603 ( .A(p_input[1407]), .B(n29033), .Z(n48774) );
  XOR U48604 ( .A(n48764), .B(n48773), .Z(n48802) );
  XOR U48605 ( .A(n48803), .B(n48770), .Z(n48773) );
  XOR U48606 ( .A(p_input[1405]), .B(p_input[2061]), .Z(n48770) );
  XOR U48607 ( .A(p_input[1406]), .B(n29035), .Z(n48803) );
  XOR U48608 ( .A(p_input[1401]), .B(p_input[2057]), .Z(n48764) );
  XOR U48609 ( .A(n48782), .B(n48780), .Z(n48762) );
  XNOR U48610 ( .A(n48804), .B(n48787), .Z(n48780) );
  XOR U48611 ( .A(p_input[1400]), .B(p_input[2056]), .Z(n48787) );
  XOR U48612 ( .A(n48777), .B(n48786), .Z(n48804) );
  XOR U48613 ( .A(n48805), .B(n48783), .Z(n48786) );
  XOR U48614 ( .A(p_input[1398]), .B(p_input[2054]), .Z(n48783) );
  XOR U48615 ( .A(p_input[1399]), .B(n30404), .Z(n48805) );
  XOR U48616 ( .A(p_input[1394]), .B(p_input[2050]), .Z(n48777) );
  XNOR U48617 ( .A(n48792), .B(n48791), .Z(n48782) );
  XOR U48618 ( .A(n48806), .B(n48788), .Z(n48791) );
  XOR U48619 ( .A(p_input[1395]), .B(p_input[2051]), .Z(n48788) );
  XOR U48620 ( .A(p_input[1396]), .B(n30406), .Z(n48806) );
  XOR U48621 ( .A(p_input[1397]), .B(p_input[2053]), .Z(n48792) );
  XNOR U48622 ( .A(n48807), .B(n48808), .Z(n48688) );
  AND U48623 ( .A(n1728), .B(n48809), .Z(n48808) );
  XNOR U48624 ( .A(n48810), .B(n48811), .Z(n1728) );
  AND U48625 ( .A(n48812), .B(n48813), .Z(n48811) );
  XOR U48626 ( .A(n48702), .B(n48810), .Z(n48813) );
  XNOR U48627 ( .A(n48814), .B(n48810), .Z(n48812) );
  XOR U48628 ( .A(n48815), .B(n48816), .Z(n48810) );
  AND U48629 ( .A(n48817), .B(n48818), .Z(n48816) );
  XOR U48630 ( .A(n48717), .B(n48815), .Z(n48818) );
  XOR U48631 ( .A(n48815), .B(n48718), .Z(n48817) );
  XOR U48632 ( .A(n48819), .B(n48820), .Z(n48815) );
  AND U48633 ( .A(n48821), .B(n48822), .Z(n48820) );
  XOR U48634 ( .A(n48745), .B(n48819), .Z(n48822) );
  XOR U48635 ( .A(n48819), .B(n48746), .Z(n48821) );
  XOR U48636 ( .A(n48823), .B(n48824), .Z(n48819) );
  AND U48637 ( .A(n48825), .B(n48826), .Z(n48824) );
  XOR U48638 ( .A(n48823), .B(n48796), .Z(n48826) );
  XNOR U48639 ( .A(n48827), .B(n48828), .Z(n48648) );
  AND U48640 ( .A(n1732), .B(n48829), .Z(n48828) );
  XNOR U48641 ( .A(n48830), .B(n48831), .Z(n1732) );
  AND U48642 ( .A(n48832), .B(n48833), .Z(n48831) );
  XOR U48643 ( .A(n48830), .B(n48658), .Z(n48833) );
  XNOR U48644 ( .A(n48830), .B(n48618), .Z(n48832) );
  XOR U48645 ( .A(n48834), .B(n48835), .Z(n48830) );
  AND U48646 ( .A(n48836), .B(n48837), .Z(n48835) );
  XOR U48647 ( .A(n48834), .B(n48626), .Z(n48836) );
  XOR U48648 ( .A(n48838), .B(n48839), .Z(n48609) );
  AND U48649 ( .A(n1736), .B(n48829), .Z(n48839) );
  XNOR U48650 ( .A(n48827), .B(n48838), .Z(n48829) );
  XNOR U48651 ( .A(n48840), .B(n48841), .Z(n1736) );
  AND U48652 ( .A(n48842), .B(n48843), .Z(n48841) );
  XNOR U48653 ( .A(n48844), .B(n48840), .Z(n48843) );
  IV U48654 ( .A(n48658), .Z(n48844) );
  XOR U48655 ( .A(n48814), .B(n48845), .Z(n48658) );
  AND U48656 ( .A(n1739), .B(n48846), .Z(n48845) );
  XOR U48657 ( .A(n48701), .B(n48698), .Z(n48846) );
  IV U48658 ( .A(n48814), .Z(n48701) );
  XNOR U48659 ( .A(n48618), .B(n48840), .Z(n48842) );
  XOR U48660 ( .A(n48847), .B(n48848), .Z(n48618) );
  AND U48661 ( .A(n1755), .B(n48849), .Z(n48848) );
  XOR U48662 ( .A(n48834), .B(n48850), .Z(n48840) );
  AND U48663 ( .A(n48851), .B(n48837), .Z(n48850) );
  XNOR U48664 ( .A(n48668), .B(n48834), .Z(n48837) );
  XOR U48665 ( .A(n48718), .B(n48852), .Z(n48668) );
  AND U48666 ( .A(n1739), .B(n48853), .Z(n48852) );
  XOR U48667 ( .A(n48714), .B(n48718), .Z(n48853) );
  XNOR U48668 ( .A(n48854), .B(n48834), .Z(n48851) );
  IV U48669 ( .A(n48626), .Z(n48854) );
  XOR U48670 ( .A(n48855), .B(n48856), .Z(n48626) );
  AND U48671 ( .A(n1755), .B(n48857), .Z(n48856) );
  XOR U48672 ( .A(n48858), .B(n48859), .Z(n48834) );
  AND U48673 ( .A(n48860), .B(n48861), .Z(n48859) );
  XNOR U48674 ( .A(n48678), .B(n48858), .Z(n48861) );
  XOR U48675 ( .A(n48746), .B(n48862), .Z(n48678) );
  AND U48676 ( .A(n1739), .B(n48863), .Z(n48862) );
  XOR U48677 ( .A(n48742), .B(n48746), .Z(n48863) );
  XOR U48678 ( .A(n48858), .B(n48635), .Z(n48860) );
  XOR U48679 ( .A(n48864), .B(n48865), .Z(n48635) );
  AND U48680 ( .A(n1755), .B(n48866), .Z(n48865) );
  XOR U48681 ( .A(n48867), .B(n48868), .Z(n48858) );
  AND U48682 ( .A(n48869), .B(n48870), .Z(n48868) );
  XNOR U48683 ( .A(n48867), .B(n48686), .Z(n48870) );
  XOR U48684 ( .A(n48797), .B(n48871), .Z(n48686) );
  AND U48685 ( .A(n1739), .B(n48872), .Z(n48871) );
  XOR U48686 ( .A(n48793), .B(n48797), .Z(n48872) );
  XNOR U48687 ( .A(n48873), .B(n48867), .Z(n48869) );
  IV U48688 ( .A(n48645), .Z(n48873) );
  XOR U48689 ( .A(n48874), .B(n48875), .Z(n48645) );
  AND U48690 ( .A(n1755), .B(n48876), .Z(n48875) );
  AND U48691 ( .A(n48838), .B(n48827), .Z(n48867) );
  XNOR U48692 ( .A(n48877), .B(n48878), .Z(n48827) );
  AND U48693 ( .A(n1739), .B(n48809), .Z(n48878) );
  XNOR U48694 ( .A(n48807), .B(n48877), .Z(n48809) );
  XNOR U48695 ( .A(n48879), .B(n48880), .Z(n1739) );
  AND U48696 ( .A(n48881), .B(n48882), .Z(n48880) );
  XNOR U48697 ( .A(n48879), .B(n48698), .Z(n48882) );
  IV U48698 ( .A(n48702), .Z(n48698) );
  XOR U48699 ( .A(n48883), .B(n48884), .Z(n48702) );
  AND U48700 ( .A(n1743), .B(n48885), .Z(n48884) );
  XOR U48701 ( .A(n48886), .B(n48883), .Z(n48885) );
  XNOR U48702 ( .A(n48879), .B(n48814), .Z(n48881) );
  XOR U48703 ( .A(n48887), .B(n48888), .Z(n48814) );
  AND U48704 ( .A(n1751), .B(n48849), .Z(n48888) );
  XOR U48705 ( .A(n48847), .B(n48887), .Z(n48849) );
  XOR U48706 ( .A(n48889), .B(n48890), .Z(n48879) );
  AND U48707 ( .A(n48891), .B(n48892), .Z(n48890) );
  XNOR U48708 ( .A(n48889), .B(n48714), .Z(n48892) );
  IV U48709 ( .A(n48717), .Z(n48714) );
  XOR U48710 ( .A(n48893), .B(n48894), .Z(n48717) );
  AND U48711 ( .A(n1743), .B(n48895), .Z(n48894) );
  XOR U48712 ( .A(n48896), .B(n48893), .Z(n48895) );
  XOR U48713 ( .A(n48718), .B(n48889), .Z(n48891) );
  XOR U48714 ( .A(n48897), .B(n48898), .Z(n48718) );
  AND U48715 ( .A(n1751), .B(n48857), .Z(n48898) );
  XOR U48716 ( .A(n48897), .B(n48855), .Z(n48857) );
  XOR U48717 ( .A(n48899), .B(n48900), .Z(n48889) );
  AND U48718 ( .A(n48901), .B(n48902), .Z(n48900) );
  XNOR U48719 ( .A(n48899), .B(n48742), .Z(n48902) );
  IV U48720 ( .A(n48745), .Z(n48742) );
  XOR U48721 ( .A(n48903), .B(n48904), .Z(n48745) );
  AND U48722 ( .A(n1743), .B(n48905), .Z(n48904) );
  XNOR U48723 ( .A(n48906), .B(n48903), .Z(n48905) );
  XOR U48724 ( .A(n48746), .B(n48899), .Z(n48901) );
  XOR U48725 ( .A(n48907), .B(n48908), .Z(n48746) );
  AND U48726 ( .A(n1751), .B(n48866), .Z(n48908) );
  XOR U48727 ( .A(n48907), .B(n48864), .Z(n48866) );
  XOR U48728 ( .A(n48823), .B(n48909), .Z(n48899) );
  AND U48729 ( .A(n48825), .B(n48910), .Z(n48909) );
  XNOR U48730 ( .A(n48823), .B(n48793), .Z(n48910) );
  IV U48731 ( .A(n48796), .Z(n48793) );
  XOR U48732 ( .A(n48911), .B(n48912), .Z(n48796) );
  AND U48733 ( .A(n1743), .B(n48913), .Z(n48912) );
  XOR U48734 ( .A(n48914), .B(n48911), .Z(n48913) );
  XOR U48735 ( .A(n48797), .B(n48823), .Z(n48825) );
  XOR U48736 ( .A(n48915), .B(n48916), .Z(n48797) );
  AND U48737 ( .A(n1751), .B(n48876), .Z(n48916) );
  XOR U48738 ( .A(n48915), .B(n48874), .Z(n48876) );
  AND U48739 ( .A(n48877), .B(n48807), .Z(n48823) );
  XNOR U48740 ( .A(n48917), .B(n48918), .Z(n48807) );
  AND U48741 ( .A(n1743), .B(n48919), .Z(n48918) );
  XNOR U48742 ( .A(n48920), .B(n48917), .Z(n48919) );
  XNOR U48743 ( .A(n48921), .B(n48922), .Z(n1743) );
  AND U48744 ( .A(n48923), .B(n48924), .Z(n48922) );
  XOR U48745 ( .A(n48886), .B(n48921), .Z(n48924) );
  AND U48746 ( .A(n48925), .B(n48926), .Z(n48886) );
  XNOR U48747 ( .A(n48883), .B(n48921), .Z(n48923) );
  XNOR U48748 ( .A(n48927), .B(n48928), .Z(n48883) );
  AND U48749 ( .A(n1747), .B(n48929), .Z(n48928) );
  XNOR U48750 ( .A(n48930), .B(n48931), .Z(n48929) );
  XOR U48751 ( .A(n48932), .B(n48933), .Z(n48921) );
  AND U48752 ( .A(n48934), .B(n48935), .Z(n48933) );
  XNOR U48753 ( .A(n48932), .B(n48925), .Z(n48935) );
  IV U48754 ( .A(n48896), .Z(n48925) );
  XOR U48755 ( .A(n48936), .B(n48937), .Z(n48896) );
  XOR U48756 ( .A(n48938), .B(n48926), .Z(n48937) );
  AND U48757 ( .A(n48906), .B(n48939), .Z(n48926) );
  AND U48758 ( .A(n48940), .B(n48941), .Z(n48938) );
  XOR U48759 ( .A(n48942), .B(n48936), .Z(n48940) );
  XNOR U48760 ( .A(n48893), .B(n48932), .Z(n48934) );
  XNOR U48761 ( .A(n48943), .B(n48944), .Z(n48893) );
  AND U48762 ( .A(n1747), .B(n48945), .Z(n48944) );
  XNOR U48763 ( .A(n48946), .B(n48947), .Z(n48945) );
  XOR U48764 ( .A(n48948), .B(n48949), .Z(n48932) );
  AND U48765 ( .A(n48950), .B(n48951), .Z(n48949) );
  XNOR U48766 ( .A(n48948), .B(n48906), .Z(n48951) );
  XOR U48767 ( .A(n48952), .B(n48941), .Z(n48906) );
  XNOR U48768 ( .A(n48953), .B(n48936), .Z(n48941) );
  XOR U48769 ( .A(n48954), .B(n48955), .Z(n48936) );
  AND U48770 ( .A(n48956), .B(n48957), .Z(n48955) );
  XOR U48771 ( .A(n48958), .B(n48954), .Z(n48956) );
  XNOR U48772 ( .A(n48959), .B(n48960), .Z(n48953) );
  AND U48773 ( .A(n48961), .B(n48962), .Z(n48960) );
  XOR U48774 ( .A(n48959), .B(n48963), .Z(n48961) );
  XNOR U48775 ( .A(n48942), .B(n48939), .Z(n48952) );
  AND U48776 ( .A(n48964), .B(n48965), .Z(n48939) );
  XOR U48777 ( .A(n48966), .B(n48967), .Z(n48942) );
  AND U48778 ( .A(n48968), .B(n48969), .Z(n48967) );
  XOR U48779 ( .A(n48966), .B(n48970), .Z(n48968) );
  XNOR U48780 ( .A(n48903), .B(n48948), .Z(n48950) );
  XNOR U48781 ( .A(n48971), .B(n48972), .Z(n48903) );
  AND U48782 ( .A(n1747), .B(n48973), .Z(n48972) );
  XNOR U48783 ( .A(n48974), .B(n48975), .Z(n48973) );
  XOR U48784 ( .A(n48976), .B(n48977), .Z(n48948) );
  AND U48785 ( .A(n48978), .B(n48979), .Z(n48977) );
  XNOR U48786 ( .A(n48976), .B(n48964), .Z(n48979) );
  IV U48787 ( .A(n48914), .Z(n48964) );
  XNOR U48788 ( .A(n48980), .B(n48957), .Z(n48914) );
  XNOR U48789 ( .A(n48981), .B(n48963), .Z(n48957) );
  XNOR U48790 ( .A(n48982), .B(n48983), .Z(n48963) );
  NOR U48791 ( .A(n48984), .B(n48985), .Z(n48983) );
  XOR U48792 ( .A(n48982), .B(n48986), .Z(n48984) );
  XNOR U48793 ( .A(n48962), .B(n48954), .Z(n48981) );
  XOR U48794 ( .A(n48987), .B(n48988), .Z(n48954) );
  AND U48795 ( .A(n48989), .B(n48990), .Z(n48988) );
  XOR U48796 ( .A(n48987), .B(n48991), .Z(n48989) );
  XNOR U48797 ( .A(n48992), .B(n48959), .Z(n48962) );
  XOR U48798 ( .A(n48993), .B(n48994), .Z(n48959) );
  AND U48799 ( .A(n48995), .B(n48996), .Z(n48994) );
  XNOR U48800 ( .A(n48997), .B(n48998), .Z(n48995) );
  IV U48801 ( .A(n48993), .Z(n48997) );
  XNOR U48802 ( .A(n48999), .B(n49000), .Z(n48992) );
  NOR U48803 ( .A(n49001), .B(n49002), .Z(n49000) );
  XNOR U48804 ( .A(n48999), .B(n49003), .Z(n49001) );
  XNOR U48805 ( .A(n48958), .B(n48965), .Z(n48980) );
  NOR U48806 ( .A(n48920), .B(n49004), .Z(n48965) );
  XOR U48807 ( .A(n48970), .B(n48969), .Z(n48958) );
  XNOR U48808 ( .A(n49005), .B(n48966), .Z(n48969) );
  XOR U48809 ( .A(n49006), .B(n49007), .Z(n48966) );
  AND U48810 ( .A(n49008), .B(n49009), .Z(n49007) );
  XNOR U48811 ( .A(n49010), .B(n49011), .Z(n49008) );
  IV U48812 ( .A(n49006), .Z(n49010) );
  XNOR U48813 ( .A(n49012), .B(n49013), .Z(n49005) );
  NOR U48814 ( .A(n49014), .B(n49015), .Z(n49013) );
  XNOR U48815 ( .A(n49012), .B(n49016), .Z(n49014) );
  XOR U48816 ( .A(n49017), .B(n49018), .Z(n48970) );
  NOR U48817 ( .A(n49019), .B(n49020), .Z(n49018) );
  XNOR U48818 ( .A(n49017), .B(n49021), .Z(n49019) );
  XNOR U48819 ( .A(n48911), .B(n48976), .Z(n48978) );
  XNOR U48820 ( .A(n49022), .B(n49023), .Z(n48911) );
  AND U48821 ( .A(n1747), .B(n49024), .Z(n49023) );
  XNOR U48822 ( .A(n49025), .B(n49026), .Z(n49024) );
  AND U48823 ( .A(n48917), .B(n48920), .Z(n48976) );
  XOR U48824 ( .A(n49027), .B(n49004), .Z(n48920) );
  XNOR U48825 ( .A(p_input[1408]), .B(p_input[2048]), .Z(n49004) );
  XNOR U48826 ( .A(n48991), .B(n48990), .Z(n49027) );
  XNOR U48827 ( .A(n49028), .B(n48998), .Z(n48990) );
  XNOR U48828 ( .A(n48986), .B(n48985), .Z(n48998) );
  XNOR U48829 ( .A(n49029), .B(n48982), .Z(n48985) );
  XNOR U48830 ( .A(p_input[1418]), .B(p_input[2058]), .Z(n48982) );
  XOR U48831 ( .A(p_input[1419]), .B(n29030), .Z(n49029) );
  XOR U48832 ( .A(p_input[1420]), .B(p_input[2060]), .Z(n48986) );
  XOR U48833 ( .A(n48996), .B(n49030), .Z(n49028) );
  IV U48834 ( .A(n48987), .Z(n49030) );
  XOR U48835 ( .A(p_input[1409]), .B(p_input[2049]), .Z(n48987) );
  XNOR U48836 ( .A(n49031), .B(n49003), .Z(n48996) );
  XNOR U48837 ( .A(p_input[1423]), .B(n29033), .Z(n49003) );
  XOR U48838 ( .A(n48993), .B(n49002), .Z(n49031) );
  XOR U48839 ( .A(n49032), .B(n48999), .Z(n49002) );
  XOR U48840 ( .A(p_input[1421]), .B(p_input[2061]), .Z(n48999) );
  XOR U48841 ( .A(p_input[1422]), .B(n29035), .Z(n49032) );
  XOR U48842 ( .A(p_input[1417]), .B(p_input[2057]), .Z(n48993) );
  XOR U48843 ( .A(n49011), .B(n49009), .Z(n48991) );
  XNOR U48844 ( .A(n49033), .B(n49016), .Z(n49009) );
  XOR U48845 ( .A(p_input[1416]), .B(p_input[2056]), .Z(n49016) );
  XOR U48846 ( .A(n49006), .B(n49015), .Z(n49033) );
  XOR U48847 ( .A(n49034), .B(n49012), .Z(n49015) );
  XOR U48848 ( .A(p_input[1414]), .B(p_input[2054]), .Z(n49012) );
  XOR U48849 ( .A(p_input[1415]), .B(n30404), .Z(n49034) );
  XOR U48850 ( .A(p_input[1410]), .B(p_input[2050]), .Z(n49006) );
  XNOR U48851 ( .A(n49021), .B(n49020), .Z(n49011) );
  XOR U48852 ( .A(n49035), .B(n49017), .Z(n49020) );
  XOR U48853 ( .A(p_input[1411]), .B(p_input[2051]), .Z(n49017) );
  XOR U48854 ( .A(p_input[1412]), .B(n30406), .Z(n49035) );
  XOR U48855 ( .A(p_input[1413]), .B(p_input[2053]), .Z(n49021) );
  XNOR U48856 ( .A(n49036), .B(n49037), .Z(n48917) );
  AND U48857 ( .A(n1747), .B(n49038), .Z(n49037) );
  XNOR U48858 ( .A(n49039), .B(n49040), .Z(n1747) );
  AND U48859 ( .A(n49041), .B(n49042), .Z(n49040) );
  XOR U48860 ( .A(n48931), .B(n49039), .Z(n49042) );
  XNOR U48861 ( .A(n49043), .B(n49039), .Z(n49041) );
  XOR U48862 ( .A(n49044), .B(n49045), .Z(n49039) );
  AND U48863 ( .A(n49046), .B(n49047), .Z(n49045) );
  XOR U48864 ( .A(n48946), .B(n49044), .Z(n49047) );
  XOR U48865 ( .A(n49044), .B(n48947), .Z(n49046) );
  XOR U48866 ( .A(n49048), .B(n49049), .Z(n49044) );
  AND U48867 ( .A(n49050), .B(n49051), .Z(n49049) );
  XOR U48868 ( .A(n48974), .B(n49048), .Z(n49051) );
  XOR U48869 ( .A(n49048), .B(n48975), .Z(n49050) );
  XOR U48870 ( .A(n49052), .B(n49053), .Z(n49048) );
  AND U48871 ( .A(n49054), .B(n49055), .Z(n49053) );
  XOR U48872 ( .A(n49052), .B(n49025), .Z(n49055) );
  XNOR U48873 ( .A(n49056), .B(n49057), .Z(n48877) );
  AND U48874 ( .A(n1751), .B(n49058), .Z(n49057) );
  XNOR U48875 ( .A(n49059), .B(n49060), .Z(n1751) );
  AND U48876 ( .A(n49061), .B(n49062), .Z(n49060) );
  XOR U48877 ( .A(n49059), .B(n48887), .Z(n49062) );
  XNOR U48878 ( .A(n49059), .B(n48847), .Z(n49061) );
  XOR U48879 ( .A(n49063), .B(n49064), .Z(n49059) );
  AND U48880 ( .A(n49065), .B(n49066), .Z(n49064) );
  XOR U48881 ( .A(n49063), .B(n48855), .Z(n49065) );
  XOR U48882 ( .A(n49067), .B(n49068), .Z(n48838) );
  AND U48883 ( .A(n1755), .B(n49058), .Z(n49068) );
  XNOR U48884 ( .A(n49056), .B(n49067), .Z(n49058) );
  XNOR U48885 ( .A(n49069), .B(n49070), .Z(n1755) );
  AND U48886 ( .A(n49071), .B(n49072), .Z(n49070) );
  XNOR U48887 ( .A(n49073), .B(n49069), .Z(n49072) );
  IV U48888 ( .A(n48887), .Z(n49073) );
  XOR U48889 ( .A(n49043), .B(n49074), .Z(n48887) );
  AND U48890 ( .A(n1758), .B(n49075), .Z(n49074) );
  XOR U48891 ( .A(n48930), .B(n48927), .Z(n49075) );
  IV U48892 ( .A(n49043), .Z(n48930) );
  XNOR U48893 ( .A(n48847), .B(n49069), .Z(n49071) );
  XOR U48894 ( .A(n49076), .B(n49077), .Z(n48847) );
  AND U48895 ( .A(n1774), .B(n49078), .Z(n49077) );
  XOR U48896 ( .A(n49063), .B(n49079), .Z(n49069) );
  AND U48897 ( .A(n49080), .B(n49066), .Z(n49079) );
  XNOR U48898 ( .A(n48897), .B(n49063), .Z(n49066) );
  XOR U48899 ( .A(n48947), .B(n49081), .Z(n48897) );
  AND U48900 ( .A(n1758), .B(n49082), .Z(n49081) );
  XOR U48901 ( .A(n48943), .B(n48947), .Z(n49082) );
  XNOR U48902 ( .A(n49083), .B(n49063), .Z(n49080) );
  IV U48903 ( .A(n48855), .Z(n49083) );
  XOR U48904 ( .A(n49084), .B(n49085), .Z(n48855) );
  AND U48905 ( .A(n1774), .B(n49086), .Z(n49085) );
  XOR U48906 ( .A(n49087), .B(n49088), .Z(n49063) );
  AND U48907 ( .A(n49089), .B(n49090), .Z(n49088) );
  XNOR U48908 ( .A(n48907), .B(n49087), .Z(n49090) );
  XOR U48909 ( .A(n48975), .B(n49091), .Z(n48907) );
  AND U48910 ( .A(n1758), .B(n49092), .Z(n49091) );
  XOR U48911 ( .A(n48971), .B(n48975), .Z(n49092) );
  XOR U48912 ( .A(n49087), .B(n48864), .Z(n49089) );
  XOR U48913 ( .A(n49093), .B(n49094), .Z(n48864) );
  AND U48914 ( .A(n1774), .B(n49095), .Z(n49094) );
  XOR U48915 ( .A(n49096), .B(n49097), .Z(n49087) );
  AND U48916 ( .A(n49098), .B(n49099), .Z(n49097) );
  XNOR U48917 ( .A(n49096), .B(n48915), .Z(n49099) );
  XOR U48918 ( .A(n49026), .B(n49100), .Z(n48915) );
  AND U48919 ( .A(n1758), .B(n49101), .Z(n49100) );
  XOR U48920 ( .A(n49022), .B(n49026), .Z(n49101) );
  XNOR U48921 ( .A(n49102), .B(n49096), .Z(n49098) );
  IV U48922 ( .A(n48874), .Z(n49102) );
  XOR U48923 ( .A(n49103), .B(n49104), .Z(n48874) );
  AND U48924 ( .A(n1774), .B(n49105), .Z(n49104) );
  AND U48925 ( .A(n49067), .B(n49056), .Z(n49096) );
  XNOR U48926 ( .A(n49106), .B(n49107), .Z(n49056) );
  AND U48927 ( .A(n1758), .B(n49038), .Z(n49107) );
  XNOR U48928 ( .A(n49036), .B(n49106), .Z(n49038) );
  XNOR U48929 ( .A(n49108), .B(n49109), .Z(n1758) );
  AND U48930 ( .A(n49110), .B(n49111), .Z(n49109) );
  XNOR U48931 ( .A(n49108), .B(n48927), .Z(n49111) );
  IV U48932 ( .A(n48931), .Z(n48927) );
  XOR U48933 ( .A(n49112), .B(n49113), .Z(n48931) );
  AND U48934 ( .A(n1762), .B(n49114), .Z(n49113) );
  XOR U48935 ( .A(n49115), .B(n49112), .Z(n49114) );
  XNOR U48936 ( .A(n49108), .B(n49043), .Z(n49110) );
  XOR U48937 ( .A(n49116), .B(n49117), .Z(n49043) );
  AND U48938 ( .A(n1770), .B(n49078), .Z(n49117) );
  XOR U48939 ( .A(n49076), .B(n49116), .Z(n49078) );
  XOR U48940 ( .A(n49118), .B(n49119), .Z(n49108) );
  AND U48941 ( .A(n49120), .B(n49121), .Z(n49119) );
  XNOR U48942 ( .A(n49118), .B(n48943), .Z(n49121) );
  IV U48943 ( .A(n48946), .Z(n48943) );
  XOR U48944 ( .A(n49122), .B(n49123), .Z(n48946) );
  AND U48945 ( .A(n1762), .B(n49124), .Z(n49123) );
  XOR U48946 ( .A(n49125), .B(n49122), .Z(n49124) );
  XOR U48947 ( .A(n48947), .B(n49118), .Z(n49120) );
  XOR U48948 ( .A(n49126), .B(n49127), .Z(n48947) );
  AND U48949 ( .A(n1770), .B(n49086), .Z(n49127) );
  XOR U48950 ( .A(n49126), .B(n49084), .Z(n49086) );
  XOR U48951 ( .A(n49128), .B(n49129), .Z(n49118) );
  AND U48952 ( .A(n49130), .B(n49131), .Z(n49129) );
  XNOR U48953 ( .A(n49128), .B(n48971), .Z(n49131) );
  IV U48954 ( .A(n48974), .Z(n48971) );
  XOR U48955 ( .A(n49132), .B(n49133), .Z(n48974) );
  AND U48956 ( .A(n1762), .B(n49134), .Z(n49133) );
  XNOR U48957 ( .A(n49135), .B(n49132), .Z(n49134) );
  XOR U48958 ( .A(n48975), .B(n49128), .Z(n49130) );
  XOR U48959 ( .A(n49136), .B(n49137), .Z(n48975) );
  AND U48960 ( .A(n1770), .B(n49095), .Z(n49137) );
  XOR U48961 ( .A(n49136), .B(n49093), .Z(n49095) );
  XOR U48962 ( .A(n49052), .B(n49138), .Z(n49128) );
  AND U48963 ( .A(n49054), .B(n49139), .Z(n49138) );
  XNOR U48964 ( .A(n49052), .B(n49022), .Z(n49139) );
  IV U48965 ( .A(n49025), .Z(n49022) );
  XOR U48966 ( .A(n49140), .B(n49141), .Z(n49025) );
  AND U48967 ( .A(n1762), .B(n49142), .Z(n49141) );
  XOR U48968 ( .A(n49143), .B(n49140), .Z(n49142) );
  XOR U48969 ( .A(n49026), .B(n49052), .Z(n49054) );
  XOR U48970 ( .A(n49144), .B(n49145), .Z(n49026) );
  AND U48971 ( .A(n1770), .B(n49105), .Z(n49145) );
  XOR U48972 ( .A(n49144), .B(n49103), .Z(n49105) );
  AND U48973 ( .A(n49106), .B(n49036), .Z(n49052) );
  XNOR U48974 ( .A(n49146), .B(n49147), .Z(n49036) );
  AND U48975 ( .A(n1762), .B(n49148), .Z(n49147) );
  XNOR U48976 ( .A(n49149), .B(n49146), .Z(n49148) );
  XNOR U48977 ( .A(n49150), .B(n49151), .Z(n1762) );
  AND U48978 ( .A(n49152), .B(n49153), .Z(n49151) );
  XOR U48979 ( .A(n49115), .B(n49150), .Z(n49153) );
  AND U48980 ( .A(n49154), .B(n49155), .Z(n49115) );
  XNOR U48981 ( .A(n49112), .B(n49150), .Z(n49152) );
  XNOR U48982 ( .A(n49156), .B(n49157), .Z(n49112) );
  AND U48983 ( .A(n1766), .B(n49158), .Z(n49157) );
  XNOR U48984 ( .A(n49159), .B(n49160), .Z(n49158) );
  XOR U48985 ( .A(n49161), .B(n49162), .Z(n49150) );
  AND U48986 ( .A(n49163), .B(n49164), .Z(n49162) );
  XNOR U48987 ( .A(n49161), .B(n49154), .Z(n49164) );
  IV U48988 ( .A(n49125), .Z(n49154) );
  XOR U48989 ( .A(n49165), .B(n49166), .Z(n49125) );
  XOR U48990 ( .A(n49167), .B(n49155), .Z(n49166) );
  AND U48991 ( .A(n49135), .B(n49168), .Z(n49155) );
  AND U48992 ( .A(n49169), .B(n49170), .Z(n49167) );
  XOR U48993 ( .A(n49171), .B(n49165), .Z(n49169) );
  XNOR U48994 ( .A(n49122), .B(n49161), .Z(n49163) );
  XNOR U48995 ( .A(n49172), .B(n49173), .Z(n49122) );
  AND U48996 ( .A(n1766), .B(n49174), .Z(n49173) );
  XNOR U48997 ( .A(n49175), .B(n49176), .Z(n49174) );
  XOR U48998 ( .A(n49177), .B(n49178), .Z(n49161) );
  AND U48999 ( .A(n49179), .B(n49180), .Z(n49178) );
  XNOR U49000 ( .A(n49177), .B(n49135), .Z(n49180) );
  XOR U49001 ( .A(n49181), .B(n49170), .Z(n49135) );
  XNOR U49002 ( .A(n49182), .B(n49165), .Z(n49170) );
  XOR U49003 ( .A(n49183), .B(n49184), .Z(n49165) );
  AND U49004 ( .A(n49185), .B(n49186), .Z(n49184) );
  XOR U49005 ( .A(n49187), .B(n49183), .Z(n49185) );
  XNOR U49006 ( .A(n49188), .B(n49189), .Z(n49182) );
  AND U49007 ( .A(n49190), .B(n49191), .Z(n49189) );
  XOR U49008 ( .A(n49188), .B(n49192), .Z(n49190) );
  XNOR U49009 ( .A(n49171), .B(n49168), .Z(n49181) );
  AND U49010 ( .A(n49193), .B(n49194), .Z(n49168) );
  XOR U49011 ( .A(n49195), .B(n49196), .Z(n49171) );
  AND U49012 ( .A(n49197), .B(n49198), .Z(n49196) );
  XOR U49013 ( .A(n49195), .B(n49199), .Z(n49197) );
  XNOR U49014 ( .A(n49132), .B(n49177), .Z(n49179) );
  XNOR U49015 ( .A(n49200), .B(n49201), .Z(n49132) );
  AND U49016 ( .A(n1766), .B(n49202), .Z(n49201) );
  XNOR U49017 ( .A(n49203), .B(n49204), .Z(n49202) );
  XOR U49018 ( .A(n49205), .B(n49206), .Z(n49177) );
  AND U49019 ( .A(n49207), .B(n49208), .Z(n49206) );
  XNOR U49020 ( .A(n49205), .B(n49193), .Z(n49208) );
  IV U49021 ( .A(n49143), .Z(n49193) );
  XNOR U49022 ( .A(n49209), .B(n49186), .Z(n49143) );
  XNOR U49023 ( .A(n49210), .B(n49192), .Z(n49186) );
  XNOR U49024 ( .A(n49211), .B(n49212), .Z(n49192) );
  NOR U49025 ( .A(n49213), .B(n49214), .Z(n49212) );
  XOR U49026 ( .A(n49211), .B(n49215), .Z(n49213) );
  XNOR U49027 ( .A(n49191), .B(n49183), .Z(n49210) );
  XOR U49028 ( .A(n49216), .B(n49217), .Z(n49183) );
  AND U49029 ( .A(n49218), .B(n49219), .Z(n49217) );
  XOR U49030 ( .A(n49216), .B(n49220), .Z(n49218) );
  XNOR U49031 ( .A(n49221), .B(n49188), .Z(n49191) );
  XOR U49032 ( .A(n49222), .B(n49223), .Z(n49188) );
  AND U49033 ( .A(n49224), .B(n49225), .Z(n49223) );
  XNOR U49034 ( .A(n49226), .B(n49227), .Z(n49224) );
  IV U49035 ( .A(n49222), .Z(n49226) );
  XNOR U49036 ( .A(n49228), .B(n49229), .Z(n49221) );
  NOR U49037 ( .A(n49230), .B(n49231), .Z(n49229) );
  XNOR U49038 ( .A(n49228), .B(n49232), .Z(n49230) );
  XNOR U49039 ( .A(n49187), .B(n49194), .Z(n49209) );
  NOR U49040 ( .A(n49149), .B(n49233), .Z(n49194) );
  XOR U49041 ( .A(n49199), .B(n49198), .Z(n49187) );
  XNOR U49042 ( .A(n49234), .B(n49195), .Z(n49198) );
  XOR U49043 ( .A(n49235), .B(n49236), .Z(n49195) );
  AND U49044 ( .A(n49237), .B(n49238), .Z(n49236) );
  XNOR U49045 ( .A(n49239), .B(n49240), .Z(n49237) );
  IV U49046 ( .A(n49235), .Z(n49239) );
  XNOR U49047 ( .A(n49241), .B(n49242), .Z(n49234) );
  NOR U49048 ( .A(n49243), .B(n49244), .Z(n49242) );
  XNOR U49049 ( .A(n49241), .B(n49245), .Z(n49243) );
  XOR U49050 ( .A(n49246), .B(n49247), .Z(n49199) );
  NOR U49051 ( .A(n49248), .B(n49249), .Z(n49247) );
  XNOR U49052 ( .A(n49246), .B(n49250), .Z(n49248) );
  XNOR U49053 ( .A(n49140), .B(n49205), .Z(n49207) );
  XNOR U49054 ( .A(n49251), .B(n49252), .Z(n49140) );
  AND U49055 ( .A(n1766), .B(n49253), .Z(n49252) );
  XNOR U49056 ( .A(n49254), .B(n49255), .Z(n49253) );
  AND U49057 ( .A(n49146), .B(n49149), .Z(n49205) );
  XOR U49058 ( .A(n49256), .B(n49233), .Z(n49149) );
  XNOR U49059 ( .A(p_input[1424]), .B(p_input[2048]), .Z(n49233) );
  XNOR U49060 ( .A(n49220), .B(n49219), .Z(n49256) );
  XNOR U49061 ( .A(n49257), .B(n49227), .Z(n49219) );
  XNOR U49062 ( .A(n49215), .B(n49214), .Z(n49227) );
  XNOR U49063 ( .A(n49258), .B(n49211), .Z(n49214) );
  XNOR U49064 ( .A(p_input[1434]), .B(p_input[2058]), .Z(n49211) );
  XOR U49065 ( .A(p_input[1435]), .B(n29030), .Z(n49258) );
  XOR U49066 ( .A(p_input[1436]), .B(p_input[2060]), .Z(n49215) );
  XOR U49067 ( .A(n49225), .B(n49259), .Z(n49257) );
  IV U49068 ( .A(n49216), .Z(n49259) );
  XOR U49069 ( .A(p_input[1425]), .B(p_input[2049]), .Z(n49216) );
  XNOR U49070 ( .A(n49260), .B(n49232), .Z(n49225) );
  XNOR U49071 ( .A(p_input[1439]), .B(n29033), .Z(n49232) );
  XOR U49072 ( .A(n49222), .B(n49231), .Z(n49260) );
  XOR U49073 ( .A(n49261), .B(n49228), .Z(n49231) );
  XOR U49074 ( .A(p_input[1437]), .B(p_input[2061]), .Z(n49228) );
  XOR U49075 ( .A(p_input[1438]), .B(n29035), .Z(n49261) );
  XOR U49076 ( .A(p_input[1433]), .B(p_input[2057]), .Z(n49222) );
  XOR U49077 ( .A(n49240), .B(n49238), .Z(n49220) );
  XNOR U49078 ( .A(n49262), .B(n49245), .Z(n49238) );
  XOR U49079 ( .A(p_input[1432]), .B(p_input[2056]), .Z(n49245) );
  XOR U49080 ( .A(n49235), .B(n49244), .Z(n49262) );
  XOR U49081 ( .A(n49263), .B(n49241), .Z(n49244) );
  XOR U49082 ( .A(p_input[1430]), .B(p_input[2054]), .Z(n49241) );
  XOR U49083 ( .A(p_input[1431]), .B(n30404), .Z(n49263) );
  XOR U49084 ( .A(p_input[1426]), .B(p_input[2050]), .Z(n49235) );
  XNOR U49085 ( .A(n49250), .B(n49249), .Z(n49240) );
  XOR U49086 ( .A(n49264), .B(n49246), .Z(n49249) );
  XOR U49087 ( .A(p_input[1427]), .B(p_input[2051]), .Z(n49246) );
  XOR U49088 ( .A(p_input[1428]), .B(n30406), .Z(n49264) );
  XOR U49089 ( .A(p_input[1429]), .B(p_input[2053]), .Z(n49250) );
  XNOR U49090 ( .A(n49265), .B(n49266), .Z(n49146) );
  AND U49091 ( .A(n1766), .B(n49267), .Z(n49266) );
  XNOR U49092 ( .A(n49268), .B(n49269), .Z(n1766) );
  AND U49093 ( .A(n49270), .B(n49271), .Z(n49269) );
  XOR U49094 ( .A(n49160), .B(n49268), .Z(n49271) );
  XNOR U49095 ( .A(n49272), .B(n49268), .Z(n49270) );
  XOR U49096 ( .A(n49273), .B(n49274), .Z(n49268) );
  AND U49097 ( .A(n49275), .B(n49276), .Z(n49274) );
  XOR U49098 ( .A(n49175), .B(n49273), .Z(n49276) );
  XOR U49099 ( .A(n49273), .B(n49176), .Z(n49275) );
  XOR U49100 ( .A(n49277), .B(n49278), .Z(n49273) );
  AND U49101 ( .A(n49279), .B(n49280), .Z(n49278) );
  XOR U49102 ( .A(n49203), .B(n49277), .Z(n49280) );
  XOR U49103 ( .A(n49277), .B(n49204), .Z(n49279) );
  XOR U49104 ( .A(n49281), .B(n49282), .Z(n49277) );
  AND U49105 ( .A(n49283), .B(n49284), .Z(n49282) );
  XOR U49106 ( .A(n49281), .B(n49254), .Z(n49284) );
  XNOR U49107 ( .A(n49285), .B(n49286), .Z(n49106) );
  AND U49108 ( .A(n1770), .B(n49287), .Z(n49286) );
  XNOR U49109 ( .A(n49288), .B(n49289), .Z(n1770) );
  AND U49110 ( .A(n49290), .B(n49291), .Z(n49289) );
  XOR U49111 ( .A(n49288), .B(n49116), .Z(n49291) );
  XNOR U49112 ( .A(n49288), .B(n49076), .Z(n49290) );
  XOR U49113 ( .A(n49292), .B(n49293), .Z(n49288) );
  AND U49114 ( .A(n49294), .B(n49295), .Z(n49293) );
  XOR U49115 ( .A(n49292), .B(n49084), .Z(n49294) );
  XOR U49116 ( .A(n49296), .B(n49297), .Z(n49067) );
  AND U49117 ( .A(n1774), .B(n49287), .Z(n49297) );
  XNOR U49118 ( .A(n49285), .B(n49296), .Z(n49287) );
  XNOR U49119 ( .A(n49298), .B(n49299), .Z(n1774) );
  AND U49120 ( .A(n49300), .B(n49301), .Z(n49299) );
  XNOR U49121 ( .A(n49302), .B(n49298), .Z(n49301) );
  IV U49122 ( .A(n49116), .Z(n49302) );
  XOR U49123 ( .A(n49272), .B(n49303), .Z(n49116) );
  AND U49124 ( .A(n1777), .B(n49304), .Z(n49303) );
  XOR U49125 ( .A(n49159), .B(n49156), .Z(n49304) );
  IV U49126 ( .A(n49272), .Z(n49159) );
  XNOR U49127 ( .A(n49076), .B(n49298), .Z(n49300) );
  XOR U49128 ( .A(n49305), .B(n49306), .Z(n49076) );
  AND U49129 ( .A(n1793), .B(n49307), .Z(n49306) );
  XOR U49130 ( .A(n49292), .B(n49308), .Z(n49298) );
  AND U49131 ( .A(n49309), .B(n49295), .Z(n49308) );
  XNOR U49132 ( .A(n49126), .B(n49292), .Z(n49295) );
  XOR U49133 ( .A(n49176), .B(n49310), .Z(n49126) );
  AND U49134 ( .A(n1777), .B(n49311), .Z(n49310) );
  XOR U49135 ( .A(n49172), .B(n49176), .Z(n49311) );
  XNOR U49136 ( .A(n49312), .B(n49292), .Z(n49309) );
  IV U49137 ( .A(n49084), .Z(n49312) );
  XOR U49138 ( .A(n49313), .B(n49314), .Z(n49084) );
  AND U49139 ( .A(n1793), .B(n49315), .Z(n49314) );
  XOR U49140 ( .A(n49316), .B(n49317), .Z(n49292) );
  AND U49141 ( .A(n49318), .B(n49319), .Z(n49317) );
  XNOR U49142 ( .A(n49136), .B(n49316), .Z(n49319) );
  XOR U49143 ( .A(n49204), .B(n49320), .Z(n49136) );
  AND U49144 ( .A(n1777), .B(n49321), .Z(n49320) );
  XOR U49145 ( .A(n49200), .B(n49204), .Z(n49321) );
  XOR U49146 ( .A(n49316), .B(n49093), .Z(n49318) );
  XOR U49147 ( .A(n49322), .B(n49323), .Z(n49093) );
  AND U49148 ( .A(n1793), .B(n49324), .Z(n49323) );
  XOR U49149 ( .A(n49325), .B(n49326), .Z(n49316) );
  AND U49150 ( .A(n49327), .B(n49328), .Z(n49326) );
  XNOR U49151 ( .A(n49325), .B(n49144), .Z(n49328) );
  XOR U49152 ( .A(n49255), .B(n49329), .Z(n49144) );
  AND U49153 ( .A(n1777), .B(n49330), .Z(n49329) );
  XOR U49154 ( .A(n49251), .B(n49255), .Z(n49330) );
  XNOR U49155 ( .A(n49331), .B(n49325), .Z(n49327) );
  IV U49156 ( .A(n49103), .Z(n49331) );
  XOR U49157 ( .A(n49332), .B(n49333), .Z(n49103) );
  AND U49158 ( .A(n1793), .B(n49334), .Z(n49333) );
  AND U49159 ( .A(n49296), .B(n49285), .Z(n49325) );
  XNOR U49160 ( .A(n49335), .B(n49336), .Z(n49285) );
  AND U49161 ( .A(n1777), .B(n49267), .Z(n49336) );
  XNOR U49162 ( .A(n49265), .B(n49335), .Z(n49267) );
  XNOR U49163 ( .A(n49337), .B(n49338), .Z(n1777) );
  AND U49164 ( .A(n49339), .B(n49340), .Z(n49338) );
  XNOR U49165 ( .A(n49337), .B(n49156), .Z(n49340) );
  IV U49166 ( .A(n49160), .Z(n49156) );
  XOR U49167 ( .A(n49341), .B(n49342), .Z(n49160) );
  AND U49168 ( .A(n1781), .B(n49343), .Z(n49342) );
  XOR U49169 ( .A(n49344), .B(n49341), .Z(n49343) );
  XNOR U49170 ( .A(n49337), .B(n49272), .Z(n49339) );
  XOR U49171 ( .A(n49345), .B(n49346), .Z(n49272) );
  AND U49172 ( .A(n1789), .B(n49307), .Z(n49346) );
  XOR U49173 ( .A(n49305), .B(n49345), .Z(n49307) );
  XOR U49174 ( .A(n49347), .B(n49348), .Z(n49337) );
  AND U49175 ( .A(n49349), .B(n49350), .Z(n49348) );
  XNOR U49176 ( .A(n49347), .B(n49172), .Z(n49350) );
  IV U49177 ( .A(n49175), .Z(n49172) );
  XOR U49178 ( .A(n49351), .B(n49352), .Z(n49175) );
  AND U49179 ( .A(n1781), .B(n49353), .Z(n49352) );
  XOR U49180 ( .A(n49354), .B(n49351), .Z(n49353) );
  XOR U49181 ( .A(n49176), .B(n49347), .Z(n49349) );
  XOR U49182 ( .A(n49355), .B(n49356), .Z(n49176) );
  AND U49183 ( .A(n1789), .B(n49315), .Z(n49356) );
  XOR U49184 ( .A(n49355), .B(n49313), .Z(n49315) );
  XOR U49185 ( .A(n49357), .B(n49358), .Z(n49347) );
  AND U49186 ( .A(n49359), .B(n49360), .Z(n49358) );
  XNOR U49187 ( .A(n49357), .B(n49200), .Z(n49360) );
  IV U49188 ( .A(n49203), .Z(n49200) );
  XOR U49189 ( .A(n49361), .B(n49362), .Z(n49203) );
  AND U49190 ( .A(n1781), .B(n49363), .Z(n49362) );
  XNOR U49191 ( .A(n49364), .B(n49361), .Z(n49363) );
  XOR U49192 ( .A(n49204), .B(n49357), .Z(n49359) );
  XOR U49193 ( .A(n49365), .B(n49366), .Z(n49204) );
  AND U49194 ( .A(n1789), .B(n49324), .Z(n49366) );
  XOR U49195 ( .A(n49365), .B(n49322), .Z(n49324) );
  XOR U49196 ( .A(n49281), .B(n49367), .Z(n49357) );
  AND U49197 ( .A(n49283), .B(n49368), .Z(n49367) );
  XNOR U49198 ( .A(n49281), .B(n49251), .Z(n49368) );
  IV U49199 ( .A(n49254), .Z(n49251) );
  XOR U49200 ( .A(n49369), .B(n49370), .Z(n49254) );
  AND U49201 ( .A(n1781), .B(n49371), .Z(n49370) );
  XOR U49202 ( .A(n49372), .B(n49369), .Z(n49371) );
  XOR U49203 ( .A(n49255), .B(n49281), .Z(n49283) );
  XOR U49204 ( .A(n49373), .B(n49374), .Z(n49255) );
  AND U49205 ( .A(n1789), .B(n49334), .Z(n49374) );
  XOR U49206 ( .A(n49373), .B(n49332), .Z(n49334) );
  AND U49207 ( .A(n49335), .B(n49265), .Z(n49281) );
  XNOR U49208 ( .A(n49375), .B(n49376), .Z(n49265) );
  AND U49209 ( .A(n1781), .B(n49377), .Z(n49376) );
  XNOR U49210 ( .A(n49378), .B(n49375), .Z(n49377) );
  XNOR U49211 ( .A(n49379), .B(n49380), .Z(n1781) );
  AND U49212 ( .A(n49381), .B(n49382), .Z(n49380) );
  XOR U49213 ( .A(n49344), .B(n49379), .Z(n49382) );
  AND U49214 ( .A(n49383), .B(n49384), .Z(n49344) );
  XNOR U49215 ( .A(n49341), .B(n49379), .Z(n49381) );
  XNOR U49216 ( .A(n49385), .B(n49386), .Z(n49341) );
  AND U49217 ( .A(n1785), .B(n49387), .Z(n49386) );
  XNOR U49218 ( .A(n49388), .B(n49389), .Z(n49387) );
  XOR U49219 ( .A(n49390), .B(n49391), .Z(n49379) );
  AND U49220 ( .A(n49392), .B(n49393), .Z(n49391) );
  XNOR U49221 ( .A(n49390), .B(n49383), .Z(n49393) );
  IV U49222 ( .A(n49354), .Z(n49383) );
  XOR U49223 ( .A(n49394), .B(n49395), .Z(n49354) );
  XOR U49224 ( .A(n49396), .B(n49384), .Z(n49395) );
  AND U49225 ( .A(n49364), .B(n49397), .Z(n49384) );
  AND U49226 ( .A(n49398), .B(n49399), .Z(n49396) );
  XOR U49227 ( .A(n49400), .B(n49394), .Z(n49398) );
  XNOR U49228 ( .A(n49351), .B(n49390), .Z(n49392) );
  XNOR U49229 ( .A(n49401), .B(n49402), .Z(n49351) );
  AND U49230 ( .A(n1785), .B(n49403), .Z(n49402) );
  XNOR U49231 ( .A(n49404), .B(n49405), .Z(n49403) );
  XOR U49232 ( .A(n49406), .B(n49407), .Z(n49390) );
  AND U49233 ( .A(n49408), .B(n49409), .Z(n49407) );
  XNOR U49234 ( .A(n49406), .B(n49364), .Z(n49409) );
  XOR U49235 ( .A(n49410), .B(n49399), .Z(n49364) );
  XNOR U49236 ( .A(n49411), .B(n49394), .Z(n49399) );
  XOR U49237 ( .A(n49412), .B(n49413), .Z(n49394) );
  AND U49238 ( .A(n49414), .B(n49415), .Z(n49413) );
  XOR U49239 ( .A(n49416), .B(n49412), .Z(n49414) );
  XNOR U49240 ( .A(n49417), .B(n49418), .Z(n49411) );
  AND U49241 ( .A(n49419), .B(n49420), .Z(n49418) );
  XOR U49242 ( .A(n49417), .B(n49421), .Z(n49419) );
  XNOR U49243 ( .A(n49400), .B(n49397), .Z(n49410) );
  AND U49244 ( .A(n49422), .B(n49423), .Z(n49397) );
  XOR U49245 ( .A(n49424), .B(n49425), .Z(n49400) );
  AND U49246 ( .A(n49426), .B(n49427), .Z(n49425) );
  XOR U49247 ( .A(n49424), .B(n49428), .Z(n49426) );
  XNOR U49248 ( .A(n49361), .B(n49406), .Z(n49408) );
  XNOR U49249 ( .A(n49429), .B(n49430), .Z(n49361) );
  AND U49250 ( .A(n1785), .B(n49431), .Z(n49430) );
  XNOR U49251 ( .A(n49432), .B(n49433), .Z(n49431) );
  XOR U49252 ( .A(n49434), .B(n49435), .Z(n49406) );
  AND U49253 ( .A(n49436), .B(n49437), .Z(n49435) );
  XNOR U49254 ( .A(n49434), .B(n49422), .Z(n49437) );
  IV U49255 ( .A(n49372), .Z(n49422) );
  XNOR U49256 ( .A(n49438), .B(n49415), .Z(n49372) );
  XNOR U49257 ( .A(n49439), .B(n49421), .Z(n49415) );
  XNOR U49258 ( .A(n49440), .B(n49441), .Z(n49421) );
  NOR U49259 ( .A(n49442), .B(n49443), .Z(n49441) );
  XOR U49260 ( .A(n49440), .B(n49444), .Z(n49442) );
  XNOR U49261 ( .A(n49420), .B(n49412), .Z(n49439) );
  XOR U49262 ( .A(n49445), .B(n49446), .Z(n49412) );
  AND U49263 ( .A(n49447), .B(n49448), .Z(n49446) );
  XOR U49264 ( .A(n49445), .B(n49449), .Z(n49447) );
  XNOR U49265 ( .A(n49450), .B(n49417), .Z(n49420) );
  XOR U49266 ( .A(n49451), .B(n49452), .Z(n49417) );
  AND U49267 ( .A(n49453), .B(n49454), .Z(n49452) );
  XNOR U49268 ( .A(n49455), .B(n49456), .Z(n49453) );
  IV U49269 ( .A(n49451), .Z(n49455) );
  XNOR U49270 ( .A(n49457), .B(n49458), .Z(n49450) );
  NOR U49271 ( .A(n49459), .B(n49460), .Z(n49458) );
  XNOR U49272 ( .A(n49457), .B(n49461), .Z(n49459) );
  XNOR U49273 ( .A(n49416), .B(n49423), .Z(n49438) );
  NOR U49274 ( .A(n49378), .B(n49462), .Z(n49423) );
  XOR U49275 ( .A(n49428), .B(n49427), .Z(n49416) );
  XNOR U49276 ( .A(n49463), .B(n49424), .Z(n49427) );
  XOR U49277 ( .A(n49464), .B(n49465), .Z(n49424) );
  AND U49278 ( .A(n49466), .B(n49467), .Z(n49465) );
  XNOR U49279 ( .A(n49468), .B(n49469), .Z(n49466) );
  IV U49280 ( .A(n49464), .Z(n49468) );
  XNOR U49281 ( .A(n49470), .B(n49471), .Z(n49463) );
  NOR U49282 ( .A(n49472), .B(n49473), .Z(n49471) );
  XNOR U49283 ( .A(n49470), .B(n49474), .Z(n49472) );
  XOR U49284 ( .A(n49475), .B(n49476), .Z(n49428) );
  NOR U49285 ( .A(n49477), .B(n49478), .Z(n49476) );
  XNOR U49286 ( .A(n49475), .B(n49479), .Z(n49477) );
  XNOR U49287 ( .A(n49369), .B(n49434), .Z(n49436) );
  XNOR U49288 ( .A(n49480), .B(n49481), .Z(n49369) );
  AND U49289 ( .A(n1785), .B(n49482), .Z(n49481) );
  XNOR U49290 ( .A(n49483), .B(n49484), .Z(n49482) );
  AND U49291 ( .A(n49375), .B(n49378), .Z(n49434) );
  XOR U49292 ( .A(n49485), .B(n49462), .Z(n49378) );
  XNOR U49293 ( .A(p_input[1440]), .B(p_input[2048]), .Z(n49462) );
  XNOR U49294 ( .A(n49449), .B(n49448), .Z(n49485) );
  XNOR U49295 ( .A(n49486), .B(n49456), .Z(n49448) );
  XNOR U49296 ( .A(n49444), .B(n49443), .Z(n49456) );
  XNOR U49297 ( .A(n49487), .B(n49440), .Z(n49443) );
  XNOR U49298 ( .A(p_input[1450]), .B(p_input[2058]), .Z(n49440) );
  XOR U49299 ( .A(p_input[1451]), .B(n29030), .Z(n49487) );
  XOR U49300 ( .A(p_input[1452]), .B(p_input[2060]), .Z(n49444) );
  XOR U49301 ( .A(n49454), .B(n49488), .Z(n49486) );
  IV U49302 ( .A(n49445), .Z(n49488) );
  XOR U49303 ( .A(p_input[1441]), .B(p_input[2049]), .Z(n49445) );
  XNOR U49304 ( .A(n49489), .B(n49461), .Z(n49454) );
  XNOR U49305 ( .A(p_input[1455]), .B(n29033), .Z(n49461) );
  XOR U49306 ( .A(n49451), .B(n49460), .Z(n49489) );
  XOR U49307 ( .A(n49490), .B(n49457), .Z(n49460) );
  XOR U49308 ( .A(p_input[1453]), .B(p_input[2061]), .Z(n49457) );
  XOR U49309 ( .A(p_input[1454]), .B(n29035), .Z(n49490) );
  XOR U49310 ( .A(p_input[1449]), .B(p_input[2057]), .Z(n49451) );
  XOR U49311 ( .A(n49469), .B(n49467), .Z(n49449) );
  XNOR U49312 ( .A(n49491), .B(n49474), .Z(n49467) );
  XOR U49313 ( .A(p_input[1448]), .B(p_input[2056]), .Z(n49474) );
  XOR U49314 ( .A(n49464), .B(n49473), .Z(n49491) );
  XOR U49315 ( .A(n49492), .B(n49470), .Z(n49473) );
  XOR U49316 ( .A(p_input[1446]), .B(p_input[2054]), .Z(n49470) );
  XOR U49317 ( .A(p_input[1447]), .B(n30404), .Z(n49492) );
  XOR U49318 ( .A(p_input[1442]), .B(p_input[2050]), .Z(n49464) );
  XNOR U49319 ( .A(n49479), .B(n49478), .Z(n49469) );
  XOR U49320 ( .A(n49493), .B(n49475), .Z(n49478) );
  XOR U49321 ( .A(p_input[1443]), .B(p_input[2051]), .Z(n49475) );
  XOR U49322 ( .A(p_input[1444]), .B(n30406), .Z(n49493) );
  XOR U49323 ( .A(p_input[1445]), .B(p_input[2053]), .Z(n49479) );
  XNOR U49324 ( .A(n49494), .B(n49495), .Z(n49375) );
  AND U49325 ( .A(n1785), .B(n49496), .Z(n49495) );
  XNOR U49326 ( .A(n49497), .B(n49498), .Z(n1785) );
  AND U49327 ( .A(n49499), .B(n49500), .Z(n49498) );
  XOR U49328 ( .A(n49389), .B(n49497), .Z(n49500) );
  XNOR U49329 ( .A(n49501), .B(n49497), .Z(n49499) );
  XOR U49330 ( .A(n49502), .B(n49503), .Z(n49497) );
  AND U49331 ( .A(n49504), .B(n49505), .Z(n49503) );
  XOR U49332 ( .A(n49404), .B(n49502), .Z(n49505) );
  XOR U49333 ( .A(n49502), .B(n49405), .Z(n49504) );
  XOR U49334 ( .A(n49506), .B(n49507), .Z(n49502) );
  AND U49335 ( .A(n49508), .B(n49509), .Z(n49507) );
  XOR U49336 ( .A(n49432), .B(n49506), .Z(n49509) );
  XOR U49337 ( .A(n49506), .B(n49433), .Z(n49508) );
  XOR U49338 ( .A(n49510), .B(n49511), .Z(n49506) );
  AND U49339 ( .A(n49512), .B(n49513), .Z(n49511) );
  XOR U49340 ( .A(n49510), .B(n49483), .Z(n49513) );
  XNOR U49341 ( .A(n49514), .B(n49515), .Z(n49335) );
  AND U49342 ( .A(n1789), .B(n49516), .Z(n49515) );
  XNOR U49343 ( .A(n49517), .B(n49518), .Z(n1789) );
  AND U49344 ( .A(n49519), .B(n49520), .Z(n49518) );
  XOR U49345 ( .A(n49517), .B(n49345), .Z(n49520) );
  XNOR U49346 ( .A(n49517), .B(n49305), .Z(n49519) );
  XOR U49347 ( .A(n49521), .B(n49522), .Z(n49517) );
  AND U49348 ( .A(n49523), .B(n49524), .Z(n49522) );
  XOR U49349 ( .A(n49521), .B(n49313), .Z(n49523) );
  XOR U49350 ( .A(n49525), .B(n49526), .Z(n49296) );
  AND U49351 ( .A(n1793), .B(n49516), .Z(n49526) );
  XNOR U49352 ( .A(n49514), .B(n49525), .Z(n49516) );
  XNOR U49353 ( .A(n49527), .B(n49528), .Z(n1793) );
  AND U49354 ( .A(n49529), .B(n49530), .Z(n49528) );
  XNOR U49355 ( .A(n49531), .B(n49527), .Z(n49530) );
  IV U49356 ( .A(n49345), .Z(n49531) );
  XOR U49357 ( .A(n49501), .B(n49532), .Z(n49345) );
  AND U49358 ( .A(n1796), .B(n49533), .Z(n49532) );
  XOR U49359 ( .A(n49388), .B(n49385), .Z(n49533) );
  IV U49360 ( .A(n49501), .Z(n49388) );
  XNOR U49361 ( .A(n49305), .B(n49527), .Z(n49529) );
  XOR U49362 ( .A(n49534), .B(n49535), .Z(n49305) );
  AND U49363 ( .A(n1812), .B(n49536), .Z(n49535) );
  XOR U49364 ( .A(n49521), .B(n49537), .Z(n49527) );
  AND U49365 ( .A(n49538), .B(n49524), .Z(n49537) );
  XNOR U49366 ( .A(n49355), .B(n49521), .Z(n49524) );
  XOR U49367 ( .A(n49405), .B(n49539), .Z(n49355) );
  AND U49368 ( .A(n1796), .B(n49540), .Z(n49539) );
  XOR U49369 ( .A(n49401), .B(n49405), .Z(n49540) );
  XNOR U49370 ( .A(n49541), .B(n49521), .Z(n49538) );
  IV U49371 ( .A(n49313), .Z(n49541) );
  XOR U49372 ( .A(n49542), .B(n49543), .Z(n49313) );
  AND U49373 ( .A(n1812), .B(n49544), .Z(n49543) );
  XOR U49374 ( .A(n49545), .B(n49546), .Z(n49521) );
  AND U49375 ( .A(n49547), .B(n49548), .Z(n49546) );
  XNOR U49376 ( .A(n49365), .B(n49545), .Z(n49548) );
  XOR U49377 ( .A(n49433), .B(n49549), .Z(n49365) );
  AND U49378 ( .A(n1796), .B(n49550), .Z(n49549) );
  XOR U49379 ( .A(n49429), .B(n49433), .Z(n49550) );
  XOR U49380 ( .A(n49545), .B(n49322), .Z(n49547) );
  XOR U49381 ( .A(n49551), .B(n49552), .Z(n49322) );
  AND U49382 ( .A(n1812), .B(n49553), .Z(n49552) );
  XOR U49383 ( .A(n49554), .B(n49555), .Z(n49545) );
  AND U49384 ( .A(n49556), .B(n49557), .Z(n49555) );
  XNOR U49385 ( .A(n49554), .B(n49373), .Z(n49557) );
  XOR U49386 ( .A(n49484), .B(n49558), .Z(n49373) );
  AND U49387 ( .A(n1796), .B(n49559), .Z(n49558) );
  XOR U49388 ( .A(n49480), .B(n49484), .Z(n49559) );
  XNOR U49389 ( .A(n49560), .B(n49554), .Z(n49556) );
  IV U49390 ( .A(n49332), .Z(n49560) );
  XOR U49391 ( .A(n49561), .B(n49562), .Z(n49332) );
  AND U49392 ( .A(n1812), .B(n49563), .Z(n49562) );
  AND U49393 ( .A(n49525), .B(n49514), .Z(n49554) );
  XNOR U49394 ( .A(n49564), .B(n49565), .Z(n49514) );
  AND U49395 ( .A(n1796), .B(n49496), .Z(n49565) );
  XNOR U49396 ( .A(n49494), .B(n49564), .Z(n49496) );
  XNOR U49397 ( .A(n49566), .B(n49567), .Z(n1796) );
  AND U49398 ( .A(n49568), .B(n49569), .Z(n49567) );
  XNOR U49399 ( .A(n49566), .B(n49385), .Z(n49569) );
  IV U49400 ( .A(n49389), .Z(n49385) );
  XOR U49401 ( .A(n49570), .B(n49571), .Z(n49389) );
  AND U49402 ( .A(n1800), .B(n49572), .Z(n49571) );
  XOR U49403 ( .A(n49573), .B(n49570), .Z(n49572) );
  XNOR U49404 ( .A(n49566), .B(n49501), .Z(n49568) );
  XOR U49405 ( .A(n49574), .B(n49575), .Z(n49501) );
  AND U49406 ( .A(n1808), .B(n49536), .Z(n49575) );
  XOR U49407 ( .A(n49534), .B(n49574), .Z(n49536) );
  XOR U49408 ( .A(n49576), .B(n49577), .Z(n49566) );
  AND U49409 ( .A(n49578), .B(n49579), .Z(n49577) );
  XNOR U49410 ( .A(n49576), .B(n49401), .Z(n49579) );
  IV U49411 ( .A(n49404), .Z(n49401) );
  XOR U49412 ( .A(n49580), .B(n49581), .Z(n49404) );
  AND U49413 ( .A(n1800), .B(n49582), .Z(n49581) );
  XOR U49414 ( .A(n49583), .B(n49580), .Z(n49582) );
  XOR U49415 ( .A(n49405), .B(n49576), .Z(n49578) );
  XOR U49416 ( .A(n49584), .B(n49585), .Z(n49405) );
  AND U49417 ( .A(n1808), .B(n49544), .Z(n49585) );
  XOR U49418 ( .A(n49584), .B(n49542), .Z(n49544) );
  XOR U49419 ( .A(n49586), .B(n49587), .Z(n49576) );
  AND U49420 ( .A(n49588), .B(n49589), .Z(n49587) );
  XNOR U49421 ( .A(n49586), .B(n49429), .Z(n49589) );
  IV U49422 ( .A(n49432), .Z(n49429) );
  XOR U49423 ( .A(n49590), .B(n49591), .Z(n49432) );
  AND U49424 ( .A(n1800), .B(n49592), .Z(n49591) );
  XNOR U49425 ( .A(n49593), .B(n49590), .Z(n49592) );
  XOR U49426 ( .A(n49433), .B(n49586), .Z(n49588) );
  XOR U49427 ( .A(n49594), .B(n49595), .Z(n49433) );
  AND U49428 ( .A(n1808), .B(n49553), .Z(n49595) );
  XOR U49429 ( .A(n49594), .B(n49551), .Z(n49553) );
  XOR U49430 ( .A(n49510), .B(n49596), .Z(n49586) );
  AND U49431 ( .A(n49512), .B(n49597), .Z(n49596) );
  XNOR U49432 ( .A(n49510), .B(n49480), .Z(n49597) );
  IV U49433 ( .A(n49483), .Z(n49480) );
  XOR U49434 ( .A(n49598), .B(n49599), .Z(n49483) );
  AND U49435 ( .A(n1800), .B(n49600), .Z(n49599) );
  XOR U49436 ( .A(n49601), .B(n49598), .Z(n49600) );
  XOR U49437 ( .A(n49484), .B(n49510), .Z(n49512) );
  XOR U49438 ( .A(n49602), .B(n49603), .Z(n49484) );
  AND U49439 ( .A(n1808), .B(n49563), .Z(n49603) );
  XOR U49440 ( .A(n49602), .B(n49561), .Z(n49563) );
  AND U49441 ( .A(n49564), .B(n49494), .Z(n49510) );
  XNOR U49442 ( .A(n49604), .B(n49605), .Z(n49494) );
  AND U49443 ( .A(n1800), .B(n49606), .Z(n49605) );
  XNOR U49444 ( .A(n49607), .B(n49604), .Z(n49606) );
  XNOR U49445 ( .A(n49608), .B(n49609), .Z(n1800) );
  AND U49446 ( .A(n49610), .B(n49611), .Z(n49609) );
  XOR U49447 ( .A(n49573), .B(n49608), .Z(n49611) );
  AND U49448 ( .A(n49612), .B(n49613), .Z(n49573) );
  XNOR U49449 ( .A(n49570), .B(n49608), .Z(n49610) );
  XNOR U49450 ( .A(n49614), .B(n49615), .Z(n49570) );
  AND U49451 ( .A(n1804), .B(n49616), .Z(n49615) );
  XNOR U49452 ( .A(n49617), .B(n49618), .Z(n49616) );
  XOR U49453 ( .A(n49619), .B(n49620), .Z(n49608) );
  AND U49454 ( .A(n49621), .B(n49622), .Z(n49620) );
  XNOR U49455 ( .A(n49619), .B(n49612), .Z(n49622) );
  IV U49456 ( .A(n49583), .Z(n49612) );
  XOR U49457 ( .A(n49623), .B(n49624), .Z(n49583) );
  XOR U49458 ( .A(n49625), .B(n49613), .Z(n49624) );
  AND U49459 ( .A(n49593), .B(n49626), .Z(n49613) );
  AND U49460 ( .A(n49627), .B(n49628), .Z(n49625) );
  XOR U49461 ( .A(n49629), .B(n49623), .Z(n49627) );
  XNOR U49462 ( .A(n49580), .B(n49619), .Z(n49621) );
  XNOR U49463 ( .A(n49630), .B(n49631), .Z(n49580) );
  AND U49464 ( .A(n1804), .B(n49632), .Z(n49631) );
  XNOR U49465 ( .A(n49633), .B(n49634), .Z(n49632) );
  XOR U49466 ( .A(n49635), .B(n49636), .Z(n49619) );
  AND U49467 ( .A(n49637), .B(n49638), .Z(n49636) );
  XNOR U49468 ( .A(n49635), .B(n49593), .Z(n49638) );
  XOR U49469 ( .A(n49639), .B(n49628), .Z(n49593) );
  XNOR U49470 ( .A(n49640), .B(n49623), .Z(n49628) );
  XOR U49471 ( .A(n49641), .B(n49642), .Z(n49623) );
  AND U49472 ( .A(n49643), .B(n49644), .Z(n49642) );
  XOR U49473 ( .A(n49645), .B(n49641), .Z(n49643) );
  XNOR U49474 ( .A(n49646), .B(n49647), .Z(n49640) );
  AND U49475 ( .A(n49648), .B(n49649), .Z(n49647) );
  XOR U49476 ( .A(n49646), .B(n49650), .Z(n49648) );
  XNOR U49477 ( .A(n49629), .B(n49626), .Z(n49639) );
  AND U49478 ( .A(n49651), .B(n49652), .Z(n49626) );
  XOR U49479 ( .A(n49653), .B(n49654), .Z(n49629) );
  AND U49480 ( .A(n49655), .B(n49656), .Z(n49654) );
  XOR U49481 ( .A(n49653), .B(n49657), .Z(n49655) );
  XNOR U49482 ( .A(n49590), .B(n49635), .Z(n49637) );
  XNOR U49483 ( .A(n49658), .B(n49659), .Z(n49590) );
  AND U49484 ( .A(n1804), .B(n49660), .Z(n49659) );
  XNOR U49485 ( .A(n49661), .B(n49662), .Z(n49660) );
  XOR U49486 ( .A(n49663), .B(n49664), .Z(n49635) );
  AND U49487 ( .A(n49665), .B(n49666), .Z(n49664) );
  XNOR U49488 ( .A(n49663), .B(n49651), .Z(n49666) );
  IV U49489 ( .A(n49601), .Z(n49651) );
  XNOR U49490 ( .A(n49667), .B(n49644), .Z(n49601) );
  XNOR U49491 ( .A(n49668), .B(n49650), .Z(n49644) );
  XNOR U49492 ( .A(n49669), .B(n49670), .Z(n49650) );
  NOR U49493 ( .A(n49671), .B(n49672), .Z(n49670) );
  XOR U49494 ( .A(n49669), .B(n49673), .Z(n49671) );
  XNOR U49495 ( .A(n49649), .B(n49641), .Z(n49668) );
  XOR U49496 ( .A(n49674), .B(n49675), .Z(n49641) );
  AND U49497 ( .A(n49676), .B(n49677), .Z(n49675) );
  XOR U49498 ( .A(n49674), .B(n49678), .Z(n49676) );
  XNOR U49499 ( .A(n49679), .B(n49646), .Z(n49649) );
  XOR U49500 ( .A(n49680), .B(n49681), .Z(n49646) );
  AND U49501 ( .A(n49682), .B(n49683), .Z(n49681) );
  XNOR U49502 ( .A(n49684), .B(n49685), .Z(n49682) );
  IV U49503 ( .A(n49680), .Z(n49684) );
  XNOR U49504 ( .A(n49686), .B(n49687), .Z(n49679) );
  NOR U49505 ( .A(n49688), .B(n49689), .Z(n49687) );
  XNOR U49506 ( .A(n49686), .B(n49690), .Z(n49688) );
  XNOR U49507 ( .A(n49645), .B(n49652), .Z(n49667) );
  NOR U49508 ( .A(n49607), .B(n49691), .Z(n49652) );
  XOR U49509 ( .A(n49657), .B(n49656), .Z(n49645) );
  XNOR U49510 ( .A(n49692), .B(n49653), .Z(n49656) );
  XOR U49511 ( .A(n49693), .B(n49694), .Z(n49653) );
  AND U49512 ( .A(n49695), .B(n49696), .Z(n49694) );
  XNOR U49513 ( .A(n49697), .B(n49698), .Z(n49695) );
  IV U49514 ( .A(n49693), .Z(n49697) );
  XNOR U49515 ( .A(n49699), .B(n49700), .Z(n49692) );
  NOR U49516 ( .A(n49701), .B(n49702), .Z(n49700) );
  XNOR U49517 ( .A(n49699), .B(n49703), .Z(n49701) );
  XOR U49518 ( .A(n49704), .B(n49705), .Z(n49657) );
  NOR U49519 ( .A(n49706), .B(n49707), .Z(n49705) );
  XNOR U49520 ( .A(n49704), .B(n49708), .Z(n49706) );
  XNOR U49521 ( .A(n49598), .B(n49663), .Z(n49665) );
  XNOR U49522 ( .A(n49709), .B(n49710), .Z(n49598) );
  AND U49523 ( .A(n1804), .B(n49711), .Z(n49710) );
  XNOR U49524 ( .A(n49712), .B(n49713), .Z(n49711) );
  AND U49525 ( .A(n49604), .B(n49607), .Z(n49663) );
  XOR U49526 ( .A(n49714), .B(n49691), .Z(n49607) );
  XNOR U49527 ( .A(p_input[1456]), .B(p_input[2048]), .Z(n49691) );
  XNOR U49528 ( .A(n49678), .B(n49677), .Z(n49714) );
  XNOR U49529 ( .A(n49715), .B(n49685), .Z(n49677) );
  XNOR U49530 ( .A(n49673), .B(n49672), .Z(n49685) );
  XNOR U49531 ( .A(n49716), .B(n49669), .Z(n49672) );
  XNOR U49532 ( .A(p_input[1466]), .B(p_input[2058]), .Z(n49669) );
  XOR U49533 ( .A(p_input[1467]), .B(n29030), .Z(n49716) );
  XOR U49534 ( .A(p_input[1468]), .B(p_input[2060]), .Z(n49673) );
  XOR U49535 ( .A(n49683), .B(n49717), .Z(n49715) );
  IV U49536 ( .A(n49674), .Z(n49717) );
  XOR U49537 ( .A(p_input[1457]), .B(p_input[2049]), .Z(n49674) );
  XNOR U49538 ( .A(n49718), .B(n49690), .Z(n49683) );
  XNOR U49539 ( .A(p_input[1471]), .B(n29033), .Z(n49690) );
  XOR U49540 ( .A(n49680), .B(n49689), .Z(n49718) );
  XOR U49541 ( .A(n49719), .B(n49686), .Z(n49689) );
  XOR U49542 ( .A(p_input[1469]), .B(p_input[2061]), .Z(n49686) );
  XOR U49543 ( .A(p_input[1470]), .B(n29035), .Z(n49719) );
  XOR U49544 ( .A(p_input[1465]), .B(p_input[2057]), .Z(n49680) );
  XOR U49545 ( .A(n49698), .B(n49696), .Z(n49678) );
  XNOR U49546 ( .A(n49720), .B(n49703), .Z(n49696) );
  XOR U49547 ( .A(p_input[1464]), .B(p_input[2056]), .Z(n49703) );
  XOR U49548 ( .A(n49693), .B(n49702), .Z(n49720) );
  XOR U49549 ( .A(n49721), .B(n49699), .Z(n49702) );
  XOR U49550 ( .A(p_input[1462]), .B(p_input[2054]), .Z(n49699) );
  XOR U49551 ( .A(p_input[1463]), .B(n30404), .Z(n49721) );
  XOR U49552 ( .A(p_input[1458]), .B(p_input[2050]), .Z(n49693) );
  XNOR U49553 ( .A(n49708), .B(n49707), .Z(n49698) );
  XOR U49554 ( .A(n49722), .B(n49704), .Z(n49707) );
  XOR U49555 ( .A(p_input[1459]), .B(p_input[2051]), .Z(n49704) );
  XOR U49556 ( .A(p_input[1460]), .B(n30406), .Z(n49722) );
  XOR U49557 ( .A(p_input[1461]), .B(p_input[2053]), .Z(n49708) );
  XNOR U49558 ( .A(n49723), .B(n49724), .Z(n49604) );
  AND U49559 ( .A(n1804), .B(n49725), .Z(n49724) );
  XNOR U49560 ( .A(n49726), .B(n49727), .Z(n1804) );
  AND U49561 ( .A(n49728), .B(n49729), .Z(n49727) );
  XOR U49562 ( .A(n49618), .B(n49726), .Z(n49729) );
  XNOR U49563 ( .A(n49730), .B(n49726), .Z(n49728) );
  XOR U49564 ( .A(n49731), .B(n49732), .Z(n49726) );
  AND U49565 ( .A(n49733), .B(n49734), .Z(n49732) );
  XOR U49566 ( .A(n49633), .B(n49731), .Z(n49734) );
  XOR U49567 ( .A(n49731), .B(n49634), .Z(n49733) );
  XOR U49568 ( .A(n49735), .B(n49736), .Z(n49731) );
  AND U49569 ( .A(n49737), .B(n49738), .Z(n49736) );
  XOR U49570 ( .A(n49661), .B(n49735), .Z(n49738) );
  XOR U49571 ( .A(n49735), .B(n49662), .Z(n49737) );
  XOR U49572 ( .A(n49739), .B(n49740), .Z(n49735) );
  AND U49573 ( .A(n49741), .B(n49742), .Z(n49740) );
  XOR U49574 ( .A(n49739), .B(n49712), .Z(n49742) );
  XNOR U49575 ( .A(n49743), .B(n49744), .Z(n49564) );
  AND U49576 ( .A(n1808), .B(n49745), .Z(n49744) );
  XNOR U49577 ( .A(n49746), .B(n49747), .Z(n1808) );
  AND U49578 ( .A(n49748), .B(n49749), .Z(n49747) );
  XOR U49579 ( .A(n49746), .B(n49574), .Z(n49749) );
  XNOR U49580 ( .A(n49746), .B(n49534), .Z(n49748) );
  XOR U49581 ( .A(n49750), .B(n49751), .Z(n49746) );
  AND U49582 ( .A(n49752), .B(n49753), .Z(n49751) );
  XOR U49583 ( .A(n49750), .B(n49542), .Z(n49752) );
  XOR U49584 ( .A(n49754), .B(n49755), .Z(n49525) );
  AND U49585 ( .A(n1812), .B(n49745), .Z(n49755) );
  XNOR U49586 ( .A(n49743), .B(n49754), .Z(n49745) );
  XNOR U49587 ( .A(n49756), .B(n49757), .Z(n1812) );
  AND U49588 ( .A(n49758), .B(n49759), .Z(n49757) );
  XNOR U49589 ( .A(n49760), .B(n49756), .Z(n49759) );
  IV U49590 ( .A(n49574), .Z(n49760) );
  XOR U49591 ( .A(n49730), .B(n49761), .Z(n49574) );
  AND U49592 ( .A(n1815), .B(n49762), .Z(n49761) );
  XOR U49593 ( .A(n49617), .B(n49614), .Z(n49762) );
  IV U49594 ( .A(n49730), .Z(n49617) );
  XNOR U49595 ( .A(n49534), .B(n49756), .Z(n49758) );
  XOR U49596 ( .A(n49763), .B(n49764), .Z(n49534) );
  AND U49597 ( .A(n1831), .B(n49765), .Z(n49764) );
  XOR U49598 ( .A(n49750), .B(n49766), .Z(n49756) );
  AND U49599 ( .A(n49767), .B(n49753), .Z(n49766) );
  XNOR U49600 ( .A(n49584), .B(n49750), .Z(n49753) );
  XOR U49601 ( .A(n49634), .B(n49768), .Z(n49584) );
  AND U49602 ( .A(n1815), .B(n49769), .Z(n49768) );
  XOR U49603 ( .A(n49630), .B(n49634), .Z(n49769) );
  XNOR U49604 ( .A(n49770), .B(n49750), .Z(n49767) );
  IV U49605 ( .A(n49542), .Z(n49770) );
  XOR U49606 ( .A(n49771), .B(n49772), .Z(n49542) );
  AND U49607 ( .A(n1831), .B(n49773), .Z(n49772) );
  XOR U49608 ( .A(n49774), .B(n49775), .Z(n49750) );
  AND U49609 ( .A(n49776), .B(n49777), .Z(n49775) );
  XNOR U49610 ( .A(n49594), .B(n49774), .Z(n49777) );
  XOR U49611 ( .A(n49662), .B(n49778), .Z(n49594) );
  AND U49612 ( .A(n1815), .B(n49779), .Z(n49778) );
  XOR U49613 ( .A(n49658), .B(n49662), .Z(n49779) );
  XOR U49614 ( .A(n49774), .B(n49551), .Z(n49776) );
  XOR U49615 ( .A(n49780), .B(n49781), .Z(n49551) );
  AND U49616 ( .A(n1831), .B(n49782), .Z(n49781) );
  XOR U49617 ( .A(n49783), .B(n49784), .Z(n49774) );
  AND U49618 ( .A(n49785), .B(n49786), .Z(n49784) );
  XNOR U49619 ( .A(n49783), .B(n49602), .Z(n49786) );
  XOR U49620 ( .A(n49713), .B(n49787), .Z(n49602) );
  AND U49621 ( .A(n1815), .B(n49788), .Z(n49787) );
  XOR U49622 ( .A(n49709), .B(n49713), .Z(n49788) );
  XNOR U49623 ( .A(n49789), .B(n49783), .Z(n49785) );
  IV U49624 ( .A(n49561), .Z(n49789) );
  XOR U49625 ( .A(n49790), .B(n49791), .Z(n49561) );
  AND U49626 ( .A(n1831), .B(n49792), .Z(n49791) );
  AND U49627 ( .A(n49754), .B(n49743), .Z(n49783) );
  XNOR U49628 ( .A(n49793), .B(n49794), .Z(n49743) );
  AND U49629 ( .A(n1815), .B(n49725), .Z(n49794) );
  XNOR U49630 ( .A(n49723), .B(n49793), .Z(n49725) );
  XNOR U49631 ( .A(n49795), .B(n49796), .Z(n1815) );
  AND U49632 ( .A(n49797), .B(n49798), .Z(n49796) );
  XNOR U49633 ( .A(n49795), .B(n49614), .Z(n49798) );
  IV U49634 ( .A(n49618), .Z(n49614) );
  XOR U49635 ( .A(n49799), .B(n49800), .Z(n49618) );
  AND U49636 ( .A(n1819), .B(n49801), .Z(n49800) );
  XOR U49637 ( .A(n49802), .B(n49799), .Z(n49801) );
  XNOR U49638 ( .A(n49795), .B(n49730), .Z(n49797) );
  XOR U49639 ( .A(n49803), .B(n49804), .Z(n49730) );
  AND U49640 ( .A(n1827), .B(n49765), .Z(n49804) );
  XOR U49641 ( .A(n49763), .B(n49803), .Z(n49765) );
  XOR U49642 ( .A(n49805), .B(n49806), .Z(n49795) );
  AND U49643 ( .A(n49807), .B(n49808), .Z(n49806) );
  XNOR U49644 ( .A(n49805), .B(n49630), .Z(n49808) );
  IV U49645 ( .A(n49633), .Z(n49630) );
  XOR U49646 ( .A(n49809), .B(n49810), .Z(n49633) );
  AND U49647 ( .A(n1819), .B(n49811), .Z(n49810) );
  XOR U49648 ( .A(n49812), .B(n49809), .Z(n49811) );
  XOR U49649 ( .A(n49634), .B(n49805), .Z(n49807) );
  XOR U49650 ( .A(n49813), .B(n49814), .Z(n49634) );
  AND U49651 ( .A(n1827), .B(n49773), .Z(n49814) );
  XOR U49652 ( .A(n49813), .B(n49771), .Z(n49773) );
  XOR U49653 ( .A(n49815), .B(n49816), .Z(n49805) );
  AND U49654 ( .A(n49817), .B(n49818), .Z(n49816) );
  XNOR U49655 ( .A(n49815), .B(n49658), .Z(n49818) );
  IV U49656 ( .A(n49661), .Z(n49658) );
  XOR U49657 ( .A(n49819), .B(n49820), .Z(n49661) );
  AND U49658 ( .A(n1819), .B(n49821), .Z(n49820) );
  XNOR U49659 ( .A(n49822), .B(n49819), .Z(n49821) );
  XOR U49660 ( .A(n49662), .B(n49815), .Z(n49817) );
  XOR U49661 ( .A(n49823), .B(n49824), .Z(n49662) );
  AND U49662 ( .A(n1827), .B(n49782), .Z(n49824) );
  XOR U49663 ( .A(n49823), .B(n49780), .Z(n49782) );
  XOR U49664 ( .A(n49739), .B(n49825), .Z(n49815) );
  AND U49665 ( .A(n49741), .B(n49826), .Z(n49825) );
  XNOR U49666 ( .A(n49739), .B(n49709), .Z(n49826) );
  IV U49667 ( .A(n49712), .Z(n49709) );
  XOR U49668 ( .A(n49827), .B(n49828), .Z(n49712) );
  AND U49669 ( .A(n1819), .B(n49829), .Z(n49828) );
  XOR U49670 ( .A(n49830), .B(n49827), .Z(n49829) );
  XOR U49671 ( .A(n49713), .B(n49739), .Z(n49741) );
  XOR U49672 ( .A(n49831), .B(n49832), .Z(n49713) );
  AND U49673 ( .A(n1827), .B(n49792), .Z(n49832) );
  XOR U49674 ( .A(n49831), .B(n49790), .Z(n49792) );
  AND U49675 ( .A(n49793), .B(n49723), .Z(n49739) );
  XNOR U49676 ( .A(n49833), .B(n49834), .Z(n49723) );
  AND U49677 ( .A(n1819), .B(n49835), .Z(n49834) );
  XNOR U49678 ( .A(n49836), .B(n49833), .Z(n49835) );
  XNOR U49679 ( .A(n49837), .B(n49838), .Z(n1819) );
  AND U49680 ( .A(n49839), .B(n49840), .Z(n49838) );
  XOR U49681 ( .A(n49802), .B(n49837), .Z(n49840) );
  AND U49682 ( .A(n49841), .B(n49842), .Z(n49802) );
  XNOR U49683 ( .A(n49799), .B(n49837), .Z(n49839) );
  XNOR U49684 ( .A(n49843), .B(n49844), .Z(n49799) );
  AND U49685 ( .A(n1823), .B(n49845), .Z(n49844) );
  XNOR U49686 ( .A(n49846), .B(n49847), .Z(n49845) );
  XOR U49687 ( .A(n49848), .B(n49849), .Z(n49837) );
  AND U49688 ( .A(n49850), .B(n49851), .Z(n49849) );
  XNOR U49689 ( .A(n49848), .B(n49841), .Z(n49851) );
  IV U49690 ( .A(n49812), .Z(n49841) );
  XOR U49691 ( .A(n49852), .B(n49853), .Z(n49812) );
  XOR U49692 ( .A(n49854), .B(n49842), .Z(n49853) );
  AND U49693 ( .A(n49822), .B(n49855), .Z(n49842) );
  AND U49694 ( .A(n49856), .B(n49857), .Z(n49854) );
  XOR U49695 ( .A(n49858), .B(n49852), .Z(n49856) );
  XNOR U49696 ( .A(n49809), .B(n49848), .Z(n49850) );
  XNOR U49697 ( .A(n49859), .B(n49860), .Z(n49809) );
  AND U49698 ( .A(n1823), .B(n49861), .Z(n49860) );
  XNOR U49699 ( .A(n49862), .B(n49863), .Z(n49861) );
  XOR U49700 ( .A(n49864), .B(n49865), .Z(n49848) );
  AND U49701 ( .A(n49866), .B(n49867), .Z(n49865) );
  XNOR U49702 ( .A(n49864), .B(n49822), .Z(n49867) );
  XOR U49703 ( .A(n49868), .B(n49857), .Z(n49822) );
  XNOR U49704 ( .A(n49869), .B(n49852), .Z(n49857) );
  XOR U49705 ( .A(n49870), .B(n49871), .Z(n49852) );
  AND U49706 ( .A(n49872), .B(n49873), .Z(n49871) );
  XOR U49707 ( .A(n49874), .B(n49870), .Z(n49872) );
  XNOR U49708 ( .A(n49875), .B(n49876), .Z(n49869) );
  AND U49709 ( .A(n49877), .B(n49878), .Z(n49876) );
  XOR U49710 ( .A(n49875), .B(n49879), .Z(n49877) );
  XNOR U49711 ( .A(n49858), .B(n49855), .Z(n49868) );
  AND U49712 ( .A(n49880), .B(n49881), .Z(n49855) );
  XOR U49713 ( .A(n49882), .B(n49883), .Z(n49858) );
  AND U49714 ( .A(n49884), .B(n49885), .Z(n49883) );
  XOR U49715 ( .A(n49882), .B(n49886), .Z(n49884) );
  XNOR U49716 ( .A(n49819), .B(n49864), .Z(n49866) );
  XNOR U49717 ( .A(n49887), .B(n49888), .Z(n49819) );
  AND U49718 ( .A(n1823), .B(n49889), .Z(n49888) );
  XNOR U49719 ( .A(n49890), .B(n49891), .Z(n49889) );
  XOR U49720 ( .A(n49892), .B(n49893), .Z(n49864) );
  AND U49721 ( .A(n49894), .B(n49895), .Z(n49893) );
  XNOR U49722 ( .A(n49892), .B(n49880), .Z(n49895) );
  IV U49723 ( .A(n49830), .Z(n49880) );
  XNOR U49724 ( .A(n49896), .B(n49873), .Z(n49830) );
  XNOR U49725 ( .A(n49897), .B(n49879), .Z(n49873) );
  XNOR U49726 ( .A(n49898), .B(n49899), .Z(n49879) );
  NOR U49727 ( .A(n49900), .B(n49901), .Z(n49899) );
  XOR U49728 ( .A(n49898), .B(n49902), .Z(n49900) );
  XNOR U49729 ( .A(n49878), .B(n49870), .Z(n49897) );
  XOR U49730 ( .A(n49903), .B(n49904), .Z(n49870) );
  AND U49731 ( .A(n49905), .B(n49906), .Z(n49904) );
  XOR U49732 ( .A(n49903), .B(n49907), .Z(n49905) );
  XNOR U49733 ( .A(n49908), .B(n49875), .Z(n49878) );
  XOR U49734 ( .A(n49909), .B(n49910), .Z(n49875) );
  AND U49735 ( .A(n49911), .B(n49912), .Z(n49910) );
  XNOR U49736 ( .A(n49913), .B(n49914), .Z(n49911) );
  IV U49737 ( .A(n49909), .Z(n49913) );
  XNOR U49738 ( .A(n49915), .B(n49916), .Z(n49908) );
  NOR U49739 ( .A(n49917), .B(n49918), .Z(n49916) );
  XNOR U49740 ( .A(n49915), .B(n49919), .Z(n49917) );
  XNOR U49741 ( .A(n49874), .B(n49881), .Z(n49896) );
  NOR U49742 ( .A(n49836), .B(n49920), .Z(n49881) );
  XOR U49743 ( .A(n49886), .B(n49885), .Z(n49874) );
  XNOR U49744 ( .A(n49921), .B(n49882), .Z(n49885) );
  XOR U49745 ( .A(n49922), .B(n49923), .Z(n49882) );
  AND U49746 ( .A(n49924), .B(n49925), .Z(n49923) );
  XNOR U49747 ( .A(n49926), .B(n49927), .Z(n49924) );
  IV U49748 ( .A(n49922), .Z(n49926) );
  XNOR U49749 ( .A(n49928), .B(n49929), .Z(n49921) );
  NOR U49750 ( .A(n49930), .B(n49931), .Z(n49929) );
  XNOR U49751 ( .A(n49928), .B(n49932), .Z(n49930) );
  XOR U49752 ( .A(n49933), .B(n49934), .Z(n49886) );
  NOR U49753 ( .A(n49935), .B(n49936), .Z(n49934) );
  XNOR U49754 ( .A(n49933), .B(n49937), .Z(n49935) );
  XNOR U49755 ( .A(n49827), .B(n49892), .Z(n49894) );
  XNOR U49756 ( .A(n49938), .B(n49939), .Z(n49827) );
  AND U49757 ( .A(n1823), .B(n49940), .Z(n49939) );
  XNOR U49758 ( .A(n49941), .B(n49942), .Z(n49940) );
  AND U49759 ( .A(n49833), .B(n49836), .Z(n49892) );
  XOR U49760 ( .A(n49943), .B(n49920), .Z(n49836) );
  XNOR U49761 ( .A(p_input[1472]), .B(p_input[2048]), .Z(n49920) );
  XNOR U49762 ( .A(n49907), .B(n49906), .Z(n49943) );
  XNOR U49763 ( .A(n49944), .B(n49914), .Z(n49906) );
  XNOR U49764 ( .A(n49902), .B(n49901), .Z(n49914) );
  XNOR U49765 ( .A(n49945), .B(n49898), .Z(n49901) );
  XNOR U49766 ( .A(p_input[1482]), .B(p_input[2058]), .Z(n49898) );
  XOR U49767 ( .A(p_input[1483]), .B(n29030), .Z(n49945) );
  XOR U49768 ( .A(p_input[1484]), .B(p_input[2060]), .Z(n49902) );
  XOR U49769 ( .A(n49912), .B(n49946), .Z(n49944) );
  IV U49770 ( .A(n49903), .Z(n49946) );
  XOR U49771 ( .A(p_input[1473]), .B(p_input[2049]), .Z(n49903) );
  XNOR U49772 ( .A(n49947), .B(n49919), .Z(n49912) );
  XNOR U49773 ( .A(p_input[1487]), .B(n29033), .Z(n49919) );
  XOR U49774 ( .A(n49909), .B(n49918), .Z(n49947) );
  XOR U49775 ( .A(n49948), .B(n49915), .Z(n49918) );
  XOR U49776 ( .A(p_input[1485]), .B(p_input[2061]), .Z(n49915) );
  XOR U49777 ( .A(p_input[1486]), .B(n29035), .Z(n49948) );
  XOR U49778 ( .A(p_input[1481]), .B(p_input[2057]), .Z(n49909) );
  XOR U49779 ( .A(n49927), .B(n49925), .Z(n49907) );
  XNOR U49780 ( .A(n49949), .B(n49932), .Z(n49925) );
  XOR U49781 ( .A(p_input[1480]), .B(p_input[2056]), .Z(n49932) );
  XOR U49782 ( .A(n49922), .B(n49931), .Z(n49949) );
  XOR U49783 ( .A(n49950), .B(n49928), .Z(n49931) );
  XOR U49784 ( .A(p_input[1478]), .B(p_input[2054]), .Z(n49928) );
  XOR U49785 ( .A(p_input[1479]), .B(n30404), .Z(n49950) );
  XOR U49786 ( .A(p_input[1474]), .B(p_input[2050]), .Z(n49922) );
  XNOR U49787 ( .A(n49937), .B(n49936), .Z(n49927) );
  XOR U49788 ( .A(n49951), .B(n49933), .Z(n49936) );
  XOR U49789 ( .A(p_input[1475]), .B(p_input[2051]), .Z(n49933) );
  XOR U49790 ( .A(p_input[1476]), .B(n30406), .Z(n49951) );
  XOR U49791 ( .A(p_input[1477]), .B(p_input[2053]), .Z(n49937) );
  XNOR U49792 ( .A(n49952), .B(n49953), .Z(n49833) );
  AND U49793 ( .A(n1823), .B(n49954), .Z(n49953) );
  XNOR U49794 ( .A(n49955), .B(n49956), .Z(n1823) );
  AND U49795 ( .A(n49957), .B(n49958), .Z(n49956) );
  XOR U49796 ( .A(n49847), .B(n49955), .Z(n49958) );
  XNOR U49797 ( .A(n49959), .B(n49955), .Z(n49957) );
  XOR U49798 ( .A(n49960), .B(n49961), .Z(n49955) );
  AND U49799 ( .A(n49962), .B(n49963), .Z(n49961) );
  XOR U49800 ( .A(n49862), .B(n49960), .Z(n49963) );
  XOR U49801 ( .A(n49960), .B(n49863), .Z(n49962) );
  XOR U49802 ( .A(n49964), .B(n49965), .Z(n49960) );
  AND U49803 ( .A(n49966), .B(n49967), .Z(n49965) );
  XOR U49804 ( .A(n49890), .B(n49964), .Z(n49967) );
  XOR U49805 ( .A(n49964), .B(n49891), .Z(n49966) );
  XOR U49806 ( .A(n49968), .B(n49969), .Z(n49964) );
  AND U49807 ( .A(n49970), .B(n49971), .Z(n49969) );
  XOR U49808 ( .A(n49968), .B(n49941), .Z(n49971) );
  XNOR U49809 ( .A(n49972), .B(n49973), .Z(n49793) );
  AND U49810 ( .A(n1827), .B(n49974), .Z(n49973) );
  XNOR U49811 ( .A(n49975), .B(n49976), .Z(n1827) );
  AND U49812 ( .A(n49977), .B(n49978), .Z(n49976) );
  XOR U49813 ( .A(n49975), .B(n49803), .Z(n49978) );
  XNOR U49814 ( .A(n49975), .B(n49763), .Z(n49977) );
  XOR U49815 ( .A(n49979), .B(n49980), .Z(n49975) );
  AND U49816 ( .A(n49981), .B(n49982), .Z(n49980) );
  XOR U49817 ( .A(n49979), .B(n49771), .Z(n49981) );
  XOR U49818 ( .A(n49983), .B(n49984), .Z(n49754) );
  AND U49819 ( .A(n1831), .B(n49974), .Z(n49984) );
  XNOR U49820 ( .A(n49972), .B(n49983), .Z(n49974) );
  XNOR U49821 ( .A(n49985), .B(n49986), .Z(n1831) );
  AND U49822 ( .A(n49987), .B(n49988), .Z(n49986) );
  XNOR U49823 ( .A(n49989), .B(n49985), .Z(n49988) );
  IV U49824 ( .A(n49803), .Z(n49989) );
  XOR U49825 ( .A(n49959), .B(n49990), .Z(n49803) );
  AND U49826 ( .A(n1834), .B(n49991), .Z(n49990) );
  XOR U49827 ( .A(n49846), .B(n49843), .Z(n49991) );
  IV U49828 ( .A(n49959), .Z(n49846) );
  XNOR U49829 ( .A(n49763), .B(n49985), .Z(n49987) );
  XOR U49830 ( .A(n49992), .B(n49993), .Z(n49763) );
  AND U49831 ( .A(n1850), .B(n49994), .Z(n49993) );
  XOR U49832 ( .A(n49979), .B(n49995), .Z(n49985) );
  AND U49833 ( .A(n49996), .B(n49982), .Z(n49995) );
  XNOR U49834 ( .A(n49813), .B(n49979), .Z(n49982) );
  XOR U49835 ( .A(n49863), .B(n49997), .Z(n49813) );
  AND U49836 ( .A(n1834), .B(n49998), .Z(n49997) );
  XOR U49837 ( .A(n49859), .B(n49863), .Z(n49998) );
  XNOR U49838 ( .A(n49999), .B(n49979), .Z(n49996) );
  IV U49839 ( .A(n49771), .Z(n49999) );
  XOR U49840 ( .A(n50000), .B(n50001), .Z(n49771) );
  AND U49841 ( .A(n1850), .B(n50002), .Z(n50001) );
  XOR U49842 ( .A(n50003), .B(n50004), .Z(n49979) );
  AND U49843 ( .A(n50005), .B(n50006), .Z(n50004) );
  XNOR U49844 ( .A(n49823), .B(n50003), .Z(n50006) );
  XOR U49845 ( .A(n49891), .B(n50007), .Z(n49823) );
  AND U49846 ( .A(n1834), .B(n50008), .Z(n50007) );
  XOR U49847 ( .A(n49887), .B(n49891), .Z(n50008) );
  XOR U49848 ( .A(n50003), .B(n49780), .Z(n50005) );
  XOR U49849 ( .A(n50009), .B(n50010), .Z(n49780) );
  AND U49850 ( .A(n1850), .B(n50011), .Z(n50010) );
  XOR U49851 ( .A(n50012), .B(n50013), .Z(n50003) );
  AND U49852 ( .A(n50014), .B(n50015), .Z(n50013) );
  XNOR U49853 ( .A(n50012), .B(n49831), .Z(n50015) );
  XOR U49854 ( .A(n49942), .B(n50016), .Z(n49831) );
  AND U49855 ( .A(n1834), .B(n50017), .Z(n50016) );
  XOR U49856 ( .A(n49938), .B(n49942), .Z(n50017) );
  XNOR U49857 ( .A(n50018), .B(n50012), .Z(n50014) );
  IV U49858 ( .A(n49790), .Z(n50018) );
  XOR U49859 ( .A(n50019), .B(n50020), .Z(n49790) );
  AND U49860 ( .A(n1850), .B(n50021), .Z(n50020) );
  AND U49861 ( .A(n49983), .B(n49972), .Z(n50012) );
  XNOR U49862 ( .A(n50022), .B(n50023), .Z(n49972) );
  AND U49863 ( .A(n1834), .B(n49954), .Z(n50023) );
  XNOR U49864 ( .A(n49952), .B(n50022), .Z(n49954) );
  XNOR U49865 ( .A(n50024), .B(n50025), .Z(n1834) );
  AND U49866 ( .A(n50026), .B(n50027), .Z(n50025) );
  XNOR U49867 ( .A(n50024), .B(n49843), .Z(n50027) );
  IV U49868 ( .A(n49847), .Z(n49843) );
  XOR U49869 ( .A(n50028), .B(n50029), .Z(n49847) );
  AND U49870 ( .A(n1838), .B(n50030), .Z(n50029) );
  XOR U49871 ( .A(n50031), .B(n50028), .Z(n50030) );
  XNOR U49872 ( .A(n50024), .B(n49959), .Z(n50026) );
  XOR U49873 ( .A(n50032), .B(n50033), .Z(n49959) );
  AND U49874 ( .A(n1846), .B(n49994), .Z(n50033) );
  XOR U49875 ( .A(n49992), .B(n50032), .Z(n49994) );
  XOR U49876 ( .A(n50034), .B(n50035), .Z(n50024) );
  AND U49877 ( .A(n50036), .B(n50037), .Z(n50035) );
  XNOR U49878 ( .A(n50034), .B(n49859), .Z(n50037) );
  IV U49879 ( .A(n49862), .Z(n49859) );
  XOR U49880 ( .A(n50038), .B(n50039), .Z(n49862) );
  AND U49881 ( .A(n1838), .B(n50040), .Z(n50039) );
  XOR U49882 ( .A(n50041), .B(n50038), .Z(n50040) );
  XOR U49883 ( .A(n49863), .B(n50034), .Z(n50036) );
  XOR U49884 ( .A(n50042), .B(n50043), .Z(n49863) );
  AND U49885 ( .A(n1846), .B(n50002), .Z(n50043) );
  XOR U49886 ( .A(n50042), .B(n50000), .Z(n50002) );
  XOR U49887 ( .A(n50044), .B(n50045), .Z(n50034) );
  AND U49888 ( .A(n50046), .B(n50047), .Z(n50045) );
  XNOR U49889 ( .A(n50044), .B(n49887), .Z(n50047) );
  IV U49890 ( .A(n49890), .Z(n49887) );
  XOR U49891 ( .A(n50048), .B(n50049), .Z(n49890) );
  AND U49892 ( .A(n1838), .B(n50050), .Z(n50049) );
  XNOR U49893 ( .A(n50051), .B(n50048), .Z(n50050) );
  XOR U49894 ( .A(n49891), .B(n50044), .Z(n50046) );
  XOR U49895 ( .A(n50052), .B(n50053), .Z(n49891) );
  AND U49896 ( .A(n1846), .B(n50011), .Z(n50053) );
  XOR U49897 ( .A(n50052), .B(n50009), .Z(n50011) );
  XOR U49898 ( .A(n49968), .B(n50054), .Z(n50044) );
  AND U49899 ( .A(n49970), .B(n50055), .Z(n50054) );
  XNOR U49900 ( .A(n49968), .B(n49938), .Z(n50055) );
  IV U49901 ( .A(n49941), .Z(n49938) );
  XOR U49902 ( .A(n50056), .B(n50057), .Z(n49941) );
  AND U49903 ( .A(n1838), .B(n50058), .Z(n50057) );
  XOR U49904 ( .A(n50059), .B(n50056), .Z(n50058) );
  XOR U49905 ( .A(n49942), .B(n49968), .Z(n49970) );
  XOR U49906 ( .A(n50060), .B(n50061), .Z(n49942) );
  AND U49907 ( .A(n1846), .B(n50021), .Z(n50061) );
  XOR U49908 ( .A(n50060), .B(n50019), .Z(n50021) );
  AND U49909 ( .A(n50022), .B(n49952), .Z(n49968) );
  XNOR U49910 ( .A(n50062), .B(n50063), .Z(n49952) );
  AND U49911 ( .A(n1838), .B(n50064), .Z(n50063) );
  XNOR U49912 ( .A(n50065), .B(n50062), .Z(n50064) );
  XNOR U49913 ( .A(n50066), .B(n50067), .Z(n1838) );
  AND U49914 ( .A(n50068), .B(n50069), .Z(n50067) );
  XOR U49915 ( .A(n50031), .B(n50066), .Z(n50069) );
  AND U49916 ( .A(n50070), .B(n50071), .Z(n50031) );
  XNOR U49917 ( .A(n50028), .B(n50066), .Z(n50068) );
  XNOR U49918 ( .A(n50072), .B(n50073), .Z(n50028) );
  AND U49919 ( .A(n1842), .B(n50074), .Z(n50073) );
  XNOR U49920 ( .A(n50075), .B(n50076), .Z(n50074) );
  XOR U49921 ( .A(n50077), .B(n50078), .Z(n50066) );
  AND U49922 ( .A(n50079), .B(n50080), .Z(n50078) );
  XNOR U49923 ( .A(n50077), .B(n50070), .Z(n50080) );
  IV U49924 ( .A(n50041), .Z(n50070) );
  XOR U49925 ( .A(n50081), .B(n50082), .Z(n50041) );
  XOR U49926 ( .A(n50083), .B(n50071), .Z(n50082) );
  AND U49927 ( .A(n50051), .B(n50084), .Z(n50071) );
  AND U49928 ( .A(n50085), .B(n50086), .Z(n50083) );
  XOR U49929 ( .A(n50087), .B(n50081), .Z(n50085) );
  XNOR U49930 ( .A(n50038), .B(n50077), .Z(n50079) );
  XNOR U49931 ( .A(n50088), .B(n50089), .Z(n50038) );
  AND U49932 ( .A(n1842), .B(n50090), .Z(n50089) );
  XNOR U49933 ( .A(n50091), .B(n50092), .Z(n50090) );
  XOR U49934 ( .A(n50093), .B(n50094), .Z(n50077) );
  AND U49935 ( .A(n50095), .B(n50096), .Z(n50094) );
  XNOR U49936 ( .A(n50093), .B(n50051), .Z(n50096) );
  XOR U49937 ( .A(n50097), .B(n50086), .Z(n50051) );
  XNOR U49938 ( .A(n50098), .B(n50081), .Z(n50086) );
  XOR U49939 ( .A(n50099), .B(n50100), .Z(n50081) );
  AND U49940 ( .A(n50101), .B(n50102), .Z(n50100) );
  XOR U49941 ( .A(n50103), .B(n50099), .Z(n50101) );
  XNOR U49942 ( .A(n50104), .B(n50105), .Z(n50098) );
  AND U49943 ( .A(n50106), .B(n50107), .Z(n50105) );
  XOR U49944 ( .A(n50104), .B(n50108), .Z(n50106) );
  XNOR U49945 ( .A(n50087), .B(n50084), .Z(n50097) );
  AND U49946 ( .A(n50109), .B(n50110), .Z(n50084) );
  XOR U49947 ( .A(n50111), .B(n50112), .Z(n50087) );
  AND U49948 ( .A(n50113), .B(n50114), .Z(n50112) );
  XOR U49949 ( .A(n50111), .B(n50115), .Z(n50113) );
  XNOR U49950 ( .A(n50048), .B(n50093), .Z(n50095) );
  XNOR U49951 ( .A(n50116), .B(n50117), .Z(n50048) );
  AND U49952 ( .A(n1842), .B(n50118), .Z(n50117) );
  XNOR U49953 ( .A(n50119), .B(n50120), .Z(n50118) );
  XOR U49954 ( .A(n50121), .B(n50122), .Z(n50093) );
  AND U49955 ( .A(n50123), .B(n50124), .Z(n50122) );
  XNOR U49956 ( .A(n50121), .B(n50109), .Z(n50124) );
  IV U49957 ( .A(n50059), .Z(n50109) );
  XNOR U49958 ( .A(n50125), .B(n50102), .Z(n50059) );
  XNOR U49959 ( .A(n50126), .B(n50108), .Z(n50102) );
  XNOR U49960 ( .A(n50127), .B(n50128), .Z(n50108) );
  NOR U49961 ( .A(n50129), .B(n50130), .Z(n50128) );
  XOR U49962 ( .A(n50127), .B(n50131), .Z(n50129) );
  XNOR U49963 ( .A(n50107), .B(n50099), .Z(n50126) );
  XOR U49964 ( .A(n50132), .B(n50133), .Z(n50099) );
  AND U49965 ( .A(n50134), .B(n50135), .Z(n50133) );
  XOR U49966 ( .A(n50132), .B(n50136), .Z(n50134) );
  XNOR U49967 ( .A(n50137), .B(n50104), .Z(n50107) );
  XOR U49968 ( .A(n50138), .B(n50139), .Z(n50104) );
  AND U49969 ( .A(n50140), .B(n50141), .Z(n50139) );
  XNOR U49970 ( .A(n50142), .B(n50143), .Z(n50140) );
  IV U49971 ( .A(n50138), .Z(n50142) );
  XNOR U49972 ( .A(n50144), .B(n50145), .Z(n50137) );
  NOR U49973 ( .A(n50146), .B(n50147), .Z(n50145) );
  XNOR U49974 ( .A(n50144), .B(n50148), .Z(n50146) );
  XNOR U49975 ( .A(n50103), .B(n50110), .Z(n50125) );
  NOR U49976 ( .A(n50065), .B(n50149), .Z(n50110) );
  XOR U49977 ( .A(n50115), .B(n50114), .Z(n50103) );
  XNOR U49978 ( .A(n50150), .B(n50111), .Z(n50114) );
  XOR U49979 ( .A(n50151), .B(n50152), .Z(n50111) );
  AND U49980 ( .A(n50153), .B(n50154), .Z(n50152) );
  XNOR U49981 ( .A(n50155), .B(n50156), .Z(n50153) );
  IV U49982 ( .A(n50151), .Z(n50155) );
  XNOR U49983 ( .A(n50157), .B(n50158), .Z(n50150) );
  NOR U49984 ( .A(n50159), .B(n50160), .Z(n50158) );
  XNOR U49985 ( .A(n50157), .B(n50161), .Z(n50159) );
  XOR U49986 ( .A(n50162), .B(n50163), .Z(n50115) );
  NOR U49987 ( .A(n50164), .B(n50165), .Z(n50163) );
  XNOR U49988 ( .A(n50162), .B(n50166), .Z(n50164) );
  XNOR U49989 ( .A(n50056), .B(n50121), .Z(n50123) );
  XNOR U49990 ( .A(n50167), .B(n50168), .Z(n50056) );
  AND U49991 ( .A(n1842), .B(n50169), .Z(n50168) );
  XNOR U49992 ( .A(n50170), .B(n50171), .Z(n50169) );
  AND U49993 ( .A(n50062), .B(n50065), .Z(n50121) );
  XOR U49994 ( .A(n50172), .B(n50149), .Z(n50065) );
  XNOR U49995 ( .A(p_input[1488]), .B(p_input[2048]), .Z(n50149) );
  XNOR U49996 ( .A(n50136), .B(n50135), .Z(n50172) );
  XNOR U49997 ( .A(n50173), .B(n50143), .Z(n50135) );
  XNOR U49998 ( .A(n50131), .B(n50130), .Z(n50143) );
  XNOR U49999 ( .A(n50174), .B(n50127), .Z(n50130) );
  XNOR U50000 ( .A(p_input[1498]), .B(p_input[2058]), .Z(n50127) );
  XOR U50001 ( .A(p_input[1499]), .B(n29030), .Z(n50174) );
  XOR U50002 ( .A(p_input[1500]), .B(p_input[2060]), .Z(n50131) );
  XOR U50003 ( .A(n50141), .B(n50175), .Z(n50173) );
  IV U50004 ( .A(n50132), .Z(n50175) );
  XOR U50005 ( .A(p_input[1489]), .B(p_input[2049]), .Z(n50132) );
  XNOR U50006 ( .A(n50176), .B(n50148), .Z(n50141) );
  XNOR U50007 ( .A(p_input[1503]), .B(n29033), .Z(n50148) );
  XOR U50008 ( .A(n50138), .B(n50147), .Z(n50176) );
  XOR U50009 ( .A(n50177), .B(n50144), .Z(n50147) );
  XOR U50010 ( .A(p_input[1501]), .B(p_input[2061]), .Z(n50144) );
  XOR U50011 ( .A(p_input[1502]), .B(n29035), .Z(n50177) );
  XOR U50012 ( .A(p_input[1497]), .B(p_input[2057]), .Z(n50138) );
  XOR U50013 ( .A(n50156), .B(n50154), .Z(n50136) );
  XNOR U50014 ( .A(n50178), .B(n50161), .Z(n50154) );
  XOR U50015 ( .A(p_input[1496]), .B(p_input[2056]), .Z(n50161) );
  XOR U50016 ( .A(n50151), .B(n50160), .Z(n50178) );
  XOR U50017 ( .A(n50179), .B(n50157), .Z(n50160) );
  XOR U50018 ( .A(p_input[1494]), .B(p_input[2054]), .Z(n50157) );
  XOR U50019 ( .A(p_input[1495]), .B(n30404), .Z(n50179) );
  XOR U50020 ( .A(p_input[1490]), .B(p_input[2050]), .Z(n50151) );
  XNOR U50021 ( .A(n50166), .B(n50165), .Z(n50156) );
  XOR U50022 ( .A(n50180), .B(n50162), .Z(n50165) );
  XOR U50023 ( .A(p_input[1491]), .B(p_input[2051]), .Z(n50162) );
  XOR U50024 ( .A(p_input[1492]), .B(n30406), .Z(n50180) );
  XOR U50025 ( .A(p_input[1493]), .B(p_input[2053]), .Z(n50166) );
  XNOR U50026 ( .A(n50181), .B(n50182), .Z(n50062) );
  AND U50027 ( .A(n1842), .B(n50183), .Z(n50182) );
  XNOR U50028 ( .A(n50184), .B(n50185), .Z(n1842) );
  AND U50029 ( .A(n50186), .B(n50187), .Z(n50185) );
  XOR U50030 ( .A(n50076), .B(n50184), .Z(n50187) );
  XNOR U50031 ( .A(n50188), .B(n50184), .Z(n50186) );
  XOR U50032 ( .A(n50189), .B(n50190), .Z(n50184) );
  AND U50033 ( .A(n50191), .B(n50192), .Z(n50190) );
  XOR U50034 ( .A(n50091), .B(n50189), .Z(n50192) );
  XOR U50035 ( .A(n50189), .B(n50092), .Z(n50191) );
  XOR U50036 ( .A(n50193), .B(n50194), .Z(n50189) );
  AND U50037 ( .A(n50195), .B(n50196), .Z(n50194) );
  XOR U50038 ( .A(n50119), .B(n50193), .Z(n50196) );
  XOR U50039 ( .A(n50193), .B(n50120), .Z(n50195) );
  XOR U50040 ( .A(n50197), .B(n50198), .Z(n50193) );
  AND U50041 ( .A(n50199), .B(n50200), .Z(n50198) );
  XOR U50042 ( .A(n50197), .B(n50170), .Z(n50200) );
  XNOR U50043 ( .A(n50201), .B(n50202), .Z(n50022) );
  AND U50044 ( .A(n1846), .B(n50203), .Z(n50202) );
  XNOR U50045 ( .A(n50204), .B(n50205), .Z(n1846) );
  AND U50046 ( .A(n50206), .B(n50207), .Z(n50205) );
  XOR U50047 ( .A(n50204), .B(n50032), .Z(n50207) );
  XNOR U50048 ( .A(n50204), .B(n49992), .Z(n50206) );
  XOR U50049 ( .A(n50208), .B(n50209), .Z(n50204) );
  AND U50050 ( .A(n50210), .B(n50211), .Z(n50209) );
  XOR U50051 ( .A(n50208), .B(n50000), .Z(n50210) );
  XOR U50052 ( .A(n50212), .B(n50213), .Z(n49983) );
  AND U50053 ( .A(n1850), .B(n50203), .Z(n50213) );
  XNOR U50054 ( .A(n50201), .B(n50212), .Z(n50203) );
  XNOR U50055 ( .A(n50214), .B(n50215), .Z(n1850) );
  AND U50056 ( .A(n50216), .B(n50217), .Z(n50215) );
  XNOR U50057 ( .A(n50218), .B(n50214), .Z(n50217) );
  IV U50058 ( .A(n50032), .Z(n50218) );
  XOR U50059 ( .A(n50188), .B(n50219), .Z(n50032) );
  AND U50060 ( .A(n1853), .B(n50220), .Z(n50219) );
  XOR U50061 ( .A(n50075), .B(n50072), .Z(n50220) );
  IV U50062 ( .A(n50188), .Z(n50075) );
  XNOR U50063 ( .A(n49992), .B(n50214), .Z(n50216) );
  XOR U50064 ( .A(n50221), .B(n50222), .Z(n49992) );
  AND U50065 ( .A(n1869), .B(n50223), .Z(n50222) );
  XOR U50066 ( .A(n50208), .B(n50224), .Z(n50214) );
  AND U50067 ( .A(n50225), .B(n50211), .Z(n50224) );
  XNOR U50068 ( .A(n50042), .B(n50208), .Z(n50211) );
  XOR U50069 ( .A(n50092), .B(n50226), .Z(n50042) );
  AND U50070 ( .A(n1853), .B(n50227), .Z(n50226) );
  XOR U50071 ( .A(n50088), .B(n50092), .Z(n50227) );
  XNOR U50072 ( .A(n50228), .B(n50208), .Z(n50225) );
  IV U50073 ( .A(n50000), .Z(n50228) );
  XOR U50074 ( .A(n50229), .B(n50230), .Z(n50000) );
  AND U50075 ( .A(n1869), .B(n50231), .Z(n50230) );
  XOR U50076 ( .A(n50232), .B(n50233), .Z(n50208) );
  AND U50077 ( .A(n50234), .B(n50235), .Z(n50233) );
  XNOR U50078 ( .A(n50052), .B(n50232), .Z(n50235) );
  XOR U50079 ( .A(n50120), .B(n50236), .Z(n50052) );
  AND U50080 ( .A(n1853), .B(n50237), .Z(n50236) );
  XOR U50081 ( .A(n50116), .B(n50120), .Z(n50237) );
  XOR U50082 ( .A(n50232), .B(n50009), .Z(n50234) );
  XOR U50083 ( .A(n50238), .B(n50239), .Z(n50009) );
  AND U50084 ( .A(n1869), .B(n50240), .Z(n50239) );
  XOR U50085 ( .A(n50241), .B(n50242), .Z(n50232) );
  AND U50086 ( .A(n50243), .B(n50244), .Z(n50242) );
  XNOR U50087 ( .A(n50241), .B(n50060), .Z(n50244) );
  XOR U50088 ( .A(n50171), .B(n50245), .Z(n50060) );
  AND U50089 ( .A(n1853), .B(n50246), .Z(n50245) );
  XOR U50090 ( .A(n50167), .B(n50171), .Z(n50246) );
  XNOR U50091 ( .A(n50247), .B(n50241), .Z(n50243) );
  IV U50092 ( .A(n50019), .Z(n50247) );
  XOR U50093 ( .A(n50248), .B(n50249), .Z(n50019) );
  AND U50094 ( .A(n1869), .B(n50250), .Z(n50249) );
  AND U50095 ( .A(n50212), .B(n50201), .Z(n50241) );
  XNOR U50096 ( .A(n50251), .B(n50252), .Z(n50201) );
  AND U50097 ( .A(n1853), .B(n50183), .Z(n50252) );
  XNOR U50098 ( .A(n50181), .B(n50251), .Z(n50183) );
  XNOR U50099 ( .A(n50253), .B(n50254), .Z(n1853) );
  AND U50100 ( .A(n50255), .B(n50256), .Z(n50254) );
  XNOR U50101 ( .A(n50253), .B(n50072), .Z(n50256) );
  IV U50102 ( .A(n50076), .Z(n50072) );
  XOR U50103 ( .A(n50257), .B(n50258), .Z(n50076) );
  AND U50104 ( .A(n1857), .B(n50259), .Z(n50258) );
  XOR U50105 ( .A(n50260), .B(n50257), .Z(n50259) );
  XNOR U50106 ( .A(n50253), .B(n50188), .Z(n50255) );
  XOR U50107 ( .A(n50261), .B(n50262), .Z(n50188) );
  AND U50108 ( .A(n1865), .B(n50223), .Z(n50262) );
  XOR U50109 ( .A(n50221), .B(n50261), .Z(n50223) );
  XOR U50110 ( .A(n50263), .B(n50264), .Z(n50253) );
  AND U50111 ( .A(n50265), .B(n50266), .Z(n50264) );
  XNOR U50112 ( .A(n50263), .B(n50088), .Z(n50266) );
  IV U50113 ( .A(n50091), .Z(n50088) );
  XOR U50114 ( .A(n50267), .B(n50268), .Z(n50091) );
  AND U50115 ( .A(n1857), .B(n50269), .Z(n50268) );
  XOR U50116 ( .A(n50270), .B(n50267), .Z(n50269) );
  XOR U50117 ( .A(n50092), .B(n50263), .Z(n50265) );
  XOR U50118 ( .A(n50271), .B(n50272), .Z(n50092) );
  AND U50119 ( .A(n1865), .B(n50231), .Z(n50272) );
  XOR U50120 ( .A(n50271), .B(n50229), .Z(n50231) );
  XOR U50121 ( .A(n50273), .B(n50274), .Z(n50263) );
  AND U50122 ( .A(n50275), .B(n50276), .Z(n50274) );
  XNOR U50123 ( .A(n50273), .B(n50116), .Z(n50276) );
  IV U50124 ( .A(n50119), .Z(n50116) );
  XOR U50125 ( .A(n50277), .B(n50278), .Z(n50119) );
  AND U50126 ( .A(n1857), .B(n50279), .Z(n50278) );
  XNOR U50127 ( .A(n50280), .B(n50277), .Z(n50279) );
  XOR U50128 ( .A(n50120), .B(n50273), .Z(n50275) );
  XOR U50129 ( .A(n50281), .B(n50282), .Z(n50120) );
  AND U50130 ( .A(n1865), .B(n50240), .Z(n50282) );
  XOR U50131 ( .A(n50281), .B(n50238), .Z(n50240) );
  XOR U50132 ( .A(n50197), .B(n50283), .Z(n50273) );
  AND U50133 ( .A(n50199), .B(n50284), .Z(n50283) );
  XNOR U50134 ( .A(n50197), .B(n50167), .Z(n50284) );
  IV U50135 ( .A(n50170), .Z(n50167) );
  XOR U50136 ( .A(n50285), .B(n50286), .Z(n50170) );
  AND U50137 ( .A(n1857), .B(n50287), .Z(n50286) );
  XOR U50138 ( .A(n50288), .B(n50285), .Z(n50287) );
  XOR U50139 ( .A(n50171), .B(n50197), .Z(n50199) );
  XOR U50140 ( .A(n50289), .B(n50290), .Z(n50171) );
  AND U50141 ( .A(n1865), .B(n50250), .Z(n50290) );
  XOR U50142 ( .A(n50289), .B(n50248), .Z(n50250) );
  AND U50143 ( .A(n50251), .B(n50181), .Z(n50197) );
  XNOR U50144 ( .A(n50291), .B(n50292), .Z(n50181) );
  AND U50145 ( .A(n1857), .B(n50293), .Z(n50292) );
  XNOR U50146 ( .A(n50294), .B(n50291), .Z(n50293) );
  XNOR U50147 ( .A(n50295), .B(n50296), .Z(n1857) );
  AND U50148 ( .A(n50297), .B(n50298), .Z(n50296) );
  XOR U50149 ( .A(n50260), .B(n50295), .Z(n50298) );
  AND U50150 ( .A(n50299), .B(n50300), .Z(n50260) );
  XNOR U50151 ( .A(n50257), .B(n50295), .Z(n50297) );
  XNOR U50152 ( .A(n50301), .B(n50302), .Z(n50257) );
  AND U50153 ( .A(n1861), .B(n50303), .Z(n50302) );
  XNOR U50154 ( .A(n50304), .B(n50305), .Z(n50303) );
  XOR U50155 ( .A(n50306), .B(n50307), .Z(n50295) );
  AND U50156 ( .A(n50308), .B(n50309), .Z(n50307) );
  XNOR U50157 ( .A(n50306), .B(n50299), .Z(n50309) );
  IV U50158 ( .A(n50270), .Z(n50299) );
  XOR U50159 ( .A(n50310), .B(n50311), .Z(n50270) );
  XOR U50160 ( .A(n50312), .B(n50300), .Z(n50311) );
  AND U50161 ( .A(n50280), .B(n50313), .Z(n50300) );
  AND U50162 ( .A(n50314), .B(n50315), .Z(n50312) );
  XOR U50163 ( .A(n50316), .B(n50310), .Z(n50314) );
  XNOR U50164 ( .A(n50267), .B(n50306), .Z(n50308) );
  XNOR U50165 ( .A(n50317), .B(n50318), .Z(n50267) );
  AND U50166 ( .A(n1861), .B(n50319), .Z(n50318) );
  XNOR U50167 ( .A(n50320), .B(n50321), .Z(n50319) );
  XOR U50168 ( .A(n50322), .B(n50323), .Z(n50306) );
  AND U50169 ( .A(n50324), .B(n50325), .Z(n50323) );
  XNOR U50170 ( .A(n50322), .B(n50280), .Z(n50325) );
  XOR U50171 ( .A(n50326), .B(n50315), .Z(n50280) );
  XNOR U50172 ( .A(n50327), .B(n50310), .Z(n50315) );
  XOR U50173 ( .A(n50328), .B(n50329), .Z(n50310) );
  AND U50174 ( .A(n50330), .B(n50331), .Z(n50329) );
  XOR U50175 ( .A(n50332), .B(n50328), .Z(n50330) );
  XNOR U50176 ( .A(n50333), .B(n50334), .Z(n50327) );
  AND U50177 ( .A(n50335), .B(n50336), .Z(n50334) );
  XOR U50178 ( .A(n50333), .B(n50337), .Z(n50335) );
  XNOR U50179 ( .A(n50316), .B(n50313), .Z(n50326) );
  AND U50180 ( .A(n50338), .B(n50339), .Z(n50313) );
  XOR U50181 ( .A(n50340), .B(n50341), .Z(n50316) );
  AND U50182 ( .A(n50342), .B(n50343), .Z(n50341) );
  XOR U50183 ( .A(n50340), .B(n50344), .Z(n50342) );
  XNOR U50184 ( .A(n50277), .B(n50322), .Z(n50324) );
  XNOR U50185 ( .A(n50345), .B(n50346), .Z(n50277) );
  AND U50186 ( .A(n1861), .B(n50347), .Z(n50346) );
  XNOR U50187 ( .A(n50348), .B(n50349), .Z(n50347) );
  XOR U50188 ( .A(n50350), .B(n50351), .Z(n50322) );
  AND U50189 ( .A(n50352), .B(n50353), .Z(n50351) );
  XNOR U50190 ( .A(n50350), .B(n50338), .Z(n50353) );
  IV U50191 ( .A(n50288), .Z(n50338) );
  XNOR U50192 ( .A(n50354), .B(n50331), .Z(n50288) );
  XNOR U50193 ( .A(n50355), .B(n50337), .Z(n50331) );
  XNOR U50194 ( .A(n50356), .B(n50357), .Z(n50337) );
  NOR U50195 ( .A(n50358), .B(n50359), .Z(n50357) );
  XOR U50196 ( .A(n50356), .B(n50360), .Z(n50358) );
  XNOR U50197 ( .A(n50336), .B(n50328), .Z(n50355) );
  XOR U50198 ( .A(n50361), .B(n50362), .Z(n50328) );
  AND U50199 ( .A(n50363), .B(n50364), .Z(n50362) );
  XOR U50200 ( .A(n50361), .B(n50365), .Z(n50363) );
  XNOR U50201 ( .A(n50366), .B(n50333), .Z(n50336) );
  XOR U50202 ( .A(n50367), .B(n50368), .Z(n50333) );
  AND U50203 ( .A(n50369), .B(n50370), .Z(n50368) );
  XNOR U50204 ( .A(n50371), .B(n50372), .Z(n50369) );
  IV U50205 ( .A(n50367), .Z(n50371) );
  XNOR U50206 ( .A(n50373), .B(n50374), .Z(n50366) );
  NOR U50207 ( .A(n50375), .B(n50376), .Z(n50374) );
  XNOR U50208 ( .A(n50373), .B(n50377), .Z(n50375) );
  XNOR U50209 ( .A(n50332), .B(n50339), .Z(n50354) );
  NOR U50210 ( .A(n50294), .B(n50378), .Z(n50339) );
  XOR U50211 ( .A(n50344), .B(n50343), .Z(n50332) );
  XNOR U50212 ( .A(n50379), .B(n50340), .Z(n50343) );
  XOR U50213 ( .A(n50380), .B(n50381), .Z(n50340) );
  AND U50214 ( .A(n50382), .B(n50383), .Z(n50381) );
  XNOR U50215 ( .A(n50384), .B(n50385), .Z(n50382) );
  IV U50216 ( .A(n50380), .Z(n50384) );
  XNOR U50217 ( .A(n50386), .B(n50387), .Z(n50379) );
  NOR U50218 ( .A(n50388), .B(n50389), .Z(n50387) );
  XNOR U50219 ( .A(n50386), .B(n50390), .Z(n50388) );
  XOR U50220 ( .A(n50391), .B(n50392), .Z(n50344) );
  NOR U50221 ( .A(n50393), .B(n50394), .Z(n50392) );
  XNOR U50222 ( .A(n50391), .B(n50395), .Z(n50393) );
  XNOR U50223 ( .A(n50285), .B(n50350), .Z(n50352) );
  XNOR U50224 ( .A(n50396), .B(n50397), .Z(n50285) );
  AND U50225 ( .A(n1861), .B(n50398), .Z(n50397) );
  XNOR U50226 ( .A(n50399), .B(n50400), .Z(n50398) );
  AND U50227 ( .A(n50291), .B(n50294), .Z(n50350) );
  XOR U50228 ( .A(n50401), .B(n50378), .Z(n50294) );
  XNOR U50229 ( .A(p_input[1504]), .B(p_input[2048]), .Z(n50378) );
  XNOR U50230 ( .A(n50365), .B(n50364), .Z(n50401) );
  XNOR U50231 ( .A(n50402), .B(n50372), .Z(n50364) );
  XNOR U50232 ( .A(n50360), .B(n50359), .Z(n50372) );
  XNOR U50233 ( .A(n50403), .B(n50356), .Z(n50359) );
  XNOR U50234 ( .A(p_input[1514]), .B(p_input[2058]), .Z(n50356) );
  XOR U50235 ( .A(p_input[1515]), .B(n29030), .Z(n50403) );
  XOR U50236 ( .A(p_input[1516]), .B(p_input[2060]), .Z(n50360) );
  XOR U50237 ( .A(n50370), .B(n50404), .Z(n50402) );
  IV U50238 ( .A(n50361), .Z(n50404) );
  XOR U50239 ( .A(p_input[1505]), .B(p_input[2049]), .Z(n50361) );
  XNOR U50240 ( .A(n50405), .B(n50377), .Z(n50370) );
  XNOR U50241 ( .A(p_input[1519]), .B(n29033), .Z(n50377) );
  XOR U50242 ( .A(n50367), .B(n50376), .Z(n50405) );
  XOR U50243 ( .A(n50406), .B(n50373), .Z(n50376) );
  XOR U50244 ( .A(p_input[1517]), .B(p_input[2061]), .Z(n50373) );
  XOR U50245 ( .A(p_input[1518]), .B(n29035), .Z(n50406) );
  XOR U50246 ( .A(p_input[1513]), .B(p_input[2057]), .Z(n50367) );
  XOR U50247 ( .A(n50385), .B(n50383), .Z(n50365) );
  XNOR U50248 ( .A(n50407), .B(n50390), .Z(n50383) );
  XOR U50249 ( .A(p_input[1512]), .B(p_input[2056]), .Z(n50390) );
  XOR U50250 ( .A(n50380), .B(n50389), .Z(n50407) );
  XOR U50251 ( .A(n50408), .B(n50386), .Z(n50389) );
  XOR U50252 ( .A(p_input[1510]), .B(p_input[2054]), .Z(n50386) );
  XOR U50253 ( .A(p_input[1511]), .B(n30404), .Z(n50408) );
  XOR U50254 ( .A(p_input[1506]), .B(p_input[2050]), .Z(n50380) );
  XNOR U50255 ( .A(n50395), .B(n50394), .Z(n50385) );
  XOR U50256 ( .A(n50409), .B(n50391), .Z(n50394) );
  XOR U50257 ( .A(p_input[1507]), .B(p_input[2051]), .Z(n50391) );
  XOR U50258 ( .A(p_input[1508]), .B(n30406), .Z(n50409) );
  XOR U50259 ( .A(p_input[1509]), .B(p_input[2053]), .Z(n50395) );
  XNOR U50260 ( .A(n50410), .B(n50411), .Z(n50291) );
  AND U50261 ( .A(n1861), .B(n50412), .Z(n50411) );
  XNOR U50262 ( .A(n50413), .B(n50414), .Z(n1861) );
  AND U50263 ( .A(n50415), .B(n50416), .Z(n50414) );
  XOR U50264 ( .A(n50305), .B(n50413), .Z(n50416) );
  XNOR U50265 ( .A(n50417), .B(n50413), .Z(n50415) );
  XOR U50266 ( .A(n50418), .B(n50419), .Z(n50413) );
  AND U50267 ( .A(n50420), .B(n50421), .Z(n50419) );
  XOR U50268 ( .A(n50320), .B(n50418), .Z(n50421) );
  XOR U50269 ( .A(n50418), .B(n50321), .Z(n50420) );
  XOR U50270 ( .A(n50422), .B(n50423), .Z(n50418) );
  AND U50271 ( .A(n50424), .B(n50425), .Z(n50423) );
  XOR U50272 ( .A(n50348), .B(n50422), .Z(n50425) );
  XOR U50273 ( .A(n50422), .B(n50349), .Z(n50424) );
  XOR U50274 ( .A(n50426), .B(n50427), .Z(n50422) );
  AND U50275 ( .A(n50428), .B(n50429), .Z(n50427) );
  XOR U50276 ( .A(n50426), .B(n50399), .Z(n50429) );
  XNOR U50277 ( .A(n50430), .B(n50431), .Z(n50251) );
  AND U50278 ( .A(n1865), .B(n50432), .Z(n50431) );
  XNOR U50279 ( .A(n50433), .B(n50434), .Z(n1865) );
  AND U50280 ( .A(n50435), .B(n50436), .Z(n50434) );
  XOR U50281 ( .A(n50433), .B(n50261), .Z(n50436) );
  XNOR U50282 ( .A(n50433), .B(n50221), .Z(n50435) );
  XOR U50283 ( .A(n50437), .B(n50438), .Z(n50433) );
  AND U50284 ( .A(n50439), .B(n50440), .Z(n50438) );
  XOR U50285 ( .A(n50437), .B(n50229), .Z(n50439) );
  XOR U50286 ( .A(n50441), .B(n50442), .Z(n50212) );
  AND U50287 ( .A(n1869), .B(n50432), .Z(n50442) );
  XNOR U50288 ( .A(n50430), .B(n50441), .Z(n50432) );
  XNOR U50289 ( .A(n50443), .B(n50444), .Z(n1869) );
  AND U50290 ( .A(n50445), .B(n50446), .Z(n50444) );
  XNOR U50291 ( .A(n50447), .B(n50443), .Z(n50446) );
  IV U50292 ( .A(n50261), .Z(n50447) );
  XOR U50293 ( .A(n50417), .B(n50448), .Z(n50261) );
  AND U50294 ( .A(n1872), .B(n50449), .Z(n50448) );
  XOR U50295 ( .A(n50304), .B(n50301), .Z(n50449) );
  IV U50296 ( .A(n50417), .Z(n50304) );
  XNOR U50297 ( .A(n50221), .B(n50443), .Z(n50445) );
  XOR U50298 ( .A(n50450), .B(n50451), .Z(n50221) );
  AND U50299 ( .A(n1888), .B(n50452), .Z(n50451) );
  XOR U50300 ( .A(n50437), .B(n50453), .Z(n50443) );
  AND U50301 ( .A(n50454), .B(n50440), .Z(n50453) );
  XNOR U50302 ( .A(n50271), .B(n50437), .Z(n50440) );
  XOR U50303 ( .A(n50321), .B(n50455), .Z(n50271) );
  AND U50304 ( .A(n1872), .B(n50456), .Z(n50455) );
  XOR U50305 ( .A(n50317), .B(n50321), .Z(n50456) );
  XNOR U50306 ( .A(n50457), .B(n50437), .Z(n50454) );
  IV U50307 ( .A(n50229), .Z(n50457) );
  XOR U50308 ( .A(n50458), .B(n50459), .Z(n50229) );
  AND U50309 ( .A(n1888), .B(n50460), .Z(n50459) );
  XOR U50310 ( .A(n50461), .B(n50462), .Z(n50437) );
  AND U50311 ( .A(n50463), .B(n50464), .Z(n50462) );
  XNOR U50312 ( .A(n50281), .B(n50461), .Z(n50464) );
  XOR U50313 ( .A(n50349), .B(n50465), .Z(n50281) );
  AND U50314 ( .A(n1872), .B(n50466), .Z(n50465) );
  XOR U50315 ( .A(n50345), .B(n50349), .Z(n50466) );
  XOR U50316 ( .A(n50461), .B(n50238), .Z(n50463) );
  XOR U50317 ( .A(n50467), .B(n50468), .Z(n50238) );
  AND U50318 ( .A(n1888), .B(n50469), .Z(n50468) );
  XOR U50319 ( .A(n50470), .B(n50471), .Z(n50461) );
  AND U50320 ( .A(n50472), .B(n50473), .Z(n50471) );
  XNOR U50321 ( .A(n50470), .B(n50289), .Z(n50473) );
  XOR U50322 ( .A(n50400), .B(n50474), .Z(n50289) );
  AND U50323 ( .A(n1872), .B(n50475), .Z(n50474) );
  XOR U50324 ( .A(n50396), .B(n50400), .Z(n50475) );
  XNOR U50325 ( .A(n50476), .B(n50470), .Z(n50472) );
  IV U50326 ( .A(n50248), .Z(n50476) );
  XOR U50327 ( .A(n50477), .B(n50478), .Z(n50248) );
  AND U50328 ( .A(n1888), .B(n50479), .Z(n50478) );
  AND U50329 ( .A(n50441), .B(n50430), .Z(n50470) );
  XNOR U50330 ( .A(n50480), .B(n50481), .Z(n50430) );
  AND U50331 ( .A(n1872), .B(n50412), .Z(n50481) );
  XNOR U50332 ( .A(n50410), .B(n50480), .Z(n50412) );
  XNOR U50333 ( .A(n50482), .B(n50483), .Z(n1872) );
  AND U50334 ( .A(n50484), .B(n50485), .Z(n50483) );
  XNOR U50335 ( .A(n50482), .B(n50301), .Z(n50485) );
  IV U50336 ( .A(n50305), .Z(n50301) );
  XOR U50337 ( .A(n50486), .B(n50487), .Z(n50305) );
  AND U50338 ( .A(n1876), .B(n50488), .Z(n50487) );
  XOR U50339 ( .A(n50489), .B(n50486), .Z(n50488) );
  XNOR U50340 ( .A(n50482), .B(n50417), .Z(n50484) );
  XOR U50341 ( .A(n50490), .B(n50491), .Z(n50417) );
  AND U50342 ( .A(n1884), .B(n50452), .Z(n50491) );
  XOR U50343 ( .A(n50450), .B(n50490), .Z(n50452) );
  XOR U50344 ( .A(n50492), .B(n50493), .Z(n50482) );
  AND U50345 ( .A(n50494), .B(n50495), .Z(n50493) );
  XNOR U50346 ( .A(n50492), .B(n50317), .Z(n50495) );
  IV U50347 ( .A(n50320), .Z(n50317) );
  XOR U50348 ( .A(n50496), .B(n50497), .Z(n50320) );
  AND U50349 ( .A(n1876), .B(n50498), .Z(n50497) );
  XOR U50350 ( .A(n50499), .B(n50496), .Z(n50498) );
  XOR U50351 ( .A(n50321), .B(n50492), .Z(n50494) );
  XOR U50352 ( .A(n50500), .B(n50501), .Z(n50321) );
  AND U50353 ( .A(n1884), .B(n50460), .Z(n50501) );
  XOR U50354 ( .A(n50500), .B(n50458), .Z(n50460) );
  XOR U50355 ( .A(n50502), .B(n50503), .Z(n50492) );
  AND U50356 ( .A(n50504), .B(n50505), .Z(n50503) );
  XNOR U50357 ( .A(n50502), .B(n50345), .Z(n50505) );
  IV U50358 ( .A(n50348), .Z(n50345) );
  XOR U50359 ( .A(n50506), .B(n50507), .Z(n50348) );
  AND U50360 ( .A(n1876), .B(n50508), .Z(n50507) );
  XNOR U50361 ( .A(n50509), .B(n50506), .Z(n50508) );
  XOR U50362 ( .A(n50349), .B(n50502), .Z(n50504) );
  XOR U50363 ( .A(n50510), .B(n50511), .Z(n50349) );
  AND U50364 ( .A(n1884), .B(n50469), .Z(n50511) );
  XOR U50365 ( .A(n50510), .B(n50467), .Z(n50469) );
  XOR U50366 ( .A(n50426), .B(n50512), .Z(n50502) );
  AND U50367 ( .A(n50428), .B(n50513), .Z(n50512) );
  XNOR U50368 ( .A(n50426), .B(n50396), .Z(n50513) );
  IV U50369 ( .A(n50399), .Z(n50396) );
  XOR U50370 ( .A(n50514), .B(n50515), .Z(n50399) );
  AND U50371 ( .A(n1876), .B(n50516), .Z(n50515) );
  XOR U50372 ( .A(n50517), .B(n50514), .Z(n50516) );
  XOR U50373 ( .A(n50400), .B(n50426), .Z(n50428) );
  XOR U50374 ( .A(n50518), .B(n50519), .Z(n50400) );
  AND U50375 ( .A(n1884), .B(n50479), .Z(n50519) );
  XOR U50376 ( .A(n50518), .B(n50477), .Z(n50479) );
  AND U50377 ( .A(n50480), .B(n50410), .Z(n50426) );
  XNOR U50378 ( .A(n50520), .B(n50521), .Z(n50410) );
  AND U50379 ( .A(n1876), .B(n50522), .Z(n50521) );
  XNOR U50380 ( .A(n50523), .B(n50520), .Z(n50522) );
  XNOR U50381 ( .A(n50524), .B(n50525), .Z(n1876) );
  AND U50382 ( .A(n50526), .B(n50527), .Z(n50525) );
  XOR U50383 ( .A(n50489), .B(n50524), .Z(n50527) );
  AND U50384 ( .A(n50528), .B(n50529), .Z(n50489) );
  XNOR U50385 ( .A(n50486), .B(n50524), .Z(n50526) );
  XNOR U50386 ( .A(n50530), .B(n50531), .Z(n50486) );
  AND U50387 ( .A(n1880), .B(n50532), .Z(n50531) );
  XNOR U50388 ( .A(n50533), .B(n50534), .Z(n50532) );
  XOR U50389 ( .A(n50535), .B(n50536), .Z(n50524) );
  AND U50390 ( .A(n50537), .B(n50538), .Z(n50536) );
  XNOR U50391 ( .A(n50535), .B(n50528), .Z(n50538) );
  IV U50392 ( .A(n50499), .Z(n50528) );
  XOR U50393 ( .A(n50539), .B(n50540), .Z(n50499) );
  XOR U50394 ( .A(n50541), .B(n50529), .Z(n50540) );
  AND U50395 ( .A(n50509), .B(n50542), .Z(n50529) );
  AND U50396 ( .A(n50543), .B(n50544), .Z(n50541) );
  XOR U50397 ( .A(n50545), .B(n50539), .Z(n50543) );
  XNOR U50398 ( .A(n50496), .B(n50535), .Z(n50537) );
  XNOR U50399 ( .A(n50546), .B(n50547), .Z(n50496) );
  AND U50400 ( .A(n1880), .B(n50548), .Z(n50547) );
  XNOR U50401 ( .A(n50549), .B(n50550), .Z(n50548) );
  XOR U50402 ( .A(n50551), .B(n50552), .Z(n50535) );
  AND U50403 ( .A(n50553), .B(n50554), .Z(n50552) );
  XNOR U50404 ( .A(n50551), .B(n50509), .Z(n50554) );
  XOR U50405 ( .A(n50555), .B(n50544), .Z(n50509) );
  XNOR U50406 ( .A(n50556), .B(n50539), .Z(n50544) );
  XOR U50407 ( .A(n50557), .B(n50558), .Z(n50539) );
  AND U50408 ( .A(n50559), .B(n50560), .Z(n50558) );
  XOR U50409 ( .A(n50561), .B(n50557), .Z(n50559) );
  XNOR U50410 ( .A(n50562), .B(n50563), .Z(n50556) );
  AND U50411 ( .A(n50564), .B(n50565), .Z(n50563) );
  XOR U50412 ( .A(n50562), .B(n50566), .Z(n50564) );
  XNOR U50413 ( .A(n50545), .B(n50542), .Z(n50555) );
  AND U50414 ( .A(n50567), .B(n50568), .Z(n50542) );
  XOR U50415 ( .A(n50569), .B(n50570), .Z(n50545) );
  AND U50416 ( .A(n50571), .B(n50572), .Z(n50570) );
  XOR U50417 ( .A(n50569), .B(n50573), .Z(n50571) );
  XNOR U50418 ( .A(n50506), .B(n50551), .Z(n50553) );
  XNOR U50419 ( .A(n50574), .B(n50575), .Z(n50506) );
  AND U50420 ( .A(n1880), .B(n50576), .Z(n50575) );
  XNOR U50421 ( .A(n50577), .B(n50578), .Z(n50576) );
  XOR U50422 ( .A(n50579), .B(n50580), .Z(n50551) );
  AND U50423 ( .A(n50581), .B(n50582), .Z(n50580) );
  XNOR U50424 ( .A(n50579), .B(n50567), .Z(n50582) );
  IV U50425 ( .A(n50517), .Z(n50567) );
  XNOR U50426 ( .A(n50583), .B(n50560), .Z(n50517) );
  XNOR U50427 ( .A(n50584), .B(n50566), .Z(n50560) );
  XNOR U50428 ( .A(n50585), .B(n50586), .Z(n50566) );
  NOR U50429 ( .A(n50587), .B(n50588), .Z(n50586) );
  XOR U50430 ( .A(n50585), .B(n50589), .Z(n50587) );
  XNOR U50431 ( .A(n50565), .B(n50557), .Z(n50584) );
  XOR U50432 ( .A(n50590), .B(n50591), .Z(n50557) );
  AND U50433 ( .A(n50592), .B(n50593), .Z(n50591) );
  XOR U50434 ( .A(n50590), .B(n50594), .Z(n50592) );
  XNOR U50435 ( .A(n50595), .B(n50562), .Z(n50565) );
  XOR U50436 ( .A(n50596), .B(n50597), .Z(n50562) );
  AND U50437 ( .A(n50598), .B(n50599), .Z(n50597) );
  XNOR U50438 ( .A(n50600), .B(n50601), .Z(n50598) );
  IV U50439 ( .A(n50596), .Z(n50600) );
  XNOR U50440 ( .A(n50602), .B(n50603), .Z(n50595) );
  NOR U50441 ( .A(n50604), .B(n50605), .Z(n50603) );
  XNOR U50442 ( .A(n50602), .B(n50606), .Z(n50604) );
  XNOR U50443 ( .A(n50561), .B(n50568), .Z(n50583) );
  NOR U50444 ( .A(n50523), .B(n50607), .Z(n50568) );
  XOR U50445 ( .A(n50573), .B(n50572), .Z(n50561) );
  XNOR U50446 ( .A(n50608), .B(n50569), .Z(n50572) );
  XOR U50447 ( .A(n50609), .B(n50610), .Z(n50569) );
  AND U50448 ( .A(n50611), .B(n50612), .Z(n50610) );
  XNOR U50449 ( .A(n50613), .B(n50614), .Z(n50611) );
  IV U50450 ( .A(n50609), .Z(n50613) );
  XNOR U50451 ( .A(n50615), .B(n50616), .Z(n50608) );
  NOR U50452 ( .A(n50617), .B(n50618), .Z(n50616) );
  XNOR U50453 ( .A(n50615), .B(n50619), .Z(n50617) );
  XOR U50454 ( .A(n50620), .B(n50621), .Z(n50573) );
  NOR U50455 ( .A(n50622), .B(n50623), .Z(n50621) );
  XNOR U50456 ( .A(n50620), .B(n50624), .Z(n50622) );
  XNOR U50457 ( .A(n50514), .B(n50579), .Z(n50581) );
  XNOR U50458 ( .A(n50625), .B(n50626), .Z(n50514) );
  AND U50459 ( .A(n1880), .B(n50627), .Z(n50626) );
  XNOR U50460 ( .A(n50628), .B(n50629), .Z(n50627) );
  AND U50461 ( .A(n50520), .B(n50523), .Z(n50579) );
  XOR U50462 ( .A(n50630), .B(n50607), .Z(n50523) );
  XNOR U50463 ( .A(p_input[1520]), .B(p_input[2048]), .Z(n50607) );
  XNOR U50464 ( .A(n50594), .B(n50593), .Z(n50630) );
  XNOR U50465 ( .A(n50631), .B(n50601), .Z(n50593) );
  XNOR U50466 ( .A(n50589), .B(n50588), .Z(n50601) );
  XNOR U50467 ( .A(n50632), .B(n50585), .Z(n50588) );
  XNOR U50468 ( .A(p_input[1530]), .B(p_input[2058]), .Z(n50585) );
  XOR U50469 ( .A(p_input[1531]), .B(n29030), .Z(n50632) );
  XOR U50470 ( .A(p_input[1532]), .B(p_input[2060]), .Z(n50589) );
  XOR U50471 ( .A(n50599), .B(n50633), .Z(n50631) );
  IV U50472 ( .A(n50590), .Z(n50633) );
  XOR U50473 ( .A(p_input[1521]), .B(p_input[2049]), .Z(n50590) );
  XNOR U50474 ( .A(n50634), .B(n50606), .Z(n50599) );
  XNOR U50475 ( .A(p_input[1535]), .B(n29033), .Z(n50606) );
  XOR U50476 ( .A(n50596), .B(n50605), .Z(n50634) );
  XOR U50477 ( .A(n50635), .B(n50602), .Z(n50605) );
  XOR U50478 ( .A(p_input[1533]), .B(p_input[2061]), .Z(n50602) );
  XOR U50479 ( .A(p_input[1534]), .B(n29035), .Z(n50635) );
  XOR U50480 ( .A(p_input[1529]), .B(p_input[2057]), .Z(n50596) );
  XOR U50481 ( .A(n50614), .B(n50612), .Z(n50594) );
  XNOR U50482 ( .A(n50636), .B(n50619), .Z(n50612) );
  XOR U50483 ( .A(p_input[1528]), .B(p_input[2056]), .Z(n50619) );
  XOR U50484 ( .A(n50609), .B(n50618), .Z(n50636) );
  XOR U50485 ( .A(n50637), .B(n50615), .Z(n50618) );
  XOR U50486 ( .A(p_input[1526]), .B(p_input[2054]), .Z(n50615) );
  XOR U50487 ( .A(p_input[1527]), .B(n30404), .Z(n50637) );
  XOR U50488 ( .A(p_input[1522]), .B(p_input[2050]), .Z(n50609) );
  XNOR U50489 ( .A(n50624), .B(n50623), .Z(n50614) );
  XOR U50490 ( .A(n50638), .B(n50620), .Z(n50623) );
  XOR U50491 ( .A(p_input[1523]), .B(p_input[2051]), .Z(n50620) );
  XOR U50492 ( .A(p_input[1524]), .B(n30406), .Z(n50638) );
  XOR U50493 ( .A(p_input[1525]), .B(p_input[2053]), .Z(n50624) );
  XNOR U50494 ( .A(n50639), .B(n50640), .Z(n50520) );
  AND U50495 ( .A(n1880), .B(n50641), .Z(n50640) );
  XNOR U50496 ( .A(n50642), .B(n50643), .Z(n1880) );
  AND U50497 ( .A(n50644), .B(n50645), .Z(n50643) );
  XOR U50498 ( .A(n50534), .B(n50642), .Z(n50645) );
  XNOR U50499 ( .A(n50646), .B(n50642), .Z(n50644) );
  XOR U50500 ( .A(n50647), .B(n50648), .Z(n50642) );
  AND U50501 ( .A(n50649), .B(n50650), .Z(n50648) );
  XOR U50502 ( .A(n50549), .B(n50647), .Z(n50650) );
  XOR U50503 ( .A(n50647), .B(n50550), .Z(n50649) );
  XOR U50504 ( .A(n50651), .B(n50652), .Z(n50647) );
  AND U50505 ( .A(n50653), .B(n50654), .Z(n50652) );
  XOR U50506 ( .A(n50577), .B(n50651), .Z(n50654) );
  XOR U50507 ( .A(n50651), .B(n50578), .Z(n50653) );
  XOR U50508 ( .A(n50655), .B(n50656), .Z(n50651) );
  AND U50509 ( .A(n50657), .B(n50658), .Z(n50656) );
  XOR U50510 ( .A(n50655), .B(n50628), .Z(n50658) );
  XNOR U50511 ( .A(n50659), .B(n50660), .Z(n50480) );
  AND U50512 ( .A(n1884), .B(n50661), .Z(n50660) );
  XNOR U50513 ( .A(n50662), .B(n50663), .Z(n1884) );
  AND U50514 ( .A(n50664), .B(n50665), .Z(n50663) );
  XOR U50515 ( .A(n50662), .B(n50490), .Z(n50665) );
  XNOR U50516 ( .A(n50662), .B(n50450), .Z(n50664) );
  XOR U50517 ( .A(n50666), .B(n50667), .Z(n50662) );
  AND U50518 ( .A(n50668), .B(n50669), .Z(n50667) );
  XOR U50519 ( .A(n50666), .B(n50458), .Z(n50668) );
  XOR U50520 ( .A(n50670), .B(n50671), .Z(n50441) );
  AND U50521 ( .A(n1888), .B(n50661), .Z(n50671) );
  XNOR U50522 ( .A(n50659), .B(n50670), .Z(n50661) );
  XNOR U50523 ( .A(n50672), .B(n50673), .Z(n1888) );
  AND U50524 ( .A(n50674), .B(n50675), .Z(n50673) );
  XNOR U50525 ( .A(n50676), .B(n50672), .Z(n50675) );
  IV U50526 ( .A(n50490), .Z(n50676) );
  XOR U50527 ( .A(n50646), .B(n50677), .Z(n50490) );
  AND U50528 ( .A(n1891), .B(n50678), .Z(n50677) );
  XOR U50529 ( .A(n50533), .B(n50530), .Z(n50678) );
  IV U50530 ( .A(n50646), .Z(n50533) );
  XNOR U50531 ( .A(n50450), .B(n50672), .Z(n50674) );
  XOR U50532 ( .A(n50679), .B(n50680), .Z(n50450) );
  AND U50533 ( .A(n1907), .B(n50681), .Z(n50680) );
  XOR U50534 ( .A(n50666), .B(n50682), .Z(n50672) );
  AND U50535 ( .A(n50683), .B(n50669), .Z(n50682) );
  XNOR U50536 ( .A(n50500), .B(n50666), .Z(n50669) );
  XOR U50537 ( .A(n50550), .B(n50684), .Z(n50500) );
  AND U50538 ( .A(n1891), .B(n50685), .Z(n50684) );
  XOR U50539 ( .A(n50546), .B(n50550), .Z(n50685) );
  XNOR U50540 ( .A(n50686), .B(n50666), .Z(n50683) );
  IV U50541 ( .A(n50458), .Z(n50686) );
  XOR U50542 ( .A(n50687), .B(n50688), .Z(n50458) );
  AND U50543 ( .A(n1907), .B(n50689), .Z(n50688) );
  XOR U50544 ( .A(n50690), .B(n50691), .Z(n50666) );
  AND U50545 ( .A(n50692), .B(n50693), .Z(n50691) );
  XNOR U50546 ( .A(n50510), .B(n50690), .Z(n50693) );
  XOR U50547 ( .A(n50578), .B(n50694), .Z(n50510) );
  AND U50548 ( .A(n1891), .B(n50695), .Z(n50694) );
  XOR U50549 ( .A(n50574), .B(n50578), .Z(n50695) );
  XOR U50550 ( .A(n50690), .B(n50467), .Z(n50692) );
  XOR U50551 ( .A(n50696), .B(n50697), .Z(n50467) );
  AND U50552 ( .A(n1907), .B(n50698), .Z(n50697) );
  XOR U50553 ( .A(n50699), .B(n50700), .Z(n50690) );
  AND U50554 ( .A(n50701), .B(n50702), .Z(n50700) );
  XNOR U50555 ( .A(n50699), .B(n50518), .Z(n50702) );
  XOR U50556 ( .A(n50629), .B(n50703), .Z(n50518) );
  AND U50557 ( .A(n1891), .B(n50704), .Z(n50703) );
  XOR U50558 ( .A(n50625), .B(n50629), .Z(n50704) );
  XNOR U50559 ( .A(n50705), .B(n50699), .Z(n50701) );
  IV U50560 ( .A(n50477), .Z(n50705) );
  XOR U50561 ( .A(n50706), .B(n50707), .Z(n50477) );
  AND U50562 ( .A(n1907), .B(n50708), .Z(n50707) );
  AND U50563 ( .A(n50670), .B(n50659), .Z(n50699) );
  XNOR U50564 ( .A(n50709), .B(n50710), .Z(n50659) );
  AND U50565 ( .A(n1891), .B(n50641), .Z(n50710) );
  XNOR U50566 ( .A(n50639), .B(n50709), .Z(n50641) );
  XNOR U50567 ( .A(n50711), .B(n50712), .Z(n1891) );
  AND U50568 ( .A(n50713), .B(n50714), .Z(n50712) );
  XNOR U50569 ( .A(n50711), .B(n50530), .Z(n50714) );
  IV U50570 ( .A(n50534), .Z(n50530) );
  XOR U50571 ( .A(n50715), .B(n50716), .Z(n50534) );
  AND U50572 ( .A(n1895), .B(n50717), .Z(n50716) );
  XOR U50573 ( .A(n50718), .B(n50715), .Z(n50717) );
  XNOR U50574 ( .A(n50711), .B(n50646), .Z(n50713) );
  XOR U50575 ( .A(n50719), .B(n50720), .Z(n50646) );
  AND U50576 ( .A(n1903), .B(n50681), .Z(n50720) );
  XOR U50577 ( .A(n50679), .B(n50719), .Z(n50681) );
  XOR U50578 ( .A(n50721), .B(n50722), .Z(n50711) );
  AND U50579 ( .A(n50723), .B(n50724), .Z(n50722) );
  XNOR U50580 ( .A(n50721), .B(n50546), .Z(n50724) );
  IV U50581 ( .A(n50549), .Z(n50546) );
  XOR U50582 ( .A(n50725), .B(n50726), .Z(n50549) );
  AND U50583 ( .A(n1895), .B(n50727), .Z(n50726) );
  XOR U50584 ( .A(n50728), .B(n50725), .Z(n50727) );
  XOR U50585 ( .A(n50550), .B(n50721), .Z(n50723) );
  XOR U50586 ( .A(n50729), .B(n50730), .Z(n50550) );
  AND U50587 ( .A(n1903), .B(n50689), .Z(n50730) );
  XOR U50588 ( .A(n50729), .B(n50687), .Z(n50689) );
  XOR U50589 ( .A(n50731), .B(n50732), .Z(n50721) );
  AND U50590 ( .A(n50733), .B(n50734), .Z(n50732) );
  XNOR U50591 ( .A(n50731), .B(n50574), .Z(n50734) );
  IV U50592 ( .A(n50577), .Z(n50574) );
  XOR U50593 ( .A(n50735), .B(n50736), .Z(n50577) );
  AND U50594 ( .A(n1895), .B(n50737), .Z(n50736) );
  XNOR U50595 ( .A(n50738), .B(n50735), .Z(n50737) );
  XOR U50596 ( .A(n50578), .B(n50731), .Z(n50733) );
  XOR U50597 ( .A(n50739), .B(n50740), .Z(n50578) );
  AND U50598 ( .A(n1903), .B(n50698), .Z(n50740) );
  XOR U50599 ( .A(n50739), .B(n50696), .Z(n50698) );
  XOR U50600 ( .A(n50655), .B(n50741), .Z(n50731) );
  AND U50601 ( .A(n50657), .B(n50742), .Z(n50741) );
  XNOR U50602 ( .A(n50655), .B(n50625), .Z(n50742) );
  IV U50603 ( .A(n50628), .Z(n50625) );
  XOR U50604 ( .A(n50743), .B(n50744), .Z(n50628) );
  AND U50605 ( .A(n1895), .B(n50745), .Z(n50744) );
  XOR U50606 ( .A(n50746), .B(n50743), .Z(n50745) );
  XOR U50607 ( .A(n50629), .B(n50655), .Z(n50657) );
  XOR U50608 ( .A(n50747), .B(n50748), .Z(n50629) );
  AND U50609 ( .A(n1903), .B(n50708), .Z(n50748) );
  XOR U50610 ( .A(n50747), .B(n50706), .Z(n50708) );
  AND U50611 ( .A(n50709), .B(n50639), .Z(n50655) );
  XNOR U50612 ( .A(n50749), .B(n50750), .Z(n50639) );
  AND U50613 ( .A(n1895), .B(n50751), .Z(n50750) );
  XNOR U50614 ( .A(n50752), .B(n50749), .Z(n50751) );
  XNOR U50615 ( .A(n50753), .B(n50754), .Z(n1895) );
  AND U50616 ( .A(n50755), .B(n50756), .Z(n50754) );
  XOR U50617 ( .A(n50718), .B(n50753), .Z(n50756) );
  AND U50618 ( .A(n50757), .B(n50758), .Z(n50718) );
  XNOR U50619 ( .A(n50715), .B(n50753), .Z(n50755) );
  XNOR U50620 ( .A(n50759), .B(n50760), .Z(n50715) );
  AND U50621 ( .A(n1899), .B(n50761), .Z(n50760) );
  XNOR U50622 ( .A(n50762), .B(n50763), .Z(n50761) );
  XOR U50623 ( .A(n50764), .B(n50765), .Z(n50753) );
  AND U50624 ( .A(n50766), .B(n50767), .Z(n50765) );
  XNOR U50625 ( .A(n50764), .B(n50757), .Z(n50767) );
  IV U50626 ( .A(n50728), .Z(n50757) );
  XOR U50627 ( .A(n50768), .B(n50769), .Z(n50728) );
  XOR U50628 ( .A(n50770), .B(n50758), .Z(n50769) );
  AND U50629 ( .A(n50738), .B(n50771), .Z(n50758) );
  AND U50630 ( .A(n50772), .B(n50773), .Z(n50770) );
  XOR U50631 ( .A(n50774), .B(n50768), .Z(n50772) );
  XNOR U50632 ( .A(n50725), .B(n50764), .Z(n50766) );
  XNOR U50633 ( .A(n50775), .B(n50776), .Z(n50725) );
  AND U50634 ( .A(n1899), .B(n50777), .Z(n50776) );
  XNOR U50635 ( .A(n50778), .B(n50779), .Z(n50777) );
  XOR U50636 ( .A(n50780), .B(n50781), .Z(n50764) );
  AND U50637 ( .A(n50782), .B(n50783), .Z(n50781) );
  XNOR U50638 ( .A(n50780), .B(n50738), .Z(n50783) );
  XOR U50639 ( .A(n50784), .B(n50773), .Z(n50738) );
  XNOR U50640 ( .A(n50785), .B(n50768), .Z(n50773) );
  XOR U50641 ( .A(n50786), .B(n50787), .Z(n50768) );
  AND U50642 ( .A(n50788), .B(n50789), .Z(n50787) );
  XOR U50643 ( .A(n50790), .B(n50786), .Z(n50788) );
  XNOR U50644 ( .A(n50791), .B(n50792), .Z(n50785) );
  AND U50645 ( .A(n50793), .B(n50794), .Z(n50792) );
  XOR U50646 ( .A(n50791), .B(n50795), .Z(n50793) );
  XNOR U50647 ( .A(n50774), .B(n50771), .Z(n50784) );
  AND U50648 ( .A(n50796), .B(n50797), .Z(n50771) );
  XOR U50649 ( .A(n50798), .B(n50799), .Z(n50774) );
  AND U50650 ( .A(n50800), .B(n50801), .Z(n50799) );
  XOR U50651 ( .A(n50798), .B(n50802), .Z(n50800) );
  XNOR U50652 ( .A(n50735), .B(n50780), .Z(n50782) );
  XNOR U50653 ( .A(n50803), .B(n50804), .Z(n50735) );
  AND U50654 ( .A(n1899), .B(n50805), .Z(n50804) );
  XNOR U50655 ( .A(n50806), .B(n50807), .Z(n50805) );
  XOR U50656 ( .A(n50808), .B(n50809), .Z(n50780) );
  AND U50657 ( .A(n50810), .B(n50811), .Z(n50809) );
  XNOR U50658 ( .A(n50808), .B(n50796), .Z(n50811) );
  IV U50659 ( .A(n50746), .Z(n50796) );
  XNOR U50660 ( .A(n50812), .B(n50789), .Z(n50746) );
  XNOR U50661 ( .A(n50813), .B(n50795), .Z(n50789) );
  XNOR U50662 ( .A(n50814), .B(n50815), .Z(n50795) );
  NOR U50663 ( .A(n50816), .B(n50817), .Z(n50815) );
  XOR U50664 ( .A(n50814), .B(n50818), .Z(n50816) );
  XNOR U50665 ( .A(n50794), .B(n50786), .Z(n50813) );
  XOR U50666 ( .A(n50819), .B(n50820), .Z(n50786) );
  AND U50667 ( .A(n50821), .B(n50822), .Z(n50820) );
  XOR U50668 ( .A(n50819), .B(n50823), .Z(n50821) );
  XNOR U50669 ( .A(n50824), .B(n50791), .Z(n50794) );
  XOR U50670 ( .A(n50825), .B(n50826), .Z(n50791) );
  AND U50671 ( .A(n50827), .B(n50828), .Z(n50826) );
  XNOR U50672 ( .A(n50829), .B(n50830), .Z(n50827) );
  IV U50673 ( .A(n50825), .Z(n50829) );
  XNOR U50674 ( .A(n50831), .B(n50832), .Z(n50824) );
  NOR U50675 ( .A(n50833), .B(n50834), .Z(n50832) );
  XNOR U50676 ( .A(n50831), .B(n50835), .Z(n50833) );
  XNOR U50677 ( .A(n50790), .B(n50797), .Z(n50812) );
  NOR U50678 ( .A(n50752), .B(n50836), .Z(n50797) );
  XOR U50679 ( .A(n50802), .B(n50801), .Z(n50790) );
  XNOR U50680 ( .A(n50837), .B(n50798), .Z(n50801) );
  XOR U50681 ( .A(n50838), .B(n50839), .Z(n50798) );
  AND U50682 ( .A(n50840), .B(n50841), .Z(n50839) );
  XNOR U50683 ( .A(n50842), .B(n50843), .Z(n50840) );
  IV U50684 ( .A(n50838), .Z(n50842) );
  XNOR U50685 ( .A(n50844), .B(n50845), .Z(n50837) );
  NOR U50686 ( .A(n50846), .B(n50847), .Z(n50845) );
  XNOR U50687 ( .A(n50844), .B(n50848), .Z(n50846) );
  XOR U50688 ( .A(n50849), .B(n50850), .Z(n50802) );
  NOR U50689 ( .A(n50851), .B(n50852), .Z(n50850) );
  XNOR U50690 ( .A(n50849), .B(n50853), .Z(n50851) );
  XNOR U50691 ( .A(n50743), .B(n50808), .Z(n50810) );
  XNOR U50692 ( .A(n50854), .B(n50855), .Z(n50743) );
  AND U50693 ( .A(n1899), .B(n50856), .Z(n50855) );
  XNOR U50694 ( .A(n50857), .B(n50858), .Z(n50856) );
  AND U50695 ( .A(n50749), .B(n50752), .Z(n50808) );
  XOR U50696 ( .A(n50859), .B(n50836), .Z(n50752) );
  XNOR U50697 ( .A(p_input[1536]), .B(p_input[2048]), .Z(n50836) );
  XNOR U50698 ( .A(n50823), .B(n50822), .Z(n50859) );
  XNOR U50699 ( .A(n50860), .B(n50830), .Z(n50822) );
  XNOR U50700 ( .A(n50818), .B(n50817), .Z(n50830) );
  XNOR U50701 ( .A(n50861), .B(n50814), .Z(n50817) );
  XNOR U50702 ( .A(p_input[1546]), .B(p_input[2058]), .Z(n50814) );
  XOR U50703 ( .A(p_input[1547]), .B(n29030), .Z(n50861) );
  XOR U50704 ( .A(p_input[1548]), .B(p_input[2060]), .Z(n50818) );
  XOR U50705 ( .A(n50828), .B(n50862), .Z(n50860) );
  IV U50706 ( .A(n50819), .Z(n50862) );
  XOR U50707 ( .A(p_input[1537]), .B(p_input[2049]), .Z(n50819) );
  XNOR U50708 ( .A(n50863), .B(n50835), .Z(n50828) );
  XNOR U50709 ( .A(p_input[1551]), .B(n29033), .Z(n50835) );
  XOR U50710 ( .A(n50825), .B(n50834), .Z(n50863) );
  XOR U50711 ( .A(n50864), .B(n50831), .Z(n50834) );
  XOR U50712 ( .A(p_input[1549]), .B(p_input[2061]), .Z(n50831) );
  XOR U50713 ( .A(p_input[1550]), .B(n29035), .Z(n50864) );
  XOR U50714 ( .A(p_input[1545]), .B(p_input[2057]), .Z(n50825) );
  XOR U50715 ( .A(n50843), .B(n50841), .Z(n50823) );
  XNOR U50716 ( .A(n50865), .B(n50848), .Z(n50841) );
  XOR U50717 ( .A(p_input[1544]), .B(p_input[2056]), .Z(n50848) );
  XOR U50718 ( .A(n50838), .B(n50847), .Z(n50865) );
  XOR U50719 ( .A(n50866), .B(n50844), .Z(n50847) );
  XOR U50720 ( .A(p_input[1542]), .B(p_input[2054]), .Z(n50844) );
  XOR U50721 ( .A(p_input[1543]), .B(n30404), .Z(n50866) );
  XOR U50722 ( .A(p_input[1538]), .B(p_input[2050]), .Z(n50838) );
  XNOR U50723 ( .A(n50853), .B(n50852), .Z(n50843) );
  XOR U50724 ( .A(n50867), .B(n50849), .Z(n50852) );
  XOR U50725 ( .A(p_input[1539]), .B(p_input[2051]), .Z(n50849) );
  XOR U50726 ( .A(p_input[1540]), .B(n30406), .Z(n50867) );
  XOR U50727 ( .A(p_input[1541]), .B(p_input[2053]), .Z(n50853) );
  XNOR U50728 ( .A(n50868), .B(n50869), .Z(n50749) );
  AND U50729 ( .A(n1899), .B(n50870), .Z(n50869) );
  XNOR U50730 ( .A(n50871), .B(n50872), .Z(n1899) );
  AND U50731 ( .A(n50873), .B(n50874), .Z(n50872) );
  XOR U50732 ( .A(n50763), .B(n50871), .Z(n50874) );
  XNOR U50733 ( .A(n50875), .B(n50871), .Z(n50873) );
  XOR U50734 ( .A(n50876), .B(n50877), .Z(n50871) );
  AND U50735 ( .A(n50878), .B(n50879), .Z(n50877) );
  XOR U50736 ( .A(n50778), .B(n50876), .Z(n50879) );
  XOR U50737 ( .A(n50876), .B(n50779), .Z(n50878) );
  XOR U50738 ( .A(n50880), .B(n50881), .Z(n50876) );
  AND U50739 ( .A(n50882), .B(n50883), .Z(n50881) );
  XOR U50740 ( .A(n50806), .B(n50880), .Z(n50883) );
  XOR U50741 ( .A(n50880), .B(n50807), .Z(n50882) );
  XOR U50742 ( .A(n50884), .B(n50885), .Z(n50880) );
  AND U50743 ( .A(n50886), .B(n50887), .Z(n50885) );
  XOR U50744 ( .A(n50884), .B(n50857), .Z(n50887) );
  XNOR U50745 ( .A(n50888), .B(n50889), .Z(n50709) );
  AND U50746 ( .A(n1903), .B(n50890), .Z(n50889) );
  XNOR U50747 ( .A(n50891), .B(n50892), .Z(n1903) );
  AND U50748 ( .A(n50893), .B(n50894), .Z(n50892) );
  XOR U50749 ( .A(n50891), .B(n50719), .Z(n50894) );
  XNOR U50750 ( .A(n50891), .B(n50679), .Z(n50893) );
  XOR U50751 ( .A(n50895), .B(n50896), .Z(n50891) );
  AND U50752 ( .A(n50897), .B(n50898), .Z(n50896) );
  XOR U50753 ( .A(n50895), .B(n50687), .Z(n50897) );
  XOR U50754 ( .A(n50899), .B(n50900), .Z(n50670) );
  AND U50755 ( .A(n1907), .B(n50890), .Z(n50900) );
  XNOR U50756 ( .A(n50888), .B(n50899), .Z(n50890) );
  XNOR U50757 ( .A(n50901), .B(n50902), .Z(n1907) );
  AND U50758 ( .A(n50903), .B(n50904), .Z(n50902) );
  XNOR U50759 ( .A(n50905), .B(n50901), .Z(n50904) );
  IV U50760 ( .A(n50719), .Z(n50905) );
  XOR U50761 ( .A(n50875), .B(n50906), .Z(n50719) );
  AND U50762 ( .A(n1910), .B(n50907), .Z(n50906) );
  XOR U50763 ( .A(n50762), .B(n50759), .Z(n50907) );
  IV U50764 ( .A(n50875), .Z(n50762) );
  XNOR U50765 ( .A(n50679), .B(n50901), .Z(n50903) );
  XOR U50766 ( .A(n50908), .B(n50909), .Z(n50679) );
  AND U50767 ( .A(n1926), .B(n50910), .Z(n50909) );
  XOR U50768 ( .A(n50895), .B(n50911), .Z(n50901) );
  AND U50769 ( .A(n50912), .B(n50898), .Z(n50911) );
  XNOR U50770 ( .A(n50729), .B(n50895), .Z(n50898) );
  XOR U50771 ( .A(n50779), .B(n50913), .Z(n50729) );
  AND U50772 ( .A(n1910), .B(n50914), .Z(n50913) );
  XOR U50773 ( .A(n50775), .B(n50779), .Z(n50914) );
  XNOR U50774 ( .A(n50915), .B(n50895), .Z(n50912) );
  IV U50775 ( .A(n50687), .Z(n50915) );
  XOR U50776 ( .A(n50916), .B(n50917), .Z(n50687) );
  AND U50777 ( .A(n1926), .B(n50918), .Z(n50917) );
  XOR U50778 ( .A(n50919), .B(n50920), .Z(n50895) );
  AND U50779 ( .A(n50921), .B(n50922), .Z(n50920) );
  XNOR U50780 ( .A(n50739), .B(n50919), .Z(n50922) );
  XOR U50781 ( .A(n50807), .B(n50923), .Z(n50739) );
  AND U50782 ( .A(n1910), .B(n50924), .Z(n50923) );
  XOR U50783 ( .A(n50803), .B(n50807), .Z(n50924) );
  XOR U50784 ( .A(n50919), .B(n50696), .Z(n50921) );
  XOR U50785 ( .A(n50925), .B(n50926), .Z(n50696) );
  AND U50786 ( .A(n1926), .B(n50927), .Z(n50926) );
  XOR U50787 ( .A(n50928), .B(n50929), .Z(n50919) );
  AND U50788 ( .A(n50930), .B(n50931), .Z(n50929) );
  XNOR U50789 ( .A(n50928), .B(n50747), .Z(n50931) );
  XOR U50790 ( .A(n50858), .B(n50932), .Z(n50747) );
  AND U50791 ( .A(n1910), .B(n50933), .Z(n50932) );
  XOR U50792 ( .A(n50854), .B(n50858), .Z(n50933) );
  XNOR U50793 ( .A(n50934), .B(n50928), .Z(n50930) );
  IV U50794 ( .A(n50706), .Z(n50934) );
  XOR U50795 ( .A(n50935), .B(n50936), .Z(n50706) );
  AND U50796 ( .A(n1926), .B(n50937), .Z(n50936) );
  AND U50797 ( .A(n50899), .B(n50888), .Z(n50928) );
  XNOR U50798 ( .A(n50938), .B(n50939), .Z(n50888) );
  AND U50799 ( .A(n1910), .B(n50870), .Z(n50939) );
  XNOR U50800 ( .A(n50868), .B(n50938), .Z(n50870) );
  XNOR U50801 ( .A(n50940), .B(n50941), .Z(n1910) );
  AND U50802 ( .A(n50942), .B(n50943), .Z(n50941) );
  XNOR U50803 ( .A(n50940), .B(n50759), .Z(n50943) );
  IV U50804 ( .A(n50763), .Z(n50759) );
  XOR U50805 ( .A(n50944), .B(n50945), .Z(n50763) );
  AND U50806 ( .A(n1914), .B(n50946), .Z(n50945) );
  XOR U50807 ( .A(n50947), .B(n50944), .Z(n50946) );
  XNOR U50808 ( .A(n50940), .B(n50875), .Z(n50942) );
  XOR U50809 ( .A(n50948), .B(n50949), .Z(n50875) );
  AND U50810 ( .A(n1922), .B(n50910), .Z(n50949) );
  XOR U50811 ( .A(n50908), .B(n50948), .Z(n50910) );
  XOR U50812 ( .A(n50950), .B(n50951), .Z(n50940) );
  AND U50813 ( .A(n50952), .B(n50953), .Z(n50951) );
  XNOR U50814 ( .A(n50950), .B(n50775), .Z(n50953) );
  IV U50815 ( .A(n50778), .Z(n50775) );
  XOR U50816 ( .A(n50954), .B(n50955), .Z(n50778) );
  AND U50817 ( .A(n1914), .B(n50956), .Z(n50955) );
  XOR U50818 ( .A(n50957), .B(n50954), .Z(n50956) );
  XOR U50819 ( .A(n50779), .B(n50950), .Z(n50952) );
  XOR U50820 ( .A(n50958), .B(n50959), .Z(n50779) );
  AND U50821 ( .A(n1922), .B(n50918), .Z(n50959) );
  XOR U50822 ( .A(n50958), .B(n50916), .Z(n50918) );
  XOR U50823 ( .A(n50960), .B(n50961), .Z(n50950) );
  AND U50824 ( .A(n50962), .B(n50963), .Z(n50961) );
  XNOR U50825 ( .A(n50960), .B(n50803), .Z(n50963) );
  IV U50826 ( .A(n50806), .Z(n50803) );
  XOR U50827 ( .A(n50964), .B(n50965), .Z(n50806) );
  AND U50828 ( .A(n1914), .B(n50966), .Z(n50965) );
  XNOR U50829 ( .A(n50967), .B(n50964), .Z(n50966) );
  XOR U50830 ( .A(n50807), .B(n50960), .Z(n50962) );
  XOR U50831 ( .A(n50968), .B(n50969), .Z(n50807) );
  AND U50832 ( .A(n1922), .B(n50927), .Z(n50969) );
  XOR U50833 ( .A(n50968), .B(n50925), .Z(n50927) );
  XOR U50834 ( .A(n50884), .B(n50970), .Z(n50960) );
  AND U50835 ( .A(n50886), .B(n50971), .Z(n50970) );
  XNOR U50836 ( .A(n50884), .B(n50854), .Z(n50971) );
  IV U50837 ( .A(n50857), .Z(n50854) );
  XOR U50838 ( .A(n50972), .B(n50973), .Z(n50857) );
  AND U50839 ( .A(n1914), .B(n50974), .Z(n50973) );
  XOR U50840 ( .A(n50975), .B(n50972), .Z(n50974) );
  XOR U50841 ( .A(n50858), .B(n50884), .Z(n50886) );
  XOR U50842 ( .A(n50976), .B(n50977), .Z(n50858) );
  AND U50843 ( .A(n1922), .B(n50937), .Z(n50977) );
  XOR U50844 ( .A(n50976), .B(n50935), .Z(n50937) );
  AND U50845 ( .A(n50938), .B(n50868), .Z(n50884) );
  XNOR U50846 ( .A(n50978), .B(n50979), .Z(n50868) );
  AND U50847 ( .A(n1914), .B(n50980), .Z(n50979) );
  XNOR U50848 ( .A(n50981), .B(n50978), .Z(n50980) );
  XNOR U50849 ( .A(n50982), .B(n50983), .Z(n1914) );
  AND U50850 ( .A(n50984), .B(n50985), .Z(n50983) );
  XOR U50851 ( .A(n50947), .B(n50982), .Z(n50985) );
  AND U50852 ( .A(n50986), .B(n50987), .Z(n50947) );
  XNOR U50853 ( .A(n50944), .B(n50982), .Z(n50984) );
  XNOR U50854 ( .A(n50988), .B(n50989), .Z(n50944) );
  AND U50855 ( .A(n1918), .B(n50990), .Z(n50989) );
  XNOR U50856 ( .A(n50991), .B(n50992), .Z(n50990) );
  XOR U50857 ( .A(n50993), .B(n50994), .Z(n50982) );
  AND U50858 ( .A(n50995), .B(n50996), .Z(n50994) );
  XNOR U50859 ( .A(n50993), .B(n50986), .Z(n50996) );
  IV U50860 ( .A(n50957), .Z(n50986) );
  XOR U50861 ( .A(n50997), .B(n50998), .Z(n50957) );
  XOR U50862 ( .A(n50999), .B(n50987), .Z(n50998) );
  AND U50863 ( .A(n50967), .B(n51000), .Z(n50987) );
  AND U50864 ( .A(n51001), .B(n51002), .Z(n50999) );
  XOR U50865 ( .A(n51003), .B(n50997), .Z(n51001) );
  XNOR U50866 ( .A(n50954), .B(n50993), .Z(n50995) );
  XNOR U50867 ( .A(n51004), .B(n51005), .Z(n50954) );
  AND U50868 ( .A(n1918), .B(n51006), .Z(n51005) );
  XNOR U50869 ( .A(n51007), .B(n51008), .Z(n51006) );
  XOR U50870 ( .A(n51009), .B(n51010), .Z(n50993) );
  AND U50871 ( .A(n51011), .B(n51012), .Z(n51010) );
  XNOR U50872 ( .A(n51009), .B(n50967), .Z(n51012) );
  XOR U50873 ( .A(n51013), .B(n51002), .Z(n50967) );
  XNOR U50874 ( .A(n51014), .B(n50997), .Z(n51002) );
  XOR U50875 ( .A(n51015), .B(n51016), .Z(n50997) );
  AND U50876 ( .A(n51017), .B(n51018), .Z(n51016) );
  XOR U50877 ( .A(n51019), .B(n51015), .Z(n51017) );
  XNOR U50878 ( .A(n51020), .B(n51021), .Z(n51014) );
  AND U50879 ( .A(n51022), .B(n51023), .Z(n51021) );
  XOR U50880 ( .A(n51020), .B(n51024), .Z(n51022) );
  XNOR U50881 ( .A(n51003), .B(n51000), .Z(n51013) );
  AND U50882 ( .A(n51025), .B(n51026), .Z(n51000) );
  XOR U50883 ( .A(n51027), .B(n51028), .Z(n51003) );
  AND U50884 ( .A(n51029), .B(n51030), .Z(n51028) );
  XOR U50885 ( .A(n51027), .B(n51031), .Z(n51029) );
  XNOR U50886 ( .A(n50964), .B(n51009), .Z(n51011) );
  XNOR U50887 ( .A(n51032), .B(n51033), .Z(n50964) );
  AND U50888 ( .A(n1918), .B(n51034), .Z(n51033) );
  XNOR U50889 ( .A(n51035), .B(n51036), .Z(n51034) );
  XOR U50890 ( .A(n51037), .B(n51038), .Z(n51009) );
  AND U50891 ( .A(n51039), .B(n51040), .Z(n51038) );
  XNOR U50892 ( .A(n51037), .B(n51025), .Z(n51040) );
  IV U50893 ( .A(n50975), .Z(n51025) );
  XNOR U50894 ( .A(n51041), .B(n51018), .Z(n50975) );
  XNOR U50895 ( .A(n51042), .B(n51024), .Z(n51018) );
  XNOR U50896 ( .A(n51043), .B(n51044), .Z(n51024) );
  NOR U50897 ( .A(n51045), .B(n51046), .Z(n51044) );
  XOR U50898 ( .A(n51043), .B(n51047), .Z(n51045) );
  XNOR U50899 ( .A(n51023), .B(n51015), .Z(n51042) );
  XOR U50900 ( .A(n51048), .B(n51049), .Z(n51015) );
  AND U50901 ( .A(n51050), .B(n51051), .Z(n51049) );
  XOR U50902 ( .A(n51048), .B(n51052), .Z(n51050) );
  XNOR U50903 ( .A(n51053), .B(n51020), .Z(n51023) );
  XOR U50904 ( .A(n51054), .B(n51055), .Z(n51020) );
  AND U50905 ( .A(n51056), .B(n51057), .Z(n51055) );
  XNOR U50906 ( .A(n51058), .B(n51059), .Z(n51056) );
  IV U50907 ( .A(n51054), .Z(n51058) );
  XNOR U50908 ( .A(n51060), .B(n51061), .Z(n51053) );
  NOR U50909 ( .A(n51062), .B(n51063), .Z(n51061) );
  XNOR U50910 ( .A(n51060), .B(n51064), .Z(n51062) );
  XNOR U50911 ( .A(n51019), .B(n51026), .Z(n51041) );
  NOR U50912 ( .A(n50981), .B(n51065), .Z(n51026) );
  XOR U50913 ( .A(n51031), .B(n51030), .Z(n51019) );
  XNOR U50914 ( .A(n51066), .B(n51027), .Z(n51030) );
  XOR U50915 ( .A(n51067), .B(n51068), .Z(n51027) );
  AND U50916 ( .A(n51069), .B(n51070), .Z(n51068) );
  XNOR U50917 ( .A(n51071), .B(n51072), .Z(n51069) );
  IV U50918 ( .A(n51067), .Z(n51071) );
  XNOR U50919 ( .A(n51073), .B(n51074), .Z(n51066) );
  NOR U50920 ( .A(n51075), .B(n51076), .Z(n51074) );
  XNOR U50921 ( .A(n51073), .B(n51077), .Z(n51075) );
  XOR U50922 ( .A(n51078), .B(n51079), .Z(n51031) );
  NOR U50923 ( .A(n51080), .B(n51081), .Z(n51079) );
  XNOR U50924 ( .A(n51078), .B(n51082), .Z(n51080) );
  XNOR U50925 ( .A(n50972), .B(n51037), .Z(n51039) );
  XNOR U50926 ( .A(n51083), .B(n51084), .Z(n50972) );
  AND U50927 ( .A(n1918), .B(n51085), .Z(n51084) );
  XNOR U50928 ( .A(n51086), .B(n51087), .Z(n51085) );
  AND U50929 ( .A(n50978), .B(n50981), .Z(n51037) );
  XOR U50930 ( .A(n51088), .B(n51065), .Z(n50981) );
  XNOR U50931 ( .A(p_input[1552]), .B(p_input[2048]), .Z(n51065) );
  XNOR U50932 ( .A(n51052), .B(n51051), .Z(n51088) );
  XNOR U50933 ( .A(n51089), .B(n51059), .Z(n51051) );
  XNOR U50934 ( .A(n51047), .B(n51046), .Z(n51059) );
  XNOR U50935 ( .A(n51090), .B(n51043), .Z(n51046) );
  XNOR U50936 ( .A(p_input[1562]), .B(p_input[2058]), .Z(n51043) );
  XOR U50937 ( .A(p_input[1563]), .B(n29030), .Z(n51090) );
  XOR U50938 ( .A(p_input[1564]), .B(p_input[2060]), .Z(n51047) );
  XOR U50939 ( .A(n51057), .B(n51091), .Z(n51089) );
  IV U50940 ( .A(n51048), .Z(n51091) );
  XOR U50941 ( .A(p_input[1553]), .B(p_input[2049]), .Z(n51048) );
  XNOR U50942 ( .A(n51092), .B(n51064), .Z(n51057) );
  XNOR U50943 ( .A(p_input[1567]), .B(n29033), .Z(n51064) );
  XOR U50944 ( .A(n51054), .B(n51063), .Z(n51092) );
  XOR U50945 ( .A(n51093), .B(n51060), .Z(n51063) );
  XOR U50946 ( .A(p_input[1565]), .B(p_input[2061]), .Z(n51060) );
  XOR U50947 ( .A(p_input[1566]), .B(n29035), .Z(n51093) );
  XOR U50948 ( .A(p_input[1561]), .B(p_input[2057]), .Z(n51054) );
  XOR U50949 ( .A(n51072), .B(n51070), .Z(n51052) );
  XNOR U50950 ( .A(n51094), .B(n51077), .Z(n51070) );
  XOR U50951 ( .A(p_input[1560]), .B(p_input[2056]), .Z(n51077) );
  XOR U50952 ( .A(n51067), .B(n51076), .Z(n51094) );
  XOR U50953 ( .A(n51095), .B(n51073), .Z(n51076) );
  XOR U50954 ( .A(p_input[1558]), .B(p_input[2054]), .Z(n51073) );
  XOR U50955 ( .A(p_input[1559]), .B(n30404), .Z(n51095) );
  XOR U50956 ( .A(p_input[1554]), .B(p_input[2050]), .Z(n51067) );
  XNOR U50957 ( .A(n51082), .B(n51081), .Z(n51072) );
  XOR U50958 ( .A(n51096), .B(n51078), .Z(n51081) );
  XOR U50959 ( .A(p_input[1555]), .B(p_input[2051]), .Z(n51078) );
  XOR U50960 ( .A(p_input[1556]), .B(n30406), .Z(n51096) );
  XOR U50961 ( .A(p_input[1557]), .B(p_input[2053]), .Z(n51082) );
  XNOR U50962 ( .A(n51097), .B(n51098), .Z(n50978) );
  AND U50963 ( .A(n1918), .B(n51099), .Z(n51098) );
  XNOR U50964 ( .A(n51100), .B(n51101), .Z(n1918) );
  AND U50965 ( .A(n51102), .B(n51103), .Z(n51101) );
  XOR U50966 ( .A(n50992), .B(n51100), .Z(n51103) );
  XNOR U50967 ( .A(n51104), .B(n51100), .Z(n51102) );
  XOR U50968 ( .A(n51105), .B(n51106), .Z(n51100) );
  AND U50969 ( .A(n51107), .B(n51108), .Z(n51106) );
  XOR U50970 ( .A(n51007), .B(n51105), .Z(n51108) );
  XOR U50971 ( .A(n51105), .B(n51008), .Z(n51107) );
  XOR U50972 ( .A(n51109), .B(n51110), .Z(n51105) );
  AND U50973 ( .A(n51111), .B(n51112), .Z(n51110) );
  XOR U50974 ( .A(n51035), .B(n51109), .Z(n51112) );
  XOR U50975 ( .A(n51109), .B(n51036), .Z(n51111) );
  XOR U50976 ( .A(n51113), .B(n51114), .Z(n51109) );
  AND U50977 ( .A(n51115), .B(n51116), .Z(n51114) );
  XOR U50978 ( .A(n51113), .B(n51086), .Z(n51116) );
  XNOR U50979 ( .A(n51117), .B(n51118), .Z(n50938) );
  AND U50980 ( .A(n1922), .B(n51119), .Z(n51118) );
  XNOR U50981 ( .A(n51120), .B(n51121), .Z(n1922) );
  AND U50982 ( .A(n51122), .B(n51123), .Z(n51121) );
  XOR U50983 ( .A(n51120), .B(n50948), .Z(n51123) );
  XNOR U50984 ( .A(n51120), .B(n50908), .Z(n51122) );
  XOR U50985 ( .A(n51124), .B(n51125), .Z(n51120) );
  AND U50986 ( .A(n51126), .B(n51127), .Z(n51125) );
  XOR U50987 ( .A(n51124), .B(n50916), .Z(n51126) );
  XOR U50988 ( .A(n51128), .B(n51129), .Z(n50899) );
  AND U50989 ( .A(n1926), .B(n51119), .Z(n51129) );
  XNOR U50990 ( .A(n51117), .B(n51128), .Z(n51119) );
  XNOR U50991 ( .A(n51130), .B(n51131), .Z(n1926) );
  AND U50992 ( .A(n51132), .B(n51133), .Z(n51131) );
  XNOR U50993 ( .A(n51134), .B(n51130), .Z(n51133) );
  IV U50994 ( .A(n50948), .Z(n51134) );
  XOR U50995 ( .A(n51104), .B(n51135), .Z(n50948) );
  AND U50996 ( .A(n1929), .B(n51136), .Z(n51135) );
  XOR U50997 ( .A(n50991), .B(n50988), .Z(n51136) );
  IV U50998 ( .A(n51104), .Z(n50991) );
  XNOR U50999 ( .A(n50908), .B(n51130), .Z(n51132) );
  XOR U51000 ( .A(n51137), .B(n51138), .Z(n50908) );
  AND U51001 ( .A(n1945), .B(n51139), .Z(n51138) );
  XOR U51002 ( .A(n51124), .B(n51140), .Z(n51130) );
  AND U51003 ( .A(n51141), .B(n51127), .Z(n51140) );
  XNOR U51004 ( .A(n50958), .B(n51124), .Z(n51127) );
  XOR U51005 ( .A(n51008), .B(n51142), .Z(n50958) );
  AND U51006 ( .A(n1929), .B(n51143), .Z(n51142) );
  XOR U51007 ( .A(n51004), .B(n51008), .Z(n51143) );
  XNOR U51008 ( .A(n51144), .B(n51124), .Z(n51141) );
  IV U51009 ( .A(n50916), .Z(n51144) );
  XOR U51010 ( .A(n51145), .B(n51146), .Z(n50916) );
  AND U51011 ( .A(n1945), .B(n51147), .Z(n51146) );
  XOR U51012 ( .A(n51148), .B(n51149), .Z(n51124) );
  AND U51013 ( .A(n51150), .B(n51151), .Z(n51149) );
  XNOR U51014 ( .A(n50968), .B(n51148), .Z(n51151) );
  XOR U51015 ( .A(n51036), .B(n51152), .Z(n50968) );
  AND U51016 ( .A(n1929), .B(n51153), .Z(n51152) );
  XOR U51017 ( .A(n51032), .B(n51036), .Z(n51153) );
  XOR U51018 ( .A(n51148), .B(n50925), .Z(n51150) );
  XOR U51019 ( .A(n51154), .B(n51155), .Z(n50925) );
  AND U51020 ( .A(n1945), .B(n51156), .Z(n51155) );
  XOR U51021 ( .A(n51157), .B(n51158), .Z(n51148) );
  AND U51022 ( .A(n51159), .B(n51160), .Z(n51158) );
  XNOR U51023 ( .A(n51157), .B(n50976), .Z(n51160) );
  XOR U51024 ( .A(n51087), .B(n51161), .Z(n50976) );
  AND U51025 ( .A(n1929), .B(n51162), .Z(n51161) );
  XOR U51026 ( .A(n51083), .B(n51087), .Z(n51162) );
  XNOR U51027 ( .A(n51163), .B(n51157), .Z(n51159) );
  IV U51028 ( .A(n50935), .Z(n51163) );
  XOR U51029 ( .A(n51164), .B(n51165), .Z(n50935) );
  AND U51030 ( .A(n1945), .B(n51166), .Z(n51165) );
  AND U51031 ( .A(n51128), .B(n51117), .Z(n51157) );
  XNOR U51032 ( .A(n51167), .B(n51168), .Z(n51117) );
  AND U51033 ( .A(n1929), .B(n51099), .Z(n51168) );
  XNOR U51034 ( .A(n51097), .B(n51167), .Z(n51099) );
  XNOR U51035 ( .A(n51169), .B(n51170), .Z(n1929) );
  AND U51036 ( .A(n51171), .B(n51172), .Z(n51170) );
  XNOR U51037 ( .A(n51169), .B(n50988), .Z(n51172) );
  IV U51038 ( .A(n50992), .Z(n50988) );
  XOR U51039 ( .A(n51173), .B(n51174), .Z(n50992) );
  AND U51040 ( .A(n1933), .B(n51175), .Z(n51174) );
  XOR U51041 ( .A(n51176), .B(n51173), .Z(n51175) );
  XNOR U51042 ( .A(n51169), .B(n51104), .Z(n51171) );
  XOR U51043 ( .A(n51177), .B(n51178), .Z(n51104) );
  AND U51044 ( .A(n1941), .B(n51139), .Z(n51178) );
  XOR U51045 ( .A(n51137), .B(n51177), .Z(n51139) );
  XOR U51046 ( .A(n51179), .B(n51180), .Z(n51169) );
  AND U51047 ( .A(n51181), .B(n51182), .Z(n51180) );
  XNOR U51048 ( .A(n51179), .B(n51004), .Z(n51182) );
  IV U51049 ( .A(n51007), .Z(n51004) );
  XOR U51050 ( .A(n51183), .B(n51184), .Z(n51007) );
  AND U51051 ( .A(n1933), .B(n51185), .Z(n51184) );
  XOR U51052 ( .A(n51186), .B(n51183), .Z(n51185) );
  XOR U51053 ( .A(n51008), .B(n51179), .Z(n51181) );
  XOR U51054 ( .A(n51187), .B(n51188), .Z(n51008) );
  AND U51055 ( .A(n1941), .B(n51147), .Z(n51188) );
  XOR U51056 ( .A(n51187), .B(n51145), .Z(n51147) );
  XOR U51057 ( .A(n51189), .B(n51190), .Z(n51179) );
  AND U51058 ( .A(n51191), .B(n51192), .Z(n51190) );
  XNOR U51059 ( .A(n51189), .B(n51032), .Z(n51192) );
  IV U51060 ( .A(n51035), .Z(n51032) );
  XOR U51061 ( .A(n51193), .B(n51194), .Z(n51035) );
  AND U51062 ( .A(n1933), .B(n51195), .Z(n51194) );
  XNOR U51063 ( .A(n51196), .B(n51193), .Z(n51195) );
  XOR U51064 ( .A(n51036), .B(n51189), .Z(n51191) );
  XOR U51065 ( .A(n51197), .B(n51198), .Z(n51036) );
  AND U51066 ( .A(n1941), .B(n51156), .Z(n51198) );
  XOR U51067 ( .A(n51197), .B(n51154), .Z(n51156) );
  XOR U51068 ( .A(n51113), .B(n51199), .Z(n51189) );
  AND U51069 ( .A(n51115), .B(n51200), .Z(n51199) );
  XNOR U51070 ( .A(n51113), .B(n51083), .Z(n51200) );
  IV U51071 ( .A(n51086), .Z(n51083) );
  XOR U51072 ( .A(n51201), .B(n51202), .Z(n51086) );
  AND U51073 ( .A(n1933), .B(n51203), .Z(n51202) );
  XOR U51074 ( .A(n51204), .B(n51201), .Z(n51203) );
  XOR U51075 ( .A(n51087), .B(n51113), .Z(n51115) );
  XOR U51076 ( .A(n51205), .B(n51206), .Z(n51087) );
  AND U51077 ( .A(n1941), .B(n51166), .Z(n51206) );
  XOR U51078 ( .A(n51205), .B(n51164), .Z(n51166) );
  AND U51079 ( .A(n51167), .B(n51097), .Z(n51113) );
  XNOR U51080 ( .A(n51207), .B(n51208), .Z(n51097) );
  AND U51081 ( .A(n1933), .B(n51209), .Z(n51208) );
  XNOR U51082 ( .A(n51210), .B(n51207), .Z(n51209) );
  XNOR U51083 ( .A(n51211), .B(n51212), .Z(n1933) );
  AND U51084 ( .A(n51213), .B(n51214), .Z(n51212) );
  XOR U51085 ( .A(n51176), .B(n51211), .Z(n51214) );
  AND U51086 ( .A(n51215), .B(n51216), .Z(n51176) );
  XNOR U51087 ( .A(n51173), .B(n51211), .Z(n51213) );
  XNOR U51088 ( .A(n51217), .B(n51218), .Z(n51173) );
  AND U51089 ( .A(n1937), .B(n51219), .Z(n51218) );
  XNOR U51090 ( .A(n51220), .B(n51221), .Z(n51219) );
  XOR U51091 ( .A(n51222), .B(n51223), .Z(n51211) );
  AND U51092 ( .A(n51224), .B(n51225), .Z(n51223) );
  XNOR U51093 ( .A(n51222), .B(n51215), .Z(n51225) );
  IV U51094 ( .A(n51186), .Z(n51215) );
  XOR U51095 ( .A(n51226), .B(n51227), .Z(n51186) );
  XOR U51096 ( .A(n51228), .B(n51216), .Z(n51227) );
  AND U51097 ( .A(n51196), .B(n51229), .Z(n51216) );
  AND U51098 ( .A(n51230), .B(n51231), .Z(n51228) );
  XOR U51099 ( .A(n51232), .B(n51226), .Z(n51230) );
  XNOR U51100 ( .A(n51183), .B(n51222), .Z(n51224) );
  XNOR U51101 ( .A(n51233), .B(n51234), .Z(n51183) );
  AND U51102 ( .A(n1937), .B(n51235), .Z(n51234) );
  XNOR U51103 ( .A(n51236), .B(n51237), .Z(n51235) );
  XOR U51104 ( .A(n51238), .B(n51239), .Z(n51222) );
  AND U51105 ( .A(n51240), .B(n51241), .Z(n51239) );
  XNOR U51106 ( .A(n51238), .B(n51196), .Z(n51241) );
  XOR U51107 ( .A(n51242), .B(n51231), .Z(n51196) );
  XNOR U51108 ( .A(n51243), .B(n51226), .Z(n51231) );
  XOR U51109 ( .A(n51244), .B(n51245), .Z(n51226) );
  AND U51110 ( .A(n51246), .B(n51247), .Z(n51245) );
  XOR U51111 ( .A(n51248), .B(n51244), .Z(n51246) );
  XNOR U51112 ( .A(n51249), .B(n51250), .Z(n51243) );
  AND U51113 ( .A(n51251), .B(n51252), .Z(n51250) );
  XOR U51114 ( .A(n51249), .B(n51253), .Z(n51251) );
  XNOR U51115 ( .A(n51232), .B(n51229), .Z(n51242) );
  AND U51116 ( .A(n51254), .B(n51255), .Z(n51229) );
  XOR U51117 ( .A(n51256), .B(n51257), .Z(n51232) );
  AND U51118 ( .A(n51258), .B(n51259), .Z(n51257) );
  XOR U51119 ( .A(n51256), .B(n51260), .Z(n51258) );
  XNOR U51120 ( .A(n51193), .B(n51238), .Z(n51240) );
  XNOR U51121 ( .A(n51261), .B(n51262), .Z(n51193) );
  AND U51122 ( .A(n1937), .B(n51263), .Z(n51262) );
  XNOR U51123 ( .A(n51264), .B(n51265), .Z(n51263) );
  XOR U51124 ( .A(n51266), .B(n51267), .Z(n51238) );
  AND U51125 ( .A(n51268), .B(n51269), .Z(n51267) );
  XNOR U51126 ( .A(n51266), .B(n51254), .Z(n51269) );
  IV U51127 ( .A(n51204), .Z(n51254) );
  XNOR U51128 ( .A(n51270), .B(n51247), .Z(n51204) );
  XNOR U51129 ( .A(n51271), .B(n51253), .Z(n51247) );
  XNOR U51130 ( .A(n51272), .B(n51273), .Z(n51253) );
  NOR U51131 ( .A(n51274), .B(n51275), .Z(n51273) );
  XOR U51132 ( .A(n51272), .B(n51276), .Z(n51274) );
  XNOR U51133 ( .A(n51252), .B(n51244), .Z(n51271) );
  XOR U51134 ( .A(n51277), .B(n51278), .Z(n51244) );
  AND U51135 ( .A(n51279), .B(n51280), .Z(n51278) );
  XOR U51136 ( .A(n51277), .B(n51281), .Z(n51279) );
  XNOR U51137 ( .A(n51282), .B(n51249), .Z(n51252) );
  XOR U51138 ( .A(n51283), .B(n51284), .Z(n51249) );
  AND U51139 ( .A(n51285), .B(n51286), .Z(n51284) );
  XNOR U51140 ( .A(n51287), .B(n51288), .Z(n51285) );
  IV U51141 ( .A(n51283), .Z(n51287) );
  XNOR U51142 ( .A(n51289), .B(n51290), .Z(n51282) );
  NOR U51143 ( .A(n51291), .B(n51292), .Z(n51290) );
  XNOR U51144 ( .A(n51289), .B(n51293), .Z(n51291) );
  XNOR U51145 ( .A(n51248), .B(n51255), .Z(n51270) );
  NOR U51146 ( .A(n51210), .B(n51294), .Z(n51255) );
  XOR U51147 ( .A(n51260), .B(n51259), .Z(n51248) );
  XNOR U51148 ( .A(n51295), .B(n51256), .Z(n51259) );
  XOR U51149 ( .A(n51296), .B(n51297), .Z(n51256) );
  AND U51150 ( .A(n51298), .B(n51299), .Z(n51297) );
  XNOR U51151 ( .A(n51300), .B(n51301), .Z(n51298) );
  IV U51152 ( .A(n51296), .Z(n51300) );
  XNOR U51153 ( .A(n51302), .B(n51303), .Z(n51295) );
  NOR U51154 ( .A(n51304), .B(n51305), .Z(n51303) );
  XNOR U51155 ( .A(n51302), .B(n51306), .Z(n51304) );
  XOR U51156 ( .A(n51307), .B(n51308), .Z(n51260) );
  NOR U51157 ( .A(n51309), .B(n51310), .Z(n51308) );
  XNOR U51158 ( .A(n51307), .B(n51311), .Z(n51309) );
  XNOR U51159 ( .A(n51201), .B(n51266), .Z(n51268) );
  XNOR U51160 ( .A(n51312), .B(n51313), .Z(n51201) );
  AND U51161 ( .A(n1937), .B(n51314), .Z(n51313) );
  XNOR U51162 ( .A(n51315), .B(n51316), .Z(n51314) );
  AND U51163 ( .A(n51207), .B(n51210), .Z(n51266) );
  XOR U51164 ( .A(n51317), .B(n51294), .Z(n51210) );
  XNOR U51165 ( .A(p_input[1568]), .B(p_input[2048]), .Z(n51294) );
  XNOR U51166 ( .A(n51281), .B(n51280), .Z(n51317) );
  XNOR U51167 ( .A(n51318), .B(n51288), .Z(n51280) );
  XNOR U51168 ( .A(n51276), .B(n51275), .Z(n51288) );
  XNOR U51169 ( .A(n51319), .B(n51272), .Z(n51275) );
  XNOR U51170 ( .A(p_input[1578]), .B(p_input[2058]), .Z(n51272) );
  XOR U51171 ( .A(p_input[1579]), .B(n29030), .Z(n51319) );
  XOR U51172 ( .A(p_input[1580]), .B(p_input[2060]), .Z(n51276) );
  XOR U51173 ( .A(n51286), .B(n51320), .Z(n51318) );
  IV U51174 ( .A(n51277), .Z(n51320) );
  XOR U51175 ( .A(p_input[1569]), .B(p_input[2049]), .Z(n51277) );
  XNOR U51176 ( .A(n51321), .B(n51293), .Z(n51286) );
  XNOR U51177 ( .A(p_input[1583]), .B(n29033), .Z(n51293) );
  XOR U51178 ( .A(n51283), .B(n51292), .Z(n51321) );
  XOR U51179 ( .A(n51322), .B(n51289), .Z(n51292) );
  XOR U51180 ( .A(p_input[1581]), .B(p_input[2061]), .Z(n51289) );
  XOR U51181 ( .A(p_input[1582]), .B(n29035), .Z(n51322) );
  XOR U51182 ( .A(p_input[1577]), .B(p_input[2057]), .Z(n51283) );
  XOR U51183 ( .A(n51301), .B(n51299), .Z(n51281) );
  XNOR U51184 ( .A(n51323), .B(n51306), .Z(n51299) );
  XOR U51185 ( .A(p_input[1576]), .B(p_input[2056]), .Z(n51306) );
  XOR U51186 ( .A(n51296), .B(n51305), .Z(n51323) );
  XOR U51187 ( .A(n51324), .B(n51302), .Z(n51305) );
  XOR U51188 ( .A(p_input[1574]), .B(p_input[2054]), .Z(n51302) );
  XOR U51189 ( .A(p_input[1575]), .B(n30404), .Z(n51324) );
  XOR U51190 ( .A(p_input[1570]), .B(p_input[2050]), .Z(n51296) );
  XNOR U51191 ( .A(n51311), .B(n51310), .Z(n51301) );
  XOR U51192 ( .A(n51325), .B(n51307), .Z(n51310) );
  XOR U51193 ( .A(p_input[1571]), .B(p_input[2051]), .Z(n51307) );
  XOR U51194 ( .A(p_input[1572]), .B(n30406), .Z(n51325) );
  XOR U51195 ( .A(p_input[1573]), .B(p_input[2053]), .Z(n51311) );
  XNOR U51196 ( .A(n51326), .B(n51327), .Z(n51207) );
  AND U51197 ( .A(n1937), .B(n51328), .Z(n51327) );
  XNOR U51198 ( .A(n51329), .B(n51330), .Z(n1937) );
  AND U51199 ( .A(n51331), .B(n51332), .Z(n51330) );
  XOR U51200 ( .A(n51221), .B(n51329), .Z(n51332) );
  XNOR U51201 ( .A(n51333), .B(n51329), .Z(n51331) );
  XOR U51202 ( .A(n51334), .B(n51335), .Z(n51329) );
  AND U51203 ( .A(n51336), .B(n51337), .Z(n51335) );
  XOR U51204 ( .A(n51236), .B(n51334), .Z(n51337) );
  XOR U51205 ( .A(n51334), .B(n51237), .Z(n51336) );
  XOR U51206 ( .A(n51338), .B(n51339), .Z(n51334) );
  AND U51207 ( .A(n51340), .B(n51341), .Z(n51339) );
  XOR U51208 ( .A(n51264), .B(n51338), .Z(n51341) );
  XOR U51209 ( .A(n51338), .B(n51265), .Z(n51340) );
  XOR U51210 ( .A(n51342), .B(n51343), .Z(n51338) );
  AND U51211 ( .A(n51344), .B(n51345), .Z(n51343) );
  XOR U51212 ( .A(n51342), .B(n51315), .Z(n51345) );
  XNOR U51213 ( .A(n51346), .B(n51347), .Z(n51167) );
  AND U51214 ( .A(n1941), .B(n51348), .Z(n51347) );
  XNOR U51215 ( .A(n51349), .B(n51350), .Z(n1941) );
  AND U51216 ( .A(n51351), .B(n51352), .Z(n51350) );
  XOR U51217 ( .A(n51349), .B(n51177), .Z(n51352) );
  XNOR U51218 ( .A(n51349), .B(n51137), .Z(n51351) );
  XOR U51219 ( .A(n51353), .B(n51354), .Z(n51349) );
  AND U51220 ( .A(n51355), .B(n51356), .Z(n51354) );
  XOR U51221 ( .A(n51353), .B(n51145), .Z(n51355) );
  XOR U51222 ( .A(n51357), .B(n51358), .Z(n51128) );
  AND U51223 ( .A(n1945), .B(n51348), .Z(n51358) );
  XNOR U51224 ( .A(n51346), .B(n51357), .Z(n51348) );
  XNOR U51225 ( .A(n51359), .B(n51360), .Z(n1945) );
  AND U51226 ( .A(n51361), .B(n51362), .Z(n51360) );
  XNOR U51227 ( .A(n51363), .B(n51359), .Z(n51362) );
  IV U51228 ( .A(n51177), .Z(n51363) );
  XOR U51229 ( .A(n51333), .B(n51364), .Z(n51177) );
  AND U51230 ( .A(n1948), .B(n51365), .Z(n51364) );
  XOR U51231 ( .A(n51220), .B(n51217), .Z(n51365) );
  IV U51232 ( .A(n51333), .Z(n51220) );
  XNOR U51233 ( .A(n51137), .B(n51359), .Z(n51361) );
  XOR U51234 ( .A(n51366), .B(n51367), .Z(n51137) );
  AND U51235 ( .A(n1964), .B(n51368), .Z(n51367) );
  XOR U51236 ( .A(n51353), .B(n51369), .Z(n51359) );
  AND U51237 ( .A(n51370), .B(n51356), .Z(n51369) );
  XNOR U51238 ( .A(n51187), .B(n51353), .Z(n51356) );
  XOR U51239 ( .A(n51237), .B(n51371), .Z(n51187) );
  AND U51240 ( .A(n1948), .B(n51372), .Z(n51371) );
  XOR U51241 ( .A(n51233), .B(n51237), .Z(n51372) );
  XNOR U51242 ( .A(n51373), .B(n51353), .Z(n51370) );
  IV U51243 ( .A(n51145), .Z(n51373) );
  XOR U51244 ( .A(n51374), .B(n51375), .Z(n51145) );
  AND U51245 ( .A(n1964), .B(n51376), .Z(n51375) );
  XOR U51246 ( .A(n51377), .B(n51378), .Z(n51353) );
  AND U51247 ( .A(n51379), .B(n51380), .Z(n51378) );
  XNOR U51248 ( .A(n51197), .B(n51377), .Z(n51380) );
  XOR U51249 ( .A(n51265), .B(n51381), .Z(n51197) );
  AND U51250 ( .A(n1948), .B(n51382), .Z(n51381) );
  XOR U51251 ( .A(n51261), .B(n51265), .Z(n51382) );
  XOR U51252 ( .A(n51377), .B(n51154), .Z(n51379) );
  XOR U51253 ( .A(n51383), .B(n51384), .Z(n51154) );
  AND U51254 ( .A(n1964), .B(n51385), .Z(n51384) );
  XOR U51255 ( .A(n51386), .B(n51387), .Z(n51377) );
  AND U51256 ( .A(n51388), .B(n51389), .Z(n51387) );
  XNOR U51257 ( .A(n51386), .B(n51205), .Z(n51389) );
  XOR U51258 ( .A(n51316), .B(n51390), .Z(n51205) );
  AND U51259 ( .A(n1948), .B(n51391), .Z(n51390) );
  XOR U51260 ( .A(n51312), .B(n51316), .Z(n51391) );
  XNOR U51261 ( .A(n51392), .B(n51386), .Z(n51388) );
  IV U51262 ( .A(n51164), .Z(n51392) );
  XOR U51263 ( .A(n51393), .B(n51394), .Z(n51164) );
  AND U51264 ( .A(n1964), .B(n51395), .Z(n51394) );
  AND U51265 ( .A(n51357), .B(n51346), .Z(n51386) );
  XNOR U51266 ( .A(n51396), .B(n51397), .Z(n51346) );
  AND U51267 ( .A(n1948), .B(n51328), .Z(n51397) );
  XNOR U51268 ( .A(n51326), .B(n51396), .Z(n51328) );
  XNOR U51269 ( .A(n51398), .B(n51399), .Z(n1948) );
  AND U51270 ( .A(n51400), .B(n51401), .Z(n51399) );
  XNOR U51271 ( .A(n51398), .B(n51217), .Z(n51401) );
  IV U51272 ( .A(n51221), .Z(n51217) );
  XOR U51273 ( .A(n51402), .B(n51403), .Z(n51221) );
  AND U51274 ( .A(n1952), .B(n51404), .Z(n51403) );
  XOR U51275 ( .A(n51405), .B(n51402), .Z(n51404) );
  XNOR U51276 ( .A(n51398), .B(n51333), .Z(n51400) );
  XOR U51277 ( .A(n51406), .B(n51407), .Z(n51333) );
  AND U51278 ( .A(n1960), .B(n51368), .Z(n51407) );
  XOR U51279 ( .A(n51366), .B(n51406), .Z(n51368) );
  XOR U51280 ( .A(n51408), .B(n51409), .Z(n51398) );
  AND U51281 ( .A(n51410), .B(n51411), .Z(n51409) );
  XNOR U51282 ( .A(n51408), .B(n51233), .Z(n51411) );
  IV U51283 ( .A(n51236), .Z(n51233) );
  XOR U51284 ( .A(n51412), .B(n51413), .Z(n51236) );
  AND U51285 ( .A(n1952), .B(n51414), .Z(n51413) );
  XOR U51286 ( .A(n51415), .B(n51412), .Z(n51414) );
  XOR U51287 ( .A(n51237), .B(n51408), .Z(n51410) );
  XOR U51288 ( .A(n51416), .B(n51417), .Z(n51237) );
  AND U51289 ( .A(n1960), .B(n51376), .Z(n51417) );
  XOR U51290 ( .A(n51416), .B(n51374), .Z(n51376) );
  XOR U51291 ( .A(n51418), .B(n51419), .Z(n51408) );
  AND U51292 ( .A(n51420), .B(n51421), .Z(n51419) );
  XNOR U51293 ( .A(n51418), .B(n51261), .Z(n51421) );
  IV U51294 ( .A(n51264), .Z(n51261) );
  XOR U51295 ( .A(n51422), .B(n51423), .Z(n51264) );
  AND U51296 ( .A(n1952), .B(n51424), .Z(n51423) );
  XNOR U51297 ( .A(n51425), .B(n51422), .Z(n51424) );
  XOR U51298 ( .A(n51265), .B(n51418), .Z(n51420) );
  XOR U51299 ( .A(n51426), .B(n51427), .Z(n51265) );
  AND U51300 ( .A(n1960), .B(n51385), .Z(n51427) );
  XOR U51301 ( .A(n51426), .B(n51383), .Z(n51385) );
  XOR U51302 ( .A(n51342), .B(n51428), .Z(n51418) );
  AND U51303 ( .A(n51344), .B(n51429), .Z(n51428) );
  XNOR U51304 ( .A(n51342), .B(n51312), .Z(n51429) );
  IV U51305 ( .A(n51315), .Z(n51312) );
  XOR U51306 ( .A(n51430), .B(n51431), .Z(n51315) );
  AND U51307 ( .A(n1952), .B(n51432), .Z(n51431) );
  XOR U51308 ( .A(n51433), .B(n51430), .Z(n51432) );
  XOR U51309 ( .A(n51316), .B(n51342), .Z(n51344) );
  XOR U51310 ( .A(n51434), .B(n51435), .Z(n51316) );
  AND U51311 ( .A(n1960), .B(n51395), .Z(n51435) );
  XOR U51312 ( .A(n51434), .B(n51393), .Z(n51395) );
  AND U51313 ( .A(n51396), .B(n51326), .Z(n51342) );
  XNOR U51314 ( .A(n51436), .B(n51437), .Z(n51326) );
  AND U51315 ( .A(n1952), .B(n51438), .Z(n51437) );
  XNOR U51316 ( .A(n51439), .B(n51436), .Z(n51438) );
  XNOR U51317 ( .A(n51440), .B(n51441), .Z(n1952) );
  AND U51318 ( .A(n51442), .B(n51443), .Z(n51441) );
  XOR U51319 ( .A(n51405), .B(n51440), .Z(n51443) );
  AND U51320 ( .A(n51444), .B(n51445), .Z(n51405) );
  XNOR U51321 ( .A(n51402), .B(n51440), .Z(n51442) );
  XNOR U51322 ( .A(n51446), .B(n51447), .Z(n51402) );
  AND U51323 ( .A(n1956), .B(n51448), .Z(n51447) );
  XNOR U51324 ( .A(n51449), .B(n51450), .Z(n51448) );
  XOR U51325 ( .A(n51451), .B(n51452), .Z(n51440) );
  AND U51326 ( .A(n51453), .B(n51454), .Z(n51452) );
  XNOR U51327 ( .A(n51451), .B(n51444), .Z(n51454) );
  IV U51328 ( .A(n51415), .Z(n51444) );
  XOR U51329 ( .A(n51455), .B(n51456), .Z(n51415) );
  XOR U51330 ( .A(n51457), .B(n51445), .Z(n51456) );
  AND U51331 ( .A(n51425), .B(n51458), .Z(n51445) );
  AND U51332 ( .A(n51459), .B(n51460), .Z(n51457) );
  XOR U51333 ( .A(n51461), .B(n51455), .Z(n51459) );
  XNOR U51334 ( .A(n51412), .B(n51451), .Z(n51453) );
  XNOR U51335 ( .A(n51462), .B(n51463), .Z(n51412) );
  AND U51336 ( .A(n1956), .B(n51464), .Z(n51463) );
  XNOR U51337 ( .A(n51465), .B(n51466), .Z(n51464) );
  XOR U51338 ( .A(n51467), .B(n51468), .Z(n51451) );
  AND U51339 ( .A(n51469), .B(n51470), .Z(n51468) );
  XNOR U51340 ( .A(n51467), .B(n51425), .Z(n51470) );
  XOR U51341 ( .A(n51471), .B(n51460), .Z(n51425) );
  XNOR U51342 ( .A(n51472), .B(n51455), .Z(n51460) );
  XOR U51343 ( .A(n51473), .B(n51474), .Z(n51455) );
  AND U51344 ( .A(n51475), .B(n51476), .Z(n51474) );
  XOR U51345 ( .A(n51477), .B(n51473), .Z(n51475) );
  XNOR U51346 ( .A(n51478), .B(n51479), .Z(n51472) );
  AND U51347 ( .A(n51480), .B(n51481), .Z(n51479) );
  XOR U51348 ( .A(n51478), .B(n51482), .Z(n51480) );
  XNOR U51349 ( .A(n51461), .B(n51458), .Z(n51471) );
  AND U51350 ( .A(n51483), .B(n51484), .Z(n51458) );
  XOR U51351 ( .A(n51485), .B(n51486), .Z(n51461) );
  AND U51352 ( .A(n51487), .B(n51488), .Z(n51486) );
  XOR U51353 ( .A(n51485), .B(n51489), .Z(n51487) );
  XNOR U51354 ( .A(n51422), .B(n51467), .Z(n51469) );
  XNOR U51355 ( .A(n51490), .B(n51491), .Z(n51422) );
  AND U51356 ( .A(n1956), .B(n51492), .Z(n51491) );
  XNOR U51357 ( .A(n51493), .B(n51494), .Z(n51492) );
  XOR U51358 ( .A(n51495), .B(n51496), .Z(n51467) );
  AND U51359 ( .A(n51497), .B(n51498), .Z(n51496) );
  XNOR U51360 ( .A(n51495), .B(n51483), .Z(n51498) );
  IV U51361 ( .A(n51433), .Z(n51483) );
  XNOR U51362 ( .A(n51499), .B(n51476), .Z(n51433) );
  XNOR U51363 ( .A(n51500), .B(n51482), .Z(n51476) );
  XNOR U51364 ( .A(n51501), .B(n51502), .Z(n51482) );
  NOR U51365 ( .A(n51503), .B(n51504), .Z(n51502) );
  XOR U51366 ( .A(n51501), .B(n51505), .Z(n51503) );
  XNOR U51367 ( .A(n51481), .B(n51473), .Z(n51500) );
  XOR U51368 ( .A(n51506), .B(n51507), .Z(n51473) );
  AND U51369 ( .A(n51508), .B(n51509), .Z(n51507) );
  XOR U51370 ( .A(n51506), .B(n51510), .Z(n51508) );
  XNOR U51371 ( .A(n51511), .B(n51478), .Z(n51481) );
  XOR U51372 ( .A(n51512), .B(n51513), .Z(n51478) );
  AND U51373 ( .A(n51514), .B(n51515), .Z(n51513) );
  XNOR U51374 ( .A(n51516), .B(n51517), .Z(n51514) );
  IV U51375 ( .A(n51512), .Z(n51516) );
  XNOR U51376 ( .A(n51518), .B(n51519), .Z(n51511) );
  NOR U51377 ( .A(n51520), .B(n51521), .Z(n51519) );
  XNOR U51378 ( .A(n51518), .B(n51522), .Z(n51520) );
  XNOR U51379 ( .A(n51477), .B(n51484), .Z(n51499) );
  NOR U51380 ( .A(n51439), .B(n51523), .Z(n51484) );
  XOR U51381 ( .A(n51489), .B(n51488), .Z(n51477) );
  XNOR U51382 ( .A(n51524), .B(n51485), .Z(n51488) );
  XOR U51383 ( .A(n51525), .B(n51526), .Z(n51485) );
  AND U51384 ( .A(n51527), .B(n51528), .Z(n51526) );
  XNOR U51385 ( .A(n51529), .B(n51530), .Z(n51527) );
  IV U51386 ( .A(n51525), .Z(n51529) );
  XNOR U51387 ( .A(n51531), .B(n51532), .Z(n51524) );
  NOR U51388 ( .A(n51533), .B(n51534), .Z(n51532) );
  XNOR U51389 ( .A(n51531), .B(n51535), .Z(n51533) );
  XOR U51390 ( .A(n51536), .B(n51537), .Z(n51489) );
  NOR U51391 ( .A(n51538), .B(n51539), .Z(n51537) );
  XNOR U51392 ( .A(n51536), .B(n51540), .Z(n51538) );
  XNOR U51393 ( .A(n51430), .B(n51495), .Z(n51497) );
  XNOR U51394 ( .A(n51541), .B(n51542), .Z(n51430) );
  AND U51395 ( .A(n1956), .B(n51543), .Z(n51542) );
  XNOR U51396 ( .A(n51544), .B(n51545), .Z(n51543) );
  AND U51397 ( .A(n51436), .B(n51439), .Z(n51495) );
  XOR U51398 ( .A(n51546), .B(n51523), .Z(n51439) );
  XNOR U51399 ( .A(p_input[1584]), .B(p_input[2048]), .Z(n51523) );
  XNOR U51400 ( .A(n51510), .B(n51509), .Z(n51546) );
  XNOR U51401 ( .A(n51547), .B(n51517), .Z(n51509) );
  XNOR U51402 ( .A(n51505), .B(n51504), .Z(n51517) );
  XNOR U51403 ( .A(n51548), .B(n51501), .Z(n51504) );
  XNOR U51404 ( .A(p_input[1594]), .B(p_input[2058]), .Z(n51501) );
  XOR U51405 ( .A(p_input[1595]), .B(n29030), .Z(n51548) );
  XOR U51406 ( .A(p_input[1596]), .B(p_input[2060]), .Z(n51505) );
  XOR U51407 ( .A(n51515), .B(n51549), .Z(n51547) );
  IV U51408 ( .A(n51506), .Z(n51549) );
  XOR U51409 ( .A(p_input[1585]), .B(p_input[2049]), .Z(n51506) );
  XNOR U51410 ( .A(n51550), .B(n51522), .Z(n51515) );
  XNOR U51411 ( .A(p_input[1599]), .B(n29033), .Z(n51522) );
  XOR U51412 ( .A(n51512), .B(n51521), .Z(n51550) );
  XOR U51413 ( .A(n51551), .B(n51518), .Z(n51521) );
  XOR U51414 ( .A(p_input[1597]), .B(p_input[2061]), .Z(n51518) );
  XOR U51415 ( .A(p_input[1598]), .B(n29035), .Z(n51551) );
  XOR U51416 ( .A(p_input[1593]), .B(p_input[2057]), .Z(n51512) );
  XOR U51417 ( .A(n51530), .B(n51528), .Z(n51510) );
  XNOR U51418 ( .A(n51552), .B(n51535), .Z(n51528) );
  XOR U51419 ( .A(p_input[1592]), .B(p_input[2056]), .Z(n51535) );
  XOR U51420 ( .A(n51525), .B(n51534), .Z(n51552) );
  XOR U51421 ( .A(n51553), .B(n51531), .Z(n51534) );
  XOR U51422 ( .A(p_input[1590]), .B(p_input[2054]), .Z(n51531) );
  XOR U51423 ( .A(p_input[1591]), .B(n30404), .Z(n51553) );
  XOR U51424 ( .A(p_input[1586]), .B(p_input[2050]), .Z(n51525) );
  XNOR U51425 ( .A(n51540), .B(n51539), .Z(n51530) );
  XOR U51426 ( .A(n51554), .B(n51536), .Z(n51539) );
  XOR U51427 ( .A(p_input[1587]), .B(p_input[2051]), .Z(n51536) );
  XOR U51428 ( .A(p_input[1588]), .B(n30406), .Z(n51554) );
  XOR U51429 ( .A(p_input[1589]), .B(p_input[2053]), .Z(n51540) );
  XNOR U51430 ( .A(n51555), .B(n51556), .Z(n51436) );
  AND U51431 ( .A(n1956), .B(n51557), .Z(n51556) );
  XNOR U51432 ( .A(n51558), .B(n51559), .Z(n1956) );
  AND U51433 ( .A(n51560), .B(n51561), .Z(n51559) );
  XOR U51434 ( .A(n51450), .B(n51558), .Z(n51561) );
  XNOR U51435 ( .A(n51562), .B(n51558), .Z(n51560) );
  XOR U51436 ( .A(n51563), .B(n51564), .Z(n51558) );
  AND U51437 ( .A(n51565), .B(n51566), .Z(n51564) );
  XOR U51438 ( .A(n51465), .B(n51563), .Z(n51566) );
  XOR U51439 ( .A(n51563), .B(n51466), .Z(n51565) );
  XOR U51440 ( .A(n51567), .B(n51568), .Z(n51563) );
  AND U51441 ( .A(n51569), .B(n51570), .Z(n51568) );
  XOR U51442 ( .A(n51493), .B(n51567), .Z(n51570) );
  XOR U51443 ( .A(n51567), .B(n51494), .Z(n51569) );
  XOR U51444 ( .A(n51571), .B(n51572), .Z(n51567) );
  AND U51445 ( .A(n51573), .B(n51574), .Z(n51572) );
  XOR U51446 ( .A(n51571), .B(n51544), .Z(n51574) );
  XNOR U51447 ( .A(n51575), .B(n51576), .Z(n51396) );
  AND U51448 ( .A(n1960), .B(n51577), .Z(n51576) );
  XNOR U51449 ( .A(n51578), .B(n51579), .Z(n1960) );
  AND U51450 ( .A(n51580), .B(n51581), .Z(n51579) );
  XOR U51451 ( .A(n51578), .B(n51406), .Z(n51581) );
  XNOR U51452 ( .A(n51578), .B(n51366), .Z(n51580) );
  XOR U51453 ( .A(n51582), .B(n51583), .Z(n51578) );
  AND U51454 ( .A(n51584), .B(n51585), .Z(n51583) );
  XOR U51455 ( .A(n51582), .B(n51374), .Z(n51584) );
  XOR U51456 ( .A(n51586), .B(n51587), .Z(n51357) );
  AND U51457 ( .A(n1964), .B(n51577), .Z(n51587) );
  XNOR U51458 ( .A(n51575), .B(n51586), .Z(n51577) );
  XNOR U51459 ( .A(n51588), .B(n51589), .Z(n1964) );
  AND U51460 ( .A(n51590), .B(n51591), .Z(n51589) );
  XNOR U51461 ( .A(n51592), .B(n51588), .Z(n51591) );
  IV U51462 ( .A(n51406), .Z(n51592) );
  XOR U51463 ( .A(n51562), .B(n51593), .Z(n51406) );
  AND U51464 ( .A(n1967), .B(n51594), .Z(n51593) );
  XOR U51465 ( .A(n51449), .B(n51446), .Z(n51594) );
  IV U51466 ( .A(n51562), .Z(n51449) );
  XNOR U51467 ( .A(n51366), .B(n51588), .Z(n51590) );
  XOR U51468 ( .A(n51595), .B(n51596), .Z(n51366) );
  AND U51469 ( .A(n1983), .B(n51597), .Z(n51596) );
  XOR U51470 ( .A(n51582), .B(n51598), .Z(n51588) );
  AND U51471 ( .A(n51599), .B(n51585), .Z(n51598) );
  XNOR U51472 ( .A(n51416), .B(n51582), .Z(n51585) );
  XOR U51473 ( .A(n51466), .B(n51600), .Z(n51416) );
  AND U51474 ( .A(n1967), .B(n51601), .Z(n51600) );
  XOR U51475 ( .A(n51462), .B(n51466), .Z(n51601) );
  XNOR U51476 ( .A(n51602), .B(n51582), .Z(n51599) );
  IV U51477 ( .A(n51374), .Z(n51602) );
  XOR U51478 ( .A(n51603), .B(n51604), .Z(n51374) );
  AND U51479 ( .A(n1983), .B(n51605), .Z(n51604) );
  XOR U51480 ( .A(n51606), .B(n51607), .Z(n51582) );
  AND U51481 ( .A(n51608), .B(n51609), .Z(n51607) );
  XNOR U51482 ( .A(n51426), .B(n51606), .Z(n51609) );
  XOR U51483 ( .A(n51494), .B(n51610), .Z(n51426) );
  AND U51484 ( .A(n1967), .B(n51611), .Z(n51610) );
  XOR U51485 ( .A(n51490), .B(n51494), .Z(n51611) );
  XOR U51486 ( .A(n51606), .B(n51383), .Z(n51608) );
  XOR U51487 ( .A(n51612), .B(n51613), .Z(n51383) );
  AND U51488 ( .A(n1983), .B(n51614), .Z(n51613) );
  XOR U51489 ( .A(n51615), .B(n51616), .Z(n51606) );
  AND U51490 ( .A(n51617), .B(n51618), .Z(n51616) );
  XNOR U51491 ( .A(n51615), .B(n51434), .Z(n51618) );
  XOR U51492 ( .A(n51545), .B(n51619), .Z(n51434) );
  AND U51493 ( .A(n1967), .B(n51620), .Z(n51619) );
  XOR U51494 ( .A(n51541), .B(n51545), .Z(n51620) );
  XNOR U51495 ( .A(n51621), .B(n51615), .Z(n51617) );
  IV U51496 ( .A(n51393), .Z(n51621) );
  XOR U51497 ( .A(n51622), .B(n51623), .Z(n51393) );
  AND U51498 ( .A(n1983), .B(n51624), .Z(n51623) );
  AND U51499 ( .A(n51586), .B(n51575), .Z(n51615) );
  XNOR U51500 ( .A(n51625), .B(n51626), .Z(n51575) );
  AND U51501 ( .A(n1967), .B(n51557), .Z(n51626) );
  XNOR U51502 ( .A(n51555), .B(n51625), .Z(n51557) );
  XNOR U51503 ( .A(n51627), .B(n51628), .Z(n1967) );
  AND U51504 ( .A(n51629), .B(n51630), .Z(n51628) );
  XNOR U51505 ( .A(n51627), .B(n51446), .Z(n51630) );
  IV U51506 ( .A(n51450), .Z(n51446) );
  XOR U51507 ( .A(n51631), .B(n51632), .Z(n51450) );
  AND U51508 ( .A(n1971), .B(n51633), .Z(n51632) );
  XOR U51509 ( .A(n51634), .B(n51631), .Z(n51633) );
  XNOR U51510 ( .A(n51627), .B(n51562), .Z(n51629) );
  XOR U51511 ( .A(n51635), .B(n51636), .Z(n51562) );
  AND U51512 ( .A(n1979), .B(n51597), .Z(n51636) );
  XOR U51513 ( .A(n51595), .B(n51635), .Z(n51597) );
  XOR U51514 ( .A(n51637), .B(n51638), .Z(n51627) );
  AND U51515 ( .A(n51639), .B(n51640), .Z(n51638) );
  XNOR U51516 ( .A(n51637), .B(n51462), .Z(n51640) );
  IV U51517 ( .A(n51465), .Z(n51462) );
  XOR U51518 ( .A(n51641), .B(n51642), .Z(n51465) );
  AND U51519 ( .A(n1971), .B(n51643), .Z(n51642) );
  XOR U51520 ( .A(n51644), .B(n51641), .Z(n51643) );
  XOR U51521 ( .A(n51466), .B(n51637), .Z(n51639) );
  XOR U51522 ( .A(n51645), .B(n51646), .Z(n51466) );
  AND U51523 ( .A(n1979), .B(n51605), .Z(n51646) );
  XOR U51524 ( .A(n51645), .B(n51603), .Z(n51605) );
  XOR U51525 ( .A(n51647), .B(n51648), .Z(n51637) );
  AND U51526 ( .A(n51649), .B(n51650), .Z(n51648) );
  XNOR U51527 ( .A(n51647), .B(n51490), .Z(n51650) );
  IV U51528 ( .A(n51493), .Z(n51490) );
  XOR U51529 ( .A(n51651), .B(n51652), .Z(n51493) );
  AND U51530 ( .A(n1971), .B(n51653), .Z(n51652) );
  XNOR U51531 ( .A(n51654), .B(n51651), .Z(n51653) );
  XOR U51532 ( .A(n51494), .B(n51647), .Z(n51649) );
  XOR U51533 ( .A(n51655), .B(n51656), .Z(n51494) );
  AND U51534 ( .A(n1979), .B(n51614), .Z(n51656) );
  XOR U51535 ( .A(n51655), .B(n51612), .Z(n51614) );
  XOR U51536 ( .A(n51571), .B(n51657), .Z(n51647) );
  AND U51537 ( .A(n51573), .B(n51658), .Z(n51657) );
  XNOR U51538 ( .A(n51571), .B(n51541), .Z(n51658) );
  IV U51539 ( .A(n51544), .Z(n51541) );
  XOR U51540 ( .A(n51659), .B(n51660), .Z(n51544) );
  AND U51541 ( .A(n1971), .B(n51661), .Z(n51660) );
  XOR U51542 ( .A(n51662), .B(n51659), .Z(n51661) );
  XOR U51543 ( .A(n51545), .B(n51571), .Z(n51573) );
  XOR U51544 ( .A(n51663), .B(n51664), .Z(n51545) );
  AND U51545 ( .A(n1979), .B(n51624), .Z(n51664) );
  XOR U51546 ( .A(n51663), .B(n51622), .Z(n51624) );
  AND U51547 ( .A(n51625), .B(n51555), .Z(n51571) );
  XNOR U51548 ( .A(n51665), .B(n51666), .Z(n51555) );
  AND U51549 ( .A(n1971), .B(n51667), .Z(n51666) );
  XNOR U51550 ( .A(n51668), .B(n51665), .Z(n51667) );
  XNOR U51551 ( .A(n51669), .B(n51670), .Z(n1971) );
  AND U51552 ( .A(n51671), .B(n51672), .Z(n51670) );
  XOR U51553 ( .A(n51634), .B(n51669), .Z(n51672) );
  AND U51554 ( .A(n51673), .B(n51674), .Z(n51634) );
  XNOR U51555 ( .A(n51631), .B(n51669), .Z(n51671) );
  XNOR U51556 ( .A(n51675), .B(n51676), .Z(n51631) );
  AND U51557 ( .A(n1975), .B(n51677), .Z(n51676) );
  XNOR U51558 ( .A(n51678), .B(n51679), .Z(n51677) );
  XOR U51559 ( .A(n51680), .B(n51681), .Z(n51669) );
  AND U51560 ( .A(n51682), .B(n51683), .Z(n51681) );
  XNOR U51561 ( .A(n51680), .B(n51673), .Z(n51683) );
  IV U51562 ( .A(n51644), .Z(n51673) );
  XOR U51563 ( .A(n51684), .B(n51685), .Z(n51644) );
  XOR U51564 ( .A(n51686), .B(n51674), .Z(n51685) );
  AND U51565 ( .A(n51654), .B(n51687), .Z(n51674) );
  AND U51566 ( .A(n51688), .B(n51689), .Z(n51686) );
  XOR U51567 ( .A(n51690), .B(n51684), .Z(n51688) );
  XNOR U51568 ( .A(n51641), .B(n51680), .Z(n51682) );
  XNOR U51569 ( .A(n51691), .B(n51692), .Z(n51641) );
  AND U51570 ( .A(n1975), .B(n51693), .Z(n51692) );
  XNOR U51571 ( .A(n51694), .B(n51695), .Z(n51693) );
  XOR U51572 ( .A(n51696), .B(n51697), .Z(n51680) );
  AND U51573 ( .A(n51698), .B(n51699), .Z(n51697) );
  XNOR U51574 ( .A(n51696), .B(n51654), .Z(n51699) );
  XOR U51575 ( .A(n51700), .B(n51689), .Z(n51654) );
  XNOR U51576 ( .A(n51701), .B(n51684), .Z(n51689) );
  XOR U51577 ( .A(n51702), .B(n51703), .Z(n51684) );
  AND U51578 ( .A(n51704), .B(n51705), .Z(n51703) );
  XOR U51579 ( .A(n51706), .B(n51702), .Z(n51704) );
  XNOR U51580 ( .A(n51707), .B(n51708), .Z(n51701) );
  AND U51581 ( .A(n51709), .B(n51710), .Z(n51708) );
  XOR U51582 ( .A(n51707), .B(n51711), .Z(n51709) );
  XNOR U51583 ( .A(n51690), .B(n51687), .Z(n51700) );
  AND U51584 ( .A(n51712), .B(n51713), .Z(n51687) );
  XOR U51585 ( .A(n51714), .B(n51715), .Z(n51690) );
  AND U51586 ( .A(n51716), .B(n51717), .Z(n51715) );
  XOR U51587 ( .A(n51714), .B(n51718), .Z(n51716) );
  XNOR U51588 ( .A(n51651), .B(n51696), .Z(n51698) );
  XNOR U51589 ( .A(n51719), .B(n51720), .Z(n51651) );
  AND U51590 ( .A(n1975), .B(n51721), .Z(n51720) );
  XNOR U51591 ( .A(n51722), .B(n51723), .Z(n51721) );
  XOR U51592 ( .A(n51724), .B(n51725), .Z(n51696) );
  AND U51593 ( .A(n51726), .B(n51727), .Z(n51725) );
  XNOR U51594 ( .A(n51724), .B(n51712), .Z(n51727) );
  IV U51595 ( .A(n51662), .Z(n51712) );
  XNOR U51596 ( .A(n51728), .B(n51705), .Z(n51662) );
  XNOR U51597 ( .A(n51729), .B(n51711), .Z(n51705) );
  XNOR U51598 ( .A(n51730), .B(n51731), .Z(n51711) );
  NOR U51599 ( .A(n51732), .B(n51733), .Z(n51731) );
  XOR U51600 ( .A(n51730), .B(n51734), .Z(n51732) );
  XNOR U51601 ( .A(n51710), .B(n51702), .Z(n51729) );
  XOR U51602 ( .A(n51735), .B(n51736), .Z(n51702) );
  AND U51603 ( .A(n51737), .B(n51738), .Z(n51736) );
  XOR U51604 ( .A(n51735), .B(n51739), .Z(n51737) );
  XNOR U51605 ( .A(n51740), .B(n51707), .Z(n51710) );
  XOR U51606 ( .A(n51741), .B(n51742), .Z(n51707) );
  AND U51607 ( .A(n51743), .B(n51744), .Z(n51742) );
  XNOR U51608 ( .A(n51745), .B(n51746), .Z(n51743) );
  IV U51609 ( .A(n51741), .Z(n51745) );
  XNOR U51610 ( .A(n51747), .B(n51748), .Z(n51740) );
  NOR U51611 ( .A(n51749), .B(n51750), .Z(n51748) );
  XNOR U51612 ( .A(n51747), .B(n51751), .Z(n51749) );
  XNOR U51613 ( .A(n51706), .B(n51713), .Z(n51728) );
  NOR U51614 ( .A(n51668), .B(n51752), .Z(n51713) );
  XOR U51615 ( .A(n51718), .B(n51717), .Z(n51706) );
  XNOR U51616 ( .A(n51753), .B(n51714), .Z(n51717) );
  XOR U51617 ( .A(n51754), .B(n51755), .Z(n51714) );
  AND U51618 ( .A(n51756), .B(n51757), .Z(n51755) );
  XNOR U51619 ( .A(n51758), .B(n51759), .Z(n51756) );
  IV U51620 ( .A(n51754), .Z(n51758) );
  XNOR U51621 ( .A(n51760), .B(n51761), .Z(n51753) );
  NOR U51622 ( .A(n51762), .B(n51763), .Z(n51761) );
  XNOR U51623 ( .A(n51760), .B(n51764), .Z(n51762) );
  XOR U51624 ( .A(n51765), .B(n51766), .Z(n51718) );
  NOR U51625 ( .A(n51767), .B(n51768), .Z(n51766) );
  XNOR U51626 ( .A(n51765), .B(n51769), .Z(n51767) );
  XNOR U51627 ( .A(n51659), .B(n51724), .Z(n51726) );
  XNOR U51628 ( .A(n51770), .B(n51771), .Z(n51659) );
  AND U51629 ( .A(n1975), .B(n51772), .Z(n51771) );
  XNOR U51630 ( .A(n51773), .B(n51774), .Z(n51772) );
  AND U51631 ( .A(n51665), .B(n51668), .Z(n51724) );
  XOR U51632 ( .A(n51775), .B(n51752), .Z(n51668) );
  XNOR U51633 ( .A(p_input[1600]), .B(p_input[2048]), .Z(n51752) );
  XNOR U51634 ( .A(n51739), .B(n51738), .Z(n51775) );
  XNOR U51635 ( .A(n51776), .B(n51746), .Z(n51738) );
  XNOR U51636 ( .A(n51734), .B(n51733), .Z(n51746) );
  XNOR U51637 ( .A(n51777), .B(n51730), .Z(n51733) );
  XNOR U51638 ( .A(p_input[1610]), .B(p_input[2058]), .Z(n51730) );
  XOR U51639 ( .A(p_input[1611]), .B(n29030), .Z(n51777) );
  XOR U51640 ( .A(p_input[1612]), .B(p_input[2060]), .Z(n51734) );
  XOR U51641 ( .A(n51744), .B(n51778), .Z(n51776) );
  IV U51642 ( .A(n51735), .Z(n51778) );
  XOR U51643 ( .A(p_input[1601]), .B(p_input[2049]), .Z(n51735) );
  XNOR U51644 ( .A(n51779), .B(n51751), .Z(n51744) );
  XNOR U51645 ( .A(p_input[1615]), .B(n29033), .Z(n51751) );
  XOR U51646 ( .A(n51741), .B(n51750), .Z(n51779) );
  XOR U51647 ( .A(n51780), .B(n51747), .Z(n51750) );
  XOR U51648 ( .A(p_input[1613]), .B(p_input[2061]), .Z(n51747) );
  XOR U51649 ( .A(p_input[1614]), .B(n29035), .Z(n51780) );
  XOR U51650 ( .A(p_input[1609]), .B(p_input[2057]), .Z(n51741) );
  XOR U51651 ( .A(n51759), .B(n51757), .Z(n51739) );
  XNOR U51652 ( .A(n51781), .B(n51764), .Z(n51757) );
  XOR U51653 ( .A(p_input[1608]), .B(p_input[2056]), .Z(n51764) );
  XOR U51654 ( .A(n51754), .B(n51763), .Z(n51781) );
  XOR U51655 ( .A(n51782), .B(n51760), .Z(n51763) );
  XOR U51656 ( .A(p_input[1606]), .B(p_input[2054]), .Z(n51760) );
  XOR U51657 ( .A(p_input[1607]), .B(n30404), .Z(n51782) );
  XOR U51658 ( .A(p_input[1602]), .B(p_input[2050]), .Z(n51754) );
  XNOR U51659 ( .A(n51769), .B(n51768), .Z(n51759) );
  XOR U51660 ( .A(n51783), .B(n51765), .Z(n51768) );
  XOR U51661 ( .A(p_input[1603]), .B(p_input[2051]), .Z(n51765) );
  XOR U51662 ( .A(p_input[1604]), .B(n30406), .Z(n51783) );
  XOR U51663 ( .A(p_input[1605]), .B(p_input[2053]), .Z(n51769) );
  XNOR U51664 ( .A(n51784), .B(n51785), .Z(n51665) );
  AND U51665 ( .A(n1975), .B(n51786), .Z(n51785) );
  XNOR U51666 ( .A(n51787), .B(n51788), .Z(n1975) );
  AND U51667 ( .A(n51789), .B(n51790), .Z(n51788) );
  XOR U51668 ( .A(n51679), .B(n51787), .Z(n51790) );
  XNOR U51669 ( .A(n51791), .B(n51787), .Z(n51789) );
  XOR U51670 ( .A(n51792), .B(n51793), .Z(n51787) );
  AND U51671 ( .A(n51794), .B(n51795), .Z(n51793) );
  XOR U51672 ( .A(n51694), .B(n51792), .Z(n51795) );
  XOR U51673 ( .A(n51792), .B(n51695), .Z(n51794) );
  XOR U51674 ( .A(n51796), .B(n51797), .Z(n51792) );
  AND U51675 ( .A(n51798), .B(n51799), .Z(n51797) );
  XOR U51676 ( .A(n51722), .B(n51796), .Z(n51799) );
  XOR U51677 ( .A(n51796), .B(n51723), .Z(n51798) );
  XOR U51678 ( .A(n51800), .B(n51801), .Z(n51796) );
  AND U51679 ( .A(n51802), .B(n51803), .Z(n51801) );
  XOR U51680 ( .A(n51800), .B(n51773), .Z(n51803) );
  XNOR U51681 ( .A(n51804), .B(n51805), .Z(n51625) );
  AND U51682 ( .A(n1979), .B(n51806), .Z(n51805) );
  XNOR U51683 ( .A(n51807), .B(n51808), .Z(n1979) );
  AND U51684 ( .A(n51809), .B(n51810), .Z(n51808) );
  XOR U51685 ( .A(n51807), .B(n51635), .Z(n51810) );
  XNOR U51686 ( .A(n51807), .B(n51595), .Z(n51809) );
  XOR U51687 ( .A(n51811), .B(n51812), .Z(n51807) );
  AND U51688 ( .A(n51813), .B(n51814), .Z(n51812) );
  XOR U51689 ( .A(n51811), .B(n51603), .Z(n51813) );
  XOR U51690 ( .A(n51815), .B(n51816), .Z(n51586) );
  AND U51691 ( .A(n1983), .B(n51806), .Z(n51816) );
  XNOR U51692 ( .A(n51804), .B(n51815), .Z(n51806) );
  XNOR U51693 ( .A(n51817), .B(n51818), .Z(n1983) );
  AND U51694 ( .A(n51819), .B(n51820), .Z(n51818) );
  XNOR U51695 ( .A(n51821), .B(n51817), .Z(n51820) );
  IV U51696 ( .A(n51635), .Z(n51821) );
  XOR U51697 ( .A(n51791), .B(n51822), .Z(n51635) );
  AND U51698 ( .A(n1986), .B(n51823), .Z(n51822) );
  XOR U51699 ( .A(n51678), .B(n51675), .Z(n51823) );
  IV U51700 ( .A(n51791), .Z(n51678) );
  XNOR U51701 ( .A(n51595), .B(n51817), .Z(n51819) );
  XOR U51702 ( .A(n51824), .B(n51825), .Z(n51595) );
  AND U51703 ( .A(n2002), .B(n51826), .Z(n51825) );
  XOR U51704 ( .A(n51811), .B(n51827), .Z(n51817) );
  AND U51705 ( .A(n51828), .B(n51814), .Z(n51827) );
  XNOR U51706 ( .A(n51645), .B(n51811), .Z(n51814) );
  XOR U51707 ( .A(n51695), .B(n51829), .Z(n51645) );
  AND U51708 ( .A(n1986), .B(n51830), .Z(n51829) );
  XOR U51709 ( .A(n51691), .B(n51695), .Z(n51830) );
  XNOR U51710 ( .A(n51831), .B(n51811), .Z(n51828) );
  IV U51711 ( .A(n51603), .Z(n51831) );
  XOR U51712 ( .A(n51832), .B(n51833), .Z(n51603) );
  AND U51713 ( .A(n2002), .B(n51834), .Z(n51833) );
  XOR U51714 ( .A(n51835), .B(n51836), .Z(n51811) );
  AND U51715 ( .A(n51837), .B(n51838), .Z(n51836) );
  XNOR U51716 ( .A(n51655), .B(n51835), .Z(n51838) );
  XOR U51717 ( .A(n51723), .B(n51839), .Z(n51655) );
  AND U51718 ( .A(n1986), .B(n51840), .Z(n51839) );
  XOR U51719 ( .A(n51719), .B(n51723), .Z(n51840) );
  XOR U51720 ( .A(n51835), .B(n51612), .Z(n51837) );
  XOR U51721 ( .A(n51841), .B(n51842), .Z(n51612) );
  AND U51722 ( .A(n2002), .B(n51843), .Z(n51842) );
  XOR U51723 ( .A(n51844), .B(n51845), .Z(n51835) );
  AND U51724 ( .A(n51846), .B(n51847), .Z(n51845) );
  XNOR U51725 ( .A(n51844), .B(n51663), .Z(n51847) );
  XOR U51726 ( .A(n51774), .B(n51848), .Z(n51663) );
  AND U51727 ( .A(n1986), .B(n51849), .Z(n51848) );
  XOR U51728 ( .A(n51770), .B(n51774), .Z(n51849) );
  XNOR U51729 ( .A(n51850), .B(n51844), .Z(n51846) );
  IV U51730 ( .A(n51622), .Z(n51850) );
  XOR U51731 ( .A(n51851), .B(n51852), .Z(n51622) );
  AND U51732 ( .A(n2002), .B(n51853), .Z(n51852) );
  AND U51733 ( .A(n51815), .B(n51804), .Z(n51844) );
  XNOR U51734 ( .A(n51854), .B(n51855), .Z(n51804) );
  AND U51735 ( .A(n1986), .B(n51786), .Z(n51855) );
  XNOR U51736 ( .A(n51784), .B(n51854), .Z(n51786) );
  XNOR U51737 ( .A(n51856), .B(n51857), .Z(n1986) );
  AND U51738 ( .A(n51858), .B(n51859), .Z(n51857) );
  XNOR U51739 ( .A(n51856), .B(n51675), .Z(n51859) );
  IV U51740 ( .A(n51679), .Z(n51675) );
  XOR U51741 ( .A(n51860), .B(n51861), .Z(n51679) );
  AND U51742 ( .A(n1990), .B(n51862), .Z(n51861) );
  XOR U51743 ( .A(n51863), .B(n51860), .Z(n51862) );
  XNOR U51744 ( .A(n51856), .B(n51791), .Z(n51858) );
  XOR U51745 ( .A(n51864), .B(n51865), .Z(n51791) );
  AND U51746 ( .A(n1998), .B(n51826), .Z(n51865) );
  XOR U51747 ( .A(n51824), .B(n51864), .Z(n51826) );
  XOR U51748 ( .A(n51866), .B(n51867), .Z(n51856) );
  AND U51749 ( .A(n51868), .B(n51869), .Z(n51867) );
  XNOR U51750 ( .A(n51866), .B(n51691), .Z(n51869) );
  IV U51751 ( .A(n51694), .Z(n51691) );
  XOR U51752 ( .A(n51870), .B(n51871), .Z(n51694) );
  AND U51753 ( .A(n1990), .B(n51872), .Z(n51871) );
  XOR U51754 ( .A(n51873), .B(n51870), .Z(n51872) );
  XOR U51755 ( .A(n51695), .B(n51866), .Z(n51868) );
  XOR U51756 ( .A(n51874), .B(n51875), .Z(n51695) );
  AND U51757 ( .A(n1998), .B(n51834), .Z(n51875) );
  XOR U51758 ( .A(n51874), .B(n51832), .Z(n51834) );
  XOR U51759 ( .A(n51876), .B(n51877), .Z(n51866) );
  AND U51760 ( .A(n51878), .B(n51879), .Z(n51877) );
  XNOR U51761 ( .A(n51876), .B(n51719), .Z(n51879) );
  IV U51762 ( .A(n51722), .Z(n51719) );
  XOR U51763 ( .A(n51880), .B(n51881), .Z(n51722) );
  AND U51764 ( .A(n1990), .B(n51882), .Z(n51881) );
  XNOR U51765 ( .A(n51883), .B(n51880), .Z(n51882) );
  XOR U51766 ( .A(n51723), .B(n51876), .Z(n51878) );
  XOR U51767 ( .A(n51884), .B(n51885), .Z(n51723) );
  AND U51768 ( .A(n1998), .B(n51843), .Z(n51885) );
  XOR U51769 ( .A(n51884), .B(n51841), .Z(n51843) );
  XOR U51770 ( .A(n51800), .B(n51886), .Z(n51876) );
  AND U51771 ( .A(n51802), .B(n51887), .Z(n51886) );
  XNOR U51772 ( .A(n51800), .B(n51770), .Z(n51887) );
  IV U51773 ( .A(n51773), .Z(n51770) );
  XOR U51774 ( .A(n51888), .B(n51889), .Z(n51773) );
  AND U51775 ( .A(n1990), .B(n51890), .Z(n51889) );
  XOR U51776 ( .A(n51891), .B(n51888), .Z(n51890) );
  XOR U51777 ( .A(n51774), .B(n51800), .Z(n51802) );
  XOR U51778 ( .A(n51892), .B(n51893), .Z(n51774) );
  AND U51779 ( .A(n1998), .B(n51853), .Z(n51893) );
  XOR U51780 ( .A(n51892), .B(n51851), .Z(n51853) );
  AND U51781 ( .A(n51854), .B(n51784), .Z(n51800) );
  XNOR U51782 ( .A(n51894), .B(n51895), .Z(n51784) );
  AND U51783 ( .A(n1990), .B(n51896), .Z(n51895) );
  XNOR U51784 ( .A(n51897), .B(n51894), .Z(n51896) );
  XNOR U51785 ( .A(n51898), .B(n51899), .Z(n1990) );
  AND U51786 ( .A(n51900), .B(n51901), .Z(n51899) );
  XOR U51787 ( .A(n51863), .B(n51898), .Z(n51901) );
  AND U51788 ( .A(n51902), .B(n51903), .Z(n51863) );
  XNOR U51789 ( .A(n51860), .B(n51898), .Z(n51900) );
  XNOR U51790 ( .A(n51904), .B(n51905), .Z(n51860) );
  AND U51791 ( .A(n1994), .B(n51906), .Z(n51905) );
  XNOR U51792 ( .A(n51907), .B(n51908), .Z(n51906) );
  XOR U51793 ( .A(n51909), .B(n51910), .Z(n51898) );
  AND U51794 ( .A(n51911), .B(n51912), .Z(n51910) );
  XNOR U51795 ( .A(n51909), .B(n51902), .Z(n51912) );
  IV U51796 ( .A(n51873), .Z(n51902) );
  XOR U51797 ( .A(n51913), .B(n51914), .Z(n51873) );
  XOR U51798 ( .A(n51915), .B(n51903), .Z(n51914) );
  AND U51799 ( .A(n51883), .B(n51916), .Z(n51903) );
  AND U51800 ( .A(n51917), .B(n51918), .Z(n51915) );
  XOR U51801 ( .A(n51919), .B(n51913), .Z(n51917) );
  XNOR U51802 ( .A(n51870), .B(n51909), .Z(n51911) );
  XNOR U51803 ( .A(n51920), .B(n51921), .Z(n51870) );
  AND U51804 ( .A(n1994), .B(n51922), .Z(n51921) );
  XNOR U51805 ( .A(n51923), .B(n51924), .Z(n51922) );
  XOR U51806 ( .A(n51925), .B(n51926), .Z(n51909) );
  AND U51807 ( .A(n51927), .B(n51928), .Z(n51926) );
  XNOR U51808 ( .A(n51925), .B(n51883), .Z(n51928) );
  XOR U51809 ( .A(n51929), .B(n51918), .Z(n51883) );
  XNOR U51810 ( .A(n51930), .B(n51913), .Z(n51918) );
  XOR U51811 ( .A(n51931), .B(n51932), .Z(n51913) );
  AND U51812 ( .A(n51933), .B(n51934), .Z(n51932) );
  XOR U51813 ( .A(n51935), .B(n51931), .Z(n51933) );
  XNOR U51814 ( .A(n51936), .B(n51937), .Z(n51930) );
  AND U51815 ( .A(n51938), .B(n51939), .Z(n51937) );
  XOR U51816 ( .A(n51936), .B(n51940), .Z(n51938) );
  XNOR U51817 ( .A(n51919), .B(n51916), .Z(n51929) );
  AND U51818 ( .A(n51941), .B(n51942), .Z(n51916) );
  XOR U51819 ( .A(n51943), .B(n51944), .Z(n51919) );
  AND U51820 ( .A(n51945), .B(n51946), .Z(n51944) );
  XOR U51821 ( .A(n51943), .B(n51947), .Z(n51945) );
  XNOR U51822 ( .A(n51880), .B(n51925), .Z(n51927) );
  XNOR U51823 ( .A(n51948), .B(n51949), .Z(n51880) );
  AND U51824 ( .A(n1994), .B(n51950), .Z(n51949) );
  XNOR U51825 ( .A(n51951), .B(n51952), .Z(n51950) );
  XOR U51826 ( .A(n51953), .B(n51954), .Z(n51925) );
  AND U51827 ( .A(n51955), .B(n51956), .Z(n51954) );
  XNOR U51828 ( .A(n51953), .B(n51941), .Z(n51956) );
  IV U51829 ( .A(n51891), .Z(n51941) );
  XNOR U51830 ( .A(n51957), .B(n51934), .Z(n51891) );
  XNOR U51831 ( .A(n51958), .B(n51940), .Z(n51934) );
  XNOR U51832 ( .A(n51959), .B(n51960), .Z(n51940) );
  NOR U51833 ( .A(n51961), .B(n51962), .Z(n51960) );
  XOR U51834 ( .A(n51959), .B(n51963), .Z(n51961) );
  XNOR U51835 ( .A(n51939), .B(n51931), .Z(n51958) );
  XOR U51836 ( .A(n51964), .B(n51965), .Z(n51931) );
  AND U51837 ( .A(n51966), .B(n51967), .Z(n51965) );
  XOR U51838 ( .A(n51964), .B(n51968), .Z(n51966) );
  XNOR U51839 ( .A(n51969), .B(n51936), .Z(n51939) );
  XOR U51840 ( .A(n51970), .B(n51971), .Z(n51936) );
  AND U51841 ( .A(n51972), .B(n51973), .Z(n51971) );
  XNOR U51842 ( .A(n51974), .B(n51975), .Z(n51972) );
  IV U51843 ( .A(n51970), .Z(n51974) );
  XNOR U51844 ( .A(n51976), .B(n51977), .Z(n51969) );
  NOR U51845 ( .A(n51978), .B(n51979), .Z(n51977) );
  XNOR U51846 ( .A(n51976), .B(n51980), .Z(n51978) );
  XNOR U51847 ( .A(n51935), .B(n51942), .Z(n51957) );
  NOR U51848 ( .A(n51897), .B(n51981), .Z(n51942) );
  XOR U51849 ( .A(n51947), .B(n51946), .Z(n51935) );
  XNOR U51850 ( .A(n51982), .B(n51943), .Z(n51946) );
  XOR U51851 ( .A(n51983), .B(n51984), .Z(n51943) );
  AND U51852 ( .A(n51985), .B(n51986), .Z(n51984) );
  XNOR U51853 ( .A(n51987), .B(n51988), .Z(n51985) );
  IV U51854 ( .A(n51983), .Z(n51987) );
  XNOR U51855 ( .A(n51989), .B(n51990), .Z(n51982) );
  NOR U51856 ( .A(n51991), .B(n51992), .Z(n51990) );
  XNOR U51857 ( .A(n51989), .B(n51993), .Z(n51991) );
  XOR U51858 ( .A(n51994), .B(n51995), .Z(n51947) );
  NOR U51859 ( .A(n51996), .B(n51997), .Z(n51995) );
  XNOR U51860 ( .A(n51994), .B(n51998), .Z(n51996) );
  XNOR U51861 ( .A(n51888), .B(n51953), .Z(n51955) );
  XNOR U51862 ( .A(n51999), .B(n52000), .Z(n51888) );
  AND U51863 ( .A(n1994), .B(n52001), .Z(n52000) );
  XNOR U51864 ( .A(n52002), .B(n52003), .Z(n52001) );
  AND U51865 ( .A(n51894), .B(n51897), .Z(n51953) );
  XOR U51866 ( .A(n52004), .B(n51981), .Z(n51897) );
  XNOR U51867 ( .A(p_input[1616]), .B(p_input[2048]), .Z(n51981) );
  XNOR U51868 ( .A(n51968), .B(n51967), .Z(n52004) );
  XNOR U51869 ( .A(n52005), .B(n51975), .Z(n51967) );
  XNOR U51870 ( .A(n51963), .B(n51962), .Z(n51975) );
  XNOR U51871 ( .A(n52006), .B(n51959), .Z(n51962) );
  XNOR U51872 ( .A(p_input[1626]), .B(p_input[2058]), .Z(n51959) );
  XOR U51873 ( .A(p_input[1627]), .B(n29030), .Z(n52006) );
  XOR U51874 ( .A(p_input[1628]), .B(p_input[2060]), .Z(n51963) );
  XOR U51875 ( .A(n51973), .B(n52007), .Z(n52005) );
  IV U51876 ( .A(n51964), .Z(n52007) );
  XOR U51877 ( .A(p_input[1617]), .B(p_input[2049]), .Z(n51964) );
  XNOR U51878 ( .A(n52008), .B(n51980), .Z(n51973) );
  XNOR U51879 ( .A(p_input[1631]), .B(n29033), .Z(n51980) );
  XOR U51880 ( .A(n51970), .B(n51979), .Z(n52008) );
  XOR U51881 ( .A(n52009), .B(n51976), .Z(n51979) );
  XOR U51882 ( .A(p_input[1629]), .B(p_input[2061]), .Z(n51976) );
  XOR U51883 ( .A(p_input[1630]), .B(n29035), .Z(n52009) );
  XOR U51884 ( .A(p_input[1625]), .B(p_input[2057]), .Z(n51970) );
  XOR U51885 ( .A(n51988), .B(n51986), .Z(n51968) );
  XNOR U51886 ( .A(n52010), .B(n51993), .Z(n51986) );
  XOR U51887 ( .A(p_input[1624]), .B(p_input[2056]), .Z(n51993) );
  XOR U51888 ( .A(n51983), .B(n51992), .Z(n52010) );
  XOR U51889 ( .A(n52011), .B(n51989), .Z(n51992) );
  XOR U51890 ( .A(p_input[1622]), .B(p_input[2054]), .Z(n51989) );
  XOR U51891 ( .A(p_input[1623]), .B(n30404), .Z(n52011) );
  XOR U51892 ( .A(p_input[1618]), .B(p_input[2050]), .Z(n51983) );
  XNOR U51893 ( .A(n51998), .B(n51997), .Z(n51988) );
  XOR U51894 ( .A(n52012), .B(n51994), .Z(n51997) );
  XOR U51895 ( .A(p_input[1619]), .B(p_input[2051]), .Z(n51994) );
  XOR U51896 ( .A(p_input[1620]), .B(n30406), .Z(n52012) );
  XOR U51897 ( .A(p_input[1621]), .B(p_input[2053]), .Z(n51998) );
  XNOR U51898 ( .A(n52013), .B(n52014), .Z(n51894) );
  AND U51899 ( .A(n1994), .B(n52015), .Z(n52014) );
  XNOR U51900 ( .A(n52016), .B(n52017), .Z(n1994) );
  AND U51901 ( .A(n52018), .B(n52019), .Z(n52017) );
  XOR U51902 ( .A(n51908), .B(n52016), .Z(n52019) );
  XNOR U51903 ( .A(n52020), .B(n52016), .Z(n52018) );
  XOR U51904 ( .A(n52021), .B(n52022), .Z(n52016) );
  AND U51905 ( .A(n52023), .B(n52024), .Z(n52022) );
  XOR U51906 ( .A(n51923), .B(n52021), .Z(n52024) );
  XOR U51907 ( .A(n52021), .B(n51924), .Z(n52023) );
  XOR U51908 ( .A(n52025), .B(n52026), .Z(n52021) );
  AND U51909 ( .A(n52027), .B(n52028), .Z(n52026) );
  XOR U51910 ( .A(n51951), .B(n52025), .Z(n52028) );
  XOR U51911 ( .A(n52025), .B(n51952), .Z(n52027) );
  XOR U51912 ( .A(n52029), .B(n52030), .Z(n52025) );
  AND U51913 ( .A(n52031), .B(n52032), .Z(n52030) );
  XOR U51914 ( .A(n52029), .B(n52002), .Z(n52032) );
  XNOR U51915 ( .A(n52033), .B(n52034), .Z(n51854) );
  AND U51916 ( .A(n1998), .B(n52035), .Z(n52034) );
  XNOR U51917 ( .A(n52036), .B(n52037), .Z(n1998) );
  AND U51918 ( .A(n52038), .B(n52039), .Z(n52037) );
  XOR U51919 ( .A(n52036), .B(n51864), .Z(n52039) );
  XNOR U51920 ( .A(n52036), .B(n51824), .Z(n52038) );
  XOR U51921 ( .A(n52040), .B(n52041), .Z(n52036) );
  AND U51922 ( .A(n52042), .B(n52043), .Z(n52041) );
  XOR U51923 ( .A(n52040), .B(n51832), .Z(n52042) );
  XOR U51924 ( .A(n52044), .B(n52045), .Z(n51815) );
  AND U51925 ( .A(n2002), .B(n52035), .Z(n52045) );
  XNOR U51926 ( .A(n52033), .B(n52044), .Z(n52035) );
  XNOR U51927 ( .A(n52046), .B(n52047), .Z(n2002) );
  AND U51928 ( .A(n52048), .B(n52049), .Z(n52047) );
  XNOR U51929 ( .A(n52050), .B(n52046), .Z(n52049) );
  IV U51930 ( .A(n51864), .Z(n52050) );
  XOR U51931 ( .A(n52020), .B(n52051), .Z(n51864) );
  AND U51932 ( .A(n2005), .B(n52052), .Z(n52051) );
  XOR U51933 ( .A(n51907), .B(n51904), .Z(n52052) );
  IV U51934 ( .A(n52020), .Z(n51907) );
  XNOR U51935 ( .A(n51824), .B(n52046), .Z(n52048) );
  XOR U51936 ( .A(n52053), .B(n52054), .Z(n51824) );
  AND U51937 ( .A(n2021), .B(n52055), .Z(n52054) );
  XOR U51938 ( .A(n52040), .B(n52056), .Z(n52046) );
  AND U51939 ( .A(n52057), .B(n52043), .Z(n52056) );
  XNOR U51940 ( .A(n51874), .B(n52040), .Z(n52043) );
  XOR U51941 ( .A(n51924), .B(n52058), .Z(n51874) );
  AND U51942 ( .A(n2005), .B(n52059), .Z(n52058) );
  XOR U51943 ( .A(n51920), .B(n51924), .Z(n52059) );
  XNOR U51944 ( .A(n52060), .B(n52040), .Z(n52057) );
  IV U51945 ( .A(n51832), .Z(n52060) );
  XOR U51946 ( .A(n52061), .B(n52062), .Z(n51832) );
  AND U51947 ( .A(n2021), .B(n52063), .Z(n52062) );
  XOR U51948 ( .A(n52064), .B(n52065), .Z(n52040) );
  AND U51949 ( .A(n52066), .B(n52067), .Z(n52065) );
  XNOR U51950 ( .A(n51884), .B(n52064), .Z(n52067) );
  XOR U51951 ( .A(n51952), .B(n52068), .Z(n51884) );
  AND U51952 ( .A(n2005), .B(n52069), .Z(n52068) );
  XOR U51953 ( .A(n51948), .B(n51952), .Z(n52069) );
  XOR U51954 ( .A(n52064), .B(n51841), .Z(n52066) );
  XOR U51955 ( .A(n52070), .B(n52071), .Z(n51841) );
  AND U51956 ( .A(n2021), .B(n52072), .Z(n52071) );
  XOR U51957 ( .A(n52073), .B(n52074), .Z(n52064) );
  AND U51958 ( .A(n52075), .B(n52076), .Z(n52074) );
  XNOR U51959 ( .A(n52073), .B(n51892), .Z(n52076) );
  XOR U51960 ( .A(n52003), .B(n52077), .Z(n51892) );
  AND U51961 ( .A(n2005), .B(n52078), .Z(n52077) );
  XOR U51962 ( .A(n51999), .B(n52003), .Z(n52078) );
  XNOR U51963 ( .A(n52079), .B(n52073), .Z(n52075) );
  IV U51964 ( .A(n51851), .Z(n52079) );
  XOR U51965 ( .A(n52080), .B(n52081), .Z(n51851) );
  AND U51966 ( .A(n2021), .B(n52082), .Z(n52081) );
  AND U51967 ( .A(n52044), .B(n52033), .Z(n52073) );
  XNOR U51968 ( .A(n52083), .B(n52084), .Z(n52033) );
  AND U51969 ( .A(n2005), .B(n52015), .Z(n52084) );
  XNOR U51970 ( .A(n52013), .B(n52083), .Z(n52015) );
  XNOR U51971 ( .A(n52085), .B(n52086), .Z(n2005) );
  AND U51972 ( .A(n52087), .B(n52088), .Z(n52086) );
  XNOR U51973 ( .A(n52085), .B(n51904), .Z(n52088) );
  IV U51974 ( .A(n51908), .Z(n51904) );
  XOR U51975 ( .A(n52089), .B(n52090), .Z(n51908) );
  AND U51976 ( .A(n2009), .B(n52091), .Z(n52090) );
  XOR U51977 ( .A(n52092), .B(n52089), .Z(n52091) );
  XNOR U51978 ( .A(n52085), .B(n52020), .Z(n52087) );
  XOR U51979 ( .A(n52093), .B(n52094), .Z(n52020) );
  AND U51980 ( .A(n2017), .B(n52055), .Z(n52094) );
  XOR U51981 ( .A(n52053), .B(n52093), .Z(n52055) );
  XOR U51982 ( .A(n52095), .B(n52096), .Z(n52085) );
  AND U51983 ( .A(n52097), .B(n52098), .Z(n52096) );
  XNOR U51984 ( .A(n52095), .B(n51920), .Z(n52098) );
  IV U51985 ( .A(n51923), .Z(n51920) );
  XOR U51986 ( .A(n52099), .B(n52100), .Z(n51923) );
  AND U51987 ( .A(n2009), .B(n52101), .Z(n52100) );
  XOR U51988 ( .A(n52102), .B(n52099), .Z(n52101) );
  XOR U51989 ( .A(n51924), .B(n52095), .Z(n52097) );
  XOR U51990 ( .A(n52103), .B(n52104), .Z(n51924) );
  AND U51991 ( .A(n2017), .B(n52063), .Z(n52104) );
  XOR U51992 ( .A(n52103), .B(n52061), .Z(n52063) );
  XOR U51993 ( .A(n52105), .B(n52106), .Z(n52095) );
  AND U51994 ( .A(n52107), .B(n52108), .Z(n52106) );
  XNOR U51995 ( .A(n52105), .B(n51948), .Z(n52108) );
  IV U51996 ( .A(n51951), .Z(n51948) );
  XOR U51997 ( .A(n52109), .B(n52110), .Z(n51951) );
  AND U51998 ( .A(n2009), .B(n52111), .Z(n52110) );
  XNOR U51999 ( .A(n52112), .B(n52109), .Z(n52111) );
  XOR U52000 ( .A(n51952), .B(n52105), .Z(n52107) );
  XOR U52001 ( .A(n52113), .B(n52114), .Z(n51952) );
  AND U52002 ( .A(n2017), .B(n52072), .Z(n52114) );
  XOR U52003 ( .A(n52113), .B(n52070), .Z(n52072) );
  XOR U52004 ( .A(n52029), .B(n52115), .Z(n52105) );
  AND U52005 ( .A(n52031), .B(n52116), .Z(n52115) );
  XNOR U52006 ( .A(n52029), .B(n51999), .Z(n52116) );
  IV U52007 ( .A(n52002), .Z(n51999) );
  XOR U52008 ( .A(n52117), .B(n52118), .Z(n52002) );
  AND U52009 ( .A(n2009), .B(n52119), .Z(n52118) );
  XOR U52010 ( .A(n52120), .B(n52117), .Z(n52119) );
  XOR U52011 ( .A(n52003), .B(n52029), .Z(n52031) );
  XOR U52012 ( .A(n52121), .B(n52122), .Z(n52003) );
  AND U52013 ( .A(n2017), .B(n52082), .Z(n52122) );
  XOR U52014 ( .A(n52121), .B(n52080), .Z(n52082) );
  AND U52015 ( .A(n52083), .B(n52013), .Z(n52029) );
  XNOR U52016 ( .A(n52123), .B(n52124), .Z(n52013) );
  AND U52017 ( .A(n2009), .B(n52125), .Z(n52124) );
  XNOR U52018 ( .A(n52126), .B(n52123), .Z(n52125) );
  XNOR U52019 ( .A(n52127), .B(n52128), .Z(n2009) );
  AND U52020 ( .A(n52129), .B(n52130), .Z(n52128) );
  XOR U52021 ( .A(n52092), .B(n52127), .Z(n52130) );
  AND U52022 ( .A(n52131), .B(n52132), .Z(n52092) );
  XNOR U52023 ( .A(n52089), .B(n52127), .Z(n52129) );
  XNOR U52024 ( .A(n52133), .B(n52134), .Z(n52089) );
  AND U52025 ( .A(n2013), .B(n52135), .Z(n52134) );
  XNOR U52026 ( .A(n52136), .B(n52137), .Z(n52135) );
  XOR U52027 ( .A(n52138), .B(n52139), .Z(n52127) );
  AND U52028 ( .A(n52140), .B(n52141), .Z(n52139) );
  XNOR U52029 ( .A(n52138), .B(n52131), .Z(n52141) );
  IV U52030 ( .A(n52102), .Z(n52131) );
  XOR U52031 ( .A(n52142), .B(n52143), .Z(n52102) );
  XOR U52032 ( .A(n52144), .B(n52132), .Z(n52143) );
  AND U52033 ( .A(n52112), .B(n52145), .Z(n52132) );
  AND U52034 ( .A(n52146), .B(n52147), .Z(n52144) );
  XOR U52035 ( .A(n52148), .B(n52142), .Z(n52146) );
  XNOR U52036 ( .A(n52099), .B(n52138), .Z(n52140) );
  XNOR U52037 ( .A(n52149), .B(n52150), .Z(n52099) );
  AND U52038 ( .A(n2013), .B(n52151), .Z(n52150) );
  XNOR U52039 ( .A(n52152), .B(n52153), .Z(n52151) );
  XOR U52040 ( .A(n52154), .B(n52155), .Z(n52138) );
  AND U52041 ( .A(n52156), .B(n52157), .Z(n52155) );
  XNOR U52042 ( .A(n52154), .B(n52112), .Z(n52157) );
  XOR U52043 ( .A(n52158), .B(n52147), .Z(n52112) );
  XNOR U52044 ( .A(n52159), .B(n52142), .Z(n52147) );
  XOR U52045 ( .A(n52160), .B(n52161), .Z(n52142) );
  AND U52046 ( .A(n52162), .B(n52163), .Z(n52161) );
  XOR U52047 ( .A(n52164), .B(n52160), .Z(n52162) );
  XNOR U52048 ( .A(n52165), .B(n52166), .Z(n52159) );
  AND U52049 ( .A(n52167), .B(n52168), .Z(n52166) );
  XOR U52050 ( .A(n52165), .B(n52169), .Z(n52167) );
  XNOR U52051 ( .A(n52148), .B(n52145), .Z(n52158) );
  AND U52052 ( .A(n52170), .B(n52171), .Z(n52145) );
  XOR U52053 ( .A(n52172), .B(n52173), .Z(n52148) );
  AND U52054 ( .A(n52174), .B(n52175), .Z(n52173) );
  XOR U52055 ( .A(n52172), .B(n52176), .Z(n52174) );
  XNOR U52056 ( .A(n52109), .B(n52154), .Z(n52156) );
  XNOR U52057 ( .A(n52177), .B(n52178), .Z(n52109) );
  AND U52058 ( .A(n2013), .B(n52179), .Z(n52178) );
  XNOR U52059 ( .A(n52180), .B(n52181), .Z(n52179) );
  XOR U52060 ( .A(n52182), .B(n52183), .Z(n52154) );
  AND U52061 ( .A(n52184), .B(n52185), .Z(n52183) );
  XNOR U52062 ( .A(n52182), .B(n52170), .Z(n52185) );
  IV U52063 ( .A(n52120), .Z(n52170) );
  XNOR U52064 ( .A(n52186), .B(n52163), .Z(n52120) );
  XNOR U52065 ( .A(n52187), .B(n52169), .Z(n52163) );
  XNOR U52066 ( .A(n52188), .B(n52189), .Z(n52169) );
  NOR U52067 ( .A(n52190), .B(n52191), .Z(n52189) );
  XOR U52068 ( .A(n52188), .B(n52192), .Z(n52190) );
  XNOR U52069 ( .A(n52168), .B(n52160), .Z(n52187) );
  XOR U52070 ( .A(n52193), .B(n52194), .Z(n52160) );
  AND U52071 ( .A(n52195), .B(n52196), .Z(n52194) );
  XOR U52072 ( .A(n52193), .B(n52197), .Z(n52195) );
  XNOR U52073 ( .A(n52198), .B(n52165), .Z(n52168) );
  XOR U52074 ( .A(n52199), .B(n52200), .Z(n52165) );
  AND U52075 ( .A(n52201), .B(n52202), .Z(n52200) );
  XNOR U52076 ( .A(n52203), .B(n52204), .Z(n52201) );
  IV U52077 ( .A(n52199), .Z(n52203) );
  XNOR U52078 ( .A(n52205), .B(n52206), .Z(n52198) );
  NOR U52079 ( .A(n52207), .B(n52208), .Z(n52206) );
  XNOR U52080 ( .A(n52205), .B(n52209), .Z(n52207) );
  XNOR U52081 ( .A(n52164), .B(n52171), .Z(n52186) );
  NOR U52082 ( .A(n52126), .B(n52210), .Z(n52171) );
  XOR U52083 ( .A(n52176), .B(n52175), .Z(n52164) );
  XNOR U52084 ( .A(n52211), .B(n52172), .Z(n52175) );
  XOR U52085 ( .A(n52212), .B(n52213), .Z(n52172) );
  AND U52086 ( .A(n52214), .B(n52215), .Z(n52213) );
  XNOR U52087 ( .A(n52216), .B(n52217), .Z(n52214) );
  IV U52088 ( .A(n52212), .Z(n52216) );
  XNOR U52089 ( .A(n52218), .B(n52219), .Z(n52211) );
  NOR U52090 ( .A(n52220), .B(n52221), .Z(n52219) );
  XNOR U52091 ( .A(n52218), .B(n52222), .Z(n52220) );
  XOR U52092 ( .A(n52223), .B(n52224), .Z(n52176) );
  NOR U52093 ( .A(n52225), .B(n52226), .Z(n52224) );
  XNOR U52094 ( .A(n52223), .B(n52227), .Z(n52225) );
  XNOR U52095 ( .A(n52117), .B(n52182), .Z(n52184) );
  XNOR U52096 ( .A(n52228), .B(n52229), .Z(n52117) );
  AND U52097 ( .A(n2013), .B(n52230), .Z(n52229) );
  XNOR U52098 ( .A(n52231), .B(n52232), .Z(n52230) );
  AND U52099 ( .A(n52123), .B(n52126), .Z(n52182) );
  XOR U52100 ( .A(n52233), .B(n52210), .Z(n52126) );
  XNOR U52101 ( .A(p_input[1632]), .B(p_input[2048]), .Z(n52210) );
  XNOR U52102 ( .A(n52197), .B(n52196), .Z(n52233) );
  XNOR U52103 ( .A(n52234), .B(n52204), .Z(n52196) );
  XNOR U52104 ( .A(n52192), .B(n52191), .Z(n52204) );
  XNOR U52105 ( .A(n52235), .B(n52188), .Z(n52191) );
  XNOR U52106 ( .A(p_input[1642]), .B(p_input[2058]), .Z(n52188) );
  XOR U52107 ( .A(p_input[1643]), .B(n29030), .Z(n52235) );
  XOR U52108 ( .A(p_input[1644]), .B(p_input[2060]), .Z(n52192) );
  XOR U52109 ( .A(n52202), .B(n52236), .Z(n52234) );
  IV U52110 ( .A(n52193), .Z(n52236) );
  XOR U52111 ( .A(p_input[1633]), .B(p_input[2049]), .Z(n52193) );
  XNOR U52112 ( .A(n52237), .B(n52209), .Z(n52202) );
  XNOR U52113 ( .A(p_input[1647]), .B(n29033), .Z(n52209) );
  XOR U52114 ( .A(n52199), .B(n52208), .Z(n52237) );
  XOR U52115 ( .A(n52238), .B(n52205), .Z(n52208) );
  XOR U52116 ( .A(p_input[1645]), .B(p_input[2061]), .Z(n52205) );
  XOR U52117 ( .A(p_input[1646]), .B(n29035), .Z(n52238) );
  XOR U52118 ( .A(p_input[1641]), .B(p_input[2057]), .Z(n52199) );
  XOR U52119 ( .A(n52217), .B(n52215), .Z(n52197) );
  XNOR U52120 ( .A(n52239), .B(n52222), .Z(n52215) );
  XOR U52121 ( .A(p_input[1640]), .B(p_input[2056]), .Z(n52222) );
  XOR U52122 ( .A(n52212), .B(n52221), .Z(n52239) );
  XOR U52123 ( .A(n52240), .B(n52218), .Z(n52221) );
  XOR U52124 ( .A(p_input[1638]), .B(p_input[2054]), .Z(n52218) );
  XOR U52125 ( .A(p_input[1639]), .B(n30404), .Z(n52240) );
  XOR U52126 ( .A(p_input[1634]), .B(p_input[2050]), .Z(n52212) );
  XNOR U52127 ( .A(n52227), .B(n52226), .Z(n52217) );
  XOR U52128 ( .A(n52241), .B(n52223), .Z(n52226) );
  XOR U52129 ( .A(p_input[1635]), .B(p_input[2051]), .Z(n52223) );
  XOR U52130 ( .A(p_input[1636]), .B(n30406), .Z(n52241) );
  XOR U52131 ( .A(p_input[1637]), .B(p_input[2053]), .Z(n52227) );
  XNOR U52132 ( .A(n52242), .B(n52243), .Z(n52123) );
  AND U52133 ( .A(n2013), .B(n52244), .Z(n52243) );
  XNOR U52134 ( .A(n52245), .B(n52246), .Z(n2013) );
  AND U52135 ( .A(n52247), .B(n52248), .Z(n52246) );
  XOR U52136 ( .A(n52137), .B(n52245), .Z(n52248) );
  XNOR U52137 ( .A(n52249), .B(n52245), .Z(n52247) );
  XOR U52138 ( .A(n52250), .B(n52251), .Z(n52245) );
  AND U52139 ( .A(n52252), .B(n52253), .Z(n52251) );
  XOR U52140 ( .A(n52152), .B(n52250), .Z(n52253) );
  XOR U52141 ( .A(n52250), .B(n52153), .Z(n52252) );
  XOR U52142 ( .A(n52254), .B(n52255), .Z(n52250) );
  AND U52143 ( .A(n52256), .B(n52257), .Z(n52255) );
  XOR U52144 ( .A(n52180), .B(n52254), .Z(n52257) );
  XOR U52145 ( .A(n52254), .B(n52181), .Z(n52256) );
  XOR U52146 ( .A(n52258), .B(n52259), .Z(n52254) );
  AND U52147 ( .A(n52260), .B(n52261), .Z(n52259) );
  XOR U52148 ( .A(n52258), .B(n52231), .Z(n52261) );
  XNOR U52149 ( .A(n52262), .B(n52263), .Z(n52083) );
  AND U52150 ( .A(n2017), .B(n52264), .Z(n52263) );
  XNOR U52151 ( .A(n52265), .B(n52266), .Z(n2017) );
  AND U52152 ( .A(n52267), .B(n52268), .Z(n52266) );
  XOR U52153 ( .A(n52265), .B(n52093), .Z(n52268) );
  XNOR U52154 ( .A(n52265), .B(n52053), .Z(n52267) );
  XOR U52155 ( .A(n52269), .B(n52270), .Z(n52265) );
  AND U52156 ( .A(n52271), .B(n52272), .Z(n52270) );
  XOR U52157 ( .A(n52269), .B(n52061), .Z(n52271) );
  XOR U52158 ( .A(n52273), .B(n52274), .Z(n52044) );
  AND U52159 ( .A(n2021), .B(n52264), .Z(n52274) );
  XNOR U52160 ( .A(n52262), .B(n52273), .Z(n52264) );
  XNOR U52161 ( .A(n52275), .B(n52276), .Z(n2021) );
  AND U52162 ( .A(n52277), .B(n52278), .Z(n52276) );
  XNOR U52163 ( .A(n52279), .B(n52275), .Z(n52278) );
  IV U52164 ( .A(n52093), .Z(n52279) );
  XOR U52165 ( .A(n52249), .B(n52280), .Z(n52093) );
  AND U52166 ( .A(n2024), .B(n52281), .Z(n52280) );
  XOR U52167 ( .A(n52136), .B(n52133), .Z(n52281) );
  IV U52168 ( .A(n52249), .Z(n52136) );
  XNOR U52169 ( .A(n52053), .B(n52275), .Z(n52277) );
  XOR U52170 ( .A(n52282), .B(n52283), .Z(n52053) );
  AND U52171 ( .A(n2040), .B(n52284), .Z(n52283) );
  XOR U52172 ( .A(n52269), .B(n52285), .Z(n52275) );
  AND U52173 ( .A(n52286), .B(n52272), .Z(n52285) );
  XNOR U52174 ( .A(n52103), .B(n52269), .Z(n52272) );
  XOR U52175 ( .A(n52153), .B(n52287), .Z(n52103) );
  AND U52176 ( .A(n2024), .B(n52288), .Z(n52287) );
  XOR U52177 ( .A(n52149), .B(n52153), .Z(n52288) );
  XNOR U52178 ( .A(n52289), .B(n52269), .Z(n52286) );
  IV U52179 ( .A(n52061), .Z(n52289) );
  XOR U52180 ( .A(n52290), .B(n52291), .Z(n52061) );
  AND U52181 ( .A(n2040), .B(n52292), .Z(n52291) );
  XOR U52182 ( .A(n52293), .B(n52294), .Z(n52269) );
  AND U52183 ( .A(n52295), .B(n52296), .Z(n52294) );
  XNOR U52184 ( .A(n52113), .B(n52293), .Z(n52296) );
  XOR U52185 ( .A(n52181), .B(n52297), .Z(n52113) );
  AND U52186 ( .A(n2024), .B(n52298), .Z(n52297) );
  XOR U52187 ( .A(n52177), .B(n52181), .Z(n52298) );
  XOR U52188 ( .A(n52293), .B(n52070), .Z(n52295) );
  XOR U52189 ( .A(n52299), .B(n52300), .Z(n52070) );
  AND U52190 ( .A(n2040), .B(n52301), .Z(n52300) );
  XOR U52191 ( .A(n52302), .B(n52303), .Z(n52293) );
  AND U52192 ( .A(n52304), .B(n52305), .Z(n52303) );
  XNOR U52193 ( .A(n52302), .B(n52121), .Z(n52305) );
  XOR U52194 ( .A(n52232), .B(n52306), .Z(n52121) );
  AND U52195 ( .A(n2024), .B(n52307), .Z(n52306) );
  XOR U52196 ( .A(n52228), .B(n52232), .Z(n52307) );
  XNOR U52197 ( .A(n52308), .B(n52302), .Z(n52304) );
  IV U52198 ( .A(n52080), .Z(n52308) );
  XOR U52199 ( .A(n52309), .B(n52310), .Z(n52080) );
  AND U52200 ( .A(n2040), .B(n52311), .Z(n52310) );
  AND U52201 ( .A(n52273), .B(n52262), .Z(n52302) );
  XNOR U52202 ( .A(n52312), .B(n52313), .Z(n52262) );
  AND U52203 ( .A(n2024), .B(n52244), .Z(n52313) );
  XNOR U52204 ( .A(n52242), .B(n52312), .Z(n52244) );
  XNOR U52205 ( .A(n52314), .B(n52315), .Z(n2024) );
  AND U52206 ( .A(n52316), .B(n52317), .Z(n52315) );
  XNOR U52207 ( .A(n52314), .B(n52133), .Z(n52317) );
  IV U52208 ( .A(n52137), .Z(n52133) );
  XOR U52209 ( .A(n52318), .B(n52319), .Z(n52137) );
  AND U52210 ( .A(n2028), .B(n52320), .Z(n52319) );
  XOR U52211 ( .A(n52321), .B(n52318), .Z(n52320) );
  XNOR U52212 ( .A(n52314), .B(n52249), .Z(n52316) );
  XOR U52213 ( .A(n52322), .B(n52323), .Z(n52249) );
  AND U52214 ( .A(n2036), .B(n52284), .Z(n52323) );
  XOR U52215 ( .A(n52282), .B(n52322), .Z(n52284) );
  XOR U52216 ( .A(n52324), .B(n52325), .Z(n52314) );
  AND U52217 ( .A(n52326), .B(n52327), .Z(n52325) );
  XNOR U52218 ( .A(n52324), .B(n52149), .Z(n52327) );
  IV U52219 ( .A(n52152), .Z(n52149) );
  XOR U52220 ( .A(n52328), .B(n52329), .Z(n52152) );
  AND U52221 ( .A(n2028), .B(n52330), .Z(n52329) );
  XOR U52222 ( .A(n52331), .B(n52328), .Z(n52330) );
  XOR U52223 ( .A(n52153), .B(n52324), .Z(n52326) );
  XOR U52224 ( .A(n52332), .B(n52333), .Z(n52153) );
  AND U52225 ( .A(n2036), .B(n52292), .Z(n52333) );
  XOR U52226 ( .A(n52332), .B(n52290), .Z(n52292) );
  XOR U52227 ( .A(n52334), .B(n52335), .Z(n52324) );
  AND U52228 ( .A(n52336), .B(n52337), .Z(n52335) );
  XNOR U52229 ( .A(n52334), .B(n52177), .Z(n52337) );
  IV U52230 ( .A(n52180), .Z(n52177) );
  XOR U52231 ( .A(n52338), .B(n52339), .Z(n52180) );
  AND U52232 ( .A(n2028), .B(n52340), .Z(n52339) );
  XNOR U52233 ( .A(n52341), .B(n52338), .Z(n52340) );
  XOR U52234 ( .A(n52181), .B(n52334), .Z(n52336) );
  XOR U52235 ( .A(n52342), .B(n52343), .Z(n52181) );
  AND U52236 ( .A(n2036), .B(n52301), .Z(n52343) );
  XOR U52237 ( .A(n52342), .B(n52299), .Z(n52301) );
  XOR U52238 ( .A(n52258), .B(n52344), .Z(n52334) );
  AND U52239 ( .A(n52260), .B(n52345), .Z(n52344) );
  XNOR U52240 ( .A(n52258), .B(n52228), .Z(n52345) );
  IV U52241 ( .A(n52231), .Z(n52228) );
  XOR U52242 ( .A(n52346), .B(n52347), .Z(n52231) );
  AND U52243 ( .A(n2028), .B(n52348), .Z(n52347) );
  XOR U52244 ( .A(n52349), .B(n52346), .Z(n52348) );
  XOR U52245 ( .A(n52232), .B(n52258), .Z(n52260) );
  XOR U52246 ( .A(n52350), .B(n52351), .Z(n52232) );
  AND U52247 ( .A(n2036), .B(n52311), .Z(n52351) );
  XOR U52248 ( .A(n52350), .B(n52309), .Z(n52311) );
  AND U52249 ( .A(n52312), .B(n52242), .Z(n52258) );
  XNOR U52250 ( .A(n52352), .B(n52353), .Z(n52242) );
  AND U52251 ( .A(n2028), .B(n52354), .Z(n52353) );
  XNOR U52252 ( .A(n52355), .B(n52352), .Z(n52354) );
  XNOR U52253 ( .A(n52356), .B(n52357), .Z(n2028) );
  AND U52254 ( .A(n52358), .B(n52359), .Z(n52357) );
  XOR U52255 ( .A(n52321), .B(n52356), .Z(n52359) );
  AND U52256 ( .A(n52360), .B(n52361), .Z(n52321) );
  XNOR U52257 ( .A(n52318), .B(n52356), .Z(n52358) );
  XNOR U52258 ( .A(n52362), .B(n52363), .Z(n52318) );
  AND U52259 ( .A(n2032), .B(n52364), .Z(n52363) );
  XNOR U52260 ( .A(n52365), .B(n52366), .Z(n52364) );
  XOR U52261 ( .A(n52367), .B(n52368), .Z(n52356) );
  AND U52262 ( .A(n52369), .B(n52370), .Z(n52368) );
  XNOR U52263 ( .A(n52367), .B(n52360), .Z(n52370) );
  IV U52264 ( .A(n52331), .Z(n52360) );
  XOR U52265 ( .A(n52371), .B(n52372), .Z(n52331) );
  XOR U52266 ( .A(n52373), .B(n52361), .Z(n52372) );
  AND U52267 ( .A(n52341), .B(n52374), .Z(n52361) );
  AND U52268 ( .A(n52375), .B(n52376), .Z(n52373) );
  XOR U52269 ( .A(n52377), .B(n52371), .Z(n52375) );
  XNOR U52270 ( .A(n52328), .B(n52367), .Z(n52369) );
  XNOR U52271 ( .A(n52378), .B(n52379), .Z(n52328) );
  AND U52272 ( .A(n2032), .B(n52380), .Z(n52379) );
  XNOR U52273 ( .A(n52381), .B(n52382), .Z(n52380) );
  XOR U52274 ( .A(n52383), .B(n52384), .Z(n52367) );
  AND U52275 ( .A(n52385), .B(n52386), .Z(n52384) );
  XNOR U52276 ( .A(n52383), .B(n52341), .Z(n52386) );
  XOR U52277 ( .A(n52387), .B(n52376), .Z(n52341) );
  XNOR U52278 ( .A(n52388), .B(n52371), .Z(n52376) );
  XOR U52279 ( .A(n52389), .B(n52390), .Z(n52371) );
  AND U52280 ( .A(n52391), .B(n52392), .Z(n52390) );
  XOR U52281 ( .A(n52393), .B(n52389), .Z(n52391) );
  XNOR U52282 ( .A(n52394), .B(n52395), .Z(n52388) );
  AND U52283 ( .A(n52396), .B(n52397), .Z(n52395) );
  XOR U52284 ( .A(n52394), .B(n52398), .Z(n52396) );
  XNOR U52285 ( .A(n52377), .B(n52374), .Z(n52387) );
  AND U52286 ( .A(n52399), .B(n52400), .Z(n52374) );
  XOR U52287 ( .A(n52401), .B(n52402), .Z(n52377) );
  AND U52288 ( .A(n52403), .B(n52404), .Z(n52402) );
  XOR U52289 ( .A(n52401), .B(n52405), .Z(n52403) );
  XNOR U52290 ( .A(n52338), .B(n52383), .Z(n52385) );
  XNOR U52291 ( .A(n52406), .B(n52407), .Z(n52338) );
  AND U52292 ( .A(n2032), .B(n52408), .Z(n52407) );
  XNOR U52293 ( .A(n52409), .B(n52410), .Z(n52408) );
  XOR U52294 ( .A(n52411), .B(n52412), .Z(n52383) );
  AND U52295 ( .A(n52413), .B(n52414), .Z(n52412) );
  XNOR U52296 ( .A(n52411), .B(n52399), .Z(n52414) );
  IV U52297 ( .A(n52349), .Z(n52399) );
  XNOR U52298 ( .A(n52415), .B(n52392), .Z(n52349) );
  XNOR U52299 ( .A(n52416), .B(n52398), .Z(n52392) );
  XNOR U52300 ( .A(n52417), .B(n52418), .Z(n52398) );
  NOR U52301 ( .A(n52419), .B(n52420), .Z(n52418) );
  XOR U52302 ( .A(n52417), .B(n52421), .Z(n52419) );
  XNOR U52303 ( .A(n52397), .B(n52389), .Z(n52416) );
  XOR U52304 ( .A(n52422), .B(n52423), .Z(n52389) );
  AND U52305 ( .A(n52424), .B(n52425), .Z(n52423) );
  XOR U52306 ( .A(n52422), .B(n52426), .Z(n52424) );
  XNOR U52307 ( .A(n52427), .B(n52394), .Z(n52397) );
  XOR U52308 ( .A(n52428), .B(n52429), .Z(n52394) );
  AND U52309 ( .A(n52430), .B(n52431), .Z(n52429) );
  XNOR U52310 ( .A(n52432), .B(n52433), .Z(n52430) );
  IV U52311 ( .A(n52428), .Z(n52432) );
  XNOR U52312 ( .A(n52434), .B(n52435), .Z(n52427) );
  NOR U52313 ( .A(n52436), .B(n52437), .Z(n52435) );
  XNOR U52314 ( .A(n52434), .B(n52438), .Z(n52436) );
  XNOR U52315 ( .A(n52393), .B(n52400), .Z(n52415) );
  NOR U52316 ( .A(n52355), .B(n52439), .Z(n52400) );
  XOR U52317 ( .A(n52405), .B(n52404), .Z(n52393) );
  XNOR U52318 ( .A(n52440), .B(n52401), .Z(n52404) );
  XOR U52319 ( .A(n52441), .B(n52442), .Z(n52401) );
  AND U52320 ( .A(n52443), .B(n52444), .Z(n52442) );
  XNOR U52321 ( .A(n52445), .B(n52446), .Z(n52443) );
  IV U52322 ( .A(n52441), .Z(n52445) );
  XNOR U52323 ( .A(n52447), .B(n52448), .Z(n52440) );
  NOR U52324 ( .A(n52449), .B(n52450), .Z(n52448) );
  XNOR U52325 ( .A(n52447), .B(n52451), .Z(n52449) );
  XOR U52326 ( .A(n52452), .B(n52453), .Z(n52405) );
  NOR U52327 ( .A(n52454), .B(n52455), .Z(n52453) );
  XNOR U52328 ( .A(n52452), .B(n52456), .Z(n52454) );
  XNOR U52329 ( .A(n52346), .B(n52411), .Z(n52413) );
  XNOR U52330 ( .A(n52457), .B(n52458), .Z(n52346) );
  AND U52331 ( .A(n2032), .B(n52459), .Z(n52458) );
  XNOR U52332 ( .A(n52460), .B(n52461), .Z(n52459) );
  AND U52333 ( .A(n52352), .B(n52355), .Z(n52411) );
  XOR U52334 ( .A(n52462), .B(n52439), .Z(n52355) );
  XNOR U52335 ( .A(p_input[1648]), .B(p_input[2048]), .Z(n52439) );
  XNOR U52336 ( .A(n52426), .B(n52425), .Z(n52462) );
  XNOR U52337 ( .A(n52463), .B(n52433), .Z(n52425) );
  XNOR U52338 ( .A(n52421), .B(n52420), .Z(n52433) );
  XNOR U52339 ( .A(n52464), .B(n52417), .Z(n52420) );
  XNOR U52340 ( .A(p_input[1658]), .B(p_input[2058]), .Z(n52417) );
  XOR U52341 ( .A(p_input[1659]), .B(n29030), .Z(n52464) );
  XOR U52342 ( .A(p_input[1660]), .B(p_input[2060]), .Z(n52421) );
  XOR U52343 ( .A(n52431), .B(n52465), .Z(n52463) );
  IV U52344 ( .A(n52422), .Z(n52465) );
  XOR U52345 ( .A(p_input[1649]), .B(p_input[2049]), .Z(n52422) );
  XNOR U52346 ( .A(n52466), .B(n52438), .Z(n52431) );
  XNOR U52347 ( .A(p_input[1663]), .B(n29033), .Z(n52438) );
  XOR U52348 ( .A(n52428), .B(n52437), .Z(n52466) );
  XOR U52349 ( .A(n52467), .B(n52434), .Z(n52437) );
  XOR U52350 ( .A(p_input[1661]), .B(p_input[2061]), .Z(n52434) );
  XOR U52351 ( .A(p_input[1662]), .B(n29035), .Z(n52467) );
  XOR U52352 ( .A(p_input[1657]), .B(p_input[2057]), .Z(n52428) );
  XOR U52353 ( .A(n52446), .B(n52444), .Z(n52426) );
  XNOR U52354 ( .A(n52468), .B(n52451), .Z(n52444) );
  XOR U52355 ( .A(p_input[1656]), .B(p_input[2056]), .Z(n52451) );
  XOR U52356 ( .A(n52441), .B(n52450), .Z(n52468) );
  XOR U52357 ( .A(n52469), .B(n52447), .Z(n52450) );
  XOR U52358 ( .A(p_input[1654]), .B(p_input[2054]), .Z(n52447) );
  XOR U52359 ( .A(p_input[1655]), .B(n30404), .Z(n52469) );
  XOR U52360 ( .A(p_input[1650]), .B(p_input[2050]), .Z(n52441) );
  XNOR U52361 ( .A(n52456), .B(n52455), .Z(n52446) );
  XOR U52362 ( .A(n52470), .B(n52452), .Z(n52455) );
  XOR U52363 ( .A(p_input[1651]), .B(p_input[2051]), .Z(n52452) );
  XOR U52364 ( .A(p_input[1652]), .B(n30406), .Z(n52470) );
  XOR U52365 ( .A(p_input[1653]), .B(p_input[2053]), .Z(n52456) );
  XNOR U52366 ( .A(n52471), .B(n52472), .Z(n52352) );
  AND U52367 ( .A(n2032), .B(n52473), .Z(n52472) );
  XNOR U52368 ( .A(n52474), .B(n52475), .Z(n2032) );
  AND U52369 ( .A(n52476), .B(n52477), .Z(n52475) );
  XOR U52370 ( .A(n52366), .B(n52474), .Z(n52477) );
  XNOR U52371 ( .A(n52478), .B(n52474), .Z(n52476) );
  XOR U52372 ( .A(n52479), .B(n52480), .Z(n52474) );
  AND U52373 ( .A(n52481), .B(n52482), .Z(n52480) );
  XOR U52374 ( .A(n52381), .B(n52479), .Z(n52482) );
  XOR U52375 ( .A(n52479), .B(n52382), .Z(n52481) );
  XOR U52376 ( .A(n52483), .B(n52484), .Z(n52479) );
  AND U52377 ( .A(n52485), .B(n52486), .Z(n52484) );
  XOR U52378 ( .A(n52409), .B(n52483), .Z(n52486) );
  XOR U52379 ( .A(n52483), .B(n52410), .Z(n52485) );
  XOR U52380 ( .A(n52487), .B(n52488), .Z(n52483) );
  AND U52381 ( .A(n52489), .B(n52490), .Z(n52488) );
  XOR U52382 ( .A(n52487), .B(n52460), .Z(n52490) );
  XNOR U52383 ( .A(n52491), .B(n52492), .Z(n52312) );
  AND U52384 ( .A(n2036), .B(n52493), .Z(n52492) );
  XNOR U52385 ( .A(n52494), .B(n52495), .Z(n2036) );
  AND U52386 ( .A(n52496), .B(n52497), .Z(n52495) );
  XOR U52387 ( .A(n52494), .B(n52322), .Z(n52497) );
  XNOR U52388 ( .A(n52494), .B(n52282), .Z(n52496) );
  XOR U52389 ( .A(n52498), .B(n52499), .Z(n52494) );
  AND U52390 ( .A(n52500), .B(n52501), .Z(n52499) );
  XOR U52391 ( .A(n52498), .B(n52290), .Z(n52500) );
  XOR U52392 ( .A(n52502), .B(n52503), .Z(n52273) );
  AND U52393 ( .A(n2040), .B(n52493), .Z(n52503) );
  XNOR U52394 ( .A(n52491), .B(n52502), .Z(n52493) );
  XNOR U52395 ( .A(n52504), .B(n52505), .Z(n2040) );
  AND U52396 ( .A(n52506), .B(n52507), .Z(n52505) );
  XNOR U52397 ( .A(n52508), .B(n52504), .Z(n52507) );
  IV U52398 ( .A(n52322), .Z(n52508) );
  XOR U52399 ( .A(n52478), .B(n52509), .Z(n52322) );
  AND U52400 ( .A(n2043), .B(n52510), .Z(n52509) );
  XOR U52401 ( .A(n52365), .B(n52362), .Z(n52510) );
  IV U52402 ( .A(n52478), .Z(n52365) );
  XNOR U52403 ( .A(n52282), .B(n52504), .Z(n52506) );
  XOR U52404 ( .A(n52511), .B(n52512), .Z(n52282) );
  AND U52405 ( .A(n2059), .B(n52513), .Z(n52512) );
  XOR U52406 ( .A(n52498), .B(n52514), .Z(n52504) );
  AND U52407 ( .A(n52515), .B(n52501), .Z(n52514) );
  XNOR U52408 ( .A(n52332), .B(n52498), .Z(n52501) );
  XOR U52409 ( .A(n52382), .B(n52516), .Z(n52332) );
  AND U52410 ( .A(n2043), .B(n52517), .Z(n52516) );
  XOR U52411 ( .A(n52378), .B(n52382), .Z(n52517) );
  XNOR U52412 ( .A(n52518), .B(n52498), .Z(n52515) );
  IV U52413 ( .A(n52290), .Z(n52518) );
  XOR U52414 ( .A(n52519), .B(n52520), .Z(n52290) );
  AND U52415 ( .A(n2059), .B(n52521), .Z(n52520) );
  XOR U52416 ( .A(n52522), .B(n52523), .Z(n52498) );
  AND U52417 ( .A(n52524), .B(n52525), .Z(n52523) );
  XNOR U52418 ( .A(n52342), .B(n52522), .Z(n52525) );
  XOR U52419 ( .A(n52410), .B(n52526), .Z(n52342) );
  AND U52420 ( .A(n2043), .B(n52527), .Z(n52526) );
  XOR U52421 ( .A(n52406), .B(n52410), .Z(n52527) );
  XOR U52422 ( .A(n52522), .B(n52299), .Z(n52524) );
  XOR U52423 ( .A(n52528), .B(n52529), .Z(n52299) );
  AND U52424 ( .A(n2059), .B(n52530), .Z(n52529) );
  XOR U52425 ( .A(n52531), .B(n52532), .Z(n52522) );
  AND U52426 ( .A(n52533), .B(n52534), .Z(n52532) );
  XNOR U52427 ( .A(n52531), .B(n52350), .Z(n52534) );
  XOR U52428 ( .A(n52461), .B(n52535), .Z(n52350) );
  AND U52429 ( .A(n2043), .B(n52536), .Z(n52535) );
  XOR U52430 ( .A(n52457), .B(n52461), .Z(n52536) );
  XNOR U52431 ( .A(n52537), .B(n52531), .Z(n52533) );
  IV U52432 ( .A(n52309), .Z(n52537) );
  XOR U52433 ( .A(n52538), .B(n52539), .Z(n52309) );
  AND U52434 ( .A(n2059), .B(n52540), .Z(n52539) );
  AND U52435 ( .A(n52502), .B(n52491), .Z(n52531) );
  XNOR U52436 ( .A(n52541), .B(n52542), .Z(n52491) );
  AND U52437 ( .A(n2043), .B(n52473), .Z(n52542) );
  XNOR U52438 ( .A(n52471), .B(n52541), .Z(n52473) );
  XNOR U52439 ( .A(n52543), .B(n52544), .Z(n2043) );
  AND U52440 ( .A(n52545), .B(n52546), .Z(n52544) );
  XNOR U52441 ( .A(n52543), .B(n52362), .Z(n52546) );
  IV U52442 ( .A(n52366), .Z(n52362) );
  XOR U52443 ( .A(n52547), .B(n52548), .Z(n52366) );
  AND U52444 ( .A(n2047), .B(n52549), .Z(n52548) );
  XOR U52445 ( .A(n52550), .B(n52547), .Z(n52549) );
  XNOR U52446 ( .A(n52543), .B(n52478), .Z(n52545) );
  XOR U52447 ( .A(n52551), .B(n52552), .Z(n52478) );
  AND U52448 ( .A(n2055), .B(n52513), .Z(n52552) );
  XOR U52449 ( .A(n52511), .B(n52551), .Z(n52513) );
  XOR U52450 ( .A(n52553), .B(n52554), .Z(n52543) );
  AND U52451 ( .A(n52555), .B(n52556), .Z(n52554) );
  XNOR U52452 ( .A(n52553), .B(n52378), .Z(n52556) );
  IV U52453 ( .A(n52381), .Z(n52378) );
  XOR U52454 ( .A(n52557), .B(n52558), .Z(n52381) );
  AND U52455 ( .A(n2047), .B(n52559), .Z(n52558) );
  XOR U52456 ( .A(n52560), .B(n52557), .Z(n52559) );
  XOR U52457 ( .A(n52382), .B(n52553), .Z(n52555) );
  XOR U52458 ( .A(n52561), .B(n52562), .Z(n52382) );
  AND U52459 ( .A(n2055), .B(n52521), .Z(n52562) );
  XOR U52460 ( .A(n52561), .B(n52519), .Z(n52521) );
  XOR U52461 ( .A(n52563), .B(n52564), .Z(n52553) );
  AND U52462 ( .A(n52565), .B(n52566), .Z(n52564) );
  XNOR U52463 ( .A(n52563), .B(n52406), .Z(n52566) );
  IV U52464 ( .A(n52409), .Z(n52406) );
  XOR U52465 ( .A(n52567), .B(n52568), .Z(n52409) );
  AND U52466 ( .A(n2047), .B(n52569), .Z(n52568) );
  XNOR U52467 ( .A(n52570), .B(n52567), .Z(n52569) );
  XOR U52468 ( .A(n52410), .B(n52563), .Z(n52565) );
  XOR U52469 ( .A(n52571), .B(n52572), .Z(n52410) );
  AND U52470 ( .A(n2055), .B(n52530), .Z(n52572) );
  XOR U52471 ( .A(n52571), .B(n52528), .Z(n52530) );
  XOR U52472 ( .A(n52487), .B(n52573), .Z(n52563) );
  AND U52473 ( .A(n52489), .B(n52574), .Z(n52573) );
  XNOR U52474 ( .A(n52487), .B(n52457), .Z(n52574) );
  IV U52475 ( .A(n52460), .Z(n52457) );
  XOR U52476 ( .A(n52575), .B(n52576), .Z(n52460) );
  AND U52477 ( .A(n2047), .B(n52577), .Z(n52576) );
  XOR U52478 ( .A(n52578), .B(n52575), .Z(n52577) );
  XOR U52479 ( .A(n52461), .B(n52487), .Z(n52489) );
  XOR U52480 ( .A(n52579), .B(n52580), .Z(n52461) );
  AND U52481 ( .A(n2055), .B(n52540), .Z(n52580) );
  XOR U52482 ( .A(n52579), .B(n52538), .Z(n52540) );
  AND U52483 ( .A(n52541), .B(n52471), .Z(n52487) );
  XNOR U52484 ( .A(n52581), .B(n52582), .Z(n52471) );
  AND U52485 ( .A(n2047), .B(n52583), .Z(n52582) );
  XNOR U52486 ( .A(n52584), .B(n52581), .Z(n52583) );
  XNOR U52487 ( .A(n52585), .B(n52586), .Z(n2047) );
  AND U52488 ( .A(n52587), .B(n52588), .Z(n52586) );
  XOR U52489 ( .A(n52550), .B(n52585), .Z(n52588) );
  AND U52490 ( .A(n52589), .B(n52590), .Z(n52550) );
  XNOR U52491 ( .A(n52547), .B(n52585), .Z(n52587) );
  XNOR U52492 ( .A(n52591), .B(n52592), .Z(n52547) );
  AND U52493 ( .A(n2051), .B(n52593), .Z(n52592) );
  XNOR U52494 ( .A(n52594), .B(n52595), .Z(n52593) );
  XOR U52495 ( .A(n52596), .B(n52597), .Z(n52585) );
  AND U52496 ( .A(n52598), .B(n52599), .Z(n52597) );
  XNOR U52497 ( .A(n52596), .B(n52589), .Z(n52599) );
  IV U52498 ( .A(n52560), .Z(n52589) );
  XOR U52499 ( .A(n52600), .B(n52601), .Z(n52560) );
  XOR U52500 ( .A(n52602), .B(n52590), .Z(n52601) );
  AND U52501 ( .A(n52570), .B(n52603), .Z(n52590) );
  AND U52502 ( .A(n52604), .B(n52605), .Z(n52602) );
  XOR U52503 ( .A(n52606), .B(n52600), .Z(n52604) );
  XNOR U52504 ( .A(n52557), .B(n52596), .Z(n52598) );
  XNOR U52505 ( .A(n52607), .B(n52608), .Z(n52557) );
  AND U52506 ( .A(n2051), .B(n52609), .Z(n52608) );
  XNOR U52507 ( .A(n52610), .B(n52611), .Z(n52609) );
  XOR U52508 ( .A(n52612), .B(n52613), .Z(n52596) );
  AND U52509 ( .A(n52614), .B(n52615), .Z(n52613) );
  XNOR U52510 ( .A(n52612), .B(n52570), .Z(n52615) );
  XOR U52511 ( .A(n52616), .B(n52605), .Z(n52570) );
  XNOR U52512 ( .A(n52617), .B(n52600), .Z(n52605) );
  XOR U52513 ( .A(n52618), .B(n52619), .Z(n52600) );
  AND U52514 ( .A(n52620), .B(n52621), .Z(n52619) );
  XOR U52515 ( .A(n52622), .B(n52618), .Z(n52620) );
  XNOR U52516 ( .A(n52623), .B(n52624), .Z(n52617) );
  AND U52517 ( .A(n52625), .B(n52626), .Z(n52624) );
  XOR U52518 ( .A(n52623), .B(n52627), .Z(n52625) );
  XNOR U52519 ( .A(n52606), .B(n52603), .Z(n52616) );
  AND U52520 ( .A(n52628), .B(n52629), .Z(n52603) );
  XOR U52521 ( .A(n52630), .B(n52631), .Z(n52606) );
  AND U52522 ( .A(n52632), .B(n52633), .Z(n52631) );
  XOR U52523 ( .A(n52630), .B(n52634), .Z(n52632) );
  XNOR U52524 ( .A(n52567), .B(n52612), .Z(n52614) );
  XNOR U52525 ( .A(n52635), .B(n52636), .Z(n52567) );
  AND U52526 ( .A(n2051), .B(n52637), .Z(n52636) );
  XNOR U52527 ( .A(n52638), .B(n52639), .Z(n52637) );
  XOR U52528 ( .A(n52640), .B(n52641), .Z(n52612) );
  AND U52529 ( .A(n52642), .B(n52643), .Z(n52641) );
  XNOR U52530 ( .A(n52640), .B(n52628), .Z(n52643) );
  IV U52531 ( .A(n52578), .Z(n52628) );
  XNOR U52532 ( .A(n52644), .B(n52621), .Z(n52578) );
  XNOR U52533 ( .A(n52645), .B(n52627), .Z(n52621) );
  XNOR U52534 ( .A(n52646), .B(n52647), .Z(n52627) );
  NOR U52535 ( .A(n52648), .B(n52649), .Z(n52647) );
  XOR U52536 ( .A(n52646), .B(n52650), .Z(n52648) );
  XNOR U52537 ( .A(n52626), .B(n52618), .Z(n52645) );
  XOR U52538 ( .A(n52651), .B(n52652), .Z(n52618) );
  AND U52539 ( .A(n52653), .B(n52654), .Z(n52652) );
  XOR U52540 ( .A(n52651), .B(n52655), .Z(n52653) );
  XNOR U52541 ( .A(n52656), .B(n52623), .Z(n52626) );
  XOR U52542 ( .A(n52657), .B(n52658), .Z(n52623) );
  AND U52543 ( .A(n52659), .B(n52660), .Z(n52658) );
  XNOR U52544 ( .A(n52661), .B(n52662), .Z(n52659) );
  IV U52545 ( .A(n52657), .Z(n52661) );
  XNOR U52546 ( .A(n52663), .B(n52664), .Z(n52656) );
  NOR U52547 ( .A(n52665), .B(n52666), .Z(n52664) );
  XNOR U52548 ( .A(n52663), .B(n52667), .Z(n52665) );
  XNOR U52549 ( .A(n52622), .B(n52629), .Z(n52644) );
  NOR U52550 ( .A(n52584), .B(n52668), .Z(n52629) );
  XOR U52551 ( .A(n52634), .B(n52633), .Z(n52622) );
  XNOR U52552 ( .A(n52669), .B(n52630), .Z(n52633) );
  XOR U52553 ( .A(n52670), .B(n52671), .Z(n52630) );
  AND U52554 ( .A(n52672), .B(n52673), .Z(n52671) );
  XNOR U52555 ( .A(n52674), .B(n52675), .Z(n52672) );
  IV U52556 ( .A(n52670), .Z(n52674) );
  XNOR U52557 ( .A(n52676), .B(n52677), .Z(n52669) );
  NOR U52558 ( .A(n52678), .B(n52679), .Z(n52677) );
  XNOR U52559 ( .A(n52676), .B(n52680), .Z(n52678) );
  XOR U52560 ( .A(n52681), .B(n52682), .Z(n52634) );
  NOR U52561 ( .A(n52683), .B(n52684), .Z(n52682) );
  XNOR U52562 ( .A(n52681), .B(n52685), .Z(n52683) );
  XNOR U52563 ( .A(n52575), .B(n52640), .Z(n52642) );
  XNOR U52564 ( .A(n52686), .B(n52687), .Z(n52575) );
  AND U52565 ( .A(n2051), .B(n52688), .Z(n52687) );
  XNOR U52566 ( .A(n52689), .B(n52690), .Z(n52688) );
  AND U52567 ( .A(n52581), .B(n52584), .Z(n52640) );
  XOR U52568 ( .A(n52691), .B(n52668), .Z(n52584) );
  XNOR U52569 ( .A(p_input[1664]), .B(p_input[2048]), .Z(n52668) );
  XNOR U52570 ( .A(n52655), .B(n52654), .Z(n52691) );
  XNOR U52571 ( .A(n52692), .B(n52662), .Z(n52654) );
  XNOR U52572 ( .A(n52650), .B(n52649), .Z(n52662) );
  XNOR U52573 ( .A(n52693), .B(n52646), .Z(n52649) );
  XNOR U52574 ( .A(p_input[1674]), .B(p_input[2058]), .Z(n52646) );
  XOR U52575 ( .A(p_input[1675]), .B(n29030), .Z(n52693) );
  XOR U52576 ( .A(p_input[1676]), .B(p_input[2060]), .Z(n52650) );
  XOR U52577 ( .A(n52660), .B(n52694), .Z(n52692) );
  IV U52578 ( .A(n52651), .Z(n52694) );
  XOR U52579 ( .A(p_input[1665]), .B(p_input[2049]), .Z(n52651) );
  XNOR U52580 ( .A(n52695), .B(n52667), .Z(n52660) );
  XNOR U52581 ( .A(p_input[1679]), .B(n29033), .Z(n52667) );
  XOR U52582 ( .A(n52657), .B(n52666), .Z(n52695) );
  XOR U52583 ( .A(n52696), .B(n52663), .Z(n52666) );
  XOR U52584 ( .A(p_input[1677]), .B(p_input[2061]), .Z(n52663) );
  XOR U52585 ( .A(p_input[1678]), .B(n29035), .Z(n52696) );
  XOR U52586 ( .A(p_input[1673]), .B(p_input[2057]), .Z(n52657) );
  XOR U52587 ( .A(n52675), .B(n52673), .Z(n52655) );
  XNOR U52588 ( .A(n52697), .B(n52680), .Z(n52673) );
  XOR U52589 ( .A(p_input[1672]), .B(p_input[2056]), .Z(n52680) );
  XOR U52590 ( .A(n52670), .B(n52679), .Z(n52697) );
  XOR U52591 ( .A(n52698), .B(n52676), .Z(n52679) );
  XOR U52592 ( .A(p_input[1670]), .B(p_input[2054]), .Z(n52676) );
  XOR U52593 ( .A(p_input[1671]), .B(n30404), .Z(n52698) );
  XOR U52594 ( .A(p_input[1666]), .B(p_input[2050]), .Z(n52670) );
  XNOR U52595 ( .A(n52685), .B(n52684), .Z(n52675) );
  XOR U52596 ( .A(n52699), .B(n52681), .Z(n52684) );
  XOR U52597 ( .A(p_input[1667]), .B(p_input[2051]), .Z(n52681) );
  XOR U52598 ( .A(p_input[1668]), .B(n30406), .Z(n52699) );
  XOR U52599 ( .A(p_input[1669]), .B(p_input[2053]), .Z(n52685) );
  XNOR U52600 ( .A(n52700), .B(n52701), .Z(n52581) );
  AND U52601 ( .A(n2051), .B(n52702), .Z(n52701) );
  XNOR U52602 ( .A(n52703), .B(n52704), .Z(n2051) );
  AND U52603 ( .A(n52705), .B(n52706), .Z(n52704) );
  XOR U52604 ( .A(n52595), .B(n52703), .Z(n52706) );
  XNOR U52605 ( .A(n52707), .B(n52703), .Z(n52705) );
  XOR U52606 ( .A(n52708), .B(n52709), .Z(n52703) );
  AND U52607 ( .A(n52710), .B(n52711), .Z(n52709) );
  XOR U52608 ( .A(n52610), .B(n52708), .Z(n52711) );
  XOR U52609 ( .A(n52708), .B(n52611), .Z(n52710) );
  XOR U52610 ( .A(n52712), .B(n52713), .Z(n52708) );
  AND U52611 ( .A(n52714), .B(n52715), .Z(n52713) );
  XOR U52612 ( .A(n52638), .B(n52712), .Z(n52715) );
  XOR U52613 ( .A(n52712), .B(n52639), .Z(n52714) );
  XOR U52614 ( .A(n52716), .B(n52717), .Z(n52712) );
  AND U52615 ( .A(n52718), .B(n52719), .Z(n52717) );
  XOR U52616 ( .A(n52716), .B(n52689), .Z(n52719) );
  XNOR U52617 ( .A(n52720), .B(n52721), .Z(n52541) );
  AND U52618 ( .A(n2055), .B(n52722), .Z(n52721) );
  XNOR U52619 ( .A(n52723), .B(n52724), .Z(n2055) );
  AND U52620 ( .A(n52725), .B(n52726), .Z(n52724) );
  XOR U52621 ( .A(n52723), .B(n52551), .Z(n52726) );
  XNOR U52622 ( .A(n52723), .B(n52511), .Z(n52725) );
  XOR U52623 ( .A(n52727), .B(n52728), .Z(n52723) );
  AND U52624 ( .A(n52729), .B(n52730), .Z(n52728) );
  XOR U52625 ( .A(n52727), .B(n52519), .Z(n52729) );
  XOR U52626 ( .A(n52731), .B(n52732), .Z(n52502) );
  AND U52627 ( .A(n2059), .B(n52722), .Z(n52732) );
  XNOR U52628 ( .A(n52720), .B(n52731), .Z(n52722) );
  XNOR U52629 ( .A(n52733), .B(n52734), .Z(n2059) );
  AND U52630 ( .A(n52735), .B(n52736), .Z(n52734) );
  XNOR U52631 ( .A(n52737), .B(n52733), .Z(n52736) );
  IV U52632 ( .A(n52551), .Z(n52737) );
  XOR U52633 ( .A(n52707), .B(n52738), .Z(n52551) );
  AND U52634 ( .A(n2062), .B(n52739), .Z(n52738) );
  XOR U52635 ( .A(n52594), .B(n52591), .Z(n52739) );
  IV U52636 ( .A(n52707), .Z(n52594) );
  XNOR U52637 ( .A(n52511), .B(n52733), .Z(n52735) );
  XOR U52638 ( .A(n52740), .B(n52741), .Z(n52511) );
  AND U52639 ( .A(n2078), .B(n52742), .Z(n52741) );
  XOR U52640 ( .A(n52727), .B(n52743), .Z(n52733) );
  AND U52641 ( .A(n52744), .B(n52730), .Z(n52743) );
  XNOR U52642 ( .A(n52561), .B(n52727), .Z(n52730) );
  XOR U52643 ( .A(n52611), .B(n52745), .Z(n52561) );
  AND U52644 ( .A(n2062), .B(n52746), .Z(n52745) );
  XOR U52645 ( .A(n52607), .B(n52611), .Z(n52746) );
  XNOR U52646 ( .A(n52747), .B(n52727), .Z(n52744) );
  IV U52647 ( .A(n52519), .Z(n52747) );
  XOR U52648 ( .A(n52748), .B(n52749), .Z(n52519) );
  AND U52649 ( .A(n2078), .B(n52750), .Z(n52749) );
  XOR U52650 ( .A(n52751), .B(n52752), .Z(n52727) );
  AND U52651 ( .A(n52753), .B(n52754), .Z(n52752) );
  XNOR U52652 ( .A(n52571), .B(n52751), .Z(n52754) );
  XOR U52653 ( .A(n52639), .B(n52755), .Z(n52571) );
  AND U52654 ( .A(n2062), .B(n52756), .Z(n52755) );
  XOR U52655 ( .A(n52635), .B(n52639), .Z(n52756) );
  XOR U52656 ( .A(n52751), .B(n52528), .Z(n52753) );
  XOR U52657 ( .A(n52757), .B(n52758), .Z(n52528) );
  AND U52658 ( .A(n2078), .B(n52759), .Z(n52758) );
  XOR U52659 ( .A(n52760), .B(n52761), .Z(n52751) );
  AND U52660 ( .A(n52762), .B(n52763), .Z(n52761) );
  XNOR U52661 ( .A(n52760), .B(n52579), .Z(n52763) );
  XOR U52662 ( .A(n52690), .B(n52764), .Z(n52579) );
  AND U52663 ( .A(n2062), .B(n52765), .Z(n52764) );
  XOR U52664 ( .A(n52686), .B(n52690), .Z(n52765) );
  XNOR U52665 ( .A(n52766), .B(n52760), .Z(n52762) );
  IV U52666 ( .A(n52538), .Z(n52766) );
  XOR U52667 ( .A(n52767), .B(n52768), .Z(n52538) );
  AND U52668 ( .A(n2078), .B(n52769), .Z(n52768) );
  AND U52669 ( .A(n52731), .B(n52720), .Z(n52760) );
  XNOR U52670 ( .A(n52770), .B(n52771), .Z(n52720) );
  AND U52671 ( .A(n2062), .B(n52702), .Z(n52771) );
  XNOR U52672 ( .A(n52700), .B(n52770), .Z(n52702) );
  XNOR U52673 ( .A(n52772), .B(n52773), .Z(n2062) );
  AND U52674 ( .A(n52774), .B(n52775), .Z(n52773) );
  XNOR U52675 ( .A(n52772), .B(n52591), .Z(n52775) );
  IV U52676 ( .A(n52595), .Z(n52591) );
  XOR U52677 ( .A(n52776), .B(n52777), .Z(n52595) );
  AND U52678 ( .A(n2066), .B(n52778), .Z(n52777) );
  XOR U52679 ( .A(n52779), .B(n52776), .Z(n52778) );
  XNOR U52680 ( .A(n52772), .B(n52707), .Z(n52774) );
  XOR U52681 ( .A(n52780), .B(n52781), .Z(n52707) );
  AND U52682 ( .A(n2074), .B(n52742), .Z(n52781) );
  XOR U52683 ( .A(n52740), .B(n52780), .Z(n52742) );
  XOR U52684 ( .A(n52782), .B(n52783), .Z(n52772) );
  AND U52685 ( .A(n52784), .B(n52785), .Z(n52783) );
  XNOR U52686 ( .A(n52782), .B(n52607), .Z(n52785) );
  IV U52687 ( .A(n52610), .Z(n52607) );
  XOR U52688 ( .A(n52786), .B(n52787), .Z(n52610) );
  AND U52689 ( .A(n2066), .B(n52788), .Z(n52787) );
  XOR U52690 ( .A(n52789), .B(n52786), .Z(n52788) );
  XOR U52691 ( .A(n52611), .B(n52782), .Z(n52784) );
  XOR U52692 ( .A(n52790), .B(n52791), .Z(n52611) );
  AND U52693 ( .A(n2074), .B(n52750), .Z(n52791) );
  XOR U52694 ( .A(n52790), .B(n52748), .Z(n52750) );
  XOR U52695 ( .A(n52792), .B(n52793), .Z(n52782) );
  AND U52696 ( .A(n52794), .B(n52795), .Z(n52793) );
  XNOR U52697 ( .A(n52792), .B(n52635), .Z(n52795) );
  IV U52698 ( .A(n52638), .Z(n52635) );
  XOR U52699 ( .A(n52796), .B(n52797), .Z(n52638) );
  AND U52700 ( .A(n2066), .B(n52798), .Z(n52797) );
  XNOR U52701 ( .A(n52799), .B(n52796), .Z(n52798) );
  XOR U52702 ( .A(n52639), .B(n52792), .Z(n52794) );
  XOR U52703 ( .A(n52800), .B(n52801), .Z(n52639) );
  AND U52704 ( .A(n2074), .B(n52759), .Z(n52801) );
  XOR U52705 ( .A(n52800), .B(n52757), .Z(n52759) );
  XOR U52706 ( .A(n52716), .B(n52802), .Z(n52792) );
  AND U52707 ( .A(n52718), .B(n52803), .Z(n52802) );
  XNOR U52708 ( .A(n52716), .B(n52686), .Z(n52803) );
  IV U52709 ( .A(n52689), .Z(n52686) );
  XOR U52710 ( .A(n52804), .B(n52805), .Z(n52689) );
  AND U52711 ( .A(n2066), .B(n52806), .Z(n52805) );
  XOR U52712 ( .A(n52807), .B(n52804), .Z(n52806) );
  XOR U52713 ( .A(n52690), .B(n52716), .Z(n52718) );
  XOR U52714 ( .A(n52808), .B(n52809), .Z(n52690) );
  AND U52715 ( .A(n2074), .B(n52769), .Z(n52809) );
  XOR U52716 ( .A(n52808), .B(n52767), .Z(n52769) );
  AND U52717 ( .A(n52770), .B(n52700), .Z(n52716) );
  XNOR U52718 ( .A(n52810), .B(n52811), .Z(n52700) );
  AND U52719 ( .A(n2066), .B(n52812), .Z(n52811) );
  XNOR U52720 ( .A(n52813), .B(n52810), .Z(n52812) );
  XNOR U52721 ( .A(n52814), .B(n52815), .Z(n2066) );
  AND U52722 ( .A(n52816), .B(n52817), .Z(n52815) );
  XOR U52723 ( .A(n52779), .B(n52814), .Z(n52817) );
  AND U52724 ( .A(n52818), .B(n52819), .Z(n52779) );
  XNOR U52725 ( .A(n52776), .B(n52814), .Z(n52816) );
  XNOR U52726 ( .A(n52820), .B(n52821), .Z(n52776) );
  AND U52727 ( .A(n2070), .B(n52822), .Z(n52821) );
  XNOR U52728 ( .A(n52823), .B(n52824), .Z(n52822) );
  XOR U52729 ( .A(n52825), .B(n52826), .Z(n52814) );
  AND U52730 ( .A(n52827), .B(n52828), .Z(n52826) );
  XNOR U52731 ( .A(n52825), .B(n52818), .Z(n52828) );
  IV U52732 ( .A(n52789), .Z(n52818) );
  XOR U52733 ( .A(n52829), .B(n52830), .Z(n52789) );
  XOR U52734 ( .A(n52831), .B(n52819), .Z(n52830) );
  AND U52735 ( .A(n52799), .B(n52832), .Z(n52819) );
  AND U52736 ( .A(n52833), .B(n52834), .Z(n52831) );
  XOR U52737 ( .A(n52835), .B(n52829), .Z(n52833) );
  XNOR U52738 ( .A(n52786), .B(n52825), .Z(n52827) );
  XNOR U52739 ( .A(n52836), .B(n52837), .Z(n52786) );
  AND U52740 ( .A(n2070), .B(n52838), .Z(n52837) );
  XNOR U52741 ( .A(n52839), .B(n52840), .Z(n52838) );
  XOR U52742 ( .A(n52841), .B(n52842), .Z(n52825) );
  AND U52743 ( .A(n52843), .B(n52844), .Z(n52842) );
  XNOR U52744 ( .A(n52841), .B(n52799), .Z(n52844) );
  XOR U52745 ( .A(n52845), .B(n52834), .Z(n52799) );
  XNOR U52746 ( .A(n52846), .B(n52829), .Z(n52834) );
  XOR U52747 ( .A(n52847), .B(n52848), .Z(n52829) );
  AND U52748 ( .A(n52849), .B(n52850), .Z(n52848) );
  XOR U52749 ( .A(n52851), .B(n52847), .Z(n52849) );
  XNOR U52750 ( .A(n52852), .B(n52853), .Z(n52846) );
  AND U52751 ( .A(n52854), .B(n52855), .Z(n52853) );
  XOR U52752 ( .A(n52852), .B(n52856), .Z(n52854) );
  XNOR U52753 ( .A(n52835), .B(n52832), .Z(n52845) );
  AND U52754 ( .A(n52857), .B(n52858), .Z(n52832) );
  XOR U52755 ( .A(n52859), .B(n52860), .Z(n52835) );
  AND U52756 ( .A(n52861), .B(n52862), .Z(n52860) );
  XOR U52757 ( .A(n52859), .B(n52863), .Z(n52861) );
  XNOR U52758 ( .A(n52796), .B(n52841), .Z(n52843) );
  XNOR U52759 ( .A(n52864), .B(n52865), .Z(n52796) );
  AND U52760 ( .A(n2070), .B(n52866), .Z(n52865) );
  XNOR U52761 ( .A(n52867), .B(n52868), .Z(n52866) );
  XOR U52762 ( .A(n52869), .B(n52870), .Z(n52841) );
  AND U52763 ( .A(n52871), .B(n52872), .Z(n52870) );
  XNOR U52764 ( .A(n52869), .B(n52857), .Z(n52872) );
  IV U52765 ( .A(n52807), .Z(n52857) );
  XNOR U52766 ( .A(n52873), .B(n52850), .Z(n52807) );
  XNOR U52767 ( .A(n52874), .B(n52856), .Z(n52850) );
  XNOR U52768 ( .A(n52875), .B(n52876), .Z(n52856) );
  NOR U52769 ( .A(n52877), .B(n52878), .Z(n52876) );
  XOR U52770 ( .A(n52875), .B(n52879), .Z(n52877) );
  XNOR U52771 ( .A(n52855), .B(n52847), .Z(n52874) );
  XOR U52772 ( .A(n52880), .B(n52881), .Z(n52847) );
  AND U52773 ( .A(n52882), .B(n52883), .Z(n52881) );
  XOR U52774 ( .A(n52880), .B(n52884), .Z(n52882) );
  XNOR U52775 ( .A(n52885), .B(n52852), .Z(n52855) );
  XOR U52776 ( .A(n52886), .B(n52887), .Z(n52852) );
  AND U52777 ( .A(n52888), .B(n52889), .Z(n52887) );
  XNOR U52778 ( .A(n52890), .B(n52891), .Z(n52888) );
  IV U52779 ( .A(n52886), .Z(n52890) );
  XNOR U52780 ( .A(n52892), .B(n52893), .Z(n52885) );
  NOR U52781 ( .A(n52894), .B(n52895), .Z(n52893) );
  XNOR U52782 ( .A(n52892), .B(n52896), .Z(n52894) );
  XNOR U52783 ( .A(n52851), .B(n52858), .Z(n52873) );
  NOR U52784 ( .A(n52813), .B(n52897), .Z(n52858) );
  XOR U52785 ( .A(n52863), .B(n52862), .Z(n52851) );
  XNOR U52786 ( .A(n52898), .B(n52859), .Z(n52862) );
  XOR U52787 ( .A(n52899), .B(n52900), .Z(n52859) );
  AND U52788 ( .A(n52901), .B(n52902), .Z(n52900) );
  XNOR U52789 ( .A(n52903), .B(n52904), .Z(n52901) );
  IV U52790 ( .A(n52899), .Z(n52903) );
  XNOR U52791 ( .A(n52905), .B(n52906), .Z(n52898) );
  NOR U52792 ( .A(n52907), .B(n52908), .Z(n52906) );
  XNOR U52793 ( .A(n52905), .B(n52909), .Z(n52907) );
  XOR U52794 ( .A(n52910), .B(n52911), .Z(n52863) );
  NOR U52795 ( .A(n52912), .B(n52913), .Z(n52911) );
  XNOR U52796 ( .A(n52910), .B(n52914), .Z(n52912) );
  XNOR U52797 ( .A(n52804), .B(n52869), .Z(n52871) );
  XNOR U52798 ( .A(n52915), .B(n52916), .Z(n52804) );
  AND U52799 ( .A(n2070), .B(n52917), .Z(n52916) );
  XNOR U52800 ( .A(n52918), .B(n52919), .Z(n52917) );
  AND U52801 ( .A(n52810), .B(n52813), .Z(n52869) );
  XOR U52802 ( .A(n52920), .B(n52897), .Z(n52813) );
  XNOR U52803 ( .A(p_input[1680]), .B(p_input[2048]), .Z(n52897) );
  XNOR U52804 ( .A(n52884), .B(n52883), .Z(n52920) );
  XNOR U52805 ( .A(n52921), .B(n52891), .Z(n52883) );
  XNOR U52806 ( .A(n52879), .B(n52878), .Z(n52891) );
  XNOR U52807 ( .A(n52922), .B(n52875), .Z(n52878) );
  XNOR U52808 ( .A(p_input[1690]), .B(p_input[2058]), .Z(n52875) );
  XOR U52809 ( .A(p_input[1691]), .B(n29030), .Z(n52922) );
  XOR U52810 ( .A(p_input[1692]), .B(p_input[2060]), .Z(n52879) );
  XOR U52811 ( .A(n52889), .B(n52923), .Z(n52921) );
  IV U52812 ( .A(n52880), .Z(n52923) );
  XOR U52813 ( .A(p_input[1681]), .B(p_input[2049]), .Z(n52880) );
  XNOR U52814 ( .A(n52924), .B(n52896), .Z(n52889) );
  XNOR U52815 ( .A(p_input[1695]), .B(n29033), .Z(n52896) );
  XOR U52816 ( .A(n52886), .B(n52895), .Z(n52924) );
  XOR U52817 ( .A(n52925), .B(n52892), .Z(n52895) );
  XOR U52818 ( .A(p_input[1693]), .B(p_input[2061]), .Z(n52892) );
  XOR U52819 ( .A(p_input[1694]), .B(n29035), .Z(n52925) );
  XOR U52820 ( .A(p_input[1689]), .B(p_input[2057]), .Z(n52886) );
  XOR U52821 ( .A(n52904), .B(n52902), .Z(n52884) );
  XNOR U52822 ( .A(n52926), .B(n52909), .Z(n52902) );
  XOR U52823 ( .A(p_input[1688]), .B(p_input[2056]), .Z(n52909) );
  XOR U52824 ( .A(n52899), .B(n52908), .Z(n52926) );
  XOR U52825 ( .A(n52927), .B(n52905), .Z(n52908) );
  XOR U52826 ( .A(p_input[1686]), .B(p_input[2054]), .Z(n52905) );
  XOR U52827 ( .A(p_input[1687]), .B(n30404), .Z(n52927) );
  XOR U52828 ( .A(p_input[1682]), .B(p_input[2050]), .Z(n52899) );
  XNOR U52829 ( .A(n52914), .B(n52913), .Z(n52904) );
  XOR U52830 ( .A(n52928), .B(n52910), .Z(n52913) );
  XOR U52831 ( .A(p_input[1683]), .B(p_input[2051]), .Z(n52910) );
  XOR U52832 ( .A(p_input[1684]), .B(n30406), .Z(n52928) );
  XOR U52833 ( .A(p_input[1685]), .B(p_input[2053]), .Z(n52914) );
  XNOR U52834 ( .A(n52929), .B(n52930), .Z(n52810) );
  AND U52835 ( .A(n2070), .B(n52931), .Z(n52930) );
  XNOR U52836 ( .A(n52932), .B(n52933), .Z(n2070) );
  AND U52837 ( .A(n52934), .B(n52935), .Z(n52933) );
  XOR U52838 ( .A(n52824), .B(n52932), .Z(n52935) );
  XNOR U52839 ( .A(n52936), .B(n52932), .Z(n52934) );
  XOR U52840 ( .A(n52937), .B(n52938), .Z(n52932) );
  AND U52841 ( .A(n52939), .B(n52940), .Z(n52938) );
  XOR U52842 ( .A(n52839), .B(n52937), .Z(n52940) );
  XOR U52843 ( .A(n52937), .B(n52840), .Z(n52939) );
  XOR U52844 ( .A(n52941), .B(n52942), .Z(n52937) );
  AND U52845 ( .A(n52943), .B(n52944), .Z(n52942) );
  XOR U52846 ( .A(n52867), .B(n52941), .Z(n52944) );
  XOR U52847 ( .A(n52941), .B(n52868), .Z(n52943) );
  XOR U52848 ( .A(n52945), .B(n52946), .Z(n52941) );
  AND U52849 ( .A(n52947), .B(n52948), .Z(n52946) );
  XOR U52850 ( .A(n52945), .B(n52918), .Z(n52948) );
  XNOR U52851 ( .A(n52949), .B(n52950), .Z(n52770) );
  AND U52852 ( .A(n2074), .B(n52951), .Z(n52950) );
  XNOR U52853 ( .A(n52952), .B(n52953), .Z(n2074) );
  AND U52854 ( .A(n52954), .B(n52955), .Z(n52953) );
  XOR U52855 ( .A(n52952), .B(n52780), .Z(n52955) );
  XNOR U52856 ( .A(n52952), .B(n52740), .Z(n52954) );
  XOR U52857 ( .A(n52956), .B(n52957), .Z(n52952) );
  AND U52858 ( .A(n52958), .B(n52959), .Z(n52957) );
  XOR U52859 ( .A(n52956), .B(n52748), .Z(n52958) );
  XOR U52860 ( .A(n52960), .B(n52961), .Z(n52731) );
  AND U52861 ( .A(n2078), .B(n52951), .Z(n52961) );
  XNOR U52862 ( .A(n52949), .B(n52960), .Z(n52951) );
  XNOR U52863 ( .A(n52962), .B(n52963), .Z(n2078) );
  AND U52864 ( .A(n52964), .B(n52965), .Z(n52963) );
  XNOR U52865 ( .A(n52966), .B(n52962), .Z(n52965) );
  IV U52866 ( .A(n52780), .Z(n52966) );
  XOR U52867 ( .A(n52936), .B(n52967), .Z(n52780) );
  AND U52868 ( .A(n2081), .B(n52968), .Z(n52967) );
  XOR U52869 ( .A(n52823), .B(n52820), .Z(n52968) );
  IV U52870 ( .A(n52936), .Z(n52823) );
  XNOR U52871 ( .A(n52740), .B(n52962), .Z(n52964) );
  XOR U52872 ( .A(n52969), .B(n52970), .Z(n52740) );
  AND U52873 ( .A(n2097), .B(n52971), .Z(n52970) );
  XOR U52874 ( .A(n52956), .B(n52972), .Z(n52962) );
  AND U52875 ( .A(n52973), .B(n52959), .Z(n52972) );
  XNOR U52876 ( .A(n52790), .B(n52956), .Z(n52959) );
  XOR U52877 ( .A(n52840), .B(n52974), .Z(n52790) );
  AND U52878 ( .A(n2081), .B(n52975), .Z(n52974) );
  XOR U52879 ( .A(n52836), .B(n52840), .Z(n52975) );
  XNOR U52880 ( .A(n52976), .B(n52956), .Z(n52973) );
  IV U52881 ( .A(n52748), .Z(n52976) );
  XOR U52882 ( .A(n52977), .B(n52978), .Z(n52748) );
  AND U52883 ( .A(n2097), .B(n52979), .Z(n52978) );
  XOR U52884 ( .A(n52980), .B(n52981), .Z(n52956) );
  AND U52885 ( .A(n52982), .B(n52983), .Z(n52981) );
  XNOR U52886 ( .A(n52800), .B(n52980), .Z(n52983) );
  XOR U52887 ( .A(n52868), .B(n52984), .Z(n52800) );
  AND U52888 ( .A(n2081), .B(n52985), .Z(n52984) );
  XOR U52889 ( .A(n52864), .B(n52868), .Z(n52985) );
  XOR U52890 ( .A(n52980), .B(n52757), .Z(n52982) );
  XOR U52891 ( .A(n52986), .B(n52987), .Z(n52757) );
  AND U52892 ( .A(n2097), .B(n52988), .Z(n52987) );
  XOR U52893 ( .A(n52989), .B(n52990), .Z(n52980) );
  AND U52894 ( .A(n52991), .B(n52992), .Z(n52990) );
  XNOR U52895 ( .A(n52989), .B(n52808), .Z(n52992) );
  XOR U52896 ( .A(n52919), .B(n52993), .Z(n52808) );
  AND U52897 ( .A(n2081), .B(n52994), .Z(n52993) );
  XOR U52898 ( .A(n52915), .B(n52919), .Z(n52994) );
  XNOR U52899 ( .A(n52995), .B(n52989), .Z(n52991) );
  IV U52900 ( .A(n52767), .Z(n52995) );
  XOR U52901 ( .A(n52996), .B(n52997), .Z(n52767) );
  AND U52902 ( .A(n2097), .B(n52998), .Z(n52997) );
  AND U52903 ( .A(n52960), .B(n52949), .Z(n52989) );
  XNOR U52904 ( .A(n52999), .B(n53000), .Z(n52949) );
  AND U52905 ( .A(n2081), .B(n52931), .Z(n53000) );
  XNOR U52906 ( .A(n52929), .B(n52999), .Z(n52931) );
  XNOR U52907 ( .A(n53001), .B(n53002), .Z(n2081) );
  AND U52908 ( .A(n53003), .B(n53004), .Z(n53002) );
  XNOR U52909 ( .A(n53001), .B(n52820), .Z(n53004) );
  IV U52910 ( .A(n52824), .Z(n52820) );
  XOR U52911 ( .A(n53005), .B(n53006), .Z(n52824) );
  AND U52912 ( .A(n2085), .B(n53007), .Z(n53006) );
  XOR U52913 ( .A(n53008), .B(n53005), .Z(n53007) );
  XNOR U52914 ( .A(n53001), .B(n52936), .Z(n53003) );
  XOR U52915 ( .A(n53009), .B(n53010), .Z(n52936) );
  AND U52916 ( .A(n2093), .B(n52971), .Z(n53010) );
  XOR U52917 ( .A(n52969), .B(n53009), .Z(n52971) );
  XOR U52918 ( .A(n53011), .B(n53012), .Z(n53001) );
  AND U52919 ( .A(n53013), .B(n53014), .Z(n53012) );
  XNOR U52920 ( .A(n53011), .B(n52836), .Z(n53014) );
  IV U52921 ( .A(n52839), .Z(n52836) );
  XOR U52922 ( .A(n53015), .B(n53016), .Z(n52839) );
  AND U52923 ( .A(n2085), .B(n53017), .Z(n53016) );
  XOR U52924 ( .A(n53018), .B(n53015), .Z(n53017) );
  XOR U52925 ( .A(n52840), .B(n53011), .Z(n53013) );
  XOR U52926 ( .A(n53019), .B(n53020), .Z(n52840) );
  AND U52927 ( .A(n2093), .B(n52979), .Z(n53020) );
  XOR U52928 ( .A(n53019), .B(n52977), .Z(n52979) );
  XOR U52929 ( .A(n53021), .B(n53022), .Z(n53011) );
  AND U52930 ( .A(n53023), .B(n53024), .Z(n53022) );
  XNOR U52931 ( .A(n53021), .B(n52864), .Z(n53024) );
  IV U52932 ( .A(n52867), .Z(n52864) );
  XOR U52933 ( .A(n53025), .B(n53026), .Z(n52867) );
  AND U52934 ( .A(n2085), .B(n53027), .Z(n53026) );
  XNOR U52935 ( .A(n53028), .B(n53025), .Z(n53027) );
  XOR U52936 ( .A(n52868), .B(n53021), .Z(n53023) );
  XOR U52937 ( .A(n53029), .B(n53030), .Z(n52868) );
  AND U52938 ( .A(n2093), .B(n52988), .Z(n53030) );
  XOR U52939 ( .A(n53029), .B(n52986), .Z(n52988) );
  XOR U52940 ( .A(n52945), .B(n53031), .Z(n53021) );
  AND U52941 ( .A(n52947), .B(n53032), .Z(n53031) );
  XNOR U52942 ( .A(n52945), .B(n52915), .Z(n53032) );
  IV U52943 ( .A(n52918), .Z(n52915) );
  XOR U52944 ( .A(n53033), .B(n53034), .Z(n52918) );
  AND U52945 ( .A(n2085), .B(n53035), .Z(n53034) );
  XOR U52946 ( .A(n53036), .B(n53033), .Z(n53035) );
  XOR U52947 ( .A(n52919), .B(n52945), .Z(n52947) );
  XOR U52948 ( .A(n53037), .B(n53038), .Z(n52919) );
  AND U52949 ( .A(n2093), .B(n52998), .Z(n53038) );
  XOR U52950 ( .A(n53037), .B(n52996), .Z(n52998) );
  AND U52951 ( .A(n52999), .B(n52929), .Z(n52945) );
  XNOR U52952 ( .A(n53039), .B(n53040), .Z(n52929) );
  AND U52953 ( .A(n2085), .B(n53041), .Z(n53040) );
  XNOR U52954 ( .A(n53042), .B(n53039), .Z(n53041) );
  XNOR U52955 ( .A(n53043), .B(n53044), .Z(n2085) );
  AND U52956 ( .A(n53045), .B(n53046), .Z(n53044) );
  XOR U52957 ( .A(n53008), .B(n53043), .Z(n53046) );
  AND U52958 ( .A(n53047), .B(n53048), .Z(n53008) );
  XNOR U52959 ( .A(n53005), .B(n53043), .Z(n53045) );
  XNOR U52960 ( .A(n53049), .B(n53050), .Z(n53005) );
  AND U52961 ( .A(n2089), .B(n53051), .Z(n53050) );
  XNOR U52962 ( .A(n53052), .B(n53053), .Z(n53051) );
  XOR U52963 ( .A(n53054), .B(n53055), .Z(n53043) );
  AND U52964 ( .A(n53056), .B(n53057), .Z(n53055) );
  XNOR U52965 ( .A(n53054), .B(n53047), .Z(n53057) );
  IV U52966 ( .A(n53018), .Z(n53047) );
  XOR U52967 ( .A(n53058), .B(n53059), .Z(n53018) );
  XOR U52968 ( .A(n53060), .B(n53048), .Z(n53059) );
  AND U52969 ( .A(n53028), .B(n53061), .Z(n53048) );
  AND U52970 ( .A(n53062), .B(n53063), .Z(n53060) );
  XOR U52971 ( .A(n53064), .B(n53058), .Z(n53062) );
  XNOR U52972 ( .A(n53015), .B(n53054), .Z(n53056) );
  XNOR U52973 ( .A(n53065), .B(n53066), .Z(n53015) );
  AND U52974 ( .A(n2089), .B(n53067), .Z(n53066) );
  XNOR U52975 ( .A(n53068), .B(n53069), .Z(n53067) );
  XOR U52976 ( .A(n53070), .B(n53071), .Z(n53054) );
  AND U52977 ( .A(n53072), .B(n53073), .Z(n53071) );
  XNOR U52978 ( .A(n53070), .B(n53028), .Z(n53073) );
  XOR U52979 ( .A(n53074), .B(n53063), .Z(n53028) );
  XNOR U52980 ( .A(n53075), .B(n53058), .Z(n53063) );
  XOR U52981 ( .A(n53076), .B(n53077), .Z(n53058) );
  AND U52982 ( .A(n53078), .B(n53079), .Z(n53077) );
  XOR U52983 ( .A(n53080), .B(n53076), .Z(n53078) );
  XNOR U52984 ( .A(n53081), .B(n53082), .Z(n53075) );
  AND U52985 ( .A(n53083), .B(n53084), .Z(n53082) );
  XOR U52986 ( .A(n53081), .B(n53085), .Z(n53083) );
  XNOR U52987 ( .A(n53064), .B(n53061), .Z(n53074) );
  AND U52988 ( .A(n53086), .B(n53087), .Z(n53061) );
  XOR U52989 ( .A(n53088), .B(n53089), .Z(n53064) );
  AND U52990 ( .A(n53090), .B(n53091), .Z(n53089) );
  XOR U52991 ( .A(n53088), .B(n53092), .Z(n53090) );
  XNOR U52992 ( .A(n53025), .B(n53070), .Z(n53072) );
  XNOR U52993 ( .A(n53093), .B(n53094), .Z(n53025) );
  AND U52994 ( .A(n2089), .B(n53095), .Z(n53094) );
  XNOR U52995 ( .A(n53096), .B(n53097), .Z(n53095) );
  XOR U52996 ( .A(n53098), .B(n53099), .Z(n53070) );
  AND U52997 ( .A(n53100), .B(n53101), .Z(n53099) );
  XNOR U52998 ( .A(n53098), .B(n53086), .Z(n53101) );
  IV U52999 ( .A(n53036), .Z(n53086) );
  XNOR U53000 ( .A(n53102), .B(n53079), .Z(n53036) );
  XNOR U53001 ( .A(n53103), .B(n53085), .Z(n53079) );
  XNOR U53002 ( .A(n53104), .B(n53105), .Z(n53085) );
  NOR U53003 ( .A(n53106), .B(n53107), .Z(n53105) );
  XOR U53004 ( .A(n53104), .B(n53108), .Z(n53106) );
  XNOR U53005 ( .A(n53084), .B(n53076), .Z(n53103) );
  XOR U53006 ( .A(n53109), .B(n53110), .Z(n53076) );
  AND U53007 ( .A(n53111), .B(n53112), .Z(n53110) );
  XOR U53008 ( .A(n53109), .B(n53113), .Z(n53111) );
  XNOR U53009 ( .A(n53114), .B(n53081), .Z(n53084) );
  XOR U53010 ( .A(n53115), .B(n53116), .Z(n53081) );
  AND U53011 ( .A(n53117), .B(n53118), .Z(n53116) );
  XNOR U53012 ( .A(n53119), .B(n53120), .Z(n53117) );
  IV U53013 ( .A(n53115), .Z(n53119) );
  XNOR U53014 ( .A(n53121), .B(n53122), .Z(n53114) );
  NOR U53015 ( .A(n53123), .B(n53124), .Z(n53122) );
  XNOR U53016 ( .A(n53121), .B(n53125), .Z(n53123) );
  XNOR U53017 ( .A(n53080), .B(n53087), .Z(n53102) );
  NOR U53018 ( .A(n53042), .B(n53126), .Z(n53087) );
  XOR U53019 ( .A(n53092), .B(n53091), .Z(n53080) );
  XNOR U53020 ( .A(n53127), .B(n53088), .Z(n53091) );
  XOR U53021 ( .A(n53128), .B(n53129), .Z(n53088) );
  AND U53022 ( .A(n53130), .B(n53131), .Z(n53129) );
  XNOR U53023 ( .A(n53132), .B(n53133), .Z(n53130) );
  IV U53024 ( .A(n53128), .Z(n53132) );
  XNOR U53025 ( .A(n53134), .B(n53135), .Z(n53127) );
  NOR U53026 ( .A(n53136), .B(n53137), .Z(n53135) );
  XNOR U53027 ( .A(n53134), .B(n53138), .Z(n53136) );
  XOR U53028 ( .A(n53139), .B(n53140), .Z(n53092) );
  NOR U53029 ( .A(n53141), .B(n53142), .Z(n53140) );
  XNOR U53030 ( .A(n53139), .B(n53143), .Z(n53141) );
  XNOR U53031 ( .A(n53033), .B(n53098), .Z(n53100) );
  XNOR U53032 ( .A(n53144), .B(n53145), .Z(n53033) );
  AND U53033 ( .A(n2089), .B(n53146), .Z(n53145) );
  XNOR U53034 ( .A(n53147), .B(n53148), .Z(n53146) );
  AND U53035 ( .A(n53039), .B(n53042), .Z(n53098) );
  XOR U53036 ( .A(n53149), .B(n53126), .Z(n53042) );
  XNOR U53037 ( .A(p_input[1696]), .B(p_input[2048]), .Z(n53126) );
  XNOR U53038 ( .A(n53113), .B(n53112), .Z(n53149) );
  XNOR U53039 ( .A(n53150), .B(n53120), .Z(n53112) );
  XNOR U53040 ( .A(n53108), .B(n53107), .Z(n53120) );
  XNOR U53041 ( .A(n53151), .B(n53104), .Z(n53107) );
  XNOR U53042 ( .A(p_input[1706]), .B(p_input[2058]), .Z(n53104) );
  XOR U53043 ( .A(p_input[1707]), .B(n29030), .Z(n53151) );
  XOR U53044 ( .A(p_input[1708]), .B(p_input[2060]), .Z(n53108) );
  XOR U53045 ( .A(n53118), .B(n53152), .Z(n53150) );
  IV U53046 ( .A(n53109), .Z(n53152) );
  XOR U53047 ( .A(p_input[1697]), .B(p_input[2049]), .Z(n53109) );
  XNOR U53048 ( .A(n53153), .B(n53125), .Z(n53118) );
  XNOR U53049 ( .A(p_input[1711]), .B(n29033), .Z(n53125) );
  XOR U53050 ( .A(n53115), .B(n53124), .Z(n53153) );
  XOR U53051 ( .A(n53154), .B(n53121), .Z(n53124) );
  XOR U53052 ( .A(p_input[1709]), .B(p_input[2061]), .Z(n53121) );
  XOR U53053 ( .A(p_input[1710]), .B(n29035), .Z(n53154) );
  XOR U53054 ( .A(p_input[1705]), .B(p_input[2057]), .Z(n53115) );
  XOR U53055 ( .A(n53133), .B(n53131), .Z(n53113) );
  XNOR U53056 ( .A(n53155), .B(n53138), .Z(n53131) );
  XOR U53057 ( .A(p_input[1704]), .B(p_input[2056]), .Z(n53138) );
  XOR U53058 ( .A(n53128), .B(n53137), .Z(n53155) );
  XOR U53059 ( .A(n53156), .B(n53134), .Z(n53137) );
  XOR U53060 ( .A(p_input[1702]), .B(p_input[2054]), .Z(n53134) );
  XOR U53061 ( .A(p_input[1703]), .B(n30404), .Z(n53156) );
  XOR U53062 ( .A(p_input[1698]), .B(p_input[2050]), .Z(n53128) );
  XNOR U53063 ( .A(n53143), .B(n53142), .Z(n53133) );
  XOR U53064 ( .A(n53157), .B(n53139), .Z(n53142) );
  XOR U53065 ( .A(p_input[1699]), .B(p_input[2051]), .Z(n53139) );
  XOR U53066 ( .A(p_input[1700]), .B(n30406), .Z(n53157) );
  XOR U53067 ( .A(p_input[1701]), .B(p_input[2053]), .Z(n53143) );
  XNOR U53068 ( .A(n53158), .B(n53159), .Z(n53039) );
  AND U53069 ( .A(n2089), .B(n53160), .Z(n53159) );
  XNOR U53070 ( .A(n53161), .B(n53162), .Z(n2089) );
  AND U53071 ( .A(n53163), .B(n53164), .Z(n53162) );
  XOR U53072 ( .A(n53053), .B(n53161), .Z(n53164) );
  XNOR U53073 ( .A(n53165), .B(n53161), .Z(n53163) );
  XOR U53074 ( .A(n53166), .B(n53167), .Z(n53161) );
  AND U53075 ( .A(n53168), .B(n53169), .Z(n53167) );
  XOR U53076 ( .A(n53068), .B(n53166), .Z(n53169) );
  XOR U53077 ( .A(n53166), .B(n53069), .Z(n53168) );
  XOR U53078 ( .A(n53170), .B(n53171), .Z(n53166) );
  AND U53079 ( .A(n53172), .B(n53173), .Z(n53171) );
  XOR U53080 ( .A(n53096), .B(n53170), .Z(n53173) );
  XOR U53081 ( .A(n53170), .B(n53097), .Z(n53172) );
  XOR U53082 ( .A(n53174), .B(n53175), .Z(n53170) );
  AND U53083 ( .A(n53176), .B(n53177), .Z(n53175) );
  XOR U53084 ( .A(n53174), .B(n53147), .Z(n53177) );
  XNOR U53085 ( .A(n53178), .B(n53179), .Z(n52999) );
  AND U53086 ( .A(n2093), .B(n53180), .Z(n53179) );
  XNOR U53087 ( .A(n53181), .B(n53182), .Z(n2093) );
  AND U53088 ( .A(n53183), .B(n53184), .Z(n53182) );
  XOR U53089 ( .A(n53181), .B(n53009), .Z(n53184) );
  XNOR U53090 ( .A(n53181), .B(n52969), .Z(n53183) );
  XOR U53091 ( .A(n53185), .B(n53186), .Z(n53181) );
  AND U53092 ( .A(n53187), .B(n53188), .Z(n53186) );
  XOR U53093 ( .A(n53185), .B(n52977), .Z(n53187) );
  XOR U53094 ( .A(n53189), .B(n53190), .Z(n52960) );
  AND U53095 ( .A(n2097), .B(n53180), .Z(n53190) );
  XNOR U53096 ( .A(n53178), .B(n53189), .Z(n53180) );
  XNOR U53097 ( .A(n53191), .B(n53192), .Z(n2097) );
  AND U53098 ( .A(n53193), .B(n53194), .Z(n53192) );
  XNOR U53099 ( .A(n53195), .B(n53191), .Z(n53194) );
  IV U53100 ( .A(n53009), .Z(n53195) );
  XOR U53101 ( .A(n53165), .B(n53196), .Z(n53009) );
  AND U53102 ( .A(n2100), .B(n53197), .Z(n53196) );
  XOR U53103 ( .A(n53052), .B(n53049), .Z(n53197) );
  IV U53104 ( .A(n53165), .Z(n53052) );
  XNOR U53105 ( .A(n52969), .B(n53191), .Z(n53193) );
  XOR U53106 ( .A(n53198), .B(n53199), .Z(n52969) );
  AND U53107 ( .A(n2116), .B(n53200), .Z(n53199) );
  XOR U53108 ( .A(n53185), .B(n53201), .Z(n53191) );
  AND U53109 ( .A(n53202), .B(n53188), .Z(n53201) );
  XNOR U53110 ( .A(n53019), .B(n53185), .Z(n53188) );
  XOR U53111 ( .A(n53069), .B(n53203), .Z(n53019) );
  AND U53112 ( .A(n2100), .B(n53204), .Z(n53203) );
  XOR U53113 ( .A(n53065), .B(n53069), .Z(n53204) );
  XNOR U53114 ( .A(n53205), .B(n53185), .Z(n53202) );
  IV U53115 ( .A(n52977), .Z(n53205) );
  XOR U53116 ( .A(n53206), .B(n53207), .Z(n52977) );
  AND U53117 ( .A(n2116), .B(n53208), .Z(n53207) );
  XOR U53118 ( .A(n53209), .B(n53210), .Z(n53185) );
  AND U53119 ( .A(n53211), .B(n53212), .Z(n53210) );
  XNOR U53120 ( .A(n53029), .B(n53209), .Z(n53212) );
  XOR U53121 ( .A(n53097), .B(n53213), .Z(n53029) );
  AND U53122 ( .A(n2100), .B(n53214), .Z(n53213) );
  XOR U53123 ( .A(n53093), .B(n53097), .Z(n53214) );
  XOR U53124 ( .A(n53209), .B(n52986), .Z(n53211) );
  XOR U53125 ( .A(n53215), .B(n53216), .Z(n52986) );
  AND U53126 ( .A(n2116), .B(n53217), .Z(n53216) );
  XOR U53127 ( .A(n53218), .B(n53219), .Z(n53209) );
  AND U53128 ( .A(n53220), .B(n53221), .Z(n53219) );
  XNOR U53129 ( .A(n53218), .B(n53037), .Z(n53221) );
  XOR U53130 ( .A(n53148), .B(n53222), .Z(n53037) );
  AND U53131 ( .A(n2100), .B(n53223), .Z(n53222) );
  XOR U53132 ( .A(n53144), .B(n53148), .Z(n53223) );
  XNOR U53133 ( .A(n53224), .B(n53218), .Z(n53220) );
  IV U53134 ( .A(n52996), .Z(n53224) );
  XOR U53135 ( .A(n53225), .B(n53226), .Z(n52996) );
  AND U53136 ( .A(n2116), .B(n53227), .Z(n53226) );
  AND U53137 ( .A(n53189), .B(n53178), .Z(n53218) );
  XNOR U53138 ( .A(n53228), .B(n53229), .Z(n53178) );
  AND U53139 ( .A(n2100), .B(n53160), .Z(n53229) );
  XNOR U53140 ( .A(n53158), .B(n53228), .Z(n53160) );
  XNOR U53141 ( .A(n53230), .B(n53231), .Z(n2100) );
  AND U53142 ( .A(n53232), .B(n53233), .Z(n53231) );
  XNOR U53143 ( .A(n53230), .B(n53049), .Z(n53233) );
  IV U53144 ( .A(n53053), .Z(n53049) );
  XOR U53145 ( .A(n53234), .B(n53235), .Z(n53053) );
  AND U53146 ( .A(n2104), .B(n53236), .Z(n53235) );
  XOR U53147 ( .A(n53237), .B(n53234), .Z(n53236) );
  XNOR U53148 ( .A(n53230), .B(n53165), .Z(n53232) );
  XOR U53149 ( .A(n53238), .B(n53239), .Z(n53165) );
  AND U53150 ( .A(n2112), .B(n53200), .Z(n53239) );
  XOR U53151 ( .A(n53198), .B(n53238), .Z(n53200) );
  XOR U53152 ( .A(n53240), .B(n53241), .Z(n53230) );
  AND U53153 ( .A(n53242), .B(n53243), .Z(n53241) );
  XNOR U53154 ( .A(n53240), .B(n53065), .Z(n53243) );
  IV U53155 ( .A(n53068), .Z(n53065) );
  XOR U53156 ( .A(n53244), .B(n53245), .Z(n53068) );
  AND U53157 ( .A(n2104), .B(n53246), .Z(n53245) );
  XOR U53158 ( .A(n53247), .B(n53244), .Z(n53246) );
  XOR U53159 ( .A(n53069), .B(n53240), .Z(n53242) );
  XOR U53160 ( .A(n53248), .B(n53249), .Z(n53069) );
  AND U53161 ( .A(n2112), .B(n53208), .Z(n53249) );
  XOR U53162 ( .A(n53248), .B(n53206), .Z(n53208) );
  XOR U53163 ( .A(n53250), .B(n53251), .Z(n53240) );
  AND U53164 ( .A(n53252), .B(n53253), .Z(n53251) );
  XNOR U53165 ( .A(n53250), .B(n53093), .Z(n53253) );
  IV U53166 ( .A(n53096), .Z(n53093) );
  XOR U53167 ( .A(n53254), .B(n53255), .Z(n53096) );
  AND U53168 ( .A(n2104), .B(n53256), .Z(n53255) );
  XNOR U53169 ( .A(n53257), .B(n53254), .Z(n53256) );
  XOR U53170 ( .A(n53097), .B(n53250), .Z(n53252) );
  XOR U53171 ( .A(n53258), .B(n53259), .Z(n53097) );
  AND U53172 ( .A(n2112), .B(n53217), .Z(n53259) );
  XOR U53173 ( .A(n53258), .B(n53215), .Z(n53217) );
  XOR U53174 ( .A(n53174), .B(n53260), .Z(n53250) );
  AND U53175 ( .A(n53176), .B(n53261), .Z(n53260) );
  XNOR U53176 ( .A(n53174), .B(n53144), .Z(n53261) );
  IV U53177 ( .A(n53147), .Z(n53144) );
  XOR U53178 ( .A(n53262), .B(n53263), .Z(n53147) );
  AND U53179 ( .A(n2104), .B(n53264), .Z(n53263) );
  XOR U53180 ( .A(n53265), .B(n53262), .Z(n53264) );
  XOR U53181 ( .A(n53148), .B(n53174), .Z(n53176) );
  XOR U53182 ( .A(n53266), .B(n53267), .Z(n53148) );
  AND U53183 ( .A(n2112), .B(n53227), .Z(n53267) );
  XOR U53184 ( .A(n53266), .B(n53225), .Z(n53227) );
  AND U53185 ( .A(n53228), .B(n53158), .Z(n53174) );
  XNOR U53186 ( .A(n53268), .B(n53269), .Z(n53158) );
  AND U53187 ( .A(n2104), .B(n53270), .Z(n53269) );
  XNOR U53188 ( .A(n53271), .B(n53268), .Z(n53270) );
  XNOR U53189 ( .A(n53272), .B(n53273), .Z(n2104) );
  AND U53190 ( .A(n53274), .B(n53275), .Z(n53273) );
  XOR U53191 ( .A(n53237), .B(n53272), .Z(n53275) );
  AND U53192 ( .A(n53276), .B(n53277), .Z(n53237) );
  XNOR U53193 ( .A(n53234), .B(n53272), .Z(n53274) );
  XNOR U53194 ( .A(n53278), .B(n53279), .Z(n53234) );
  AND U53195 ( .A(n2108), .B(n53280), .Z(n53279) );
  XNOR U53196 ( .A(n53281), .B(n53282), .Z(n53280) );
  XOR U53197 ( .A(n53283), .B(n53284), .Z(n53272) );
  AND U53198 ( .A(n53285), .B(n53286), .Z(n53284) );
  XNOR U53199 ( .A(n53283), .B(n53276), .Z(n53286) );
  IV U53200 ( .A(n53247), .Z(n53276) );
  XOR U53201 ( .A(n53287), .B(n53288), .Z(n53247) );
  XOR U53202 ( .A(n53289), .B(n53277), .Z(n53288) );
  AND U53203 ( .A(n53257), .B(n53290), .Z(n53277) );
  AND U53204 ( .A(n53291), .B(n53292), .Z(n53289) );
  XOR U53205 ( .A(n53293), .B(n53287), .Z(n53291) );
  XNOR U53206 ( .A(n53244), .B(n53283), .Z(n53285) );
  XNOR U53207 ( .A(n53294), .B(n53295), .Z(n53244) );
  AND U53208 ( .A(n2108), .B(n53296), .Z(n53295) );
  XNOR U53209 ( .A(n53297), .B(n53298), .Z(n53296) );
  XOR U53210 ( .A(n53299), .B(n53300), .Z(n53283) );
  AND U53211 ( .A(n53301), .B(n53302), .Z(n53300) );
  XNOR U53212 ( .A(n53299), .B(n53257), .Z(n53302) );
  XOR U53213 ( .A(n53303), .B(n53292), .Z(n53257) );
  XNOR U53214 ( .A(n53304), .B(n53287), .Z(n53292) );
  XOR U53215 ( .A(n53305), .B(n53306), .Z(n53287) );
  AND U53216 ( .A(n53307), .B(n53308), .Z(n53306) );
  XOR U53217 ( .A(n53309), .B(n53305), .Z(n53307) );
  XNOR U53218 ( .A(n53310), .B(n53311), .Z(n53304) );
  AND U53219 ( .A(n53312), .B(n53313), .Z(n53311) );
  XOR U53220 ( .A(n53310), .B(n53314), .Z(n53312) );
  XNOR U53221 ( .A(n53293), .B(n53290), .Z(n53303) );
  AND U53222 ( .A(n53315), .B(n53316), .Z(n53290) );
  XOR U53223 ( .A(n53317), .B(n53318), .Z(n53293) );
  AND U53224 ( .A(n53319), .B(n53320), .Z(n53318) );
  XOR U53225 ( .A(n53317), .B(n53321), .Z(n53319) );
  XNOR U53226 ( .A(n53254), .B(n53299), .Z(n53301) );
  XNOR U53227 ( .A(n53322), .B(n53323), .Z(n53254) );
  AND U53228 ( .A(n2108), .B(n53324), .Z(n53323) );
  XNOR U53229 ( .A(n53325), .B(n53326), .Z(n53324) );
  XOR U53230 ( .A(n53327), .B(n53328), .Z(n53299) );
  AND U53231 ( .A(n53329), .B(n53330), .Z(n53328) );
  XNOR U53232 ( .A(n53327), .B(n53315), .Z(n53330) );
  IV U53233 ( .A(n53265), .Z(n53315) );
  XNOR U53234 ( .A(n53331), .B(n53308), .Z(n53265) );
  XNOR U53235 ( .A(n53332), .B(n53314), .Z(n53308) );
  XNOR U53236 ( .A(n53333), .B(n53334), .Z(n53314) );
  NOR U53237 ( .A(n53335), .B(n53336), .Z(n53334) );
  XOR U53238 ( .A(n53333), .B(n53337), .Z(n53335) );
  XNOR U53239 ( .A(n53313), .B(n53305), .Z(n53332) );
  XOR U53240 ( .A(n53338), .B(n53339), .Z(n53305) );
  AND U53241 ( .A(n53340), .B(n53341), .Z(n53339) );
  XOR U53242 ( .A(n53338), .B(n53342), .Z(n53340) );
  XNOR U53243 ( .A(n53343), .B(n53310), .Z(n53313) );
  XOR U53244 ( .A(n53344), .B(n53345), .Z(n53310) );
  AND U53245 ( .A(n53346), .B(n53347), .Z(n53345) );
  XNOR U53246 ( .A(n53348), .B(n53349), .Z(n53346) );
  IV U53247 ( .A(n53344), .Z(n53348) );
  XNOR U53248 ( .A(n53350), .B(n53351), .Z(n53343) );
  NOR U53249 ( .A(n53352), .B(n53353), .Z(n53351) );
  XNOR U53250 ( .A(n53350), .B(n53354), .Z(n53352) );
  XNOR U53251 ( .A(n53309), .B(n53316), .Z(n53331) );
  NOR U53252 ( .A(n53271), .B(n53355), .Z(n53316) );
  XOR U53253 ( .A(n53321), .B(n53320), .Z(n53309) );
  XNOR U53254 ( .A(n53356), .B(n53317), .Z(n53320) );
  XOR U53255 ( .A(n53357), .B(n53358), .Z(n53317) );
  AND U53256 ( .A(n53359), .B(n53360), .Z(n53358) );
  XNOR U53257 ( .A(n53361), .B(n53362), .Z(n53359) );
  IV U53258 ( .A(n53357), .Z(n53361) );
  XNOR U53259 ( .A(n53363), .B(n53364), .Z(n53356) );
  NOR U53260 ( .A(n53365), .B(n53366), .Z(n53364) );
  XNOR U53261 ( .A(n53363), .B(n53367), .Z(n53365) );
  XOR U53262 ( .A(n53368), .B(n53369), .Z(n53321) );
  NOR U53263 ( .A(n53370), .B(n53371), .Z(n53369) );
  XNOR U53264 ( .A(n53368), .B(n53372), .Z(n53370) );
  XNOR U53265 ( .A(n53262), .B(n53327), .Z(n53329) );
  XNOR U53266 ( .A(n53373), .B(n53374), .Z(n53262) );
  AND U53267 ( .A(n2108), .B(n53375), .Z(n53374) );
  XNOR U53268 ( .A(n53376), .B(n53377), .Z(n53375) );
  AND U53269 ( .A(n53268), .B(n53271), .Z(n53327) );
  XOR U53270 ( .A(n53378), .B(n53355), .Z(n53271) );
  XNOR U53271 ( .A(p_input[1712]), .B(p_input[2048]), .Z(n53355) );
  XNOR U53272 ( .A(n53342), .B(n53341), .Z(n53378) );
  XNOR U53273 ( .A(n53379), .B(n53349), .Z(n53341) );
  XNOR U53274 ( .A(n53337), .B(n53336), .Z(n53349) );
  XNOR U53275 ( .A(n53380), .B(n53333), .Z(n53336) );
  XNOR U53276 ( .A(p_input[1722]), .B(p_input[2058]), .Z(n53333) );
  XOR U53277 ( .A(p_input[1723]), .B(n29030), .Z(n53380) );
  XOR U53278 ( .A(p_input[1724]), .B(p_input[2060]), .Z(n53337) );
  XOR U53279 ( .A(n53347), .B(n53381), .Z(n53379) );
  IV U53280 ( .A(n53338), .Z(n53381) );
  XOR U53281 ( .A(p_input[1713]), .B(p_input[2049]), .Z(n53338) );
  XNOR U53282 ( .A(n53382), .B(n53354), .Z(n53347) );
  XNOR U53283 ( .A(p_input[1727]), .B(n29033), .Z(n53354) );
  XOR U53284 ( .A(n53344), .B(n53353), .Z(n53382) );
  XOR U53285 ( .A(n53383), .B(n53350), .Z(n53353) );
  XOR U53286 ( .A(p_input[1725]), .B(p_input[2061]), .Z(n53350) );
  XOR U53287 ( .A(p_input[1726]), .B(n29035), .Z(n53383) );
  XOR U53288 ( .A(p_input[1721]), .B(p_input[2057]), .Z(n53344) );
  XOR U53289 ( .A(n53362), .B(n53360), .Z(n53342) );
  XNOR U53290 ( .A(n53384), .B(n53367), .Z(n53360) );
  XOR U53291 ( .A(p_input[1720]), .B(p_input[2056]), .Z(n53367) );
  XOR U53292 ( .A(n53357), .B(n53366), .Z(n53384) );
  XOR U53293 ( .A(n53385), .B(n53363), .Z(n53366) );
  XOR U53294 ( .A(p_input[1718]), .B(p_input[2054]), .Z(n53363) );
  XOR U53295 ( .A(p_input[1719]), .B(n30404), .Z(n53385) );
  XOR U53296 ( .A(p_input[1714]), .B(p_input[2050]), .Z(n53357) );
  XNOR U53297 ( .A(n53372), .B(n53371), .Z(n53362) );
  XOR U53298 ( .A(n53386), .B(n53368), .Z(n53371) );
  XOR U53299 ( .A(p_input[1715]), .B(p_input[2051]), .Z(n53368) );
  XOR U53300 ( .A(p_input[1716]), .B(n30406), .Z(n53386) );
  XOR U53301 ( .A(p_input[1717]), .B(p_input[2053]), .Z(n53372) );
  XNOR U53302 ( .A(n53387), .B(n53388), .Z(n53268) );
  AND U53303 ( .A(n2108), .B(n53389), .Z(n53388) );
  XNOR U53304 ( .A(n53390), .B(n53391), .Z(n2108) );
  AND U53305 ( .A(n53392), .B(n53393), .Z(n53391) );
  XOR U53306 ( .A(n53282), .B(n53390), .Z(n53393) );
  XNOR U53307 ( .A(n53394), .B(n53390), .Z(n53392) );
  XOR U53308 ( .A(n53395), .B(n53396), .Z(n53390) );
  AND U53309 ( .A(n53397), .B(n53398), .Z(n53396) );
  XOR U53310 ( .A(n53297), .B(n53395), .Z(n53398) );
  XOR U53311 ( .A(n53395), .B(n53298), .Z(n53397) );
  XOR U53312 ( .A(n53399), .B(n53400), .Z(n53395) );
  AND U53313 ( .A(n53401), .B(n53402), .Z(n53400) );
  XOR U53314 ( .A(n53325), .B(n53399), .Z(n53402) );
  XOR U53315 ( .A(n53399), .B(n53326), .Z(n53401) );
  XOR U53316 ( .A(n53403), .B(n53404), .Z(n53399) );
  AND U53317 ( .A(n53405), .B(n53406), .Z(n53404) );
  XOR U53318 ( .A(n53403), .B(n53376), .Z(n53406) );
  XNOR U53319 ( .A(n53407), .B(n53408), .Z(n53228) );
  AND U53320 ( .A(n2112), .B(n53409), .Z(n53408) );
  XNOR U53321 ( .A(n53410), .B(n53411), .Z(n2112) );
  AND U53322 ( .A(n53412), .B(n53413), .Z(n53411) );
  XOR U53323 ( .A(n53410), .B(n53238), .Z(n53413) );
  XNOR U53324 ( .A(n53410), .B(n53198), .Z(n53412) );
  XOR U53325 ( .A(n53414), .B(n53415), .Z(n53410) );
  AND U53326 ( .A(n53416), .B(n53417), .Z(n53415) );
  XOR U53327 ( .A(n53414), .B(n53206), .Z(n53416) );
  XOR U53328 ( .A(n53418), .B(n53419), .Z(n53189) );
  AND U53329 ( .A(n2116), .B(n53409), .Z(n53419) );
  XNOR U53330 ( .A(n53407), .B(n53418), .Z(n53409) );
  XNOR U53331 ( .A(n53420), .B(n53421), .Z(n2116) );
  AND U53332 ( .A(n53422), .B(n53423), .Z(n53421) );
  XNOR U53333 ( .A(n53424), .B(n53420), .Z(n53423) );
  IV U53334 ( .A(n53238), .Z(n53424) );
  XOR U53335 ( .A(n53394), .B(n53425), .Z(n53238) );
  AND U53336 ( .A(n2119), .B(n53426), .Z(n53425) );
  XOR U53337 ( .A(n53281), .B(n53278), .Z(n53426) );
  IV U53338 ( .A(n53394), .Z(n53281) );
  XNOR U53339 ( .A(n53198), .B(n53420), .Z(n53422) );
  XOR U53340 ( .A(n53427), .B(n53428), .Z(n53198) );
  AND U53341 ( .A(n2135), .B(n53429), .Z(n53428) );
  XOR U53342 ( .A(n53414), .B(n53430), .Z(n53420) );
  AND U53343 ( .A(n53431), .B(n53417), .Z(n53430) );
  XNOR U53344 ( .A(n53248), .B(n53414), .Z(n53417) );
  XOR U53345 ( .A(n53298), .B(n53432), .Z(n53248) );
  AND U53346 ( .A(n2119), .B(n53433), .Z(n53432) );
  XOR U53347 ( .A(n53294), .B(n53298), .Z(n53433) );
  XNOR U53348 ( .A(n53434), .B(n53414), .Z(n53431) );
  IV U53349 ( .A(n53206), .Z(n53434) );
  XOR U53350 ( .A(n53435), .B(n53436), .Z(n53206) );
  AND U53351 ( .A(n2135), .B(n53437), .Z(n53436) );
  XOR U53352 ( .A(n53438), .B(n53439), .Z(n53414) );
  AND U53353 ( .A(n53440), .B(n53441), .Z(n53439) );
  XNOR U53354 ( .A(n53258), .B(n53438), .Z(n53441) );
  XOR U53355 ( .A(n53326), .B(n53442), .Z(n53258) );
  AND U53356 ( .A(n2119), .B(n53443), .Z(n53442) );
  XOR U53357 ( .A(n53322), .B(n53326), .Z(n53443) );
  XOR U53358 ( .A(n53438), .B(n53215), .Z(n53440) );
  XOR U53359 ( .A(n53444), .B(n53445), .Z(n53215) );
  AND U53360 ( .A(n2135), .B(n53446), .Z(n53445) );
  XOR U53361 ( .A(n53447), .B(n53448), .Z(n53438) );
  AND U53362 ( .A(n53449), .B(n53450), .Z(n53448) );
  XNOR U53363 ( .A(n53447), .B(n53266), .Z(n53450) );
  XOR U53364 ( .A(n53377), .B(n53451), .Z(n53266) );
  AND U53365 ( .A(n2119), .B(n53452), .Z(n53451) );
  XOR U53366 ( .A(n53373), .B(n53377), .Z(n53452) );
  XNOR U53367 ( .A(n53453), .B(n53447), .Z(n53449) );
  IV U53368 ( .A(n53225), .Z(n53453) );
  XOR U53369 ( .A(n53454), .B(n53455), .Z(n53225) );
  AND U53370 ( .A(n2135), .B(n53456), .Z(n53455) );
  AND U53371 ( .A(n53418), .B(n53407), .Z(n53447) );
  XNOR U53372 ( .A(n53457), .B(n53458), .Z(n53407) );
  AND U53373 ( .A(n2119), .B(n53389), .Z(n53458) );
  XNOR U53374 ( .A(n53387), .B(n53457), .Z(n53389) );
  XNOR U53375 ( .A(n53459), .B(n53460), .Z(n2119) );
  AND U53376 ( .A(n53461), .B(n53462), .Z(n53460) );
  XNOR U53377 ( .A(n53459), .B(n53278), .Z(n53462) );
  IV U53378 ( .A(n53282), .Z(n53278) );
  XOR U53379 ( .A(n53463), .B(n53464), .Z(n53282) );
  AND U53380 ( .A(n2123), .B(n53465), .Z(n53464) );
  XOR U53381 ( .A(n53466), .B(n53463), .Z(n53465) );
  XNOR U53382 ( .A(n53459), .B(n53394), .Z(n53461) );
  XOR U53383 ( .A(n53467), .B(n53468), .Z(n53394) );
  AND U53384 ( .A(n2131), .B(n53429), .Z(n53468) );
  XOR U53385 ( .A(n53427), .B(n53467), .Z(n53429) );
  XOR U53386 ( .A(n53469), .B(n53470), .Z(n53459) );
  AND U53387 ( .A(n53471), .B(n53472), .Z(n53470) );
  XNOR U53388 ( .A(n53469), .B(n53294), .Z(n53472) );
  IV U53389 ( .A(n53297), .Z(n53294) );
  XOR U53390 ( .A(n53473), .B(n53474), .Z(n53297) );
  AND U53391 ( .A(n2123), .B(n53475), .Z(n53474) );
  XOR U53392 ( .A(n53476), .B(n53473), .Z(n53475) );
  XOR U53393 ( .A(n53298), .B(n53469), .Z(n53471) );
  XOR U53394 ( .A(n53477), .B(n53478), .Z(n53298) );
  AND U53395 ( .A(n2131), .B(n53437), .Z(n53478) );
  XOR U53396 ( .A(n53477), .B(n53435), .Z(n53437) );
  XOR U53397 ( .A(n53479), .B(n53480), .Z(n53469) );
  AND U53398 ( .A(n53481), .B(n53482), .Z(n53480) );
  XNOR U53399 ( .A(n53479), .B(n53322), .Z(n53482) );
  IV U53400 ( .A(n53325), .Z(n53322) );
  XOR U53401 ( .A(n53483), .B(n53484), .Z(n53325) );
  AND U53402 ( .A(n2123), .B(n53485), .Z(n53484) );
  XNOR U53403 ( .A(n53486), .B(n53483), .Z(n53485) );
  XOR U53404 ( .A(n53326), .B(n53479), .Z(n53481) );
  XOR U53405 ( .A(n53487), .B(n53488), .Z(n53326) );
  AND U53406 ( .A(n2131), .B(n53446), .Z(n53488) );
  XOR U53407 ( .A(n53487), .B(n53444), .Z(n53446) );
  XOR U53408 ( .A(n53403), .B(n53489), .Z(n53479) );
  AND U53409 ( .A(n53405), .B(n53490), .Z(n53489) );
  XNOR U53410 ( .A(n53403), .B(n53373), .Z(n53490) );
  IV U53411 ( .A(n53376), .Z(n53373) );
  XOR U53412 ( .A(n53491), .B(n53492), .Z(n53376) );
  AND U53413 ( .A(n2123), .B(n53493), .Z(n53492) );
  XOR U53414 ( .A(n53494), .B(n53491), .Z(n53493) );
  XOR U53415 ( .A(n53377), .B(n53403), .Z(n53405) );
  XOR U53416 ( .A(n53495), .B(n53496), .Z(n53377) );
  AND U53417 ( .A(n2131), .B(n53456), .Z(n53496) );
  XOR U53418 ( .A(n53495), .B(n53454), .Z(n53456) );
  AND U53419 ( .A(n53457), .B(n53387), .Z(n53403) );
  XNOR U53420 ( .A(n53497), .B(n53498), .Z(n53387) );
  AND U53421 ( .A(n2123), .B(n53499), .Z(n53498) );
  XNOR U53422 ( .A(n53500), .B(n53497), .Z(n53499) );
  XNOR U53423 ( .A(n53501), .B(n53502), .Z(n2123) );
  AND U53424 ( .A(n53503), .B(n53504), .Z(n53502) );
  XOR U53425 ( .A(n53466), .B(n53501), .Z(n53504) );
  AND U53426 ( .A(n53505), .B(n53506), .Z(n53466) );
  XNOR U53427 ( .A(n53463), .B(n53501), .Z(n53503) );
  XNOR U53428 ( .A(n53507), .B(n53508), .Z(n53463) );
  AND U53429 ( .A(n2127), .B(n53509), .Z(n53508) );
  XNOR U53430 ( .A(n53510), .B(n53511), .Z(n53509) );
  XOR U53431 ( .A(n53512), .B(n53513), .Z(n53501) );
  AND U53432 ( .A(n53514), .B(n53515), .Z(n53513) );
  XNOR U53433 ( .A(n53512), .B(n53505), .Z(n53515) );
  IV U53434 ( .A(n53476), .Z(n53505) );
  XOR U53435 ( .A(n53516), .B(n53517), .Z(n53476) );
  XOR U53436 ( .A(n53518), .B(n53506), .Z(n53517) );
  AND U53437 ( .A(n53486), .B(n53519), .Z(n53506) );
  AND U53438 ( .A(n53520), .B(n53521), .Z(n53518) );
  XOR U53439 ( .A(n53522), .B(n53516), .Z(n53520) );
  XNOR U53440 ( .A(n53473), .B(n53512), .Z(n53514) );
  XNOR U53441 ( .A(n53523), .B(n53524), .Z(n53473) );
  AND U53442 ( .A(n2127), .B(n53525), .Z(n53524) );
  XNOR U53443 ( .A(n53526), .B(n53527), .Z(n53525) );
  XOR U53444 ( .A(n53528), .B(n53529), .Z(n53512) );
  AND U53445 ( .A(n53530), .B(n53531), .Z(n53529) );
  XNOR U53446 ( .A(n53528), .B(n53486), .Z(n53531) );
  XOR U53447 ( .A(n53532), .B(n53521), .Z(n53486) );
  XNOR U53448 ( .A(n53533), .B(n53516), .Z(n53521) );
  XOR U53449 ( .A(n53534), .B(n53535), .Z(n53516) );
  AND U53450 ( .A(n53536), .B(n53537), .Z(n53535) );
  XOR U53451 ( .A(n53538), .B(n53534), .Z(n53536) );
  XNOR U53452 ( .A(n53539), .B(n53540), .Z(n53533) );
  AND U53453 ( .A(n53541), .B(n53542), .Z(n53540) );
  XOR U53454 ( .A(n53539), .B(n53543), .Z(n53541) );
  XNOR U53455 ( .A(n53522), .B(n53519), .Z(n53532) );
  AND U53456 ( .A(n53544), .B(n53545), .Z(n53519) );
  XOR U53457 ( .A(n53546), .B(n53547), .Z(n53522) );
  AND U53458 ( .A(n53548), .B(n53549), .Z(n53547) );
  XOR U53459 ( .A(n53546), .B(n53550), .Z(n53548) );
  XNOR U53460 ( .A(n53483), .B(n53528), .Z(n53530) );
  XNOR U53461 ( .A(n53551), .B(n53552), .Z(n53483) );
  AND U53462 ( .A(n2127), .B(n53553), .Z(n53552) );
  XNOR U53463 ( .A(n53554), .B(n53555), .Z(n53553) );
  XOR U53464 ( .A(n53556), .B(n53557), .Z(n53528) );
  AND U53465 ( .A(n53558), .B(n53559), .Z(n53557) );
  XNOR U53466 ( .A(n53556), .B(n53544), .Z(n53559) );
  IV U53467 ( .A(n53494), .Z(n53544) );
  XNOR U53468 ( .A(n53560), .B(n53537), .Z(n53494) );
  XNOR U53469 ( .A(n53561), .B(n53543), .Z(n53537) );
  XNOR U53470 ( .A(n53562), .B(n53563), .Z(n53543) );
  NOR U53471 ( .A(n53564), .B(n53565), .Z(n53563) );
  XOR U53472 ( .A(n53562), .B(n53566), .Z(n53564) );
  XNOR U53473 ( .A(n53542), .B(n53534), .Z(n53561) );
  XOR U53474 ( .A(n53567), .B(n53568), .Z(n53534) );
  AND U53475 ( .A(n53569), .B(n53570), .Z(n53568) );
  XOR U53476 ( .A(n53567), .B(n53571), .Z(n53569) );
  XNOR U53477 ( .A(n53572), .B(n53539), .Z(n53542) );
  XOR U53478 ( .A(n53573), .B(n53574), .Z(n53539) );
  AND U53479 ( .A(n53575), .B(n53576), .Z(n53574) );
  XNOR U53480 ( .A(n53577), .B(n53578), .Z(n53575) );
  IV U53481 ( .A(n53573), .Z(n53577) );
  XNOR U53482 ( .A(n53579), .B(n53580), .Z(n53572) );
  NOR U53483 ( .A(n53581), .B(n53582), .Z(n53580) );
  XNOR U53484 ( .A(n53579), .B(n53583), .Z(n53581) );
  XNOR U53485 ( .A(n53538), .B(n53545), .Z(n53560) );
  NOR U53486 ( .A(n53500), .B(n53584), .Z(n53545) );
  XOR U53487 ( .A(n53550), .B(n53549), .Z(n53538) );
  XNOR U53488 ( .A(n53585), .B(n53546), .Z(n53549) );
  XOR U53489 ( .A(n53586), .B(n53587), .Z(n53546) );
  AND U53490 ( .A(n53588), .B(n53589), .Z(n53587) );
  XNOR U53491 ( .A(n53590), .B(n53591), .Z(n53588) );
  IV U53492 ( .A(n53586), .Z(n53590) );
  XNOR U53493 ( .A(n53592), .B(n53593), .Z(n53585) );
  NOR U53494 ( .A(n53594), .B(n53595), .Z(n53593) );
  XNOR U53495 ( .A(n53592), .B(n53596), .Z(n53594) );
  XOR U53496 ( .A(n53597), .B(n53598), .Z(n53550) );
  NOR U53497 ( .A(n53599), .B(n53600), .Z(n53598) );
  XNOR U53498 ( .A(n53597), .B(n53601), .Z(n53599) );
  XNOR U53499 ( .A(n53491), .B(n53556), .Z(n53558) );
  XNOR U53500 ( .A(n53602), .B(n53603), .Z(n53491) );
  AND U53501 ( .A(n2127), .B(n53604), .Z(n53603) );
  XNOR U53502 ( .A(n53605), .B(n53606), .Z(n53604) );
  AND U53503 ( .A(n53497), .B(n53500), .Z(n53556) );
  XOR U53504 ( .A(n53607), .B(n53584), .Z(n53500) );
  XNOR U53505 ( .A(p_input[1728]), .B(p_input[2048]), .Z(n53584) );
  XNOR U53506 ( .A(n53571), .B(n53570), .Z(n53607) );
  XNOR U53507 ( .A(n53608), .B(n53578), .Z(n53570) );
  XNOR U53508 ( .A(n53566), .B(n53565), .Z(n53578) );
  XNOR U53509 ( .A(n53609), .B(n53562), .Z(n53565) );
  XNOR U53510 ( .A(p_input[1738]), .B(p_input[2058]), .Z(n53562) );
  XOR U53511 ( .A(p_input[1739]), .B(n29030), .Z(n53609) );
  XOR U53512 ( .A(p_input[1740]), .B(p_input[2060]), .Z(n53566) );
  XOR U53513 ( .A(n53576), .B(n53610), .Z(n53608) );
  IV U53514 ( .A(n53567), .Z(n53610) );
  XOR U53515 ( .A(p_input[1729]), .B(p_input[2049]), .Z(n53567) );
  XNOR U53516 ( .A(n53611), .B(n53583), .Z(n53576) );
  XNOR U53517 ( .A(p_input[1743]), .B(n29033), .Z(n53583) );
  XOR U53518 ( .A(n53573), .B(n53582), .Z(n53611) );
  XOR U53519 ( .A(n53612), .B(n53579), .Z(n53582) );
  XOR U53520 ( .A(p_input[1741]), .B(p_input[2061]), .Z(n53579) );
  XOR U53521 ( .A(p_input[1742]), .B(n29035), .Z(n53612) );
  XOR U53522 ( .A(p_input[1737]), .B(p_input[2057]), .Z(n53573) );
  XOR U53523 ( .A(n53591), .B(n53589), .Z(n53571) );
  XNOR U53524 ( .A(n53613), .B(n53596), .Z(n53589) );
  XOR U53525 ( .A(p_input[1736]), .B(p_input[2056]), .Z(n53596) );
  XOR U53526 ( .A(n53586), .B(n53595), .Z(n53613) );
  XOR U53527 ( .A(n53614), .B(n53592), .Z(n53595) );
  XOR U53528 ( .A(p_input[1734]), .B(p_input[2054]), .Z(n53592) );
  XOR U53529 ( .A(p_input[1735]), .B(n30404), .Z(n53614) );
  XOR U53530 ( .A(p_input[1730]), .B(p_input[2050]), .Z(n53586) );
  XNOR U53531 ( .A(n53601), .B(n53600), .Z(n53591) );
  XOR U53532 ( .A(n53615), .B(n53597), .Z(n53600) );
  XOR U53533 ( .A(p_input[1731]), .B(p_input[2051]), .Z(n53597) );
  XOR U53534 ( .A(p_input[1732]), .B(n30406), .Z(n53615) );
  XOR U53535 ( .A(p_input[1733]), .B(p_input[2053]), .Z(n53601) );
  XNOR U53536 ( .A(n53616), .B(n53617), .Z(n53497) );
  AND U53537 ( .A(n2127), .B(n53618), .Z(n53617) );
  XNOR U53538 ( .A(n53619), .B(n53620), .Z(n2127) );
  AND U53539 ( .A(n53621), .B(n53622), .Z(n53620) );
  XOR U53540 ( .A(n53511), .B(n53619), .Z(n53622) );
  XNOR U53541 ( .A(n53623), .B(n53619), .Z(n53621) );
  XOR U53542 ( .A(n53624), .B(n53625), .Z(n53619) );
  AND U53543 ( .A(n53626), .B(n53627), .Z(n53625) );
  XOR U53544 ( .A(n53526), .B(n53624), .Z(n53627) );
  XOR U53545 ( .A(n53624), .B(n53527), .Z(n53626) );
  XOR U53546 ( .A(n53628), .B(n53629), .Z(n53624) );
  AND U53547 ( .A(n53630), .B(n53631), .Z(n53629) );
  XOR U53548 ( .A(n53554), .B(n53628), .Z(n53631) );
  XOR U53549 ( .A(n53628), .B(n53555), .Z(n53630) );
  XOR U53550 ( .A(n53632), .B(n53633), .Z(n53628) );
  AND U53551 ( .A(n53634), .B(n53635), .Z(n53633) );
  XOR U53552 ( .A(n53632), .B(n53605), .Z(n53635) );
  XNOR U53553 ( .A(n53636), .B(n53637), .Z(n53457) );
  AND U53554 ( .A(n2131), .B(n53638), .Z(n53637) );
  XNOR U53555 ( .A(n53639), .B(n53640), .Z(n2131) );
  AND U53556 ( .A(n53641), .B(n53642), .Z(n53640) );
  XOR U53557 ( .A(n53639), .B(n53467), .Z(n53642) );
  XNOR U53558 ( .A(n53639), .B(n53427), .Z(n53641) );
  XOR U53559 ( .A(n53643), .B(n53644), .Z(n53639) );
  AND U53560 ( .A(n53645), .B(n53646), .Z(n53644) );
  XOR U53561 ( .A(n53643), .B(n53435), .Z(n53645) );
  XOR U53562 ( .A(n53647), .B(n53648), .Z(n53418) );
  AND U53563 ( .A(n2135), .B(n53638), .Z(n53648) );
  XNOR U53564 ( .A(n53636), .B(n53647), .Z(n53638) );
  XNOR U53565 ( .A(n53649), .B(n53650), .Z(n2135) );
  AND U53566 ( .A(n53651), .B(n53652), .Z(n53650) );
  XNOR U53567 ( .A(n53653), .B(n53649), .Z(n53652) );
  IV U53568 ( .A(n53467), .Z(n53653) );
  XOR U53569 ( .A(n53623), .B(n53654), .Z(n53467) );
  AND U53570 ( .A(n2138), .B(n53655), .Z(n53654) );
  XOR U53571 ( .A(n53510), .B(n53507), .Z(n53655) );
  IV U53572 ( .A(n53623), .Z(n53510) );
  XNOR U53573 ( .A(n53427), .B(n53649), .Z(n53651) );
  XOR U53574 ( .A(n53656), .B(n53657), .Z(n53427) );
  AND U53575 ( .A(n2154), .B(n53658), .Z(n53657) );
  XOR U53576 ( .A(n53643), .B(n53659), .Z(n53649) );
  AND U53577 ( .A(n53660), .B(n53646), .Z(n53659) );
  XNOR U53578 ( .A(n53477), .B(n53643), .Z(n53646) );
  XOR U53579 ( .A(n53527), .B(n53661), .Z(n53477) );
  AND U53580 ( .A(n2138), .B(n53662), .Z(n53661) );
  XOR U53581 ( .A(n53523), .B(n53527), .Z(n53662) );
  XNOR U53582 ( .A(n53663), .B(n53643), .Z(n53660) );
  IV U53583 ( .A(n53435), .Z(n53663) );
  XOR U53584 ( .A(n53664), .B(n53665), .Z(n53435) );
  AND U53585 ( .A(n2154), .B(n53666), .Z(n53665) );
  XOR U53586 ( .A(n53667), .B(n53668), .Z(n53643) );
  AND U53587 ( .A(n53669), .B(n53670), .Z(n53668) );
  XNOR U53588 ( .A(n53487), .B(n53667), .Z(n53670) );
  XOR U53589 ( .A(n53555), .B(n53671), .Z(n53487) );
  AND U53590 ( .A(n2138), .B(n53672), .Z(n53671) );
  XOR U53591 ( .A(n53551), .B(n53555), .Z(n53672) );
  XOR U53592 ( .A(n53667), .B(n53444), .Z(n53669) );
  XOR U53593 ( .A(n53673), .B(n53674), .Z(n53444) );
  AND U53594 ( .A(n2154), .B(n53675), .Z(n53674) );
  XOR U53595 ( .A(n53676), .B(n53677), .Z(n53667) );
  AND U53596 ( .A(n53678), .B(n53679), .Z(n53677) );
  XNOR U53597 ( .A(n53676), .B(n53495), .Z(n53679) );
  XOR U53598 ( .A(n53606), .B(n53680), .Z(n53495) );
  AND U53599 ( .A(n2138), .B(n53681), .Z(n53680) );
  XOR U53600 ( .A(n53602), .B(n53606), .Z(n53681) );
  XNOR U53601 ( .A(n53682), .B(n53676), .Z(n53678) );
  IV U53602 ( .A(n53454), .Z(n53682) );
  XOR U53603 ( .A(n53683), .B(n53684), .Z(n53454) );
  AND U53604 ( .A(n2154), .B(n53685), .Z(n53684) );
  AND U53605 ( .A(n53647), .B(n53636), .Z(n53676) );
  XNOR U53606 ( .A(n53686), .B(n53687), .Z(n53636) );
  AND U53607 ( .A(n2138), .B(n53618), .Z(n53687) );
  XNOR U53608 ( .A(n53616), .B(n53686), .Z(n53618) );
  XNOR U53609 ( .A(n53688), .B(n53689), .Z(n2138) );
  AND U53610 ( .A(n53690), .B(n53691), .Z(n53689) );
  XNOR U53611 ( .A(n53688), .B(n53507), .Z(n53691) );
  IV U53612 ( .A(n53511), .Z(n53507) );
  XOR U53613 ( .A(n53692), .B(n53693), .Z(n53511) );
  AND U53614 ( .A(n2142), .B(n53694), .Z(n53693) );
  XOR U53615 ( .A(n53695), .B(n53692), .Z(n53694) );
  XNOR U53616 ( .A(n53688), .B(n53623), .Z(n53690) );
  XOR U53617 ( .A(n53696), .B(n53697), .Z(n53623) );
  AND U53618 ( .A(n2150), .B(n53658), .Z(n53697) );
  XOR U53619 ( .A(n53656), .B(n53696), .Z(n53658) );
  XOR U53620 ( .A(n53698), .B(n53699), .Z(n53688) );
  AND U53621 ( .A(n53700), .B(n53701), .Z(n53699) );
  XNOR U53622 ( .A(n53698), .B(n53523), .Z(n53701) );
  IV U53623 ( .A(n53526), .Z(n53523) );
  XOR U53624 ( .A(n53702), .B(n53703), .Z(n53526) );
  AND U53625 ( .A(n2142), .B(n53704), .Z(n53703) );
  XOR U53626 ( .A(n53705), .B(n53702), .Z(n53704) );
  XOR U53627 ( .A(n53527), .B(n53698), .Z(n53700) );
  XOR U53628 ( .A(n53706), .B(n53707), .Z(n53527) );
  AND U53629 ( .A(n2150), .B(n53666), .Z(n53707) );
  XOR U53630 ( .A(n53706), .B(n53664), .Z(n53666) );
  XOR U53631 ( .A(n53708), .B(n53709), .Z(n53698) );
  AND U53632 ( .A(n53710), .B(n53711), .Z(n53709) );
  XNOR U53633 ( .A(n53708), .B(n53551), .Z(n53711) );
  IV U53634 ( .A(n53554), .Z(n53551) );
  XOR U53635 ( .A(n53712), .B(n53713), .Z(n53554) );
  AND U53636 ( .A(n2142), .B(n53714), .Z(n53713) );
  XNOR U53637 ( .A(n53715), .B(n53712), .Z(n53714) );
  XOR U53638 ( .A(n53555), .B(n53708), .Z(n53710) );
  XOR U53639 ( .A(n53716), .B(n53717), .Z(n53555) );
  AND U53640 ( .A(n2150), .B(n53675), .Z(n53717) );
  XOR U53641 ( .A(n53716), .B(n53673), .Z(n53675) );
  XOR U53642 ( .A(n53632), .B(n53718), .Z(n53708) );
  AND U53643 ( .A(n53634), .B(n53719), .Z(n53718) );
  XNOR U53644 ( .A(n53632), .B(n53602), .Z(n53719) );
  IV U53645 ( .A(n53605), .Z(n53602) );
  XOR U53646 ( .A(n53720), .B(n53721), .Z(n53605) );
  AND U53647 ( .A(n2142), .B(n53722), .Z(n53721) );
  XOR U53648 ( .A(n53723), .B(n53720), .Z(n53722) );
  XOR U53649 ( .A(n53606), .B(n53632), .Z(n53634) );
  XOR U53650 ( .A(n53724), .B(n53725), .Z(n53606) );
  AND U53651 ( .A(n2150), .B(n53685), .Z(n53725) );
  XOR U53652 ( .A(n53724), .B(n53683), .Z(n53685) );
  AND U53653 ( .A(n53686), .B(n53616), .Z(n53632) );
  XNOR U53654 ( .A(n53726), .B(n53727), .Z(n53616) );
  AND U53655 ( .A(n2142), .B(n53728), .Z(n53727) );
  XNOR U53656 ( .A(n53729), .B(n53726), .Z(n53728) );
  XNOR U53657 ( .A(n53730), .B(n53731), .Z(n2142) );
  AND U53658 ( .A(n53732), .B(n53733), .Z(n53731) );
  XOR U53659 ( .A(n53695), .B(n53730), .Z(n53733) );
  AND U53660 ( .A(n53734), .B(n53735), .Z(n53695) );
  XNOR U53661 ( .A(n53692), .B(n53730), .Z(n53732) );
  XNOR U53662 ( .A(n53736), .B(n53737), .Z(n53692) );
  AND U53663 ( .A(n2146), .B(n53738), .Z(n53737) );
  XNOR U53664 ( .A(n53739), .B(n53740), .Z(n53738) );
  XOR U53665 ( .A(n53741), .B(n53742), .Z(n53730) );
  AND U53666 ( .A(n53743), .B(n53744), .Z(n53742) );
  XNOR U53667 ( .A(n53741), .B(n53734), .Z(n53744) );
  IV U53668 ( .A(n53705), .Z(n53734) );
  XOR U53669 ( .A(n53745), .B(n53746), .Z(n53705) );
  XOR U53670 ( .A(n53747), .B(n53735), .Z(n53746) );
  AND U53671 ( .A(n53715), .B(n53748), .Z(n53735) );
  AND U53672 ( .A(n53749), .B(n53750), .Z(n53747) );
  XOR U53673 ( .A(n53751), .B(n53745), .Z(n53749) );
  XNOR U53674 ( .A(n53702), .B(n53741), .Z(n53743) );
  XNOR U53675 ( .A(n53752), .B(n53753), .Z(n53702) );
  AND U53676 ( .A(n2146), .B(n53754), .Z(n53753) );
  XNOR U53677 ( .A(n53755), .B(n53756), .Z(n53754) );
  XOR U53678 ( .A(n53757), .B(n53758), .Z(n53741) );
  AND U53679 ( .A(n53759), .B(n53760), .Z(n53758) );
  XNOR U53680 ( .A(n53757), .B(n53715), .Z(n53760) );
  XOR U53681 ( .A(n53761), .B(n53750), .Z(n53715) );
  XNOR U53682 ( .A(n53762), .B(n53745), .Z(n53750) );
  XOR U53683 ( .A(n53763), .B(n53764), .Z(n53745) );
  AND U53684 ( .A(n53765), .B(n53766), .Z(n53764) );
  XOR U53685 ( .A(n53767), .B(n53763), .Z(n53765) );
  XNOR U53686 ( .A(n53768), .B(n53769), .Z(n53762) );
  AND U53687 ( .A(n53770), .B(n53771), .Z(n53769) );
  XOR U53688 ( .A(n53768), .B(n53772), .Z(n53770) );
  XNOR U53689 ( .A(n53751), .B(n53748), .Z(n53761) );
  AND U53690 ( .A(n53773), .B(n53774), .Z(n53748) );
  XOR U53691 ( .A(n53775), .B(n53776), .Z(n53751) );
  AND U53692 ( .A(n53777), .B(n53778), .Z(n53776) );
  XOR U53693 ( .A(n53775), .B(n53779), .Z(n53777) );
  XNOR U53694 ( .A(n53712), .B(n53757), .Z(n53759) );
  XNOR U53695 ( .A(n53780), .B(n53781), .Z(n53712) );
  AND U53696 ( .A(n2146), .B(n53782), .Z(n53781) );
  XNOR U53697 ( .A(n53783), .B(n53784), .Z(n53782) );
  XOR U53698 ( .A(n53785), .B(n53786), .Z(n53757) );
  AND U53699 ( .A(n53787), .B(n53788), .Z(n53786) );
  XNOR U53700 ( .A(n53785), .B(n53773), .Z(n53788) );
  IV U53701 ( .A(n53723), .Z(n53773) );
  XNOR U53702 ( .A(n53789), .B(n53766), .Z(n53723) );
  XNOR U53703 ( .A(n53790), .B(n53772), .Z(n53766) );
  XNOR U53704 ( .A(n53791), .B(n53792), .Z(n53772) );
  NOR U53705 ( .A(n53793), .B(n53794), .Z(n53792) );
  XOR U53706 ( .A(n53791), .B(n53795), .Z(n53793) );
  XNOR U53707 ( .A(n53771), .B(n53763), .Z(n53790) );
  XOR U53708 ( .A(n53796), .B(n53797), .Z(n53763) );
  AND U53709 ( .A(n53798), .B(n53799), .Z(n53797) );
  XOR U53710 ( .A(n53796), .B(n53800), .Z(n53798) );
  XNOR U53711 ( .A(n53801), .B(n53768), .Z(n53771) );
  XOR U53712 ( .A(n53802), .B(n53803), .Z(n53768) );
  AND U53713 ( .A(n53804), .B(n53805), .Z(n53803) );
  XNOR U53714 ( .A(n53806), .B(n53807), .Z(n53804) );
  IV U53715 ( .A(n53802), .Z(n53806) );
  XNOR U53716 ( .A(n53808), .B(n53809), .Z(n53801) );
  NOR U53717 ( .A(n53810), .B(n53811), .Z(n53809) );
  XNOR U53718 ( .A(n53808), .B(n53812), .Z(n53810) );
  XNOR U53719 ( .A(n53767), .B(n53774), .Z(n53789) );
  NOR U53720 ( .A(n53729), .B(n53813), .Z(n53774) );
  XOR U53721 ( .A(n53779), .B(n53778), .Z(n53767) );
  XNOR U53722 ( .A(n53814), .B(n53775), .Z(n53778) );
  XOR U53723 ( .A(n53815), .B(n53816), .Z(n53775) );
  AND U53724 ( .A(n53817), .B(n53818), .Z(n53816) );
  XNOR U53725 ( .A(n53819), .B(n53820), .Z(n53817) );
  IV U53726 ( .A(n53815), .Z(n53819) );
  XNOR U53727 ( .A(n53821), .B(n53822), .Z(n53814) );
  NOR U53728 ( .A(n53823), .B(n53824), .Z(n53822) );
  XNOR U53729 ( .A(n53821), .B(n53825), .Z(n53823) );
  XOR U53730 ( .A(n53826), .B(n53827), .Z(n53779) );
  NOR U53731 ( .A(n53828), .B(n53829), .Z(n53827) );
  XNOR U53732 ( .A(n53826), .B(n53830), .Z(n53828) );
  XNOR U53733 ( .A(n53720), .B(n53785), .Z(n53787) );
  XNOR U53734 ( .A(n53831), .B(n53832), .Z(n53720) );
  AND U53735 ( .A(n2146), .B(n53833), .Z(n53832) );
  XNOR U53736 ( .A(n53834), .B(n53835), .Z(n53833) );
  AND U53737 ( .A(n53726), .B(n53729), .Z(n53785) );
  XOR U53738 ( .A(n53836), .B(n53813), .Z(n53729) );
  XNOR U53739 ( .A(p_input[1744]), .B(p_input[2048]), .Z(n53813) );
  XNOR U53740 ( .A(n53800), .B(n53799), .Z(n53836) );
  XNOR U53741 ( .A(n53837), .B(n53807), .Z(n53799) );
  XNOR U53742 ( .A(n53795), .B(n53794), .Z(n53807) );
  XNOR U53743 ( .A(n53838), .B(n53791), .Z(n53794) );
  XNOR U53744 ( .A(p_input[1754]), .B(p_input[2058]), .Z(n53791) );
  XOR U53745 ( .A(p_input[1755]), .B(n29030), .Z(n53838) );
  XOR U53746 ( .A(p_input[1756]), .B(p_input[2060]), .Z(n53795) );
  XOR U53747 ( .A(n53805), .B(n53839), .Z(n53837) );
  IV U53748 ( .A(n53796), .Z(n53839) );
  XOR U53749 ( .A(p_input[1745]), .B(p_input[2049]), .Z(n53796) );
  XNOR U53750 ( .A(n53840), .B(n53812), .Z(n53805) );
  XNOR U53751 ( .A(p_input[1759]), .B(n29033), .Z(n53812) );
  XOR U53752 ( .A(n53802), .B(n53811), .Z(n53840) );
  XOR U53753 ( .A(n53841), .B(n53808), .Z(n53811) );
  XOR U53754 ( .A(p_input[1757]), .B(p_input[2061]), .Z(n53808) );
  XOR U53755 ( .A(p_input[1758]), .B(n29035), .Z(n53841) );
  XOR U53756 ( .A(p_input[1753]), .B(p_input[2057]), .Z(n53802) );
  XOR U53757 ( .A(n53820), .B(n53818), .Z(n53800) );
  XNOR U53758 ( .A(n53842), .B(n53825), .Z(n53818) );
  XOR U53759 ( .A(p_input[1752]), .B(p_input[2056]), .Z(n53825) );
  XOR U53760 ( .A(n53815), .B(n53824), .Z(n53842) );
  XOR U53761 ( .A(n53843), .B(n53821), .Z(n53824) );
  XOR U53762 ( .A(p_input[1750]), .B(p_input[2054]), .Z(n53821) );
  XOR U53763 ( .A(p_input[1751]), .B(n30404), .Z(n53843) );
  XOR U53764 ( .A(p_input[1746]), .B(p_input[2050]), .Z(n53815) );
  XNOR U53765 ( .A(n53830), .B(n53829), .Z(n53820) );
  XOR U53766 ( .A(n53844), .B(n53826), .Z(n53829) );
  XOR U53767 ( .A(p_input[1747]), .B(p_input[2051]), .Z(n53826) );
  XOR U53768 ( .A(p_input[1748]), .B(n30406), .Z(n53844) );
  XOR U53769 ( .A(p_input[1749]), .B(p_input[2053]), .Z(n53830) );
  XNOR U53770 ( .A(n53845), .B(n53846), .Z(n53726) );
  AND U53771 ( .A(n2146), .B(n53847), .Z(n53846) );
  XNOR U53772 ( .A(n53848), .B(n53849), .Z(n2146) );
  AND U53773 ( .A(n53850), .B(n53851), .Z(n53849) );
  XOR U53774 ( .A(n53740), .B(n53848), .Z(n53851) );
  XNOR U53775 ( .A(n53852), .B(n53848), .Z(n53850) );
  XOR U53776 ( .A(n53853), .B(n53854), .Z(n53848) );
  AND U53777 ( .A(n53855), .B(n53856), .Z(n53854) );
  XOR U53778 ( .A(n53755), .B(n53853), .Z(n53856) );
  XOR U53779 ( .A(n53853), .B(n53756), .Z(n53855) );
  XOR U53780 ( .A(n53857), .B(n53858), .Z(n53853) );
  AND U53781 ( .A(n53859), .B(n53860), .Z(n53858) );
  XOR U53782 ( .A(n53783), .B(n53857), .Z(n53860) );
  XOR U53783 ( .A(n53857), .B(n53784), .Z(n53859) );
  XOR U53784 ( .A(n53861), .B(n53862), .Z(n53857) );
  AND U53785 ( .A(n53863), .B(n53864), .Z(n53862) );
  XOR U53786 ( .A(n53861), .B(n53834), .Z(n53864) );
  XNOR U53787 ( .A(n53865), .B(n53866), .Z(n53686) );
  AND U53788 ( .A(n2150), .B(n53867), .Z(n53866) );
  XNOR U53789 ( .A(n53868), .B(n53869), .Z(n2150) );
  AND U53790 ( .A(n53870), .B(n53871), .Z(n53869) );
  XOR U53791 ( .A(n53868), .B(n53696), .Z(n53871) );
  XNOR U53792 ( .A(n53868), .B(n53656), .Z(n53870) );
  XOR U53793 ( .A(n53872), .B(n53873), .Z(n53868) );
  AND U53794 ( .A(n53874), .B(n53875), .Z(n53873) );
  XOR U53795 ( .A(n53872), .B(n53664), .Z(n53874) );
  XOR U53796 ( .A(n53876), .B(n53877), .Z(n53647) );
  AND U53797 ( .A(n2154), .B(n53867), .Z(n53877) );
  XNOR U53798 ( .A(n53865), .B(n53876), .Z(n53867) );
  XNOR U53799 ( .A(n53878), .B(n53879), .Z(n2154) );
  AND U53800 ( .A(n53880), .B(n53881), .Z(n53879) );
  XNOR U53801 ( .A(n53882), .B(n53878), .Z(n53881) );
  IV U53802 ( .A(n53696), .Z(n53882) );
  XOR U53803 ( .A(n53852), .B(n53883), .Z(n53696) );
  AND U53804 ( .A(n2157), .B(n53884), .Z(n53883) );
  XOR U53805 ( .A(n53739), .B(n53736), .Z(n53884) );
  IV U53806 ( .A(n53852), .Z(n53739) );
  XNOR U53807 ( .A(n53656), .B(n53878), .Z(n53880) );
  XOR U53808 ( .A(n53885), .B(n53886), .Z(n53656) );
  AND U53809 ( .A(n2173), .B(n53887), .Z(n53886) );
  XOR U53810 ( .A(n53872), .B(n53888), .Z(n53878) );
  AND U53811 ( .A(n53889), .B(n53875), .Z(n53888) );
  XNOR U53812 ( .A(n53706), .B(n53872), .Z(n53875) );
  XOR U53813 ( .A(n53756), .B(n53890), .Z(n53706) );
  AND U53814 ( .A(n2157), .B(n53891), .Z(n53890) );
  XOR U53815 ( .A(n53752), .B(n53756), .Z(n53891) );
  XNOR U53816 ( .A(n53892), .B(n53872), .Z(n53889) );
  IV U53817 ( .A(n53664), .Z(n53892) );
  XOR U53818 ( .A(n53893), .B(n53894), .Z(n53664) );
  AND U53819 ( .A(n2173), .B(n53895), .Z(n53894) );
  XOR U53820 ( .A(n53896), .B(n53897), .Z(n53872) );
  AND U53821 ( .A(n53898), .B(n53899), .Z(n53897) );
  XNOR U53822 ( .A(n53716), .B(n53896), .Z(n53899) );
  XOR U53823 ( .A(n53784), .B(n53900), .Z(n53716) );
  AND U53824 ( .A(n2157), .B(n53901), .Z(n53900) );
  XOR U53825 ( .A(n53780), .B(n53784), .Z(n53901) );
  XOR U53826 ( .A(n53896), .B(n53673), .Z(n53898) );
  XOR U53827 ( .A(n53902), .B(n53903), .Z(n53673) );
  AND U53828 ( .A(n2173), .B(n53904), .Z(n53903) );
  XOR U53829 ( .A(n53905), .B(n53906), .Z(n53896) );
  AND U53830 ( .A(n53907), .B(n53908), .Z(n53906) );
  XNOR U53831 ( .A(n53905), .B(n53724), .Z(n53908) );
  XOR U53832 ( .A(n53835), .B(n53909), .Z(n53724) );
  AND U53833 ( .A(n2157), .B(n53910), .Z(n53909) );
  XOR U53834 ( .A(n53831), .B(n53835), .Z(n53910) );
  XNOR U53835 ( .A(n53911), .B(n53905), .Z(n53907) );
  IV U53836 ( .A(n53683), .Z(n53911) );
  XOR U53837 ( .A(n53912), .B(n53913), .Z(n53683) );
  AND U53838 ( .A(n2173), .B(n53914), .Z(n53913) );
  AND U53839 ( .A(n53876), .B(n53865), .Z(n53905) );
  XNOR U53840 ( .A(n53915), .B(n53916), .Z(n53865) );
  AND U53841 ( .A(n2157), .B(n53847), .Z(n53916) );
  XNOR U53842 ( .A(n53845), .B(n53915), .Z(n53847) );
  XNOR U53843 ( .A(n53917), .B(n53918), .Z(n2157) );
  AND U53844 ( .A(n53919), .B(n53920), .Z(n53918) );
  XNOR U53845 ( .A(n53917), .B(n53736), .Z(n53920) );
  IV U53846 ( .A(n53740), .Z(n53736) );
  XOR U53847 ( .A(n53921), .B(n53922), .Z(n53740) );
  AND U53848 ( .A(n2161), .B(n53923), .Z(n53922) );
  XOR U53849 ( .A(n53924), .B(n53921), .Z(n53923) );
  XNOR U53850 ( .A(n53917), .B(n53852), .Z(n53919) );
  XOR U53851 ( .A(n53925), .B(n53926), .Z(n53852) );
  AND U53852 ( .A(n2169), .B(n53887), .Z(n53926) );
  XOR U53853 ( .A(n53885), .B(n53925), .Z(n53887) );
  XOR U53854 ( .A(n53927), .B(n53928), .Z(n53917) );
  AND U53855 ( .A(n53929), .B(n53930), .Z(n53928) );
  XNOR U53856 ( .A(n53927), .B(n53752), .Z(n53930) );
  IV U53857 ( .A(n53755), .Z(n53752) );
  XOR U53858 ( .A(n53931), .B(n53932), .Z(n53755) );
  AND U53859 ( .A(n2161), .B(n53933), .Z(n53932) );
  XOR U53860 ( .A(n53934), .B(n53931), .Z(n53933) );
  XOR U53861 ( .A(n53756), .B(n53927), .Z(n53929) );
  XOR U53862 ( .A(n53935), .B(n53936), .Z(n53756) );
  AND U53863 ( .A(n2169), .B(n53895), .Z(n53936) );
  XOR U53864 ( .A(n53935), .B(n53893), .Z(n53895) );
  XOR U53865 ( .A(n53937), .B(n53938), .Z(n53927) );
  AND U53866 ( .A(n53939), .B(n53940), .Z(n53938) );
  XNOR U53867 ( .A(n53937), .B(n53780), .Z(n53940) );
  IV U53868 ( .A(n53783), .Z(n53780) );
  XOR U53869 ( .A(n53941), .B(n53942), .Z(n53783) );
  AND U53870 ( .A(n2161), .B(n53943), .Z(n53942) );
  XNOR U53871 ( .A(n53944), .B(n53941), .Z(n53943) );
  XOR U53872 ( .A(n53784), .B(n53937), .Z(n53939) );
  XOR U53873 ( .A(n53945), .B(n53946), .Z(n53784) );
  AND U53874 ( .A(n2169), .B(n53904), .Z(n53946) );
  XOR U53875 ( .A(n53945), .B(n53902), .Z(n53904) );
  XOR U53876 ( .A(n53861), .B(n53947), .Z(n53937) );
  AND U53877 ( .A(n53863), .B(n53948), .Z(n53947) );
  XNOR U53878 ( .A(n53861), .B(n53831), .Z(n53948) );
  IV U53879 ( .A(n53834), .Z(n53831) );
  XOR U53880 ( .A(n53949), .B(n53950), .Z(n53834) );
  AND U53881 ( .A(n2161), .B(n53951), .Z(n53950) );
  XOR U53882 ( .A(n53952), .B(n53949), .Z(n53951) );
  XOR U53883 ( .A(n53835), .B(n53861), .Z(n53863) );
  XOR U53884 ( .A(n53953), .B(n53954), .Z(n53835) );
  AND U53885 ( .A(n2169), .B(n53914), .Z(n53954) );
  XOR U53886 ( .A(n53953), .B(n53912), .Z(n53914) );
  AND U53887 ( .A(n53915), .B(n53845), .Z(n53861) );
  XNOR U53888 ( .A(n53955), .B(n53956), .Z(n53845) );
  AND U53889 ( .A(n2161), .B(n53957), .Z(n53956) );
  XNOR U53890 ( .A(n53958), .B(n53955), .Z(n53957) );
  XNOR U53891 ( .A(n53959), .B(n53960), .Z(n2161) );
  AND U53892 ( .A(n53961), .B(n53962), .Z(n53960) );
  XOR U53893 ( .A(n53924), .B(n53959), .Z(n53962) );
  AND U53894 ( .A(n53963), .B(n53964), .Z(n53924) );
  XNOR U53895 ( .A(n53921), .B(n53959), .Z(n53961) );
  XNOR U53896 ( .A(n53965), .B(n53966), .Z(n53921) );
  AND U53897 ( .A(n2165), .B(n53967), .Z(n53966) );
  XNOR U53898 ( .A(n53968), .B(n53969), .Z(n53967) );
  XOR U53899 ( .A(n53970), .B(n53971), .Z(n53959) );
  AND U53900 ( .A(n53972), .B(n53973), .Z(n53971) );
  XNOR U53901 ( .A(n53970), .B(n53963), .Z(n53973) );
  IV U53902 ( .A(n53934), .Z(n53963) );
  XOR U53903 ( .A(n53974), .B(n53975), .Z(n53934) );
  XOR U53904 ( .A(n53976), .B(n53964), .Z(n53975) );
  AND U53905 ( .A(n53944), .B(n53977), .Z(n53964) );
  AND U53906 ( .A(n53978), .B(n53979), .Z(n53976) );
  XOR U53907 ( .A(n53980), .B(n53974), .Z(n53978) );
  XNOR U53908 ( .A(n53931), .B(n53970), .Z(n53972) );
  XNOR U53909 ( .A(n53981), .B(n53982), .Z(n53931) );
  AND U53910 ( .A(n2165), .B(n53983), .Z(n53982) );
  XNOR U53911 ( .A(n53984), .B(n53985), .Z(n53983) );
  XOR U53912 ( .A(n53986), .B(n53987), .Z(n53970) );
  AND U53913 ( .A(n53988), .B(n53989), .Z(n53987) );
  XNOR U53914 ( .A(n53986), .B(n53944), .Z(n53989) );
  XOR U53915 ( .A(n53990), .B(n53979), .Z(n53944) );
  XNOR U53916 ( .A(n53991), .B(n53974), .Z(n53979) );
  XOR U53917 ( .A(n53992), .B(n53993), .Z(n53974) );
  AND U53918 ( .A(n53994), .B(n53995), .Z(n53993) );
  XOR U53919 ( .A(n53996), .B(n53992), .Z(n53994) );
  XNOR U53920 ( .A(n53997), .B(n53998), .Z(n53991) );
  AND U53921 ( .A(n53999), .B(n54000), .Z(n53998) );
  XOR U53922 ( .A(n53997), .B(n54001), .Z(n53999) );
  XNOR U53923 ( .A(n53980), .B(n53977), .Z(n53990) );
  AND U53924 ( .A(n54002), .B(n54003), .Z(n53977) );
  XOR U53925 ( .A(n54004), .B(n54005), .Z(n53980) );
  AND U53926 ( .A(n54006), .B(n54007), .Z(n54005) );
  XOR U53927 ( .A(n54004), .B(n54008), .Z(n54006) );
  XNOR U53928 ( .A(n53941), .B(n53986), .Z(n53988) );
  XNOR U53929 ( .A(n54009), .B(n54010), .Z(n53941) );
  AND U53930 ( .A(n2165), .B(n54011), .Z(n54010) );
  XNOR U53931 ( .A(n54012), .B(n54013), .Z(n54011) );
  XOR U53932 ( .A(n54014), .B(n54015), .Z(n53986) );
  AND U53933 ( .A(n54016), .B(n54017), .Z(n54015) );
  XNOR U53934 ( .A(n54014), .B(n54002), .Z(n54017) );
  IV U53935 ( .A(n53952), .Z(n54002) );
  XNOR U53936 ( .A(n54018), .B(n53995), .Z(n53952) );
  XNOR U53937 ( .A(n54019), .B(n54001), .Z(n53995) );
  XNOR U53938 ( .A(n54020), .B(n54021), .Z(n54001) );
  NOR U53939 ( .A(n54022), .B(n54023), .Z(n54021) );
  XOR U53940 ( .A(n54020), .B(n54024), .Z(n54022) );
  XNOR U53941 ( .A(n54000), .B(n53992), .Z(n54019) );
  XOR U53942 ( .A(n54025), .B(n54026), .Z(n53992) );
  AND U53943 ( .A(n54027), .B(n54028), .Z(n54026) );
  XOR U53944 ( .A(n54025), .B(n54029), .Z(n54027) );
  XNOR U53945 ( .A(n54030), .B(n53997), .Z(n54000) );
  XOR U53946 ( .A(n54031), .B(n54032), .Z(n53997) );
  AND U53947 ( .A(n54033), .B(n54034), .Z(n54032) );
  XNOR U53948 ( .A(n54035), .B(n54036), .Z(n54033) );
  IV U53949 ( .A(n54031), .Z(n54035) );
  XNOR U53950 ( .A(n54037), .B(n54038), .Z(n54030) );
  NOR U53951 ( .A(n54039), .B(n54040), .Z(n54038) );
  XNOR U53952 ( .A(n54037), .B(n54041), .Z(n54039) );
  XNOR U53953 ( .A(n53996), .B(n54003), .Z(n54018) );
  NOR U53954 ( .A(n53958), .B(n54042), .Z(n54003) );
  XOR U53955 ( .A(n54008), .B(n54007), .Z(n53996) );
  XNOR U53956 ( .A(n54043), .B(n54004), .Z(n54007) );
  XOR U53957 ( .A(n54044), .B(n54045), .Z(n54004) );
  AND U53958 ( .A(n54046), .B(n54047), .Z(n54045) );
  XNOR U53959 ( .A(n54048), .B(n54049), .Z(n54046) );
  IV U53960 ( .A(n54044), .Z(n54048) );
  XNOR U53961 ( .A(n54050), .B(n54051), .Z(n54043) );
  NOR U53962 ( .A(n54052), .B(n54053), .Z(n54051) );
  XNOR U53963 ( .A(n54050), .B(n54054), .Z(n54052) );
  XOR U53964 ( .A(n54055), .B(n54056), .Z(n54008) );
  NOR U53965 ( .A(n54057), .B(n54058), .Z(n54056) );
  XNOR U53966 ( .A(n54055), .B(n54059), .Z(n54057) );
  XNOR U53967 ( .A(n53949), .B(n54014), .Z(n54016) );
  XNOR U53968 ( .A(n54060), .B(n54061), .Z(n53949) );
  AND U53969 ( .A(n2165), .B(n54062), .Z(n54061) );
  XNOR U53970 ( .A(n54063), .B(n54064), .Z(n54062) );
  AND U53971 ( .A(n53955), .B(n53958), .Z(n54014) );
  XOR U53972 ( .A(n54065), .B(n54042), .Z(n53958) );
  XNOR U53973 ( .A(p_input[1760]), .B(p_input[2048]), .Z(n54042) );
  XNOR U53974 ( .A(n54029), .B(n54028), .Z(n54065) );
  XNOR U53975 ( .A(n54066), .B(n54036), .Z(n54028) );
  XNOR U53976 ( .A(n54024), .B(n54023), .Z(n54036) );
  XNOR U53977 ( .A(n54067), .B(n54020), .Z(n54023) );
  XNOR U53978 ( .A(p_input[1770]), .B(p_input[2058]), .Z(n54020) );
  XOR U53979 ( .A(p_input[1771]), .B(n29030), .Z(n54067) );
  XOR U53980 ( .A(p_input[1772]), .B(p_input[2060]), .Z(n54024) );
  XOR U53981 ( .A(n54034), .B(n54068), .Z(n54066) );
  IV U53982 ( .A(n54025), .Z(n54068) );
  XOR U53983 ( .A(p_input[1761]), .B(p_input[2049]), .Z(n54025) );
  XNOR U53984 ( .A(n54069), .B(n54041), .Z(n54034) );
  XNOR U53985 ( .A(p_input[1775]), .B(n29033), .Z(n54041) );
  XOR U53986 ( .A(n54031), .B(n54040), .Z(n54069) );
  XOR U53987 ( .A(n54070), .B(n54037), .Z(n54040) );
  XOR U53988 ( .A(p_input[1773]), .B(p_input[2061]), .Z(n54037) );
  XOR U53989 ( .A(p_input[1774]), .B(n29035), .Z(n54070) );
  XOR U53990 ( .A(p_input[1769]), .B(p_input[2057]), .Z(n54031) );
  XOR U53991 ( .A(n54049), .B(n54047), .Z(n54029) );
  XNOR U53992 ( .A(n54071), .B(n54054), .Z(n54047) );
  XOR U53993 ( .A(p_input[1768]), .B(p_input[2056]), .Z(n54054) );
  XOR U53994 ( .A(n54044), .B(n54053), .Z(n54071) );
  XOR U53995 ( .A(n54072), .B(n54050), .Z(n54053) );
  XOR U53996 ( .A(p_input[1766]), .B(p_input[2054]), .Z(n54050) );
  XOR U53997 ( .A(p_input[1767]), .B(n30404), .Z(n54072) );
  XOR U53998 ( .A(p_input[1762]), .B(p_input[2050]), .Z(n54044) );
  XNOR U53999 ( .A(n54059), .B(n54058), .Z(n54049) );
  XOR U54000 ( .A(n54073), .B(n54055), .Z(n54058) );
  XOR U54001 ( .A(p_input[1763]), .B(p_input[2051]), .Z(n54055) );
  XOR U54002 ( .A(p_input[1764]), .B(n30406), .Z(n54073) );
  XOR U54003 ( .A(p_input[1765]), .B(p_input[2053]), .Z(n54059) );
  XNOR U54004 ( .A(n54074), .B(n54075), .Z(n53955) );
  AND U54005 ( .A(n2165), .B(n54076), .Z(n54075) );
  XNOR U54006 ( .A(n54077), .B(n54078), .Z(n2165) );
  AND U54007 ( .A(n54079), .B(n54080), .Z(n54078) );
  XOR U54008 ( .A(n53969), .B(n54077), .Z(n54080) );
  XNOR U54009 ( .A(n54081), .B(n54077), .Z(n54079) );
  XOR U54010 ( .A(n54082), .B(n54083), .Z(n54077) );
  AND U54011 ( .A(n54084), .B(n54085), .Z(n54083) );
  XOR U54012 ( .A(n53984), .B(n54082), .Z(n54085) );
  XOR U54013 ( .A(n54082), .B(n53985), .Z(n54084) );
  XOR U54014 ( .A(n54086), .B(n54087), .Z(n54082) );
  AND U54015 ( .A(n54088), .B(n54089), .Z(n54087) );
  XOR U54016 ( .A(n54012), .B(n54086), .Z(n54089) );
  XOR U54017 ( .A(n54086), .B(n54013), .Z(n54088) );
  XOR U54018 ( .A(n54090), .B(n54091), .Z(n54086) );
  AND U54019 ( .A(n54092), .B(n54093), .Z(n54091) );
  XOR U54020 ( .A(n54090), .B(n54063), .Z(n54093) );
  XNOR U54021 ( .A(n54094), .B(n54095), .Z(n53915) );
  AND U54022 ( .A(n2169), .B(n54096), .Z(n54095) );
  XNOR U54023 ( .A(n54097), .B(n54098), .Z(n2169) );
  AND U54024 ( .A(n54099), .B(n54100), .Z(n54098) );
  XOR U54025 ( .A(n54097), .B(n53925), .Z(n54100) );
  XNOR U54026 ( .A(n54097), .B(n53885), .Z(n54099) );
  XOR U54027 ( .A(n54101), .B(n54102), .Z(n54097) );
  AND U54028 ( .A(n54103), .B(n54104), .Z(n54102) );
  XOR U54029 ( .A(n54101), .B(n53893), .Z(n54103) );
  XOR U54030 ( .A(n54105), .B(n54106), .Z(n53876) );
  AND U54031 ( .A(n2173), .B(n54096), .Z(n54106) );
  XNOR U54032 ( .A(n54094), .B(n54105), .Z(n54096) );
  XNOR U54033 ( .A(n54107), .B(n54108), .Z(n2173) );
  AND U54034 ( .A(n54109), .B(n54110), .Z(n54108) );
  XNOR U54035 ( .A(n54111), .B(n54107), .Z(n54110) );
  IV U54036 ( .A(n53925), .Z(n54111) );
  XOR U54037 ( .A(n54081), .B(n54112), .Z(n53925) );
  AND U54038 ( .A(n2176), .B(n54113), .Z(n54112) );
  XOR U54039 ( .A(n53968), .B(n53965), .Z(n54113) );
  IV U54040 ( .A(n54081), .Z(n53968) );
  XNOR U54041 ( .A(n53885), .B(n54107), .Z(n54109) );
  XOR U54042 ( .A(n54114), .B(n54115), .Z(n53885) );
  AND U54043 ( .A(n2192), .B(n54116), .Z(n54115) );
  XOR U54044 ( .A(n54101), .B(n54117), .Z(n54107) );
  AND U54045 ( .A(n54118), .B(n54104), .Z(n54117) );
  XNOR U54046 ( .A(n53935), .B(n54101), .Z(n54104) );
  XOR U54047 ( .A(n53985), .B(n54119), .Z(n53935) );
  AND U54048 ( .A(n2176), .B(n54120), .Z(n54119) );
  XOR U54049 ( .A(n53981), .B(n53985), .Z(n54120) );
  XNOR U54050 ( .A(n54121), .B(n54101), .Z(n54118) );
  IV U54051 ( .A(n53893), .Z(n54121) );
  XOR U54052 ( .A(n54122), .B(n54123), .Z(n53893) );
  AND U54053 ( .A(n2192), .B(n54124), .Z(n54123) );
  XOR U54054 ( .A(n54125), .B(n54126), .Z(n54101) );
  AND U54055 ( .A(n54127), .B(n54128), .Z(n54126) );
  XNOR U54056 ( .A(n53945), .B(n54125), .Z(n54128) );
  XOR U54057 ( .A(n54013), .B(n54129), .Z(n53945) );
  AND U54058 ( .A(n2176), .B(n54130), .Z(n54129) );
  XOR U54059 ( .A(n54009), .B(n54013), .Z(n54130) );
  XOR U54060 ( .A(n54125), .B(n53902), .Z(n54127) );
  XOR U54061 ( .A(n54131), .B(n54132), .Z(n53902) );
  AND U54062 ( .A(n2192), .B(n54133), .Z(n54132) );
  XOR U54063 ( .A(n54134), .B(n54135), .Z(n54125) );
  AND U54064 ( .A(n54136), .B(n54137), .Z(n54135) );
  XNOR U54065 ( .A(n54134), .B(n53953), .Z(n54137) );
  XOR U54066 ( .A(n54064), .B(n54138), .Z(n53953) );
  AND U54067 ( .A(n2176), .B(n54139), .Z(n54138) );
  XOR U54068 ( .A(n54060), .B(n54064), .Z(n54139) );
  XNOR U54069 ( .A(n54140), .B(n54134), .Z(n54136) );
  IV U54070 ( .A(n53912), .Z(n54140) );
  XOR U54071 ( .A(n54141), .B(n54142), .Z(n53912) );
  AND U54072 ( .A(n2192), .B(n54143), .Z(n54142) );
  AND U54073 ( .A(n54105), .B(n54094), .Z(n54134) );
  XNOR U54074 ( .A(n54144), .B(n54145), .Z(n54094) );
  AND U54075 ( .A(n2176), .B(n54076), .Z(n54145) );
  XNOR U54076 ( .A(n54074), .B(n54144), .Z(n54076) );
  XNOR U54077 ( .A(n54146), .B(n54147), .Z(n2176) );
  AND U54078 ( .A(n54148), .B(n54149), .Z(n54147) );
  XNOR U54079 ( .A(n54146), .B(n53965), .Z(n54149) );
  IV U54080 ( .A(n53969), .Z(n53965) );
  XOR U54081 ( .A(n54150), .B(n54151), .Z(n53969) );
  AND U54082 ( .A(n2180), .B(n54152), .Z(n54151) );
  XOR U54083 ( .A(n54153), .B(n54150), .Z(n54152) );
  XNOR U54084 ( .A(n54146), .B(n54081), .Z(n54148) );
  XOR U54085 ( .A(n54154), .B(n54155), .Z(n54081) );
  AND U54086 ( .A(n2188), .B(n54116), .Z(n54155) );
  XOR U54087 ( .A(n54114), .B(n54154), .Z(n54116) );
  XOR U54088 ( .A(n54156), .B(n54157), .Z(n54146) );
  AND U54089 ( .A(n54158), .B(n54159), .Z(n54157) );
  XNOR U54090 ( .A(n54156), .B(n53981), .Z(n54159) );
  IV U54091 ( .A(n53984), .Z(n53981) );
  XOR U54092 ( .A(n54160), .B(n54161), .Z(n53984) );
  AND U54093 ( .A(n2180), .B(n54162), .Z(n54161) );
  XOR U54094 ( .A(n54163), .B(n54160), .Z(n54162) );
  XOR U54095 ( .A(n53985), .B(n54156), .Z(n54158) );
  XOR U54096 ( .A(n54164), .B(n54165), .Z(n53985) );
  AND U54097 ( .A(n2188), .B(n54124), .Z(n54165) );
  XOR U54098 ( .A(n54164), .B(n54122), .Z(n54124) );
  XOR U54099 ( .A(n54166), .B(n54167), .Z(n54156) );
  AND U54100 ( .A(n54168), .B(n54169), .Z(n54167) );
  XNOR U54101 ( .A(n54166), .B(n54009), .Z(n54169) );
  IV U54102 ( .A(n54012), .Z(n54009) );
  XOR U54103 ( .A(n54170), .B(n54171), .Z(n54012) );
  AND U54104 ( .A(n2180), .B(n54172), .Z(n54171) );
  XNOR U54105 ( .A(n54173), .B(n54170), .Z(n54172) );
  XOR U54106 ( .A(n54013), .B(n54166), .Z(n54168) );
  XOR U54107 ( .A(n54174), .B(n54175), .Z(n54013) );
  AND U54108 ( .A(n2188), .B(n54133), .Z(n54175) );
  XOR U54109 ( .A(n54174), .B(n54131), .Z(n54133) );
  XOR U54110 ( .A(n54090), .B(n54176), .Z(n54166) );
  AND U54111 ( .A(n54092), .B(n54177), .Z(n54176) );
  XNOR U54112 ( .A(n54090), .B(n54060), .Z(n54177) );
  IV U54113 ( .A(n54063), .Z(n54060) );
  XOR U54114 ( .A(n54178), .B(n54179), .Z(n54063) );
  AND U54115 ( .A(n2180), .B(n54180), .Z(n54179) );
  XOR U54116 ( .A(n54181), .B(n54178), .Z(n54180) );
  XOR U54117 ( .A(n54064), .B(n54090), .Z(n54092) );
  XOR U54118 ( .A(n54182), .B(n54183), .Z(n54064) );
  AND U54119 ( .A(n2188), .B(n54143), .Z(n54183) );
  XOR U54120 ( .A(n54182), .B(n54141), .Z(n54143) );
  AND U54121 ( .A(n54144), .B(n54074), .Z(n54090) );
  XNOR U54122 ( .A(n54184), .B(n54185), .Z(n54074) );
  AND U54123 ( .A(n2180), .B(n54186), .Z(n54185) );
  XNOR U54124 ( .A(n54187), .B(n54184), .Z(n54186) );
  XNOR U54125 ( .A(n54188), .B(n54189), .Z(n2180) );
  AND U54126 ( .A(n54190), .B(n54191), .Z(n54189) );
  XOR U54127 ( .A(n54153), .B(n54188), .Z(n54191) );
  AND U54128 ( .A(n54192), .B(n54193), .Z(n54153) );
  XNOR U54129 ( .A(n54150), .B(n54188), .Z(n54190) );
  XNOR U54130 ( .A(n54194), .B(n54195), .Z(n54150) );
  AND U54131 ( .A(n2184), .B(n54196), .Z(n54195) );
  XNOR U54132 ( .A(n54197), .B(n54198), .Z(n54196) );
  XOR U54133 ( .A(n54199), .B(n54200), .Z(n54188) );
  AND U54134 ( .A(n54201), .B(n54202), .Z(n54200) );
  XNOR U54135 ( .A(n54199), .B(n54192), .Z(n54202) );
  IV U54136 ( .A(n54163), .Z(n54192) );
  XOR U54137 ( .A(n54203), .B(n54204), .Z(n54163) );
  XOR U54138 ( .A(n54205), .B(n54193), .Z(n54204) );
  AND U54139 ( .A(n54173), .B(n54206), .Z(n54193) );
  AND U54140 ( .A(n54207), .B(n54208), .Z(n54205) );
  XOR U54141 ( .A(n54209), .B(n54203), .Z(n54207) );
  XNOR U54142 ( .A(n54160), .B(n54199), .Z(n54201) );
  XNOR U54143 ( .A(n54210), .B(n54211), .Z(n54160) );
  AND U54144 ( .A(n2184), .B(n54212), .Z(n54211) );
  XNOR U54145 ( .A(n54213), .B(n54214), .Z(n54212) );
  XOR U54146 ( .A(n54215), .B(n54216), .Z(n54199) );
  AND U54147 ( .A(n54217), .B(n54218), .Z(n54216) );
  XNOR U54148 ( .A(n54215), .B(n54173), .Z(n54218) );
  XOR U54149 ( .A(n54219), .B(n54208), .Z(n54173) );
  XNOR U54150 ( .A(n54220), .B(n54203), .Z(n54208) );
  XOR U54151 ( .A(n54221), .B(n54222), .Z(n54203) );
  AND U54152 ( .A(n54223), .B(n54224), .Z(n54222) );
  XOR U54153 ( .A(n54225), .B(n54221), .Z(n54223) );
  XNOR U54154 ( .A(n54226), .B(n54227), .Z(n54220) );
  AND U54155 ( .A(n54228), .B(n54229), .Z(n54227) );
  XOR U54156 ( .A(n54226), .B(n54230), .Z(n54228) );
  XNOR U54157 ( .A(n54209), .B(n54206), .Z(n54219) );
  AND U54158 ( .A(n54231), .B(n54232), .Z(n54206) );
  XOR U54159 ( .A(n54233), .B(n54234), .Z(n54209) );
  AND U54160 ( .A(n54235), .B(n54236), .Z(n54234) );
  XOR U54161 ( .A(n54233), .B(n54237), .Z(n54235) );
  XNOR U54162 ( .A(n54170), .B(n54215), .Z(n54217) );
  XNOR U54163 ( .A(n54238), .B(n54239), .Z(n54170) );
  AND U54164 ( .A(n2184), .B(n54240), .Z(n54239) );
  XNOR U54165 ( .A(n54241), .B(n54242), .Z(n54240) );
  XOR U54166 ( .A(n54243), .B(n54244), .Z(n54215) );
  AND U54167 ( .A(n54245), .B(n54246), .Z(n54244) );
  XNOR U54168 ( .A(n54243), .B(n54231), .Z(n54246) );
  IV U54169 ( .A(n54181), .Z(n54231) );
  XNOR U54170 ( .A(n54247), .B(n54224), .Z(n54181) );
  XNOR U54171 ( .A(n54248), .B(n54230), .Z(n54224) );
  XNOR U54172 ( .A(n54249), .B(n54250), .Z(n54230) );
  NOR U54173 ( .A(n54251), .B(n54252), .Z(n54250) );
  XOR U54174 ( .A(n54249), .B(n54253), .Z(n54251) );
  XNOR U54175 ( .A(n54229), .B(n54221), .Z(n54248) );
  XOR U54176 ( .A(n54254), .B(n54255), .Z(n54221) );
  AND U54177 ( .A(n54256), .B(n54257), .Z(n54255) );
  XOR U54178 ( .A(n54254), .B(n54258), .Z(n54256) );
  XNOR U54179 ( .A(n54259), .B(n54226), .Z(n54229) );
  XOR U54180 ( .A(n54260), .B(n54261), .Z(n54226) );
  AND U54181 ( .A(n54262), .B(n54263), .Z(n54261) );
  XNOR U54182 ( .A(n54264), .B(n54265), .Z(n54262) );
  IV U54183 ( .A(n54260), .Z(n54264) );
  XNOR U54184 ( .A(n54266), .B(n54267), .Z(n54259) );
  NOR U54185 ( .A(n54268), .B(n54269), .Z(n54267) );
  XNOR U54186 ( .A(n54266), .B(n54270), .Z(n54268) );
  XNOR U54187 ( .A(n54225), .B(n54232), .Z(n54247) );
  NOR U54188 ( .A(n54187), .B(n54271), .Z(n54232) );
  XOR U54189 ( .A(n54237), .B(n54236), .Z(n54225) );
  XNOR U54190 ( .A(n54272), .B(n54233), .Z(n54236) );
  XOR U54191 ( .A(n54273), .B(n54274), .Z(n54233) );
  AND U54192 ( .A(n54275), .B(n54276), .Z(n54274) );
  XNOR U54193 ( .A(n54277), .B(n54278), .Z(n54275) );
  IV U54194 ( .A(n54273), .Z(n54277) );
  XNOR U54195 ( .A(n54279), .B(n54280), .Z(n54272) );
  NOR U54196 ( .A(n54281), .B(n54282), .Z(n54280) );
  XNOR U54197 ( .A(n54279), .B(n54283), .Z(n54281) );
  XOR U54198 ( .A(n54284), .B(n54285), .Z(n54237) );
  NOR U54199 ( .A(n54286), .B(n54287), .Z(n54285) );
  XNOR U54200 ( .A(n54284), .B(n54288), .Z(n54286) );
  XNOR U54201 ( .A(n54178), .B(n54243), .Z(n54245) );
  XNOR U54202 ( .A(n54289), .B(n54290), .Z(n54178) );
  AND U54203 ( .A(n2184), .B(n54291), .Z(n54290) );
  XNOR U54204 ( .A(n54292), .B(n54293), .Z(n54291) );
  AND U54205 ( .A(n54184), .B(n54187), .Z(n54243) );
  XOR U54206 ( .A(n54294), .B(n54271), .Z(n54187) );
  XNOR U54207 ( .A(p_input[1776]), .B(p_input[2048]), .Z(n54271) );
  XNOR U54208 ( .A(n54258), .B(n54257), .Z(n54294) );
  XNOR U54209 ( .A(n54295), .B(n54265), .Z(n54257) );
  XNOR U54210 ( .A(n54253), .B(n54252), .Z(n54265) );
  XNOR U54211 ( .A(n54296), .B(n54249), .Z(n54252) );
  XNOR U54212 ( .A(p_input[1786]), .B(p_input[2058]), .Z(n54249) );
  XOR U54213 ( .A(p_input[1787]), .B(n29030), .Z(n54296) );
  XOR U54214 ( .A(p_input[1788]), .B(p_input[2060]), .Z(n54253) );
  XOR U54215 ( .A(n54263), .B(n54297), .Z(n54295) );
  IV U54216 ( .A(n54254), .Z(n54297) );
  XOR U54217 ( .A(p_input[1777]), .B(p_input[2049]), .Z(n54254) );
  XNOR U54218 ( .A(n54298), .B(n54270), .Z(n54263) );
  XNOR U54219 ( .A(p_input[1791]), .B(n29033), .Z(n54270) );
  XOR U54220 ( .A(n54260), .B(n54269), .Z(n54298) );
  XOR U54221 ( .A(n54299), .B(n54266), .Z(n54269) );
  XOR U54222 ( .A(p_input[1789]), .B(p_input[2061]), .Z(n54266) );
  XOR U54223 ( .A(p_input[1790]), .B(n29035), .Z(n54299) );
  XOR U54224 ( .A(p_input[1785]), .B(p_input[2057]), .Z(n54260) );
  XOR U54225 ( .A(n54278), .B(n54276), .Z(n54258) );
  XNOR U54226 ( .A(n54300), .B(n54283), .Z(n54276) );
  XOR U54227 ( .A(p_input[1784]), .B(p_input[2056]), .Z(n54283) );
  XOR U54228 ( .A(n54273), .B(n54282), .Z(n54300) );
  XOR U54229 ( .A(n54301), .B(n54279), .Z(n54282) );
  XOR U54230 ( .A(p_input[1782]), .B(p_input[2054]), .Z(n54279) );
  XOR U54231 ( .A(p_input[1783]), .B(n30404), .Z(n54301) );
  XOR U54232 ( .A(p_input[1778]), .B(p_input[2050]), .Z(n54273) );
  XNOR U54233 ( .A(n54288), .B(n54287), .Z(n54278) );
  XOR U54234 ( .A(n54302), .B(n54284), .Z(n54287) );
  XOR U54235 ( .A(p_input[1779]), .B(p_input[2051]), .Z(n54284) );
  XOR U54236 ( .A(p_input[1780]), .B(n30406), .Z(n54302) );
  XOR U54237 ( .A(p_input[1781]), .B(p_input[2053]), .Z(n54288) );
  XNOR U54238 ( .A(n54303), .B(n54304), .Z(n54184) );
  AND U54239 ( .A(n2184), .B(n54305), .Z(n54304) );
  XNOR U54240 ( .A(n54306), .B(n54307), .Z(n2184) );
  AND U54241 ( .A(n54308), .B(n54309), .Z(n54307) );
  XOR U54242 ( .A(n54198), .B(n54306), .Z(n54309) );
  XNOR U54243 ( .A(n54310), .B(n54306), .Z(n54308) );
  XOR U54244 ( .A(n54311), .B(n54312), .Z(n54306) );
  AND U54245 ( .A(n54313), .B(n54314), .Z(n54312) );
  XOR U54246 ( .A(n54213), .B(n54311), .Z(n54314) );
  XOR U54247 ( .A(n54311), .B(n54214), .Z(n54313) );
  XOR U54248 ( .A(n54315), .B(n54316), .Z(n54311) );
  AND U54249 ( .A(n54317), .B(n54318), .Z(n54316) );
  XOR U54250 ( .A(n54241), .B(n54315), .Z(n54318) );
  XOR U54251 ( .A(n54315), .B(n54242), .Z(n54317) );
  XOR U54252 ( .A(n54319), .B(n54320), .Z(n54315) );
  AND U54253 ( .A(n54321), .B(n54322), .Z(n54320) );
  XOR U54254 ( .A(n54319), .B(n54292), .Z(n54322) );
  XNOR U54255 ( .A(n54323), .B(n54324), .Z(n54144) );
  AND U54256 ( .A(n2188), .B(n54325), .Z(n54324) );
  XNOR U54257 ( .A(n54326), .B(n54327), .Z(n2188) );
  AND U54258 ( .A(n54328), .B(n54329), .Z(n54327) );
  XOR U54259 ( .A(n54326), .B(n54154), .Z(n54329) );
  XNOR U54260 ( .A(n54326), .B(n54114), .Z(n54328) );
  XOR U54261 ( .A(n54330), .B(n54331), .Z(n54326) );
  AND U54262 ( .A(n54332), .B(n54333), .Z(n54331) );
  XOR U54263 ( .A(n54330), .B(n54122), .Z(n54332) );
  XOR U54264 ( .A(n54334), .B(n54335), .Z(n54105) );
  AND U54265 ( .A(n2192), .B(n54325), .Z(n54335) );
  XNOR U54266 ( .A(n54323), .B(n54334), .Z(n54325) );
  XNOR U54267 ( .A(n54336), .B(n54337), .Z(n2192) );
  AND U54268 ( .A(n54338), .B(n54339), .Z(n54337) );
  XNOR U54269 ( .A(n54340), .B(n54336), .Z(n54339) );
  IV U54270 ( .A(n54154), .Z(n54340) );
  XOR U54271 ( .A(n54310), .B(n54341), .Z(n54154) );
  AND U54272 ( .A(n2195), .B(n54342), .Z(n54341) );
  XOR U54273 ( .A(n54197), .B(n54194), .Z(n54342) );
  IV U54274 ( .A(n54310), .Z(n54197) );
  XNOR U54275 ( .A(n54114), .B(n54336), .Z(n54338) );
  XOR U54276 ( .A(n54343), .B(n54344), .Z(n54114) );
  AND U54277 ( .A(n2211), .B(n54345), .Z(n54344) );
  XOR U54278 ( .A(n54330), .B(n54346), .Z(n54336) );
  AND U54279 ( .A(n54347), .B(n54333), .Z(n54346) );
  XNOR U54280 ( .A(n54164), .B(n54330), .Z(n54333) );
  XOR U54281 ( .A(n54214), .B(n54348), .Z(n54164) );
  AND U54282 ( .A(n2195), .B(n54349), .Z(n54348) );
  XOR U54283 ( .A(n54210), .B(n54214), .Z(n54349) );
  XNOR U54284 ( .A(n54350), .B(n54330), .Z(n54347) );
  IV U54285 ( .A(n54122), .Z(n54350) );
  XOR U54286 ( .A(n54351), .B(n54352), .Z(n54122) );
  AND U54287 ( .A(n2211), .B(n54353), .Z(n54352) );
  XOR U54288 ( .A(n54354), .B(n54355), .Z(n54330) );
  AND U54289 ( .A(n54356), .B(n54357), .Z(n54355) );
  XNOR U54290 ( .A(n54174), .B(n54354), .Z(n54357) );
  XOR U54291 ( .A(n54242), .B(n54358), .Z(n54174) );
  AND U54292 ( .A(n2195), .B(n54359), .Z(n54358) );
  XOR U54293 ( .A(n54238), .B(n54242), .Z(n54359) );
  XOR U54294 ( .A(n54354), .B(n54131), .Z(n54356) );
  XOR U54295 ( .A(n54360), .B(n54361), .Z(n54131) );
  AND U54296 ( .A(n2211), .B(n54362), .Z(n54361) );
  XOR U54297 ( .A(n54363), .B(n54364), .Z(n54354) );
  AND U54298 ( .A(n54365), .B(n54366), .Z(n54364) );
  XNOR U54299 ( .A(n54363), .B(n54182), .Z(n54366) );
  XOR U54300 ( .A(n54293), .B(n54367), .Z(n54182) );
  AND U54301 ( .A(n2195), .B(n54368), .Z(n54367) );
  XOR U54302 ( .A(n54289), .B(n54293), .Z(n54368) );
  XNOR U54303 ( .A(n54369), .B(n54363), .Z(n54365) );
  IV U54304 ( .A(n54141), .Z(n54369) );
  XOR U54305 ( .A(n54370), .B(n54371), .Z(n54141) );
  AND U54306 ( .A(n2211), .B(n54372), .Z(n54371) );
  AND U54307 ( .A(n54334), .B(n54323), .Z(n54363) );
  XNOR U54308 ( .A(n54373), .B(n54374), .Z(n54323) );
  AND U54309 ( .A(n2195), .B(n54305), .Z(n54374) );
  XNOR U54310 ( .A(n54303), .B(n54373), .Z(n54305) );
  XNOR U54311 ( .A(n54375), .B(n54376), .Z(n2195) );
  AND U54312 ( .A(n54377), .B(n54378), .Z(n54376) );
  XNOR U54313 ( .A(n54375), .B(n54194), .Z(n54378) );
  IV U54314 ( .A(n54198), .Z(n54194) );
  XOR U54315 ( .A(n54379), .B(n54380), .Z(n54198) );
  AND U54316 ( .A(n2199), .B(n54381), .Z(n54380) );
  XOR U54317 ( .A(n54382), .B(n54379), .Z(n54381) );
  XNOR U54318 ( .A(n54375), .B(n54310), .Z(n54377) );
  XOR U54319 ( .A(n54383), .B(n54384), .Z(n54310) );
  AND U54320 ( .A(n2207), .B(n54345), .Z(n54384) );
  XOR U54321 ( .A(n54343), .B(n54383), .Z(n54345) );
  XOR U54322 ( .A(n54385), .B(n54386), .Z(n54375) );
  AND U54323 ( .A(n54387), .B(n54388), .Z(n54386) );
  XNOR U54324 ( .A(n54385), .B(n54210), .Z(n54388) );
  IV U54325 ( .A(n54213), .Z(n54210) );
  XOR U54326 ( .A(n54389), .B(n54390), .Z(n54213) );
  AND U54327 ( .A(n2199), .B(n54391), .Z(n54390) );
  XOR U54328 ( .A(n54392), .B(n54389), .Z(n54391) );
  XOR U54329 ( .A(n54214), .B(n54385), .Z(n54387) );
  XOR U54330 ( .A(n54393), .B(n54394), .Z(n54214) );
  AND U54331 ( .A(n2207), .B(n54353), .Z(n54394) );
  XOR U54332 ( .A(n54393), .B(n54351), .Z(n54353) );
  XOR U54333 ( .A(n54395), .B(n54396), .Z(n54385) );
  AND U54334 ( .A(n54397), .B(n54398), .Z(n54396) );
  XNOR U54335 ( .A(n54395), .B(n54238), .Z(n54398) );
  IV U54336 ( .A(n54241), .Z(n54238) );
  XOR U54337 ( .A(n54399), .B(n54400), .Z(n54241) );
  AND U54338 ( .A(n2199), .B(n54401), .Z(n54400) );
  XNOR U54339 ( .A(n54402), .B(n54399), .Z(n54401) );
  XOR U54340 ( .A(n54242), .B(n54395), .Z(n54397) );
  XOR U54341 ( .A(n54403), .B(n54404), .Z(n54242) );
  AND U54342 ( .A(n2207), .B(n54362), .Z(n54404) );
  XOR U54343 ( .A(n54403), .B(n54360), .Z(n54362) );
  XOR U54344 ( .A(n54319), .B(n54405), .Z(n54395) );
  AND U54345 ( .A(n54321), .B(n54406), .Z(n54405) );
  XNOR U54346 ( .A(n54319), .B(n54289), .Z(n54406) );
  IV U54347 ( .A(n54292), .Z(n54289) );
  XOR U54348 ( .A(n54407), .B(n54408), .Z(n54292) );
  AND U54349 ( .A(n2199), .B(n54409), .Z(n54408) );
  XOR U54350 ( .A(n54410), .B(n54407), .Z(n54409) );
  XOR U54351 ( .A(n54293), .B(n54319), .Z(n54321) );
  XOR U54352 ( .A(n54411), .B(n54412), .Z(n54293) );
  AND U54353 ( .A(n2207), .B(n54372), .Z(n54412) );
  XOR U54354 ( .A(n54411), .B(n54370), .Z(n54372) );
  AND U54355 ( .A(n54373), .B(n54303), .Z(n54319) );
  XNOR U54356 ( .A(n54413), .B(n54414), .Z(n54303) );
  AND U54357 ( .A(n2199), .B(n54415), .Z(n54414) );
  XNOR U54358 ( .A(n54416), .B(n54413), .Z(n54415) );
  XNOR U54359 ( .A(n54417), .B(n54418), .Z(n2199) );
  AND U54360 ( .A(n54419), .B(n54420), .Z(n54418) );
  XOR U54361 ( .A(n54382), .B(n54417), .Z(n54420) );
  AND U54362 ( .A(n54421), .B(n54422), .Z(n54382) );
  XNOR U54363 ( .A(n54379), .B(n54417), .Z(n54419) );
  XNOR U54364 ( .A(n54423), .B(n54424), .Z(n54379) );
  AND U54365 ( .A(n2203), .B(n54425), .Z(n54424) );
  XNOR U54366 ( .A(n54426), .B(n54427), .Z(n54425) );
  XOR U54367 ( .A(n54428), .B(n54429), .Z(n54417) );
  AND U54368 ( .A(n54430), .B(n54431), .Z(n54429) );
  XNOR U54369 ( .A(n54428), .B(n54421), .Z(n54431) );
  IV U54370 ( .A(n54392), .Z(n54421) );
  XOR U54371 ( .A(n54432), .B(n54433), .Z(n54392) );
  XOR U54372 ( .A(n54434), .B(n54422), .Z(n54433) );
  AND U54373 ( .A(n54402), .B(n54435), .Z(n54422) );
  AND U54374 ( .A(n54436), .B(n54437), .Z(n54434) );
  XOR U54375 ( .A(n54438), .B(n54432), .Z(n54436) );
  XNOR U54376 ( .A(n54389), .B(n54428), .Z(n54430) );
  XNOR U54377 ( .A(n54439), .B(n54440), .Z(n54389) );
  AND U54378 ( .A(n2203), .B(n54441), .Z(n54440) );
  XNOR U54379 ( .A(n54442), .B(n54443), .Z(n54441) );
  XOR U54380 ( .A(n54444), .B(n54445), .Z(n54428) );
  AND U54381 ( .A(n54446), .B(n54447), .Z(n54445) );
  XNOR U54382 ( .A(n54444), .B(n54402), .Z(n54447) );
  XOR U54383 ( .A(n54448), .B(n54437), .Z(n54402) );
  XNOR U54384 ( .A(n54449), .B(n54432), .Z(n54437) );
  XOR U54385 ( .A(n54450), .B(n54451), .Z(n54432) );
  AND U54386 ( .A(n54452), .B(n54453), .Z(n54451) );
  XOR U54387 ( .A(n54454), .B(n54450), .Z(n54452) );
  XNOR U54388 ( .A(n54455), .B(n54456), .Z(n54449) );
  AND U54389 ( .A(n54457), .B(n54458), .Z(n54456) );
  XOR U54390 ( .A(n54455), .B(n54459), .Z(n54457) );
  XNOR U54391 ( .A(n54438), .B(n54435), .Z(n54448) );
  AND U54392 ( .A(n54460), .B(n54461), .Z(n54435) );
  XOR U54393 ( .A(n54462), .B(n54463), .Z(n54438) );
  AND U54394 ( .A(n54464), .B(n54465), .Z(n54463) );
  XOR U54395 ( .A(n54462), .B(n54466), .Z(n54464) );
  XNOR U54396 ( .A(n54399), .B(n54444), .Z(n54446) );
  XNOR U54397 ( .A(n54467), .B(n54468), .Z(n54399) );
  AND U54398 ( .A(n2203), .B(n54469), .Z(n54468) );
  XNOR U54399 ( .A(n54470), .B(n54471), .Z(n54469) );
  XOR U54400 ( .A(n54472), .B(n54473), .Z(n54444) );
  AND U54401 ( .A(n54474), .B(n54475), .Z(n54473) );
  XNOR U54402 ( .A(n54472), .B(n54460), .Z(n54475) );
  IV U54403 ( .A(n54410), .Z(n54460) );
  XNOR U54404 ( .A(n54476), .B(n54453), .Z(n54410) );
  XNOR U54405 ( .A(n54477), .B(n54459), .Z(n54453) );
  XNOR U54406 ( .A(n54478), .B(n54479), .Z(n54459) );
  NOR U54407 ( .A(n54480), .B(n54481), .Z(n54479) );
  XOR U54408 ( .A(n54478), .B(n54482), .Z(n54480) );
  XNOR U54409 ( .A(n54458), .B(n54450), .Z(n54477) );
  XOR U54410 ( .A(n54483), .B(n54484), .Z(n54450) );
  AND U54411 ( .A(n54485), .B(n54486), .Z(n54484) );
  XOR U54412 ( .A(n54483), .B(n54487), .Z(n54485) );
  XNOR U54413 ( .A(n54488), .B(n54455), .Z(n54458) );
  XOR U54414 ( .A(n54489), .B(n54490), .Z(n54455) );
  AND U54415 ( .A(n54491), .B(n54492), .Z(n54490) );
  XNOR U54416 ( .A(n54493), .B(n54494), .Z(n54491) );
  IV U54417 ( .A(n54489), .Z(n54493) );
  XNOR U54418 ( .A(n54495), .B(n54496), .Z(n54488) );
  NOR U54419 ( .A(n54497), .B(n54498), .Z(n54496) );
  XNOR U54420 ( .A(n54495), .B(n54499), .Z(n54497) );
  XNOR U54421 ( .A(n54454), .B(n54461), .Z(n54476) );
  NOR U54422 ( .A(n54416), .B(n54500), .Z(n54461) );
  XOR U54423 ( .A(n54466), .B(n54465), .Z(n54454) );
  XNOR U54424 ( .A(n54501), .B(n54462), .Z(n54465) );
  XOR U54425 ( .A(n54502), .B(n54503), .Z(n54462) );
  AND U54426 ( .A(n54504), .B(n54505), .Z(n54503) );
  XNOR U54427 ( .A(n54506), .B(n54507), .Z(n54504) );
  IV U54428 ( .A(n54502), .Z(n54506) );
  XNOR U54429 ( .A(n54508), .B(n54509), .Z(n54501) );
  NOR U54430 ( .A(n54510), .B(n54511), .Z(n54509) );
  XNOR U54431 ( .A(n54508), .B(n54512), .Z(n54510) );
  XOR U54432 ( .A(n54513), .B(n54514), .Z(n54466) );
  NOR U54433 ( .A(n54515), .B(n54516), .Z(n54514) );
  XNOR U54434 ( .A(n54513), .B(n54517), .Z(n54515) );
  XNOR U54435 ( .A(n54407), .B(n54472), .Z(n54474) );
  XNOR U54436 ( .A(n54518), .B(n54519), .Z(n54407) );
  AND U54437 ( .A(n2203), .B(n54520), .Z(n54519) );
  XNOR U54438 ( .A(n54521), .B(n54522), .Z(n54520) );
  AND U54439 ( .A(n54413), .B(n54416), .Z(n54472) );
  XOR U54440 ( .A(n54523), .B(n54500), .Z(n54416) );
  XNOR U54441 ( .A(p_input[1792]), .B(p_input[2048]), .Z(n54500) );
  XNOR U54442 ( .A(n54487), .B(n54486), .Z(n54523) );
  XNOR U54443 ( .A(n54524), .B(n54494), .Z(n54486) );
  XNOR U54444 ( .A(n54482), .B(n54481), .Z(n54494) );
  XNOR U54445 ( .A(n54525), .B(n54478), .Z(n54481) );
  XNOR U54446 ( .A(p_input[1802]), .B(p_input[2058]), .Z(n54478) );
  XOR U54447 ( .A(p_input[1803]), .B(n29030), .Z(n54525) );
  XOR U54448 ( .A(p_input[1804]), .B(p_input[2060]), .Z(n54482) );
  XOR U54449 ( .A(n54492), .B(n54526), .Z(n54524) );
  IV U54450 ( .A(n54483), .Z(n54526) );
  XOR U54451 ( .A(p_input[1793]), .B(p_input[2049]), .Z(n54483) );
  XNOR U54452 ( .A(n54527), .B(n54499), .Z(n54492) );
  XNOR U54453 ( .A(p_input[1807]), .B(n29033), .Z(n54499) );
  XOR U54454 ( .A(n54489), .B(n54498), .Z(n54527) );
  XOR U54455 ( .A(n54528), .B(n54495), .Z(n54498) );
  XOR U54456 ( .A(p_input[1805]), .B(p_input[2061]), .Z(n54495) );
  XOR U54457 ( .A(p_input[1806]), .B(n29035), .Z(n54528) );
  XOR U54458 ( .A(p_input[1801]), .B(p_input[2057]), .Z(n54489) );
  XOR U54459 ( .A(n54507), .B(n54505), .Z(n54487) );
  XNOR U54460 ( .A(n54529), .B(n54512), .Z(n54505) );
  XOR U54461 ( .A(p_input[1800]), .B(p_input[2056]), .Z(n54512) );
  XOR U54462 ( .A(n54502), .B(n54511), .Z(n54529) );
  XOR U54463 ( .A(n54530), .B(n54508), .Z(n54511) );
  XOR U54464 ( .A(p_input[1798]), .B(p_input[2054]), .Z(n54508) );
  XOR U54465 ( .A(p_input[1799]), .B(n30404), .Z(n54530) );
  XOR U54466 ( .A(p_input[1794]), .B(p_input[2050]), .Z(n54502) );
  XNOR U54467 ( .A(n54517), .B(n54516), .Z(n54507) );
  XOR U54468 ( .A(n54531), .B(n54513), .Z(n54516) );
  XOR U54469 ( .A(p_input[1795]), .B(p_input[2051]), .Z(n54513) );
  XOR U54470 ( .A(p_input[1796]), .B(n30406), .Z(n54531) );
  XOR U54471 ( .A(p_input[1797]), .B(p_input[2053]), .Z(n54517) );
  XNOR U54472 ( .A(n54532), .B(n54533), .Z(n54413) );
  AND U54473 ( .A(n2203), .B(n54534), .Z(n54533) );
  XNOR U54474 ( .A(n54535), .B(n54536), .Z(n2203) );
  AND U54475 ( .A(n54537), .B(n54538), .Z(n54536) );
  XOR U54476 ( .A(n54427), .B(n54535), .Z(n54538) );
  XNOR U54477 ( .A(n54539), .B(n54535), .Z(n54537) );
  XOR U54478 ( .A(n54540), .B(n54541), .Z(n54535) );
  AND U54479 ( .A(n54542), .B(n54543), .Z(n54541) );
  XOR U54480 ( .A(n54442), .B(n54540), .Z(n54543) );
  XOR U54481 ( .A(n54540), .B(n54443), .Z(n54542) );
  XOR U54482 ( .A(n54544), .B(n54545), .Z(n54540) );
  AND U54483 ( .A(n54546), .B(n54547), .Z(n54545) );
  XOR U54484 ( .A(n54470), .B(n54544), .Z(n54547) );
  XOR U54485 ( .A(n54544), .B(n54471), .Z(n54546) );
  XOR U54486 ( .A(n54548), .B(n54549), .Z(n54544) );
  AND U54487 ( .A(n54550), .B(n54551), .Z(n54549) );
  XOR U54488 ( .A(n54548), .B(n54521), .Z(n54551) );
  XNOR U54489 ( .A(n54552), .B(n54553), .Z(n54373) );
  AND U54490 ( .A(n2207), .B(n54554), .Z(n54553) );
  XNOR U54491 ( .A(n54555), .B(n54556), .Z(n2207) );
  AND U54492 ( .A(n54557), .B(n54558), .Z(n54556) );
  XOR U54493 ( .A(n54555), .B(n54383), .Z(n54558) );
  XNOR U54494 ( .A(n54555), .B(n54343), .Z(n54557) );
  XOR U54495 ( .A(n54559), .B(n54560), .Z(n54555) );
  AND U54496 ( .A(n54561), .B(n54562), .Z(n54560) );
  XOR U54497 ( .A(n54559), .B(n54351), .Z(n54561) );
  XOR U54498 ( .A(n54563), .B(n54564), .Z(n54334) );
  AND U54499 ( .A(n2211), .B(n54554), .Z(n54564) );
  XNOR U54500 ( .A(n54552), .B(n54563), .Z(n54554) );
  XNOR U54501 ( .A(n54565), .B(n54566), .Z(n2211) );
  AND U54502 ( .A(n54567), .B(n54568), .Z(n54566) );
  XNOR U54503 ( .A(n54569), .B(n54565), .Z(n54568) );
  IV U54504 ( .A(n54383), .Z(n54569) );
  XOR U54505 ( .A(n54539), .B(n54570), .Z(n54383) );
  AND U54506 ( .A(n2214), .B(n54571), .Z(n54570) );
  XOR U54507 ( .A(n54426), .B(n54423), .Z(n54571) );
  IV U54508 ( .A(n54539), .Z(n54426) );
  XNOR U54509 ( .A(n54343), .B(n54565), .Z(n54567) );
  XOR U54510 ( .A(n54572), .B(n54573), .Z(n54343) );
  AND U54511 ( .A(n2230), .B(n54574), .Z(n54573) );
  XOR U54512 ( .A(n54559), .B(n54575), .Z(n54565) );
  AND U54513 ( .A(n54576), .B(n54562), .Z(n54575) );
  XNOR U54514 ( .A(n54393), .B(n54559), .Z(n54562) );
  XOR U54515 ( .A(n54443), .B(n54577), .Z(n54393) );
  AND U54516 ( .A(n2214), .B(n54578), .Z(n54577) );
  XOR U54517 ( .A(n54439), .B(n54443), .Z(n54578) );
  XNOR U54518 ( .A(n54579), .B(n54559), .Z(n54576) );
  IV U54519 ( .A(n54351), .Z(n54579) );
  XOR U54520 ( .A(n54580), .B(n54581), .Z(n54351) );
  AND U54521 ( .A(n2230), .B(n54582), .Z(n54581) );
  XOR U54522 ( .A(n54583), .B(n54584), .Z(n54559) );
  AND U54523 ( .A(n54585), .B(n54586), .Z(n54584) );
  XNOR U54524 ( .A(n54403), .B(n54583), .Z(n54586) );
  XOR U54525 ( .A(n54471), .B(n54587), .Z(n54403) );
  AND U54526 ( .A(n2214), .B(n54588), .Z(n54587) );
  XOR U54527 ( .A(n54467), .B(n54471), .Z(n54588) );
  XOR U54528 ( .A(n54583), .B(n54360), .Z(n54585) );
  XOR U54529 ( .A(n54589), .B(n54590), .Z(n54360) );
  AND U54530 ( .A(n2230), .B(n54591), .Z(n54590) );
  XOR U54531 ( .A(n54592), .B(n54593), .Z(n54583) );
  AND U54532 ( .A(n54594), .B(n54595), .Z(n54593) );
  XNOR U54533 ( .A(n54592), .B(n54411), .Z(n54595) );
  XOR U54534 ( .A(n54522), .B(n54596), .Z(n54411) );
  AND U54535 ( .A(n2214), .B(n54597), .Z(n54596) );
  XOR U54536 ( .A(n54518), .B(n54522), .Z(n54597) );
  XNOR U54537 ( .A(n54598), .B(n54592), .Z(n54594) );
  IV U54538 ( .A(n54370), .Z(n54598) );
  XOR U54539 ( .A(n54599), .B(n54600), .Z(n54370) );
  AND U54540 ( .A(n2230), .B(n54601), .Z(n54600) );
  AND U54541 ( .A(n54563), .B(n54552), .Z(n54592) );
  XNOR U54542 ( .A(n54602), .B(n54603), .Z(n54552) );
  AND U54543 ( .A(n2214), .B(n54534), .Z(n54603) );
  XNOR U54544 ( .A(n54532), .B(n54602), .Z(n54534) );
  XNOR U54545 ( .A(n54604), .B(n54605), .Z(n2214) );
  AND U54546 ( .A(n54606), .B(n54607), .Z(n54605) );
  XNOR U54547 ( .A(n54604), .B(n54423), .Z(n54607) );
  IV U54548 ( .A(n54427), .Z(n54423) );
  XOR U54549 ( .A(n54608), .B(n54609), .Z(n54427) );
  AND U54550 ( .A(n2218), .B(n54610), .Z(n54609) );
  XOR U54551 ( .A(n54611), .B(n54608), .Z(n54610) );
  XNOR U54552 ( .A(n54604), .B(n54539), .Z(n54606) );
  XOR U54553 ( .A(n54612), .B(n54613), .Z(n54539) );
  AND U54554 ( .A(n2226), .B(n54574), .Z(n54613) );
  XOR U54555 ( .A(n54572), .B(n54612), .Z(n54574) );
  XOR U54556 ( .A(n54614), .B(n54615), .Z(n54604) );
  AND U54557 ( .A(n54616), .B(n54617), .Z(n54615) );
  XNOR U54558 ( .A(n54614), .B(n54439), .Z(n54617) );
  IV U54559 ( .A(n54442), .Z(n54439) );
  XOR U54560 ( .A(n54618), .B(n54619), .Z(n54442) );
  AND U54561 ( .A(n2218), .B(n54620), .Z(n54619) );
  XOR U54562 ( .A(n54621), .B(n54618), .Z(n54620) );
  XOR U54563 ( .A(n54443), .B(n54614), .Z(n54616) );
  XOR U54564 ( .A(n54622), .B(n54623), .Z(n54443) );
  AND U54565 ( .A(n2226), .B(n54582), .Z(n54623) );
  XOR U54566 ( .A(n54622), .B(n54580), .Z(n54582) );
  XOR U54567 ( .A(n54624), .B(n54625), .Z(n54614) );
  AND U54568 ( .A(n54626), .B(n54627), .Z(n54625) );
  XNOR U54569 ( .A(n54624), .B(n54467), .Z(n54627) );
  IV U54570 ( .A(n54470), .Z(n54467) );
  XOR U54571 ( .A(n54628), .B(n54629), .Z(n54470) );
  AND U54572 ( .A(n2218), .B(n54630), .Z(n54629) );
  XNOR U54573 ( .A(n54631), .B(n54628), .Z(n54630) );
  XOR U54574 ( .A(n54471), .B(n54624), .Z(n54626) );
  XOR U54575 ( .A(n54632), .B(n54633), .Z(n54471) );
  AND U54576 ( .A(n2226), .B(n54591), .Z(n54633) );
  XOR U54577 ( .A(n54632), .B(n54589), .Z(n54591) );
  XOR U54578 ( .A(n54548), .B(n54634), .Z(n54624) );
  AND U54579 ( .A(n54550), .B(n54635), .Z(n54634) );
  XNOR U54580 ( .A(n54548), .B(n54518), .Z(n54635) );
  IV U54581 ( .A(n54521), .Z(n54518) );
  XOR U54582 ( .A(n54636), .B(n54637), .Z(n54521) );
  AND U54583 ( .A(n2218), .B(n54638), .Z(n54637) );
  XOR U54584 ( .A(n54639), .B(n54636), .Z(n54638) );
  XOR U54585 ( .A(n54522), .B(n54548), .Z(n54550) );
  XOR U54586 ( .A(n54640), .B(n54641), .Z(n54522) );
  AND U54587 ( .A(n2226), .B(n54601), .Z(n54641) );
  XOR U54588 ( .A(n54640), .B(n54599), .Z(n54601) );
  AND U54589 ( .A(n54602), .B(n54532), .Z(n54548) );
  XNOR U54590 ( .A(n54642), .B(n54643), .Z(n54532) );
  AND U54591 ( .A(n2218), .B(n54644), .Z(n54643) );
  XNOR U54592 ( .A(n54645), .B(n54642), .Z(n54644) );
  XNOR U54593 ( .A(n54646), .B(n54647), .Z(n2218) );
  AND U54594 ( .A(n54648), .B(n54649), .Z(n54647) );
  XOR U54595 ( .A(n54611), .B(n54646), .Z(n54649) );
  AND U54596 ( .A(n54650), .B(n54651), .Z(n54611) );
  XNOR U54597 ( .A(n54608), .B(n54646), .Z(n54648) );
  XNOR U54598 ( .A(n54652), .B(n54653), .Z(n54608) );
  AND U54599 ( .A(n2222), .B(n54654), .Z(n54653) );
  XNOR U54600 ( .A(n54655), .B(n54656), .Z(n54654) );
  XOR U54601 ( .A(n54657), .B(n54658), .Z(n54646) );
  AND U54602 ( .A(n54659), .B(n54660), .Z(n54658) );
  XNOR U54603 ( .A(n54657), .B(n54650), .Z(n54660) );
  IV U54604 ( .A(n54621), .Z(n54650) );
  XOR U54605 ( .A(n54661), .B(n54662), .Z(n54621) );
  XOR U54606 ( .A(n54663), .B(n54651), .Z(n54662) );
  AND U54607 ( .A(n54631), .B(n54664), .Z(n54651) );
  AND U54608 ( .A(n54665), .B(n54666), .Z(n54663) );
  XOR U54609 ( .A(n54667), .B(n54661), .Z(n54665) );
  XNOR U54610 ( .A(n54618), .B(n54657), .Z(n54659) );
  XNOR U54611 ( .A(n54668), .B(n54669), .Z(n54618) );
  AND U54612 ( .A(n2222), .B(n54670), .Z(n54669) );
  XNOR U54613 ( .A(n54671), .B(n54672), .Z(n54670) );
  XOR U54614 ( .A(n54673), .B(n54674), .Z(n54657) );
  AND U54615 ( .A(n54675), .B(n54676), .Z(n54674) );
  XNOR U54616 ( .A(n54673), .B(n54631), .Z(n54676) );
  XOR U54617 ( .A(n54677), .B(n54666), .Z(n54631) );
  XNOR U54618 ( .A(n54678), .B(n54661), .Z(n54666) );
  XOR U54619 ( .A(n54679), .B(n54680), .Z(n54661) );
  AND U54620 ( .A(n54681), .B(n54682), .Z(n54680) );
  XOR U54621 ( .A(n54683), .B(n54679), .Z(n54681) );
  XNOR U54622 ( .A(n54684), .B(n54685), .Z(n54678) );
  AND U54623 ( .A(n54686), .B(n54687), .Z(n54685) );
  XOR U54624 ( .A(n54684), .B(n54688), .Z(n54686) );
  XNOR U54625 ( .A(n54667), .B(n54664), .Z(n54677) );
  AND U54626 ( .A(n54689), .B(n54690), .Z(n54664) );
  XOR U54627 ( .A(n54691), .B(n54692), .Z(n54667) );
  AND U54628 ( .A(n54693), .B(n54694), .Z(n54692) );
  XOR U54629 ( .A(n54691), .B(n54695), .Z(n54693) );
  XNOR U54630 ( .A(n54628), .B(n54673), .Z(n54675) );
  XNOR U54631 ( .A(n54696), .B(n54697), .Z(n54628) );
  AND U54632 ( .A(n2222), .B(n54698), .Z(n54697) );
  XNOR U54633 ( .A(n54699), .B(n54700), .Z(n54698) );
  XOR U54634 ( .A(n54701), .B(n54702), .Z(n54673) );
  AND U54635 ( .A(n54703), .B(n54704), .Z(n54702) );
  XNOR U54636 ( .A(n54701), .B(n54689), .Z(n54704) );
  IV U54637 ( .A(n54639), .Z(n54689) );
  XNOR U54638 ( .A(n54705), .B(n54682), .Z(n54639) );
  XNOR U54639 ( .A(n54706), .B(n54688), .Z(n54682) );
  XNOR U54640 ( .A(n54707), .B(n54708), .Z(n54688) );
  NOR U54641 ( .A(n54709), .B(n54710), .Z(n54708) );
  XOR U54642 ( .A(n54707), .B(n54711), .Z(n54709) );
  XNOR U54643 ( .A(n54687), .B(n54679), .Z(n54706) );
  XOR U54644 ( .A(n54712), .B(n54713), .Z(n54679) );
  AND U54645 ( .A(n54714), .B(n54715), .Z(n54713) );
  XOR U54646 ( .A(n54712), .B(n54716), .Z(n54714) );
  XNOR U54647 ( .A(n54717), .B(n54684), .Z(n54687) );
  XOR U54648 ( .A(n54718), .B(n54719), .Z(n54684) );
  AND U54649 ( .A(n54720), .B(n54721), .Z(n54719) );
  XNOR U54650 ( .A(n54722), .B(n54723), .Z(n54720) );
  IV U54651 ( .A(n54718), .Z(n54722) );
  XNOR U54652 ( .A(n54724), .B(n54725), .Z(n54717) );
  NOR U54653 ( .A(n54726), .B(n54727), .Z(n54725) );
  XNOR U54654 ( .A(n54724), .B(n54728), .Z(n54726) );
  XNOR U54655 ( .A(n54683), .B(n54690), .Z(n54705) );
  NOR U54656 ( .A(n54645), .B(n54729), .Z(n54690) );
  XOR U54657 ( .A(n54695), .B(n54694), .Z(n54683) );
  XNOR U54658 ( .A(n54730), .B(n54691), .Z(n54694) );
  XOR U54659 ( .A(n54731), .B(n54732), .Z(n54691) );
  AND U54660 ( .A(n54733), .B(n54734), .Z(n54732) );
  XNOR U54661 ( .A(n54735), .B(n54736), .Z(n54733) );
  IV U54662 ( .A(n54731), .Z(n54735) );
  XNOR U54663 ( .A(n54737), .B(n54738), .Z(n54730) );
  NOR U54664 ( .A(n54739), .B(n54740), .Z(n54738) );
  XNOR U54665 ( .A(n54737), .B(n54741), .Z(n54739) );
  XOR U54666 ( .A(n54742), .B(n54743), .Z(n54695) );
  NOR U54667 ( .A(n54744), .B(n54745), .Z(n54743) );
  XNOR U54668 ( .A(n54742), .B(n54746), .Z(n54744) );
  XNOR U54669 ( .A(n54636), .B(n54701), .Z(n54703) );
  XNOR U54670 ( .A(n54747), .B(n54748), .Z(n54636) );
  AND U54671 ( .A(n2222), .B(n54749), .Z(n54748) );
  XNOR U54672 ( .A(n54750), .B(n54751), .Z(n54749) );
  AND U54673 ( .A(n54642), .B(n54645), .Z(n54701) );
  XOR U54674 ( .A(n54752), .B(n54729), .Z(n54645) );
  XNOR U54675 ( .A(p_input[1808]), .B(p_input[2048]), .Z(n54729) );
  XNOR U54676 ( .A(n54716), .B(n54715), .Z(n54752) );
  XNOR U54677 ( .A(n54753), .B(n54723), .Z(n54715) );
  XNOR U54678 ( .A(n54711), .B(n54710), .Z(n54723) );
  XNOR U54679 ( .A(n54754), .B(n54707), .Z(n54710) );
  XNOR U54680 ( .A(p_input[1818]), .B(p_input[2058]), .Z(n54707) );
  XOR U54681 ( .A(p_input[1819]), .B(n29030), .Z(n54754) );
  XOR U54682 ( .A(p_input[1820]), .B(p_input[2060]), .Z(n54711) );
  XOR U54683 ( .A(n54721), .B(n54755), .Z(n54753) );
  IV U54684 ( .A(n54712), .Z(n54755) );
  XOR U54685 ( .A(p_input[1809]), .B(p_input[2049]), .Z(n54712) );
  XNOR U54686 ( .A(n54756), .B(n54728), .Z(n54721) );
  XNOR U54687 ( .A(p_input[1823]), .B(n29033), .Z(n54728) );
  XOR U54688 ( .A(n54718), .B(n54727), .Z(n54756) );
  XOR U54689 ( .A(n54757), .B(n54724), .Z(n54727) );
  XOR U54690 ( .A(p_input[1821]), .B(p_input[2061]), .Z(n54724) );
  XOR U54691 ( .A(p_input[1822]), .B(n29035), .Z(n54757) );
  XOR U54692 ( .A(p_input[1817]), .B(p_input[2057]), .Z(n54718) );
  XOR U54693 ( .A(n54736), .B(n54734), .Z(n54716) );
  XNOR U54694 ( .A(n54758), .B(n54741), .Z(n54734) );
  XOR U54695 ( .A(p_input[1816]), .B(p_input[2056]), .Z(n54741) );
  XOR U54696 ( .A(n54731), .B(n54740), .Z(n54758) );
  XOR U54697 ( .A(n54759), .B(n54737), .Z(n54740) );
  XOR U54698 ( .A(p_input[1814]), .B(p_input[2054]), .Z(n54737) );
  XOR U54699 ( .A(p_input[1815]), .B(n30404), .Z(n54759) );
  XOR U54700 ( .A(p_input[1810]), .B(p_input[2050]), .Z(n54731) );
  XNOR U54701 ( .A(n54746), .B(n54745), .Z(n54736) );
  XOR U54702 ( .A(n54760), .B(n54742), .Z(n54745) );
  XOR U54703 ( .A(p_input[1811]), .B(p_input[2051]), .Z(n54742) );
  XOR U54704 ( .A(p_input[1812]), .B(n30406), .Z(n54760) );
  XOR U54705 ( .A(p_input[1813]), .B(p_input[2053]), .Z(n54746) );
  XNOR U54706 ( .A(n54761), .B(n54762), .Z(n54642) );
  AND U54707 ( .A(n2222), .B(n54763), .Z(n54762) );
  XNOR U54708 ( .A(n54764), .B(n54765), .Z(n2222) );
  AND U54709 ( .A(n54766), .B(n54767), .Z(n54765) );
  XOR U54710 ( .A(n54656), .B(n54764), .Z(n54767) );
  XNOR U54711 ( .A(n54768), .B(n54764), .Z(n54766) );
  XOR U54712 ( .A(n54769), .B(n54770), .Z(n54764) );
  AND U54713 ( .A(n54771), .B(n54772), .Z(n54770) );
  XOR U54714 ( .A(n54671), .B(n54769), .Z(n54772) );
  XOR U54715 ( .A(n54769), .B(n54672), .Z(n54771) );
  XOR U54716 ( .A(n54773), .B(n54774), .Z(n54769) );
  AND U54717 ( .A(n54775), .B(n54776), .Z(n54774) );
  XOR U54718 ( .A(n54699), .B(n54773), .Z(n54776) );
  XOR U54719 ( .A(n54773), .B(n54700), .Z(n54775) );
  XOR U54720 ( .A(n54777), .B(n54778), .Z(n54773) );
  AND U54721 ( .A(n54779), .B(n54780), .Z(n54778) );
  XOR U54722 ( .A(n54777), .B(n54750), .Z(n54780) );
  XNOR U54723 ( .A(n54781), .B(n54782), .Z(n54602) );
  AND U54724 ( .A(n2226), .B(n54783), .Z(n54782) );
  XNOR U54725 ( .A(n54784), .B(n54785), .Z(n2226) );
  AND U54726 ( .A(n54786), .B(n54787), .Z(n54785) );
  XOR U54727 ( .A(n54784), .B(n54612), .Z(n54787) );
  XNOR U54728 ( .A(n54784), .B(n54572), .Z(n54786) );
  XOR U54729 ( .A(n54788), .B(n54789), .Z(n54784) );
  AND U54730 ( .A(n54790), .B(n54791), .Z(n54789) );
  XOR U54731 ( .A(n54788), .B(n54580), .Z(n54790) );
  XOR U54732 ( .A(n54792), .B(n54793), .Z(n54563) );
  AND U54733 ( .A(n2230), .B(n54783), .Z(n54793) );
  XNOR U54734 ( .A(n54781), .B(n54792), .Z(n54783) );
  XNOR U54735 ( .A(n54794), .B(n54795), .Z(n2230) );
  AND U54736 ( .A(n54796), .B(n54797), .Z(n54795) );
  XNOR U54737 ( .A(n54798), .B(n54794), .Z(n54797) );
  IV U54738 ( .A(n54612), .Z(n54798) );
  XOR U54739 ( .A(n54768), .B(n54799), .Z(n54612) );
  AND U54740 ( .A(n2233), .B(n54800), .Z(n54799) );
  XOR U54741 ( .A(n54655), .B(n54652), .Z(n54800) );
  IV U54742 ( .A(n54768), .Z(n54655) );
  XNOR U54743 ( .A(n54572), .B(n54794), .Z(n54796) );
  XOR U54744 ( .A(n54801), .B(n54802), .Z(n54572) );
  AND U54745 ( .A(n2249), .B(n54803), .Z(n54802) );
  XOR U54746 ( .A(n54788), .B(n54804), .Z(n54794) );
  AND U54747 ( .A(n54805), .B(n54791), .Z(n54804) );
  XNOR U54748 ( .A(n54622), .B(n54788), .Z(n54791) );
  XOR U54749 ( .A(n54672), .B(n54806), .Z(n54622) );
  AND U54750 ( .A(n2233), .B(n54807), .Z(n54806) );
  XOR U54751 ( .A(n54668), .B(n54672), .Z(n54807) );
  XNOR U54752 ( .A(n54808), .B(n54788), .Z(n54805) );
  IV U54753 ( .A(n54580), .Z(n54808) );
  XOR U54754 ( .A(n54809), .B(n54810), .Z(n54580) );
  AND U54755 ( .A(n2249), .B(n54811), .Z(n54810) );
  XOR U54756 ( .A(n54812), .B(n54813), .Z(n54788) );
  AND U54757 ( .A(n54814), .B(n54815), .Z(n54813) );
  XNOR U54758 ( .A(n54632), .B(n54812), .Z(n54815) );
  XOR U54759 ( .A(n54700), .B(n54816), .Z(n54632) );
  AND U54760 ( .A(n2233), .B(n54817), .Z(n54816) );
  XOR U54761 ( .A(n54696), .B(n54700), .Z(n54817) );
  XOR U54762 ( .A(n54812), .B(n54589), .Z(n54814) );
  XOR U54763 ( .A(n54818), .B(n54819), .Z(n54589) );
  AND U54764 ( .A(n2249), .B(n54820), .Z(n54819) );
  XOR U54765 ( .A(n54821), .B(n54822), .Z(n54812) );
  AND U54766 ( .A(n54823), .B(n54824), .Z(n54822) );
  XNOR U54767 ( .A(n54821), .B(n54640), .Z(n54824) );
  XOR U54768 ( .A(n54751), .B(n54825), .Z(n54640) );
  AND U54769 ( .A(n2233), .B(n54826), .Z(n54825) );
  XOR U54770 ( .A(n54747), .B(n54751), .Z(n54826) );
  XNOR U54771 ( .A(n54827), .B(n54821), .Z(n54823) );
  IV U54772 ( .A(n54599), .Z(n54827) );
  XOR U54773 ( .A(n54828), .B(n54829), .Z(n54599) );
  AND U54774 ( .A(n2249), .B(n54830), .Z(n54829) );
  AND U54775 ( .A(n54792), .B(n54781), .Z(n54821) );
  XNOR U54776 ( .A(n54831), .B(n54832), .Z(n54781) );
  AND U54777 ( .A(n2233), .B(n54763), .Z(n54832) );
  XNOR U54778 ( .A(n54761), .B(n54831), .Z(n54763) );
  XNOR U54779 ( .A(n54833), .B(n54834), .Z(n2233) );
  AND U54780 ( .A(n54835), .B(n54836), .Z(n54834) );
  XNOR U54781 ( .A(n54833), .B(n54652), .Z(n54836) );
  IV U54782 ( .A(n54656), .Z(n54652) );
  XOR U54783 ( .A(n54837), .B(n54838), .Z(n54656) );
  AND U54784 ( .A(n2237), .B(n54839), .Z(n54838) );
  XOR U54785 ( .A(n54840), .B(n54837), .Z(n54839) );
  XNOR U54786 ( .A(n54833), .B(n54768), .Z(n54835) );
  XOR U54787 ( .A(n54841), .B(n54842), .Z(n54768) );
  AND U54788 ( .A(n2245), .B(n54803), .Z(n54842) );
  XOR U54789 ( .A(n54801), .B(n54841), .Z(n54803) );
  XOR U54790 ( .A(n54843), .B(n54844), .Z(n54833) );
  AND U54791 ( .A(n54845), .B(n54846), .Z(n54844) );
  XNOR U54792 ( .A(n54843), .B(n54668), .Z(n54846) );
  IV U54793 ( .A(n54671), .Z(n54668) );
  XOR U54794 ( .A(n54847), .B(n54848), .Z(n54671) );
  AND U54795 ( .A(n2237), .B(n54849), .Z(n54848) );
  XOR U54796 ( .A(n54850), .B(n54847), .Z(n54849) );
  XOR U54797 ( .A(n54672), .B(n54843), .Z(n54845) );
  XOR U54798 ( .A(n54851), .B(n54852), .Z(n54672) );
  AND U54799 ( .A(n2245), .B(n54811), .Z(n54852) );
  XOR U54800 ( .A(n54851), .B(n54809), .Z(n54811) );
  XOR U54801 ( .A(n54853), .B(n54854), .Z(n54843) );
  AND U54802 ( .A(n54855), .B(n54856), .Z(n54854) );
  XNOR U54803 ( .A(n54853), .B(n54696), .Z(n54856) );
  IV U54804 ( .A(n54699), .Z(n54696) );
  XOR U54805 ( .A(n54857), .B(n54858), .Z(n54699) );
  AND U54806 ( .A(n2237), .B(n54859), .Z(n54858) );
  XNOR U54807 ( .A(n54860), .B(n54857), .Z(n54859) );
  XOR U54808 ( .A(n54700), .B(n54853), .Z(n54855) );
  XOR U54809 ( .A(n54861), .B(n54862), .Z(n54700) );
  AND U54810 ( .A(n2245), .B(n54820), .Z(n54862) );
  XOR U54811 ( .A(n54861), .B(n54818), .Z(n54820) );
  XOR U54812 ( .A(n54777), .B(n54863), .Z(n54853) );
  AND U54813 ( .A(n54779), .B(n54864), .Z(n54863) );
  XNOR U54814 ( .A(n54777), .B(n54747), .Z(n54864) );
  IV U54815 ( .A(n54750), .Z(n54747) );
  XOR U54816 ( .A(n54865), .B(n54866), .Z(n54750) );
  AND U54817 ( .A(n2237), .B(n54867), .Z(n54866) );
  XOR U54818 ( .A(n54868), .B(n54865), .Z(n54867) );
  XOR U54819 ( .A(n54751), .B(n54777), .Z(n54779) );
  XOR U54820 ( .A(n54869), .B(n54870), .Z(n54751) );
  AND U54821 ( .A(n2245), .B(n54830), .Z(n54870) );
  XOR U54822 ( .A(n54869), .B(n54828), .Z(n54830) );
  AND U54823 ( .A(n54831), .B(n54761), .Z(n54777) );
  XNOR U54824 ( .A(n54871), .B(n54872), .Z(n54761) );
  AND U54825 ( .A(n2237), .B(n54873), .Z(n54872) );
  XNOR U54826 ( .A(n54874), .B(n54871), .Z(n54873) );
  XNOR U54827 ( .A(n54875), .B(n54876), .Z(n2237) );
  AND U54828 ( .A(n54877), .B(n54878), .Z(n54876) );
  XOR U54829 ( .A(n54840), .B(n54875), .Z(n54878) );
  AND U54830 ( .A(n54879), .B(n54880), .Z(n54840) );
  XNOR U54831 ( .A(n54837), .B(n54875), .Z(n54877) );
  XNOR U54832 ( .A(n54881), .B(n54882), .Z(n54837) );
  AND U54833 ( .A(n2241), .B(n54883), .Z(n54882) );
  XNOR U54834 ( .A(n54884), .B(n54885), .Z(n54883) );
  XOR U54835 ( .A(n54886), .B(n54887), .Z(n54875) );
  AND U54836 ( .A(n54888), .B(n54889), .Z(n54887) );
  XNOR U54837 ( .A(n54886), .B(n54879), .Z(n54889) );
  IV U54838 ( .A(n54850), .Z(n54879) );
  XOR U54839 ( .A(n54890), .B(n54891), .Z(n54850) );
  XOR U54840 ( .A(n54892), .B(n54880), .Z(n54891) );
  AND U54841 ( .A(n54860), .B(n54893), .Z(n54880) );
  AND U54842 ( .A(n54894), .B(n54895), .Z(n54892) );
  XOR U54843 ( .A(n54896), .B(n54890), .Z(n54894) );
  XNOR U54844 ( .A(n54847), .B(n54886), .Z(n54888) );
  XNOR U54845 ( .A(n54897), .B(n54898), .Z(n54847) );
  AND U54846 ( .A(n2241), .B(n54899), .Z(n54898) );
  XNOR U54847 ( .A(n54900), .B(n54901), .Z(n54899) );
  XOR U54848 ( .A(n54902), .B(n54903), .Z(n54886) );
  AND U54849 ( .A(n54904), .B(n54905), .Z(n54903) );
  XNOR U54850 ( .A(n54902), .B(n54860), .Z(n54905) );
  XOR U54851 ( .A(n54906), .B(n54895), .Z(n54860) );
  XNOR U54852 ( .A(n54907), .B(n54890), .Z(n54895) );
  XOR U54853 ( .A(n54908), .B(n54909), .Z(n54890) );
  AND U54854 ( .A(n54910), .B(n54911), .Z(n54909) );
  XOR U54855 ( .A(n54912), .B(n54908), .Z(n54910) );
  XNOR U54856 ( .A(n54913), .B(n54914), .Z(n54907) );
  AND U54857 ( .A(n54915), .B(n54916), .Z(n54914) );
  XOR U54858 ( .A(n54913), .B(n54917), .Z(n54915) );
  XNOR U54859 ( .A(n54896), .B(n54893), .Z(n54906) );
  AND U54860 ( .A(n54918), .B(n54919), .Z(n54893) );
  XOR U54861 ( .A(n54920), .B(n54921), .Z(n54896) );
  AND U54862 ( .A(n54922), .B(n54923), .Z(n54921) );
  XOR U54863 ( .A(n54920), .B(n54924), .Z(n54922) );
  XNOR U54864 ( .A(n54857), .B(n54902), .Z(n54904) );
  XNOR U54865 ( .A(n54925), .B(n54926), .Z(n54857) );
  AND U54866 ( .A(n2241), .B(n54927), .Z(n54926) );
  XNOR U54867 ( .A(n54928), .B(n54929), .Z(n54927) );
  XOR U54868 ( .A(n54930), .B(n54931), .Z(n54902) );
  AND U54869 ( .A(n54932), .B(n54933), .Z(n54931) );
  XNOR U54870 ( .A(n54930), .B(n54918), .Z(n54933) );
  IV U54871 ( .A(n54868), .Z(n54918) );
  XNOR U54872 ( .A(n54934), .B(n54911), .Z(n54868) );
  XNOR U54873 ( .A(n54935), .B(n54917), .Z(n54911) );
  XNOR U54874 ( .A(n54936), .B(n54937), .Z(n54917) );
  NOR U54875 ( .A(n54938), .B(n54939), .Z(n54937) );
  XOR U54876 ( .A(n54936), .B(n54940), .Z(n54938) );
  XNOR U54877 ( .A(n54916), .B(n54908), .Z(n54935) );
  XOR U54878 ( .A(n54941), .B(n54942), .Z(n54908) );
  AND U54879 ( .A(n54943), .B(n54944), .Z(n54942) );
  XOR U54880 ( .A(n54941), .B(n54945), .Z(n54943) );
  XNOR U54881 ( .A(n54946), .B(n54913), .Z(n54916) );
  XOR U54882 ( .A(n54947), .B(n54948), .Z(n54913) );
  AND U54883 ( .A(n54949), .B(n54950), .Z(n54948) );
  XNOR U54884 ( .A(n54951), .B(n54952), .Z(n54949) );
  IV U54885 ( .A(n54947), .Z(n54951) );
  XNOR U54886 ( .A(n54953), .B(n54954), .Z(n54946) );
  NOR U54887 ( .A(n54955), .B(n54956), .Z(n54954) );
  XNOR U54888 ( .A(n54953), .B(n54957), .Z(n54955) );
  XNOR U54889 ( .A(n54912), .B(n54919), .Z(n54934) );
  NOR U54890 ( .A(n54874), .B(n54958), .Z(n54919) );
  XOR U54891 ( .A(n54924), .B(n54923), .Z(n54912) );
  XNOR U54892 ( .A(n54959), .B(n54920), .Z(n54923) );
  XOR U54893 ( .A(n54960), .B(n54961), .Z(n54920) );
  AND U54894 ( .A(n54962), .B(n54963), .Z(n54961) );
  XNOR U54895 ( .A(n54964), .B(n54965), .Z(n54962) );
  IV U54896 ( .A(n54960), .Z(n54964) );
  XNOR U54897 ( .A(n54966), .B(n54967), .Z(n54959) );
  NOR U54898 ( .A(n54968), .B(n54969), .Z(n54967) );
  XNOR U54899 ( .A(n54966), .B(n54970), .Z(n54968) );
  XOR U54900 ( .A(n54971), .B(n54972), .Z(n54924) );
  NOR U54901 ( .A(n54973), .B(n54974), .Z(n54972) );
  XNOR U54902 ( .A(n54971), .B(n54975), .Z(n54973) );
  XNOR U54903 ( .A(n54865), .B(n54930), .Z(n54932) );
  XNOR U54904 ( .A(n54976), .B(n54977), .Z(n54865) );
  AND U54905 ( .A(n2241), .B(n54978), .Z(n54977) );
  XNOR U54906 ( .A(n54979), .B(n54980), .Z(n54978) );
  AND U54907 ( .A(n54871), .B(n54874), .Z(n54930) );
  XOR U54908 ( .A(n54981), .B(n54958), .Z(n54874) );
  XNOR U54909 ( .A(p_input[1824]), .B(p_input[2048]), .Z(n54958) );
  XNOR U54910 ( .A(n54945), .B(n54944), .Z(n54981) );
  XNOR U54911 ( .A(n54982), .B(n54952), .Z(n54944) );
  XNOR U54912 ( .A(n54940), .B(n54939), .Z(n54952) );
  XNOR U54913 ( .A(n54983), .B(n54936), .Z(n54939) );
  XNOR U54914 ( .A(p_input[1834]), .B(p_input[2058]), .Z(n54936) );
  XOR U54915 ( .A(p_input[1835]), .B(n29030), .Z(n54983) );
  XOR U54916 ( .A(p_input[1836]), .B(p_input[2060]), .Z(n54940) );
  XOR U54917 ( .A(n54950), .B(n54984), .Z(n54982) );
  IV U54918 ( .A(n54941), .Z(n54984) );
  XOR U54919 ( .A(p_input[1825]), .B(p_input[2049]), .Z(n54941) );
  XNOR U54920 ( .A(n54985), .B(n54957), .Z(n54950) );
  XNOR U54921 ( .A(p_input[1839]), .B(n29033), .Z(n54957) );
  XOR U54922 ( .A(n54947), .B(n54956), .Z(n54985) );
  XOR U54923 ( .A(n54986), .B(n54953), .Z(n54956) );
  XOR U54924 ( .A(p_input[1837]), .B(p_input[2061]), .Z(n54953) );
  XOR U54925 ( .A(p_input[1838]), .B(n29035), .Z(n54986) );
  XOR U54926 ( .A(p_input[1833]), .B(p_input[2057]), .Z(n54947) );
  XOR U54927 ( .A(n54965), .B(n54963), .Z(n54945) );
  XNOR U54928 ( .A(n54987), .B(n54970), .Z(n54963) );
  XOR U54929 ( .A(p_input[1832]), .B(p_input[2056]), .Z(n54970) );
  XOR U54930 ( .A(n54960), .B(n54969), .Z(n54987) );
  XOR U54931 ( .A(n54988), .B(n54966), .Z(n54969) );
  XOR U54932 ( .A(p_input[1830]), .B(p_input[2054]), .Z(n54966) );
  XOR U54933 ( .A(p_input[1831]), .B(n30404), .Z(n54988) );
  XOR U54934 ( .A(p_input[1826]), .B(p_input[2050]), .Z(n54960) );
  XNOR U54935 ( .A(n54975), .B(n54974), .Z(n54965) );
  XOR U54936 ( .A(n54989), .B(n54971), .Z(n54974) );
  XOR U54937 ( .A(p_input[1827]), .B(p_input[2051]), .Z(n54971) );
  XOR U54938 ( .A(p_input[1828]), .B(n30406), .Z(n54989) );
  XOR U54939 ( .A(p_input[1829]), .B(p_input[2053]), .Z(n54975) );
  XNOR U54940 ( .A(n54990), .B(n54991), .Z(n54871) );
  AND U54941 ( .A(n2241), .B(n54992), .Z(n54991) );
  XNOR U54942 ( .A(n54993), .B(n54994), .Z(n2241) );
  AND U54943 ( .A(n54995), .B(n54996), .Z(n54994) );
  XOR U54944 ( .A(n54885), .B(n54993), .Z(n54996) );
  XNOR U54945 ( .A(n54997), .B(n54993), .Z(n54995) );
  XOR U54946 ( .A(n54998), .B(n54999), .Z(n54993) );
  AND U54947 ( .A(n55000), .B(n55001), .Z(n54999) );
  XOR U54948 ( .A(n54900), .B(n54998), .Z(n55001) );
  XOR U54949 ( .A(n54998), .B(n54901), .Z(n55000) );
  XOR U54950 ( .A(n55002), .B(n55003), .Z(n54998) );
  AND U54951 ( .A(n55004), .B(n55005), .Z(n55003) );
  XOR U54952 ( .A(n54928), .B(n55002), .Z(n55005) );
  XOR U54953 ( .A(n55002), .B(n54929), .Z(n55004) );
  XOR U54954 ( .A(n55006), .B(n55007), .Z(n55002) );
  AND U54955 ( .A(n55008), .B(n55009), .Z(n55007) );
  XOR U54956 ( .A(n55006), .B(n54979), .Z(n55009) );
  XNOR U54957 ( .A(n55010), .B(n55011), .Z(n54831) );
  AND U54958 ( .A(n2245), .B(n55012), .Z(n55011) );
  XNOR U54959 ( .A(n55013), .B(n55014), .Z(n2245) );
  AND U54960 ( .A(n55015), .B(n55016), .Z(n55014) );
  XOR U54961 ( .A(n55013), .B(n54841), .Z(n55016) );
  XNOR U54962 ( .A(n55013), .B(n54801), .Z(n55015) );
  XOR U54963 ( .A(n55017), .B(n55018), .Z(n55013) );
  AND U54964 ( .A(n55019), .B(n55020), .Z(n55018) );
  XOR U54965 ( .A(n55017), .B(n54809), .Z(n55019) );
  XOR U54966 ( .A(n55021), .B(n55022), .Z(n54792) );
  AND U54967 ( .A(n2249), .B(n55012), .Z(n55022) );
  XNOR U54968 ( .A(n55010), .B(n55021), .Z(n55012) );
  XNOR U54969 ( .A(n55023), .B(n55024), .Z(n2249) );
  AND U54970 ( .A(n55025), .B(n55026), .Z(n55024) );
  XNOR U54971 ( .A(n55027), .B(n55023), .Z(n55026) );
  IV U54972 ( .A(n54841), .Z(n55027) );
  XOR U54973 ( .A(n54997), .B(n55028), .Z(n54841) );
  AND U54974 ( .A(n2252), .B(n55029), .Z(n55028) );
  XOR U54975 ( .A(n54884), .B(n54881), .Z(n55029) );
  IV U54976 ( .A(n54997), .Z(n54884) );
  XNOR U54977 ( .A(n54801), .B(n55023), .Z(n55025) );
  XOR U54978 ( .A(n55030), .B(n55031), .Z(n54801) );
  AND U54979 ( .A(n2268), .B(n55032), .Z(n55031) );
  XOR U54980 ( .A(n55017), .B(n55033), .Z(n55023) );
  AND U54981 ( .A(n55034), .B(n55020), .Z(n55033) );
  XNOR U54982 ( .A(n54851), .B(n55017), .Z(n55020) );
  XOR U54983 ( .A(n54901), .B(n55035), .Z(n54851) );
  AND U54984 ( .A(n2252), .B(n55036), .Z(n55035) );
  XOR U54985 ( .A(n54897), .B(n54901), .Z(n55036) );
  XNOR U54986 ( .A(n55037), .B(n55017), .Z(n55034) );
  IV U54987 ( .A(n54809), .Z(n55037) );
  XOR U54988 ( .A(n55038), .B(n55039), .Z(n54809) );
  AND U54989 ( .A(n2268), .B(n55040), .Z(n55039) );
  XOR U54990 ( .A(n55041), .B(n55042), .Z(n55017) );
  AND U54991 ( .A(n55043), .B(n55044), .Z(n55042) );
  XNOR U54992 ( .A(n54861), .B(n55041), .Z(n55044) );
  XOR U54993 ( .A(n54929), .B(n55045), .Z(n54861) );
  AND U54994 ( .A(n2252), .B(n55046), .Z(n55045) );
  XOR U54995 ( .A(n54925), .B(n54929), .Z(n55046) );
  XOR U54996 ( .A(n55041), .B(n54818), .Z(n55043) );
  XOR U54997 ( .A(n55047), .B(n55048), .Z(n54818) );
  AND U54998 ( .A(n2268), .B(n55049), .Z(n55048) );
  XOR U54999 ( .A(n55050), .B(n55051), .Z(n55041) );
  AND U55000 ( .A(n55052), .B(n55053), .Z(n55051) );
  XNOR U55001 ( .A(n55050), .B(n54869), .Z(n55053) );
  XOR U55002 ( .A(n54980), .B(n55054), .Z(n54869) );
  AND U55003 ( .A(n2252), .B(n55055), .Z(n55054) );
  XOR U55004 ( .A(n54976), .B(n54980), .Z(n55055) );
  XNOR U55005 ( .A(n55056), .B(n55050), .Z(n55052) );
  IV U55006 ( .A(n54828), .Z(n55056) );
  XOR U55007 ( .A(n55057), .B(n55058), .Z(n54828) );
  AND U55008 ( .A(n2268), .B(n55059), .Z(n55058) );
  AND U55009 ( .A(n55021), .B(n55010), .Z(n55050) );
  XNOR U55010 ( .A(n55060), .B(n55061), .Z(n55010) );
  AND U55011 ( .A(n2252), .B(n54992), .Z(n55061) );
  XNOR U55012 ( .A(n54990), .B(n55060), .Z(n54992) );
  XNOR U55013 ( .A(n55062), .B(n55063), .Z(n2252) );
  AND U55014 ( .A(n55064), .B(n55065), .Z(n55063) );
  XNOR U55015 ( .A(n55062), .B(n54881), .Z(n55065) );
  IV U55016 ( .A(n54885), .Z(n54881) );
  XOR U55017 ( .A(n55066), .B(n55067), .Z(n54885) );
  AND U55018 ( .A(n2256), .B(n55068), .Z(n55067) );
  XOR U55019 ( .A(n55069), .B(n55066), .Z(n55068) );
  XNOR U55020 ( .A(n55062), .B(n54997), .Z(n55064) );
  XOR U55021 ( .A(n55070), .B(n55071), .Z(n54997) );
  AND U55022 ( .A(n2264), .B(n55032), .Z(n55071) );
  XOR U55023 ( .A(n55030), .B(n55070), .Z(n55032) );
  XOR U55024 ( .A(n55072), .B(n55073), .Z(n55062) );
  AND U55025 ( .A(n55074), .B(n55075), .Z(n55073) );
  XNOR U55026 ( .A(n55072), .B(n54897), .Z(n55075) );
  IV U55027 ( .A(n54900), .Z(n54897) );
  XOR U55028 ( .A(n55076), .B(n55077), .Z(n54900) );
  AND U55029 ( .A(n2256), .B(n55078), .Z(n55077) );
  XOR U55030 ( .A(n55079), .B(n55076), .Z(n55078) );
  XOR U55031 ( .A(n54901), .B(n55072), .Z(n55074) );
  XOR U55032 ( .A(n55080), .B(n55081), .Z(n54901) );
  AND U55033 ( .A(n2264), .B(n55040), .Z(n55081) );
  XOR U55034 ( .A(n55080), .B(n55038), .Z(n55040) );
  XOR U55035 ( .A(n55082), .B(n55083), .Z(n55072) );
  AND U55036 ( .A(n55084), .B(n55085), .Z(n55083) );
  XNOR U55037 ( .A(n55082), .B(n54925), .Z(n55085) );
  IV U55038 ( .A(n54928), .Z(n54925) );
  XOR U55039 ( .A(n55086), .B(n55087), .Z(n54928) );
  AND U55040 ( .A(n2256), .B(n55088), .Z(n55087) );
  XNOR U55041 ( .A(n55089), .B(n55086), .Z(n55088) );
  XOR U55042 ( .A(n54929), .B(n55082), .Z(n55084) );
  XOR U55043 ( .A(n55090), .B(n55091), .Z(n54929) );
  AND U55044 ( .A(n2264), .B(n55049), .Z(n55091) );
  XOR U55045 ( .A(n55090), .B(n55047), .Z(n55049) );
  XOR U55046 ( .A(n55006), .B(n55092), .Z(n55082) );
  AND U55047 ( .A(n55008), .B(n55093), .Z(n55092) );
  XNOR U55048 ( .A(n55006), .B(n54976), .Z(n55093) );
  IV U55049 ( .A(n54979), .Z(n54976) );
  XOR U55050 ( .A(n55094), .B(n55095), .Z(n54979) );
  AND U55051 ( .A(n2256), .B(n55096), .Z(n55095) );
  XOR U55052 ( .A(n55097), .B(n55094), .Z(n55096) );
  XOR U55053 ( .A(n54980), .B(n55006), .Z(n55008) );
  XOR U55054 ( .A(n55098), .B(n55099), .Z(n54980) );
  AND U55055 ( .A(n2264), .B(n55059), .Z(n55099) );
  XOR U55056 ( .A(n55098), .B(n55057), .Z(n55059) );
  AND U55057 ( .A(n55060), .B(n54990), .Z(n55006) );
  XNOR U55058 ( .A(n55100), .B(n55101), .Z(n54990) );
  AND U55059 ( .A(n2256), .B(n55102), .Z(n55101) );
  XNOR U55060 ( .A(n55103), .B(n55100), .Z(n55102) );
  XNOR U55061 ( .A(n55104), .B(n55105), .Z(n2256) );
  AND U55062 ( .A(n55106), .B(n55107), .Z(n55105) );
  XOR U55063 ( .A(n55069), .B(n55104), .Z(n55107) );
  AND U55064 ( .A(n55108), .B(n55109), .Z(n55069) );
  XNOR U55065 ( .A(n55066), .B(n55104), .Z(n55106) );
  XNOR U55066 ( .A(n55110), .B(n55111), .Z(n55066) );
  AND U55067 ( .A(n2260), .B(n55112), .Z(n55111) );
  XNOR U55068 ( .A(n55113), .B(n55114), .Z(n55112) );
  XOR U55069 ( .A(n55115), .B(n55116), .Z(n55104) );
  AND U55070 ( .A(n55117), .B(n55118), .Z(n55116) );
  XNOR U55071 ( .A(n55115), .B(n55108), .Z(n55118) );
  IV U55072 ( .A(n55079), .Z(n55108) );
  XOR U55073 ( .A(n55119), .B(n55120), .Z(n55079) );
  XOR U55074 ( .A(n55121), .B(n55109), .Z(n55120) );
  AND U55075 ( .A(n55089), .B(n55122), .Z(n55109) );
  AND U55076 ( .A(n55123), .B(n55124), .Z(n55121) );
  XOR U55077 ( .A(n55125), .B(n55119), .Z(n55123) );
  XNOR U55078 ( .A(n55076), .B(n55115), .Z(n55117) );
  XNOR U55079 ( .A(n55126), .B(n55127), .Z(n55076) );
  AND U55080 ( .A(n2260), .B(n55128), .Z(n55127) );
  XNOR U55081 ( .A(n55129), .B(n55130), .Z(n55128) );
  XOR U55082 ( .A(n55131), .B(n55132), .Z(n55115) );
  AND U55083 ( .A(n55133), .B(n55134), .Z(n55132) );
  XNOR U55084 ( .A(n55131), .B(n55089), .Z(n55134) );
  XOR U55085 ( .A(n55135), .B(n55124), .Z(n55089) );
  XNOR U55086 ( .A(n55136), .B(n55119), .Z(n55124) );
  XOR U55087 ( .A(n55137), .B(n55138), .Z(n55119) );
  AND U55088 ( .A(n55139), .B(n55140), .Z(n55138) );
  XOR U55089 ( .A(n55141), .B(n55137), .Z(n55139) );
  XNOR U55090 ( .A(n55142), .B(n55143), .Z(n55136) );
  AND U55091 ( .A(n55144), .B(n55145), .Z(n55143) );
  XOR U55092 ( .A(n55142), .B(n55146), .Z(n55144) );
  XNOR U55093 ( .A(n55125), .B(n55122), .Z(n55135) );
  AND U55094 ( .A(n55147), .B(n55148), .Z(n55122) );
  XOR U55095 ( .A(n55149), .B(n55150), .Z(n55125) );
  AND U55096 ( .A(n55151), .B(n55152), .Z(n55150) );
  XOR U55097 ( .A(n55149), .B(n55153), .Z(n55151) );
  XNOR U55098 ( .A(n55086), .B(n55131), .Z(n55133) );
  XNOR U55099 ( .A(n55154), .B(n55155), .Z(n55086) );
  AND U55100 ( .A(n2260), .B(n55156), .Z(n55155) );
  XNOR U55101 ( .A(n55157), .B(n55158), .Z(n55156) );
  XOR U55102 ( .A(n55159), .B(n55160), .Z(n55131) );
  AND U55103 ( .A(n55161), .B(n55162), .Z(n55160) );
  XNOR U55104 ( .A(n55159), .B(n55147), .Z(n55162) );
  IV U55105 ( .A(n55097), .Z(n55147) );
  XNOR U55106 ( .A(n55163), .B(n55140), .Z(n55097) );
  XNOR U55107 ( .A(n55164), .B(n55146), .Z(n55140) );
  XNOR U55108 ( .A(n55165), .B(n55166), .Z(n55146) );
  NOR U55109 ( .A(n55167), .B(n55168), .Z(n55166) );
  XOR U55110 ( .A(n55165), .B(n55169), .Z(n55167) );
  XNOR U55111 ( .A(n55145), .B(n55137), .Z(n55164) );
  XOR U55112 ( .A(n55170), .B(n55171), .Z(n55137) );
  AND U55113 ( .A(n55172), .B(n55173), .Z(n55171) );
  XOR U55114 ( .A(n55170), .B(n55174), .Z(n55172) );
  XNOR U55115 ( .A(n55175), .B(n55142), .Z(n55145) );
  XOR U55116 ( .A(n55176), .B(n55177), .Z(n55142) );
  AND U55117 ( .A(n55178), .B(n55179), .Z(n55177) );
  XNOR U55118 ( .A(n55180), .B(n55181), .Z(n55178) );
  IV U55119 ( .A(n55176), .Z(n55180) );
  XNOR U55120 ( .A(n55182), .B(n55183), .Z(n55175) );
  NOR U55121 ( .A(n55184), .B(n55185), .Z(n55183) );
  XNOR U55122 ( .A(n55182), .B(n55186), .Z(n55184) );
  XNOR U55123 ( .A(n55141), .B(n55148), .Z(n55163) );
  NOR U55124 ( .A(n55103), .B(n55187), .Z(n55148) );
  XOR U55125 ( .A(n55153), .B(n55152), .Z(n55141) );
  XNOR U55126 ( .A(n55188), .B(n55149), .Z(n55152) );
  XOR U55127 ( .A(n55189), .B(n55190), .Z(n55149) );
  AND U55128 ( .A(n55191), .B(n55192), .Z(n55190) );
  XNOR U55129 ( .A(n55193), .B(n55194), .Z(n55191) );
  IV U55130 ( .A(n55189), .Z(n55193) );
  XNOR U55131 ( .A(n55195), .B(n55196), .Z(n55188) );
  NOR U55132 ( .A(n55197), .B(n55198), .Z(n55196) );
  XNOR U55133 ( .A(n55195), .B(n55199), .Z(n55197) );
  XOR U55134 ( .A(n55200), .B(n55201), .Z(n55153) );
  NOR U55135 ( .A(n55202), .B(n55203), .Z(n55201) );
  XNOR U55136 ( .A(n55200), .B(n55204), .Z(n55202) );
  XNOR U55137 ( .A(n55094), .B(n55159), .Z(n55161) );
  XNOR U55138 ( .A(n55205), .B(n55206), .Z(n55094) );
  AND U55139 ( .A(n2260), .B(n55207), .Z(n55206) );
  XNOR U55140 ( .A(n55208), .B(n55209), .Z(n55207) );
  AND U55141 ( .A(n55100), .B(n55103), .Z(n55159) );
  XOR U55142 ( .A(n55210), .B(n55187), .Z(n55103) );
  XNOR U55143 ( .A(p_input[1840]), .B(p_input[2048]), .Z(n55187) );
  XNOR U55144 ( .A(n55174), .B(n55173), .Z(n55210) );
  XNOR U55145 ( .A(n55211), .B(n55181), .Z(n55173) );
  XNOR U55146 ( .A(n55169), .B(n55168), .Z(n55181) );
  XNOR U55147 ( .A(n55212), .B(n55165), .Z(n55168) );
  XNOR U55148 ( .A(p_input[1850]), .B(p_input[2058]), .Z(n55165) );
  XOR U55149 ( .A(p_input[1851]), .B(n29030), .Z(n55212) );
  XOR U55150 ( .A(p_input[1852]), .B(p_input[2060]), .Z(n55169) );
  XOR U55151 ( .A(n55179), .B(n55213), .Z(n55211) );
  IV U55152 ( .A(n55170), .Z(n55213) );
  XOR U55153 ( .A(p_input[1841]), .B(p_input[2049]), .Z(n55170) );
  XNOR U55154 ( .A(n55214), .B(n55186), .Z(n55179) );
  XNOR U55155 ( .A(p_input[1855]), .B(n29033), .Z(n55186) );
  XOR U55156 ( .A(n55176), .B(n55185), .Z(n55214) );
  XOR U55157 ( .A(n55215), .B(n55182), .Z(n55185) );
  XOR U55158 ( .A(p_input[1853]), .B(p_input[2061]), .Z(n55182) );
  XOR U55159 ( .A(p_input[1854]), .B(n29035), .Z(n55215) );
  XOR U55160 ( .A(p_input[1849]), .B(p_input[2057]), .Z(n55176) );
  XOR U55161 ( .A(n55194), .B(n55192), .Z(n55174) );
  XNOR U55162 ( .A(n55216), .B(n55199), .Z(n55192) );
  XOR U55163 ( .A(p_input[1848]), .B(p_input[2056]), .Z(n55199) );
  XOR U55164 ( .A(n55189), .B(n55198), .Z(n55216) );
  XOR U55165 ( .A(n55217), .B(n55195), .Z(n55198) );
  XOR U55166 ( .A(p_input[1846]), .B(p_input[2054]), .Z(n55195) );
  XOR U55167 ( .A(p_input[1847]), .B(n30404), .Z(n55217) );
  XOR U55168 ( .A(p_input[1842]), .B(p_input[2050]), .Z(n55189) );
  XNOR U55169 ( .A(n55204), .B(n55203), .Z(n55194) );
  XOR U55170 ( .A(n55218), .B(n55200), .Z(n55203) );
  XOR U55171 ( .A(p_input[1843]), .B(p_input[2051]), .Z(n55200) );
  XOR U55172 ( .A(p_input[1844]), .B(n30406), .Z(n55218) );
  XOR U55173 ( .A(p_input[1845]), .B(p_input[2053]), .Z(n55204) );
  XNOR U55174 ( .A(n55219), .B(n55220), .Z(n55100) );
  AND U55175 ( .A(n2260), .B(n55221), .Z(n55220) );
  XNOR U55176 ( .A(n55222), .B(n55223), .Z(n2260) );
  AND U55177 ( .A(n55224), .B(n55225), .Z(n55223) );
  XOR U55178 ( .A(n55114), .B(n55222), .Z(n55225) );
  XNOR U55179 ( .A(n55226), .B(n55222), .Z(n55224) );
  XOR U55180 ( .A(n55227), .B(n55228), .Z(n55222) );
  AND U55181 ( .A(n55229), .B(n55230), .Z(n55228) );
  XOR U55182 ( .A(n55129), .B(n55227), .Z(n55230) );
  XOR U55183 ( .A(n55227), .B(n55130), .Z(n55229) );
  XOR U55184 ( .A(n55231), .B(n55232), .Z(n55227) );
  AND U55185 ( .A(n55233), .B(n55234), .Z(n55232) );
  XOR U55186 ( .A(n55157), .B(n55231), .Z(n55234) );
  XOR U55187 ( .A(n55231), .B(n55158), .Z(n55233) );
  XOR U55188 ( .A(n55235), .B(n55236), .Z(n55231) );
  AND U55189 ( .A(n55237), .B(n55238), .Z(n55236) );
  XOR U55190 ( .A(n55235), .B(n55208), .Z(n55238) );
  XNOR U55191 ( .A(n55239), .B(n55240), .Z(n55060) );
  AND U55192 ( .A(n2264), .B(n55241), .Z(n55240) );
  XNOR U55193 ( .A(n55242), .B(n55243), .Z(n2264) );
  AND U55194 ( .A(n55244), .B(n55245), .Z(n55243) );
  XOR U55195 ( .A(n55242), .B(n55070), .Z(n55245) );
  XNOR U55196 ( .A(n55242), .B(n55030), .Z(n55244) );
  XOR U55197 ( .A(n55246), .B(n55247), .Z(n55242) );
  AND U55198 ( .A(n55248), .B(n55249), .Z(n55247) );
  XOR U55199 ( .A(n55246), .B(n55038), .Z(n55248) );
  XOR U55200 ( .A(n55250), .B(n55251), .Z(n55021) );
  AND U55201 ( .A(n2268), .B(n55241), .Z(n55251) );
  XNOR U55202 ( .A(n55239), .B(n55250), .Z(n55241) );
  XNOR U55203 ( .A(n55252), .B(n55253), .Z(n2268) );
  AND U55204 ( .A(n55254), .B(n55255), .Z(n55253) );
  XNOR U55205 ( .A(n55256), .B(n55252), .Z(n55255) );
  IV U55206 ( .A(n55070), .Z(n55256) );
  XOR U55207 ( .A(n55226), .B(n55257), .Z(n55070) );
  AND U55208 ( .A(n2271), .B(n55258), .Z(n55257) );
  XOR U55209 ( .A(n55113), .B(n55110), .Z(n55258) );
  IV U55210 ( .A(n55226), .Z(n55113) );
  XNOR U55211 ( .A(n55030), .B(n55252), .Z(n55254) );
  XOR U55212 ( .A(n55259), .B(n55260), .Z(n55030) );
  AND U55213 ( .A(n2287), .B(n55261), .Z(n55260) );
  XOR U55214 ( .A(n55246), .B(n55262), .Z(n55252) );
  AND U55215 ( .A(n55263), .B(n55249), .Z(n55262) );
  XNOR U55216 ( .A(n55080), .B(n55246), .Z(n55249) );
  XOR U55217 ( .A(n55130), .B(n55264), .Z(n55080) );
  AND U55218 ( .A(n2271), .B(n55265), .Z(n55264) );
  XOR U55219 ( .A(n55126), .B(n55130), .Z(n55265) );
  XNOR U55220 ( .A(n55266), .B(n55246), .Z(n55263) );
  IV U55221 ( .A(n55038), .Z(n55266) );
  XOR U55222 ( .A(n55267), .B(n55268), .Z(n55038) );
  AND U55223 ( .A(n2287), .B(n55269), .Z(n55268) );
  XOR U55224 ( .A(n55270), .B(n55271), .Z(n55246) );
  AND U55225 ( .A(n55272), .B(n55273), .Z(n55271) );
  XNOR U55226 ( .A(n55090), .B(n55270), .Z(n55273) );
  XOR U55227 ( .A(n55158), .B(n55274), .Z(n55090) );
  AND U55228 ( .A(n2271), .B(n55275), .Z(n55274) );
  XOR U55229 ( .A(n55154), .B(n55158), .Z(n55275) );
  XOR U55230 ( .A(n55270), .B(n55047), .Z(n55272) );
  XOR U55231 ( .A(n55276), .B(n55277), .Z(n55047) );
  AND U55232 ( .A(n2287), .B(n55278), .Z(n55277) );
  XOR U55233 ( .A(n55279), .B(n55280), .Z(n55270) );
  AND U55234 ( .A(n55281), .B(n55282), .Z(n55280) );
  XNOR U55235 ( .A(n55279), .B(n55098), .Z(n55282) );
  XOR U55236 ( .A(n55209), .B(n55283), .Z(n55098) );
  AND U55237 ( .A(n2271), .B(n55284), .Z(n55283) );
  XOR U55238 ( .A(n55205), .B(n55209), .Z(n55284) );
  XNOR U55239 ( .A(n55285), .B(n55279), .Z(n55281) );
  IV U55240 ( .A(n55057), .Z(n55285) );
  XOR U55241 ( .A(n55286), .B(n55287), .Z(n55057) );
  AND U55242 ( .A(n2287), .B(n55288), .Z(n55287) );
  AND U55243 ( .A(n55250), .B(n55239), .Z(n55279) );
  XNOR U55244 ( .A(n55289), .B(n55290), .Z(n55239) );
  AND U55245 ( .A(n2271), .B(n55221), .Z(n55290) );
  XNOR U55246 ( .A(n55219), .B(n55289), .Z(n55221) );
  XNOR U55247 ( .A(n55291), .B(n55292), .Z(n2271) );
  AND U55248 ( .A(n55293), .B(n55294), .Z(n55292) );
  XNOR U55249 ( .A(n55291), .B(n55110), .Z(n55294) );
  IV U55250 ( .A(n55114), .Z(n55110) );
  XOR U55251 ( .A(n55295), .B(n55296), .Z(n55114) );
  AND U55252 ( .A(n2275), .B(n55297), .Z(n55296) );
  XOR U55253 ( .A(n55298), .B(n55295), .Z(n55297) );
  XNOR U55254 ( .A(n55291), .B(n55226), .Z(n55293) );
  XOR U55255 ( .A(n55299), .B(n55300), .Z(n55226) );
  AND U55256 ( .A(n2283), .B(n55261), .Z(n55300) );
  XOR U55257 ( .A(n55259), .B(n55299), .Z(n55261) );
  XOR U55258 ( .A(n55301), .B(n55302), .Z(n55291) );
  AND U55259 ( .A(n55303), .B(n55304), .Z(n55302) );
  XNOR U55260 ( .A(n55301), .B(n55126), .Z(n55304) );
  IV U55261 ( .A(n55129), .Z(n55126) );
  XOR U55262 ( .A(n55305), .B(n55306), .Z(n55129) );
  AND U55263 ( .A(n2275), .B(n55307), .Z(n55306) );
  XOR U55264 ( .A(n55308), .B(n55305), .Z(n55307) );
  XOR U55265 ( .A(n55130), .B(n55301), .Z(n55303) );
  XOR U55266 ( .A(n55309), .B(n55310), .Z(n55130) );
  AND U55267 ( .A(n2283), .B(n55269), .Z(n55310) );
  XOR U55268 ( .A(n55309), .B(n55267), .Z(n55269) );
  XOR U55269 ( .A(n55311), .B(n55312), .Z(n55301) );
  AND U55270 ( .A(n55313), .B(n55314), .Z(n55312) );
  XNOR U55271 ( .A(n55311), .B(n55154), .Z(n55314) );
  IV U55272 ( .A(n55157), .Z(n55154) );
  XOR U55273 ( .A(n55315), .B(n55316), .Z(n55157) );
  AND U55274 ( .A(n2275), .B(n55317), .Z(n55316) );
  XNOR U55275 ( .A(n55318), .B(n55315), .Z(n55317) );
  XOR U55276 ( .A(n55158), .B(n55311), .Z(n55313) );
  XOR U55277 ( .A(n55319), .B(n55320), .Z(n55158) );
  AND U55278 ( .A(n2283), .B(n55278), .Z(n55320) );
  XOR U55279 ( .A(n55319), .B(n55276), .Z(n55278) );
  XOR U55280 ( .A(n55235), .B(n55321), .Z(n55311) );
  AND U55281 ( .A(n55237), .B(n55322), .Z(n55321) );
  XNOR U55282 ( .A(n55235), .B(n55205), .Z(n55322) );
  IV U55283 ( .A(n55208), .Z(n55205) );
  XOR U55284 ( .A(n55323), .B(n55324), .Z(n55208) );
  AND U55285 ( .A(n2275), .B(n55325), .Z(n55324) );
  XOR U55286 ( .A(n55326), .B(n55323), .Z(n55325) );
  XOR U55287 ( .A(n55209), .B(n55235), .Z(n55237) );
  XOR U55288 ( .A(n55327), .B(n55328), .Z(n55209) );
  AND U55289 ( .A(n2283), .B(n55288), .Z(n55328) );
  XOR U55290 ( .A(n55327), .B(n55286), .Z(n55288) );
  AND U55291 ( .A(n55289), .B(n55219), .Z(n55235) );
  XNOR U55292 ( .A(n55329), .B(n55330), .Z(n55219) );
  AND U55293 ( .A(n2275), .B(n55331), .Z(n55330) );
  XNOR U55294 ( .A(n55332), .B(n55329), .Z(n55331) );
  XNOR U55295 ( .A(n55333), .B(n55334), .Z(n2275) );
  AND U55296 ( .A(n55335), .B(n55336), .Z(n55334) );
  XOR U55297 ( .A(n55298), .B(n55333), .Z(n55336) );
  AND U55298 ( .A(n55337), .B(n55338), .Z(n55298) );
  XNOR U55299 ( .A(n55295), .B(n55333), .Z(n55335) );
  XNOR U55300 ( .A(n55339), .B(n55340), .Z(n55295) );
  AND U55301 ( .A(n2279), .B(n55341), .Z(n55340) );
  XNOR U55302 ( .A(n55342), .B(n55343), .Z(n55341) );
  XOR U55303 ( .A(n55344), .B(n55345), .Z(n55333) );
  AND U55304 ( .A(n55346), .B(n55347), .Z(n55345) );
  XNOR U55305 ( .A(n55344), .B(n55337), .Z(n55347) );
  IV U55306 ( .A(n55308), .Z(n55337) );
  XOR U55307 ( .A(n55348), .B(n55349), .Z(n55308) );
  XOR U55308 ( .A(n55350), .B(n55338), .Z(n55349) );
  AND U55309 ( .A(n55318), .B(n55351), .Z(n55338) );
  AND U55310 ( .A(n55352), .B(n55353), .Z(n55350) );
  XOR U55311 ( .A(n55354), .B(n55348), .Z(n55352) );
  XNOR U55312 ( .A(n55305), .B(n55344), .Z(n55346) );
  XNOR U55313 ( .A(n55355), .B(n55356), .Z(n55305) );
  AND U55314 ( .A(n2279), .B(n55357), .Z(n55356) );
  XNOR U55315 ( .A(n55358), .B(n55359), .Z(n55357) );
  XOR U55316 ( .A(n55360), .B(n55361), .Z(n55344) );
  AND U55317 ( .A(n55362), .B(n55363), .Z(n55361) );
  XNOR U55318 ( .A(n55360), .B(n55318), .Z(n55363) );
  XOR U55319 ( .A(n55364), .B(n55353), .Z(n55318) );
  XNOR U55320 ( .A(n55365), .B(n55348), .Z(n55353) );
  XOR U55321 ( .A(n55366), .B(n55367), .Z(n55348) );
  AND U55322 ( .A(n55368), .B(n55369), .Z(n55367) );
  XOR U55323 ( .A(n55370), .B(n55366), .Z(n55368) );
  XNOR U55324 ( .A(n55371), .B(n55372), .Z(n55365) );
  AND U55325 ( .A(n55373), .B(n55374), .Z(n55372) );
  XOR U55326 ( .A(n55371), .B(n55375), .Z(n55373) );
  XNOR U55327 ( .A(n55354), .B(n55351), .Z(n55364) );
  AND U55328 ( .A(n55376), .B(n55377), .Z(n55351) );
  XOR U55329 ( .A(n55378), .B(n55379), .Z(n55354) );
  AND U55330 ( .A(n55380), .B(n55381), .Z(n55379) );
  XOR U55331 ( .A(n55378), .B(n55382), .Z(n55380) );
  XNOR U55332 ( .A(n55315), .B(n55360), .Z(n55362) );
  XNOR U55333 ( .A(n55383), .B(n55384), .Z(n55315) );
  AND U55334 ( .A(n2279), .B(n55385), .Z(n55384) );
  XNOR U55335 ( .A(n55386), .B(n55387), .Z(n55385) );
  XOR U55336 ( .A(n55388), .B(n55389), .Z(n55360) );
  AND U55337 ( .A(n55390), .B(n55391), .Z(n55389) );
  XNOR U55338 ( .A(n55388), .B(n55376), .Z(n55391) );
  IV U55339 ( .A(n55326), .Z(n55376) );
  XNOR U55340 ( .A(n55392), .B(n55369), .Z(n55326) );
  XNOR U55341 ( .A(n55393), .B(n55375), .Z(n55369) );
  XNOR U55342 ( .A(n55394), .B(n55395), .Z(n55375) );
  NOR U55343 ( .A(n55396), .B(n55397), .Z(n55395) );
  XOR U55344 ( .A(n55394), .B(n55398), .Z(n55396) );
  XNOR U55345 ( .A(n55374), .B(n55366), .Z(n55393) );
  XOR U55346 ( .A(n55399), .B(n55400), .Z(n55366) );
  AND U55347 ( .A(n55401), .B(n55402), .Z(n55400) );
  XOR U55348 ( .A(n55399), .B(n55403), .Z(n55401) );
  XNOR U55349 ( .A(n55404), .B(n55371), .Z(n55374) );
  XOR U55350 ( .A(n55405), .B(n55406), .Z(n55371) );
  AND U55351 ( .A(n55407), .B(n55408), .Z(n55406) );
  XNOR U55352 ( .A(n55409), .B(n55410), .Z(n55407) );
  IV U55353 ( .A(n55405), .Z(n55409) );
  XNOR U55354 ( .A(n55411), .B(n55412), .Z(n55404) );
  NOR U55355 ( .A(n55413), .B(n55414), .Z(n55412) );
  XNOR U55356 ( .A(n55411), .B(n55415), .Z(n55413) );
  XNOR U55357 ( .A(n55370), .B(n55377), .Z(n55392) );
  NOR U55358 ( .A(n55332), .B(n55416), .Z(n55377) );
  XOR U55359 ( .A(n55382), .B(n55381), .Z(n55370) );
  XNOR U55360 ( .A(n55417), .B(n55378), .Z(n55381) );
  XOR U55361 ( .A(n55418), .B(n55419), .Z(n55378) );
  AND U55362 ( .A(n55420), .B(n55421), .Z(n55419) );
  XNOR U55363 ( .A(n55422), .B(n55423), .Z(n55420) );
  IV U55364 ( .A(n55418), .Z(n55422) );
  XNOR U55365 ( .A(n55424), .B(n55425), .Z(n55417) );
  NOR U55366 ( .A(n55426), .B(n55427), .Z(n55425) );
  XNOR U55367 ( .A(n55424), .B(n55428), .Z(n55426) );
  XOR U55368 ( .A(n55429), .B(n55430), .Z(n55382) );
  NOR U55369 ( .A(n55431), .B(n55432), .Z(n55430) );
  XNOR U55370 ( .A(n55429), .B(n55433), .Z(n55431) );
  XNOR U55371 ( .A(n55323), .B(n55388), .Z(n55390) );
  XNOR U55372 ( .A(n55434), .B(n55435), .Z(n55323) );
  AND U55373 ( .A(n2279), .B(n55436), .Z(n55435) );
  XNOR U55374 ( .A(n55437), .B(n55438), .Z(n55436) );
  AND U55375 ( .A(n55329), .B(n55332), .Z(n55388) );
  XOR U55376 ( .A(n55439), .B(n55416), .Z(n55332) );
  XNOR U55377 ( .A(p_input[1856]), .B(p_input[2048]), .Z(n55416) );
  XNOR U55378 ( .A(n55403), .B(n55402), .Z(n55439) );
  XNOR U55379 ( .A(n55440), .B(n55410), .Z(n55402) );
  XNOR U55380 ( .A(n55398), .B(n55397), .Z(n55410) );
  XNOR U55381 ( .A(n55441), .B(n55394), .Z(n55397) );
  XNOR U55382 ( .A(p_input[1866]), .B(p_input[2058]), .Z(n55394) );
  XOR U55383 ( .A(p_input[1867]), .B(n29030), .Z(n55441) );
  XOR U55384 ( .A(p_input[1868]), .B(p_input[2060]), .Z(n55398) );
  XOR U55385 ( .A(n55408), .B(n55442), .Z(n55440) );
  IV U55386 ( .A(n55399), .Z(n55442) );
  XOR U55387 ( .A(p_input[1857]), .B(p_input[2049]), .Z(n55399) );
  XNOR U55388 ( .A(n55443), .B(n55415), .Z(n55408) );
  XNOR U55389 ( .A(p_input[1871]), .B(n29033), .Z(n55415) );
  XOR U55390 ( .A(n55405), .B(n55414), .Z(n55443) );
  XOR U55391 ( .A(n55444), .B(n55411), .Z(n55414) );
  XOR U55392 ( .A(p_input[1869]), .B(p_input[2061]), .Z(n55411) );
  XOR U55393 ( .A(p_input[1870]), .B(n29035), .Z(n55444) );
  XOR U55394 ( .A(p_input[1865]), .B(p_input[2057]), .Z(n55405) );
  XOR U55395 ( .A(n55423), .B(n55421), .Z(n55403) );
  XNOR U55396 ( .A(n55445), .B(n55428), .Z(n55421) );
  XOR U55397 ( .A(p_input[1864]), .B(p_input[2056]), .Z(n55428) );
  XOR U55398 ( .A(n55418), .B(n55427), .Z(n55445) );
  XOR U55399 ( .A(n55446), .B(n55424), .Z(n55427) );
  XOR U55400 ( .A(p_input[1862]), .B(p_input[2054]), .Z(n55424) );
  XOR U55401 ( .A(p_input[1863]), .B(n30404), .Z(n55446) );
  XOR U55402 ( .A(p_input[1858]), .B(p_input[2050]), .Z(n55418) );
  XNOR U55403 ( .A(n55433), .B(n55432), .Z(n55423) );
  XOR U55404 ( .A(n55447), .B(n55429), .Z(n55432) );
  XOR U55405 ( .A(p_input[1859]), .B(p_input[2051]), .Z(n55429) );
  XOR U55406 ( .A(p_input[1860]), .B(n30406), .Z(n55447) );
  XOR U55407 ( .A(p_input[1861]), .B(p_input[2053]), .Z(n55433) );
  XNOR U55408 ( .A(n55448), .B(n55449), .Z(n55329) );
  AND U55409 ( .A(n2279), .B(n55450), .Z(n55449) );
  XNOR U55410 ( .A(n55451), .B(n55452), .Z(n2279) );
  AND U55411 ( .A(n55453), .B(n55454), .Z(n55452) );
  XOR U55412 ( .A(n55343), .B(n55451), .Z(n55454) );
  XNOR U55413 ( .A(n55455), .B(n55451), .Z(n55453) );
  XOR U55414 ( .A(n55456), .B(n55457), .Z(n55451) );
  AND U55415 ( .A(n55458), .B(n55459), .Z(n55457) );
  XOR U55416 ( .A(n55358), .B(n55456), .Z(n55459) );
  XOR U55417 ( .A(n55456), .B(n55359), .Z(n55458) );
  XOR U55418 ( .A(n55460), .B(n55461), .Z(n55456) );
  AND U55419 ( .A(n55462), .B(n55463), .Z(n55461) );
  XOR U55420 ( .A(n55386), .B(n55460), .Z(n55463) );
  XOR U55421 ( .A(n55460), .B(n55387), .Z(n55462) );
  XOR U55422 ( .A(n55464), .B(n55465), .Z(n55460) );
  AND U55423 ( .A(n55466), .B(n55467), .Z(n55465) );
  XOR U55424 ( .A(n55464), .B(n55437), .Z(n55467) );
  XNOR U55425 ( .A(n55468), .B(n55469), .Z(n55289) );
  AND U55426 ( .A(n2283), .B(n55470), .Z(n55469) );
  XNOR U55427 ( .A(n55471), .B(n55472), .Z(n2283) );
  AND U55428 ( .A(n55473), .B(n55474), .Z(n55472) );
  XOR U55429 ( .A(n55471), .B(n55299), .Z(n55474) );
  XNOR U55430 ( .A(n55471), .B(n55259), .Z(n55473) );
  XOR U55431 ( .A(n55475), .B(n55476), .Z(n55471) );
  AND U55432 ( .A(n55477), .B(n55478), .Z(n55476) );
  XOR U55433 ( .A(n55475), .B(n55267), .Z(n55477) );
  XOR U55434 ( .A(n55479), .B(n55480), .Z(n55250) );
  AND U55435 ( .A(n2287), .B(n55470), .Z(n55480) );
  XNOR U55436 ( .A(n55468), .B(n55479), .Z(n55470) );
  XNOR U55437 ( .A(n55481), .B(n55482), .Z(n2287) );
  AND U55438 ( .A(n55483), .B(n55484), .Z(n55482) );
  XNOR U55439 ( .A(n55485), .B(n55481), .Z(n55484) );
  IV U55440 ( .A(n55299), .Z(n55485) );
  XOR U55441 ( .A(n55455), .B(n55486), .Z(n55299) );
  AND U55442 ( .A(n2290), .B(n55487), .Z(n55486) );
  XOR U55443 ( .A(n55342), .B(n55339), .Z(n55487) );
  IV U55444 ( .A(n55455), .Z(n55342) );
  XNOR U55445 ( .A(n55259), .B(n55481), .Z(n55483) );
  XOR U55446 ( .A(n55488), .B(n55489), .Z(n55259) );
  AND U55447 ( .A(n2306), .B(n55490), .Z(n55489) );
  XOR U55448 ( .A(n55475), .B(n55491), .Z(n55481) );
  AND U55449 ( .A(n55492), .B(n55478), .Z(n55491) );
  XNOR U55450 ( .A(n55309), .B(n55475), .Z(n55478) );
  XOR U55451 ( .A(n55359), .B(n55493), .Z(n55309) );
  AND U55452 ( .A(n2290), .B(n55494), .Z(n55493) );
  XOR U55453 ( .A(n55355), .B(n55359), .Z(n55494) );
  XNOR U55454 ( .A(n55495), .B(n55475), .Z(n55492) );
  IV U55455 ( .A(n55267), .Z(n55495) );
  XOR U55456 ( .A(n55496), .B(n55497), .Z(n55267) );
  AND U55457 ( .A(n2306), .B(n55498), .Z(n55497) );
  XOR U55458 ( .A(n55499), .B(n55500), .Z(n55475) );
  AND U55459 ( .A(n55501), .B(n55502), .Z(n55500) );
  XNOR U55460 ( .A(n55319), .B(n55499), .Z(n55502) );
  XOR U55461 ( .A(n55387), .B(n55503), .Z(n55319) );
  AND U55462 ( .A(n2290), .B(n55504), .Z(n55503) );
  XOR U55463 ( .A(n55383), .B(n55387), .Z(n55504) );
  XOR U55464 ( .A(n55499), .B(n55276), .Z(n55501) );
  XOR U55465 ( .A(n55505), .B(n55506), .Z(n55276) );
  AND U55466 ( .A(n2306), .B(n55507), .Z(n55506) );
  XOR U55467 ( .A(n55508), .B(n55509), .Z(n55499) );
  AND U55468 ( .A(n55510), .B(n55511), .Z(n55509) );
  XNOR U55469 ( .A(n55508), .B(n55327), .Z(n55511) );
  XOR U55470 ( .A(n55438), .B(n55512), .Z(n55327) );
  AND U55471 ( .A(n2290), .B(n55513), .Z(n55512) );
  XOR U55472 ( .A(n55434), .B(n55438), .Z(n55513) );
  XNOR U55473 ( .A(n55514), .B(n55508), .Z(n55510) );
  IV U55474 ( .A(n55286), .Z(n55514) );
  XOR U55475 ( .A(n55515), .B(n55516), .Z(n55286) );
  AND U55476 ( .A(n2306), .B(n55517), .Z(n55516) );
  AND U55477 ( .A(n55479), .B(n55468), .Z(n55508) );
  XNOR U55478 ( .A(n55518), .B(n55519), .Z(n55468) );
  AND U55479 ( .A(n2290), .B(n55450), .Z(n55519) );
  XNOR U55480 ( .A(n55448), .B(n55518), .Z(n55450) );
  XNOR U55481 ( .A(n55520), .B(n55521), .Z(n2290) );
  AND U55482 ( .A(n55522), .B(n55523), .Z(n55521) );
  XNOR U55483 ( .A(n55520), .B(n55339), .Z(n55523) );
  IV U55484 ( .A(n55343), .Z(n55339) );
  XOR U55485 ( .A(n55524), .B(n55525), .Z(n55343) );
  AND U55486 ( .A(n2294), .B(n55526), .Z(n55525) );
  XOR U55487 ( .A(n55527), .B(n55524), .Z(n55526) );
  XNOR U55488 ( .A(n55520), .B(n55455), .Z(n55522) );
  XOR U55489 ( .A(n55528), .B(n55529), .Z(n55455) );
  AND U55490 ( .A(n2302), .B(n55490), .Z(n55529) );
  XOR U55491 ( .A(n55488), .B(n55528), .Z(n55490) );
  XOR U55492 ( .A(n55530), .B(n55531), .Z(n55520) );
  AND U55493 ( .A(n55532), .B(n55533), .Z(n55531) );
  XNOR U55494 ( .A(n55530), .B(n55355), .Z(n55533) );
  IV U55495 ( .A(n55358), .Z(n55355) );
  XOR U55496 ( .A(n55534), .B(n55535), .Z(n55358) );
  AND U55497 ( .A(n2294), .B(n55536), .Z(n55535) );
  XOR U55498 ( .A(n55537), .B(n55534), .Z(n55536) );
  XOR U55499 ( .A(n55359), .B(n55530), .Z(n55532) );
  XOR U55500 ( .A(n55538), .B(n55539), .Z(n55359) );
  AND U55501 ( .A(n2302), .B(n55498), .Z(n55539) );
  XOR U55502 ( .A(n55538), .B(n55496), .Z(n55498) );
  XOR U55503 ( .A(n55540), .B(n55541), .Z(n55530) );
  AND U55504 ( .A(n55542), .B(n55543), .Z(n55541) );
  XNOR U55505 ( .A(n55540), .B(n55383), .Z(n55543) );
  IV U55506 ( .A(n55386), .Z(n55383) );
  XOR U55507 ( .A(n55544), .B(n55545), .Z(n55386) );
  AND U55508 ( .A(n2294), .B(n55546), .Z(n55545) );
  XNOR U55509 ( .A(n55547), .B(n55544), .Z(n55546) );
  XOR U55510 ( .A(n55387), .B(n55540), .Z(n55542) );
  XOR U55511 ( .A(n55548), .B(n55549), .Z(n55387) );
  AND U55512 ( .A(n2302), .B(n55507), .Z(n55549) );
  XOR U55513 ( .A(n55548), .B(n55505), .Z(n55507) );
  XOR U55514 ( .A(n55464), .B(n55550), .Z(n55540) );
  AND U55515 ( .A(n55466), .B(n55551), .Z(n55550) );
  XNOR U55516 ( .A(n55464), .B(n55434), .Z(n55551) );
  IV U55517 ( .A(n55437), .Z(n55434) );
  XOR U55518 ( .A(n55552), .B(n55553), .Z(n55437) );
  AND U55519 ( .A(n2294), .B(n55554), .Z(n55553) );
  XOR U55520 ( .A(n55555), .B(n55552), .Z(n55554) );
  XOR U55521 ( .A(n55438), .B(n55464), .Z(n55466) );
  XOR U55522 ( .A(n55556), .B(n55557), .Z(n55438) );
  AND U55523 ( .A(n2302), .B(n55517), .Z(n55557) );
  XOR U55524 ( .A(n55556), .B(n55515), .Z(n55517) );
  AND U55525 ( .A(n55518), .B(n55448), .Z(n55464) );
  XNOR U55526 ( .A(n55558), .B(n55559), .Z(n55448) );
  AND U55527 ( .A(n2294), .B(n55560), .Z(n55559) );
  XNOR U55528 ( .A(n55561), .B(n55558), .Z(n55560) );
  XNOR U55529 ( .A(n55562), .B(n55563), .Z(n2294) );
  AND U55530 ( .A(n55564), .B(n55565), .Z(n55563) );
  XOR U55531 ( .A(n55527), .B(n55562), .Z(n55565) );
  AND U55532 ( .A(n55566), .B(n55567), .Z(n55527) );
  XNOR U55533 ( .A(n55524), .B(n55562), .Z(n55564) );
  XNOR U55534 ( .A(n55568), .B(n55569), .Z(n55524) );
  AND U55535 ( .A(n2298), .B(n55570), .Z(n55569) );
  XNOR U55536 ( .A(n55571), .B(n55572), .Z(n55570) );
  XOR U55537 ( .A(n55573), .B(n55574), .Z(n55562) );
  AND U55538 ( .A(n55575), .B(n55576), .Z(n55574) );
  XNOR U55539 ( .A(n55573), .B(n55566), .Z(n55576) );
  IV U55540 ( .A(n55537), .Z(n55566) );
  XOR U55541 ( .A(n55577), .B(n55578), .Z(n55537) );
  XOR U55542 ( .A(n55579), .B(n55567), .Z(n55578) );
  AND U55543 ( .A(n55547), .B(n55580), .Z(n55567) );
  AND U55544 ( .A(n55581), .B(n55582), .Z(n55579) );
  XOR U55545 ( .A(n55583), .B(n55577), .Z(n55581) );
  XNOR U55546 ( .A(n55534), .B(n55573), .Z(n55575) );
  XNOR U55547 ( .A(n55584), .B(n55585), .Z(n55534) );
  AND U55548 ( .A(n2298), .B(n55586), .Z(n55585) );
  XNOR U55549 ( .A(n55587), .B(n55588), .Z(n55586) );
  XOR U55550 ( .A(n55589), .B(n55590), .Z(n55573) );
  AND U55551 ( .A(n55591), .B(n55592), .Z(n55590) );
  XNOR U55552 ( .A(n55589), .B(n55547), .Z(n55592) );
  XOR U55553 ( .A(n55593), .B(n55582), .Z(n55547) );
  XNOR U55554 ( .A(n55594), .B(n55577), .Z(n55582) );
  XOR U55555 ( .A(n55595), .B(n55596), .Z(n55577) );
  AND U55556 ( .A(n55597), .B(n55598), .Z(n55596) );
  XOR U55557 ( .A(n55599), .B(n55595), .Z(n55597) );
  XNOR U55558 ( .A(n55600), .B(n55601), .Z(n55594) );
  AND U55559 ( .A(n55602), .B(n55603), .Z(n55601) );
  XOR U55560 ( .A(n55600), .B(n55604), .Z(n55602) );
  XNOR U55561 ( .A(n55583), .B(n55580), .Z(n55593) );
  AND U55562 ( .A(n55605), .B(n55606), .Z(n55580) );
  XOR U55563 ( .A(n55607), .B(n55608), .Z(n55583) );
  AND U55564 ( .A(n55609), .B(n55610), .Z(n55608) );
  XOR U55565 ( .A(n55607), .B(n55611), .Z(n55609) );
  XNOR U55566 ( .A(n55544), .B(n55589), .Z(n55591) );
  XNOR U55567 ( .A(n55612), .B(n55613), .Z(n55544) );
  AND U55568 ( .A(n2298), .B(n55614), .Z(n55613) );
  XNOR U55569 ( .A(n55615), .B(n55616), .Z(n55614) );
  XOR U55570 ( .A(n55617), .B(n55618), .Z(n55589) );
  AND U55571 ( .A(n55619), .B(n55620), .Z(n55618) );
  XNOR U55572 ( .A(n55617), .B(n55605), .Z(n55620) );
  IV U55573 ( .A(n55555), .Z(n55605) );
  XNOR U55574 ( .A(n55621), .B(n55598), .Z(n55555) );
  XNOR U55575 ( .A(n55622), .B(n55604), .Z(n55598) );
  XNOR U55576 ( .A(n55623), .B(n55624), .Z(n55604) );
  NOR U55577 ( .A(n55625), .B(n55626), .Z(n55624) );
  XOR U55578 ( .A(n55623), .B(n55627), .Z(n55625) );
  XNOR U55579 ( .A(n55603), .B(n55595), .Z(n55622) );
  XOR U55580 ( .A(n55628), .B(n55629), .Z(n55595) );
  AND U55581 ( .A(n55630), .B(n55631), .Z(n55629) );
  XOR U55582 ( .A(n55628), .B(n55632), .Z(n55630) );
  XNOR U55583 ( .A(n55633), .B(n55600), .Z(n55603) );
  XOR U55584 ( .A(n55634), .B(n55635), .Z(n55600) );
  AND U55585 ( .A(n55636), .B(n55637), .Z(n55635) );
  XNOR U55586 ( .A(n55638), .B(n55639), .Z(n55636) );
  IV U55587 ( .A(n55634), .Z(n55638) );
  XNOR U55588 ( .A(n55640), .B(n55641), .Z(n55633) );
  NOR U55589 ( .A(n55642), .B(n55643), .Z(n55641) );
  XNOR U55590 ( .A(n55640), .B(n55644), .Z(n55642) );
  XNOR U55591 ( .A(n55599), .B(n55606), .Z(n55621) );
  NOR U55592 ( .A(n55561), .B(n55645), .Z(n55606) );
  XOR U55593 ( .A(n55611), .B(n55610), .Z(n55599) );
  XNOR U55594 ( .A(n55646), .B(n55607), .Z(n55610) );
  XOR U55595 ( .A(n55647), .B(n55648), .Z(n55607) );
  AND U55596 ( .A(n55649), .B(n55650), .Z(n55648) );
  XNOR U55597 ( .A(n55651), .B(n55652), .Z(n55649) );
  IV U55598 ( .A(n55647), .Z(n55651) );
  XNOR U55599 ( .A(n55653), .B(n55654), .Z(n55646) );
  NOR U55600 ( .A(n55655), .B(n55656), .Z(n55654) );
  XNOR U55601 ( .A(n55653), .B(n55657), .Z(n55655) );
  XOR U55602 ( .A(n55658), .B(n55659), .Z(n55611) );
  NOR U55603 ( .A(n55660), .B(n55661), .Z(n55659) );
  XNOR U55604 ( .A(n55658), .B(n55662), .Z(n55660) );
  XNOR U55605 ( .A(n55552), .B(n55617), .Z(n55619) );
  XNOR U55606 ( .A(n55663), .B(n55664), .Z(n55552) );
  AND U55607 ( .A(n2298), .B(n55665), .Z(n55664) );
  XNOR U55608 ( .A(n55666), .B(n55667), .Z(n55665) );
  AND U55609 ( .A(n55558), .B(n55561), .Z(n55617) );
  XOR U55610 ( .A(n55668), .B(n55645), .Z(n55561) );
  XNOR U55611 ( .A(p_input[1872]), .B(p_input[2048]), .Z(n55645) );
  XNOR U55612 ( .A(n55632), .B(n55631), .Z(n55668) );
  XNOR U55613 ( .A(n55669), .B(n55639), .Z(n55631) );
  XNOR U55614 ( .A(n55627), .B(n55626), .Z(n55639) );
  XNOR U55615 ( .A(n55670), .B(n55623), .Z(n55626) );
  XNOR U55616 ( .A(p_input[1882]), .B(p_input[2058]), .Z(n55623) );
  XOR U55617 ( .A(p_input[1883]), .B(n29030), .Z(n55670) );
  XOR U55618 ( .A(p_input[1884]), .B(p_input[2060]), .Z(n55627) );
  XOR U55619 ( .A(n55637), .B(n55671), .Z(n55669) );
  IV U55620 ( .A(n55628), .Z(n55671) );
  XOR U55621 ( .A(p_input[1873]), .B(p_input[2049]), .Z(n55628) );
  XNOR U55622 ( .A(n55672), .B(n55644), .Z(n55637) );
  XNOR U55623 ( .A(p_input[1887]), .B(n29033), .Z(n55644) );
  XOR U55624 ( .A(n55634), .B(n55643), .Z(n55672) );
  XOR U55625 ( .A(n55673), .B(n55640), .Z(n55643) );
  XOR U55626 ( .A(p_input[1885]), .B(p_input[2061]), .Z(n55640) );
  XOR U55627 ( .A(p_input[1886]), .B(n29035), .Z(n55673) );
  XOR U55628 ( .A(p_input[1881]), .B(p_input[2057]), .Z(n55634) );
  XOR U55629 ( .A(n55652), .B(n55650), .Z(n55632) );
  XNOR U55630 ( .A(n55674), .B(n55657), .Z(n55650) );
  XOR U55631 ( .A(p_input[1880]), .B(p_input[2056]), .Z(n55657) );
  XOR U55632 ( .A(n55647), .B(n55656), .Z(n55674) );
  XOR U55633 ( .A(n55675), .B(n55653), .Z(n55656) );
  XOR U55634 ( .A(p_input[1878]), .B(p_input[2054]), .Z(n55653) );
  XOR U55635 ( .A(p_input[1879]), .B(n30404), .Z(n55675) );
  XOR U55636 ( .A(p_input[1874]), .B(p_input[2050]), .Z(n55647) );
  XNOR U55637 ( .A(n55662), .B(n55661), .Z(n55652) );
  XOR U55638 ( .A(n55676), .B(n55658), .Z(n55661) );
  XOR U55639 ( .A(p_input[1875]), .B(p_input[2051]), .Z(n55658) );
  XOR U55640 ( .A(p_input[1876]), .B(n30406), .Z(n55676) );
  XOR U55641 ( .A(p_input[1877]), .B(p_input[2053]), .Z(n55662) );
  XNOR U55642 ( .A(n55677), .B(n55678), .Z(n55558) );
  AND U55643 ( .A(n2298), .B(n55679), .Z(n55678) );
  XNOR U55644 ( .A(n55680), .B(n55681), .Z(n2298) );
  AND U55645 ( .A(n55682), .B(n55683), .Z(n55681) );
  XOR U55646 ( .A(n55572), .B(n55680), .Z(n55683) );
  XNOR U55647 ( .A(n55684), .B(n55680), .Z(n55682) );
  XOR U55648 ( .A(n55685), .B(n55686), .Z(n55680) );
  AND U55649 ( .A(n55687), .B(n55688), .Z(n55686) );
  XOR U55650 ( .A(n55587), .B(n55685), .Z(n55688) );
  XOR U55651 ( .A(n55685), .B(n55588), .Z(n55687) );
  XOR U55652 ( .A(n55689), .B(n55690), .Z(n55685) );
  AND U55653 ( .A(n55691), .B(n55692), .Z(n55690) );
  XOR U55654 ( .A(n55615), .B(n55689), .Z(n55692) );
  XOR U55655 ( .A(n55689), .B(n55616), .Z(n55691) );
  XOR U55656 ( .A(n55693), .B(n55694), .Z(n55689) );
  AND U55657 ( .A(n55695), .B(n55696), .Z(n55694) );
  XOR U55658 ( .A(n55693), .B(n55666), .Z(n55696) );
  XNOR U55659 ( .A(n55697), .B(n55698), .Z(n55518) );
  AND U55660 ( .A(n2302), .B(n55699), .Z(n55698) );
  XNOR U55661 ( .A(n55700), .B(n55701), .Z(n2302) );
  AND U55662 ( .A(n55702), .B(n55703), .Z(n55701) );
  XOR U55663 ( .A(n55700), .B(n55528), .Z(n55703) );
  XNOR U55664 ( .A(n55700), .B(n55488), .Z(n55702) );
  XOR U55665 ( .A(n55704), .B(n55705), .Z(n55700) );
  AND U55666 ( .A(n55706), .B(n55707), .Z(n55705) );
  XOR U55667 ( .A(n55704), .B(n55496), .Z(n55706) );
  XOR U55668 ( .A(n55708), .B(n55709), .Z(n55479) );
  AND U55669 ( .A(n2306), .B(n55699), .Z(n55709) );
  XNOR U55670 ( .A(n55697), .B(n55708), .Z(n55699) );
  XNOR U55671 ( .A(n55710), .B(n55711), .Z(n2306) );
  AND U55672 ( .A(n55712), .B(n55713), .Z(n55711) );
  XNOR U55673 ( .A(n55714), .B(n55710), .Z(n55713) );
  IV U55674 ( .A(n55528), .Z(n55714) );
  XOR U55675 ( .A(n55684), .B(n55715), .Z(n55528) );
  AND U55676 ( .A(n2309), .B(n55716), .Z(n55715) );
  XOR U55677 ( .A(n55571), .B(n55568), .Z(n55716) );
  IV U55678 ( .A(n55684), .Z(n55571) );
  XNOR U55679 ( .A(n55488), .B(n55710), .Z(n55712) );
  XOR U55680 ( .A(n55717), .B(n55718), .Z(n55488) );
  AND U55681 ( .A(n2325), .B(n55719), .Z(n55718) );
  XOR U55682 ( .A(n55704), .B(n55720), .Z(n55710) );
  AND U55683 ( .A(n55721), .B(n55707), .Z(n55720) );
  XNOR U55684 ( .A(n55538), .B(n55704), .Z(n55707) );
  XOR U55685 ( .A(n55588), .B(n55722), .Z(n55538) );
  AND U55686 ( .A(n2309), .B(n55723), .Z(n55722) );
  XOR U55687 ( .A(n55584), .B(n55588), .Z(n55723) );
  XNOR U55688 ( .A(n55724), .B(n55704), .Z(n55721) );
  IV U55689 ( .A(n55496), .Z(n55724) );
  XOR U55690 ( .A(n55725), .B(n55726), .Z(n55496) );
  AND U55691 ( .A(n2325), .B(n55727), .Z(n55726) );
  XOR U55692 ( .A(n55728), .B(n55729), .Z(n55704) );
  AND U55693 ( .A(n55730), .B(n55731), .Z(n55729) );
  XNOR U55694 ( .A(n55548), .B(n55728), .Z(n55731) );
  XOR U55695 ( .A(n55616), .B(n55732), .Z(n55548) );
  AND U55696 ( .A(n2309), .B(n55733), .Z(n55732) );
  XOR U55697 ( .A(n55612), .B(n55616), .Z(n55733) );
  XOR U55698 ( .A(n55728), .B(n55505), .Z(n55730) );
  XOR U55699 ( .A(n55734), .B(n55735), .Z(n55505) );
  AND U55700 ( .A(n2325), .B(n55736), .Z(n55735) );
  XOR U55701 ( .A(n55737), .B(n55738), .Z(n55728) );
  AND U55702 ( .A(n55739), .B(n55740), .Z(n55738) );
  XNOR U55703 ( .A(n55737), .B(n55556), .Z(n55740) );
  XOR U55704 ( .A(n55667), .B(n55741), .Z(n55556) );
  AND U55705 ( .A(n2309), .B(n55742), .Z(n55741) );
  XOR U55706 ( .A(n55663), .B(n55667), .Z(n55742) );
  XNOR U55707 ( .A(n55743), .B(n55737), .Z(n55739) );
  IV U55708 ( .A(n55515), .Z(n55743) );
  XOR U55709 ( .A(n55744), .B(n55745), .Z(n55515) );
  AND U55710 ( .A(n2325), .B(n55746), .Z(n55745) );
  AND U55711 ( .A(n55708), .B(n55697), .Z(n55737) );
  XNOR U55712 ( .A(n55747), .B(n55748), .Z(n55697) );
  AND U55713 ( .A(n2309), .B(n55679), .Z(n55748) );
  XNOR U55714 ( .A(n55677), .B(n55747), .Z(n55679) );
  XNOR U55715 ( .A(n55749), .B(n55750), .Z(n2309) );
  AND U55716 ( .A(n55751), .B(n55752), .Z(n55750) );
  XNOR U55717 ( .A(n55749), .B(n55568), .Z(n55752) );
  IV U55718 ( .A(n55572), .Z(n55568) );
  XOR U55719 ( .A(n55753), .B(n55754), .Z(n55572) );
  AND U55720 ( .A(n2313), .B(n55755), .Z(n55754) );
  XOR U55721 ( .A(n55756), .B(n55753), .Z(n55755) );
  XNOR U55722 ( .A(n55749), .B(n55684), .Z(n55751) );
  XOR U55723 ( .A(n55757), .B(n55758), .Z(n55684) );
  AND U55724 ( .A(n2321), .B(n55719), .Z(n55758) );
  XOR U55725 ( .A(n55717), .B(n55757), .Z(n55719) );
  XOR U55726 ( .A(n55759), .B(n55760), .Z(n55749) );
  AND U55727 ( .A(n55761), .B(n55762), .Z(n55760) );
  XNOR U55728 ( .A(n55759), .B(n55584), .Z(n55762) );
  IV U55729 ( .A(n55587), .Z(n55584) );
  XOR U55730 ( .A(n55763), .B(n55764), .Z(n55587) );
  AND U55731 ( .A(n2313), .B(n55765), .Z(n55764) );
  XOR U55732 ( .A(n55766), .B(n55763), .Z(n55765) );
  XOR U55733 ( .A(n55588), .B(n55759), .Z(n55761) );
  XOR U55734 ( .A(n55767), .B(n55768), .Z(n55588) );
  AND U55735 ( .A(n2321), .B(n55727), .Z(n55768) );
  XOR U55736 ( .A(n55767), .B(n55725), .Z(n55727) );
  XOR U55737 ( .A(n55769), .B(n55770), .Z(n55759) );
  AND U55738 ( .A(n55771), .B(n55772), .Z(n55770) );
  XNOR U55739 ( .A(n55769), .B(n55612), .Z(n55772) );
  IV U55740 ( .A(n55615), .Z(n55612) );
  XOR U55741 ( .A(n55773), .B(n55774), .Z(n55615) );
  AND U55742 ( .A(n2313), .B(n55775), .Z(n55774) );
  XNOR U55743 ( .A(n55776), .B(n55773), .Z(n55775) );
  XOR U55744 ( .A(n55616), .B(n55769), .Z(n55771) );
  XOR U55745 ( .A(n55777), .B(n55778), .Z(n55616) );
  AND U55746 ( .A(n2321), .B(n55736), .Z(n55778) );
  XOR U55747 ( .A(n55777), .B(n55734), .Z(n55736) );
  XOR U55748 ( .A(n55693), .B(n55779), .Z(n55769) );
  AND U55749 ( .A(n55695), .B(n55780), .Z(n55779) );
  XNOR U55750 ( .A(n55693), .B(n55663), .Z(n55780) );
  IV U55751 ( .A(n55666), .Z(n55663) );
  XOR U55752 ( .A(n55781), .B(n55782), .Z(n55666) );
  AND U55753 ( .A(n2313), .B(n55783), .Z(n55782) );
  XOR U55754 ( .A(n55784), .B(n55781), .Z(n55783) );
  XOR U55755 ( .A(n55667), .B(n55693), .Z(n55695) );
  XOR U55756 ( .A(n55785), .B(n55786), .Z(n55667) );
  AND U55757 ( .A(n2321), .B(n55746), .Z(n55786) );
  XOR U55758 ( .A(n55785), .B(n55744), .Z(n55746) );
  AND U55759 ( .A(n55747), .B(n55677), .Z(n55693) );
  XNOR U55760 ( .A(n55787), .B(n55788), .Z(n55677) );
  AND U55761 ( .A(n2313), .B(n55789), .Z(n55788) );
  XNOR U55762 ( .A(n55790), .B(n55787), .Z(n55789) );
  XNOR U55763 ( .A(n55791), .B(n55792), .Z(n2313) );
  AND U55764 ( .A(n55793), .B(n55794), .Z(n55792) );
  XOR U55765 ( .A(n55756), .B(n55791), .Z(n55794) );
  AND U55766 ( .A(n55795), .B(n55796), .Z(n55756) );
  XNOR U55767 ( .A(n55753), .B(n55791), .Z(n55793) );
  XNOR U55768 ( .A(n55797), .B(n55798), .Z(n55753) );
  AND U55769 ( .A(n2317), .B(n55799), .Z(n55798) );
  XNOR U55770 ( .A(n55800), .B(n55801), .Z(n55799) );
  XOR U55771 ( .A(n55802), .B(n55803), .Z(n55791) );
  AND U55772 ( .A(n55804), .B(n55805), .Z(n55803) );
  XNOR U55773 ( .A(n55802), .B(n55795), .Z(n55805) );
  IV U55774 ( .A(n55766), .Z(n55795) );
  XOR U55775 ( .A(n55806), .B(n55807), .Z(n55766) );
  XOR U55776 ( .A(n55808), .B(n55796), .Z(n55807) );
  AND U55777 ( .A(n55776), .B(n55809), .Z(n55796) );
  AND U55778 ( .A(n55810), .B(n55811), .Z(n55808) );
  XOR U55779 ( .A(n55812), .B(n55806), .Z(n55810) );
  XNOR U55780 ( .A(n55763), .B(n55802), .Z(n55804) );
  XNOR U55781 ( .A(n55813), .B(n55814), .Z(n55763) );
  AND U55782 ( .A(n2317), .B(n55815), .Z(n55814) );
  XNOR U55783 ( .A(n55816), .B(n55817), .Z(n55815) );
  XOR U55784 ( .A(n55818), .B(n55819), .Z(n55802) );
  AND U55785 ( .A(n55820), .B(n55821), .Z(n55819) );
  XNOR U55786 ( .A(n55818), .B(n55776), .Z(n55821) );
  XOR U55787 ( .A(n55822), .B(n55811), .Z(n55776) );
  XNOR U55788 ( .A(n55823), .B(n55806), .Z(n55811) );
  XOR U55789 ( .A(n55824), .B(n55825), .Z(n55806) );
  AND U55790 ( .A(n55826), .B(n55827), .Z(n55825) );
  XOR U55791 ( .A(n55828), .B(n55824), .Z(n55826) );
  XNOR U55792 ( .A(n55829), .B(n55830), .Z(n55823) );
  AND U55793 ( .A(n55831), .B(n55832), .Z(n55830) );
  XOR U55794 ( .A(n55829), .B(n55833), .Z(n55831) );
  XNOR U55795 ( .A(n55812), .B(n55809), .Z(n55822) );
  AND U55796 ( .A(n55834), .B(n55835), .Z(n55809) );
  XOR U55797 ( .A(n55836), .B(n55837), .Z(n55812) );
  AND U55798 ( .A(n55838), .B(n55839), .Z(n55837) );
  XOR U55799 ( .A(n55836), .B(n55840), .Z(n55838) );
  XNOR U55800 ( .A(n55773), .B(n55818), .Z(n55820) );
  XNOR U55801 ( .A(n55841), .B(n55842), .Z(n55773) );
  AND U55802 ( .A(n2317), .B(n55843), .Z(n55842) );
  XNOR U55803 ( .A(n55844), .B(n55845), .Z(n55843) );
  XOR U55804 ( .A(n55846), .B(n55847), .Z(n55818) );
  AND U55805 ( .A(n55848), .B(n55849), .Z(n55847) );
  XNOR U55806 ( .A(n55846), .B(n55834), .Z(n55849) );
  IV U55807 ( .A(n55784), .Z(n55834) );
  XNOR U55808 ( .A(n55850), .B(n55827), .Z(n55784) );
  XNOR U55809 ( .A(n55851), .B(n55833), .Z(n55827) );
  XNOR U55810 ( .A(n55852), .B(n55853), .Z(n55833) );
  NOR U55811 ( .A(n55854), .B(n55855), .Z(n55853) );
  XOR U55812 ( .A(n55852), .B(n55856), .Z(n55854) );
  XNOR U55813 ( .A(n55832), .B(n55824), .Z(n55851) );
  XOR U55814 ( .A(n55857), .B(n55858), .Z(n55824) );
  AND U55815 ( .A(n55859), .B(n55860), .Z(n55858) );
  XOR U55816 ( .A(n55857), .B(n55861), .Z(n55859) );
  XNOR U55817 ( .A(n55862), .B(n55829), .Z(n55832) );
  XOR U55818 ( .A(n55863), .B(n55864), .Z(n55829) );
  AND U55819 ( .A(n55865), .B(n55866), .Z(n55864) );
  XNOR U55820 ( .A(n55867), .B(n55868), .Z(n55865) );
  IV U55821 ( .A(n55863), .Z(n55867) );
  XNOR U55822 ( .A(n55869), .B(n55870), .Z(n55862) );
  NOR U55823 ( .A(n55871), .B(n55872), .Z(n55870) );
  XNOR U55824 ( .A(n55869), .B(n55873), .Z(n55871) );
  XNOR U55825 ( .A(n55828), .B(n55835), .Z(n55850) );
  NOR U55826 ( .A(n55790), .B(n55874), .Z(n55835) );
  XOR U55827 ( .A(n55840), .B(n55839), .Z(n55828) );
  XNOR U55828 ( .A(n55875), .B(n55836), .Z(n55839) );
  XOR U55829 ( .A(n55876), .B(n55877), .Z(n55836) );
  AND U55830 ( .A(n55878), .B(n55879), .Z(n55877) );
  XNOR U55831 ( .A(n55880), .B(n55881), .Z(n55878) );
  IV U55832 ( .A(n55876), .Z(n55880) );
  XNOR U55833 ( .A(n55882), .B(n55883), .Z(n55875) );
  NOR U55834 ( .A(n55884), .B(n55885), .Z(n55883) );
  XNOR U55835 ( .A(n55882), .B(n55886), .Z(n55884) );
  XOR U55836 ( .A(n55887), .B(n55888), .Z(n55840) );
  NOR U55837 ( .A(n55889), .B(n55890), .Z(n55888) );
  XNOR U55838 ( .A(n55887), .B(n55891), .Z(n55889) );
  XNOR U55839 ( .A(n55781), .B(n55846), .Z(n55848) );
  XNOR U55840 ( .A(n55892), .B(n55893), .Z(n55781) );
  AND U55841 ( .A(n2317), .B(n55894), .Z(n55893) );
  XNOR U55842 ( .A(n55895), .B(n55896), .Z(n55894) );
  AND U55843 ( .A(n55787), .B(n55790), .Z(n55846) );
  XOR U55844 ( .A(n55897), .B(n55874), .Z(n55790) );
  XNOR U55845 ( .A(p_input[1888]), .B(p_input[2048]), .Z(n55874) );
  XNOR U55846 ( .A(n55861), .B(n55860), .Z(n55897) );
  XNOR U55847 ( .A(n55898), .B(n55868), .Z(n55860) );
  XNOR U55848 ( .A(n55856), .B(n55855), .Z(n55868) );
  XNOR U55849 ( .A(n55899), .B(n55852), .Z(n55855) );
  XNOR U55850 ( .A(p_input[1898]), .B(p_input[2058]), .Z(n55852) );
  XOR U55851 ( .A(p_input[1899]), .B(n29030), .Z(n55899) );
  XOR U55852 ( .A(p_input[1900]), .B(p_input[2060]), .Z(n55856) );
  XOR U55853 ( .A(n55866), .B(n55900), .Z(n55898) );
  IV U55854 ( .A(n55857), .Z(n55900) );
  XOR U55855 ( .A(p_input[1889]), .B(p_input[2049]), .Z(n55857) );
  XNOR U55856 ( .A(n55901), .B(n55873), .Z(n55866) );
  XNOR U55857 ( .A(p_input[1903]), .B(n29033), .Z(n55873) );
  XOR U55858 ( .A(n55863), .B(n55872), .Z(n55901) );
  XOR U55859 ( .A(n55902), .B(n55869), .Z(n55872) );
  XOR U55860 ( .A(p_input[1901]), .B(p_input[2061]), .Z(n55869) );
  XOR U55861 ( .A(p_input[1902]), .B(n29035), .Z(n55902) );
  XOR U55862 ( .A(p_input[1897]), .B(p_input[2057]), .Z(n55863) );
  XOR U55863 ( .A(n55881), .B(n55879), .Z(n55861) );
  XNOR U55864 ( .A(n55903), .B(n55886), .Z(n55879) );
  XOR U55865 ( .A(p_input[1896]), .B(p_input[2056]), .Z(n55886) );
  XOR U55866 ( .A(n55876), .B(n55885), .Z(n55903) );
  XOR U55867 ( .A(n55904), .B(n55882), .Z(n55885) );
  XOR U55868 ( .A(p_input[1894]), .B(p_input[2054]), .Z(n55882) );
  XOR U55869 ( .A(p_input[1895]), .B(n30404), .Z(n55904) );
  XOR U55870 ( .A(p_input[1890]), .B(p_input[2050]), .Z(n55876) );
  XNOR U55871 ( .A(n55891), .B(n55890), .Z(n55881) );
  XOR U55872 ( .A(n55905), .B(n55887), .Z(n55890) );
  XOR U55873 ( .A(p_input[1891]), .B(p_input[2051]), .Z(n55887) );
  XOR U55874 ( .A(p_input[1892]), .B(n30406), .Z(n55905) );
  XOR U55875 ( .A(p_input[1893]), .B(p_input[2053]), .Z(n55891) );
  XNOR U55876 ( .A(n55906), .B(n55907), .Z(n55787) );
  AND U55877 ( .A(n2317), .B(n55908), .Z(n55907) );
  XNOR U55878 ( .A(n55909), .B(n55910), .Z(n2317) );
  AND U55879 ( .A(n55911), .B(n55912), .Z(n55910) );
  XOR U55880 ( .A(n55801), .B(n55909), .Z(n55912) );
  XNOR U55881 ( .A(n55913), .B(n55909), .Z(n55911) );
  XOR U55882 ( .A(n55914), .B(n55915), .Z(n55909) );
  AND U55883 ( .A(n55916), .B(n55917), .Z(n55915) );
  XOR U55884 ( .A(n55816), .B(n55914), .Z(n55917) );
  XOR U55885 ( .A(n55914), .B(n55817), .Z(n55916) );
  XOR U55886 ( .A(n55918), .B(n55919), .Z(n55914) );
  AND U55887 ( .A(n55920), .B(n55921), .Z(n55919) );
  XOR U55888 ( .A(n55844), .B(n55918), .Z(n55921) );
  XOR U55889 ( .A(n55918), .B(n55845), .Z(n55920) );
  XOR U55890 ( .A(n55922), .B(n55923), .Z(n55918) );
  AND U55891 ( .A(n55924), .B(n55925), .Z(n55923) );
  XOR U55892 ( .A(n55922), .B(n55895), .Z(n55925) );
  XNOR U55893 ( .A(n55926), .B(n55927), .Z(n55747) );
  AND U55894 ( .A(n2321), .B(n55928), .Z(n55927) );
  XNOR U55895 ( .A(n55929), .B(n55930), .Z(n2321) );
  AND U55896 ( .A(n55931), .B(n55932), .Z(n55930) );
  XOR U55897 ( .A(n55929), .B(n55757), .Z(n55932) );
  XNOR U55898 ( .A(n55929), .B(n55717), .Z(n55931) );
  XOR U55899 ( .A(n55933), .B(n55934), .Z(n55929) );
  AND U55900 ( .A(n55935), .B(n55936), .Z(n55934) );
  XOR U55901 ( .A(n55933), .B(n55725), .Z(n55935) );
  XOR U55902 ( .A(n55937), .B(n55938), .Z(n55708) );
  AND U55903 ( .A(n2325), .B(n55928), .Z(n55938) );
  XNOR U55904 ( .A(n55926), .B(n55937), .Z(n55928) );
  XNOR U55905 ( .A(n55939), .B(n55940), .Z(n2325) );
  AND U55906 ( .A(n55941), .B(n55942), .Z(n55940) );
  XNOR U55907 ( .A(n55943), .B(n55939), .Z(n55942) );
  IV U55908 ( .A(n55757), .Z(n55943) );
  XOR U55909 ( .A(n55913), .B(n55944), .Z(n55757) );
  AND U55910 ( .A(n2328), .B(n55945), .Z(n55944) );
  XOR U55911 ( .A(n55800), .B(n55797), .Z(n55945) );
  IV U55912 ( .A(n55913), .Z(n55800) );
  XNOR U55913 ( .A(n55717), .B(n55939), .Z(n55941) );
  XOR U55914 ( .A(n55946), .B(n55947), .Z(n55717) );
  AND U55915 ( .A(n2344), .B(n55948), .Z(n55947) );
  XOR U55916 ( .A(n55933), .B(n55949), .Z(n55939) );
  AND U55917 ( .A(n55950), .B(n55936), .Z(n55949) );
  XNOR U55918 ( .A(n55767), .B(n55933), .Z(n55936) );
  XOR U55919 ( .A(n55817), .B(n55951), .Z(n55767) );
  AND U55920 ( .A(n2328), .B(n55952), .Z(n55951) );
  XOR U55921 ( .A(n55813), .B(n55817), .Z(n55952) );
  XNOR U55922 ( .A(n55953), .B(n55933), .Z(n55950) );
  IV U55923 ( .A(n55725), .Z(n55953) );
  XOR U55924 ( .A(n55954), .B(n55955), .Z(n55725) );
  AND U55925 ( .A(n2344), .B(n55956), .Z(n55955) );
  XOR U55926 ( .A(n55957), .B(n55958), .Z(n55933) );
  AND U55927 ( .A(n55959), .B(n55960), .Z(n55958) );
  XNOR U55928 ( .A(n55777), .B(n55957), .Z(n55960) );
  XOR U55929 ( .A(n55845), .B(n55961), .Z(n55777) );
  AND U55930 ( .A(n2328), .B(n55962), .Z(n55961) );
  XOR U55931 ( .A(n55841), .B(n55845), .Z(n55962) );
  XOR U55932 ( .A(n55957), .B(n55734), .Z(n55959) );
  XOR U55933 ( .A(n55963), .B(n55964), .Z(n55734) );
  AND U55934 ( .A(n2344), .B(n55965), .Z(n55964) );
  XOR U55935 ( .A(n55966), .B(n55967), .Z(n55957) );
  AND U55936 ( .A(n55968), .B(n55969), .Z(n55967) );
  XNOR U55937 ( .A(n55966), .B(n55785), .Z(n55969) );
  XOR U55938 ( .A(n55896), .B(n55970), .Z(n55785) );
  AND U55939 ( .A(n2328), .B(n55971), .Z(n55970) );
  XOR U55940 ( .A(n55892), .B(n55896), .Z(n55971) );
  XNOR U55941 ( .A(n55972), .B(n55966), .Z(n55968) );
  IV U55942 ( .A(n55744), .Z(n55972) );
  XOR U55943 ( .A(n55973), .B(n55974), .Z(n55744) );
  AND U55944 ( .A(n2344), .B(n55975), .Z(n55974) );
  AND U55945 ( .A(n55937), .B(n55926), .Z(n55966) );
  XNOR U55946 ( .A(n55976), .B(n55977), .Z(n55926) );
  AND U55947 ( .A(n2328), .B(n55908), .Z(n55977) );
  XNOR U55948 ( .A(n55906), .B(n55976), .Z(n55908) );
  XNOR U55949 ( .A(n55978), .B(n55979), .Z(n2328) );
  AND U55950 ( .A(n55980), .B(n55981), .Z(n55979) );
  XNOR U55951 ( .A(n55978), .B(n55797), .Z(n55981) );
  IV U55952 ( .A(n55801), .Z(n55797) );
  XOR U55953 ( .A(n55982), .B(n55983), .Z(n55801) );
  AND U55954 ( .A(n2332), .B(n55984), .Z(n55983) );
  XOR U55955 ( .A(n55985), .B(n55982), .Z(n55984) );
  XNOR U55956 ( .A(n55978), .B(n55913), .Z(n55980) );
  XOR U55957 ( .A(n55986), .B(n55987), .Z(n55913) );
  AND U55958 ( .A(n2340), .B(n55948), .Z(n55987) );
  XOR U55959 ( .A(n55946), .B(n55986), .Z(n55948) );
  XOR U55960 ( .A(n55988), .B(n55989), .Z(n55978) );
  AND U55961 ( .A(n55990), .B(n55991), .Z(n55989) );
  XNOR U55962 ( .A(n55988), .B(n55813), .Z(n55991) );
  IV U55963 ( .A(n55816), .Z(n55813) );
  XOR U55964 ( .A(n55992), .B(n55993), .Z(n55816) );
  AND U55965 ( .A(n2332), .B(n55994), .Z(n55993) );
  XOR U55966 ( .A(n55995), .B(n55992), .Z(n55994) );
  XOR U55967 ( .A(n55817), .B(n55988), .Z(n55990) );
  XOR U55968 ( .A(n55996), .B(n55997), .Z(n55817) );
  AND U55969 ( .A(n2340), .B(n55956), .Z(n55997) );
  XOR U55970 ( .A(n55996), .B(n55954), .Z(n55956) );
  XOR U55971 ( .A(n55998), .B(n55999), .Z(n55988) );
  AND U55972 ( .A(n56000), .B(n56001), .Z(n55999) );
  XNOR U55973 ( .A(n55998), .B(n55841), .Z(n56001) );
  IV U55974 ( .A(n55844), .Z(n55841) );
  XOR U55975 ( .A(n56002), .B(n56003), .Z(n55844) );
  AND U55976 ( .A(n2332), .B(n56004), .Z(n56003) );
  XNOR U55977 ( .A(n56005), .B(n56002), .Z(n56004) );
  XOR U55978 ( .A(n55845), .B(n55998), .Z(n56000) );
  XOR U55979 ( .A(n56006), .B(n56007), .Z(n55845) );
  AND U55980 ( .A(n2340), .B(n55965), .Z(n56007) );
  XOR U55981 ( .A(n56006), .B(n55963), .Z(n55965) );
  XOR U55982 ( .A(n55922), .B(n56008), .Z(n55998) );
  AND U55983 ( .A(n55924), .B(n56009), .Z(n56008) );
  XNOR U55984 ( .A(n55922), .B(n55892), .Z(n56009) );
  IV U55985 ( .A(n55895), .Z(n55892) );
  XOR U55986 ( .A(n56010), .B(n56011), .Z(n55895) );
  AND U55987 ( .A(n2332), .B(n56012), .Z(n56011) );
  XOR U55988 ( .A(n56013), .B(n56010), .Z(n56012) );
  XOR U55989 ( .A(n55896), .B(n55922), .Z(n55924) );
  XOR U55990 ( .A(n56014), .B(n56015), .Z(n55896) );
  AND U55991 ( .A(n2340), .B(n55975), .Z(n56015) );
  XOR U55992 ( .A(n56014), .B(n55973), .Z(n55975) );
  AND U55993 ( .A(n55976), .B(n55906), .Z(n55922) );
  XNOR U55994 ( .A(n56016), .B(n56017), .Z(n55906) );
  AND U55995 ( .A(n2332), .B(n56018), .Z(n56017) );
  XNOR U55996 ( .A(n56019), .B(n56016), .Z(n56018) );
  XNOR U55997 ( .A(n56020), .B(n56021), .Z(n2332) );
  AND U55998 ( .A(n56022), .B(n56023), .Z(n56021) );
  XOR U55999 ( .A(n55985), .B(n56020), .Z(n56023) );
  AND U56000 ( .A(n56024), .B(n56025), .Z(n55985) );
  XNOR U56001 ( .A(n55982), .B(n56020), .Z(n56022) );
  XNOR U56002 ( .A(n56026), .B(n56027), .Z(n55982) );
  AND U56003 ( .A(n2336), .B(n56028), .Z(n56027) );
  XNOR U56004 ( .A(n56029), .B(n56030), .Z(n56028) );
  XOR U56005 ( .A(n56031), .B(n56032), .Z(n56020) );
  AND U56006 ( .A(n56033), .B(n56034), .Z(n56032) );
  XNOR U56007 ( .A(n56031), .B(n56024), .Z(n56034) );
  IV U56008 ( .A(n55995), .Z(n56024) );
  XOR U56009 ( .A(n56035), .B(n56036), .Z(n55995) );
  XOR U56010 ( .A(n56037), .B(n56025), .Z(n56036) );
  AND U56011 ( .A(n56005), .B(n56038), .Z(n56025) );
  AND U56012 ( .A(n56039), .B(n56040), .Z(n56037) );
  XOR U56013 ( .A(n56041), .B(n56035), .Z(n56039) );
  XNOR U56014 ( .A(n55992), .B(n56031), .Z(n56033) );
  XNOR U56015 ( .A(n56042), .B(n56043), .Z(n55992) );
  AND U56016 ( .A(n2336), .B(n56044), .Z(n56043) );
  XNOR U56017 ( .A(n56045), .B(n56046), .Z(n56044) );
  XOR U56018 ( .A(n56047), .B(n56048), .Z(n56031) );
  AND U56019 ( .A(n56049), .B(n56050), .Z(n56048) );
  XNOR U56020 ( .A(n56047), .B(n56005), .Z(n56050) );
  XOR U56021 ( .A(n56051), .B(n56040), .Z(n56005) );
  XNOR U56022 ( .A(n56052), .B(n56035), .Z(n56040) );
  XOR U56023 ( .A(n56053), .B(n56054), .Z(n56035) );
  AND U56024 ( .A(n56055), .B(n56056), .Z(n56054) );
  XOR U56025 ( .A(n56057), .B(n56053), .Z(n56055) );
  XNOR U56026 ( .A(n56058), .B(n56059), .Z(n56052) );
  AND U56027 ( .A(n56060), .B(n56061), .Z(n56059) );
  XOR U56028 ( .A(n56058), .B(n56062), .Z(n56060) );
  XNOR U56029 ( .A(n56041), .B(n56038), .Z(n56051) );
  AND U56030 ( .A(n56063), .B(n56064), .Z(n56038) );
  XOR U56031 ( .A(n56065), .B(n56066), .Z(n56041) );
  AND U56032 ( .A(n56067), .B(n56068), .Z(n56066) );
  XOR U56033 ( .A(n56065), .B(n56069), .Z(n56067) );
  XNOR U56034 ( .A(n56002), .B(n56047), .Z(n56049) );
  XNOR U56035 ( .A(n56070), .B(n56071), .Z(n56002) );
  AND U56036 ( .A(n2336), .B(n56072), .Z(n56071) );
  XNOR U56037 ( .A(n56073), .B(n56074), .Z(n56072) );
  XOR U56038 ( .A(n56075), .B(n56076), .Z(n56047) );
  AND U56039 ( .A(n56077), .B(n56078), .Z(n56076) );
  XNOR U56040 ( .A(n56075), .B(n56063), .Z(n56078) );
  IV U56041 ( .A(n56013), .Z(n56063) );
  XNOR U56042 ( .A(n56079), .B(n56056), .Z(n56013) );
  XNOR U56043 ( .A(n56080), .B(n56062), .Z(n56056) );
  XNOR U56044 ( .A(n56081), .B(n56082), .Z(n56062) );
  NOR U56045 ( .A(n56083), .B(n56084), .Z(n56082) );
  XOR U56046 ( .A(n56081), .B(n56085), .Z(n56083) );
  XNOR U56047 ( .A(n56061), .B(n56053), .Z(n56080) );
  XOR U56048 ( .A(n56086), .B(n56087), .Z(n56053) );
  AND U56049 ( .A(n56088), .B(n56089), .Z(n56087) );
  XOR U56050 ( .A(n56086), .B(n56090), .Z(n56088) );
  XNOR U56051 ( .A(n56091), .B(n56058), .Z(n56061) );
  XOR U56052 ( .A(n56092), .B(n56093), .Z(n56058) );
  AND U56053 ( .A(n56094), .B(n56095), .Z(n56093) );
  XNOR U56054 ( .A(n56096), .B(n56097), .Z(n56094) );
  IV U56055 ( .A(n56092), .Z(n56096) );
  XNOR U56056 ( .A(n56098), .B(n56099), .Z(n56091) );
  NOR U56057 ( .A(n56100), .B(n56101), .Z(n56099) );
  XNOR U56058 ( .A(n56098), .B(n56102), .Z(n56100) );
  XNOR U56059 ( .A(n56057), .B(n56064), .Z(n56079) );
  NOR U56060 ( .A(n56019), .B(n56103), .Z(n56064) );
  XOR U56061 ( .A(n56069), .B(n56068), .Z(n56057) );
  XNOR U56062 ( .A(n56104), .B(n56065), .Z(n56068) );
  XOR U56063 ( .A(n56105), .B(n56106), .Z(n56065) );
  AND U56064 ( .A(n56107), .B(n56108), .Z(n56106) );
  XNOR U56065 ( .A(n56109), .B(n56110), .Z(n56107) );
  IV U56066 ( .A(n56105), .Z(n56109) );
  XNOR U56067 ( .A(n56111), .B(n56112), .Z(n56104) );
  NOR U56068 ( .A(n56113), .B(n56114), .Z(n56112) );
  XNOR U56069 ( .A(n56111), .B(n56115), .Z(n56113) );
  XOR U56070 ( .A(n56116), .B(n56117), .Z(n56069) );
  NOR U56071 ( .A(n56118), .B(n56119), .Z(n56117) );
  XNOR U56072 ( .A(n56116), .B(n56120), .Z(n56118) );
  XNOR U56073 ( .A(n56010), .B(n56075), .Z(n56077) );
  XNOR U56074 ( .A(n56121), .B(n56122), .Z(n56010) );
  AND U56075 ( .A(n2336), .B(n56123), .Z(n56122) );
  XNOR U56076 ( .A(n56124), .B(n56125), .Z(n56123) );
  AND U56077 ( .A(n56016), .B(n56019), .Z(n56075) );
  XOR U56078 ( .A(n56126), .B(n56103), .Z(n56019) );
  XNOR U56079 ( .A(p_input[1904]), .B(p_input[2048]), .Z(n56103) );
  XNOR U56080 ( .A(n56090), .B(n56089), .Z(n56126) );
  XNOR U56081 ( .A(n56127), .B(n56097), .Z(n56089) );
  XNOR U56082 ( .A(n56085), .B(n56084), .Z(n56097) );
  XNOR U56083 ( .A(n56128), .B(n56081), .Z(n56084) );
  XNOR U56084 ( .A(p_input[1914]), .B(p_input[2058]), .Z(n56081) );
  XOR U56085 ( .A(p_input[1915]), .B(n29030), .Z(n56128) );
  XOR U56086 ( .A(p_input[1916]), .B(p_input[2060]), .Z(n56085) );
  XOR U56087 ( .A(n56095), .B(n56129), .Z(n56127) );
  IV U56088 ( .A(n56086), .Z(n56129) );
  XOR U56089 ( .A(p_input[1905]), .B(p_input[2049]), .Z(n56086) );
  XNOR U56090 ( .A(n56130), .B(n56102), .Z(n56095) );
  XNOR U56091 ( .A(p_input[1919]), .B(n29033), .Z(n56102) );
  XOR U56092 ( .A(n56092), .B(n56101), .Z(n56130) );
  XOR U56093 ( .A(n56131), .B(n56098), .Z(n56101) );
  XOR U56094 ( .A(p_input[1917]), .B(p_input[2061]), .Z(n56098) );
  XOR U56095 ( .A(p_input[1918]), .B(n29035), .Z(n56131) );
  XOR U56096 ( .A(p_input[1913]), .B(p_input[2057]), .Z(n56092) );
  XOR U56097 ( .A(n56110), .B(n56108), .Z(n56090) );
  XNOR U56098 ( .A(n56132), .B(n56115), .Z(n56108) );
  XOR U56099 ( .A(p_input[1912]), .B(p_input[2056]), .Z(n56115) );
  XOR U56100 ( .A(n56105), .B(n56114), .Z(n56132) );
  XOR U56101 ( .A(n56133), .B(n56111), .Z(n56114) );
  XOR U56102 ( .A(p_input[1910]), .B(p_input[2054]), .Z(n56111) );
  XOR U56103 ( .A(p_input[1911]), .B(n30404), .Z(n56133) );
  XOR U56104 ( .A(p_input[1906]), .B(p_input[2050]), .Z(n56105) );
  XNOR U56105 ( .A(n56120), .B(n56119), .Z(n56110) );
  XOR U56106 ( .A(n56134), .B(n56116), .Z(n56119) );
  XOR U56107 ( .A(p_input[1907]), .B(p_input[2051]), .Z(n56116) );
  XOR U56108 ( .A(p_input[1908]), .B(n30406), .Z(n56134) );
  XOR U56109 ( .A(p_input[1909]), .B(p_input[2053]), .Z(n56120) );
  XNOR U56110 ( .A(n56135), .B(n56136), .Z(n56016) );
  AND U56111 ( .A(n2336), .B(n56137), .Z(n56136) );
  XNOR U56112 ( .A(n56138), .B(n56139), .Z(n2336) );
  AND U56113 ( .A(n56140), .B(n56141), .Z(n56139) );
  XOR U56114 ( .A(n56030), .B(n56138), .Z(n56141) );
  XNOR U56115 ( .A(n56142), .B(n56138), .Z(n56140) );
  XOR U56116 ( .A(n56143), .B(n56144), .Z(n56138) );
  AND U56117 ( .A(n56145), .B(n56146), .Z(n56144) );
  XOR U56118 ( .A(n56045), .B(n56143), .Z(n56146) );
  XOR U56119 ( .A(n56143), .B(n56046), .Z(n56145) );
  XOR U56120 ( .A(n56147), .B(n56148), .Z(n56143) );
  AND U56121 ( .A(n56149), .B(n56150), .Z(n56148) );
  XOR U56122 ( .A(n56073), .B(n56147), .Z(n56150) );
  XOR U56123 ( .A(n56147), .B(n56074), .Z(n56149) );
  XOR U56124 ( .A(n56151), .B(n56152), .Z(n56147) );
  AND U56125 ( .A(n56153), .B(n56154), .Z(n56152) );
  XOR U56126 ( .A(n56151), .B(n56124), .Z(n56154) );
  XNOR U56127 ( .A(n56155), .B(n56156), .Z(n55976) );
  AND U56128 ( .A(n2340), .B(n56157), .Z(n56156) );
  XNOR U56129 ( .A(n56158), .B(n56159), .Z(n2340) );
  AND U56130 ( .A(n56160), .B(n56161), .Z(n56159) );
  XOR U56131 ( .A(n56158), .B(n55986), .Z(n56161) );
  XNOR U56132 ( .A(n56158), .B(n55946), .Z(n56160) );
  XOR U56133 ( .A(n56162), .B(n56163), .Z(n56158) );
  AND U56134 ( .A(n56164), .B(n56165), .Z(n56163) );
  XOR U56135 ( .A(n56162), .B(n55954), .Z(n56164) );
  XOR U56136 ( .A(n56166), .B(n56167), .Z(n55937) );
  AND U56137 ( .A(n2344), .B(n56157), .Z(n56167) );
  XNOR U56138 ( .A(n56155), .B(n56166), .Z(n56157) );
  XNOR U56139 ( .A(n56168), .B(n56169), .Z(n2344) );
  AND U56140 ( .A(n56170), .B(n56171), .Z(n56169) );
  XNOR U56141 ( .A(n56172), .B(n56168), .Z(n56171) );
  IV U56142 ( .A(n55986), .Z(n56172) );
  XOR U56143 ( .A(n56142), .B(n56173), .Z(n55986) );
  AND U56144 ( .A(n2347), .B(n56174), .Z(n56173) );
  XOR U56145 ( .A(n56029), .B(n56026), .Z(n56174) );
  XNOR U56146 ( .A(n55946), .B(n56168), .Z(n56170) );
  XNOR U56147 ( .A(n56175), .B(n56176), .Z(n55946) );
  AND U56148 ( .A(n2363), .B(n56177), .Z(n56176) );
  XNOR U56149 ( .A(n56178), .B(n56179), .Z(n56177) );
  XOR U56150 ( .A(n56162), .B(n56180), .Z(n56168) );
  AND U56151 ( .A(n56181), .B(n56165), .Z(n56180) );
  XNOR U56152 ( .A(n55996), .B(n56162), .Z(n56165) );
  XOR U56153 ( .A(n56046), .B(n56182), .Z(n55996) );
  AND U56154 ( .A(n2347), .B(n56183), .Z(n56182) );
  XOR U56155 ( .A(n56042), .B(n56046), .Z(n56183) );
  XNOR U56156 ( .A(n56184), .B(n56162), .Z(n56181) );
  IV U56157 ( .A(n55954), .Z(n56184) );
  XOR U56158 ( .A(n56185), .B(n56186), .Z(n55954) );
  AND U56159 ( .A(n2363), .B(n56187), .Z(n56186) );
  XOR U56160 ( .A(n56188), .B(n56189), .Z(n56162) );
  AND U56161 ( .A(n56190), .B(n56191), .Z(n56189) );
  XNOR U56162 ( .A(n56006), .B(n56188), .Z(n56191) );
  XOR U56163 ( .A(n56074), .B(n56192), .Z(n56006) );
  AND U56164 ( .A(n2347), .B(n56193), .Z(n56192) );
  XOR U56165 ( .A(n56070), .B(n56074), .Z(n56193) );
  XOR U56166 ( .A(n56188), .B(n55963), .Z(n56190) );
  XOR U56167 ( .A(n56194), .B(n56195), .Z(n55963) );
  AND U56168 ( .A(n2363), .B(n56196), .Z(n56195) );
  XOR U56169 ( .A(n56197), .B(n56198), .Z(n56188) );
  AND U56170 ( .A(n56199), .B(n56200), .Z(n56198) );
  XNOR U56171 ( .A(n56197), .B(n56014), .Z(n56200) );
  XOR U56172 ( .A(n56125), .B(n56201), .Z(n56014) );
  AND U56173 ( .A(n2347), .B(n56202), .Z(n56201) );
  XOR U56174 ( .A(n56121), .B(n56125), .Z(n56202) );
  XNOR U56175 ( .A(n56203), .B(n56197), .Z(n56199) );
  IV U56176 ( .A(n55973), .Z(n56203) );
  XOR U56177 ( .A(n56204), .B(n56205), .Z(n55973) );
  AND U56178 ( .A(n2363), .B(n56206), .Z(n56205) );
  AND U56179 ( .A(n56166), .B(n56155), .Z(n56197) );
  XNOR U56180 ( .A(n56207), .B(n56208), .Z(n56155) );
  AND U56181 ( .A(n2347), .B(n56137), .Z(n56208) );
  XNOR U56182 ( .A(n56135), .B(n56207), .Z(n56137) );
  XNOR U56183 ( .A(n56209), .B(n56210), .Z(n2347) );
  AND U56184 ( .A(n56211), .B(n56212), .Z(n56210) );
  XNOR U56185 ( .A(n56209), .B(n56026), .Z(n56212) );
  IV U56186 ( .A(n56030), .Z(n56026) );
  XOR U56187 ( .A(n56213), .B(n56214), .Z(n56030) );
  AND U56188 ( .A(n2351), .B(n56215), .Z(n56214) );
  XOR U56189 ( .A(n56216), .B(n56213), .Z(n56215) );
  XNOR U56190 ( .A(n56209), .B(n56142), .Z(n56211) );
  IV U56191 ( .A(n56029), .Z(n56142) );
  XOR U56192 ( .A(n56178), .B(n56217), .Z(n56029) );
  AND U56193 ( .A(n2359), .B(n56218), .Z(n56217) );
  XOR U56194 ( .A(n56178), .B(n56175), .Z(n56218) );
  XOR U56195 ( .A(n56219), .B(n56220), .Z(n56209) );
  AND U56196 ( .A(n56221), .B(n56222), .Z(n56220) );
  XNOR U56197 ( .A(n56219), .B(n56042), .Z(n56222) );
  IV U56198 ( .A(n56045), .Z(n56042) );
  XOR U56199 ( .A(n56223), .B(n56224), .Z(n56045) );
  AND U56200 ( .A(n2351), .B(n56225), .Z(n56224) );
  XOR U56201 ( .A(n56226), .B(n56223), .Z(n56225) );
  XOR U56202 ( .A(n56046), .B(n56219), .Z(n56221) );
  XOR U56203 ( .A(n56227), .B(n56228), .Z(n56046) );
  AND U56204 ( .A(n2359), .B(n56187), .Z(n56228) );
  XOR U56205 ( .A(n56227), .B(n56185), .Z(n56187) );
  XOR U56206 ( .A(n56229), .B(n56230), .Z(n56219) );
  AND U56207 ( .A(n56231), .B(n56232), .Z(n56230) );
  XNOR U56208 ( .A(n56229), .B(n56070), .Z(n56232) );
  IV U56209 ( .A(n56073), .Z(n56070) );
  XOR U56210 ( .A(n56233), .B(n56234), .Z(n56073) );
  AND U56211 ( .A(n2351), .B(n56235), .Z(n56234) );
  XNOR U56212 ( .A(n56236), .B(n56233), .Z(n56235) );
  XOR U56213 ( .A(n56074), .B(n56229), .Z(n56231) );
  XOR U56214 ( .A(n56237), .B(n56238), .Z(n56074) );
  AND U56215 ( .A(n2359), .B(n56196), .Z(n56238) );
  XOR U56216 ( .A(n56237), .B(n56194), .Z(n56196) );
  XOR U56217 ( .A(n56151), .B(n56239), .Z(n56229) );
  AND U56218 ( .A(n56153), .B(n56240), .Z(n56239) );
  XNOR U56219 ( .A(n56151), .B(n56121), .Z(n56240) );
  IV U56220 ( .A(n56124), .Z(n56121) );
  XOR U56221 ( .A(n56241), .B(n56242), .Z(n56124) );
  AND U56222 ( .A(n2351), .B(n56243), .Z(n56242) );
  XOR U56223 ( .A(n56244), .B(n56241), .Z(n56243) );
  XOR U56224 ( .A(n56125), .B(n56151), .Z(n56153) );
  XOR U56225 ( .A(n56245), .B(n56246), .Z(n56125) );
  AND U56226 ( .A(n2359), .B(n56206), .Z(n56246) );
  XOR U56227 ( .A(n56245), .B(n56204), .Z(n56206) );
  AND U56228 ( .A(n56207), .B(n56135), .Z(n56151) );
  XNOR U56229 ( .A(n56247), .B(n56248), .Z(n56135) );
  AND U56230 ( .A(n2351), .B(n56249), .Z(n56248) );
  XNOR U56231 ( .A(n56250), .B(n56247), .Z(n56249) );
  XNOR U56232 ( .A(n56251), .B(n56252), .Z(n2351) );
  AND U56233 ( .A(n56253), .B(n56254), .Z(n56252) );
  XOR U56234 ( .A(n56216), .B(n56251), .Z(n56254) );
  AND U56235 ( .A(n56255), .B(n56256), .Z(n56216) );
  XNOR U56236 ( .A(n56213), .B(n56251), .Z(n56253) );
  XNOR U56237 ( .A(n56257), .B(n56258), .Z(n56213) );
  AND U56238 ( .A(n56259), .B(n2355), .Z(n56258) );
  AND U56239 ( .A(n56257), .B(n56260), .Z(n56259) );
  XOR U56240 ( .A(n56261), .B(n56262), .Z(n56251) );
  AND U56241 ( .A(n56263), .B(n56264), .Z(n56262) );
  XNOR U56242 ( .A(n56261), .B(n56255), .Z(n56264) );
  IV U56243 ( .A(n56226), .Z(n56255) );
  XOR U56244 ( .A(n56265), .B(n56266), .Z(n56226) );
  XOR U56245 ( .A(n56267), .B(n56256), .Z(n56266) );
  AND U56246 ( .A(n56236), .B(n56268), .Z(n56256) );
  AND U56247 ( .A(n56269), .B(n56270), .Z(n56267) );
  XOR U56248 ( .A(n56271), .B(n56265), .Z(n56269) );
  XNOR U56249 ( .A(n56223), .B(n56261), .Z(n56263) );
  XNOR U56250 ( .A(n56272), .B(n56273), .Z(n56223) );
  AND U56251 ( .A(n2355), .B(n56274), .Z(n56273) );
  XNOR U56252 ( .A(n56275), .B(n56276), .Z(n56274) );
  XOR U56253 ( .A(n56277), .B(n56278), .Z(n56261) );
  AND U56254 ( .A(n56279), .B(n56280), .Z(n56278) );
  XNOR U56255 ( .A(n56277), .B(n56236), .Z(n56280) );
  XOR U56256 ( .A(n56281), .B(n56270), .Z(n56236) );
  XNOR U56257 ( .A(n56282), .B(n56265), .Z(n56270) );
  XOR U56258 ( .A(n56283), .B(n56284), .Z(n56265) );
  AND U56259 ( .A(n56285), .B(n56286), .Z(n56284) );
  XOR U56260 ( .A(n56287), .B(n56283), .Z(n56285) );
  XNOR U56261 ( .A(n56288), .B(n56289), .Z(n56282) );
  AND U56262 ( .A(n56290), .B(n56291), .Z(n56289) );
  XOR U56263 ( .A(n56288), .B(n56292), .Z(n56290) );
  XNOR U56264 ( .A(n56271), .B(n56268), .Z(n56281) );
  AND U56265 ( .A(n56293), .B(n56294), .Z(n56268) );
  XOR U56266 ( .A(n56295), .B(n56296), .Z(n56271) );
  AND U56267 ( .A(n56297), .B(n56298), .Z(n56296) );
  XOR U56268 ( .A(n56295), .B(n56299), .Z(n56297) );
  XNOR U56269 ( .A(n56233), .B(n56277), .Z(n56279) );
  XNOR U56270 ( .A(n56300), .B(n56301), .Z(n56233) );
  AND U56271 ( .A(n2355), .B(n56302), .Z(n56301) );
  XNOR U56272 ( .A(n56303), .B(n56304), .Z(n56302) );
  XOR U56273 ( .A(n56305), .B(n56306), .Z(n56277) );
  AND U56274 ( .A(n56307), .B(n56308), .Z(n56306) );
  XNOR U56275 ( .A(n56305), .B(n56293), .Z(n56308) );
  IV U56276 ( .A(n56244), .Z(n56293) );
  XNOR U56277 ( .A(n56309), .B(n56286), .Z(n56244) );
  XNOR U56278 ( .A(n56310), .B(n56292), .Z(n56286) );
  XNOR U56279 ( .A(n56311), .B(n56312), .Z(n56292) );
  NOR U56280 ( .A(n56313), .B(n56314), .Z(n56312) );
  XOR U56281 ( .A(n56311), .B(n56315), .Z(n56313) );
  XNOR U56282 ( .A(n56291), .B(n56283), .Z(n56310) );
  XOR U56283 ( .A(n56316), .B(n56317), .Z(n56283) );
  AND U56284 ( .A(n56318), .B(n56319), .Z(n56317) );
  XOR U56285 ( .A(n56316), .B(n56320), .Z(n56318) );
  XNOR U56286 ( .A(n56321), .B(n56288), .Z(n56291) );
  XOR U56287 ( .A(n56322), .B(n56323), .Z(n56288) );
  AND U56288 ( .A(n56324), .B(n56325), .Z(n56323) );
  XNOR U56289 ( .A(n56326), .B(n56327), .Z(n56324) );
  IV U56290 ( .A(n56322), .Z(n56326) );
  XNOR U56291 ( .A(n56328), .B(n56329), .Z(n56321) );
  NOR U56292 ( .A(n56330), .B(n56331), .Z(n56329) );
  XNOR U56293 ( .A(n56328), .B(n56332), .Z(n56330) );
  XNOR U56294 ( .A(n56287), .B(n56294), .Z(n56309) );
  NOR U56295 ( .A(n56250), .B(n56333), .Z(n56294) );
  XOR U56296 ( .A(n56299), .B(n56298), .Z(n56287) );
  XNOR U56297 ( .A(n56334), .B(n56295), .Z(n56298) );
  XOR U56298 ( .A(n56335), .B(n56336), .Z(n56295) );
  AND U56299 ( .A(n56337), .B(n56338), .Z(n56336) );
  XNOR U56300 ( .A(n56339), .B(n56340), .Z(n56337) );
  IV U56301 ( .A(n56335), .Z(n56339) );
  XNOR U56302 ( .A(n56341), .B(n56342), .Z(n56334) );
  NOR U56303 ( .A(n56343), .B(n56344), .Z(n56342) );
  XNOR U56304 ( .A(n56341), .B(n56345), .Z(n56343) );
  XOR U56305 ( .A(n56346), .B(n56347), .Z(n56299) );
  NOR U56306 ( .A(n56348), .B(n56349), .Z(n56347) );
  XNOR U56307 ( .A(n56346), .B(n56350), .Z(n56348) );
  XNOR U56308 ( .A(n56241), .B(n56305), .Z(n56307) );
  XNOR U56309 ( .A(n56351), .B(n56352), .Z(n56241) );
  AND U56310 ( .A(n2355), .B(n56353), .Z(n56352) );
  XNOR U56311 ( .A(n56354), .B(n56355), .Z(n56353) );
  AND U56312 ( .A(n56247), .B(n56250), .Z(n56305) );
  XOR U56313 ( .A(n56356), .B(n56333), .Z(n56250) );
  XNOR U56314 ( .A(p_input[1920]), .B(p_input[2048]), .Z(n56333) );
  XNOR U56315 ( .A(n56320), .B(n56319), .Z(n56356) );
  XNOR U56316 ( .A(n56357), .B(n56327), .Z(n56319) );
  XNOR U56317 ( .A(n56315), .B(n56314), .Z(n56327) );
  XNOR U56318 ( .A(n56358), .B(n56311), .Z(n56314) );
  XNOR U56319 ( .A(p_input[1930]), .B(p_input[2058]), .Z(n56311) );
  XOR U56320 ( .A(p_input[1931]), .B(n29030), .Z(n56358) );
  XOR U56321 ( .A(p_input[1932]), .B(p_input[2060]), .Z(n56315) );
  XOR U56322 ( .A(n56325), .B(n56359), .Z(n56357) );
  IV U56323 ( .A(n56316), .Z(n56359) );
  XOR U56324 ( .A(p_input[1921]), .B(p_input[2049]), .Z(n56316) );
  XNOR U56325 ( .A(n56360), .B(n56332), .Z(n56325) );
  XNOR U56326 ( .A(p_input[1935]), .B(n29033), .Z(n56332) );
  XOR U56327 ( .A(n56322), .B(n56331), .Z(n56360) );
  XOR U56328 ( .A(n56361), .B(n56328), .Z(n56331) );
  XOR U56329 ( .A(p_input[1933]), .B(p_input[2061]), .Z(n56328) );
  XOR U56330 ( .A(p_input[1934]), .B(n29035), .Z(n56361) );
  XOR U56331 ( .A(p_input[1929]), .B(p_input[2057]), .Z(n56322) );
  XOR U56332 ( .A(n56340), .B(n56338), .Z(n56320) );
  XNOR U56333 ( .A(n56362), .B(n56345), .Z(n56338) );
  XOR U56334 ( .A(p_input[1928]), .B(p_input[2056]), .Z(n56345) );
  XOR U56335 ( .A(n56335), .B(n56344), .Z(n56362) );
  XOR U56336 ( .A(n56363), .B(n56341), .Z(n56344) );
  XOR U56337 ( .A(p_input[1926]), .B(p_input[2054]), .Z(n56341) );
  XOR U56338 ( .A(p_input[1927]), .B(n30404), .Z(n56363) );
  XOR U56339 ( .A(p_input[1922]), .B(p_input[2050]), .Z(n56335) );
  XNOR U56340 ( .A(n56350), .B(n56349), .Z(n56340) );
  XOR U56341 ( .A(n56364), .B(n56346), .Z(n56349) );
  XOR U56342 ( .A(p_input[1923]), .B(p_input[2051]), .Z(n56346) );
  XOR U56343 ( .A(p_input[1924]), .B(n30406), .Z(n56364) );
  XOR U56344 ( .A(p_input[1925]), .B(p_input[2053]), .Z(n56350) );
  XNOR U56345 ( .A(n56365), .B(n56366), .Z(n56247) );
  AND U56346 ( .A(n2355), .B(n56367), .Z(n56366) );
  XNOR U56347 ( .A(n56368), .B(n56369), .Z(n2355) );
  AND U56348 ( .A(n56370), .B(n56371), .Z(n56369) );
  XNOR U56349 ( .A(n56257), .B(n56368), .Z(n56371) );
  XNOR U56350 ( .A(n56260), .B(n56368), .Z(n56370) );
  XOR U56351 ( .A(n56372), .B(n56373), .Z(n56368) );
  AND U56352 ( .A(n56374), .B(n56375), .Z(n56373) );
  XOR U56353 ( .A(n56275), .B(n56372), .Z(n56375) );
  XOR U56354 ( .A(n56372), .B(n56276), .Z(n56374) );
  XOR U56355 ( .A(n56376), .B(n56377), .Z(n56372) );
  AND U56356 ( .A(n56378), .B(n56379), .Z(n56377) );
  XOR U56357 ( .A(n56303), .B(n56376), .Z(n56379) );
  XOR U56358 ( .A(n56376), .B(n56304), .Z(n56378) );
  XOR U56359 ( .A(n56380), .B(n56381), .Z(n56376) );
  AND U56360 ( .A(n56382), .B(n56383), .Z(n56381) );
  XOR U56361 ( .A(n56380), .B(n56354), .Z(n56383) );
  XNOR U56362 ( .A(n56384), .B(n56385), .Z(n56207) );
  AND U56363 ( .A(n2359), .B(n56386), .Z(n56385) );
  XNOR U56364 ( .A(n56387), .B(n56388), .Z(n2359) );
  AND U56365 ( .A(n56389), .B(n56390), .Z(n56388) );
  XNOR U56366 ( .A(n56387), .B(n56178), .Z(n56390) );
  XOR U56367 ( .A(n56387), .B(n56175), .Z(n56389) );
  XOR U56368 ( .A(n56391), .B(n56392), .Z(n56387) );
  AND U56369 ( .A(n56393), .B(n56394), .Z(n56392) );
  XOR U56370 ( .A(n56391), .B(n56185), .Z(n56393) );
  XOR U56371 ( .A(n56395), .B(n56396), .Z(n56166) );
  AND U56372 ( .A(n2363), .B(n56386), .Z(n56396) );
  XNOR U56373 ( .A(n56384), .B(n56395), .Z(n56386) );
  XNOR U56374 ( .A(n56397), .B(n56398), .Z(n2363) );
  AND U56375 ( .A(n56399), .B(n56400), .Z(n56398) );
  XNOR U56376 ( .A(n56178), .B(n56397), .Z(n56400) );
  XNOR U56377 ( .A(n56260), .B(n56401), .Z(n56178) );
  AND U56378 ( .A(n56402), .B(n2366), .Z(n56401) );
  NOR U56379 ( .A(n56403), .B(n56404), .Z(n56402) );
  XOR U56380 ( .A(n56397), .B(n56175), .Z(n56399) );
  IV U56381 ( .A(n56179), .Z(n56175) );
  AND U56382 ( .A(n56405), .B(n56406), .Z(n56179) );
  XOR U56383 ( .A(n56391), .B(n56407), .Z(n56397) );
  AND U56384 ( .A(n56408), .B(n56394), .Z(n56407) );
  XNOR U56385 ( .A(n56227), .B(n56391), .Z(n56394) );
  XOR U56386 ( .A(n56276), .B(n56409), .Z(n56227) );
  AND U56387 ( .A(n2366), .B(n56410), .Z(n56409) );
  XOR U56388 ( .A(n56272), .B(n56276), .Z(n56410) );
  XNOR U56389 ( .A(n56411), .B(n56391), .Z(n56408) );
  IV U56390 ( .A(n56185), .Z(n56411) );
  XOR U56391 ( .A(n56412), .B(n56413), .Z(n56185) );
  AND U56392 ( .A(n2382), .B(n56414), .Z(n56413) );
  XOR U56393 ( .A(n56415), .B(n56416), .Z(n56391) );
  AND U56394 ( .A(n56417), .B(n56418), .Z(n56416) );
  XNOR U56395 ( .A(n56237), .B(n56415), .Z(n56418) );
  XOR U56396 ( .A(n56304), .B(n56419), .Z(n56237) );
  AND U56397 ( .A(n2366), .B(n56420), .Z(n56419) );
  XOR U56398 ( .A(n56300), .B(n56304), .Z(n56420) );
  XOR U56399 ( .A(n56415), .B(n56194), .Z(n56417) );
  XOR U56400 ( .A(n56421), .B(n56422), .Z(n56194) );
  AND U56401 ( .A(n2382), .B(n56423), .Z(n56422) );
  XOR U56402 ( .A(n56424), .B(n56425), .Z(n56415) );
  AND U56403 ( .A(n56426), .B(n56427), .Z(n56425) );
  XNOR U56404 ( .A(n56424), .B(n56245), .Z(n56427) );
  XOR U56405 ( .A(n56355), .B(n56428), .Z(n56245) );
  AND U56406 ( .A(n2366), .B(n56429), .Z(n56428) );
  XOR U56407 ( .A(n56351), .B(n56355), .Z(n56429) );
  XNOR U56408 ( .A(n56430), .B(n56424), .Z(n56426) );
  IV U56409 ( .A(n56204), .Z(n56430) );
  XOR U56410 ( .A(n56431), .B(n56432), .Z(n56204) );
  AND U56411 ( .A(n2382), .B(n56433), .Z(n56432) );
  AND U56412 ( .A(n56395), .B(n56384), .Z(n56424) );
  XNOR U56413 ( .A(n56434), .B(n56435), .Z(n56384) );
  AND U56414 ( .A(n2366), .B(n56367), .Z(n56435) );
  XNOR U56415 ( .A(n56365), .B(n56434), .Z(n56367) );
  XNOR U56416 ( .A(n56436), .B(n56437), .Z(n2366) );
  AND U56417 ( .A(n56438), .B(n56439), .Z(n56437) );
  XNOR U56418 ( .A(n56257), .B(n56436), .Z(n56439) );
  IV U56419 ( .A(n56403), .Z(n56257) );
  AND U56420 ( .A(n56440), .B(n56441), .Z(n56403) );
  IV U56421 ( .A(n56442), .Z(n56440) );
  XNOR U56422 ( .A(n56260), .B(n56436), .Z(n56438) );
  IV U56423 ( .A(n56404), .Z(n56260) );
  NOR U56424 ( .A(n56405), .B(n56406), .Z(n56404) );
  XOR U56425 ( .A(n56443), .B(n56444), .Z(n56436) );
  AND U56426 ( .A(n56445), .B(n56446), .Z(n56444) );
  XNOR U56427 ( .A(n56443), .B(n56272), .Z(n56446) );
  IV U56428 ( .A(n56275), .Z(n56272) );
  XOR U56429 ( .A(n56447), .B(n56448), .Z(n56275) );
  AND U56430 ( .A(n2370), .B(n56449), .Z(n56448) );
  XOR U56431 ( .A(n56450), .B(n56447), .Z(n56449) );
  XOR U56432 ( .A(n56276), .B(n56443), .Z(n56445) );
  XOR U56433 ( .A(n56451), .B(n56452), .Z(n56276) );
  AND U56434 ( .A(n2378), .B(n56414), .Z(n56452) );
  XOR U56435 ( .A(n56451), .B(n56412), .Z(n56414) );
  XOR U56436 ( .A(n56453), .B(n56454), .Z(n56443) );
  AND U56437 ( .A(n56455), .B(n56456), .Z(n56454) );
  XNOR U56438 ( .A(n56453), .B(n56300), .Z(n56456) );
  IV U56439 ( .A(n56303), .Z(n56300) );
  XOR U56440 ( .A(n56457), .B(n56458), .Z(n56303) );
  AND U56441 ( .A(n2370), .B(n56459), .Z(n56458) );
  XNOR U56442 ( .A(n56460), .B(n56457), .Z(n56459) );
  XOR U56443 ( .A(n56304), .B(n56453), .Z(n56455) );
  XOR U56444 ( .A(n56461), .B(n56462), .Z(n56304) );
  AND U56445 ( .A(n2378), .B(n56423), .Z(n56462) );
  XOR U56446 ( .A(n56461), .B(n56421), .Z(n56423) );
  XOR U56447 ( .A(n56380), .B(n56463), .Z(n56453) );
  AND U56448 ( .A(n56382), .B(n56464), .Z(n56463) );
  XNOR U56449 ( .A(n56380), .B(n56351), .Z(n56464) );
  IV U56450 ( .A(n56354), .Z(n56351) );
  XOR U56451 ( .A(n56465), .B(n56466), .Z(n56354) );
  AND U56452 ( .A(n2370), .B(n56467), .Z(n56466) );
  XOR U56453 ( .A(n56468), .B(n56465), .Z(n56467) );
  XOR U56454 ( .A(n56355), .B(n56380), .Z(n56382) );
  XOR U56455 ( .A(n56469), .B(n56470), .Z(n56355) );
  AND U56456 ( .A(n2378), .B(n56433), .Z(n56470) );
  XOR U56457 ( .A(n56469), .B(n56431), .Z(n56433) );
  AND U56458 ( .A(n56434), .B(n56365), .Z(n56380) );
  XNOR U56459 ( .A(n56471), .B(n56472), .Z(n56365) );
  AND U56460 ( .A(n2370), .B(n56473), .Z(n56472) );
  XNOR U56461 ( .A(n56474), .B(n56471), .Z(n56473) );
  XNOR U56462 ( .A(n56475), .B(n56476), .Z(n2370) );
  NOR U56463 ( .A(n56477), .B(n56478), .Z(n56476) );
  XNOR U56464 ( .A(n56475), .B(n56442), .Z(n56478) );
  NOR U56465 ( .A(n56479), .B(n56480), .Z(n56442) );
  NOR U56466 ( .A(n56475), .B(n56441), .Z(n56477) );
  AND U56467 ( .A(n56481), .B(n56482), .Z(n56441) );
  XOR U56468 ( .A(n56483), .B(n56484), .Z(n56475) );
  AND U56469 ( .A(n56485), .B(n56486), .Z(n56484) );
  XNOR U56470 ( .A(n56483), .B(n56481), .Z(n56486) );
  IV U56471 ( .A(n56450), .Z(n56481) );
  XOR U56472 ( .A(n56487), .B(n56488), .Z(n56450) );
  XOR U56473 ( .A(n56489), .B(n56482), .Z(n56488) );
  AND U56474 ( .A(n56460), .B(n56490), .Z(n56482) );
  AND U56475 ( .A(n56491), .B(n56492), .Z(n56489) );
  XOR U56476 ( .A(n56493), .B(n56487), .Z(n56491) );
  XNOR U56477 ( .A(n56447), .B(n56483), .Z(n56485) );
  XNOR U56478 ( .A(n56494), .B(n56495), .Z(n56447) );
  AND U56479 ( .A(n2374), .B(n56496), .Z(n56495) );
  XNOR U56480 ( .A(n56497), .B(n56498), .Z(n56496) );
  XOR U56481 ( .A(n56499), .B(n56500), .Z(n56483) );
  AND U56482 ( .A(n56501), .B(n56502), .Z(n56500) );
  XNOR U56483 ( .A(n56499), .B(n56460), .Z(n56502) );
  XOR U56484 ( .A(n56503), .B(n56492), .Z(n56460) );
  XNOR U56485 ( .A(n56504), .B(n56487), .Z(n56492) );
  XOR U56486 ( .A(n56505), .B(n56506), .Z(n56487) );
  AND U56487 ( .A(n56507), .B(n56508), .Z(n56506) );
  XOR U56488 ( .A(n56509), .B(n56505), .Z(n56507) );
  XNOR U56489 ( .A(n56510), .B(n56511), .Z(n56504) );
  AND U56490 ( .A(n56512), .B(n56513), .Z(n56511) );
  XOR U56491 ( .A(n56510), .B(n56514), .Z(n56512) );
  XNOR U56492 ( .A(n56493), .B(n56490), .Z(n56503) );
  AND U56493 ( .A(n56515), .B(n56516), .Z(n56490) );
  XOR U56494 ( .A(n56517), .B(n56518), .Z(n56493) );
  AND U56495 ( .A(n56519), .B(n56520), .Z(n56518) );
  XOR U56496 ( .A(n56517), .B(n56521), .Z(n56519) );
  XNOR U56497 ( .A(n56457), .B(n56499), .Z(n56501) );
  XNOR U56498 ( .A(n56522), .B(n56523), .Z(n56457) );
  AND U56499 ( .A(n2374), .B(n56524), .Z(n56523) );
  XNOR U56500 ( .A(n56525), .B(n56526), .Z(n56524) );
  XOR U56501 ( .A(n56527), .B(n56528), .Z(n56499) );
  AND U56502 ( .A(n56529), .B(n56530), .Z(n56528) );
  XNOR U56503 ( .A(n56527), .B(n56515), .Z(n56530) );
  IV U56504 ( .A(n56468), .Z(n56515) );
  XNOR U56505 ( .A(n56531), .B(n56508), .Z(n56468) );
  XNOR U56506 ( .A(n56532), .B(n56514), .Z(n56508) );
  XNOR U56507 ( .A(n56533), .B(n56534), .Z(n56514) );
  NOR U56508 ( .A(n56535), .B(n56536), .Z(n56534) );
  XOR U56509 ( .A(n56533), .B(n56537), .Z(n56535) );
  XNOR U56510 ( .A(n56513), .B(n56505), .Z(n56532) );
  XOR U56511 ( .A(n56538), .B(n56539), .Z(n56505) );
  AND U56512 ( .A(n56540), .B(n56541), .Z(n56539) );
  XOR U56513 ( .A(n56538), .B(n56542), .Z(n56540) );
  XNOR U56514 ( .A(n56543), .B(n56510), .Z(n56513) );
  XOR U56515 ( .A(n56544), .B(n56545), .Z(n56510) );
  AND U56516 ( .A(n56546), .B(n56547), .Z(n56545) );
  XNOR U56517 ( .A(n56548), .B(n56549), .Z(n56546) );
  IV U56518 ( .A(n56544), .Z(n56548) );
  XNOR U56519 ( .A(n56550), .B(n56551), .Z(n56543) );
  NOR U56520 ( .A(n56552), .B(n56553), .Z(n56551) );
  XNOR U56521 ( .A(n56550), .B(n56554), .Z(n56552) );
  XNOR U56522 ( .A(n56509), .B(n56516), .Z(n56531) );
  NOR U56523 ( .A(n56474), .B(n56555), .Z(n56516) );
  XOR U56524 ( .A(n56521), .B(n56520), .Z(n56509) );
  XNOR U56525 ( .A(n56556), .B(n56517), .Z(n56520) );
  XOR U56526 ( .A(n56557), .B(n56558), .Z(n56517) );
  AND U56527 ( .A(n56559), .B(n56560), .Z(n56558) );
  XNOR U56528 ( .A(n56561), .B(n56562), .Z(n56559) );
  IV U56529 ( .A(n56557), .Z(n56561) );
  XNOR U56530 ( .A(n56563), .B(n56564), .Z(n56556) );
  NOR U56531 ( .A(n56565), .B(n56566), .Z(n56564) );
  XNOR U56532 ( .A(n56563), .B(n56567), .Z(n56565) );
  XOR U56533 ( .A(n56568), .B(n56569), .Z(n56521) );
  NOR U56534 ( .A(n56570), .B(n56571), .Z(n56569) );
  XNOR U56535 ( .A(n56568), .B(n56572), .Z(n56570) );
  XNOR U56536 ( .A(n56465), .B(n56527), .Z(n56529) );
  XNOR U56537 ( .A(n56573), .B(n56574), .Z(n56465) );
  AND U56538 ( .A(n2374), .B(n56575), .Z(n56574) );
  XNOR U56539 ( .A(n56576), .B(n56577), .Z(n56575) );
  AND U56540 ( .A(n56471), .B(n56474), .Z(n56527) );
  XOR U56541 ( .A(n56578), .B(n56555), .Z(n56474) );
  XNOR U56542 ( .A(p_input[1936]), .B(p_input[2048]), .Z(n56555) );
  XNOR U56543 ( .A(n56542), .B(n56541), .Z(n56578) );
  XNOR U56544 ( .A(n56579), .B(n56549), .Z(n56541) );
  XNOR U56545 ( .A(n56537), .B(n56536), .Z(n56549) );
  XNOR U56546 ( .A(n56580), .B(n56533), .Z(n56536) );
  XNOR U56547 ( .A(p_input[1946]), .B(p_input[2058]), .Z(n56533) );
  XOR U56548 ( .A(p_input[1947]), .B(n29030), .Z(n56580) );
  XOR U56549 ( .A(p_input[1948]), .B(p_input[2060]), .Z(n56537) );
  XOR U56550 ( .A(n56547), .B(n56581), .Z(n56579) );
  IV U56551 ( .A(n56538), .Z(n56581) );
  XOR U56552 ( .A(p_input[1937]), .B(p_input[2049]), .Z(n56538) );
  XNOR U56553 ( .A(n56582), .B(n56554), .Z(n56547) );
  XNOR U56554 ( .A(p_input[1951]), .B(n29033), .Z(n56554) );
  XOR U56555 ( .A(n56544), .B(n56553), .Z(n56582) );
  XOR U56556 ( .A(n56583), .B(n56550), .Z(n56553) );
  XOR U56557 ( .A(p_input[1949]), .B(p_input[2061]), .Z(n56550) );
  XOR U56558 ( .A(p_input[1950]), .B(n29035), .Z(n56583) );
  XOR U56559 ( .A(p_input[1945]), .B(p_input[2057]), .Z(n56544) );
  XOR U56560 ( .A(n56562), .B(n56560), .Z(n56542) );
  XNOR U56561 ( .A(n56584), .B(n56567), .Z(n56560) );
  XOR U56562 ( .A(p_input[1944]), .B(p_input[2056]), .Z(n56567) );
  XOR U56563 ( .A(n56557), .B(n56566), .Z(n56584) );
  XOR U56564 ( .A(n56585), .B(n56563), .Z(n56566) );
  XOR U56565 ( .A(p_input[1942]), .B(p_input[2054]), .Z(n56563) );
  XOR U56566 ( .A(p_input[1943]), .B(n30404), .Z(n56585) );
  XOR U56567 ( .A(p_input[1938]), .B(p_input[2050]), .Z(n56557) );
  XNOR U56568 ( .A(n56572), .B(n56571), .Z(n56562) );
  XOR U56569 ( .A(n56586), .B(n56568), .Z(n56571) );
  XOR U56570 ( .A(p_input[1939]), .B(p_input[2051]), .Z(n56568) );
  XOR U56571 ( .A(p_input[1940]), .B(n30406), .Z(n56586) );
  XOR U56572 ( .A(p_input[1941]), .B(p_input[2053]), .Z(n56572) );
  XNOR U56573 ( .A(n56587), .B(n56588), .Z(n56471) );
  AND U56574 ( .A(n2374), .B(n56589), .Z(n56588) );
  XNOR U56575 ( .A(n56590), .B(n56591), .Z(n2374) );
  NOR U56576 ( .A(n56592), .B(n56593), .Z(n56591) );
  XNOR U56577 ( .A(n56590), .B(n56594), .Z(n56593) );
  NOR U56578 ( .A(n56590), .B(n56480), .Z(n56592) );
  XOR U56579 ( .A(n56595), .B(n56596), .Z(n56590) );
  AND U56580 ( .A(n56597), .B(n56598), .Z(n56596) );
  XOR U56581 ( .A(n56497), .B(n56595), .Z(n56598) );
  XOR U56582 ( .A(n56595), .B(n56498), .Z(n56597) );
  XOR U56583 ( .A(n56599), .B(n56600), .Z(n56595) );
  AND U56584 ( .A(n56601), .B(n56602), .Z(n56600) );
  XOR U56585 ( .A(n56525), .B(n56599), .Z(n56602) );
  XOR U56586 ( .A(n56599), .B(n56526), .Z(n56601) );
  XOR U56587 ( .A(n56603), .B(n56604), .Z(n56599) );
  AND U56588 ( .A(n56605), .B(n56606), .Z(n56604) );
  XOR U56589 ( .A(n56603), .B(n56576), .Z(n56606) );
  XNOR U56590 ( .A(n56607), .B(n56608), .Z(n56434) );
  AND U56591 ( .A(n2378), .B(n56609), .Z(n56608) );
  XNOR U56592 ( .A(n56610), .B(n56611), .Z(n2378) );
  NOR U56593 ( .A(n56612), .B(n56613), .Z(n56611) );
  XOR U56594 ( .A(n56406), .B(n56610), .Z(n56613) );
  NOR U56595 ( .A(n56610), .B(n56405), .Z(n56612) );
  XOR U56596 ( .A(n56614), .B(n56615), .Z(n56610) );
  AND U56597 ( .A(n56616), .B(n56617), .Z(n56615) );
  XOR U56598 ( .A(n56614), .B(n56412), .Z(n56616) );
  XOR U56599 ( .A(n56618), .B(n56619), .Z(n56395) );
  AND U56600 ( .A(n2382), .B(n56609), .Z(n56619) );
  XNOR U56601 ( .A(n56607), .B(n56618), .Z(n56609) );
  XNOR U56602 ( .A(n56620), .B(n56621), .Z(n2382) );
  NOR U56603 ( .A(n56622), .B(n56623), .Z(n56621) );
  XNOR U56604 ( .A(n56406), .B(n56624), .Z(n56623) );
  IV U56605 ( .A(n56620), .Z(n56624) );
  AND U56606 ( .A(n56625), .B(n56626), .Z(n56406) );
  NOR U56607 ( .A(n56620), .B(n56405), .Z(n56622) );
  AND U56608 ( .A(n56480), .B(n56479), .Z(n56405) );
  IV U56609 ( .A(n56594), .Z(n56479) );
  XOR U56610 ( .A(n56614), .B(n56627), .Z(n56620) );
  AND U56611 ( .A(n56628), .B(n56617), .Z(n56627) );
  XNOR U56612 ( .A(n56451), .B(n56614), .Z(n56617) );
  XOR U56613 ( .A(n56498), .B(n56629), .Z(n56451) );
  AND U56614 ( .A(n2385), .B(n56630), .Z(n56629) );
  XOR U56615 ( .A(n56494), .B(n56498), .Z(n56630) );
  XNOR U56616 ( .A(n56631), .B(n56614), .Z(n56628) );
  IV U56617 ( .A(n56412), .Z(n56631) );
  XOR U56618 ( .A(n56632), .B(n56633), .Z(n56412) );
  AND U56619 ( .A(n2401), .B(n56634), .Z(n56633) );
  XOR U56620 ( .A(n56635), .B(n56636), .Z(n56614) );
  AND U56621 ( .A(n56637), .B(n56638), .Z(n56636) );
  XNOR U56622 ( .A(n56461), .B(n56635), .Z(n56638) );
  XOR U56623 ( .A(n56526), .B(n56639), .Z(n56461) );
  AND U56624 ( .A(n2385), .B(n56640), .Z(n56639) );
  XOR U56625 ( .A(n56522), .B(n56526), .Z(n56640) );
  XOR U56626 ( .A(n56635), .B(n56421), .Z(n56637) );
  XOR U56627 ( .A(n56641), .B(n56642), .Z(n56421) );
  AND U56628 ( .A(n2401), .B(n56643), .Z(n56642) );
  XOR U56629 ( .A(n56644), .B(n56645), .Z(n56635) );
  AND U56630 ( .A(n56646), .B(n56647), .Z(n56645) );
  XNOR U56631 ( .A(n56644), .B(n56469), .Z(n56647) );
  XOR U56632 ( .A(n56577), .B(n56648), .Z(n56469) );
  AND U56633 ( .A(n2385), .B(n56649), .Z(n56648) );
  XOR U56634 ( .A(n56573), .B(n56577), .Z(n56649) );
  XNOR U56635 ( .A(n56650), .B(n56644), .Z(n56646) );
  IV U56636 ( .A(n56431), .Z(n56650) );
  XOR U56637 ( .A(n56651), .B(n56652), .Z(n56431) );
  AND U56638 ( .A(n2401), .B(n56653), .Z(n56652) );
  AND U56639 ( .A(n56618), .B(n56607), .Z(n56644) );
  XNOR U56640 ( .A(n56654), .B(n56655), .Z(n56607) );
  AND U56641 ( .A(n2385), .B(n56589), .Z(n56655) );
  XNOR U56642 ( .A(n56587), .B(n56654), .Z(n56589) );
  XNOR U56643 ( .A(n56656), .B(n56657), .Z(n2385) );
  NOR U56644 ( .A(n56658), .B(n56659), .Z(n56657) );
  XNOR U56645 ( .A(n56656), .B(n56594), .Z(n56659) );
  NOR U56646 ( .A(n56625), .B(n56626), .Z(n56594) );
  NOR U56647 ( .A(n56656), .B(n56480), .Z(n56658) );
  AND U56648 ( .A(n56660), .B(n56661), .Z(n56480) );
  IV U56649 ( .A(n56662), .Z(n56660) );
  XOR U56650 ( .A(n56663), .B(n56664), .Z(n56656) );
  AND U56651 ( .A(n56665), .B(n56666), .Z(n56664) );
  XNOR U56652 ( .A(n56663), .B(n56494), .Z(n56666) );
  IV U56653 ( .A(n56497), .Z(n56494) );
  XOR U56654 ( .A(n56667), .B(n56668), .Z(n56497) );
  AND U56655 ( .A(n2389), .B(n56669), .Z(n56668) );
  XOR U56656 ( .A(n56670), .B(n56667), .Z(n56669) );
  XOR U56657 ( .A(n56498), .B(n56663), .Z(n56665) );
  XOR U56658 ( .A(n56671), .B(n56672), .Z(n56498) );
  AND U56659 ( .A(n2397), .B(n56634), .Z(n56672) );
  XOR U56660 ( .A(n56671), .B(n56632), .Z(n56634) );
  XOR U56661 ( .A(n56673), .B(n56674), .Z(n56663) );
  AND U56662 ( .A(n56675), .B(n56676), .Z(n56674) );
  XNOR U56663 ( .A(n56673), .B(n56522), .Z(n56676) );
  IV U56664 ( .A(n56525), .Z(n56522) );
  XOR U56665 ( .A(n56677), .B(n56678), .Z(n56525) );
  AND U56666 ( .A(n2389), .B(n56679), .Z(n56678) );
  XNOR U56667 ( .A(n56680), .B(n56677), .Z(n56679) );
  XOR U56668 ( .A(n56526), .B(n56673), .Z(n56675) );
  XOR U56669 ( .A(n56681), .B(n56682), .Z(n56526) );
  AND U56670 ( .A(n2397), .B(n56643), .Z(n56682) );
  XOR U56671 ( .A(n56681), .B(n56641), .Z(n56643) );
  XOR U56672 ( .A(n56603), .B(n56683), .Z(n56673) );
  AND U56673 ( .A(n56605), .B(n56684), .Z(n56683) );
  XNOR U56674 ( .A(n56603), .B(n56573), .Z(n56684) );
  IV U56675 ( .A(n56576), .Z(n56573) );
  XOR U56676 ( .A(n56685), .B(n56686), .Z(n56576) );
  AND U56677 ( .A(n2389), .B(n56687), .Z(n56686) );
  XOR U56678 ( .A(n56688), .B(n56685), .Z(n56687) );
  XOR U56679 ( .A(n56577), .B(n56603), .Z(n56605) );
  XOR U56680 ( .A(n56689), .B(n56690), .Z(n56577) );
  AND U56681 ( .A(n2397), .B(n56653), .Z(n56690) );
  XOR U56682 ( .A(n56689), .B(n56651), .Z(n56653) );
  AND U56683 ( .A(n56654), .B(n56587), .Z(n56603) );
  XNOR U56684 ( .A(n56691), .B(n56692), .Z(n56587) );
  AND U56685 ( .A(n2389), .B(n56693), .Z(n56692) );
  XNOR U56686 ( .A(n56694), .B(n56691), .Z(n56693) );
  XNOR U56687 ( .A(n56695), .B(n56696), .Z(n2389) );
  NOR U56688 ( .A(n56697), .B(n56698), .Z(n56696) );
  XNOR U56689 ( .A(n56695), .B(n56662), .Z(n56698) );
  NOR U56690 ( .A(n56699), .B(n56700), .Z(n56662) );
  NOR U56691 ( .A(n56695), .B(n56661), .Z(n56697) );
  AND U56692 ( .A(n56701), .B(n56702), .Z(n56661) );
  XOR U56693 ( .A(n56703), .B(n56704), .Z(n56695) );
  AND U56694 ( .A(n56705), .B(n56706), .Z(n56704) );
  XNOR U56695 ( .A(n56703), .B(n56701), .Z(n56706) );
  IV U56696 ( .A(n56670), .Z(n56701) );
  XOR U56697 ( .A(n56707), .B(n56708), .Z(n56670) );
  XOR U56698 ( .A(n56709), .B(n56702), .Z(n56708) );
  AND U56699 ( .A(n56680), .B(n56710), .Z(n56702) );
  AND U56700 ( .A(n56711), .B(n56712), .Z(n56709) );
  XOR U56701 ( .A(n56713), .B(n56707), .Z(n56711) );
  XNOR U56702 ( .A(n56667), .B(n56703), .Z(n56705) );
  XNOR U56703 ( .A(n56714), .B(n56715), .Z(n56667) );
  AND U56704 ( .A(n2393), .B(n56716), .Z(n56715) );
  XNOR U56705 ( .A(n56717), .B(n56718), .Z(n56716) );
  XOR U56706 ( .A(n56719), .B(n56720), .Z(n56703) );
  AND U56707 ( .A(n56721), .B(n56722), .Z(n56720) );
  XNOR U56708 ( .A(n56719), .B(n56680), .Z(n56722) );
  XOR U56709 ( .A(n56723), .B(n56712), .Z(n56680) );
  XNOR U56710 ( .A(n56724), .B(n56707), .Z(n56712) );
  XOR U56711 ( .A(n56725), .B(n56726), .Z(n56707) );
  AND U56712 ( .A(n56727), .B(n56728), .Z(n56726) );
  XOR U56713 ( .A(n56729), .B(n56725), .Z(n56727) );
  XNOR U56714 ( .A(n56730), .B(n56731), .Z(n56724) );
  AND U56715 ( .A(n56732), .B(n56733), .Z(n56731) );
  XOR U56716 ( .A(n56730), .B(n56734), .Z(n56732) );
  XNOR U56717 ( .A(n56713), .B(n56710), .Z(n56723) );
  AND U56718 ( .A(n56735), .B(n56736), .Z(n56710) );
  XOR U56719 ( .A(n56737), .B(n56738), .Z(n56713) );
  AND U56720 ( .A(n56739), .B(n56740), .Z(n56738) );
  XOR U56721 ( .A(n56737), .B(n56741), .Z(n56739) );
  XNOR U56722 ( .A(n56677), .B(n56719), .Z(n56721) );
  XNOR U56723 ( .A(n56742), .B(n56743), .Z(n56677) );
  AND U56724 ( .A(n2393), .B(n56744), .Z(n56743) );
  XNOR U56725 ( .A(n56745), .B(n56746), .Z(n56744) );
  XOR U56726 ( .A(n56747), .B(n56748), .Z(n56719) );
  AND U56727 ( .A(n56749), .B(n56750), .Z(n56748) );
  XNOR U56728 ( .A(n56747), .B(n56735), .Z(n56750) );
  IV U56729 ( .A(n56688), .Z(n56735) );
  XNOR U56730 ( .A(n56751), .B(n56728), .Z(n56688) );
  XNOR U56731 ( .A(n56752), .B(n56734), .Z(n56728) );
  XNOR U56732 ( .A(n56753), .B(n56754), .Z(n56734) );
  NOR U56733 ( .A(n56755), .B(n56756), .Z(n56754) );
  XOR U56734 ( .A(n56753), .B(n56757), .Z(n56755) );
  XNOR U56735 ( .A(n56733), .B(n56725), .Z(n56752) );
  XOR U56736 ( .A(n56758), .B(n56759), .Z(n56725) );
  AND U56737 ( .A(n56760), .B(n56761), .Z(n56759) );
  XOR U56738 ( .A(n56758), .B(n56762), .Z(n56760) );
  XNOR U56739 ( .A(n56763), .B(n56730), .Z(n56733) );
  XOR U56740 ( .A(n56764), .B(n56765), .Z(n56730) );
  AND U56741 ( .A(n56766), .B(n56767), .Z(n56765) );
  XNOR U56742 ( .A(n56768), .B(n56769), .Z(n56766) );
  IV U56743 ( .A(n56764), .Z(n56768) );
  XNOR U56744 ( .A(n56770), .B(n56771), .Z(n56763) );
  NOR U56745 ( .A(n56772), .B(n56773), .Z(n56771) );
  XNOR U56746 ( .A(n56770), .B(n56774), .Z(n56772) );
  XNOR U56747 ( .A(n56729), .B(n56736), .Z(n56751) );
  NOR U56748 ( .A(n56694), .B(n56775), .Z(n56736) );
  XOR U56749 ( .A(n56741), .B(n56740), .Z(n56729) );
  XNOR U56750 ( .A(n56776), .B(n56737), .Z(n56740) );
  XOR U56751 ( .A(n56777), .B(n56778), .Z(n56737) );
  AND U56752 ( .A(n56779), .B(n56780), .Z(n56778) );
  XNOR U56753 ( .A(n56781), .B(n56782), .Z(n56779) );
  IV U56754 ( .A(n56777), .Z(n56781) );
  XNOR U56755 ( .A(n56783), .B(n56784), .Z(n56776) );
  NOR U56756 ( .A(n56785), .B(n56786), .Z(n56784) );
  XNOR U56757 ( .A(n56783), .B(n56787), .Z(n56785) );
  XOR U56758 ( .A(n56788), .B(n56789), .Z(n56741) );
  NOR U56759 ( .A(n56790), .B(n56791), .Z(n56789) );
  XNOR U56760 ( .A(n56788), .B(n56792), .Z(n56790) );
  XNOR U56761 ( .A(n56685), .B(n56747), .Z(n56749) );
  XNOR U56762 ( .A(n56793), .B(n56794), .Z(n56685) );
  AND U56763 ( .A(n2393), .B(n56795), .Z(n56794) );
  XNOR U56764 ( .A(n56796), .B(n56797), .Z(n56795) );
  AND U56765 ( .A(n56691), .B(n56694), .Z(n56747) );
  XOR U56766 ( .A(n56798), .B(n56775), .Z(n56694) );
  XNOR U56767 ( .A(p_input[1952]), .B(p_input[2048]), .Z(n56775) );
  XNOR U56768 ( .A(n56762), .B(n56761), .Z(n56798) );
  XNOR U56769 ( .A(n56799), .B(n56769), .Z(n56761) );
  XNOR U56770 ( .A(n56757), .B(n56756), .Z(n56769) );
  XNOR U56771 ( .A(n56800), .B(n56753), .Z(n56756) );
  XNOR U56772 ( .A(p_input[1962]), .B(p_input[2058]), .Z(n56753) );
  XOR U56773 ( .A(p_input[1963]), .B(n29030), .Z(n56800) );
  XOR U56774 ( .A(p_input[1964]), .B(p_input[2060]), .Z(n56757) );
  XOR U56775 ( .A(n56767), .B(n56801), .Z(n56799) );
  IV U56776 ( .A(n56758), .Z(n56801) );
  XOR U56777 ( .A(p_input[1953]), .B(p_input[2049]), .Z(n56758) );
  XNOR U56778 ( .A(n56802), .B(n56774), .Z(n56767) );
  XNOR U56779 ( .A(p_input[1967]), .B(n29033), .Z(n56774) );
  XOR U56780 ( .A(n56764), .B(n56773), .Z(n56802) );
  XOR U56781 ( .A(n56803), .B(n56770), .Z(n56773) );
  XOR U56782 ( .A(p_input[1965]), .B(p_input[2061]), .Z(n56770) );
  XOR U56783 ( .A(p_input[1966]), .B(n29035), .Z(n56803) );
  XOR U56784 ( .A(p_input[1961]), .B(p_input[2057]), .Z(n56764) );
  XOR U56785 ( .A(n56782), .B(n56780), .Z(n56762) );
  XNOR U56786 ( .A(n56804), .B(n56787), .Z(n56780) );
  XOR U56787 ( .A(p_input[1960]), .B(p_input[2056]), .Z(n56787) );
  XOR U56788 ( .A(n56777), .B(n56786), .Z(n56804) );
  XOR U56789 ( .A(n56805), .B(n56783), .Z(n56786) );
  XOR U56790 ( .A(p_input[1958]), .B(p_input[2054]), .Z(n56783) );
  XOR U56791 ( .A(p_input[1959]), .B(n30404), .Z(n56805) );
  XOR U56792 ( .A(p_input[1954]), .B(p_input[2050]), .Z(n56777) );
  XNOR U56793 ( .A(n56792), .B(n56791), .Z(n56782) );
  XOR U56794 ( .A(n56806), .B(n56788), .Z(n56791) );
  XOR U56795 ( .A(p_input[1955]), .B(p_input[2051]), .Z(n56788) );
  XOR U56796 ( .A(p_input[1956]), .B(n30406), .Z(n56806) );
  XOR U56797 ( .A(p_input[1957]), .B(p_input[2053]), .Z(n56792) );
  XNOR U56798 ( .A(n56807), .B(n56808), .Z(n56691) );
  AND U56799 ( .A(n2393), .B(n56809), .Z(n56808) );
  XNOR U56800 ( .A(n56810), .B(n56811), .Z(n2393) );
  NOR U56801 ( .A(n56812), .B(n56813), .Z(n56811) );
  XNOR U56802 ( .A(n56810), .B(n56814), .Z(n56813) );
  NOR U56803 ( .A(n56810), .B(n56700), .Z(n56812) );
  XOR U56804 ( .A(n56815), .B(n56816), .Z(n56810) );
  AND U56805 ( .A(n56817), .B(n56818), .Z(n56816) );
  XOR U56806 ( .A(n56717), .B(n56815), .Z(n56818) );
  XOR U56807 ( .A(n56815), .B(n56718), .Z(n56817) );
  XOR U56808 ( .A(n56819), .B(n56820), .Z(n56815) );
  AND U56809 ( .A(n56821), .B(n56822), .Z(n56820) );
  XOR U56810 ( .A(n56745), .B(n56819), .Z(n56822) );
  XOR U56811 ( .A(n56819), .B(n56746), .Z(n56821) );
  XOR U56812 ( .A(n56823), .B(n56824), .Z(n56819) );
  AND U56813 ( .A(n56825), .B(n56826), .Z(n56824) );
  XOR U56814 ( .A(n56823), .B(n56796), .Z(n56826) );
  XNOR U56815 ( .A(n56827), .B(n56828), .Z(n56654) );
  AND U56816 ( .A(n2397), .B(n56829), .Z(n56828) );
  XNOR U56817 ( .A(n56830), .B(n56831), .Z(n2397) );
  NOR U56818 ( .A(n56832), .B(n56833), .Z(n56831) );
  XOR U56819 ( .A(n56626), .B(n56830), .Z(n56833) );
  NOR U56820 ( .A(n56830), .B(n56625), .Z(n56832) );
  XOR U56821 ( .A(n56834), .B(n56835), .Z(n56830) );
  AND U56822 ( .A(n56836), .B(n56837), .Z(n56835) );
  XOR U56823 ( .A(n56834), .B(n56632), .Z(n56836) );
  XOR U56824 ( .A(n56838), .B(n56839), .Z(n56618) );
  AND U56825 ( .A(n2401), .B(n56829), .Z(n56839) );
  XNOR U56826 ( .A(n56827), .B(n56838), .Z(n56829) );
  XNOR U56827 ( .A(n56840), .B(n56841), .Z(n2401) );
  NOR U56828 ( .A(n56842), .B(n56843), .Z(n56841) );
  XNOR U56829 ( .A(n56626), .B(n56844), .Z(n56843) );
  IV U56830 ( .A(n56840), .Z(n56844) );
  AND U56831 ( .A(n56845), .B(n56846), .Z(n56626) );
  NOR U56832 ( .A(n56840), .B(n56625), .Z(n56842) );
  AND U56833 ( .A(n56700), .B(n56699), .Z(n56625) );
  IV U56834 ( .A(n56814), .Z(n56699) );
  XOR U56835 ( .A(n56834), .B(n56847), .Z(n56840) );
  AND U56836 ( .A(n56848), .B(n56837), .Z(n56847) );
  XNOR U56837 ( .A(n56671), .B(n56834), .Z(n56837) );
  XOR U56838 ( .A(n56718), .B(n56849), .Z(n56671) );
  AND U56839 ( .A(n2404), .B(n56850), .Z(n56849) );
  XOR U56840 ( .A(n56714), .B(n56718), .Z(n56850) );
  XNOR U56841 ( .A(n56851), .B(n56834), .Z(n56848) );
  IV U56842 ( .A(n56632), .Z(n56851) );
  XOR U56843 ( .A(n56852), .B(n56853), .Z(n56632) );
  AND U56844 ( .A(n2420), .B(n56854), .Z(n56853) );
  XOR U56845 ( .A(n56855), .B(n56856), .Z(n56834) );
  AND U56846 ( .A(n56857), .B(n56858), .Z(n56856) );
  XNOR U56847 ( .A(n56681), .B(n56855), .Z(n56858) );
  XOR U56848 ( .A(n56746), .B(n56859), .Z(n56681) );
  AND U56849 ( .A(n2404), .B(n56860), .Z(n56859) );
  XOR U56850 ( .A(n56742), .B(n56746), .Z(n56860) );
  XOR U56851 ( .A(n56855), .B(n56641), .Z(n56857) );
  XOR U56852 ( .A(n56861), .B(n56862), .Z(n56641) );
  AND U56853 ( .A(n2420), .B(n56863), .Z(n56862) );
  XOR U56854 ( .A(n56864), .B(n56865), .Z(n56855) );
  AND U56855 ( .A(n56866), .B(n56867), .Z(n56865) );
  XNOR U56856 ( .A(n56864), .B(n56689), .Z(n56867) );
  XOR U56857 ( .A(n56797), .B(n56868), .Z(n56689) );
  AND U56858 ( .A(n2404), .B(n56869), .Z(n56868) );
  XOR U56859 ( .A(n56793), .B(n56797), .Z(n56869) );
  XNOR U56860 ( .A(n56870), .B(n56864), .Z(n56866) );
  IV U56861 ( .A(n56651), .Z(n56870) );
  XOR U56862 ( .A(n56871), .B(n56872), .Z(n56651) );
  AND U56863 ( .A(n2420), .B(n56873), .Z(n56872) );
  AND U56864 ( .A(n56838), .B(n56827), .Z(n56864) );
  XNOR U56865 ( .A(n56874), .B(n56875), .Z(n56827) );
  AND U56866 ( .A(n2404), .B(n56809), .Z(n56875) );
  XNOR U56867 ( .A(n56807), .B(n56874), .Z(n56809) );
  XNOR U56868 ( .A(n56876), .B(n56877), .Z(n2404) );
  NOR U56869 ( .A(n56878), .B(n56879), .Z(n56877) );
  XNOR U56870 ( .A(n56876), .B(n56814), .Z(n56879) );
  NOR U56871 ( .A(n56845), .B(n56846), .Z(n56814) );
  NOR U56872 ( .A(n56876), .B(n56700), .Z(n56878) );
  AND U56873 ( .A(n56880), .B(n56881), .Z(n56700) );
  IV U56874 ( .A(n56882), .Z(n56880) );
  XOR U56875 ( .A(n56883), .B(n56884), .Z(n56876) );
  AND U56876 ( .A(n56885), .B(n56886), .Z(n56884) );
  XNOR U56877 ( .A(n56883), .B(n56714), .Z(n56886) );
  IV U56878 ( .A(n56717), .Z(n56714) );
  XOR U56879 ( .A(n56887), .B(n56888), .Z(n56717) );
  AND U56880 ( .A(n2408), .B(n56889), .Z(n56888) );
  XOR U56881 ( .A(n56890), .B(n56887), .Z(n56889) );
  XOR U56882 ( .A(n56718), .B(n56883), .Z(n56885) );
  XOR U56883 ( .A(n56891), .B(n56892), .Z(n56718) );
  AND U56884 ( .A(n2416), .B(n56854), .Z(n56892) );
  XOR U56885 ( .A(n56891), .B(n56852), .Z(n56854) );
  XOR U56886 ( .A(n56893), .B(n56894), .Z(n56883) );
  AND U56887 ( .A(n56895), .B(n56896), .Z(n56894) );
  XNOR U56888 ( .A(n56893), .B(n56742), .Z(n56896) );
  IV U56889 ( .A(n56745), .Z(n56742) );
  XOR U56890 ( .A(n56897), .B(n56898), .Z(n56745) );
  AND U56891 ( .A(n2408), .B(n56899), .Z(n56898) );
  XNOR U56892 ( .A(n56900), .B(n56897), .Z(n56899) );
  XOR U56893 ( .A(n56746), .B(n56893), .Z(n56895) );
  XOR U56894 ( .A(n56901), .B(n56902), .Z(n56746) );
  AND U56895 ( .A(n2416), .B(n56863), .Z(n56902) );
  XOR U56896 ( .A(n56901), .B(n56861), .Z(n56863) );
  XOR U56897 ( .A(n56823), .B(n56903), .Z(n56893) );
  AND U56898 ( .A(n56825), .B(n56904), .Z(n56903) );
  XNOR U56899 ( .A(n56823), .B(n56793), .Z(n56904) );
  IV U56900 ( .A(n56796), .Z(n56793) );
  XOR U56901 ( .A(n56905), .B(n56906), .Z(n56796) );
  AND U56902 ( .A(n2408), .B(n56907), .Z(n56906) );
  XOR U56903 ( .A(n56908), .B(n56905), .Z(n56907) );
  XOR U56904 ( .A(n56797), .B(n56823), .Z(n56825) );
  XOR U56905 ( .A(n56909), .B(n56910), .Z(n56797) );
  AND U56906 ( .A(n2416), .B(n56873), .Z(n56910) );
  XOR U56907 ( .A(n56909), .B(n56871), .Z(n56873) );
  AND U56908 ( .A(n56874), .B(n56807), .Z(n56823) );
  XNOR U56909 ( .A(n56911), .B(n56912), .Z(n56807) );
  AND U56910 ( .A(n2408), .B(n56913), .Z(n56912) );
  XNOR U56911 ( .A(n56914), .B(n56911), .Z(n56913) );
  XNOR U56912 ( .A(n56915), .B(n56916), .Z(n2408) );
  NOR U56913 ( .A(n56917), .B(n56918), .Z(n56916) );
  XNOR U56914 ( .A(n56915), .B(n56882), .Z(n56918) );
  NOR U56915 ( .A(n56919), .B(n56920), .Z(n56882) );
  NOR U56916 ( .A(n56915), .B(n56881), .Z(n56917) );
  AND U56917 ( .A(n56921), .B(n56922), .Z(n56881) );
  XOR U56918 ( .A(n56923), .B(n56924), .Z(n56915) );
  AND U56919 ( .A(n56925), .B(n56926), .Z(n56924) );
  XNOR U56920 ( .A(n56923), .B(n56921), .Z(n56926) );
  IV U56921 ( .A(n56890), .Z(n56921) );
  XOR U56922 ( .A(n56927), .B(n56928), .Z(n56890) );
  XOR U56923 ( .A(n56929), .B(n56922), .Z(n56928) );
  AND U56924 ( .A(n56900), .B(n56930), .Z(n56922) );
  AND U56925 ( .A(n56931), .B(n56932), .Z(n56929) );
  XOR U56926 ( .A(n56933), .B(n56927), .Z(n56931) );
  XNOR U56927 ( .A(n56887), .B(n56923), .Z(n56925) );
  XNOR U56928 ( .A(n56934), .B(n56935), .Z(n56887) );
  AND U56929 ( .A(n2412), .B(n56936), .Z(n56935) );
  XNOR U56930 ( .A(n56937), .B(n56938), .Z(n56936) );
  XOR U56931 ( .A(n56939), .B(n56940), .Z(n56923) );
  AND U56932 ( .A(n56941), .B(n56942), .Z(n56940) );
  XNOR U56933 ( .A(n56939), .B(n56900), .Z(n56942) );
  XOR U56934 ( .A(n56943), .B(n56932), .Z(n56900) );
  XNOR U56935 ( .A(n56944), .B(n56927), .Z(n56932) );
  XOR U56936 ( .A(n56945), .B(n56946), .Z(n56927) );
  AND U56937 ( .A(n56947), .B(n56948), .Z(n56946) );
  XOR U56938 ( .A(n56949), .B(n56945), .Z(n56947) );
  XNOR U56939 ( .A(n56950), .B(n56951), .Z(n56944) );
  AND U56940 ( .A(n56952), .B(n56953), .Z(n56951) );
  XOR U56941 ( .A(n56950), .B(n56954), .Z(n56952) );
  XNOR U56942 ( .A(n56933), .B(n56930), .Z(n56943) );
  AND U56943 ( .A(n56955), .B(n56956), .Z(n56930) );
  XOR U56944 ( .A(n56957), .B(n56958), .Z(n56933) );
  AND U56945 ( .A(n56959), .B(n56960), .Z(n56958) );
  XOR U56946 ( .A(n56957), .B(n56961), .Z(n56959) );
  XNOR U56947 ( .A(n56897), .B(n56939), .Z(n56941) );
  XNOR U56948 ( .A(n56962), .B(n56963), .Z(n56897) );
  AND U56949 ( .A(n2412), .B(n56964), .Z(n56963) );
  XNOR U56950 ( .A(n56965), .B(n56966), .Z(n56964) );
  XOR U56951 ( .A(n56967), .B(n56968), .Z(n56939) );
  AND U56952 ( .A(n56969), .B(n56970), .Z(n56968) );
  XNOR U56953 ( .A(n56967), .B(n56955), .Z(n56970) );
  IV U56954 ( .A(n56908), .Z(n56955) );
  XNOR U56955 ( .A(n56971), .B(n56948), .Z(n56908) );
  XNOR U56956 ( .A(n56972), .B(n56954), .Z(n56948) );
  XNOR U56957 ( .A(n56973), .B(n56974), .Z(n56954) );
  NOR U56958 ( .A(n56975), .B(n56976), .Z(n56974) );
  XOR U56959 ( .A(n56973), .B(n56977), .Z(n56975) );
  XNOR U56960 ( .A(n56953), .B(n56945), .Z(n56972) );
  XOR U56961 ( .A(n56978), .B(n56979), .Z(n56945) );
  AND U56962 ( .A(n56980), .B(n56981), .Z(n56979) );
  XOR U56963 ( .A(n56978), .B(n56982), .Z(n56980) );
  XNOR U56964 ( .A(n56983), .B(n56950), .Z(n56953) );
  XOR U56965 ( .A(n56984), .B(n56985), .Z(n56950) );
  AND U56966 ( .A(n56986), .B(n56987), .Z(n56985) );
  XNOR U56967 ( .A(n56988), .B(n56989), .Z(n56986) );
  IV U56968 ( .A(n56984), .Z(n56988) );
  XNOR U56969 ( .A(n56990), .B(n56991), .Z(n56983) );
  NOR U56970 ( .A(n56992), .B(n56993), .Z(n56991) );
  XNOR U56971 ( .A(n56990), .B(n56994), .Z(n56992) );
  XNOR U56972 ( .A(n56949), .B(n56956), .Z(n56971) );
  NOR U56973 ( .A(n56914), .B(n56995), .Z(n56956) );
  XOR U56974 ( .A(n56961), .B(n56960), .Z(n56949) );
  XNOR U56975 ( .A(n56996), .B(n56957), .Z(n56960) );
  XOR U56976 ( .A(n56997), .B(n56998), .Z(n56957) );
  AND U56977 ( .A(n56999), .B(n57000), .Z(n56998) );
  XNOR U56978 ( .A(n57001), .B(n57002), .Z(n56999) );
  IV U56979 ( .A(n56997), .Z(n57001) );
  XNOR U56980 ( .A(n57003), .B(n57004), .Z(n56996) );
  NOR U56981 ( .A(n57005), .B(n57006), .Z(n57004) );
  XNOR U56982 ( .A(n57003), .B(n57007), .Z(n57005) );
  XOR U56983 ( .A(n57008), .B(n57009), .Z(n56961) );
  NOR U56984 ( .A(n57010), .B(n57011), .Z(n57009) );
  XNOR U56985 ( .A(n57008), .B(n57012), .Z(n57010) );
  XNOR U56986 ( .A(n56905), .B(n56967), .Z(n56969) );
  XNOR U56987 ( .A(n57013), .B(n57014), .Z(n56905) );
  AND U56988 ( .A(n2412), .B(n57015), .Z(n57014) );
  XNOR U56989 ( .A(n57016), .B(n57017), .Z(n57015) );
  AND U56990 ( .A(n56911), .B(n56914), .Z(n56967) );
  XOR U56991 ( .A(n57018), .B(n56995), .Z(n56914) );
  XNOR U56992 ( .A(p_input[1968]), .B(p_input[2048]), .Z(n56995) );
  XNOR U56993 ( .A(n56982), .B(n56981), .Z(n57018) );
  XNOR U56994 ( .A(n57019), .B(n56989), .Z(n56981) );
  XNOR U56995 ( .A(n56977), .B(n56976), .Z(n56989) );
  XNOR U56996 ( .A(n57020), .B(n56973), .Z(n56976) );
  XNOR U56997 ( .A(p_input[1978]), .B(p_input[2058]), .Z(n56973) );
  XOR U56998 ( .A(p_input[1979]), .B(n29030), .Z(n57020) );
  XOR U56999 ( .A(p_input[1980]), .B(p_input[2060]), .Z(n56977) );
  XOR U57000 ( .A(n56987), .B(n57021), .Z(n57019) );
  IV U57001 ( .A(n56978), .Z(n57021) );
  XOR U57002 ( .A(p_input[1969]), .B(p_input[2049]), .Z(n56978) );
  XNOR U57003 ( .A(n57022), .B(n56994), .Z(n56987) );
  XNOR U57004 ( .A(p_input[1983]), .B(n29033), .Z(n56994) );
  XOR U57005 ( .A(n56984), .B(n56993), .Z(n57022) );
  XOR U57006 ( .A(n57023), .B(n56990), .Z(n56993) );
  XOR U57007 ( .A(p_input[1981]), .B(p_input[2061]), .Z(n56990) );
  XOR U57008 ( .A(p_input[1982]), .B(n29035), .Z(n57023) );
  XOR U57009 ( .A(p_input[1977]), .B(p_input[2057]), .Z(n56984) );
  XOR U57010 ( .A(n57002), .B(n57000), .Z(n56982) );
  XNOR U57011 ( .A(n57024), .B(n57007), .Z(n57000) );
  XOR U57012 ( .A(p_input[1976]), .B(p_input[2056]), .Z(n57007) );
  XOR U57013 ( .A(n56997), .B(n57006), .Z(n57024) );
  XOR U57014 ( .A(n57025), .B(n57003), .Z(n57006) );
  XOR U57015 ( .A(p_input[1974]), .B(p_input[2054]), .Z(n57003) );
  XOR U57016 ( .A(p_input[1975]), .B(n30404), .Z(n57025) );
  XOR U57017 ( .A(p_input[1970]), .B(p_input[2050]), .Z(n56997) );
  XNOR U57018 ( .A(n57012), .B(n57011), .Z(n57002) );
  XOR U57019 ( .A(n57026), .B(n57008), .Z(n57011) );
  XOR U57020 ( .A(p_input[1971]), .B(p_input[2051]), .Z(n57008) );
  XOR U57021 ( .A(p_input[1972]), .B(n30406), .Z(n57026) );
  XOR U57022 ( .A(p_input[1973]), .B(p_input[2053]), .Z(n57012) );
  XNOR U57023 ( .A(n57027), .B(n57028), .Z(n56911) );
  AND U57024 ( .A(n2412), .B(n57029), .Z(n57028) );
  XNOR U57025 ( .A(n57030), .B(n57031), .Z(n2412) );
  NOR U57026 ( .A(n57032), .B(n57033), .Z(n57031) );
  XNOR U57027 ( .A(n57030), .B(n57034), .Z(n57033) );
  NOR U57028 ( .A(n57030), .B(n56920), .Z(n57032) );
  XOR U57029 ( .A(n57035), .B(n57036), .Z(n57030) );
  AND U57030 ( .A(n57037), .B(n57038), .Z(n57036) );
  XOR U57031 ( .A(n56937), .B(n57035), .Z(n57038) );
  XOR U57032 ( .A(n57035), .B(n56938), .Z(n57037) );
  XOR U57033 ( .A(n57039), .B(n57040), .Z(n57035) );
  AND U57034 ( .A(n57041), .B(n57042), .Z(n57040) );
  XOR U57035 ( .A(n56965), .B(n57039), .Z(n57042) );
  XOR U57036 ( .A(n57039), .B(n56966), .Z(n57041) );
  XOR U57037 ( .A(n57043), .B(n57044), .Z(n57039) );
  AND U57038 ( .A(n57045), .B(n57046), .Z(n57044) );
  XOR U57039 ( .A(n57043), .B(n57016), .Z(n57046) );
  XNOR U57040 ( .A(n57047), .B(n57048), .Z(n56874) );
  AND U57041 ( .A(n2416), .B(n57049), .Z(n57048) );
  XNOR U57042 ( .A(n57050), .B(n57051), .Z(n2416) );
  NOR U57043 ( .A(n57052), .B(n57053), .Z(n57051) );
  XOR U57044 ( .A(n56846), .B(n57050), .Z(n57053) );
  NOR U57045 ( .A(n57050), .B(n56845), .Z(n57052) );
  XOR U57046 ( .A(n57054), .B(n57055), .Z(n57050) );
  AND U57047 ( .A(n57056), .B(n57057), .Z(n57055) );
  XOR U57048 ( .A(n57054), .B(n56852), .Z(n57056) );
  XOR U57049 ( .A(n57058), .B(n57059), .Z(n56838) );
  AND U57050 ( .A(n2420), .B(n57049), .Z(n57059) );
  XNOR U57051 ( .A(n57047), .B(n57058), .Z(n57049) );
  XNOR U57052 ( .A(n57060), .B(n57061), .Z(n2420) );
  NOR U57053 ( .A(n57062), .B(n57063), .Z(n57061) );
  XNOR U57054 ( .A(n56846), .B(n57064), .Z(n57063) );
  IV U57055 ( .A(n57060), .Z(n57064) );
  AND U57056 ( .A(n57065), .B(n57066), .Z(n56846) );
  NOR U57057 ( .A(n57060), .B(n56845), .Z(n57062) );
  AND U57058 ( .A(n56920), .B(n56919), .Z(n56845) );
  IV U57059 ( .A(n57034), .Z(n56919) );
  XOR U57060 ( .A(n57054), .B(n57067), .Z(n57060) );
  AND U57061 ( .A(n57068), .B(n57057), .Z(n57067) );
  XNOR U57062 ( .A(n56891), .B(n57054), .Z(n57057) );
  XOR U57063 ( .A(n56938), .B(n57069), .Z(n56891) );
  AND U57064 ( .A(n2423), .B(n57070), .Z(n57069) );
  XOR U57065 ( .A(n56934), .B(n56938), .Z(n57070) );
  XNOR U57066 ( .A(n57071), .B(n57054), .Z(n57068) );
  IV U57067 ( .A(n56852), .Z(n57071) );
  XOR U57068 ( .A(n57072), .B(n57073), .Z(n56852) );
  AND U57069 ( .A(n2438), .B(n57074), .Z(n57073) );
  XOR U57070 ( .A(n57075), .B(n57076), .Z(n57054) );
  AND U57071 ( .A(n57077), .B(n57078), .Z(n57076) );
  XNOR U57072 ( .A(n56901), .B(n57075), .Z(n57078) );
  XOR U57073 ( .A(n56966), .B(n57079), .Z(n56901) );
  AND U57074 ( .A(n2423), .B(n57080), .Z(n57079) );
  XOR U57075 ( .A(n56962), .B(n56966), .Z(n57080) );
  XOR U57076 ( .A(n57075), .B(n56861), .Z(n57077) );
  XOR U57077 ( .A(n57081), .B(n57082), .Z(n56861) );
  AND U57078 ( .A(n2438), .B(n57083), .Z(n57082) );
  XOR U57079 ( .A(n57084), .B(n57085), .Z(n57075) );
  AND U57080 ( .A(n57086), .B(n57087), .Z(n57085) );
  XNOR U57081 ( .A(n57084), .B(n56909), .Z(n57087) );
  XOR U57082 ( .A(n57017), .B(n57088), .Z(n56909) );
  AND U57083 ( .A(n2423), .B(n57089), .Z(n57088) );
  XOR U57084 ( .A(n57013), .B(n57017), .Z(n57089) );
  XNOR U57085 ( .A(n57090), .B(n57084), .Z(n57086) );
  IV U57086 ( .A(n56871), .Z(n57090) );
  XOR U57087 ( .A(n57091), .B(n57092), .Z(n56871) );
  AND U57088 ( .A(n2438), .B(n57093), .Z(n57092) );
  AND U57089 ( .A(n57058), .B(n57047), .Z(n57084) );
  XNOR U57090 ( .A(n57094), .B(n57095), .Z(n57047) );
  AND U57091 ( .A(n2423), .B(n57029), .Z(n57095) );
  XNOR U57092 ( .A(n57027), .B(n57094), .Z(n57029) );
  XNOR U57093 ( .A(n57096), .B(n57097), .Z(n2423) );
  NOR U57094 ( .A(n57098), .B(n57099), .Z(n57097) );
  XNOR U57095 ( .A(n57096), .B(n57034), .Z(n57099) );
  NOR U57096 ( .A(n57065), .B(n57066), .Z(n57034) );
  NOR U57097 ( .A(n57096), .B(n56920), .Z(n57098) );
  AND U57098 ( .A(n57100), .B(n57101), .Z(n56920) );
  IV U57099 ( .A(n57102), .Z(n57100) );
  XOR U57100 ( .A(n57103), .B(n57104), .Z(n57096) );
  AND U57101 ( .A(n57105), .B(n57106), .Z(n57104) );
  XNOR U57102 ( .A(n57103), .B(n56934), .Z(n57106) );
  IV U57103 ( .A(n56937), .Z(n56934) );
  XOR U57104 ( .A(n57107), .B(n57108), .Z(n56937) );
  AND U57105 ( .A(n2427), .B(n57109), .Z(n57108) );
  XOR U57106 ( .A(n57110), .B(n57107), .Z(n57109) );
  XOR U57107 ( .A(n56938), .B(n57103), .Z(n57105) );
  XOR U57108 ( .A(n57111), .B(n57112), .Z(n56938) );
  AND U57109 ( .A(n2434), .B(n57074), .Z(n57112) );
  XOR U57110 ( .A(n57111), .B(n57072), .Z(n57074) );
  XOR U57111 ( .A(n57113), .B(n57114), .Z(n57103) );
  AND U57112 ( .A(n57115), .B(n57116), .Z(n57114) );
  XNOR U57113 ( .A(n57113), .B(n56962), .Z(n57116) );
  IV U57114 ( .A(n56965), .Z(n56962) );
  XOR U57115 ( .A(n57117), .B(n57118), .Z(n56965) );
  AND U57116 ( .A(n2427), .B(n57119), .Z(n57118) );
  XNOR U57117 ( .A(n57120), .B(n57117), .Z(n57119) );
  XOR U57118 ( .A(n56966), .B(n57113), .Z(n57115) );
  XOR U57119 ( .A(n57121), .B(n57122), .Z(n56966) );
  AND U57120 ( .A(n2434), .B(n57083), .Z(n57122) );
  XOR U57121 ( .A(n57121), .B(n57081), .Z(n57083) );
  XOR U57122 ( .A(n57043), .B(n57123), .Z(n57113) );
  AND U57123 ( .A(n57045), .B(n57124), .Z(n57123) );
  XNOR U57124 ( .A(n57043), .B(n57013), .Z(n57124) );
  IV U57125 ( .A(n57016), .Z(n57013) );
  XOR U57126 ( .A(n57125), .B(n57126), .Z(n57016) );
  AND U57127 ( .A(n2427), .B(n57127), .Z(n57126) );
  XOR U57128 ( .A(n57128), .B(n57125), .Z(n57127) );
  XOR U57129 ( .A(n57017), .B(n57043), .Z(n57045) );
  XOR U57130 ( .A(n57129), .B(n57130), .Z(n57017) );
  AND U57131 ( .A(n2434), .B(n57093), .Z(n57130) );
  XOR U57132 ( .A(n57129), .B(n57091), .Z(n57093) );
  AND U57133 ( .A(n57094), .B(n57027), .Z(n57043) );
  XNOR U57134 ( .A(n57131), .B(n57132), .Z(n57027) );
  AND U57135 ( .A(n2427), .B(n57133), .Z(n57132) );
  XNOR U57136 ( .A(n57134), .B(n57131), .Z(n57133) );
  XNOR U57137 ( .A(n57135), .B(n57136), .Z(n2427) );
  NOR U57138 ( .A(n57137), .B(n57138), .Z(n57136) );
  XNOR U57139 ( .A(n57135), .B(n57102), .Z(n57138) );
  NOR U57140 ( .A(n57139), .B(n57140), .Z(n57102) );
  NOR U57141 ( .A(n57135), .B(n57101), .Z(n57137) );
  AND U57142 ( .A(n57141), .B(n57142), .Z(n57101) );
  XOR U57143 ( .A(n57143), .B(n57144), .Z(n57135) );
  AND U57144 ( .A(n57145), .B(n57146), .Z(n57144) );
  XNOR U57145 ( .A(n57143), .B(n57141), .Z(n57146) );
  IV U57146 ( .A(n57110), .Z(n57141) );
  XOR U57147 ( .A(n57147), .B(n57148), .Z(n57110) );
  XOR U57148 ( .A(n57149), .B(n57142), .Z(n57148) );
  AND U57149 ( .A(n57120), .B(n57150), .Z(n57142) );
  AND U57150 ( .A(n57151), .B(n57152), .Z(n57149) );
  XOR U57151 ( .A(n57153), .B(n57147), .Z(n57151) );
  XNOR U57152 ( .A(n57107), .B(n57143), .Z(n57145) );
  XNOR U57153 ( .A(n57154), .B(n57155), .Z(n57107) );
  AND U57154 ( .A(n2430), .B(n57156), .Z(n57155) );
  XOR U57155 ( .A(n57157), .B(n57158), .Z(n57143) );
  AND U57156 ( .A(n57159), .B(n57160), .Z(n57158) );
  XNOR U57157 ( .A(n57157), .B(n57120), .Z(n57160) );
  XOR U57158 ( .A(n57161), .B(n57152), .Z(n57120) );
  XNOR U57159 ( .A(n57162), .B(n57147), .Z(n57152) );
  XOR U57160 ( .A(n57163), .B(n57164), .Z(n57147) );
  AND U57161 ( .A(n57165), .B(n57166), .Z(n57164) );
  XOR U57162 ( .A(n57167), .B(n57163), .Z(n57165) );
  XNOR U57163 ( .A(n57168), .B(n57169), .Z(n57162) );
  AND U57164 ( .A(n57170), .B(n57171), .Z(n57169) );
  XOR U57165 ( .A(n57168), .B(n57172), .Z(n57170) );
  XNOR U57166 ( .A(n57153), .B(n57150), .Z(n57161) );
  AND U57167 ( .A(n57173), .B(n57174), .Z(n57150) );
  XOR U57168 ( .A(n57175), .B(n57176), .Z(n57153) );
  AND U57169 ( .A(n57177), .B(n57178), .Z(n57176) );
  XOR U57170 ( .A(n57175), .B(n57179), .Z(n57177) );
  XNOR U57171 ( .A(n57117), .B(n57157), .Z(n57159) );
  XNOR U57172 ( .A(n57180), .B(n57181), .Z(n57117) );
  AND U57173 ( .A(n2430), .B(n57182), .Z(n57181) );
  XOR U57174 ( .A(n57183), .B(n57184), .Z(n57157) );
  AND U57175 ( .A(n57185), .B(n57186), .Z(n57184) );
  XNOR U57176 ( .A(n57183), .B(n57173), .Z(n57186) );
  IV U57177 ( .A(n57128), .Z(n57173) );
  XNOR U57178 ( .A(n57187), .B(n57166), .Z(n57128) );
  XNOR U57179 ( .A(n57188), .B(n57172), .Z(n57166) );
  XNOR U57180 ( .A(n57189), .B(n57190), .Z(n57172) );
  NOR U57181 ( .A(n57191), .B(n57192), .Z(n57190) );
  XOR U57182 ( .A(n57189), .B(n57193), .Z(n57191) );
  XNOR U57183 ( .A(n57171), .B(n57163), .Z(n57188) );
  XOR U57184 ( .A(n57194), .B(n57195), .Z(n57163) );
  AND U57185 ( .A(n57196), .B(n57197), .Z(n57195) );
  XOR U57186 ( .A(n57194), .B(n57198), .Z(n57196) );
  XNOR U57187 ( .A(n57199), .B(n57168), .Z(n57171) );
  XOR U57188 ( .A(n57200), .B(n57201), .Z(n57168) );
  AND U57189 ( .A(n57202), .B(n57203), .Z(n57201) );
  XNOR U57190 ( .A(n57204), .B(n57205), .Z(n57202) );
  IV U57191 ( .A(n57200), .Z(n57204) );
  XNOR U57192 ( .A(n57206), .B(n57207), .Z(n57199) );
  NOR U57193 ( .A(n57208), .B(n57209), .Z(n57207) );
  XNOR U57194 ( .A(n57206), .B(n57210), .Z(n57208) );
  XNOR U57195 ( .A(n57167), .B(n57174), .Z(n57187) );
  NOR U57196 ( .A(n57134), .B(n57211), .Z(n57174) );
  XOR U57197 ( .A(n57179), .B(n57178), .Z(n57167) );
  XNOR U57198 ( .A(n57212), .B(n57175), .Z(n57178) );
  XOR U57199 ( .A(n57213), .B(n57214), .Z(n57175) );
  AND U57200 ( .A(n57215), .B(n57216), .Z(n57214) );
  XNOR U57201 ( .A(n57217), .B(n57218), .Z(n57215) );
  IV U57202 ( .A(n57213), .Z(n57217) );
  XNOR U57203 ( .A(n57219), .B(n57220), .Z(n57212) );
  NOR U57204 ( .A(n57221), .B(n57222), .Z(n57220) );
  XNOR U57205 ( .A(n57219), .B(n57223), .Z(n57221) );
  XOR U57206 ( .A(n57224), .B(n57225), .Z(n57179) );
  NOR U57207 ( .A(n57226), .B(n57227), .Z(n57225) );
  XNOR U57208 ( .A(n57224), .B(n57228), .Z(n57226) );
  XNOR U57209 ( .A(n57125), .B(n57183), .Z(n57185) );
  XNOR U57210 ( .A(n57229), .B(n57230), .Z(n57125) );
  AND U57211 ( .A(n2430), .B(n57231), .Z(n57230) );
  XNOR U57212 ( .A(n57232), .B(n57233), .Z(n57231) );
  AND U57213 ( .A(n57131), .B(n57134), .Z(n57183) );
  XOR U57214 ( .A(n57234), .B(n57211), .Z(n57134) );
  XNOR U57215 ( .A(p_input[1984]), .B(p_input[2048]), .Z(n57211) );
  XNOR U57216 ( .A(n57198), .B(n57197), .Z(n57234) );
  XNOR U57217 ( .A(n57235), .B(n57205), .Z(n57197) );
  XNOR U57218 ( .A(n57193), .B(n57192), .Z(n57205) );
  XNOR U57219 ( .A(n57236), .B(n57189), .Z(n57192) );
  XNOR U57220 ( .A(p_input[1994]), .B(p_input[2058]), .Z(n57189) );
  XOR U57221 ( .A(p_input[1995]), .B(n29030), .Z(n57236) );
  XOR U57222 ( .A(p_input[1996]), .B(p_input[2060]), .Z(n57193) );
  XOR U57223 ( .A(n57203), .B(n57237), .Z(n57235) );
  IV U57224 ( .A(n57194), .Z(n57237) );
  XOR U57225 ( .A(p_input[1985]), .B(p_input[2049]), .Z(n57194) );
  XNOR U57226 ( .A(n57238), .B(n57210), .Z(n57203) );
  XNOR U57227 ( .A(p_input[1999]), .B(n29033), .Z(n57210) );
  IV U57228 ( .A(p_input[2063]), .Z(n29033) );
  XOR U57229 ( .A(n57200), .B(n57209), .Z(n57238) );
  XOR U57230 ( .A(n57239), .B(n57206), .Z(n57209) );
  XOR U57231 ( .A(p_input[1997]), .B(p_input[2061]), .Z(n57206) );
  XOR U57232 ( .A(p_input[1998]), .B(n29035), .Z(n57239) );
  XOR U57233 ( .A(p_input[1993]), .B(p_input[2057]), .Z(n57200) );
  XOR U57234 ( .A(n57218), .B(n57216), .Z(n57198) );
  XNOR U57235 ( .A(n57240), .B(n57223), .Z(n57216) );
  XOR U57236 ( .A(p_input[1992]), .B(p_input[2056]), .Z(n57223) );
  XOR U57237 ( .A(n57213), .B(n57222), .Z(n57240) );
  XOR U57238 ( .A(n57241), .B(n57219), .Z(n57222) );
  XOR U57239 ( .A(p_input[1990]), .B(p_input[2054]), .Z(n57219) );
  XOR U57240 ( .A(p_input[1991]), .B(n30404), .Z(n57241) );
  XOR U57241 ( .A(p_input[1986]), .B(p_input[2050]), .Z(n57213) );
  XNOR U57242 ( .A(n57228), .B(n57227), .Z(n57218) );
  XOR U57243 ( .A(n57242), .B(n57224), .Z(n57227) );
  XOR U57244 ( .A(p_input[1987]), .B(p_input[2051]), .Z(n57224) );
  XOR U57245 ( .A(p_input[1988]), .B(n30406), .Z(n57242) );
  XOR U57246 ( .A(p_input[1989]), .B(p_input[2053]), .Z(n57228) );
  XNOR U57247 ( .A(n57243), .B(n57244), .Z(n57131) );
  AND U57248 ( .A(n2430), .B(n57245), .Z(n57244) );
  XNOR U57249 ( .A(n57246), .B(n57247), .Z(n2430) );
  NOR U57250 ( .A(n57248), .B(n57249), .Z(n57247) );
  XOR U57251 ( .A(n57246), .B(n57139), .Z(n57249) );
  XNOR U57252 ( .A(n57250), .B(n57251), .Z(n57094) );
  AND U57253 ( .A(n2434), .B(n57252), .Z(n57251) );
  XNOR U57254 ( .A(n57253), .B(n57254), .Z(n2434) );
  NOR U57255 ( .A(n57255), .B(n57256), .Z(n57254) );
  XOR U57256 ( .A(n57066), .B(n57253), .Z(n57256) );
  NOR U57257 ( .A(n57253), .B(n57065), .Z(n57255) );
  XOR U57258 ( .A(n57257), .B(n57258), .Z(n57253) );
  AND U57259 ( .A(n57259), .B(n57260), .Z(n57258) );
  XOR U57260 ( .A(n57257), .B(n57072), .Z(n57259) );
  XOR U57261 ( .A(n57261), .B(n57262), .Z(n57058) );
  AND U57262 ( .A(n2438), .B(n57252), .Z(n57262) );
  XNOR U57263 ( .A(n57250), .B(n57261), .Z(n57252) );
  XNOR U57264 ( .A(n57263), .B(n57264), .Z(n2438) );
  NOR U57265 ( .A(n57265), .B(n57266), .Z(n57264) );
  XNOR U57266 ( .A(n57066), .B(n57267), .Z(n57266) );
  IV U57267 ( .A(n57263), .Z(n57267) );
  AND U57268 ( .A(n57268), .B(n57269), .Z(n57066) );
  NOR U57269 ( .A(n57263), .B(n57065), .Z(n57265) );
  AND U57270 ( .A(n57139), .B(n57140), .Z(n57065) );
  IV U57271 ( .A(n57270), .Z(n57139) );
  XOR U57272 ( .A(n57257), .B(n57271), .Z(n57263) );
  AND U57273 ( .A(n57272), .B(n57260), .Z(n57271) );
  XNOR U57274 ( .A(n57111), .B(n57257), .Z(n57260) );
  XOR U57275 ( .A(n57273), .B(n57274), .Z(n57111) );
  AND U57276 ( .A(n2441), .B(n57156), .Z(n57274) );
  XOR U57277 ( .A(n57154), .B(n57273), .Z(n57156) );
  XNOR U57278 ( .A(n57275), .B(n57257), .Z(n57272) );
  IV U57279 ( .A(n57072), .Z(n57275) );
  XOR U57280 ( .A(n57276), .B(n57277), .Z(n57072) );
  AND U57281 ( .A(n2446), .B(n57278), .Z(n57277) );
  XOR U57282 ( .A(n57279), .B(n57280), .Z(n57257) );
  AND U57283 ( .A(n57281), .B(n57282), .Z(n57280) );
  XNOR U57284 ( .A(n57121), .B(n57279), .Z(n57282) );
  XOR U57285 ( .A(n57283), .B(n57284), .Z(n57121) );
  AND U57286 ( .A(n2441), .B(n57182), .Z(n57284) );
  XOR U57287 ( .A(n57180), .B(n57283), .Z(n57182) );
  XOR U57288 ( .A(n57279), .B(n57081), .Z(n57281) );
  XOR U57289 ( .A(n57285), .B(n57286), .Z(n57081) );
  AND U57290 ( .A(n2446), .B(n57287), .Z(n57286) );
  XOR U57291 ( .A(n57288), .B(n57289), .Z(n57279) );
  AND U57292 ( .A(n57290), .B(n57291), .Z(n57289) );
  XNOR U57293 ( .A(n57288), .B(n57129), .Z(n57291) );
  XOR U57294 ( .A(n57233), .B(n57292), .Z(n57129) );
  AND U57295 ( .A(n2441), .B(n57293), .Z(n57292) );
  XOR U57296 ( .A(n57229), .B(n57233), .Z(n57293) );
  XNOR U57297 ( .A(n57294), .B(n57288), .Z(n57290) );
  IV U57298 ( .A(n57091), .Z(n57294) );
  XOR U57299 ( .A(n57295), .B(n57296), .Z(n57091) );
  AND U57300 ( .A(n2446), .B(n57297), .Z(n57296) );
  AND U57301 ( .A(n57261), .B(n57250), .Z(n57288) );
  XNOR U57302 ( .A(n57298), .B(n57299), .Z(n57250) );
  AND U57303 ( .A(n2441), .B(n57245), .Z(n57299) );
  XOR U57304 ( .A(n57300), .B(n57298), .Z(n57245) );
  XNOR U57305 ( .A(n57246), .B(n57301), .Z(n2441) );
  NOR U57306 ( .A(n57248), .B(n57302), .Z(n57301) );
  XNOR U57307 ( .A(n57246), .B(n57270), .Z(n57302) );
  NOR U57308 ( .A(n57268), .B(n57269), .Z(n57270) );
  NOR U57309 ( .A(n57246), .B(n57140), .Z(n57248) );
  AND U57310 ( .A(n57154), .B(n57303), .Z(n57140) );
  XOR U57311 ( .A(n57304), .B(n57305), .Z(n57246) );
  AND U57312 ( .A(n57306), .B(n57307), .Z(n57305) );
  XNOR U57313 ( .A(n57154), .B(n57304), .Z(n57307) );
  XNOR U57314 ( .A(n57308), .B(n57309), .Z(n57154) );
  XOR U57315 ( .A(n57310), .B(n57303), .Z(n57309) );
  AND U57316 ( .A(n57180), .B(n57311), .Z(n57303) );
  AND U57317 ( .A(n57312), .B(n57313), .Z(n57310) );
  XOR U57318 ( .A(n57314), .B(n57308), .Z(n57312) );
  XOR U57319 ( .A(n57304), .B(n57273), .Z(n57306) );
  XOR U57320 ( .A(n57315), .B(n57316), .Z(n57273) );
  AND U57321 ( .A(n2443), .B(n57278), .Z(n57316) );
  XOR U57322 ( .A(n57315), .B(n57276), .Z(n57278) );
  XOR U57323 ( .A(n57317), .B(n57318), .Z(n57304) );
  AND U57324 ( .A(n57319), .B(n57320), .Z(n57318) );
  XNOR U57325 ( .A(n57180), .B(n57317), .Z(n57320) );
  XOR U57326 ( .A(n57321), .B(n57313), .Z(n57180) );
  XNOR U57327 ( .A(n57322), .B(n57308), .Z(n57313) );
  XOR U57328 ( .A(n57323), .B(n57324), .Z(n57308) );
  AND U57329 ( .A(n57325), .B(n57326), .Z(n57324) );
  XOR U57330 ( .A(n57327), .B(n57323), .Z(n57325) );
  XNOR U57331 ( .A(n57328), .B(n57329), .Z(n57322) );
  AND U57332 ( .A(n57330), .B(n57331), .Z(n57329) );
  XOR U57333 ( .A(n57328), .B(n57332), .Z(n57330) );
  XNOR U57334 ( .A(n57314), .B(n57311), .Z(n57321) );
  AND U57335 ( .A(n57229), .B(n57333), .Z(n57311) );
  XOR U57336 ( .A(n57334), .B(n57335), .Z(n57314) );
  AND U57337 ( .A(n57336), .B(n57337), .Z(n57335) );
  XOR U57338 ( .A(n57334), .B(n57338), .Z(n57336) );
  XOR U57339 ( .A(n57317), .B(n57283), .Z(n57319) );
  XOR U57340 ( .A(n57339), .B(n57340), .Z(n57283) );
  AND U57341 ( .A(n2443), .B(n57287), .Z(n57340) );
  XOR U57342 ( .A(n57339), .B(n57285), .Z(n57287) );
  XOR U57343 ( .A(n57341), .B(n57342), .Z(n57317) );
  AND U57344 ( .A(n57343), .B(n57344), .Z(n57342) );
  XNOR U57345 ( .A(n57341), .B(n57229), .Z(n57344) );
  IV U57346 ( .A(n57232), .Z(n57229) );
  XNOR U57347 ( .A(n57345), .B(n57326), .Z(n57232) );
  XNOR U57348 ( .A(n57346), .B(n57332), .Z(n57326) );
  XOR U57349 ( .A(n57347), .B(n57348), .Z(n57332) );
  NOR U57350 ( .A(n57349), .B(n57350), .Z(n57348) );
  XNOR U57351 ( .A(n57347), .B(n57351), .Z(n57349) );
  XNOR U57352 ( .A(n57331), .B(n57323), .Z(n57346) );
  XOR U57353 ( .A(n57352), .B(n57353), .Z(n57323) );
  AND U57354 ( .A(n57354), .B(n57355), .Z(n57353) );
  XNOR U57355 ( .A(n57352), .B(n57356), .Z(n57354) );
  XNOR U57356 ( .A(n57357), .B(n57328), .Z(n57331) );
  XOR U57357 ( .A(n57358), .B(n57359), .Z(n57328) );
  AND U57358 ( .A(n57360), .B(n57361), .Z(n57359) );
  XOR U57359 ( .A(n57358), .B(n57362), .Z(n57360) );
  XNOR U57360 ( .A(n57363), .B(n57364), .Z(n57357) );
  NOR U57361 ( .A(n57365), .B(n57366), .Z(n57364) );
  XOR U57362 ( .A(n57363), .B(n57367), .Z(n57365) );
  XNOR U57363 ( .A(n57327), .B(n57333), .Z(n57345) );
  AND U57364 ( .A(n57300), .B(n57368), .Z(n57333) );
  IV U57365 ( .A(n57243), .Z(n57300) );
  XOR U57366 ( .A(n57338), .B(n57337), .Z(n57327) );
  XNOR U57367 ( .A(n57369), .B(n57334), .Z(n57337) );
  XOR U57368 ( .A(n57370), .B(n57371), .Z(n57334) );
  AND U57369 ( .A(n57372), .B(n57373), .Z(n57371) );
  XOR U57370 ( .A(n57370), .B(n57374), .Z(n57372) );
  XNOR U57371 ( .A(n57375), .B(n57376), .Z(n57369) );
  NOR U57372 ( .A(n57377), .B(n57378), .Z(n57376) );
  XNOR U57373 ( .A(n57375), .B(n57379), .Z(n57377) );
  XOR U57374 ( .A(n57380), .B(n57381), .Z(n57338) );
  NOR U57375 ( .A(n57382), .B(n57383), .Z(n57381) );
  XNOR U57376 ( .A(n57380), .B(n57384), .Z(n57382) );
  XOR U57377 ( .A(n57233), .B(n57341), .Z(n57343) );
  XOR U57378 ( .A(n57385), .B(n57386), .Z(n57233) );
  AND U57379 ( .A(n2443), .B(n57297), .Z(n57386) );
  XOR U57380 ( .A(n57385), .B(n57295), .Z(n57297) );
  AND U57381 ( .A(n57298), .B(n57243), .Z(n57341) );
  XNOR U57382 ( .A(n57387), .B(n57368), .Z(n57243) );
  XOR U57383 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[2048]), .Z(n57368) );
  XOR U57384 ( .A(n57356), .B(n57355), .Z(n57387) );
  XNOR U57385 ( .A(n57388), .B(n57362), .Z(n57355) );
  XNOR U57386 ( .A(n57351), .B(n57350), .Z(n57362) );
  XOR U57387 ( .A(n57389), .B(n57347), .Z(n57350) );
  XNOR U57388 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n29266), 
        .Z(n57347) );
  XOR U57389 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n29030), 
        .Z(n57389) );
  XOR U57390 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(
        p_input[2060]), .Z(n57351) );
  XNOR U57391 ( .A(n57361), .B(n57352), .Z(n57388) );
  XNOR U57392 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n29494), 
        .Z(n57352) );
  XOR U57393 ( .A(n57390), .B(n57367), .Z(n57361) );
  XNOR U57394 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(
        p_input[2063]), .Z(n57367) );
  XOR U57395 ( .A(n57358), .B(n57366), .Z(n57390) );
  XOR U57396 ( .A(n57391), .B(n57363), .Z(n57366) );
  XOR U57397 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[2061]), .Z(n57363) );
  XOR U57398 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n29035), 
        .Z(n57391) );
  XNOR U57399 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n29036), 
        .Z(n57358) );
  IV U57400 ( .A(p_input[2057]), .Z(n29036) );
  XNOR U57401 ( .A(n57374), .B(n57373), .Z(n57356) );
  XNOR U57402 ( .A(n57392), .B(n57379), .Z(n57373) );
  XOR U57403 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(
        p_input[2056]), .Z(n57379) );
  XOR U57404 ( .A(n57370), .B(n57378), .Z(n57392) );
  XOR U57405 ( .A(n57393), .B(n57375), .Z(n57378) );
  XOR U57406 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[2054]), .Z(n57375) );
  XOR U57407 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n30404), 
        .Z(n57393) );
  XNOR U57408 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n29039), 
        .Z(n57370) );
  XNOR U57409 ( .A(n57384), .B(n57383), .Z(n57374) );
  XOR U57410 ( .A(n57394), .B(n57380), .Z(n57383) );
  XOR U57411 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(
        p_input[2051]), .Z(n57380) );
  XOR U57412 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n30406), 
        .Z(n57394) );
  XOR U57413 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(
        p_input[2053]), .Z(n57384) );
  XNOR U57414 ( .A(n57395), .B(n57396), .Z(n57298) );
  AND U57415 ( .A(n2443), .B(n57397), .Z(n57396) );
  XNOR U57416 ( .A(n57398), .B(n57399), .Z(n2443) );
  NOR U57417 ( .A(n57400), .B(n57401), .Z(n57399) );
  XOR U57418 ( .A(n57269), .B(n57398), .Z(n57401) );
  NOR U57419 ( .A(n57398), .B(n57268), .Z(n57400) );
  XOR U57420 ( .A(n57402), .B(n57403), .Z(n57398) );
  AND U57421 ( .A(n57404), .B(n57405), .Z(n57403) );
  XOR U57422 ( .A(n57402), .B(n57276), .Z(n57404) );
  XOR U57423 ( .A(n57406), .B(n57407), .Z(n57261) );
  AND U57424 ( .A(n2446), .B(n57397), .Z(n57407) );
  XOR U57425 ( .A(n57408), .B(n57406), .Z(n57397) );
  XNOR U57426 ( .A(n57409), .B(n57410), .Z(n2446) );
  NOR U57427 ( .A(n57411), .B(n57412), .Z(n57410) );
  XNOR U57428 ( .A(n57269), .B(n57413), .Z(n57412) );
  IV U57429 ( .A(n57409), .Z(n57413) );
  AND U57430 ( .A(n57276), .B(n57414), .Z(n57269) );
  NOR U57431 ( .A(n57409), .B(n57268), .Z(n57411) );
  AND U57432 ( .A(n57315), .B(n57415), .Z(n57268) );
  XOR U57433 ( .A(n57402), .B(n57416), .Z(n57409) );
  AND U57434 ( .A(n57417), .B(n57405), .Z(n57416) );
  XNOR U57435 ( .A(n57315), .B(n57402), .Z(n57405) );
  XNOR U57436 ( .A(n57418), .B(n57419), .Z(n57315) );
  XOR U57437 ( .A(n57420), .B(n57415), .Z(n57419) );
  AND U57438 ( .A(n57339), .B(n57421), .Z(n57415) );
  AND U57439 ( .A(n57422), .B(n57423), .Z(n57420) );
  XOR U57440 ( .A(n57424), .B(n57418), .Z(n57422) );
  XNOR U57441 ( .A(n57425), .B(n57402), .Z(n57417) );
  IV U57442 ( .A(n57276), .Z(n57425) );
  XNOR U57443 ( .A(n57426), .B(n57427), .Z(n57276) );
  XOR U57444 ( .A(n57428), .B(n57414), .Z(n57427) );
  AND U57445 ( .A(n57285), .B(n57429), .Z(n57414) );
  AND U57446 ( .A(n57430), .B(n57431), .Z(n57428) );
  XNOR U57447 ( .A(n57426), .B(n57432), .Z(n57430) );
  XOR U57448 ( .A(n57433), .B(n57434), .Z(n57402) );
  AND U57449 ( .A(n57435), .B(n57436), .Z(n57434) );
  XNOR U57450 ( .A(n57339), .B(n57433), .Z(n57436) );
  XOR U57451 ( .A(n57437), .B(n57423), .Z(n57339) );
  XNOR U57452 ( .A(n57438), .B(n57418), .Z(n57423) );
  XOR U57453 ( .A(n57439), .B(n57440), .Z(n57418) );
  AND U57454 ( .A(n57441), .B(n57442), .Z(n57440) );
  XOR U57455 ( .A(n57443), .B(n57439), .Z(n57441) );
  XNOR U57456 ( .A(n57444), .B(n57445), .Z(n57438) );
  AND U57457 ( .A(n57446), .B(n57447), .Z(n57445) );
  XOR U57458 ( .A(n57444), .B(n57448), .Z(n57446) );
  XNOR U57459 ( .A(n57424), .B(n57421), .Z(n57437) );
  AND U57460 ( .A(n57385), .B(n57449), .Z(n57421) );
  XOR U57461 ( .A(n57450), .B(n57451), .Z(n57424) );
  AND U57462 ( .A(n57452), .B(n57453), .Z(n57451) );
  XOR U57463 ( .A(n57450), .B(n57454), .Z(n57452) );
  XOR U57464 ( .A(n57433), .B(n57285), .Z(n57435) );
  XNOR U57465 ( .A(n57455), .B(n57432), .Z(n57285) );
  XNOR U57466 ( .A(n57456), .B(n57457), .Z(n57432) );
  AND U57467 ( .A(n57458), .B(n57459), .Z(n57457) );
  XOR U57468 ( .A(n57456), .B(n57460), .Z(n57458) );
  XNOR U57469 ( .A(n57431), .B(n57429), .Z(n57455) );
  AND U57470 ( .A(n57295), .B(n57461), .Z(n57429) );
  XNOR U57471 ( .A(n57462), .B(n57426), .Z(n57431) );
  XOR U57472 ( .A(n57463), .B(n57464), .Z(n57426) );
  AND U57473 ( .A(n57465), .B(n57466), .Z(n57464) );
  XOR U57474 ( .A(n57463), .B(n57467), .Z(n57465) );
  XNOR U57475 ( .A(n57468), .B(n57469), .Z(n57462) );
  AND U57476 ( .A(n57470), .B(n57471), .Z(n57469) );
  XNOR U57477 ( .A(n57468), .B(n57472), .Z(n57470) );
  XOR U57478 ( .A(n57473), .B(n57474), .Z(n57433) );
  AND U57479 ( .A(n57475), .B(n57476), .Z(n57474) );
  XNOR U57480 ( .A(n57473), .B(n57385), .Z(n57476) );
  XOR U57481 ( .A(n57477), .B(n57442), .Z(n57385) );
  XNOR U57482 ( .A(n57478), .B(n57448), .Z(n57442) );
  XOR U57483 ( .A(n57479), .B(n57480), .Z(n57448) );
  NOR U57484 ( .A(n57481), .B(n57482), .Z(n57480) );
  XNOR U57485 ( .A(n57479), .B(n57483), .Z(n57481) );
  XNOR U57486 ( .A(n57447), .B(n57439), .Z(n57478) );
  XOR U57487 ( .A(n57484), .B(n57485), .Z(n57439) );
  AND U57488 ( .A(n57486), .B(n57487), .Z(n57485) );
  XNOR U57489 ( .A(n57484), .B(n57488), .Z(n57486) );
  XNOR U57490 ( .A(n57489), .B(n57444), .Z(n57447) );
  XOR U57491 ( .A(n57490), .B(n57491), .Z(n57444) );
  AND U57492 ( .A(n57492), .B(n57493), .Z(n57491) );
  XOR U57493 ( .A(n57490), .B(n57494), .Z(n57492) );
  XNOR U57494 ( .A(n57495), .B(n57496), .Z(n57489) );
  NOR U57495 ( .A(n57497), .B(n57498), .Z(n57496) );
  XOR U57496 ( .A(n57495), .B(n57499), .Z(n57497) );
  XNOR U57497 ( .A(n57443), .B(n57449), .Z(n57477) );
  AND U57498 ( .A(n57408), .B(n57500), .Z(n57449) );
  IV U57499 ( .A(n57395), .Z(n57408) );
  XOR U57500 ( .A(n57454), .B(n57453), .Z(n57443) );
  XNOR U57501 ( .A(n57501), .B(n57450), .Z(n57453) );
  XOR U57502 ( .A(n57502), .B(n57503), .Z(n57450) );
  AND U57503 ( .A(n57504), .B(n57505), .Z(n57503) );
  XOR U57504 ( .A(n57502), .B(n57506), .Z(n57504) );
  XNOR U57505 ( .A(n57507), .B(n57508), .Z(n57501) );
  NOR U57506 ( .A(n57509), .B(n57510), .Z(n57508) );
  XNOR U57507 ( .A(n57507), .B(n57511), .Z(n57509) );
  XOR U57508 ( .A(n57512), .B(n57513), .Z(n57454) );
  NOR U57509 ( .A(n57514), .B(n57515), .Z(n57513) );
  XNOR U57510 ( .A(n57512), .B(n57516), .Z(n57514) );
  XNOR U57511 ( .A(n57517), .B(n57473), .Z(n57475) );
  IV U57512 ( .A(n57295), .Z(n57517) );
  XOR U57513 ( .A(n57518), .B(n57467), .Z(n57295) );
  XOR U57514 ( .A(n57460), .B(n57459), .Z(n57467) );
  XNOR U57515 ( .A(n57519), .B(n57456), .Z(n57459) );
  XOR U57516 ( .A(n57520), .B(n57521), .Z(n57456) );
  AND U57517 ( .A(n57522), .B(n57523), .Z(n57521) );
  XOR U57518 ( .A(n57520), .B(n57524), .Z(n57522) );
  XNOR U57519 ( .A(n57525), .B(n57526), .Z(n57519) );
  NOR U57520 ( .A(n57527), .B(n57528), .Z(n57526) );
  XNOR U57521 ( .A(n57525), .B(n57529), .Z(n57527) );
  XOR U57522 ( .A(n57530), .B(n57531), .Z(n57460) );
  NOR U57523 ( .A(n57532), .B(n57533), .Z(n57531) );
  XNOR U57524 ( .A(n57530), .B(n57534), .Z(n57532) );
  XNOR U57525 ( .A(n57466), .B(n57461), .Z(n57518) );
  AND U57526 ( .A(n57406), .B(n57535), .Z(n57461) );
  XOR U57527 ( .A(n57536), .B(n57472), .Z(n57466) );
  XNOR U57528 ( .A(n57537), .B(n57538), .Z(n57472) );
  NOR U57529 ( .A(n57539), .B(n57540), .Z(n57538) );
  XNOR U57530 ( .A(n57537), .B(n57541), .Z(n57539) );
  XNOR U57531 ( .A(n57471), .B(n57463), .Z(n57536) );
  XOR U57532 ( .A(n57542), .B(n57543), .Z(n57463) );
  AND U57533 ( .A(n57544), .B(n57545), .Z(n57543) );
  XOR U57534 ( .A(n57542), .B(n57546), .Z(n57544) );
  XNOR U57535 ( .A(n57547), .B(n57468), .Z(n57471) );
  XOR U57536 ( .A(n57548), .B(n57549), .Z(n57468) );
  AND U57537 ( .A(n57550), .B(n57551), .Z(n57549) );
  XOR U57538 ( .A(n57548), .B(n57552), .Z(n57550) );
  XNOR U57539 ( .A(n57553), .B(n57554), .Z(n57547) );
  NOR U57540 ( .A(n57555), .B(n57556), .Z(n57554) );
  XOR U57541 ( .A(n57553), .B(n57557), .Z(n57555) );
  AND U57542 ( .A(n57406), .B(n57395), .Z(n57473) );
  XNOR U57543 ( .A(n57558), .B(n57500), .Z(n57395) );
  XOR U57544 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[2048]), .Z(n57500) );
  XOR U57545 ( .A(n57488), .B(n57487), .Z(n57558) );
  XNOR U57546 ( .A(n57559), .B(n57494), .Z(n57487) );
  XNOR U57547 ( .A(n57483), .B(n57482), .Z(n57494) );
  XOR U57548 ( .A(n57560), .B(n57479), .Z(n57482) );
  XNOR U57549 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n29266), 
        .Z(n57479) );
  XOR U57550 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n29030), 
        .Z(n57560) );
  XOR U57551 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(
        p_input[2060]), .Z(n57483) );
  XNOR U57552 ( .A(n57493), .B(n57484), .Z(n57559) );
  XNOR U57553 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n29494), 
        .Z(n57484) );
  XOR U57554 ( .A(n57561), .B(n57499), .Z(n57493) );
  XNOR U57555 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(
        p_input[2063]), .Z(n57499) );
  XOR U57556 ( .A(n57490), .B(n57498), .Z(n57561) );
  XOR U57557 ( .A(n57562), .B(n57495), .Z(n57498) );
  XOR U57558 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[2061]), .Z(n57495) );
  XOR U57559 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n29035), 
        .Z(n57562) );
  XNOR U57560 ( .A(n2448), .B(p_input[2057]), .Z(n57490) );
  IV U57561 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n2448) );
  XNOR U57562 ( .A(n57506), .B(n57505), .Z(n57488) );
  XNOR U57563 ( .A(n57563), .B(n57511), .Z(n57505) );
  XNOR U57564 ( .A(n4207), .B(p_input[2056]), .Z(n57511) );
  IV U57565 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n4207) );
  XOR U57566 ( .A(n57502), .B(n57510), .Z(n57563) );
  XOR U57567 ( .A(n57564), .B(n57507), .Z(n57510) );
  XNOR U57568 ( .A(n7725), .B(p_input[2054]), .Z(n57507) );
  IV U57569 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n7725) );
  XOR U57570 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n30404), 
        .Z(n57564) );
  XNOR U57571 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n29039), 
        .Z(n57502) );
  XNOR U57572 ( .A(n57516), .B(n57515), .Z(n57506) );
  XOR U57573 ( .A(n57565), .B(n57512), .Z(n57515) );
  XNOR U57574 ( .A(n13004), .B(p_input[2051]), .Z(n57512) );
  IV U57575 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n13004) );
  XOR U57576 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n30406), 
        .Z(n57565) );
  XNOR U57577 ( .A(n9484), .B(p_input[2053]), .Z(n57516) );
  IV U57578 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n9484) );
  XOR U57579 ( .A(n57566), .B(n57546), .Z(n57406) );
  XOR U57580 ( .A(n57524), .B(n57523), .Z(n57546) );
  XNOR U57581 ( .A(n57567), .B(n57529), .Z(n57523) );
  XNOR U57582 ( .A(n4206), .B(p_input[2056]), .Z(n57529) );
  IV U57583 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n4206) );
  XOR U57584 ( .A(n57520), .B(n57528), .Z(n57567) );
  XOR U57585 ( .A(n57568), .B(n57525), .Z(n57528) );
  XNOR U57586 ( .A(n7724), .B(p_input[2054]), .Z(n57525) );
  IV U57587 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n7724) );
  XOR U57588 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n30404), .Z(n57568) );
  IV U57589 ( .A(p_input[2055]), .Z(n30404) );
  XNOR U57590 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n29039), .Z(n57520) );
  IV U57591 ( .A(p_input[2050]), .Z(n29039) );
  XNOR U57592 ( .A(n57534), .B(n57533), .Z(n57524) );
  XOR U57593 ( .A(n57569), .B(n57530), .Z(n57533) );
  XNOR U57594 ( .A(n13003), .B(p_input[2051]), .Z(n57530) );
  IV U57595 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n13003) );
  XOR U57596 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n30406), .Z(n57569) );
  IV U57597 ( .A(p_input[2052]), .Z(n30406) );
  XNOR U57598 ( .A(n9483), .B(p_input[2053]), .Z(n57534) );
  IV U57599 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n9483) );
  XNOR U57600 ( .A(n57545), .B(n57535), .Z(n57566) );
  XOR U57601 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[2048]), .Z(n57535) );
  XNOR U57602 ( .A(n57570), .B(n57552), .Z(n57545) );
  XNOR U57603 ( .A(n57541), .B(n57540), .Z(n57552) );
  XOR U57604 ( .A(n57571), .B(n57537), .Z(n57540) );
  XNOR U57605 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n29266), .Z(n57537) );
  IV U57606 ( .A(p_input[2058]), .Z(n29266) );
  XOR U57607 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n29030), .Z(n57571) );
  IV U57608 ( .A(p_input[2059]), .Z(n29030) );
  XOR U57609 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[2060]), .Z(
        n57541) );
  XNOR U57610 ( .A(n57551), .B(n57542), .Z(n57570) );
  XNOR U57611 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n29494), .Z(n57542) );
  IV U57612 ( .A(p_input[2049]), .Z(n29494) );
  XOR U57613 ( .A(n57572), .B(n57557), .Z(n57551) );
  XNOR U57614 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[2063]), .Z(
        n57557) );
  XOR U57615 ( .A(n57548), .B(n57556), .Z(n57572) );
  XOR U57616 ( .A(n57573), .B(n57553), .Z(n57556) );
  XOR U57617 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[2061]), .Z(
        n57553) );
  XOR U57618 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n29035), .Z(n57573) );
  IV U57619 ( .A(p_input[2062]), .Z(n29035) );
  XNOR U57620 ( .A(n2447), .B(p_input[2057]), .Z(n57548) );
  IV U57621 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n2447) );
endmodule

