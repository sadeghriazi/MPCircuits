
module knn_comb_BMR_W16_K1_N128 ( p_input, o );
  input [2063:0] p_input;
  output [15:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703;
  assign \knn_comb_/min_val_out[0][0]  = p_input[2032];
  assign \knn_comb_/min_val_out[0][1]  = p_input[2033];
  assign \knn_comb_/min_val_out[0][2]  = p_input[2034];
  assign \knn_comb_/min_val_out[0][3]  = p_input[2035];
  assign \knn_comb_/min_val_out[0][4]  = p_input[2036];
  assign \knn_comb_/min_val_out[0][5]  = p_input[2037];
  assign \knn_comb_/min_val_out[0][6]  = p_input[2038];
  assign \knn_comb_/min_val_out[0][7]  = p_input[2039];
  assign \knn_comb_/min_val_out[0][8]  = p_input[2040];
  assign \knn_comb_/min_val_out[0][9]  = p_input[2041];
  assign \knn_comb_/min_val_out[0][10]  = p_input[2042];
  assign \knn_comb_/min_val_out[0][11]  = p_input[2043];
  assign \knn_comb_/min_val_out[0][12]  = p_input[2044];
  assign \knn_comb_/min_val_out[0][13]  = p_input[2045];
  assign \knn_comb_/min_val_out[0][14]  = p_input[2046];
  assign \knn_comb_/min_val_out[0][15]  = p_input[2047];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[25]), .B(n5), .Z(n8) );
  XOR U7 ( .A(n9), .B(n10), .Z(n5) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(p_input[41]), .B(n9), .Z(n12) );
  XOR U10 ( .A(n13), .B(n14), .Z(n9) );
  AND U11 ( .A(n15), .B(n16), .Z(n14) );
  XNOR U12 ( .A(p_input[57]), .B(n13), .Z(n16) );
  XOR U13 ( .A(n17), .B(n18), .Z(n13) );
  AND U14 ( .A(n19), .B(n20), .Z(n18) );
  XNOR U15 ( .A(p_input[73]), .B(n17), .Z(n20) );
  XOR U16 ( .A(n21), .B(n22), .Z(n17) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U18 ( .A(p_input[89]), .B(n21), .Z(n24) );
  XOR U19 ( .A(n25), .B(n26), .Z(n21) );
  AND U20 ( .A(n27), .B(n28), .Z(n26) );
  XNOR U21 ( .A(p_input[105]), .B(n25), .Z(n28) );
  XOR U22 ( .A(n29), .B(n30), .Z(n25) );
  AND U23 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U24 ( .A(p_input[121]), .B(n29), .Z(n32) );
  XOR U25 ( .A(n33), .B(n34), .Z(n29) );
  AND U26 ( .A(n35), .B(n36), .Z(n34) );
  XNOR U27 ( .A(p_input[137]), .B(n33), .Z(n36) );
  XOR U28 ( .A(n37), .B(n38), .Z(n33) );
  AND U29 ( .A(n39), .B(n40), .Z(n38) );
  XNOR U30 ( .A(p_input[153]), .B(n37), .Z(n40) );
  XOR U31 ( .A(n41), .B(n42), .Z(n37) );
  AND U32 ( .A(n43), .B(n44), .Z(n42) );
  XNOR U33 ( .A(p_input[169]), .B(n41), .Z(n44) );
  XOR U34 ( .A(n45), .B(n46), .Z(n41) );
  AND U35 ( .A(n47), .B(n48), .Z(n46) );
  XNOR U36 ( .A(p_input[185]), .B(n45), .Z(n48) );
  XOR U37 ( .A(n49), .B(n50), .Z(n45) );
  AND U38 ( .A(n51), .B(n52), .Z(n50) );
  XNOR U39 ( .A(p_input[201]), .B(n49), .Z(n52) );
  XOR U40 ( .A(n53), .B(n54), .Z(n49) );
  AND U41 ( .A(n55), .B(n56), .Z(n54) );
  XNOR U42 ( .A(p_input[217]), .B(n53), .Z(n56) );
  XOR U43 ( .A(n57), .B(n58), .Z(n53) );
  AND U44 ( .A(n59), .B(n60), .Z(n58) );
  XNOR U45 ( .A(p_input[233]), .B(n57), .Z(n60) );
  XOR U46 ( .A(n61), .B(n62), .Z(n57) );
  AND U47 ( .A(n63), .B(n64), .Z(n62) );
  XNOR U48 ( .A(p_input[249]), .B(n61), .Z(n64) );
  XOR U49 ( .A(n65), .B(n66), .Z(n61) );
  AND U50 ( .A(n67), .B(n68), .Z(n66) );
  XNOR U51 ( .A(p_input[265]), .B(n65), .Z(n68) );
  XOR U52 ( .A(n69), .B(n70), .Z(n65) );
  AND U53 ( .A(n71), .B(n72), .Z(n70) );
  XNOR U54 ( .A(p_input[281]), .B(n69), .Z(n72) );
  XOR U55 ( .A(n73), .B(n74), .Z(n69) );
  AND U56 ( .A(n75), .B(n76), .Z(n74) );
  XNOR U57 ( .A(p_input[297]), .B(n73), .Z(n76) );
  XOR U58 ( .A(n77), .B(n78), .Z(n73) );
  AND U59 ( .A(n79), .B(n80), .Z(n78) );
  XNOR U60 ( .A(p_input[313]), .B(n77), .Z(n80) );
  XOR U61 ( .A(n81), .B(n82), .Z(n77) );
  AND U62 ( .A(n83), .B(n84), .Z(n82) );
  XNOR U63 ( .A(p_input[329]), .B(n81), .Z(n84) );
  XOR U64 ( .A(n85), .B(n86), .Z(n81) );
  AND U65 ( .A(n87), .B(n88), .Z(n86) );
  XNOR U66 ( .A(p_input[345]), .B(n85), .Z(n88) );
  XOR U67 ( .A(n89), .B(n90), .Z(n85) );
  AND U68 ( .A(n91), .B(n92), .Z(n90) );
  XNOR U69 ( .A(p_input[361]), .B(n89), .Z(n92) );
  XOR U70 ( .A(n93), .B(n94), .Z(n89) );
  AND U71 ( .A(n95), .B(n96), .Z(n94) );
  XNOR U72 ( .A(p_input[377]), .B(n93), .Z(n96) );
  XOR U73 ( .A(n97), .B(n98), .Z(n93) );
  AND U74 ( .A(n99), .B(n100), .Z(n98) );
  XNOR U75 ( .A(p_input[393]), .B(n97), .Z(n100) );
  XOR U76 ( .A(n101), .B(n102), .Z(n97) );
  AND U77 ( .A(n103), .B(n104), .Z(n102) );
  XNOR U78 ( .A(p_input[409]), .B(n101), .Z(n104) );
  XOR U79 ( .A(n105), .B(n106), .Z(n101) );
  AND U80 ( .A(n107), .B(n108), .Z(n106) );
  XNOR U81 ( .A(p_input[425]), .B(n105), .Z(n108) );
  XOR U82 ( .A(n109), .B(n110), .Z(n105) );
  AND U83 ( .A(n111), .B(n112), .Z(n110) );
  XNOR U84 ( .A(p_input[441]), .B(n109), .Z(n112) );
  XOR U85 ( .A(n113), .B(n114), .Z(n109) );
  AND U86 ( .A(n115), .B(n116), .Z(n114) );
  XNOR U87 ( .A(p_input[457]), .B(n113), .Z(n116) );
  XOR U88 ( .A(n117), .B(n118), .Z(n113) );
  AND U89 ( .A(n119), .B(n120), .Z(n118) );
  XNOR U90 ( .A(p_input[473]), .B(n117), .Z(n120) );
  XOR U91 ( .A(n121), .B(n122), .Z(n117) );
  AND U92 ( .A(n123), .B(n124), .Z(n122) );
  XNOR U93 ( .A(p_input[489]), .B(n121), .Z(n124) );
  XOR U94 ( .A(n125), .B(n126), .Z(n121) );
  AND U95 ( .A(n127), .B(n128), .Z(n126) );
  XNOR U96 ( .A(p_input[505]), .B(n125), .Z(n128) );
  XOR U97 ( .A(n129), .B(n130), .Z(n125) );
  AND U98 ( .A(n131), .B(n132), .Z(n130) );
  XNOR U99 ( .A(p_input[521]), .B(n129), .Z(n132) );
  XOR U100 ( .A(n133), .B(n134), .Z(n129) );
  AND U101 ( .A(n135), .B(n136), .Z(n134) );
  XNOR U102 ( .A(p_input[537]), .B(n133), .Z(n136) );
  XOR U103 ( .A(n137), .B(n138), .Z(n133) );
  AND U104 ( .A(n139), .B(n140), .Z(n138) );
  XNOR U105 ( .A(p_input[553]), .B(n137), .Z(n140) );
  XOR U106 ( .A(n141), .B(n142), .Z(n137) );
  AND U107 ( .A(n143), .B(n144), .Z(n142) );
  XNOR U108 ( .A(p_input[569]), .B(n141), .Z(n144) );
  XOR U109 ( .A(n145), .B(n146), .Z(n141) );
  AND U110 ( .A(n147), .B(n148), .Z(n146) );
  XNOR U111 ( .A(p_input[585]), .B(n145), .Z(n148) );
  XOR U112 ( .A(n149), .B(n150), .Z(n145) );
  AND U113 ( .A(n151), .B(n152), .Z(n150) );
  XNOR U114 ( .A(p_input[601]), .B(n149), .Z(n152) );
  XOR U115 ( .A(n153), .B(n154), .Z(n149) );
  AND U116 ( .A(n155), .B(n156), .Z(n154) );
  XNOR U117 ( .A(p_input[617]), .B(n153), .Z(n156) );
  XOR U118 ( .A(n157), .B(n158), .Z(n153) );
  AND U119 ( .A(n159), .B(n160), .Z(n158) );
  XNOR U120 ( .A(p_input[633]), .B(n157), .Z(n160) );
  XOR U121 ( .A(n161), .B(n162), .Z(n157) );
  AND U122 ( .A(n163), .B(n164), .Z(n162) );
  XNOR U123 ( .A(p_input[649]), .B(n161), .Z(n164) );
  XOR U124 ( .A(n165), .B(n166), .Z(n161) );
  AND U125 ( .A(n167), .B(n168), .Z(n166) );
  XNOR U126 ( .A(p_input[665]), .B(n165), .Z(n168) );
  XOR U127 ( .A(n169), .B(n170), .Z(n165) );
  AND U128 ( .A(n171), .B(n172), .Z(n170) );
  XNOR U129 ( .A(p_input[681]), .B(n169), .Z(n172) );
  XOR U130 ( .A(n173), .B(n174), .Z(n169) );
  AND U131 ( .A(n175), .B(n176), .Z(n174) );
  XNOR U132 ( .A(p_input[697]), .B(n173), .Z(n176) );
  XOR U133 ( .A(n177), .B(n178), .Z(n173) );
  AND U134 ( .A(n179), .B(n180), .Z(n178) );
  XNOR U135 ( .A(p_input[713]), .B(n177), .Z(n180) );
  XOR U136 ( .A(n181), .B(n182), .Z(n177) );
  AND U137 ( .A(n183), .B(n184), .Z(n182) );
  XNOR U138 ( .A(p_input[729]), .B(n181), .Z(n184) );
  XOR U139 ( .A(n185), .B(n186), .Z(n181) );
  AND U140 ( .A(n187), .B(n188), .Z(n186) );
  XNOR U141 ( .A(p_input[745]), .B(n185), .Z(n188) );
  XOR U142 ( .A(n189), .B(n190), .Z(n185) );
  AND U143 ( .A(n191), .B(n192), .Z(n190) );
  XNOR U144 ( .A(p_input[761]), .B(n189), .Z(n192) );
  XOR U145 ( .A(n193), .B(n194), .Z(n189) );
  AND U146 ( .A(n195), .B(n196), .Z(n194) );
  XNOR U147 ( .A(p_input[777]), .B(n193), .Z(n196) );
  XOR U148 ( .A(n197), .B(n198), .Z(n193) );
  AND U149 ( .A(n199), .B(n200), .Z(n198) );
  XNOR U150 ( .A(p_input[793]), .B(n197), .Z(n200) );
  XOR U151 ( .A(n201), .B(n202), .Z(n197) );
  AND U152 ( .A(n203), .B(n204), .Z(n202) );
  XNOR U153 ( .A(p_input[809]), .B(n201), .Z(n204) );
  XOR U154 ( .A(n205), .B(n206), .Z(n201) );
  AND U155 ( .A(n207), .B(n208), .Z(n206) );
  XNOR U156 ( .A(p_input[825]), .B(n205), .Z(n208) );
  XOR U157 ( .A(n209), .B(n210), .Z(n205) );
  AND U158 ( .A(n211), .B(n212), .Z(n210) );
  XNOR U159 ( .A(p_input[841]), .B(n209), .Z(n212) );
  XOR U160 ( .A(n213), .B(n214), .Z(n209) );
  AND U161 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U162 ( .A(p_input[857]), .B(n213), .Z(n216) );
  XOR U163 ( .A(n217), .B(n218), .Z(n213) );
  AND U164 ( .A(n219), .B(n220), .Z(n218) );
  XNOR U165 ( .A(p_input[873]), .B(n217), .Z(n220) );
  XOR U166 ( .A(n221), .B(n222), .Z(n217) );
  AND U167 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U168 ( .A(p_input[889]), .B(n221), .Z(n224) );
  XOR U169 ( .A(n225), .B(n226), .Z(n221) );
  AND U170 ( .A(n227), .B(n228), .Z(n226) );
  XNOR U171 ( .A(p_input[905]), .B(n225), .Z(n228) );
  XOR U172 ( .A(n229), .B(n230), .Z(n225) );
  AND U173 ( .A(n231), .B(n232), .Z(n230) );
  XNOR U174 ( .A(p_input[921]), .B(n229), .Z(n232) );
  XOR U175 ( .A(n233), .B(n234), .Z(n229) );
  AND U176 ( .A(n235), .B(n236), .Z(n234) );
  XNOR U177 ( .A(p_input[937]), .B(n233), .Z(n236) );
  XOR U178 ( .A(n237), .B(n238), .Z(n233) );
  AND U179 ( .A(n239), .B(n240), .Z(n238) );
  XNOR U180 ( .A(p_input[953]), .B(n237), .Z(n240) );
  XOR U181 ( .A(n241), .B(n242), .Z(n237) );
  AND U182 ( .A(n243), .B(n244), .Z(n242) );
  XNOR U183 ( .A(p_input[969]), .B(n241), .Z(n244) );
  XOR U184 ( .A(n245), .B(n246), .Z(n241) );
  AND U185 ( .A(n247), .B(n248), .Z(n246) );
  XNOR U186 ( .A(p_input[985]), .B(n245), .Z(n248) );
  XOR U187 ( .A(n249), .B(n250), .Z(n245) );
  AND U188 ( .A(n251), .B(n252), .Z(n250) );
  XNOR U189 ( .A(p_input[1001]), .B(n249), .Z(n252) );
  XOR U190 ( .A(n253), .B(n254), .Z(n249) );
  AND U191 ( .A(n255), .B(n256), .Z(n254) );
  XNOR U192 ( .A(p_input[1017]), .B(n253), .Z(n256) );
  XOR U193 ( .A(n257), .B(n258), .Z(n253) );
  AND U194 ( .A(n259), .B(n260), .Z(n258) );
  XNOR U195 ( .A(p_input[1033]), .B(n257), .Z(n260) );
  XOR U196 ( .A(n261), .B(n262), .Z(n257) );
  AND U197 ( .A(n263), .B(n264), .Z(n262) );
  XNOR U198 ( .A(p_input[1049]), .B(n261), .Z(n264) );
  XOR U199 ( .A(n265), .B(n266), .Z(n261) );
  AND U200 ( .A(n267), .B(n268), .Z(n266) );
  XNOR U201 ( .A(p_input[1065]), .B(n265), .Z(n268) );
  XOR U202 ( .A(n269), .B(n270), .Z(n265) );
  AND U203 ( .A(n271), .B(n272), .Z(n270) );
  XNOR U204 ( .A(p_input[1081]), .B(n269), .Z(n272) );
  XOR U205 ( .A(n273), .B(n274), .Z(n269) );
  AND U206 ( .A(n275), .B(n276), .Z(n274) );
  XNOR U207 ( .A(p_input[1097]), .B(n273), .Z(n276) );
  XOR U208 ( .A(n277), .B(n278), .Z(n273) );
  AND U209 ( .A(n279), .B(n280), .Z(n278) );
  XNOR U210 ( .A(p_input[1113]), .B(n277), .Z(n280) );
  XOR U211 ( .A(n281), .B(n282), .Z(n277) );
  AND U212 ( .A(n283), .B(n284), .Z(n282) );
  XNOR U213 ( .A(p_input[1129]), .B(n281), .Z(n284) );
  XOR U214 ( .A(n285), .B(n286), .Z(n281) );
  AND U215 ( .A(n287), .B(n288), .Z(n286) );
  XNOR U216 ( .A(p_input[1145]), .B(n285), .Z(n288) );
  XOR U217 ( .A(n289), .B(n290), .Z(n285) );
  AND U218 ( .A(n291), .B(n292), .Z(n290) );
  XNOR U219 ( .A(p_input[1161]), .B(n289), .Z(n292) );
  XOR U220 ( .A(n293), .B(n294), .Z(n289) );
  AND U221 ( .A(n295), .B(n296), .Z(n294) );
  XNOR U222 ( .A(p_input[1177]), .B(n293), .Z(n296) );
  XOR U223 ( .A(n297), .B(n298), .Z(n293) );
  AND U224 ( .A(n299), .B(n300), .Z(n298) );
  XNOR U225 ( .A(p_input[1193]), .B(n297), .Z(n300) );
  XOR U226 ( .A(n301), .B(n302), .Z(n297) );
  AND U227 ( .A(n303), .B(n304), .Z(n302) );
  XNOR U228 ( .A(p_input[1209]), .B(n301), .Z(n304) );
  XOR U229 ( .A(n305), .B(n306), .Z(n301) );
  AND U230 ( .A(n307), .B(n308), .Z(n306) );
  XNOR U231 ( .A(p_input[1225]), .B(n305), .Z(n308) );
  XOR U232 ( .A(n309), .B(n310), .Z(n305) );
  AND U233 ( .A(n311), .B(n312), .Z(n310) );
  XNOR U234 ( .A(p_input[1241]), .B(n309), .Z(n312) );
  XOR U235 ( .A(n313), .B(n314), .Z(n309) );
  AND U236 ( .A(n315), .B(n316), .Z(n314) );
  XNOR U237 ( .A(p_input[1257]), .B(n313), .Z(n316) );
  XOR U238 ( .A(n317), .B(n318), .Z(n313) );
  AND U239 ( .A(n319), .B(n320), .Z(n318) );
  XNOR U240 ( .A(p_input[1273]), .B(n317), .Z(n320) );
  XOR U241 ( .A(n321), .B(n322), .Z(n317) );
  AND U242 ( .A(n323), .B(n324), .Z(n322) );
  XNOR U243 ( .A(p_input[1289]), .B(n321), .Z(n324) );
  XOR U244 ( .A(n325), .B(n326), .Z(n321) );
  AND U245 ( .A(n327), .B(n328), .Z(n326) );
  XNOR U246 ( .A(p_input[1305]), .B(n325), .Z(n328) );
  XOR U247 ( .A(n329), .B(n330), .Z(n325) );
  AND U248 ( .A(n331), .B(n332), .Z(n330) );
  XNOR U249 ( .A(p_input[1321]), .B(n329), .Z(n332) );
  XOR U250 ( .A(n333), .B(n334), .Z(n329) );
  AND U251 ( .A(n335), .B(n336), .Z(n334) );
  XNOR U252 ( .A(p_input[1337]), .B(n333), .Z(n336) );
  XOR U253 ( .A(n337), .B(n338), .Z(n333) );
  AND U254 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U255 ( .A(p_input[1353]), .B(n337), .Z(n340) );
  XOR U256 ( .A(n341), .B(n342), .Z(n337) );
  AND U257 ( .A(n343), .B(n344), .Z(n342) );
  XNOR U258 ( .A(p_input[1369]), .B(n341), .Z(n344) );
  XOR U259 ( .A(n345), .B(n346), .Z(n341) );
  AND U260 ( .A(n347), .B(n348), .Z(n346) );
  XNOR U261 ( .A(p_input[1385]), .B(n345), .Z(n348) );
  XOR U262 ( .A(n349), .B(n350), .Z(n345) );
  AND U263 ( .A(n351), .B(n352), .Z(n350) );
  XNOR U264 ( .A(p_input[1401]), .B(n349), .Z(n352) );
  XOR U265 ( .A(n353), .B(n354), .Z(n349) );
  AND U266 ( .A(n355), .B(n356), .Z(n354) );
  XNOR U267 ( .A(p_input[1417]), .B(n353), .Z(n356) );
  XOR U268 ( .A(n357), .B(n358), .Z(n353) );
  AND U269 ( .A(n359), .B(n360), .Z(n358) );
  XNOR U270 ( .A(p_input[1433]), .B(n357), .Z(n360) );
  XOR U271 ( .A(n361), .B(n362), .Z(n357) );
  AND U272 ( .A(n363), .B(n364), .Z(n362) );
  XNOR U273 ( .A(p_input[1449]), .B(n361), .Z(n364) );
  XOR U274 ( .A(n365), .B(n366), .Z(n361) );
  AND U275 ( .A(n367), .B(n368), .Z(n366) );
  XNOR U276 ( .A(p_input[1465]), .B(n365), .Z(n368) );
  XOR U277 ( .A(n369), .B(n370), .Z(n365) );
  AND U278 ( .A(n371), .B(n372), .Z(n370) );
  XNOR U279 ( .A(p_input[1481]), .B(n369), .Z(n372) );
  XOR U280 ( .A(n373), .B(n374), .Z(n369) );
  AND U281 ( .A(n375), .B(n376), .Z(n374) );
  XNOR U282 ( .A(p_input[1497]), .B(n373), .Z(n376) );
  XOR U283 ( .A(n377), .B(n378), .Z(n373) );
  AND U284 ( .A(n379), .B(n380), .Z(n378) );
  XNOR U285 ( .A(p_input[1513]), .B(n377), .Z(n380) );
  XOR U286 ( .A(n381), .B(n382), .Z(n377) );
  AND U287 ( .A(n383), .B(n384), .Z(n382) );
  XNOR U288 ( .A(p_input[1529]), .B(n381), .Z(n384) );
  XOR U289 ( .A(n385), .B(n386), .Z(n381) );
  AND U290 ( .A(n387), .B(n388), .Z(n386) );
  XNOR U291 ( .A(p_input[1545]), .B(n385), .Z(n388) );
  XOR U292 ( .A(n389), .B(n390), .Z(n385) );
  AND U293 ( .A(n391), .B(n392), .Z(n390) );
  XNOR U294 ( .A(p_input[1561]), .B(n389), .Z(n392) );
  XOR U295 ( .A(n393), .B(n394), .Z(n389) );
  AND U296 ( .A(n395), .B(n396), .Z(n394) );
  XNOR U297 ( .A(p_input[1577]), .B(n393), .Z(n396) );
  XOR U298 ( .A(n397), .B(n398), .Z(n393) );
  AND U299 ( .A(n399), .B(n400), .Z(n398) );
  XNOR U300 ( .A(p_input[1593]), .B(n397), .Z(n400) );
  XOR U301 ( .A(n401), .B(n402), .Z(n397) );
  AND U302 ( .A(n403), .B(n404), .Z(n402) );
  XNOR U303 ( .A(p_input[1609]), .B(n401), .Z(n404) );
  XOR U304 ( .A(n405), .B(n406), .Z(n401) );
  AND U305 ( .A(n407), .B(n408), .Z(n406) );
  XNOR U306 ( .A(p_input[1625]), .B(n405), .Z(n408) );
  XOR U307 ( .A(n409), .B(n410), .Z(n405) );
  AND U308 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U309 ( .A(p_input[1641]), .B(n409), .Z(n412) );
  XOR U310 ( .A(n413), .B(n414), .Z(n409) );
  AND U311 ( .A(n415), .B(n416), .Z(n414) );
  XNOR U312 ( .A(p_input[1657]), .B(n413), .Z(n416) );
  XOR U313 ( .A(n417), .B(n418), .Z(n413) );
  AND U314 ( .A(n419), .B(n420), .Z(n418) );
  XNOR U315 ( .A(p_input[1673]), .B(n417), .Z(n420) );
  XOR U316 ( .A(n421), .B(n422), .Z(n417) );
  AND U317 ( .A(n423), .B(n424), .Z(n422) );
  XNOR U318 ( .A(p_input[1689]), .B(n421), .Z(n424) );
  XOR U319 ( .A(n425), .B(n426), .Z(n421) );
  AND U320 ( .A(n427), .B(n428), .Z(n426) );
  XNOR U321 ( .A(p_input[1705]), .B(n425), .Z(n428) );
  XOR U322 ( .A(n429), .B(n430), .Z(n425) );
  AND U323 ( .A(n431), .B(n432), .Z(n430) );
  XNOR U324 ( .A(p_input[1721]), .B(n429), .Z(n432) );
  XOR U325 ( .A(n433), .B(n434), .Z(n429) );
  AND U326 ( .A(n435), .B(n436), .Z(n434) );
  XNOR U327 ( .A(p_input[1737]), .B(n433), .Z(n436) );
  XOR U328 ( .A(n437), .B(n438), .Z(n433) );
  AND U329 ( .A(n439), .B(n440), .Z(n438) );
  XNOR U330 ( .A(p_input[1753]), .B(n437), .Z(n440) );
  XOR U331 ( .A(n441), .B(n442), .Z(n437) );
  AND U332 ( .A(n443), .B(n444), .Z(n442) );
  XNOR U333 ( .A(p_input[1769]), .B(n441), .Z(n444) );
  XOR U334 ( .A(n445), .B(n446), .Z(n441) );
  AND U335 ( .A(n447), .B(n448), .Z(n446) );
  XNOR U336 ( .A(p_input[1785]), .B(n445), .Z(n448) );
  XOR U337 ( .A(n449), .B(n450), .Z(n445) );
  AND U338 ( .A(n451), .B(n452), .Z(n450) );
  XNOR U339 ( .A(p_input[1801]), .B(n449), .Z(n452) );
  XOR U340 ( .A(n453), .B(n454), .Z(n449) );
  AND U341 ( .A(n455), .B(n456), .Z(n454) );
  XNOR U342 ( .A(p_input[1817]), .B(n453), .Z(n456) );
  XOR U343 ( .A(n457), .B(n458), .Z(n453) );
  AND U344 ( .A(n459), .B(n460), .Z(n458) );
  XNOR U345 ( .A(p_input[1833]), .B(n457), .Z(n460) );
  XOR U346 ( .A(n461), .B(n462), .Z(n457) );
  AND U347 ( .A(n463), .B(n464), .Z(n462) );
  XNOR U348 ( .A(p_input[1849]), .B(n461), .Z(n464) );
  XOR U349 ( .A(n465), .B(n466), .Z(n461) );
  AND U350 ( .A(n467), .B(n468), .Z(n466) );
  XNOR U351 ( .A(p_input[1865]), .B(n465), .Z(n468) );
  XOR U352 ( .A(n469), .B(n470), .Z(n465) );
  AND U353 ( .A(n471), .B(n472), .Z(n470) );
  XNOR U354 ( .A(p_input[1881]), .B(n469), .Z(n472) );
  XOR U355 ( .A(n473), .B(n474), .Z(n469) );
  AND U356 ( .A(n475), .B(n476), .Z(n474) );
  XNOR U357 ( .A(p_input[1897]), .B(n473), .Z(n476) );
  XOR U358 ( .A(n477), .B(n478), .Z(n473) );
  AND U359 ( .A(n479), .B(n480), .Z(n478) );
  XNOR U360 ( .A(p_input[1913]), .B(n477), .Z(n480) );
  XOR U361 ( .A(n481), .B(n482), .Z(n477) );
  AND U362 ( .A(n483), .B(n484), .Z(n482) );
  XNOR U363 ( .A(p_input[1929]), .B(n481), .Z(n484) );
  XOR U364 ( .A(n485), .B(n486), .Z(n481) );
  AND U365 ( .A(n487), .B(n488), .Z(n486) );
  XNOR U366 ( .A(p_input[1945]), .B(n485), .Z(n488) );
  XOR U367 ( .A(n489), .B(n490), .Z(n485) );
  AND U368 ( .A(n491), .B(n492), .Z(n490) );
  XNOR U369 ( .A(p_input[1961]), .B(n489), .Z(n492) );
  XOR U370 ( .A(n493), .B(n494), .Z(n489) );
  AND U371 ( .A(n495), .B(n496), .Z(n494) );
  XNOR U372 ( .A(p_input[1977]), .B(n493), .Z(n496) );
  XOR U373 ( .A(n497), .B(n498), .Z(n493) );
  AND U374 ( .A(n499), .B(n500), .Z(n498) );
  XNOR U375 ( .A(p_input[1993]), .B(n497), .Z(n500) );
  XNOR U376 ( .A(n501), .B(n502), .Z(n497) );
  AND U377 ( .A(n503), .B(n504), .Z(n502) );
  XOR U378 ( .A(p_input[2009]), .B(n501), .Z(n504) );
  XOR U379 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n505), .Z(n501) );
  AND U380 ( .A(n506), .B(n507), .Z(n505) );
  XOR U381 ( .A(p_input[2025]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n507) );
  XNOR U382 ( .A(n508), .B(n509), .Z(o[8]) );
  AND U383 ( .A(n3), .B(n510), .Z(n508) );
  XNOR U384 ( .A(p_input[8]), .B(n509), .Z(n510) );
  XOR U385 ( .A(n511), .B(n512), .Z(n509) );
  AND U386 ( .A(n7), .B(n513), .Z(n512) );
  XNOR U387 ( .A(p_input[24]), .B(n511), .Z(n513) );
  XOR U388 ( .A(n514), .B(n515), .Z(n511) );
  AND U389 ( .A(n11), .B(n516), .Z(n515) );
  XNOR U390 ( .A(p_input[40]), .B(n514), .Z(n516) );
  XOR U391 ( .A(n517), .B(n518), .Z(n514) );
  AND U392 ( .A(n15), .B(n519), .Z(n518) );
  XNOR U393 ( .A(p_input[56]), .B(n517), .Z(n519) );
  XOR U394 ( .A(n520), .B(n521), .Z(n517) );
  AND U395 ( .A(n19), .B(n522), .Z(n521) );
  XNOR U396 ( .A(p_input[72]), .B(n520), .Z(n522) );
  XOR U397 ( .A(n523), .B(n524), .Z(n520) );
  AND U398 ( .A(n23), .B(n525), .Z(n524) );
  XNOR U399 ( .A(p_input[88]), .B(n523), .Z(n525) );
  XOR U400 ( .A(n526), .B(n527), .Z(n523) );
  AND U401 ( .A(n27), .B(n528), .Z(n527) );
  XNOR U402 ( .A(p_input[104]), .B(n526), .Z(n528) );
  XOR U403 ( .A(n529), .B(n530), .Z(n526) );
  AND U404 ( .A(n31), .B(n531), .Z(n530) );
  XNOR U405 ( .A(p_input[120]), .B(n529), .Z(n531) );
  XOR U406 ( .A(n532), .B(n533), .Z(n529) );
  AND U407 ( .A(n35), .B(n534), .Z(n533) );
  XNOR U408 ( .A(p_input[136]), .B(n532), .Z(n534) );
  XOR U409 ( .A(n535), .B(n536), .Z(n532) );
  AND U410 ( .A(n39), .B(n537), .Z(n536) );
  XNOR U411 ( .A(p_input[152]), .B(n535), .Z(n537) );
  XOR U412 ( .A(n538), .B(n539), .Z(n535) );
  AND U413 ( .A(n43), .B(n540), .Z(n539) );
  XNOR U414 ( .A(p_input[168]), .B(n538), .Z(n540) );
  XOR U415 ( .A(n541), .B(n542), .Z(n538) );
  AND U416 ( .A(n47), .B(n543), .Z(n542) );
  XNOR U417 ( .A(p_input[184]), .B(n541), .Z(n543) );
  XOR U418 ( .A(n544), .B(n545), .Z(n541) );
  AND U419 ( .A(n51), .B(n546), .Z(n545) );
  XNOR U420 ( .A(p_input[200]), .B(n544), .Z(n546) );
  XOR U421 ( .A(n547), .B(n548), .Z(n544) );
  AND U422 ( .A(n55), .B(n549), .Z(n548) );
  XNOR U423 ( .A(p_input[216]), .B(n547), .Z(n549) );
  XOR U424 ( .A(n550), .B(n551), .Z(n547) );
  AND U425 ( .A(n59), .B(n552), .Z(n551) );
  XNOR U426 ( .A(p_input[232]), .B(n550), .Z(n552) );
  XOR U427 ( .A(n553), .B(n554), .Z(n550) );
  AND U428 ( .A(n63), .B(n555), .Z(n554) );
  XNOR U429 ( .A(p_input[248]), .B(n553), .Z(n555) );
  XOR U430 ( .A(n556), .B(n557), .Z(n553) );
  AND U431 ( .A(n67), .B(n558), .Z(n557) );
  XNOR U432 ( .A(p_input[264]), .B(n556), .Z(n558) );
  XOR U433 ( .A(n559), .B(n560), .Z(n556) );
  AND U434 ( .A(n71), .B(n561), .Z(n560) );
  XNOR U435 ( .A(p_input[280]), .B(n559), .Z(n561) );
  XOR U436 ( .A(n562), .B(n563), .Z(n559) );
  AND U437 ( .A(n75), .B(n564), .Z(n563) );
  XNOR U438 ( .A(p_input[296]), .B(n562), .Z(n564) );
  XOR U439 ( .A(n565), .B(n566), .Z(n562) );
  AND U440 ( .A(n79), .B(n567), .Z(n566) );
  XNOR U441 ( .A(p_input[312]), .B(n565), .Z(n567) );
  XOR U442 ( .A(n568), .B(n569), .Z(n565) );
  AND U443 ( .A(n83), .B(n570), .Z(n569) );
  XNOR U444 ( .A(p_input[328]), .B(n568), .Z(n570) );
  XOR U445 ( .A(n571), .B(n572), .Z(n568) );
  AND U446 ( .A(n87), .B(n573), .Z(n572) );
  XNOR U447 ( .A(p_input[344]), .B(n571), .Z(n573) );
  XOR U448 ( .A(n574), .B(n575), .Z(n571) );
  AND U449 ( .A(n91), .B(n576), .Z(n575) );
  XNOR U450 ( .A(p_input[360]), .B(n574), .Z(n576) );
  XOR U451 ( .A(n577), .B(n578), .Z(n574) );
  AND U452 ( .A(n95), .B(n579), .Z(n578) );
  XNOR U453 ( .A(p_input[376]), .B(n577), .Z(n579) );
  XOR U454 ( .A(n580), .B(n581), .Z(n577) );
  AND U455 ( .A(n99), .B(n582), .Z(n581) );
  XNOR U456 ( .A(p_input[392]), .B(n580), .Z(n582) );
  XOR U457 ( .A(n583), .B(n584), .Z(n580) );
  AND U458 ( .A(n103), .B(n585), .Z(n584) );
  XNOR U459 ( .A(p_input[408]), .B(n583), .Z(n585) );
  XOR U460 ( .A(n586), .B(n587), .Z(n583) );
  AND U461 ( .A(n107), .B(n588), .Z(n587) );
  XNOR U462 ( .A(p_input[424]), .B(n586), .Z(n588) );
  XOR U463 ( .A(n589), .B(n590), .Z(n586) );
  AND U464 ( .A(n111), .B(n591), .Z(n590) );
  XNOR U465 ( .A(p_input[440]), .B(n589), .Z(n591) );
  XOR U466 ( .A(n592), .B(n593), .Z(n589) );
  AND U467 ( .A(n115), .B(n594), .Z(n593) );
  XNOR U468 ( .A(p_input[456]), .B(n592), .Z(n594) );
  XOR U469 ( .A(n595), .B(n596), .Z(n592) );
  AND U470 ( .A(n119), .B(n597), .Z(n596) );
  XNOR U471 ( .A(p_input[472]), .B(n595), .Z(n597) );
  XOR U472 ( .A(n598), .B(n599), .Z(n595) );
  AND U473 ( .A(n123), .B(n600), .Z(n599) );
  XNOR U474 ( .A(p_input[488]), .B(n598), .Z(n600) );
  XOR U475 ( .A(n601), .B(n602), .Z(n598) );
  AND U476 ( .A(n127), .B(n603), .Z(n602) );
  XNOR U477 ( .A(p_input[504]), .B(n601), .Z(n603) );
  XOR U478 ( .A(n604), .B(n605), .Z(n601) );
  AND U479 ( .A(n131), .B(n606), .Z(n605) );
  XNOR U480 ( .A(p_input[520]), .B(n604), .Z(n606) );
  XOR U481 ( .A(n607), .B(n608), .Z(n604) );
  AND U482 ( .A(n135), .B(n609), .Z(n608) );
  XNOR U483 ( .A(p_input[536]), .B(n607), .Z(n609) );
  XOR U484 ( .A(n610), .B(n611), .Z(n607) );
  AND U485 ( .A(n139), .B(n612), .Z(n611) );
  XNOR U486 ( .A(p_input[552]), .B(n610), .Z(n612) );
  XOR U487 ( .A(n613), .B(n614), .Z(n610) );
  AND U488 ( .A(n143), .B(n615), .Z(n614) );
  XNOR U489 ( .A(p_input[568]), .B(n613), .Z(n615) );
  XOR U490 ( .A(n616), .B(n617), .Z(n613) );
  AND U491 ( .A(n147), .B(n618), .Z(n617) );
  XNOR U492 ( .A(p_input[584]), .B(n616), .Z(n618) );
  XOR U493 ( .A(n619), .B(n620), .Z(n616) );
  AND U494 ( .A(n151), .B(n621), .Z(n620) );
  XNOR U495 ( .A(p_input[600]), .B(n619), .Z(n621) );
  XOR U496 ( .A(n622), .B(n623), .Z(n619) );
  AND U497 ( .A(n155), .B(n624), .Z(n623) );
  XNOR U498 ( .A(p_input[616]), .B(n622), .Z(n624) );
  XOR U499 ( .A(n625), .B(n626), .Z(n622) );
  AND U500 ( .A(n159), .B(n627), .Z(n626) );
  XNOR U501 ( .A(p_input[632]), .B(n625), .Z(n627) );
  XOR U502 ( .A(n628), .B(n629), .Z(n625) );
  AND U503 ( .A(n163), .B(n630), .Z(n629) );
  XNOR U504 ( .A(p_input[648]), .B(n628), .Z(n630) );
  XOR U505 ( .A(n631), .B(n632), .Z(n628) );
  AND U506 ( .A(n167), .B(n633), .Z(n632) );
  XNOR U507 ( .A(p_input[664]), .B(n631), .Z(n633) );
  XOR U508 ( .A(n634), .B(n635), .Z(n631) );
  AND U509 ( .A(n171), .B(n636), .Z(n635) );
  XNOR U510 ( .A(p_input[680]), .B(n634), .Z(n636) );
  XOR U511 ( .A(n637), .B(n638), .Z(n634) );
  AND U512 ( .A(n175), .B(n639), .Z(n638) );
  XNOR U513 ( .A(p_input[696]), .B(n637), .Z(n639) );
  XOR U514 ( .A(n640), .B(n641), .Z(n637) );
  AND U515 ( .A(n179), .B(n642), .Z(n641) );
  XNOR U516 ( .A(p_input[712]), .B(n640), .Z(n642) );
  XOR U517 ( .A(n643), .B(n644), .Z(n640) );
  AND U518 ( .A(n183), .B(n645), .Z(n644) );
  XNOR U519 ( .A(p_input[728]), .B(n643), .Z(n645) );
  XOR U520 ( .A(n646), .B(n647), .Z(n643) );
  AND U521 ( .A(n187), .B(n648), .Z(n647) );
  XNOR U522 ( .A(p_input[744]), .B(n646), .Z(n648) );
  XOR U523 ( .A(n649), .B(n650), .Z(n646) );
  AND U524 ( .A(n191), .B(n651), .Z(n650) );
  XNOR U525 ( .A(p_input[760]), .B(n649), .Z(n651) );
  XOR U526 ( .A(n652), .B(n653), .Z(n649) );
  AND U527 ( .A(n195), .B(n654), .Z(n653) );
  XNOR U528 ( .A(p_input[776]), .B(n652), .Z(n654) );
  XOR U529 ( .A(n655), .B(n656), .Z(n652) );
  AND U530 ( .A(n199), .B(n657), .Z(n656) );
  XNOR U531 ( .A(p_input[792]), .B(n655), .Z(n657) );
  XOR U532 ( .A(n658), .B(n659), .Z(n655) );
  AND U533 ( .A(n203), .B(n660), .Z(n659) );
  XNOR U534 ( .A(p_input[808]), .B(n658), .Z(n660) );
  XOR U535 ( .A(n661), .B(n662), .Z(n658) );
  AND U536 ( .A(n207), .B(n663), .Z(n662) );
  XNOR U537 ( .A(p_input[824]), .B(n661), .Z(n663) );
  XOR U538 ( .A(n664), .B(n665), .Z(n661) );
  AND U539 ( .A(n211), .B(n666), .Z(n665) );
  XNOR U540 ( .A(p_input[840]), .B(n664), .Z(n666) );
  XOR U541 ( .A(n667), .B(n668), .Z(n664) );
  AND U542 ( .A(n215), .B(n669), .Z(n668) );
  XNOR U543 ( .A(p_input[856]), .B(n667), .Z(n669) );
  XOR U544 ( .A(n670), .B(n671), .Z(n667) );
  AND U545 ( .A(n219), .B(n672), .Z(n671) );
  XNOR U546 ( .A(p_input[872]), .B(n670), .Z(n672) );
  XOR U547 ( .A(n673), .B(n674), .Z(n670) );
  AND U548 ( .A(n223), .B(n675), .Z(n674) );
  XNOR U549 ( .A(p_input[888]), .B(n673), .Z(n675) );
  XOR U550 ( .A(n676), .B(n677), .Z(n673) );
  AND U551 ( .A(n227), .B(n678), .Z(n677) );
  XNOR U552 ( .A(p_input[904]), .B(n676), .Z(n678) );
  XOR U553 ( .A(n679), .B(n680), .Z(n676) );
  AND U554 ( .A(n231), .B(n681), .Z(n680) );
  XNOR U555 ( .A(p_input[920]), .B(n679), .Z(n681) );
  XOR U556 ( .A(n682), .B(n683), .Z(n679) );
  AND U557 ( .A(n235), .B(n684), .Z(n683) );
  XNOR U558 ( .A(p_input[936]), .B(n682), .Z(n684) );
  XOR U559 ( .A(n685), .B(n686), .Z(n682) );
  AND U560 ( .A(n239), .B(n687), .Z(n686) );
  XNOR U561 ( .A(p_input[952]), .B(n685), .Z(n687) );
  XOR U562 ( .A(n688), .B(n689), .Z(n685) );
  AND U563 ( .A(n243), .B(n690), .Z(n689) );
  XNOR U564 ( .A(p_input[968]), .B(n688), .Z(n690) );
  XOR U565 ( .A(n691), .B(n692), .Z(n688) );
  AND U566 ( .A(n247), .B(n693), .Z(n692) );
  XNOR U567 ( .A(p_input[984]), .B(n691), .Z(n693) );
  XOR U568 ( .A(n694), .B(n695), .Z(n691) );
  AND U569 ( .A(n251), .B(n696), .Z(n695) );
  XNOR U570 ( .A(p_input[1000]), .B(n694), .Z(n696) );
  XOR U571 ( .A(n697), .B(n698), .Z(n694) );
  AND U572 ( .A(n255), .B(n699), .Z(n698) );
  XNOR U573 ( .A(p_input[1016]), .B(n697), .Z(n699) );
  XOR U574 ( .A(n700), .B(n701), .Z(n697) );
  AND U575 ( .A(n259), .B(n702), .Z(n701) );
  XNOR U576 ( .A(p_input[1032]), .B(n700), .Z(n702) );
  XOR U577 ( .A(n703), .B(n704), .Z(n700) );
  AND U578 ( .A(n263), .B(n705), .Z(n704) );
  XNOR U579 ( .A(p_input[1048]), .B(n703), .Z(n705) );
  XOR U580 ( .A(n706), .B(n707), .Z(n703) );
  AND U581 ( .A(n267), .B(n708), .Z(n707) );
  XNOR U582 ( .A(p_input[1064]), .B(n706), .Z(n708) );
  XOR U583 ( .A(n709), .B(n710), .Z(n706) );
  AND U584 ( .A(n271), .B(n711), .Z(n710) );
  XNOR U585 ( .A(p_input[1080]), .B(n709), .Z(n711) );
  XOR U586 ( .A(n712), .B(n713), .Z(n709) );
  AND U587 ( .A(n275), .B(n714), .Z(n713) );
  XNOR U588 ( .A(p_input[1096]), .B(n712), .Z(n714) );
  XOR U589 ( .A(n715), .B(n716), .Z(n712) );
  AND U590 ( .A(n279), .B(n717), .Z(n716) );
  XNOR U591 ( .A(p_input[1112]), .B(n715), .Z(n717) );
  XOR U592 ( .A(n718), .B(n719), .Z(n715) );
  AND U593 ( .A(n283), .B(n720), .Z(n719) );
  XNOR U594 ( .A(p_input[1128]), .B(n718), .Z(n720) );
  XOR U595 ( .A(n721), .B(n722), .Z(n718) );
  AND U596 ( .A(n287), .B(n723), .Z(n722) );
  XNOR U597 ( .A(p_input[1144]), .B(n721), .Z(n723) );
  XOR U598 ( .A(n724), .B(n725), .Z(n721) );
  AND U599 ( .A(n291), .B(n726), .Z(n725) );
  XNOR U600 ( .A(p_input[1160]), .B(n724), .Z(n726) );
  XOR U601 ( .A(n727), .B(n728), .Z(n724) );
  AND U602 ( .A(n295), .B(n729), .Z(n728) );
  XNOR U603 ( .A(p_input[1176]), .B(n727), .Z(n729) );
  XOR U604 ( .A(n730), .B(n731), .Z(n727) );
  AND U605 ( .A(n299), .B(n732), .Z(n731) );
  XNOR U606 ( .A(p_input[1192]), .B(n730), .Z(n732) );
  XOR U607 ( .A(n733), .B(n734), .Z(n730) );
  AND U608 ( .A(n303), .B(n735), .Z(n734) );
  XNOR U609 ( .A(p_input[1208]), .B(n733), .Z(n735) );
  XOR U610 ( .A(n736), .B(n737), .Z(n733) );
  AND U611 ( .A(n307), .B(n738), .Z(n737) );
  XNOR U612 ( .A(p_input[1224]), .B(n736), .Z(n738) );
  XOR U613 ( .A(n739), .B(n740), .Z(n736) );
  AND U614 ( .A(n311), .B(n741), .Z(n740) );
  XNOR U615 ( .A(p_input[1240]), .B(n739), .Z(n741) );
  XOR U616 ( .A(n742), .B(n743), .Z(n739) );
  AND U617 ( .A(n315), .B(n744), .Z(n743) );
  XNOR U618 ( .A(p_input[1256]), .B(n742), .Z(n744) );
  XOR U619 ( .A(n745), .B(n746), .Z(n742) );
  AND U620 ( .A(n319), .B(n747), .Z(n746) );
  XNOR U621 ( .A(p_input[1272]), .B(n745), .Z(n747) );
  XOR U622 ( .A(n748), .B(n749), .Z(n745) );
  AND U623 ( .A(n323), .B(n750), .Z(n749) );
  XNOR U624 ( .A(p_input[1288]), .B(n748), .Z(n750) );
  XOR U625 ( .A(n751), .B(n752), .Z(n748) );
  AND U626 ( .A(n327), .B(n753), .Z(n752) );
  XNOR U627 ( .A(p_input[1304]), .B(n751), .Z(n753) );
  XOR U628 ( .A(n754), .B(n755), .Z(n751) );
  AND U629 ( .A(n331), .B(n756), .Z(n755) );
  XNOR U630 ( .A(p_input[1320]), .B(n754), .Z(n756) );
  XOR U631 ( .A(n757), .B(n758), .Z(n754) );
  AND U632 ( .A(n335), .B(n759), .Z(n758) );
  XNOR U633 ( .A(p_input[1336]), .B(n757), .Z(n759) );
  XOR U634 ( .A(n760), .B(n761), .Z(n757) );
  AND U635 ( .A(n339), .B(n762), .Z(n761) );
  XNOR U636 ( .A(p_input[1352]), .B(n760), .Z(n762) );
  XOR U637 ( .A(n763), .B(n764), .Z(n760) );
  AND U638 ( .A(n343), .B(n765), .Z(n764) );
  XNOR U639 ( .A(p_input[1368]), .B(n763), .Z(n765) );
  XOR U640 ( .A(n766), .B(n767), .Z(n763) );
  AND U641 ( .A(n347), .B(n768), .Z(n767) );
  XNOR U642 ( .A(p_input[1384]), .B(n766), .Z(n768) );
  XOR U643 ( .A(n769), .B(n770), .Z(n766) );
  AND U644 ( .A(n351), .B(n771), .Z(n770) );
  XNOR U645 ( .A(p_input[1400]), .B(n769), .Z(n771) );
  XOR U646 ( .A(n772), .B(n773), .Z(n769) );
  AND U647 ( .A(n355), .B(n774), .Z(n773) );
  XNOR U648 ( .A(p_input[1416]), .B(n772), .Z(n774) );
  XOR U649 ( .A(n775), .B(n776), .Z(n772) );
  AND U650 ( .A(n359), .B(n777), .Z(n776) );
  XNOR U651 ( .A(p_input[1432]), .B(n775), .Z(n777) );
  XOR U652 ( .A(n778), .B(n779), .Z(n775) );
  AND U653 ( .A(n363), .B(n780), .Z(n779) );
  XNOR U654 ( .A(p_input[1448]), .B(n778), .Z(n780) );
  XOR U655 ( .A(n781), .B(n782), .Z(n778) );
  AND U656 ( .A(n367), .B(n783), .Z(n782) );
  XNOR U657 ( .A(p_input[1464]), .B(n781), .Z(n783) );
  XOR U658 ( .A(n784), .B(n785), .Z(n781) );
  AND U659 ( .A(n371), .B(n786), .Z(n785) );
  XNOR U660 ( .A(p_input[1480]), .B(n784), .Z(n786) );
  XOR U661 ( .A(n787), .B(n788), .Z(n784) );
  AND U662 ( .A(n375), .B(n789), .Z(n788) );
  XNOR U663 ( .A(p_input[1496]), .B(n787), .Z(n789) );
  XOR U664 ( .A(n790), .B(n791), .Z(n787) );
  AND U665 ( .A(n379), .B(n792), .Z(n791) );
  XNOR U666 ( .A(p_input[1512]), .B(n790), .Z(n792) );
  XOR U667 ( .A(n793), .B(n794), .Z(n790) );
  AND U668 ( .A(n383), .B(n795), .Z(n794) );
  XNOR U669 ( .A(p_input[1528]), .B(n793), .Z(n795) );
  XOR U670 ( .A(n796), .B(n797), .Z(n793) );
  AND U671 ( .A(n387), .B(n798), .Z(n797) );
  XNOR U672 ( .A(p_input[1544]), .B(n796), .Z(n798) );
  XOR U673 ( .A(n799), .B(n800), .Z(n796) );
  AND U674 ( .A(n391), .B(n801), .Z(n800) );
  XNOR U675 ( .A(p_input[1560]), .B(n799), .Z(n801) );
  XOR U676 ( .A(n802), .B(n803), .Z(n799) );
  AND U677 ( .A(n395), .B(n804), .Z(n803) );
  XNOR U678 ( .A(p_input[1576]), .B(n802), .Z(n804) );
  XOR U679 ( .A(n805), .B(n806), .Z(n802) );
  AND U680 ( .A(n399), .B(n807), .Z(n806) );
  XNOR U681 ( .A(p_input[1592]), .B(n805), .Z(n807) );
  XOR U682 ( .A(n808), .B(n809), .Z(n805) );
  AND U683 ( .A(n403), .B(n810), .Z(n809) );
  XNOR U684 ( .A(p_input[1608]), .B(n808), .Z(n810) );
  XOR U685 ( .A(n811), .B(n812), .Z(n808) );
  AND U686 ( .A(n407), .B(n813), .Z(n812) );
  XNOR U687 ( .A(p_input[1624]), .B(n811), .Z(n813) );
  XOR U688 ( .A(n814), .B(n815), .Z(n811) );
  AND U689 ( .A(n411), .B(n816), .Z(n815) );
  XNOR U690 ( .A(p_input[1640]), .B(n814), .Z(n816) );
  XOR U691 ( .A(n817), .B(n818), .Z(n814) );
  AND U692 ( .A(n415), .B(n819), .Z(n818) );
  XNOR U693 ( .A(p_input[1656]), .B(n817), .Z(n819) );
  XOR U694 ( .A(n820), .B(n821), .Z(n817) );
  AND U695 ( .A(n419), .B(n822), .Z(n821) );
  XNOR U696 ( .A(p_input[1672]), .B(n820), .Z(n822) );
  XOR U697 ( .A(n823), .B(n824), .Z(n820) );
  AND U698 ( .A(n423), .B(n825), .Z(n824) );
  XNOR U699 ( .A(p_input[1688]), .B(n823), .Z(n825) );
  XOR U700 ( .A(n826), .B(n827), .Z(n823) );
  AND U701 ( .A(n427), .B(n828), .Z(n827) );
  XNOR U702 ( .A(p_input[1704]), .B(n826), .Z(n828) );
  XOR U703 ( .A(n829), .B(n830), .Z(n826) );
  AND U704 ( .A(n431), .B(n831), .Z(n830) );
  XNOR U705 ( .A(p_input[1720]), .B(n829), .Z(n831) );
  XOR U706 ( .A(n832), .B(n833), .Z(n829) );
  AND U707 ( .A(n435), .B(n834), .Z(n833) );
  XNOR U708 ( .A(p_input[1736]), .B(n832), .Z(n834) );
  XOR U709 ( .A(n835), .B(n836), .Z(n832) );
  AND U710 ( .A(n439), .B(n837), .Z(n836) );
  XNOR U711 ( .A(p_input[1752]), .B(n835), .Z(n837) );
  XOR U712 ( .A(n838), .B(n839), .Z(n835) );
  AND U713 ( .A(n443), .B(n840), .Z(n839) );
  XNOR U714 ( .A(p_input[1768]), .B(n838), .Z(n840) );
  XOR U715 ( .A(n841), .B(n842), .Z(n838) );
  AND U716 ( .A(n447), .B(n843), .Z(n842) );
  XNOR U717 ( .A(p_input[1784]), .B(n841), .Z(n843) );
  XOR U718 ( .A(n844), .B(n845), .Z(n841) );
  AND U719 ( .A(n451), .B(n846), .Z(n845) );
  XNOR U720 ( .A(p_input[1800]), .B(n844), .Z(n846) );
  XOR U721 ( .A(n847), .B(n848), .Z(n844) );
  AND U722 ( .A(n455), .B(n849), .Z(n848) );
  XNOR U723 ( .A(p_input[1816]), .B(n847), .Z(n849) );
  XOR U724 ( .A(n850), .B(n851), .Z(n847) );
  AND U725 ( .A(n459), .B(n852), .Z(n851) );
  XNOR U726 ( .A(p_input[1832]), .B(n850), .Z(n852) );
  XOR U727 ( .A(n853), .B(n854), .Z(n850) );
  AND U728 ( .A(n463), .B(n855), .Z(n854) );
  XNOR U729 ( .A(p_input[1848]), .B(n853), .Z(n855) );
  XOR U730 ( .A(n856), .B(n857), .Z(n853) );
  AND U731 ( .A(n467), .B(n858), .Z(n857) );
  XNOR U732 ( .A(p_input[1864]), .B(n856), .Z(n858) );
  XOR U733 ( .A(n859), .B(n860), .Z(n856) );
  AND U734 ( .A(n471), .B(n861), .Z(n860) );
  XNOR U735 ( .A(p_input[1880]), .B(n859), .Z(n861) );
  XOR U736 ( .A(n862), .B(n863), .Z(n859) );
  AND U737 ( .A(n475), .B(n864), .Z(n863) );
  XNOR U738 ( .A(p_input[1896]), .B(n862), .Z(n864) );
  XOR U739 ( .A(n865), .B(n866), .Z(n862) );
  AND U740 ( .A(n479), .B(n867), .Z(n866) );
  XNOR U741 ( .A(p_input[1912]), .B(n865), .Z(n867) );
  XOR U742 ( .A(n868), .B(n869), .Z(n865) );
  AND U743 ( .A(n483), .B(n870), .Z(n869) );
  XNOR U744 ( .A(p_input[1928]), .B(n868), .Z(n870) );
  XOR U745 ( .A(n871), .B(n872), .Z(n868) );
  AND U746 ( .A(n487), .B(n873), .Z(n872) );
  XNOR U747 ( .A(p_input[1944]), .B(n871), .Z(n873) );
  XOR U748 ( .A(n874), .B(n875), .Z(n871) );
  AND U749 ( .A(n491), .B(n876), .Z(n875) );
  XNOR U750 ( .A(p_input[1960]), .B(n874), .Z(n876) );
  XOR U751 ( .A(n877), .B(n878), .Z(n874) );
  AND U752 ( .A(n495), .B(n879), .Z(n878) );
  XNOR U753 ( .A(p_input[1976]), .B(n877), .Z(n879) );
  XOR U754 ( .A(n880), .B(n881), .Z(n877) );
  AND U755 ( .A(n499), .B(n882), .Z(n881) );
  XNOR U756 ( .A(p_input[1992]), .B(n880), .Z(n882) );
  XNOR U757 ( .A(n883), .B(n884), .Z(n880) );
  AND U758 ( .A(n503), .B(n885), .Z(n884) );
  XOR U759 ( .A(p_input[2008]), .B(n883), .Z(n885) );
  XOR U760 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n886), .Z(n883) );
  AND U761 ( .A(n506), .B(n887), .Z(n886) );
  XOR U762 ( .A(p_input[2024]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n887) );
  XNOR U763 ( .A(n888), .B(n889), .Z(o[7]) );
  AND U764 ( .A(n3), .B(n890), .Z(n888) );
  XNOR U765 ( .A(p_input[7]), .B(n889), .Z(n890) );
  XOR U766 ( .A(n891), .B(n892), .Z(n889) );
  AND U767 ( .A(n7), .B(n893), .Z(n892) );
  XNOR U768 ( .A(p_input[23]), .B(n891), .Z(n893) );
  XOR U769 ( .A(n894), .B(n895), .Z(n891) );
  AND U770 ( .A(n11), .B(n896), .Z(n895) );
  XNOR U771 ( .A(p_input[39]), .B(n894), .Z(n896) );
  XOR U772 ( .A(n897), .B(n898), .Z(n894) );
  AND U773 ( .A(n15), .B(n899), .Z(n898) );
  XNOR U774 ( .A(p_input[55]), .B(n897), .Z(n899) );
  XOR U775 ( .A(n900), .B(n901), .Z(n897) );
  AND U776 ( .A(n19), .B(n902), .Z(n901) );
  XNOR U777 ( .A(p_input[71]), .B(n900), .Z(n902) );
  XOR U778 ( .A(n903), .B(n904), .Z(n900) );
  AND U779 ( .A(n23), .B(n905), .Z(n904) );
  XNOR U780 ( .A(p_input[87]), .B(n903), .Z(n905) );
  XOR U781 ( .A(n906), .B(n907), .Z(n903) );
  AND U782 ( .A(n27), .B(n908), .Z(n907) );
  XNOR U783 ( .A(p_input[103]), .B(n906), .Z(n908) );
  XOR U784 ( .A(n909), .B(n910), .Z(n906) );
  AND U785 ( .A(n31), .B(n911), .Z(n910) );
  XNOR U786 ( .A(p_input[119]), .B(n909), .Z(n911) );
  XOR U787 ( .A(n912), .B(n913), .Z(n909) );
  AND U788 ( .A(n35), .B(n914), .Z(n913) );
  XNOR U789 ( .A(p_input[135]), .B(n912), .Z(n914) );
  XOR U790 ( .A(n915), .B(n916), .Z(n912) );
  AND U791 ( .A(n39), .B(n917), .Z(n916) );
  XNOR U792 ( .A(p_input[151]), .B(n915), .Z(n917) );
  XOR U793 ( .A(n918), .B(n919), .Z(n915) );
  AND U794 ( .A(n43), .B(n920), .Z(n919) );
  XNOR U795 ( .A(p_input[167]), .B(n918), .Z(n920) );
  XOR U796 ( .A(n921), .B(n922), .Z(n918) );
  AND U797 ( .A(n47), .B(n923), .Z(n922) );
  XNOR U798 ( .A(p_input[183]), .B(n921), .Z(n923) );
  XOR U799 ( .A(n924), .B(n925), .Z(n921) );
  AND U800 ( .A(n51), .B(n926), .Z(n925) );
  XNOR U801 ( .A(p_input[199]), .B(n924), .Z(n926) );
  XOR U802 ( .A(n927), .B(n928), .Z(n924) );
  AND U803 ( .A(n55), .B(n929), .Z(n928) );
  XNOR U804 ( .A(p_input[215]), .B(n927), .Z(n929) );
  XOR U805 ( .A(n930), .B(n931), .Z(n927) );
  AND U806 ( .A(n59), .B(n932), .Z(n931) );
  XNOR U807 ( .A(p_input[231]), .B(n930), .Z(n932) );
  XOR U808 ( .A(n933), .B(n934), .Z(n930) );
  AND U809 ( .A(n63), .B(n935), .Z(n934) );
  XNOR U810 ( .A(p_input[247]), .B(n933), .Z(n935) );
  XOR U811 ( .A(n936), .B(n937), .Z(n933) );
  AND U812 ( .A(n67), .B(n938), .Z(n937) );
  XNOR U813 ( .A(p_input[263]), .B(n936), .Z(n938) );
  XOR U814 ( .A(n939), .B(n940), .Z(n936) );
  AND U815 ( .A(n71), .B(n941), .Z(n940) );
  XNOR U816 ( .A(p_input[279]), .B(n939), .Z(n941) );
  XOR U817 ( .A(n942), .B(n943), .Z(n939) );
  AND U818 ( .A(n75), .B(n944), .Z(n943) );
  XNOR U819 ( .A(p_input[295]), .B(n942), .Z(n944) );
  XOR U820 ( .A(n945), .B(n946), .Z(n942) );
  AND U821 ( .A(n79), .B(n947), .Z(n946) );
  XNOR U822 ( .A(p_input[311]), .B(n945), .Z(n947) );
  XOR U823 ( .A(n948), .B(n949), .Z(n945) );
  AND U824 ( .A(n83), .B(n950), .Z(n949) );
  XNOR U825 ( .A(p_input[327]), .B(n948), .Z(n950) );
  XOR U826 ( .A(n951), .B(n952), .Z(n948) );
  AND U827 ( .A(n87), .B(n953), .Z(n952) );
  XNOR U828 ( .A(p_input[343]), .B(n951), .Z(n953) );
  XOR U829 ( .A(n954), .B(n955), .Z(n951) );
  AND U830 ( .A(n91), .B(n956), .Z(n955) );
  XNOR U831 ( .A(p_input[359]), .B(n954), .Z(n956) );
  XOR U832 ( .A(n957), .B(n958), .Z(n954) );
  AND U833 ( .A(n95), .B(n959), .Z(n958) );
  XNOR U834 ( .A(p_input[375]), .B(n957), .Z(n959) );
  XOR U835 ( .A(n960), .B(n961), .Z(n957) );
  AND U836 ( .A(n99), .B(n962), .Z(n961) );
  XNOR U837 ( .A(p_input[391]), .B(n960), .Z(n962) );
  XOR U838 ( .A(n963), .B(n964), .Z(n960) );
  AND U839 ( .A(n103), .B(n965), .Z(n964) );
  XNOR U840 ( .A(p_input[407]), .B(n963), .Z(n965) );
  XOR U841 ( .A(n966), .B(n967), .Z(n963) );
  AND U842 ( .A(n107), .B(n968), .Z(n967) );
  XNOR U843 ( .A(p_input[423]), .B(n966), .Z(n968) );
  XOR U844 ( .A(n969), .B(n970), .Z(n966) );
  AND U845 ( .A(n111), .B(n971), .Z(n970) );
  XNOR U846 ( .A(p_input[439]), .B(n969), .Z(n971) );
  XOR U847 ( .A(n972), .B(n973), .Z(n969) );
  AND U848 ( .A(n115), .B(n974), .Z(n973) );
  XNOR U849 ( .A(p_input[455]), .B(n972), .Z(n974) );
  XOR U850 ( .A(n975), .B(n976), .Z(n972) );
  AND U851 ( .A(n119), .B(n977), .Z(n976) );
  XNOR U852 ( .A(p_input[471]), .B(n975), .Z(n977) );
  XOR U853 ( .A(n978), .B(n979), .Z(n975) );
  AND U854 ( .A(n123), .B(n980), .Z(n979) );
  XNOR U855 ( .A(p_input[487]), .B(n978), .Z(n980) );
  XOR U856 ( .A(n981), .B(n982), .Z(n978) );
  AND U857 ( .A(n127), .B(n983), .Z(n982) );
  XNOR U858 ( .A(p_input[503]), .B(n981), .Z(n983) );
  XOR U859 ( .A(n984), .B(n985), .Z(n981) );
  AND U860 ( .A(n131), .B(n986), .Z(n985) );
  XNOR U861 ( .A(p_input[519]), .B(n984), .Z(n986) );
  XOR U862 ( .A(n987), .B(n988), .Z(n984) );
  AND U863 ( .A(n135), .B(n989), .Z(n988) );
  XNOR U864 ( .A(p_input[535]), .B(n987), .Z(n989) );
  XOR U865 ( .A(n990), .B(n991), .Z(n987) );
  AND U866 ( .A(n139), .B(n992), .Z(n991) );
  XNOR U867 ( .A(p_input[551]), .B(n990), .Z(n992) );
  XOR U868 ( .A(n993), .B(n994), .Z(n990) );
  AND U869 ( .A(n143), .B(n995), .Z(n994) );
  XNOR U870 ( .A(p_input[567]), .B(n993), .Z(n995) );
  XOR U871 ( .A(n996), .B(n997), .Z(n993) );
  AND U872 ( .A(n147), .B(n998), .Z(n997) );
  XNOR U873 ( .A(p_input[583]), .B(n996), .Z(n998) );
  XOR U874 ( .A(n999), .B(n1000), .Z(n996) );
  AND U875 ( .A(n151), .B(n1001), .Z(n1000) );
  XNOR U876 ( .A(p_input[599]), .B(n999), .Z(n1001) );
  XOR U877 ( .A(n1002), .B(n1003), .Z(n999) );
  AND U878 ( .A(n155), .B(n1004), .Z(n1003) );
  XNOR U879 ( .A(p_input[615]), .B(n1002), .Z(n1004) );
  XOR U880 ( .A(n1005), .B(n1006), .Z(n1002) );
  AND U881 ( .A(n159), .B(n1007), .Z(n1006) );
  XNOR U882 ( .A(p_input[631]), .B(n1005), .Z(n1007) );
  XOR U883 ( .A(n1008), .B(n1009), .Z(n1005) );
  AND U884 ( .A(n163), .B(n1010), .Z(n1009) );
  XNOR U885 ( .A(p_input[647]), .B(n1008), .Z(n1010) );
  XOR U886 ( .A(n1011), .B(n1012), .Z(n1008) );
  AND U887 ( .A(n167), .B(n1013), .Z(n1012) );
  XNOR U888 ( .A(p_input[663]), .B(n1011), .Z(n1013) );
  XOR U889 ( .A(n1014), .B(n1015), .Z(n1011) );
  AND U890 ( .A(n171), .B(n1016), .Z(n1015) );
  XNOR U891 ( .A(p_input[679]), .B(n1014), .Z(n1016) );
  XOR U892 ( .A(n1017), .B(n1018), .Z(n1014) );
  AND U893 ( .A(n175), .B(n1019), .Z(n1018) );
  XNOR U894 ( .A(p_input[695]), .B(n1017), .Z(n1019) );
  XOR U895 ( .A(n1020), .B(n1021), .Z(n1017) );
  AND U896 ( .A(n179), .B(n1022), .Z(n1021) );
  XNOR U897 ( .A(p_input[711]), .B(n1020), .Z(n1022) );
  XOR U898 ( .A(n1023), .B(n1024), .Z(n1020) );
  AND U899 ( .A(n183), .B(n1025), .Z(n1024) );
  XNOR U900 ( .A(p_input[727]), .B(n1023), .Z(n1025) );
  XOR U901 ( .A(n1026), .B(n1027), .Z(n1023) );
  AND U902 ( .A(n187), .B(n1028), .Z(n1027) );
  XNOR U903 ( .A(p_input[743]), .B(n1026), .Z(n1028) );
  XOR U904 ( .A(n1029), .B(n1030), .Z(n1026) );
  AND U905 ( .A(n191), .B(n1031), .Z(n1030) );
  XNOR U906 ( .A(p_input[759]), .B(n1029), .Z(n1031) );
  XOR U907 ( .A(n1032), .B(n1033), .Z(n1029) );
  AND U908 ( .A(n195), .B(n1034), .Z(n1033) );
  XNOR U909 ( .A(p_input[775]), .B(n1032), .Z(n1034) );
  XOR U910 ( .A(n1035), .B(n1036), .Z(n1032) );
  AND U911 ( .A(n199), .B(n1037), .Z(n1036) );
  XNOR U912 ( .A(p_input[791]), .B(n1035), .Z(n1037) );
  XOR U913 ( .A(n1038), .B(n1039), .Z(n1035) );
  AND U914 ( .A(n203), .B(n1040), .Z(n1039) );
  XNOR U915 ( .A(p_input[807]), .B(n1038), .Z(n1040) );
  XOR U916 ( .A(n1041), .B(n1042), .Z(n1038) );
  AND U917 ( .A(n207), .B(n1043), .Z(n1042) );
  XNOR U918 ( .A(p_input[823]), .B(n1041), .Z(n1043) );
  XOR U919 ( .A(n1044), .B(n1045), .Z(n1041) );
  AND U920 ( .A(n211), .B(n1046), .Z(n1045) );
  XNOR U921 ( .A(p_input[839]), .B(n1044), .Z(n1046) );
  XOR U922 ( .A(n1047), .B(n1048), .Z(n1044) );
  AND U923 ( .A(n215), .B(n1049), .Z(n1048) );
  XNOR U924 ( .A(p_input[855]), .B(n1047), .Z(n1049) );
  XOR U925 ( .A(n1050), .B(n1051), .Z(n1047) );
  AND U926 ( .A(n219), .B(n1052), .Z(n1051) );
  XNOR U927 ( .A(p_input[871]), .B(n1050), .Z(n1052) );
  XOR U928 ( .A(n1053), .B(n1054), .Z(n1050) );
  AND U929 ( .A(n223), .B(n1055), .Z(n1054) );
  XNOR U930 ( .A(p_input[887]), .B(n1053), .Z(n1055) );
  XOR U931 ( .A(n1056), .B(n1057), .Z(n1053) );
  AND U932 ( .A(n227), .B(n1058), .Z(n1057) );
  XNOR U933 ( .A(p_input[903]), .B(n1056), .Z(n1058) );
  XOR U934 ( .A(n1059), .B(n1060), .Z(n1056) );
  AND U935 ( .A(n231), .B(n1061), .Z(n1060) );
  XNOR U936 ( .A(p_input[919]), .B(n1059), .Z(n1061) );
  XOR U937 ( .A(n1062), .B(n1063), .Z(n1059) );
  AND U938 ( .A(n235), .B(n1064), .Z(n1063) );
  XNOR U939 ( .A(p_input[935]), .B(n1062), .Z(n1064) );
  XOR U940 ( .A(n1065), .B(n1066), .Z(n1062) );
  AND U941 ( .A(n239), .B(n1067), .Z(n1066) );
  XNOR U942 ( .A(p_input[951]), .B(n1065), .Z(n1067) );
  XOR U943 ( .A(n1068), .B(n1069), .Z(n1065) );
  AND U944 ( .A(n243), .B(n1070), .Z(n1069) );
  XNOR U945 ( .A(p_input[967]), .B(n1068), .Z(n1070) );
  XOR U946 ( .A(n1071), .B(n1072), .Z(n1068) );
  AND U947 ( .A(n247), .B(n1073), .Z(n1072) );
  XNOR U948 ( .A(p_input[983]), .B(n1071), .Z(n1073) );
  XOR U949 ( .A(n1074), .B(n1075), .Z(n1071) );
  AND U950 ( .A(n251), .B(n1076), .Z(n1075) );
  XNOR U951 ( .A(p_input[999]), .B(n1074), .Z(n1076) );
  XOR U952 ( .A(n1077), .B(n1078), .Z(n1074) );
  AND U953 ( .A(n255), .B(n1079), .Z(n1078) );
  XNOR U954 ( .A(p_input[1015]), .B(n1077), .Z(n1079) );
  XOR U955 ( .A(n1080), .B(n1081), .Z(n1077) );
  AND U956 ( .A(n259), .B(n1082), .Z(n1081) );
  XNOR U957 ( .A(p_input[1031]), .B(n1080), .Z(n1082) );
  XOR U958 ( .A(n1083), .B(n1084), .Z(n1080) );
  AND U959 ( .A(n263), .B(n1085), .Z(n1084) );
  XNOR U960 ( .A(p_input[1047]), .B(n1083), .Z(n1085) );
  XOR U961 ( .A(n1086), .B(n1087), .Z(n1083) );
  AND U962 ( .A(n267), .B(n1088), .Z(n1087) );
  XNOR U963 ( .A(p_input[1063]), .B(n1086), .Z(n1088) );
  XOR U964 ( .A(n1089), .B(n1090), .Z(n1086) );
  AND U965 ( .A(n271), .B(n1091), .Z(n1090) );
  XNOR U966 ( .A(p_input[1079]), .B(n1089), .Z(n1091) );
  XOR U967 ( .A(n1092), .B(n1093), .Z(n1089) );
  AND U968 ( .A(n275), .B(n1094), .Z(n1093) );
  XNOR U969 ( .A(p_input[1095]), .B(n1092), .Z(n1094) );
  XOR U970 ( .A(n1095), .B(n1096), .Z(n1092) );
  AND U971 ( .A(n279), .B(n1097), .Z(n1096) );
  XNOR U972 ( .A(p_input[1111]), .B(n1095), .Z(n1097) );
  XOR U973 ( .A(n1098), .B(n1099), .Z(n1095) );
  AND U974 ( .A(n283), .B(n1100), .Z(n1099) );
  XNOR U975 ( .A(p_input[1127]), .B(n1098), .Z(n1100) );
  XOR U976 ( .A(n1101), .B(n1102), .Z(n1098) );
  AND U977 ( .A(n287), .B(n1103), .Z(n1102) );
  XNOR U978 ( .A(p_input[1143]), .B(n1101), .Z(n1103) );
  XOR U979 ( .A(n1104), .B(n1105), .Z(n1101) );
  AND U980 ( .A(n291), .B(n1106), .Z(n1105) );
  XNOR U981 ( .A(p_input[1159]), .B(n1104), .Z(n1106) );
  XOR U982 ( .A(n1107), .B(n1108), .Z(n1104) );
  AND U983 ( .A(n295), .B(n1109), .Z(n1108) );
  XNOR U984 ( .A(p_input[1175]), .B(n1107), .Z(n1109) );
  XOR U985 ( .A(n1110), .B(n1111), .Z(n1107) );
  AND U986 ( .A(n299), .B(n1112), .Z(n1111) );
  XNOR U987 ( .A(p_input[1191]), .B(n1110), .Z(n1112) );
  XOR U988 ( .A(n1113), .B(n1114), .Z(n1110) );
  AND U989 ( .A(n303), .B(n1115), .Z(n1114) );
  XNOR U990 ( .A(p_input[1207]), .B(n1113), .Z(n1115) );
  XOR U991 ( .A(n1116), .B(n1117), .Z(n1113) );
  AND U992 ( .A(n307), .B(n1118), .Z(n1117) );
  XNOR U993 ( .A(p_input[1223]), .B(n1116), .Z(n1118) );
  XOR U994 ( .A(n1119), .B(n1120), .Z(n1116) );
  AND U995 ( .A(n311), .B(n1121), .Z(n1120) );
  XNOR U996 ( .A(p_input[1239]), .B(n1119), .Z(n1121) );
  XOR U997 ( .A(n1122), .B(n1123), .Z(n1119) );
  AND U998 ( .A(n315), .B(n1124), .Z(n1123) );
  XNOR U999 ( .A(p_input[1255]), .B(n1122), .Z(n1124) );
  XOR U1000 ( .A(n1125), .B(n1126), .Z(n1122) );
  AND U1001 ( .A(n319), .B(n1127), .Z(n1126) );
  XNOR U1002 ( .A(p_input[1271]), .B(n1125), .Z(n1127) );
  XOR U1003 ( .A(n1128), .B(n1129), .Z(n1125) );
  AND U1004 ( .A(n323), .B(n1130), .Z(n1129) );
  XNOR U1005 ( .A(p_input[1287]), .B(n1128), .Z(n1130) );
  XOR U1006 ( .A(n1131), .B(n1132), .Z(n1128) );
  AND U1007 ( .A(n327), .B(n1133), .Z(n1132) );
  XNOR U1008 ( .A(p_input[1303]), .B(n1131), .Z(n1133) );
  XOR U1009 ( .A(n1134), .B(n1135), .Z(n1131) );
  AND U1010 ( .A(n331), .B(n1136), .Z(n1135) );
  XNOR U1011 ( .A(p_input[1319]), .B(n1134), .Z(n1136) );
  XOR U1012 ( .A(n1137), .B(n1138), .Z(n1134) );
  AND U1013 ( .A(n335), .B(n1139), .Z(n1138) );
  XNOR U1014 ( .A(p_input[1335]), .B(n1137), .Z(n1139) );
  XOR U1015 ( .A(n1140), .B(n1141), .Z(n1137) );
  AND U1016 ( .A(n339), .B(n1142), .Z(n1141) );
  XNOR U1017 ( .A(p_input[1351]), .B(n1140), .Z(n1142) );
  XOR U1018 ( .A(n1143), .B(n1144), .Z(n1140) );
  AND U1019 ( .A(n343), .B(n1145), .Z(n1144) );
  XNOR U1020 ( .A(p_input[1367]), .B(n1143), .Z(n1145) );
  XOR U1021 ( .A(n1146), .B(n1147), .Z(n1143) );
  AND U1022 ( .A(n347), .B(n1148), .Z(n1147) );
  XNOR U1023 ( .A(p_input[1383]), .B(n1146), .Z(n1148) );
  XOR U1024 ( .A(n1149), .B(n1150), .Z(n1146) );
  AND U1025 ( .A(n351), .B(n1151), .Z(n1150) );
  XNOR U1026 ( .A(p_input[1399]), .B(n1149), .Z(n1151) );
  XOR U1027 ( .A(n1152), .B(n1153), .Z(n1149) );
  AND U1028 ( .A(n355), .B(n1154), .Z(n1153) );
  XNOR U1029 ( .A(p_input[1415]), .B(n1152), .Z(n1154) );
  XOR U1030 ( .A(n1155), .B(n1156), .Z(n1152) );
  AND U1031 ( .A(n359), .B(n1157), .Z(n1156) );
  XNOR U1032 ( .A(p_input[1431]), .B(n1155), .Z(n1157) );
  XOR U1033 ( .A(n1158), .B(n1159), .Z(n1155) );
  AND U1034 ( .A(n363), .B(n1160), .Z(n1159) );
  XNOR U1035 ( .A(p_input[1447]), .B(n1158), .Z(n1160) );
  XOR U1036 ( .A(n1161), .B(n1162), .Z(n1158) );
  AND U1037 ( .A(n367), .B(n1163), .Z(n1162) );
  XNOR U1038 ( .A(p_input[1463]), .B(n1161), .Z(n1163) );
  XOR U1039 ( .A(n1164), .B(n1165), .Z(n1161) );
  AND U1040 ( .A(n371), .B(n1166), .Z(n1165) );
  XNOR U1041 ( .A(p_input[1479]), .B(n1164), .Z(n1166) );
  XOR U1042 ( .A(n1167), .B(n1168), .Z(n1164) );
  AND U1043 ( .A(n375), .B(n1169), .Z(n1168) );
  XNOR U1044 ( .A(p_input[1495]), .B(n1167), .Z(n1169) );
  XOR U1045 ( .A(n1170), .B(n1171), .Z(n1167) );
  AND U1046 ( .A(n379), .B(n1172), .Z(n1171) );
  XNOR U1047 ( .A(p_input[1511]), .B(n1170), .Z(n1172) );
  XOR U1048 ( .A(n1173), .B(n1174), .Z(n1170) );
  AND U1049 ( .A(n383), .B(n1175), .Z(n1174) );
  XNOR U1050 ( .A(p_input[1527]), .B(n1173), .Z(n1175) );
  XOR U1051 ( .A(n1176), .B(n1177), .Z(n1173) );
  AND U1052 ( .A(n387), .B(n1178), .Z(n1177) );
  XNOR U1053 ( .A(p_input[1543]), .B(n1176), .Z(n1178) );
  XOR U1054 ( .A(n1179), .B(n1180), .Z(n1176) );
  AND U1055 ( .A(n391), .B(n1181), .Z(n1180) );
  XNOR U1056 ( .A(p_input[1559]), .B(n1179), .Z(n1181) );
  XOR U1057 ( .A(n1182), .B(n1183), .Z(n1179) );
  AND U1058 ( .A(n395), .B(n1184), .Z(n1183) );
  XNOR U1059 ( .A(p_input[1575]), .B(n1182), .Z(n1184) );
  XOR U1060 ( .A(n1185), .B(n1186), .Z(n1182) );
  AND U1061 ( .A(n399), .B(n1187), .Z(n1186) );
  XNOR U1062 ( .A(p_input[1591]), .B(n1185), .Z(n1187) );
  XOR U1063 ( .A(n1188), .B(n1189), .Z(n1185) );
  AND U1064 ( .A(n403), .B(n1190), .Z(n1189) );
  XNOR U1065 ( .A(p_input[1607]), .B(n1188), .Z(n1190) );
  XOR U1066 ( .A(n1191), .B(n1192), .Z(n1188) );
  AND U1067 ( .A(n407), .B(n1193), .Z(n1192) );
  XNOR U1068 ( .A(p_input[1623]), .B(n1191), .Z(n1193) );
  XOR U1069 ( .A(n1194), .B(n1195), .Z(n1191) );
  AND U1070 ( .A(n411), .B(n1196), .Z(n1195) );
  XNOR U1071 ( .A(p_input[1639]), .B(n1194), .Z(n1196) );
  XOR U1072 ( .A(n1197), .B(n1198), .Z(n1194) );
  AND U1073 ( .A(n415), .B(n1199), .Z(n1198) );
  XNOR U1074 ( .A(p_input[1655]), .B(n1197), .Z(n1199) );
  XOR U1075 ( .A(n1200), .B(n1201), .Z(n1197) );
  AND U1076 ( .A(n419), .B(n1202), .Z(n1201) );
  XNOR U1077 ( .A(p_input[1671]), .B(n1200), .Z(n1202) );
  XOR U1078 ( .A(n1203), .B(n1204), .Z(n1200) );
  AND U1079 ( .A(n423), .B(n1205), .Z(n1204) );
  XNOR U1080 ( .A(p_input[1687]), .B(n1203), .Z(n1205) );
  XOR U1081 ( .A(n1206), .B(n1207), .Z(n1203) );
  AND U1082 ( .A(n427), .B(n1208), .Z(n1207) );
  XNOR U1083 ( .A(p_input[1703]), .B(n1206), .Z(n1208) );
  XOR U1084 ( .A(n1209), .B(n1210), .Z(n1206) );
  AND U1085 ( .A(n431), .B(n1211), .Z(n1210) );
  XNOR U1086 ( .A(p_input[1719]), .B(n1209), .Z(n1211) );
  XOR U1087 ( .A(n1212), .B(n1213), .Z(n1209) );
  AND U1088 ( .A(n435), .B(n1214), .Z(n1213) );
  XNOR U1089 ( .A(p_input[1735]), .B(n1212), .Z(n1214) );
  XOR U1090 ( .A(n1215), .B(n1216), .Z(n1212) );
  AND U1091 ( .A(n439), .B(n1217), .Z(n1216) );
  XNOR U1092 ( .A(p_input[1751]), .B(n1215), .Z(n1217) );
  XOR U1093 ( .A(n1218), .B(n1219), .Z(n1215) );
  AND U1094 ( .A(n443), .B(n1220), .Z(n1219) );
  XNOR U1095 ( .A(p_input[1767]), .B(n1218), .Z(n1220) );
  XOR U1096 ( .A(n1221), .B(n1222), .Z(n1218) );
  AND U1097 ( .A(n447), .B(n1223), .Z(n1222) );
  XNOR U1098 ( .A(p_input[1783]), .B(n1221), .Z(n1223) );
  XOR U1099 ( .A(n1224), .B(n1225), .Z(n1221) );
  AND U1100 ( .A(n451), .B(n1226), .Z(n1225) );
  XNOR U1101 ( .A(p_input[1799]), .B(n1224), .Z(n1226) );
  XOR U1102 ( .A(n1227), .B(n1228), .Z(n1224) );
  AND U1103 ( .A(n455), .B(n1229), .Z(n1228) );
  XNOR U1104 ( .A(p_input[1815]), .B(n1227), .Z(n1229) );
  XOR U1105 ( .A(n1230), .B(n1231), .Z(n1227) );
  AND U1106 ( .A(n459), .B(n1232), .Z(n1231) );
  XNOR U1107 ( .A(p_input[1831]), .B(n1230), .Z(n1232) );
  XOR U1108 ( .A(n1233), .B(n1234), .Z(n1230) );
  AND U1109 ( .A(n463), .B(n1235), .Z(n1234) );
  XNOR U1110 ( .A(p_input[1847]), .B(n1233), .Z(n1235) );
  XOR U1111 ( .A(n1236), .B(n1237), .Z(n1233) );
  AND U1112 ( .A(n467), .B(n1238), .Z(n1237) );
  XNOR U1113 ( .A(p_input[1863]), .B(n1236), .Z(n1238) );
  XOR U1114 ( .A(n1239), .B(n1240), .Z(n1236) );
  AND U1115 ( .A(n471), .B(n1241), .Z(n1240) );
  XNOR U1116 ( .A(p_input[1879]), .B(n1239), .Z(n1241) );
  XOR U1117 ( .A(n1242), .B(n1243), .Z(n1239) );
  AND U1118 ( .A(n475), .B(n1244), .Z(n1243) );
  XNOR U1119 ( .A(p_input[1895]), .B(n1242), .Z(n1244) );
  XOR U1120 ( .A(n1245), .B(n1246), .Z(n1242) );
  AND U1121 ( .A(n479), .B(n1247), .Z(n1246) );
  XNOR U1122 ( .A(p_input[1911]), .B(n1245), .Z(n1247) );
  XOR U1123 ( .A(n1248), .B(n1249), .Z(n1245) );
  AND U1124 ( .A(n483), .B(n1250), .Z(n1249) );
  XNOR U1125 ( .A(p_input[1927]), .B(n1248), .Z(n1250) );
  XOR U1126 ( .A(n1251), .B(n1252), .Z(n1248) );
  AND U1127 ( .A(n487), .B(n1253), .Z(n1252) );
  XNOR U1128 ( .A(p_input[1943]), .B(n1251), .Z(n1253) );
  XOR U1129 ( .A(n1254), .B(n1255), .Z(n1251) );
  AND U1130 ( .A(n491), .B(n1256), .Z(n1255) );
  XNOR U1131 ( .A(p_input[1959]), .B(n1254), .Z(n1256) );
  XOR U1132 ( .A(n1257), .B(n1258), .Z(n1254) );
  AND U1133 ( .A(n495), .B(n1259), .Z(n1258) );
  XNOR U1134 ( .A(p_input[1975]), .B(n1257), .Z(n1259) );
  XOR U1135 ( .A(n1260), .B(n1261), .Z(n1257) );
  AND U1136 ( .A(n499), .B(n1262), .Z(n1261) );
  XNOR U1137 ( .A(p_input[1991]), .B(n1260), .Z(n1262) );
  XNOR U1138 ( .A(n1263), .B(n1264), .Z(n1260) );
  AND U1139 ( .A(n503), .B(n1265), .Z(n1264) );
  XOR U1140 ( .A(p_input[2007]), .B(n1263), .Z(n1265) );
  XOR U1141 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n1266), .Z(n1263) );
  AND U1142 ( .A(n506), .B(n1267), .Z(n1266) );
  XOR U1143 ( .A(p_input[2023]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n1267)
         );
  XNOR U1144 ( .A(n1268), .B(n1269), .Z(o[6]) );
  AND U1145 ( .A(n3), .B(n1270), .Z(n1268) );
  XNOR U1146 ( .A(p_input[6]), .B(n1269), .Z(n1270) );
  XOR U1147 ( .A(n1271), .B(n1272), .Z(n1269) );
  AND U1148 ( .A(n7), .B(n1273), .Z(n1272) );
  XNOR U1149 ( .A(p_input[22]), .B(n1271), .Z(n1273) );
  XOR U1150 ( .A(n1274), .B(n1275), .Z(n1271) );
  AND U1151 ( .A(n11), .B(n1276), .Z(n1275) );
  XNOR U1152 ( .A(p_input[38]), .B(n1274), .Z(n1276) );
  XOR U1153 ( .A(n1277), .B(n1278), .Z(n1274) );
  AND U1154 ( .A(n15), .B(n1279), .Z(n1278) );
  XNOR U1155 ( .A(p_input[54]), .B(n1277), .Z(n1279) );
  XOR U1156 ( .A(n1280), .B(n1281), .Z(n1277) );
  AND U1157 ( .A(n19), .B(n1282), .Z(n1281) );
  XNOR U1158 ( .A(p_input[70]), .B(n1280), .Z(n1282) );
  XOR U1159 ( .A(n1283), .B(n1284), .Z(n1280) );
  AND U1160 ( .A(n23), .B(n1285), .Z(n1284) );
  XNOR U1161 ( .A(p_input[86]), .B(n1283), .Z(n1285) );
  XOR U1162 ( .A(n1286), .B(n1287), .Z(n1283) );
  AND U1163 ( .A(n27), .B(n1288), .Z(n1287) );
  XNOR U1164 ( .A(p_input[102]), .B(n1286), .Z(n1288) );
  XOR U1165 ( .A(n1289), .B(n1290), .Z(n1286) );
  AND U1166 ( .A(n31), .B(n1291), .Z(n1290) );
  XNOR U1167 ( .A(p_input[118]), .B(n1289), .Z(n1291) );
  XOR U1168 ( .A(n1292), .B(n1293), .Z(n1289) );
  AND U1169 ( .A(n35), .B(n1294), .Z(n1293) );
  XNOR U1170 ( .A(p_input[134]), .B(n1292), .Z(n1294) );
  XOR U1171 ( .A(n1295), .B(n1296), .Z(n1292) );
  AND U1172 ( .A(n39), .B(n1297), .Z(n1296) );
  XNOR U1173 ( .A(p_input[150]), .B(n1295), .Z(n1297) );
  XOR U1174 ( .A(n1298), .B(n1299), .Z(n1295) );
  AND U1175 ( .A(n43), .B(n1300), .Z(n1299) );
  XNOR U1176 ( .A(p_input[166]), .B(n1298), .Z(n1300) );
  XOR U1177 ( .A(n1301), .B(n1302), .Z(n1298) );
  AND U1178 ( .A(n47), .B(n1303), .Z(n1302) );
  XNOR U1179 ( .A(p_input[182]), .B(n1301), .Z(n1303) );
  XOR U1180 ( .A(n1304), .B(n1305), .Z(n1301) );
  AND U1181 ( .A(n51), .B(n1306), .Z(n1305) );
  XNOR U1182 ( .A(p_input[198]), .B(n1304), .Z(n1306) );
  XOR U1183 ( .A(n1307), .B(n1308), .Z(n1304) );
  AND U1184 ( .A(n55), .B(n1309), .Z(n1308) );
  XNOR U1185 ( .A(p_input[214]), .B(n1307), .Z(n1309) );
  XOR U1186 ( .A(n1310), .B(n1311), .Z(n1307) );
  AND U1187 ( .A(n59), .B(n1312), .Z(n1311) );
  XNOR U1188 ( .A(p_input[230]), .B(n1310), .Z(n1312) );
  XOR U1189 ( .A(n1313), .B(n1314), .Z(n1310) );
  AND U1190 ( .A(n63), .B(n1315), .Z(n1314) );
  XNOR U1191 ( .A(p_input[246]), .B(n1313), .Z(n1315) );
  XOR U1192 ( .A(n1316), .B(n1317), .Z(n1313) );
  AND U1193 ( .A(n67), .B(n1318), .Z(n1317) );
  XNOR U1194 ( .A(p_input[262]), .B(n1316), .Z(n1318) );
  XOR U1195 ( .A(n1319), .B(n1320), .Z(n1316) );
  AND U1196 ( .A(n71), .B(n1321), .Z(n1320) );
  XNOR U1197 ( .A(p_input[278]), .B(n1319), .Z(n1321) );
  XOR U1198 ( .A(n1322), .B(n1323), .Z(n1319) );
  AND U1199 ( .A(n75), .B(n1324), .Z(n1323) );
  XNOR U1200 ( .A(p_input[294]), .B(n1322), .Z(n1324) );
  XOR U1201 ( .A(n1325), .B(n1326), .Z(n1322) );
  AND U1202 ( .A(n79), .B(n1327), .Z(n1326) );
  XNOR U1203 ( .A(p_input[310]), .B(n1325), .Z(n1327) );
  XOR U1204 ( .A(n1328), .B(n1329), .Z(n1325) );
  AND U1205 ( .A(n83), .B(n1330), .Z(n1329) );
  XNOR U1206 ( .A(p_input[326]), .B(n1328), .Z(n1330) );
  XOR U1207 ( .A(n1331), .B(n1332), .Z(n1328) );
  AND U1208 ( .A(n87), .B(n1333), .Z(n1332) );
  XNOR U1209 ( .A(p_input[342]), .B(n1331), .Z(n1333) );
  XOR U1210 ( .A(n1334), .B(n1335), .Z(n1331) );
  AND U1211 ( .A(n91), .B(n1336), .Z(n1335) );
  XNOR U1212 ( .A(p_input[358]), .B(n1334), .Z(n1336) );
  XOR U1213 ( .A(n1337), .B(n1338), .Z(n1334) );
  AND U1214 ( .A(n95), .B(n1339), .Z(n1338) );
  XNOR U1215 ( .A(p_input[374]), .B(n1337), .Z(n1339) );
  XOR U1216 ( .A(n1340), .B(n1341), .Z(n1337) );
  AND U1217 ( .A(n99), .B(n1342), .Z(n1341) );
  XNOR U1218 ( .A(p_input[390]), .B(n1340), .Z(n1342) );
  XOR U1219 ( .A(n1343), .B(n1344), .Z(n1340) );
  AND U1220 ( .A(n103), .B(n1345), .Z(n1344) );
  XNOR U1221 ( .A(p_input[406]), .B(n1343), .Z(n1345) );
  XOR U1222 ( .A(n1346), .B(n1347), .Z(n1343) );
  AND U1223 ( .A(n107), .B(n1348), .Z(n1347) );
  XNOR U1224 ( .A(p_input[422]), .B(n1346), .Z(n1348) );
  XOR U1225 ( .A(n1349), .B(n1350), .Z(n1346) );
  AND U1226 ( .A(n111), .B(n1351), .Z(n1350) );
  XNOR U1227 ( .A(p_input[438]), .B(n1349), .Z(n1351) );
  XOR U1228 ( .A(n1352), .B(n1353), .Z(n1349) );
  AND U1229 ( .A(n115), .B(n1354), .Z(n1353) );
  XNOR U1230 ( .A(p_input[454]), .B(n1352), .Z(n1354) );
  XOR U1231 ( .A(n1355), .B(n1356), .Z(n1352) );
  AND U1232 ( .A(n119), .B(n1357), .Z(n1356) );
  XNOR U1233 ( .A(p_input[470]), .B(n1355), .Z(n1357) );
  XOR U1234 ( .A(n1358), .B(n1359), .Z(n1355) );
  AND U1235 ( .A(n123), .B(n1360), .Z(n1359) );
  XNOR U1236 ( .A(p_input[486]), .B(n1358), .Z(n1360) );
  XOR U1237 ( .A(n1361), .B(n1362), .Z(n1358) );
  AND U1238 ( .A(n127), .B(n1363), .Z(n1362) );
  XNOR U1239 ( .A(p_input[502]), .B(n1361), .Z(n1363) );
  XOR U1240 ( .A(n1364), .B(n1365), .Z(n1361) );
  AND U1241 ( .A(n131), .B(n1366), .Z(n1365) );
  XNOR U1242 ( .A(p_input[518]), .B(n1364), .Z(n1366) );
  XOR U1243 ( .A(n1367), .B(n1368), .Z(n1364) );
  AND U1244 ( .A(n135), .B(n1369), .Z(n1368) );
  XNOR U1245 ( .A(p_input[534]), .B(n1367), .Z(n1369) );
  XOR U1246 ( .A(n1370), .B(n1371), .Z(n1367) );
  AND U1247 ( .A(n139), .B(n1372), .Z(n1371) );
  XNOR U1248 ( .A(p_input[550]), .B(n1370), .Z(n1372) );
  XOR U1249 ( .A(n1373), .B(n1374), .Z(n1370) );
  AND U1250 ( .A(n143), .B(n1375), .Z(n1374) );
  XNOR U1251 ( .A(p_input[566]), .B(n1373), .Z(n1375) );
  XOR U1252 ( .A(n1376), .B(n1377), .Z(n1373) );
  AND U1253 ( .A(n147), .B(n1378), .Z(n1377) );
  XNOR U1254 ( .A(p_input[582]), .B(n1376), .Z(n1378) );
  XOR U1255 ( .A(n1379), .B(n1380), .Z(n1376) );
  AND U1256 ( .A(n151), .B(n1381), .Z(n1380) );
  XNOR U1257 ( .A(p_input[598]), .B(n1379), .Z(n1381) );
  XOR U1258 ( .A(n1382), .B(n1383), .Z(n1379) );
  AND U1259 ( .A(n155), .B(n1384), .Z(n1383) );
  XNOR U1260 ( .A(p_input[614]), .B(n1382), .Z(n1384) );
  XOR U1261 ( .A(n1385), .B(n1386), .Z(n1382) );
  AND U1262 ( .A(n159), .B(n1387), .Z(n1386) );
  XNOR U1263 ( .A(p_input[630]), .B(n1385), .Z(n1387) );
  XOR U1264 ( .A(n1388), .B(n1389), .Z(n1385) );
  AND U1265 ( .A(n163), .B(n1390), .Z(n1389) );
  XNOR U1266 ( .A(p_input[646]), .B(n1388), .Z(n1390) );
  XOR U1267 ( .A(n1391), .B(n1392), .Z(n1388) );
  AND U1268 ( .A(n167), .B(n1393), .Z(n1392) );
  XNOR U1269 ( .A(p_input[662]), .B(n1391), .Z(n1393) );
  XOR U1270 ( .A(n1394), .B(n1395), .Z(n1391) );
  AND U1271 ( .A(n171), .B(n1396), .Z(n1395) );
  XNOR U1272 ( .A(p_input[678]), .B(n1394), .Z(n1396) );
  XOR U1273 ( .A(n1397), .B(n1398), .Z(n1394) );
  AND U1274 ( .A(n175), .B(n1399), .Z(n1398) );
  XNOR U1275 ( .A(p_input[694]), .B(n1397), .Z(n1399) );
  XOR U1276 ( .A(n1400), .B(n1401), .Z(n1397) );
  AND U1277 ( .A(n179), .B(n1402), .Z(n1401) );
  XNOR U1278 ( .A(p_input[710]), .B(n1400), .Z(n1402) );
  XOR U1279 ( .A(n1403), .B(n1404), .Z(n1400) );
  AND U1280 ( .A(n183), .B(n1405), .Z(n1404) );
  XNOR U1281 ( .A(p_input[726]), .B(n1403), .Z(n1405) );
  XOR U1282 ( .A(n1406), .B(n1407), .Z(n1403) );
  AND U1283 ( .A(n187), .B(n1408), .Z(n1407) );
  XNOR U1284 ( .A(p_input[742]), .B(n1406), .Z(n1408) );
  XOR U1285 ( .A(n1409), .B(n1410), .Z(n1406) );
  AND U1286 ( .A(n191), .B(n1411), .Z(n1410) );
  XNOR U1287 ( .A(p_input[758]), .B(n1409), .Z(n1411) );
  XOR U1288 ( .A(n1412), .B(n1413), .Z(n1409) );
  AND U1289 ( .A(n195), .B(n1414), .Z(n1413) );
  XNOR U1290 ( .A(p_input[774]), .B(n1412), .Z(n1414) );
  XOR U1291 ( .A(n1415), .B(n1416), .Z(n1412) );
  AND U1292 ( .A(n199), .B(n1417), .Z(n1416) );
  XNOR U1293 ( .A(p_input[790]), .B(n1415), .Z(n1417) );
  XOR U1294 ( .A(n1418), .B(n1419), .Z(n1415) );
  AND U1295 ( .A(n203), .B(n1420), .Z(n1419) );
  XNOR U1296 ( .A(p_input[806]), .B(n1418), .Z(n1420) );
  XOR U1297 ( .A(n1421), .B(n1422), .Z(n1418) );
  AND U1298 ( .A(n207), .B(n1423), .Z(n1422) );
  XNOR U1299 ( .A(p_input[822]), .B(n1421), .Z(n1423) );
  XOR U1300 ( .A(n1424), .B(n1425), .Z(n1421) );
  AND U1301 ( .A(n211), .B(n1426), .Z(n1425) );
  XNOR U1302 ( .A(p_input[838]), .B(n1424), .Z(n1426) );
  XOR U1303 ( .A(n1427), .B(n1428), .Z(n1424) );
  AND U1304 ( .A(n215), .B(n1429), .Z(n1428) );
  XNOR U1305 ( .A(p_input[854]), .B(n1427), .Z(n1429) );
  XOR U1306 ( .A(n1430), .B(n1431), .Z(n1427) );
  AND U1307 ( .A(n219), .B(n1432), .Z(n1431) );
  XNOR U1308 ( .A(p_input[870]), .B(n1430), .Z(n1432) );
  XOR U1309 ( .A(n1433), .B(n1434), .Z(n1430) );
  AND U1310 ( .A(n223), .B(n1435), .Z(n1434) );
  XNOR U1311 ( .A(p_input[886]), .B(n1433), .Z(n1435) );
  XOR U1312 ( .A(n1436), .B(n1437), .Z(n1433) );
  AND U1313 ( .A(n227), .B(n1438), .Z(n1437) );
  XNOR U1314 ( .A(p_input[902]), .B(n1436), .Z(n1438) );
  XOR U1315 ( .A(n1439), .B(n1440), .Z(n1436) );
  AND U1316 ( .A(n231), .B(n1441), .Z(n1440) );
  XNOR U1317 ( .A(p_input[918]), .B(n1439), .Z(n1441) );
  XOR U1318 ( .A(n1442), .B(n1443), .Z(n1439) );
  AND U1319 ( .A(n235), .B(n1444), .Z(n1443) );
  XNOR U1320 ( .A(p_input[934]), .B(n1442), .Z(n1444) );
  XOR U1321 ( .A(n1445), .B(n1446), .Z(n1442) );
  AND U1322 ( .A(n239), .B(n1447), .Z(n1446) );
  XNOR U1323 ( .A(p_input[950]), .B(n1445), .Z(n1447) );
  XOR U1324 ( .A(n1448), .B(n1449), .Z(n1445) );
  AND U1325 ( .A(n243), .B(n1450), .Z(n1449) );
  XNOR U1326 ( .A(p_input[966]), .B(n1448), .Z(n1450) );
  XOR U1327 ( .A(n1451), .B(n1452), .Z(n1448) );
  AND U1328 ( .A(n247), .B(n1453), .Z(n1452) );
  XNOR U1329 ( .A(p_input[982]), .B(n1451), .Z(n1453) );
  XOR U1330 ( .A(n1454), .B(n1455), .Z(n1451) );
  AND U1331 ( .A(n251), .B(n1456), .Z(n1455) );
  XNOR U1332 ( .A(p_input[998]), .B(n1454), .Z(n1456) );
  XOR U1333 ( .A(n1457), .B(n1458), .Z(n1454) );
  AND U1334 ( .A(n255), .B(n1459), .Z(n1458) );
  XNOR U1335 ( .A(p_input[1014]), .B(n1457), .Z(n1459) );
  XOR U1336 ( .A(n1460), .B(n1461), .Z(n1457) );
  AND U1337 ( .A(n259), .B(n1462), .Z(n1461) );
  XNOR U1338 ( .A(p_input[1030]), .B(n1460), .Z(n1462) );
  XOR U1339 ( .A(n1463), .B(n1464), .Z(n1460) );
  AND U1340 ( .A(n263), .B(n1465), .Z(n1464) );
  XNOR U1341 ( .A(p_input[1046]), .B(n1463), .Z(n1465) );
  XOR U1342 ( .A(n1466), .B(n1467), .Z(n1463) );
  AND U1343 ( .A(n267), .B(n1468), .Z(n1467) );
  XNOR U1344 ( .A(p_input[1062]), .B(n1466), .Z(n1468) );
  XOR U1345 ( .A(n1469), .B(n1470), .Z(n1466) );
  AND U1346 ( .A(n271), .B(n1471), .Z(n1470) );
  XNOR U1347 ( .A(p_input[1078]), .B(n1469), .Z(n1471) );
  XOR U1348 ( .A(n1472), .B(n1473), .Z(n1469) );
  AND U1349 ( .A(n275), .B(n1474), .Z(n1473) );
  XNOR U1350 ( .A(p_input[1094]), .B(n1472), .Z(n1474) );
  XOR U1351 ( .A(n1475), .B(n1476), .Z(n1472) );
  AND U1352 ( .A(n279), .B(n1477), .Z(n1476) );
  XNOR U1353 ( .A(p_input[1110]), .B(n1475), .Z(n1477) );
  XOR U1354 ( .A(n1478), .B(n1479), .Z(n1475) );
  AND U1355 ( .A(n283), .B(n1480), .Z(n1479) );
  XNOR U1356 ( .A(p_input[1126]), .B(n1478), .Z(n1480) );
  XOR U1357 ( .A(n1481), .B(n1482), .Z(n1478) );
  AND U1358 ( .A(n287), .B(n1483), .Z(n1482) );
  XNOR U1359 ( .A(p_input[1142]), .B(n1481), .Z(n1483) );
  XOR U1360 ( .A(n1484), .B(n1485), .Z(n1481) );
  AND U1361 ( .A(n291), .B(n1486), .Z(n1485) );
  XNOR U1362 ( .A(p_input[1158]), .B(n1484), .Z(n1486) );
  XOR U1363 ( .A(n1487), .B(n1488), .Z(n1484) );
  AND U1364 ( .A(n295), .B(n1489), .Z(n1488) );
  XNOR U1365 ( .A(p_input[1174]), .B(n1487), .Z(n1489) );
  XOR U1366 ( .A(n1490), .B(n1491), .Z(n1487) );
  AND U1367 ( .A(n299), .B(n1492), .Z(n1491) );
  XNOR U1368 ( .A(p_input[1190]), .B(n1490), .Z(n1492) );
  XOR U1369 ( .A(n1493), .B(n1494), .Z(n1490) );
  AND U1370 ( .A(n303), .B(n1495), .Z(n1494) );
  XNOR U1371 ( .A(p_input[1206]), .B(n1493), .Z(n1495) );
  XOR U1372 ( .A(n1496), .B(n1497), .Z(n1493) );
  AND U1373 ( .A(n307), .B(n1498), .Z(n1497) );
  XNOR U1374 ( .A(p_input[1222]), .B(n1496), .Z(n1498) );
  XOR U1375 ( .A(n1499), .B(n1500), .Z(n1496) );
  AND U1376 ( .A(n311), .B(n1501), .Z(n1500) );
  XNOR U1377 ( .A(p_input[1238]), .B(n1499), .Z(n1501) );
  XOR U1378 ( .A(n1502), .B(n1503), .Z(n1499) );
  AND U1379 ( .A(n315), .B(n1504), .Z(n1503) );
  XNOR U1380 ( .A(p_input[1254]), .B(n1502), .Z(n1504) );
  XOR U1381 ( .A(n1505), .B(n1506), .Z(n1502) );
  AND U1382 ( .A(n319), .B(n1507), .Z(n1506) );
  XNOR U1383 ( .A(p_input[1270]), .B(n1505), .Z(n1507) );
  XOR U1384 ( .A(n1508), .B(n1509), .Z(n1505) );
  AND U1385 ( .A(n323), .B(n1510), .Z(n1509) );
  XNOR U1386 ( .A(p_input[1286]), .B(n1508), .Z(n1510) );
  XOR U1387 ( .A(n1511), .B(n1512), .Z(n1508) );
  AND U1388 ( .A(n327), .B(n1513), .Z(n1512) );
  XNOR U1389 ( .A(p_input[1302]), .B(n1511), .Z(n1513) );
  XOR U1390 ( .A(n1514), .B(n1515), .Z(n1511) );
  AND U1391 ( .A(n331), .B(n1516), .Z(n1515) );
  XNOR U1392 ( .A(p_input[1318]), .B(n1514), .Z(n1516) );
  XOR U1393 ( .A(n1517), .B(n1518), .Z(n1514) );
  AND U1394 ( .A(n335), .B(n1519), .Z(n1518) );
  XNOR U1395 ( .A(p_input[1334]), .B(n1517), .Z(n1519) );
  XOR U1396 ( .A(n1520), .B(n1521), .Z(n1517) );
  AND U1397 ( .A(n339), .B(n1522), .Z(n1521) );
  XNOR U1398 ( .A(p_input[1350]), .B(n1520), .Z(n1522) );
  XOR U1399 ( .A(n1523), .B(n1524), .Z(n1520) );
  AND U1400 ( .A(n343), .B(n1525), .Z(n1524) );
  XNOR U1401 ( .A(p_input[1366]), .B(n1523), .Z(n1525) );
  XOR U1402 ( .A(n1526), .B(n1527), .Z(n1523) );
  AND U1403 ( .A(n347), .B(n1528), .Z(n1527) );
  XNOR U1404 ( .A(p_input[1382]), .B(n1526), .Z(n1528) );
  XOR U1405 ( .A(n1529), .B(n1530), .Z(n1526) );
  AND U1406 ( .A(n351), .B(n1531), .Z(n1530) );
  XNOR U1407 ( .A(p_input[1398]), .B(n1529), .Z(n1531) );
  XOR U1408 ( .A(n1532), .B(n1533), .Z(n1529) );
  AND U1409 ( .A(n355), .B(n1534), .Z(n1533) );
  XNOR U1410 ( .A(p_input[1414]), .B(n1532), .Z(n1534) );
  XOR U1411 ( .A(n1535), .B(n1536), .Z(n1532) );
  AND U1412 ( .A(n359), .B(n1537), .Z(n1536) );
  XNOR U1413 ( .A(p_input[1430]), .B(n1535), .Z(n1537) );
  XOR U1414 ( .A(n1538), .B(n1539), .Z(n1535) );
  AND U1415 ( .A(n363), .B(n1540), .Z(n1539) );
  XNOR U1416 ( .A(p_input[1446]), .B(n1538), .Z(n1540) );
  XOR U1417 ( .A(n1541), .B(n1542), .Z(n1538) );
  AND U1418 ( .A(n367), .B(n1543), .Z(n1542) );
  XNOR U1419 ( .A(p_input[1462]), .B(n1541), .Z(n1543) );
  XOR U1420 ( .A(n1544), .B(n1545), .Z(n1541) );
  AND U1421 ( .A(n371), .B(n1546), .Z(n1545) );
  XNOR U1422 ( .A(p_input[1478]), .B(n1544), .Z(n1546) );
  XOR U1423 ( .A(n1547), .B(n1548), .Z(n1544) );
  AND U1424 ( .A(n375), .B(n1549), .Z(n1548) );
  XNOR U1425 ( .A(p_input[1494]), .B(n1547), .Z(n1549) );
  XOR U1426 ( .A(n1550), .B(n1551), .Z(n1547) );
  AND U1427 ( .A(n379), .B(n1552), .Z(n1551) );
  XNOR U1428 ( .A(p_input[1510]), .B(n1550), .Z(n1552) );
  XOR U1429 ( .A(n1553), .B(n1554), .Z(n1550) );
  AND U1430 ( .A(n383), .B(n1555), .Z(n1554) );
  XNOR U1431 ( .A(p_input[1526]), .B(n1553), .Z(n1555) );
  XOR U1432 ( .A(n1556), .B(n1557), .Z(n1553) );
  AND U1433 ( .A(n387), .B(n1558), .Z(n1557) );
  XNOR U1434 ( .A(p_input[1542]), .B(n1556), .Z(n1558) );
  XOR U1435 ( .A(n1559), .B(n1560), .Z(n1556) );
  AND U1436 ( .A(n391), .B(n1561), .Z(n1560) );
  XNOR U1437 ( .A(p_input[1558]), .B(n1559), .Z(n1561) );
  XOR U1438 ( .A(n1562), .B(n1563), .Z(n1559) );
  AND U1439 ( .A(n395), .B(n1564), .Z(n1563) );
  XNOR U1440 ( .A(p_input[1574]), .B(n1562), .Z(n1564) );
  XOR U1441 ( .A(n1565), .B(n1566), .Z(n1562) );
  AND U1442 ( .A(n399), .B(n1567), .Z(n1566) );
  XNOR U1443 ( .A(p_input[1590]), .B(n1565), .Z(n1567) );
  XOR U1444 ( .A(n1568), .B(n1569), .Z(n1565) );
  AND U1445 ( .A(n403), .B(n1570), .Z(n1569) );
  XNOR U1446 ( .A(p_input[1606]), .B(n1568), .Z(n1570) );
  XOR U1447 ( .A(n1571), .B(n1572), .Z(n1568) );
  AND U1448 ( .A(n407), .B(n1573), .Z(n1572) );
  XNOR U1449 ( .A(p_input[1622]), .B(n1571), .Z(n1573) );
  XOR U1450 ( .A(n1574), .B(n1575), .Z(n1571) );
  AND U1451 ( .A(n411), .B(n1576), .Z(n1575) );
  XNOR U1452 ( .A(p_input[1638]), .B(n1574), .Z(n1576) );
  XOR U1453 ( .A(n1577), .B(n1578), .Z(n1574) );
  AND U1454 ( .A(n415), .B(n1579), .Z(n1578) );
  XNOR U1455 ( .A(p_input[1654]), .B(n1577), .Z(n1579) );
  XOR U1456 ( .A(n1580), .B(n1581), .Z(n1577) );
  AND U1457 ( .A(n419), .B(n1582), .Z(n1581) );
  XNOR U1458 ( .A(p_input[1670]), .B(n1580), .Z(n1582) );
  XOR U1459 ( .A(n1583), .B(n1584), .Z(n1580) );
  AND U1460 ( .A(n423), .B(n1585), .Z(n1584) );
  XNOR U1461 ( .A(p_input[1686]), .B(n1583), .Z(n1585) );
  XOR U1462 ( .A(n1586), .B(n1587), .Z(n1583) );
  AND U1463 ( .A(n427), .B(n1588), .Z(n1587) );
  XNOR U1464 ( .A(p_input[1702]), .B(n1586), .Z(n1588) );
  XOR U1465 ( .A(n1589), .B(n1590), .Z(n1586) );
  AND U1466 ( .A(n431), .B(n1591), .Z(n1590) );
  XNOR U1467 ( .A(p_input[1718]), .B(n1589), .Z(n1591) );
  XOR U1468 ( .A(n1592), .B(n1593), .Z(n1589) );
  AND U1469 ( .A(n435), .B(n1594), .Z(n1593) );
  XNOR U1470 ( .A(p_input[1734]), .B(n1592), .Z(n1594) );
  XOR U1471 ( .A(n1595), .B(n1596), .Z(n1592) );
  AND U1472 ( .A(n439), .B(n1597), .Z(n1596) );
  XNOR U1473 ( .A(p_input[1750]), .B(n1595), .Z(n1597) );
  XOR U1474 ( .A(n1598), .B(n1599), .Z(n1595) );
  AND U1475 ( .A(n443), .B(n1600), .Z(n1599) );
  XNOR U1476 ( .A(p_input[1766]), .B(n1598), .Z(n1600) );
  XOR U1477 ( .A(n1601), .B(n1602), .Z(n1598) );
  AND U1478 ( .A(n447), .B(n1603), .Z(n1602) );
  XNOR U1479 ( .A(p_input[1782]), .B(n1601), .Z(n1603) );
  XOR U1480 ( .A(n1604), .B(n1605), .Z(n1601) );
  AND U1481 ( .A(n451), .B(n1606), .Z(n1605) );
  XNOR U1482 ( .A(p_input[1798]), .B(n1604), .Z(n1606) );
  XOR U1483 ( .A(n1607), .B(n1608), .Z(n1604) );
  AND U1484 ( .A(n455), .B(n1609), .Z(n1608) );
  XNOR U1485 ( .A(p_input[1814]), .B(n1607), .Z(n1609) );
  XOR U1486 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U1487 ( .A(n459), .B(n1612), .Z(n1611) );
  XNOR U1488 ( .A(p_input[1830]), .B(n1610), .Z(n1612) );
  XOR U1489 ( .A(n1613), .B(n1614), .Z(n1610) );
  AND U1490 ( .A(n463), .B(n1615), .Z(n1614) );
  XNOR U1491 ( .A(p_input[1846]), .B(n1613), .Z(n1615) );
  XOR U1492 ( .A(n1616), .B(n1617), .Z(n1613) );
  AND U1493 ( .A(n467), .B(n1618), .Z(n1617) );
  XNOR U1494 ( .A(p_input[1862]), .B(n1616), .Z(n1618) );
  XOR U1495 ( .A(n1619), .B(n1620), .Z(n1616) );
  AND U1496 ( .A(n471), .B(n1621), .Z(n1620) );
  XNOR U1497 ( .A(p_input[1878]), .B(n1619), .Z(n1621) );
  XOR U1498 ( .A(n1622), .B(n1623), .Z(n1619) );
  AND U1499 ( .A(n475), .B(n1624), .Z(n1623) );
  XNOR U1500 ( .A(p_input[1894]), .B(n1622), .Z(n1624) );
  XOR U1501 ( .A(n1625), .B(n1626), .Z(n1622) );
  AND U1502 ( .A(n479), .B(n1627), .Z(n1626) );
  XNOR U1503 ( .A(p_input[1910]), .B(n1625), .Z(n1627) );
  XOR U1504 ( .A(n1628), .B(n1629), .Z(n1625) );
  AND U1505 ( .A(n483), .B(n1630), .Z(n1629) );
  XNOR U1506 ( .A(p_input[1926]), .B(n1628), .Z(n1630) );
  XOR U1507 ( .A(n1631), .B(n1632), .Z(n1628) );
  AND U1508 ( .A(n487), .B(n1633), .Z(n1632) );
  XNOR U1509 ( .A(p_input[1942]), .B(n1631), .Z(n1633) );
  XOR U1510 ( .A(n1634), .B(n1635), .Z(n1631) );
  AND U1511 ( .A(n491), .B(n1636), .Z(n1635) );
  XNOR U1512 ( .A(p_input[1958]), .B(n1634), .Z(n1636) );
  XOR U1513 ( .A(n1637), .B(n1638), .Z(n1634) );
  AND U1514 ( .A(n495), .B(n1639), .Z(n1638) );
  XNOR U1515 ( .A(p_input[1974]), .B(n1637), .Z(n1639) );
  XOR U1516 ( .A(n1640), .B(n1641), .Z(n1637) );
  AND U1517 ( .A(n499), .B(n1642), .Z(n1641) );
  XNOR U1518 ( .A(p_input[1990]), .B(n1640), .Z(n1642) );
  XNOR U1519 ( .A(n1643), .B(n1644), .Z(n1640) );
  AND U1520 ( .A(n503), .B(n1645), .Z(n1644) );
  XOR U1521 ( .A(p_input[2006]), .B(n1643), .Z(n1645) );
  XOR U1522 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n1646), .Z(n1643) );
  AND U1523 ( .A(n506), .B(n1647), .Z(n1646) );
  XOR U1524 ( .A(p_input[2022]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n1647)
         );
  XNOR U1525 ( .A(n1648), .B(n1649), .Z(o[5]) );
  AND U1526 ( .A(n3), .B(n1650), .Z(n1648) );
  XNOR U1527 ( .A(p_input[5]), .B(n1649), .Z(n1650) );
  XOR U1528 ( .A(n1651), .B(n1652), .Z(n1649) );
  AND U1529 ( .A(n7), .B(n1653), .Z(n1652) );
  XNOR U1530 ( .A(p_input[21]), .B(n1651), .Z(n1653) );
  XOR U1531 ( .A(n1654), .B(n1655), .Z(n1651) );
  AND U1532 ( .A(n11), .B(n1656), .Z(n1655) );
  XNOR U1533 ( .A(p_input[37]), .B(n1654), .Z(n1656) );
  XOR U1534 ( .A(n1657), .B(n1658), .Z(n1654) );
  AND U1535 ( .A(n15), .B(n1659), .Z(n1658) );
  XNOR U1536 ( .A(p_input[53]), .B(n1657), .Z(n1659) );
  XOR U1537 ( .A(n1660), .B(n1661), .Z(n1657) );
  AND U1538 ( .A(n19), .B(n1662), .Z(n1661) );
  XNOR U1539 ( .A(p_input[69]), .B(n1660), .Z(n1662) );
  XOR U1540 ( .A(n1663), .B(n1664), .Z(n1660) );
  AND U1541 ( .A(n23), .B(n1665), .Z(n1664) );
  XNOR U1542 ( .A(p_input[85]), .B(n1663), .Z(n1665) );
  XOR U1543 ( .A(n1666), .B(n1667), .Z(n1663) );
  AND U1544 ( .A(n27), .B(n1668), .Z(n1667) );
  XNOR U1545 ( .A(p_input[101]), .B(n1666), .Z(n1668) );
  XOR U1546 ( .A(n1669), .B(n1670), .Z(n1666) );
  AND U1547 ( .A(n31), .B(n1671), .Z(n1670) );
  XNOR U1548 ( .A(p_input[117]), .B(n1669), .Z(n1671) );
  XOR U1549 ( .A(n1672), .B(n1673), .Z(n1669) );
  AND U1550 ( .A(n35), .B(n1674), .Z(n1673) );
  XNOR U1551 ( .A(p_input[133]), .B(n1672), .Z(n1674) );
  XOR U1552 ( .A(n1675), .B(n1676), .Z(n1672) );
  AND U1553 ( .A(n39), .B(n1677), .Z(n1676) );
  XNOR U1554 ( .A(p_input[149]), .B(n1675), .Z(n1677) );
  XOR U1555 ( .A(n1678), .B(n1679), .Z(n1675) );
  AND U1556 ( .A(n43), .B(n1680), .Z(n1679) );
  XNOR U1557 ( .A(p_input[165]), .B(n1678), .Z(n1680) );
  XOR U1558 ( .A(n1681), .B(n1682), .Z(n1678) );
  AND U1559 ( .A(n47), .B(n1683), .Z(n1682) );
  XNOR U1560 ( .A(p_input[181]), .B(n1681), .Z(n1683) );
  XOR U1561 ( .A(n1684), .B(n1685), .Z(n1681) );
  AND U1562 ( .A(n51), .B(n1686), .Z(n1685) );
  XNOR U1563 ( .A(p_input[197]), .B(n1684), .Z(n1686) );
  XOR U1564 ( .A(n1687), .B(n1688), .Z(n1684) );
  AND U1565 ( .A(n55), .B(n1689), .Z(n1688) );
  XNOR U1566 ( .A(p_input[213]), .B(n1687), .Z(n1689) );
  XOR U1567 ( .A(n1690), .B(n1691), .Z(n1687) );
  AND U1568 ( .A(n59), .B(n1692), .Z(n1691) );
  XNOR U1569 ( .A(p_input[229]), .B(n1690), .Z(n1692) );
  XOR U1570 ( .A(n1693), .B(n1694), .Z(n1690) );
  AND U1571 ( .A(n63), .B(n1695), .Z(n1694) );
  XNOR U1572 ( .A(p_input[245]), .B(n1693), .Z(n1695) );
  XOR U1573 ( .A(n1696), .B(n1697), .Z(n1693) );
  AND U1574 ( .A(n67), .B(n1698), .Z(n1697) );
  XNOR U1575 ( .A(p_input[261]), .B(n1696), .Z(n1698) );
  XOR U1576 ( .A(n1699), .B(n1700), .Z(n1696) );
  AND U1577 ( .A(n71), .B(n1701), .Z(n1700) );
  XNOR U1578 ( .A(p_input[277]), .B(n1699), .Z(n1701) );
  XOR U1579 ( .A(n1702), .B(n1703), .Z(n1699) );
  AND U1580 ( .A(n75), .B(n1704), .Z(n1703) );
  XNOR U1581 ( .A(p_input[293]), .B(n1702), .Z(n1704) );
  XOR U1582 ( .A(n1705), .B(n1706), .Z(n1702) );
  AND U1583 ( .A(n79), .B(n1707), .Z(n1706) );
  XNOR U1584 ( .A(p_input[309]), .B(n1705), .Z(n1707) );
  XOR U1585 ( .A(n1708), .B(n1709), .Z(n1705) );
  AND U1586 ( .A(n83), .B(n1710), .Z(n1709) );
  XNOR U1587 ( .A(p_input[325]), .B(n1708), .Z(n1710) );
  XOR U1588 ( .A(n1711), .B(n1712), .Z(n1708) );
  AND U1589 ( .A(n87), .B(n1713), .Z(n1712) );
  XNOR U1590 ( .A(p_input[341]), .B(n1711), .Z(n1713) );
  XOR U1591 ( .A(n1714), .B(n1715), .Z(n1711) );
  AND U1592 ( .A(n91), .B(n1716), .Z(n1715) );
  XNOR U1593 ( .A(p_input[357]), .B(n1714), .Z(n1716) );
  XOR U1594 ( .A(n1717), .B(n1718), .Z(n1714) );
  AND U1595 ( .A(n95), .B(n1719), .Z(n1718) );
  XNOR U1596 ( .A(p_input[373]), .B(n1717), .Z(n1719) );
  XOR U1597 ( .A(n1720), .B(n1721), .Z(n1717) );
  AND U1598 ( .A(n99), .B(n1722), .Z(n1721) );
  XNOR U1599 ( .A(p_input[389]), .B(n1720), .Z(n1722) );
  XOR U1600 ( .A(n1723), .B(n1724), .Z(n1720) );
  AND U1601 ( .A(n103), .B(n1725), .Z(n1724) );
  XNOR U1602 ( .A(p_input[405]), .B(n1723), .Z(n1725) );
  XOR U1603 ( .A(n1726), .B(n1727), .Z(n1723) );
  AND U1604 ( .A(n107), .B(n1728), .Z(n1727) );
  XNOR U1605 ( .A(p_input[421]), .B(n1726), .Z(n1728) );
  XOR U1606 ( .A(n1729), .B(n1730), .Z(n1726) );
  AND U1607 ( .A(n111), .B(n1731), .Z(n1730) );
  XNOR U1608 ( .A(p_input[437]), .B(n1729), .Z(n1731) );
  XOR U1609 ( .A(n1732), .B(n1733), .Z(n1729) );
  AND U1610 ( .A(n115), .B(n1734), .Z(n1733) );
  XNOR U1611 ( .A(p_input[453]), .B(n1732), .Z(n1734) );
  XOR U1612 ( .A(n1735), .B(n1736), .Z(n1732) );
  AND U1613 ( .A(n119), .B(n1737), .Z(n1736) );
  XNOR U1614 ( .A(p_input[469]), .B(n1735), .Z(n1737) );
  XOR U1615 ( .A(n1738), .B(n1739), .Z(n1735) );
  AND U1616 ( .A(n123), .B(n1740), .Z(n1739) );
  XNOR U1617 ( .A(p_input[485]), .B(n1738), .Z(n1740) );
  XOR U1618 ( .A(n1741), .B(n1742), .Z(n1738) );
  AND U1619 ( .A(n127), .B(n1743), .Z(n1742) );
  XNOR U1620 ( .A(p_input[501]), .B(n1741), .Z(n1743) );
  XOR U1621 ( .A(n1744), .B(n1745), .Z(n1741) );
  AND U1622 ( .A(n131), .B(n1746), .Z(n1745) );
  XNOR U1623 ( .A(p_input[517]), .B(n1744), .Z(n1746) );
  XOR U1624 ( .A(n1747), .B(n1748), .Z(n1744) );
  AND U1625 ( .A(n135), .B(n1749), .Z(n1748) );
  XNOR U1626 ( .A(p_input[533]), .B(n1747), .Z(n1749) );
  XOR U1627 ( .A(n1750), .B(n1751), .Z(n1747) );
  AND U1628 ( .A(n139), .B(n1752), .Z(n1751) );
  XNOR U1629 ( .A(p_input[549]), .B(n1750), .Z(n1752) );
  XOR U1630 ( .A(n1753), .B(n1754), .Z(n1750) );
  AND U1631 ( .A(n143), .B(n1755), .Z(n1754) );
  XNOR U1632 ( .A(p_input[565]), .B(n1753), .Z(n1755) );
  XOR U1633 ( .A(n1756), .B(n1757), .Z(n1753) );
  AND U1634 ( .A(n147), .B(n1758), .Z(n1757) );
  XNOR U1635 ( .A(p_input[581]), .B(n1756), .Z(n1758) );
  XOR U1636 ( .A(n1759), .B(n1760), .Z(n1756) );
  AND U1637 ( .A(n151), .B(n1761), .Z(n1760) );
  XNOR U1638 ( .A(p_input[597]), .B(n1759), .Z(n1761) );
  XOR U1639 ( .A(n1762), .B(n1763), .Z(n1759) );
  AND U1640 ( .A(n155), .B(n1764), .Z(n1763) );
  XNOR U1641 ( .A(p_input[613]), .B(n1762), .Z(n1764) );
  XOR U1642 ( .A(n1765), .B(n1766), .Z(n1762) );
  AND U1643 ( .A(n159), .B(n1767), .Z(n1766) );
  XNOR U1644 ( .A(p_input[629]), .B(n1765), .Z(n1767) );
  XOR U1645 ( .A(n1768), .B(n1769), .Z(n1765) );
  AND U1646 ( .A(n163), .B(n1770), .Z(n1769) );
  XNOR U1647 ( .A(p_input[645]), .B(n1768), .Z(n1770) );
  XOR U1648 ( .A(n1771), .B(n1772), .Z(n1768) );
  AND U1649 ( .A(n167), .B(n1773), .Z(n1772) );
  XNOR U1650 ( .A(p_input[661]), .B(n1771), .Z(n1773) );
  XOR U1651 ( .A(n1774), .B(n1775), .Z(n1771) );
  AND U1652 ( .A(n171), .B(n1776), .Z(n1775) );
  XNOR U1653 ( .A(p_input[677]), .B(n1774), .Z(n1776) );
  XOR U1654 ( .A(n1777), .B(n1778), .Z(n1774) );
  AND U1655 ( .A(n175), .B(n1779), .Z(n1778) );
  XNOR U1656 ( .A(p_input[693]), .B(n1777), .Z(n1779) );
  XOR U1657 ( .A(n1780), .B(n1781), .Z(n1777) );
  AND U1658 ( .A(n179), .B(n1782), .Z(n1781) );
  XNOR U1659 ( .A(p_input[709]), .B(n1780), .Z(n1782) );
  XOR U1660 ( .A(n1783), .B(n1784), .Z(n1780) );
  AND U1661 ( .A(n183), .B(n1785), .Z(n1784) );
  XNOR U1662 ( .A(p_input[725]), .B(n1783), .Z(n1785) );
  XOR U1663 ( .A(n1786), .B(n1787), .Z(n1783) );
  AND U1664 ( .A(n187), .B(n1788), .Z(n1787) );
  XNOR U1665 ( .A(p_input[741]), .B(n1786), .Z(n1788) );
  XOR U1666 ( .A(n1789), .B(n1790), .Z(n1786) );
  AND U1667 ( .A(n191), .B(n1791), .Z(n1790) );
  XNOR U1668 ( .A(p_input[757]), .B(n1789), .Z(n1791) );
  XOR U1669 ( .A(n1792), .B(n1793), .Z(n1789) );
  AND U1670 ( .A(n195), .B(n1794), .Z(n1793) );
  XNOR U1671 ( .A(p_input[773]), .B(n1792), .Z(n1794) );
  XOR U1672 ( .A(n1795), .B(n1796), .Z(n1792) );
  AND U1673 ( .A(n199), .B(n1797), .Z(n1796) );
  XNOR U1674 ( .A(p_input[789]), .B(n1795), .Z(n1797) );
  XOR U1675 ( .A(n1798), .B(n1799), .Z(n1795) );
  AND U1676 ( .A(n203), .B(n1800), .Z(n1799) );
  XNOR U1677 ( .A(p_input[805]), .B(n1798), .Z(n1800) );
  XOR U1678 ( .A(n1801), .B(n1802), .Z(n1798) );
  AND U1679 ( .A(n207), .B(n1803), .Z(n1802) );
  XNOR U1680 ( .A(p_input[821]), .B(n1801), .Z(n1803) );
  XOR U1681 ( .A(n1804), .B(n1805), .Z(n1801) );
  AND U1682 ( .A(n211), .B(n1806), .Z(n1805) );
  XNOR U1683 ( .A(p_input[837]), .B(n1804), .Z(n1806) );
  XOR U1684 ( .A(n1807), .B(n1808), .Z(n1804) );
  AND U1685 ( .A(n215), .B(n1809), .Z(n1808) );
  XNOR U1686 ( .A(p_input[853]), .B(n1807), .Z(n1809) );
  XOR U1687 ( .A(n1810), .B(n1811), .Z(n1807) );
  AND U1688 ( .A(n219), .B(n1812), .Z(n1811) );
  XNOR U1689 ( .A(p_input[869]), .B(n1810), .Z(n1812) );
  XOR U1690 ( .A(n1813), .B(n1814), .Z(n1810) );
  AND U1691 ( .A(n223), .B(n1815), .Z(n1814) );
  XNOR U1692 ( .A(p_input[885]), .B(n1813), .Z(n1815) );
  XOR U1693 ( .A(n1816), .B(n1817), .Z(n1813) );
  AND U1694 ( .A(n227), .B(n1818), .Z(n1817) );
  XNOR U1695 ( .A(p_input[901]), .B(n1816), .Z(n1818) );
  XOR U1696 ( .A(n1819), .B(n1820), .Z(n1816) );
  AND U1697 ( .A(n231), .B(n1821), .Z(n1820) );
  XNOR U1698 ( .A(p_input[917]), .B(n1819), .Z(n1821) );
  XOR U1699 ( .A(n1822), .B(n1823), .Z(n1819) );
  AND U1700 ( .A(n235), .B(n1824), .Z(n1823) );
  XNOR U1701 ( .A(p_input[933]), .B(n1822), .Z(n1824) );
  XOR U1702 ( .A(n1825), .B(n1826), .Z(n1822) );
  AND U1703 ( .A(n239), .B(n1827), .Z(n1826) );
  XNOR U1704 ( .A(p_input[949]), .B(n1825), .Z(n1827) );
  XOR U1705 ( .A(n1828), .B(n1829), .Z(n1825) );
  AND U1706 ( .A(n243), .B(n1830), .Z(n1829) );
  XNOR U1707 ( .A(p_input[965]), .B(n1828), .Z(n1830) );
  XOR U1708 ( .A(n1831), .B(n1832), .Z(n1828) );
  AND U1709 ( .A(n247), .B(n1833), .Z(n1832) );
  XNOR U1710 ( .A(p_input[981]), .B(n1831), .Z(n1833) );
  XOR U1711 ( .A(n1834), .B(n1835), .Z(n1831) );
  AND U1712 ( .A(n251), .B(n1836), .Z(n1835) );
  XNOR U1713 ( .A(p_input[997]), .B(n1834), .Z(n1836) );
  XOR U1714 ( .A(n1837), .B(n1838), .Z(n1834) );
  AND U1715 ( .A(n255), .B(n1839), .Z(n1838) );
  XNOR U1716 ( .A(p_input[1013]), .B(n1837), .Z(n1839) );
  XOR U1717 ( .A(n1840), .B(n1841), .Z(n1837) );
  AND U1718 ( .A(n259), .B(n1842), .Z(n1841) );
  XNOR U1719 ( .A(p_input[1029]), .B(n1840), .Z(n1842) );
  XOR U1720 ( .A(n1843), .B(n1844), .Z(n1840) );
  AND U1721 ( .A(n263), .B(n1845), .Z(n1844) );
  XNOR U1722 ( .A(p_input[1045]), .B(n1843), .Z(n1845) );
  XOR U1723 ( .A(n1846), .B(n1847), .Z(n1843) );
  AND U1724 ( .A(n267), .B(n1848), .Z(n1847) );
  XNOR U1725 ( .A(p_input[1061]), .B(n1846), .Z(n1848) );
  XOR U1726 ( .A(n1849), .B(n1850), .Z(n1846) );
  AND U1727 ( .A(n271), .B(n1851), .Z(n1850) );
  XNOR U1728 ( .A(p_input[1077]), .B(n1849), .Z(n1851) );
  XOR U1729 ( .A(n1852), .B(n1853), .Z(n1849) );
  AND U1730 ( .A(n275), .B(n1854), .Z(n1853) );
  XNOR U1731 ( .A(p_input[1093]), .B(n1852), .Z(n1854) );
  XOR U1732 ( .A(n1855), .B(n1856), .Z(n1852) );
  AND U1733 ( .A(n279), .B(n1857), .Z(n1856) );
  XNOR U1734 ( .A(p_input[1109]), .B(n1855), .Z(n1857) );
  XOR U1735 ( .A(n1858), .B(n1859), .Z(n1855) );
  AND U1736 ( .A(n283), .B(n1860), .Z(n1859) );
  XNOR U1737 ( .A(p_input[1125]), .B(n1858), .Z(n1860) );
  XOR U1738 ( .A(n1861), .B(n1862), .Z(n1858) );
  AND U1739 ( .A(n287), .B(n1863), .Z(n1862) );
  XNOR U1740 ( .A(p_input[1141]), .B(n1861), .Z(n1863) );
  XOR U1741 ( .A(n1864), .B(n1865), .Z(n1861) );
  AND U1742 ( .A(n291), .B(n1866), .Z(n1865) );
  XNOR U1743 ( .A(p_input[1157]), .B(n1864), .Z(n1866) );
  XOR U1744 ( .A(n1867), .B(n1868), .Z(n1864) );
  AND U1745 ( .A(n295), .B(n1869), .Z(n1868) );
  XNOR U1746 ( .A(p_input[1173]), .B(n1867), .Z(n1869) );
  XOR U1747 ( .A(n1870), .B(n1871), .Z(n1867) );
  AND U1748 ( .A(n299), .B(n1872), .Z(n1871) );
  XNOR U1749 ( .A(p_input[1189]), .B(n1870), .Z(n1872) );
  XOR U1750 ( .A(n1873), .B(n1874), .Z(n1870) );
  AND U1751 ( .A(n303), .B(n1875), .Z(n1874) );
  XNOR U1752 ( .A(p_input[1205]), .B(n1873), .Z(n1875) );
  XOR U1753 ( .A(n1876), .B(n1877), .Z(n1873) );
  AND U1754 ( .A(n307), .B(n1878), .Z(n1877) );
  XNOR U1755 ( .A(p_input[1221]), .B(n1876), .Z(n1878) );
  XOR U1756 ( .A(n1879), .B(n1880), .Z(n1876) );
  AND U1757 ( .A(n311), .B(n1881), .Z(n1880) );
  XNOR U1758 ( .A(p_input[1237]), .B(n1879), .Z(n1881) );
  XOR U1759 ( .A(n1882), .B(n1883), .Z(n1879) );
  AND U1760 ( .A(n315), .B(n1884), .Z(n1883) );
  XNOR U1761 ( .A(p_input[1253]), .B(n1882), .Z(n1884) );
  XOR U1762 ( .A(n1885), .B(n1886), .Z(n1882) );
  AND U1763 ( .A(n319), .B(n1887), .Z(n1886) );
  XNOR U1764 ( .A(p_input[1269]), .B(n1885), .Z(n1887) );
  XOR U1765 ( .A(n1888), .B(n1889), .Z(n1885) );
  AND U1766 ( .A(n323), .B(n1890), .Z(n1889) );
  XNOR U1767 ( .A(p_input[1285]), .B(n1888), .Z(n1890) );
  XOR U1768 ( .A(n1891), .B(n1892), .Z(n1888) );
  AND U1769 ( .A(n327), .B(n1893), .Z(n1892) );
  XNOR U1770 ( .A(p_input[1301]), .B(n1891), .Z(n1893) );
  XOR U1771 ( .A(n1894), .B(n1895), .Z(n1891) );
  AND U1772 ( .A(n331), .B(n1896), .Z(n1895) );
  XNOR U1773 ( .A(p_input[1317]), .B(n1894), .Z(n1896) );
  XOR U1774 ( .A(n1897), .B(n1898), .Z(n1894) );
  AND U1775 ( .A(n335), .B(n1899), .Z(n1898) );
  XNOR U1776 ( .A(p_input[1333]), .B(n1897), .Z(n1899) );
  XOR U1777 ( .A(n1900), .B(n1901), .Z(n1897) );
  AND U1778 ( .A(n339), .B(n1902), .Z(n1901) );
  XNOR U1779 ( .A(p_input[1349]), .B(n1900), .Z(n1902) );
  XOR U1780 ( .A(n1903), .B(n1904), .Z(n1900) );
  AND U1781 ( .A(n343), .B(n1905), .Z(n1904) );
  XNOR U1782 ( .A(p_input[1365]), .B(n1903), .Z(n1905) );
  XOR U1783 ( .A(n1906), .B(n1907), .Z(n1903) );
  AND U1784 ( .A(n347), .B(n1908), .Z(n1907) );
  XNOR U1785 ( .A(p_input[1381]), .B(n1906), .Z(n1908) );
  XOR U1786 ( .A(n1909), .B(n1910), .Z(n1906) );
  AND U1787 ( .A(n351), .B(n1911), .Z(n1910) );
  XNOR U1788 ( .A(p_input[1397]), .B(n1909), .Z(n1911) );
  XOR U1789 ( .A(n1912), .B(n1913), .Z(n1909) );
  AND U1790 ( .A(n355), .B(n1914), .Z(n1913) );
  XNOR U1791 ( .A(p_input[1413]), .B(n1912), .Z(n1914) );
  XOR U1792 ( .A(n1915), .B(n1916), .Z(n1912) );
  AND U1793 ( .A(n359), .B(n1917), .Z(n1916) );
  XNOR U1794 ( .A(p_input[1429]), .B(n1915), .Z(n1917) );
  XOR U1795 ( .A(n1918), .B(n1919), .Z(n1915) );
  AND U1796 ( .A(n363), .B(n1920), .Z(n1919) );
  XNOR U1797 ( .A(p_input[1445]), .B(n1918), .Z(n1920) );
  XOR U1798 ( .A(n1921), .B(n1922), .Z(n1918) );
  AND U1799 ( .A(n367), .B(n1923), .Z(n1922) );
  XNOR U1800 ( .A(p_input[1461]), .B(n1921), .Z(n1923) );
  XOR U1801 ( .A(n1924), .B(n1925), .Z(n1921) );
  AND U1802 ( .A(n371), .B(n1926), .Z(n1925) );
  XNOR U1803 ( .A(p_input[1477]), .B(n1924), .Z(n1926) );
  XOR U1804 ( .A(n1927), .B(n1928), .Z(n1924) );
  AND U1805 ( .A(n375), .B(n1929), .Z(n1928) );
  XNOR U1806 ( .A(p_input[1493]), .B(n1927), .Z(n1929) );
  XOR U1807 ( .A(n1930), .B(n1931), .Z(n1927) );
  AND U1808 ( .A(n379), .B(n1932), .Z(n1931) );
  XNOR U1809 ( .A(p_input[1509]), .B(n1930), .Z(n1932) );
  XOR U1810 ( .A(n1933), .B(n1934), .Z(n1930) );
  AND U1811 ( .A(n383), .B(n1935), .Z(n1934) );
  XNOR U1812 ( .A(p_input[1525]), .B(n1933), .Z(n1935) );
  XOR U1813 ( .A(n1936), .B(n1937), .Z(n1933) );
  AND U1814 ( .A(n387), .B(n1938), .Z(n1937) );
  XNOR U1815 ( .A(p_input[1541]), .B(n1936), .Z(n1938) );
  XOR U1816 ( .A(n1939), .B(n1940), .Z(n1936) );
  AND U1817 ( .A(n391), .B(n1941), .Z(n1940) );
  XNOR U1818 ( .A(p_input[1557]), .B(n1939), .Z(n1941) );
  XOR U1819 ( .A(n1942), .B(n1943), .Z(n1939) );
  AND U1820 ( .A(n395), .B(n1944), .Z(n1943) );
  XNOR U1821 ( .A(p_input[1573]), .B(n1942), .Z(n1944) );
  XOR U1822 ( .A(n1945), .B(n1946), .Z(n1942) );
  AND U1823 ( .A(n399), .B(n1947), .Z(n1946) );
  XNOR U1824 ( .A(p_input[1589]), .B(n1945), .Z(n1947) );
  XOR U1825 ( .A(n1948), .B(n1949), .Z(n1945) );
  AND U1826 ( .A(n403), .B(n1950), .Z(n1949) );
  XNOR U1827 ( .A(p_input[1605]), .B(n1948), .Z(n1950) );
  XOR U1828 ( .A(n1951), .B(n1952), .Z(n1948) );
  AND U1829 ( .A(n407), .B(n1953), .Z(n1952) );
  XNOR U1830 ( .A(p_input[1621]), .B(n1951), .Z(n1953) );
  XOR U1831 ( .A(n1954), .B(n1955), .Z(n1951) );
  AND U1832 ( .A(n411), .B(n1956), .Z(n1955) );
  XNOR U1833 ( .A(p_input[1637]), .B(n1954), .Z(n1956) );
  XOR U1834 ( .A(n1957), .B(n1958), .Z(n1954) );
  AND U1835 ( .A(n415), .B(n1959), .Z(n1958) );
  XNOR U1836 ( .A(p_input[1653]), .B(n1957), .Z(n1959) );
  XOR U1837 ( .A(n1960), .B(n1961), .Z(n1957) );
  AND U1838 ( .A(n419), .B(n1962), .Z(n1961) );
  XNOR U1839 ( .A(p_input[1669]), .B(n1960), .Z(n1962) );
  XOR U1840 ( .A(n1963), .B(n1964), .Z(n1960) );
  AND U1841 ( .A(n423), .B(n1965), .Z(n1964) );
  XNOR U1842 ( .A(p_input[1685]), .B(n1963), .Z(n1965) );
  XOR U1843 ( .A(n1966), .B(n1967), .Z(n1963) );
  AND U1844 ( .A(n427), .B(n1968), .Z(n1967) );
  XNOR U1845 ( .A(p_input[1701]), .B(n1966), .Z(n1968) );
  XOR U1846 ( .A(n1969), .B(n1970), .Z(n1966) );
  AND U1847 ( .A(n431), .B(n1971), .Z(n1970) );
  XNOR U1848 ( .A(p_input[1717]), .B(n1969), .Z(n1971) );
  XOR U1849 ( .A(n1972), .B(n1973), .Z(n1969) );
  AND U1850 ( .A(n435), .B(n1974), .Z(n1973) );
  XNOR U1851 ( .A(p_input[1733]), .B(n1972), .Z(n1974) );
  XOR U1852 ( .A(n1975), .B(n1976), .Z(n1972) );
  AND U1853 ( .A(n439), .B(n1977), .Z(n1976) );
  XNOR U1854 ( .A(p_input[1749]), .B(n1975), .Z(n1977) );
  XOR U1855 ( .A(n1978), .B(n1979), .Z(n1975) );
  AND U1856 ( .A(n443), .B(n1980), .Z(n1979) );
  XNOR U1857 ( .A(p_input[1765]), .B(n1978), .Z(n1980) );
  XOR U1858 ( .A(n1981), .B(n1982), .Z(n1978) );
  AND U1859 ( .A(n447), .B(n1983), .Z(n1982) );
  XNOR U1860 ( .A(p_input[1781]), .B(n1981), .Z(n1983) );
  XOR U1861 ( .A(n1984), .B(n1985), .Z(n1981) );
  AND U1862 ( .A(n451), .B(n1986), .Z(n1985) );
  XNOR U1863 ( .A(p_input[1797]), .B(n1984), .Z(n1986) );
  XOR U1864 ( .A(n1987), .B(n1988), .Z(n1984) );
  AND U1865 ( .A(n455), .B(n1989), .Z(n1988) );
  XNOR U1866 ( .A(p_input[1813]), .B(n1987), .Z(n1989) );
  XOR U1867 ( .A(n1990), .B(n1991), .Z(n1987) );
  AND U1868 ( .A(n459), .B(n1992), .Z(n1991) );
  XNOR U1869 ( .A(p_input[1829]), .B(n1990), .Z(n1992) );
  XOR U1870 ( .A(n1993), .B(n1994), .Z(n1990) );
  AND U1871 ( .A(n463), .B(n1995), .Z(n1994) );
  XNOR U1872 ( .A(p_input[1845]), .B(n1993), .Z(n1995) );
  XOR U1873 ( .A(n1996), .B(n1997), .Z(n1993) );
  AND U1874 ( .A(n467), .B(n1998), .Z(n1997) );
  XNOR U1875 ( .A(p_input[1861]), .B(n1996), .Z(n1998) );
  XOR U1876 ( .A(n1999), .B(n2000), .Z(n1996) );
  AND U1877 ( .A(n471), .B(n2001), .Z(n2000) );
  XNOR U1878 ( .A(p_input[1877]), .B(n1999), .Z(n2001) );
  XOR U1879 ( .A(n2002), .B(n2003), .Z(n1999) );
  AND U1880 ( .A(n475), .B(n2004), .Z(n2003) );
  XNOR U1881 ( .A(p_input[1893]), .B(n2002), .Z(n2004) );
  XOR U1882 ( .A(n2005), .B(n2006), .Z(n2002) );
  AND U1883 ( .A(n479), .B(n2007), .Z(n2006) );
  XNOR U1884 ( .A(p_input[1909]), .B(n2005), .Z(n2007) );
  XOR U1885 ( .A(n2008), .B(n2009), .Z(n2005) );
  AND U1886 ( .A(n483), .B(n2010), .Z(n2009) );
  XNOR U1887 ( .A(p_input[1925]), .B(n2008), .Z(n2010) );
  XOR U1888 ( .A(n2011), .B(n2012), .Z(n2008) );
  AND U1889 ( .A(n487), .B(n2013), .Z(n2012) );
  XNOR U1890 ( .A(p_input[1941]), .B(n2011), .Z(n2013) );
  XOR U1891 ( .A(n2014), .B(n2015), .Z(n2011) );
  AND U1892 ( .A(n491), .B(n2016), .Z(n2015) );
  XNOR U1893 ( .A(p_input[1957]), .B(n2014), .Z(n2016) );
  XOR U1894 ( .A(n2017), .B(n2018), .Z(n2014) );
  AND U1895 ( .A(n495), .B(n2019), .Z(n2018) );
  XNOR U1896 ( .A(p_input[1973]), .B(n2017), .Z(n2019) );
  XOR U1897 ( .A(n2020), .B(n2021), .Z(n2017) );
  AND U1898 ( .A(n499), .B(n2022), .Z(n2021) );
  XNOR U1899 ( .A(p_input[1989]), .B(n2020), .Z(n2022) );
  XNOR U1900 ( .A(n2023), .B(n2024), .Z(n2020) );
  AND U1901 ( .A(n503), .B(n2025), .Z(n2024) );
  XOR U1902 ( .A(p_input[2005]), .B(n2023), .Z(n2025) );
  XOR U1903 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n2026), .Z(n2023) );
  AND U1904 ( .A(n506), .B(n2027), .Z(n2026) );
  XOR U1905 ( .A(p_input[2021]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n2027)
         );
  XNOR U1906 ( .A(n2028), .B(n2029), .Z(o[4]) );
  AND U1907 ( .A(n3), .B(n2030), .Z(n2028) );
  XNOR U1908 ( .A(p_input[4]), .B(n2029), .Z(n2030) );
  XOR U1909 ( .A(n2031), .B(n2032), .Z(n2029) );
  AND U1910 ( .A(n7), .B(n2033), .Z(n2032) );
  XNOR U1911 ( .A(p_input[20]), .B(n2031), .Z(n2033) );
  XOR U1912 ( .A(n2034), .B(n2035), .Z(n2031) );
  AND U1913 ( .A(n11), .B(n2036), .Z(n2035) );
  XNOR U1914 ( .A(p_input[36]), .B(n2034), .Z(n2036) );
  XOR U1915 ( .A(n2037), .B(n2038), .Z(n2034) );
  AND U1916 ( .A(n15), .B(n2039), .Z(n2038) );
  XNOR U1917 ( .A(p_input[52]), .B(n2037), .Z(n2039) );
  XOR U1918 ( .A(n2040), .B(n2041), .Z(n2037) );
  AND U1919 ( .A(n19), .B(n2042), .Z(n2041) );
  XNOR U1920 ( .A(p_input[68]), .B(n2040), .Z(n2042) );
  XOR U1921 ( .A(n2043), .B(n2044), .Z(n2040) );
  AND U1922 ( .A(n23), .B(n2045), .Z(n2044) );
  XNOR U1923 ( .A(p_input[84]), .B(n2043), .Z(n2045) );
  XOR U1924 ( .A(n2046), .B(n2047), .Z(n2043) );
  AND U1925 ( .A(n27), .B(n2048), .Z(n2047) );
  XNOR U1926 ( .A(p_input[100]), .B(n2046), .Z(n2048) );
  XOR U1927 ( .A(n2049), .B(n2050), .Z(n2046) );
  AND U1928 ( .A(n31), .B(n2051), .Z(n2050) );
  XNOR U1929 ( .A(p_input[116]), .B(n2049), .Z(n2051) );
  XOR U1930 ( .A(n2052), .B(n2053), .Z(n2049) );
  AND U1931 ( .A(n35), .B(n2054), .Z(n2053) );
  XNOR U1932 ( .A(p_input[132]), .B(n2052), .Z(n2054) );
  XOR U1933 ( .A(n2055), .B(n2056), .Z(n2052) );
  AND U1934 ( .A(n39), .B(n2057), .Z(n2056) );
  XNOR U1935 ( .A(p_input[148]), .B(n2055), .Z(n2057) );
  XOR U1936 ( .A(n2058), .B(n2059), .Z(n2055) );
  AND U1937 ( .A(n43), .B(n2060), .Z(n2059) );
  XNOR U1938 ( .A(p_input[164]), .B(n2058), .Z(n2060) );
  XOR U1939 ( .A(n2061), .B(n2062), .Z(n2058) );
  AND U1940 ( .A(n47), .B(n2063), .Z(n2062) );
  XNOR U1941 ( .A(p_input[180]), .B(n2061), .Z(n2063) );
  XOR U1942 ( .A(n2064), .B(n2065), .Z(n2061) );
  AND U1943 ( .A(n51), .B(n2066), .Z(n2065) );
  XNOR U1944 ( .A(p_input[196]), .B(n2064), .Z(n2066) );
  XOR U1945 ( .A(n2067), .B(n2068), .Z(n2064) );
  AND U1946 ( .A(n55), .B(n2069), .Z(n2068) );
  XNOR U1947 ( .A(p_input[212]), .B(n2067), .Z(n2069) );
  XOR U1948 ( .A(n2070), .B(n2071), .Z(n2067) );
  AND U1949 ( .A(n59), .B(n2072), .Z(n2071) );
  XNOR U1950 ( .A(p_input[228]), .B(n2070), .Z(n2072) );
  XOR U1951 ( .A(n2073), .B(n2074), .Z(n2070) );
  AND U1952 ( .A(n63), .B(n2075), .Z(n2074) );
  XNOR U1953 ( .A(p_input[244]), .B(n2073), .Z(n2075) );
  XOR U1954 ( .A(n2076), .B(n2077), .Z(n2073) );
  AND U1955 ( .A(n67), .B(n2078), .Z(n2077) );
  XNOR U1956 ( .A(p_input[260]), .B(n2076), .Z(n2078) );
  XOR U1957 ( .A(n2079), .B(n2080), .Z(n2076) );
  AND U1958 ( .A(n71), .B(n2081), .Z(n2080) );
  XNOR U1959 ( .A(p_input[276]), .B(n2079), .Z(n2081) );
  XOR U1960 ( .A(n2082), .B(n2083), .Z(n2079) );
  AND U1961 ( .A(n75), .B(n2084), .Z(n2083) );
  XNOR U1962 ( .A(p_input[292]), .B(n2082), .Z(n2084) );
  XOR U1963 ( .A(n2085), .B(n2086), .Z(n2082) );
  AND U1964 ( .A(n79), .B(n2087), .Z(n2086) );
  XNOR U1965 ( .A(p_input[308]), .B(n2085), .Z(n2087) );
  XOR U1966 ( .A(n2088), .B(n2089), .Z(n2085) );
  AND U1967 ( .A(n83), .B(n2090), .Z(n2089) );
  XNOR U1968 ( .A(p_input[324]), .B(n2088), .Z(n2090) );
  XOR U1969 ( .A(n2091), .B(n2092), .Z(n2088) );
  AND U1970 ( .A(n87), .B(n2093), .Z(n2092) );
  XNOR U1971 ( .A(p_input[340]), .B(n2091), .Z(n2093) );
  XOR U1972 ( .A(n2094), .B(n2095), .Z(n2091) );
  AND U1973 ( .A(n91), .B(n2096), .Z(n2095) );
  XNOR U1974 ( .A(p_input[356]), .B(n2094), .Z(n2096) );
  XOR U1975 ( .A(n2097), .B(n2098), .Z(n2094) );
  AND U1976 ( .A(n95), .B(n2099), .Z(n2098) );
  XNOR U1977 ( .A(p_input[372]), .B(n2097), .Z(n2099) );
  XOR U1978 ( .A(n2100), .B(n2101), .Z(n2097) );
  AND U1979 ( .A(n99), .B(n2102), .Z(n2101) );
  XNOR U1980 ( .A(p_input[388]), .B(n2100), .Z(n2102) );
  XOR U1981 ( .A(n2103), .B(n2104), .Z(n2100) );
  AND U1982 ( .A(n103), .B(n2105), .Z(n2104) );
  XNOR U1983 ( .A(p_input[404]), .B(n2103), .Z(n2105) );
  XOR U1984 ( .A(n2106), .B(n2107), .Z(n2103) );
  AND U1985 ( .A(n107), .B(n2108), .Z(n2107) );
  XNOR U1986 ( .A(p_input[420]), .B(n2106), .Z(n2108) );
  XOR U1987 ( .A(n2109), .B(n2110), .Z(n2106) );
  AND U1988 ( .A(n111), .B(n2111), .Z(n2110) );
  XNOR U1989 ( .A(p_input[436]), .B(n2109), .Z(n2111) );
  XOR U1990 ( .A(n2112), .B(n2113), .Z(n2109) );
  AND U1991 ( .A(n115), .B(n2114), .Z(n2113) );
  XNOR U1992 ( .A(p_input[452]), .B(n2112), .Z(n2114) );
  XOR U1993 ( .A(n2115), .B(n2116), .Z(n2112) );
  AND U1994 ( .A(n119), .B(n2117), .Z(n2116) );
  XNOR U1995 ( .A(p_input[468]), .B(n2115), .Z(n2117) );
  XOR U1996 ( .A(n2118), .B(n2119), .Z(n2115) );
  AND U1997 ( .A(n123), .B(n2120), .Z(n2119) );
  XNOR U1998 ( .A(p_input[484]), .B(n2118), .Z(n2120) );
  XOR U1999 ( .A(n2121), .B(n2122), .Z(n2118) );
  AND U2000 ( .A(n127), .B(n2123), .Z(n2122) );
  XNOR U2001 ( .A(p_input[500]), .B(n2121), .Z(n2123) );
  XOR U2002 ( .A(n2124), .B(n2125), .Z(n2121) );
  AND U2003 ( .A(n131), .B(n2126), .Z(n2125) );
  XNOR U2004 ( .A(p_input[516]), .B(n2124), .Z(n2126) );
  XOR U2005 ( .A(n2127), .B(n2128), .Z(n2124) );
  AND U2006 ( .A(n135), .B(n2129), .Z(n2128) );
  XNOR U2007 ( .A(p_input[532]), .B(n2127), .Z(n2129) );
  XOR U2008 ( .A(n2130), .B(n2131), .Z(n2127) );
  AND U2009 ( .A(n139), .B(n2132), .Z(n2131) );
  XNOR U2010 ( .A(p_input[548]), .B(n2130), .Z(n2132) );
  XOR U2011 ( .A(n2133), .B(n2134), .Z(n2130) );
  AND U2012 ( .A(n143), .B(n2135), .Z(n2134) );
  XNOR U2013 ( .A(p_input[564]), .B(n2133), .Z(n2135) );
  XOR U2014 ( .A(n2136), .B(n2137), .Z(n2133) );
  AND U2015 ( .A(n147), .B(n2138), .Z(n2137) );
  XNOR U2016 ( .A(p_input[580]), .B(n2136), .Z(n2138) );
  XOR U2017 ( .A(n2139), .B(n2140), .Z(n2136) );
  AND U2018 ( .A(n151), .B(n2141), .Z(n2140) );
  XNOR U2019 ( .A(p_input[596]), .B(n2139), .Z(n2141) );
  XOR U2020 ( .A(n2142), .B(n2143), .Z(n2139) );
  AND U2021 ( .A(n155), .B(n2144), .Z(n2143) );
  XNOR U2022 ( .A(p_input[612]), .B(n2142), .Z(n2144) );
  XOR U2023 ( .A(n2145), .B(n2146), .Z(n2142) );
  AND U2024 ( .A(n159), .B(n2147), .Z(n2146) );
  XNOR U2025 ( .A(p_input[628]), .B(n2145), .Z(n2147) );
  XOR U2026 ( .A(n2148), .B(n2149), .Z(n2145) );
  AND U2027 ( .A(n163), .B(n2150), .Z(n2149) );
  XNOR U2028 ( .A(p_input[644]), .B(n2148), .Z(n2150) );
  XOR U2029 ( .A(n2151), .B(n2152), .Z(n2148) );
  AND U2030 ( .A(n167), .B(n2153), .Z(n2152) );
  XNOR U2031 ( .A(p_input[660]), .B(n2151), .Z(n2153) );
  XOR U2032 ( .A(n2154), .B(n2155), .Z(n2151) );
  AND U2033 ( .A(n171), .B(n2156), .Z(n2155) );
  XNOR U2034 ( .A(p_input[676]), .B(n2154), .Z(n2156) );
  XOR U2035 ( .A(n2157), .B(n2158), .Z(n2154) );
  AND U2036 ( .A(n175), .B(n2159), .Z(n2158) );
  XNOR U2037 ( .A(p_input[692]), .B(n2157), .Z(n2159) );
  XOR U2038 ( .A(n2160), .B(n2161), .Z(n2157) );
  AND U2039 ( .A(n179), .B(n2162), .Z(n2161) );
  XNOR U2040 ( .A(p_input[708]), .B(n2160), .Z(n2162) );
  XOR U2041 ( .A(n2163), .B(n2164), .Z(n2160) );
  AND U2042 ( .A(n183), .B(n2165), .Z(n2164) );
  XNOR U2043 ( .A(p_input[724]), .B(n2163), .Z(n2165) );
  XOR U2044 ( .A(n2166), .B(n2167), .Z(n2163) );
  AND U2045 ( .A(n187), .B(n2168), .Z(n2167) );
  XNOR U2046 ( .A(p_input[740]), .B(n2166), .Z(n2168) );
  XOR U2047 ( .A(n2169), .B(n2170), .Z(n2166) );
  AND U2048 ( .A(n191), .B(n2171), .Z(n2170) );
  XNOR U2049 ( .A(p_input[756]), .B(n2169), .Z(n2171) );
  XOR U2050 ( .A(n2172), .B(n2173), .Z(n2169) );
  AND U2051 ( .A(n195), .B(n2174), .Z(n2173) );
  XNOR U2052 ( .A(p_input[772]), .B(n2172), .Z(n2174) );
  XOR U2053 ( .A(n2175), .B(n2176), .Z(n2172) );
  AND U2054 ( .A(n199), .B(n2177), .Z(n2176) );
  XNOR U2055 ( .A(p_input[788]), .B(n2175), .Z(n2177) );
  XOR U2056 ( .A(n2178), .B(n2179), .Z(n2175) );
  AND U2057 ( .A(n203), .B(n2180), .Z(n2179) );
  XNOR U2058 ( .A(p_input[804]), .B(n2178), .Z(n2180) );
  XOR U2059 ( .A(n2181), .B(n2182), .Z(n2178) );
  AND U2060 ( .A(n207), .B(n2183), .Z(n2182) );
  XNOR U2061 ( .A(p_input[820]), .B(n2181), .Z(n2183) );
  XOR U2062 ( .A(n2184), .B(n2185), .Z(n2181) );
  AND U2063 ( .A(n211), .B(n2186), .Z(n2185) );
  XNOR U2064 ( .A(p_input[836]), .B(n2184), .Z(n2186) );
  XOR U2065 ( .A(n2187), .B(n2188), .Z(n2184) );
  AND U2066 ( .A(n215), .B(n2189), .Z(n2188) );
  XNOR U2067 ( .A(p_input[852]), .B(n2187), .Z(n2189) );
  XOR U2068 ( .A(n2190), .B(n2191), .Z(n2187) );
  AND U2069 ( .A(n219), .B(n2192), .Z(n2191) );
  XNOR U2070 ( .A(p_input[868]), .B(n2190), .Z(n2192) );
  XOR U2071 ( .A(n2193), .B(n2194), .Z(n2190) );
  AND U2072 ( .A(n223), .B(n2195), .Z(n2194) );
  XNOR U2073 ( .A(p_input[884]), .B(n2193), .Z(n2195) );
  XOR U2074 ( .A(n2196), .B(n2197), .Z(n2193) );
  AND U2075 ( .A(n227), .B(n2198), .Z(n2197) );
  XNOR U2076 ( .A(p_input[900]), .B(n2196), .Z(n2198) );
  XOR U2077 ( .A(n2199), .B(n2200), .Z(n2196) );
  AND U2078 ( .A(n231), .B(n2201), .Z(n2200) );
  XNOR U2079 ( .A(p_input[916]), .B(n2199), .Z(n2201) );
  XOR U2080 ( .A(n2202), .B(n2203), .Z(n2199) );
  AND U2081 ( .A(n235), .B(n2204), .Z(n2203) );
  XNOR U2082 ( .A(p_input[932]), .B(n2202), .Z(n2204) );
  XOR U2083 ( .A(n2205), .B(n2206), .Z(n2202) );
  AND U2084 ( .A(n239), .B(n2207), .Z(n2206) );
  XNOR U2085 ( .A(p_input[948]), .B(n2205), .Z(n2207) );
  XOR U2086 ( .A(n2208), .B(n2209), .Z(n2205) );
  AND U2087 ( .A(n243), .B(n2210), .Z(n2209) );
  XNOR U2088 ( .A(p_input[964]), .B(n2208), .Z(n2210) );
  XOR U2089 ( .A(n2211), .B(n2212), .Z(n2208) );
  AND U2090 ( .A(n247), .B(n2213), .Z(n2212) );
  XNOR U2091 ( .A(p_input[980]), .B(n2211), .Z(n2213) );
  XOR U2092 ( .A(n2214), .B(n2215), .Z(n2211) );
  AND U2093 ( .A(n251), .B(n2216), .Z(n2215) );
  XNOR U2094 ( .A(p_input[996]), .B(n2214), .Z(n2216) );
  XOR U2095 ( .A(n2217), .B(n2218), .Z(n2214) );
  AND U2096 ( .A(n255), .B(n2219), .Z(n2218) );
  XNOR U2097 ( .A(p_input[1012]), .B(n2217), .Z(n2219) );
  XOR U2098 ( .A(n2220), .B(n2221), .Z(n2217) );
  AND U2099 ( .A(n259), .B(n2222), .Z(n2221) );
  XNOR U2100 ( .A(p_input[1028]), .B(n2220), .Z(n2222) );
  XOR U2101 ( .A(n2223), .B(n2224), .Z(n2220) );
  AND U2102 ( .A(n263), .B(n2225), .Z(n2224) );
  XNOR U2103 ( .A(p_input[1044]), .B(n2223), .Z(n2225) );
  XOR U2104 ( .A(n2226), .B(n2227), .Z(n2223) );
  AND U2105 ( .A(n267), .B(n2228), .Z(n2227) );
  XNOR U2106 ( .A(p_input[1060]), .B(n2226), .Z(n2228) );
  XOR U2107 ( .A(n2229), .B(n2230), .Z(n2226) );
  AND U2108 ( .A(n271), .B(n2231), .Z(n2230) );
  XNOR U2109 ( .A(p_input[1076]), .B(n2229), .Z(n2231) );
  XOR U2110 ( .A(n2232), .B(n2233), .Z(n2229) );
  AND U2111 ( .A(n275), .B(n2234), .Z(n2233) );
  XNOR U2112 ( .A(p_input[1092]), .B(n2232), .Z(n2234) );
  XOR U2113 ( .A(n2235), .B(n2236), .Z(n2232) );
  AND U2114 ( .A(n279), .B(n2237), .Z(n2236) );
  XNOR U2115 ( .A(p_input[1108]), .B(n2235), .Z(n2237) );
  XOR U2116 ( .A(n2238), .B(n2239), .Z(n2235) );
  AND U2117 ( .A(n283), .B(n2240), .Z(n2239) );
  XNOR U2118 ( .A(p_input[1124]), .B(n2238), .Z(n2240) );
  XOR U2119 ( .A(n2241), .B(n2242), .Z(n2238) );
  AND U2120 ( .A(n287), .B(n2243), .Z(n2242) );
  XNOR U2121 ( .A(p_input[1140]), .B(n2241), .Z(n2243) );
  XOR U2122 ( .A(n2244), .B(n2245), .Z(n2241) );
  AND U2123 ( .A(n291), .B(n2246), .Z(n2245) );
  XNOR U2124 ( .A(p_input[1156]), .B(n2244), .Z(n2246) );
  XOR U2125 ( .A(n2247), .B(n2248), .Z(n2244) );
  AND U2126 ( .A(n295), .B(n2249), .Z(n2248) );
  XNOR U2127 ( .A(p_input[1172]), .B(n2247), .Z(n2249) );
  XOR U2128 ( .A(n2250), .B(n2251), .Z(n2247) );
  AND U2129 ( .A(n299), .B(n2252), .Z(n2251) );
  XNOR U2130 ( .A(p_input[1188]), .B(n2250), .Z(n2252) );
  XOR U2131 ( .A(n2253), .B(n2254), .Z(n2250) );
  AND U2132 ( .A(n303), .B(n2255), .Z(n2254) );
  XNOR U2133 ( .A(p_input[1204]), .B(n2253), .Z(n2255) );
  XOR U2134 ( .A(n2256), .B(n2257), .Z(n2253) );
  AND U2135 ( .A(n307), .B(n2258), .Z(n2257) );
  XNOR U2136 ( .A(p_input[1220]), .B(n2256), .Z(n2258) );
  XOR U2137 ( .A(n2259), .B(n2260), .Z(n2256) );
  AND U2138 ( .A(n311), .B(n2261), .Z(n2260) );
  XNOR U2139 ( .A(p_input[1236]), .B(n2259), .Z(n2261) );
  XOR U2140 ( .A(n2262), .B(n2263), .Z(n2259) );
  AND U2141 ( .A(n315), .B(n2264), .Z(n2263) );
  XNOR U2142 ( .A(p_input[1252]), .B(n2262), .Z(n2264) );
  XOR U2143 ( .A(n2265), .B(n2266), .Z(n2262) );
  AND U2144 ( .A(n319), .B(n2267), .Z(n2266) );
  XNOR U2145 ( .A(p_input[1268]), .B(n2265), .Z(n2267) );
  XOR U2146 ( .A(n2268), .B(n2269), .Z(n2265) );
  AND U2147 ( .A(n323), .B(n2270), .Z(n2269) );
  XNOR U2148 ( .A(p_input[1284]), .B(n2268), .Z(n2270) );
  XOR U2149 ( .A(n2271), .B(n2272), .Z(n2268) );
  AND U2150 ( .A(n327), .B(n2273), .Z(n2272) );
  XNOR U2151 ( .A(p_input[1300]), .B(n2271), .Z(n2273) );
  XOR U2152 ( .A(n2274), .B(n2275), .Z(n2271) );
  AND U2153 ( .A(n331), .B(n2276), .Z(n2275) );
  XNOR U2154 ( .A(p_input[1316]), .B(n2274), .Z(n2276) );
  XOR U2155 ( .A(n2277), .B(n2278), .Z(n2274) );
  AND U2156 ( .A(n335), .B(n2279), .Z(n2278) );
  XNOR U2157 ( .A(p_input[1332]), .B(n2277), .Z(n2279) );
  XOR U2158 ( .A(n2280), .B(n2281), .Z(n2277) );
  AND U2159 ( .A(n339), .B(n2282), .Z(n2281) );
  XNOR U2160 ( .A(p_input[1348]), .B(n2280), .Z(n2282) );
  XOR U2161 ( .A(n2283), .B(n2284), .Z(n2280) );
  AND U2162 ( .A(n343), .B(n2285), .Z(n2284) );
  XNOR U2163 ( .A(p_input[1364]), .B(n2283), .Z(n2285) );
  XOR U2164 ( .A(n2286), .B(n2287), .Z(n2283) );
  AND U2165 ( .A(n347), .B(n2288), .Z(n2287) );
  XNOR U2166 ( .A(p_input[1380]), .B(n2286), .Z(n2288) );
  XOR U2167 ( .A(n2289), .B(n2290), .Z(n2286) );
  AND U2168 ( .A(n351), .B(n2291), .Z(n2290) );
  XNOR U2169 ( .A(p_input[1396]), .B(n2289), .Z(n2291) );
  XOR U2170 ( .A(n2292), .B(n2293), .Z(n2289) );
  AND U2171 ( .A(n355), .B(n2294), .Z(n2293) );
  XNOR U2172 ( .A(p_input[1412]), .B(n2292), .Z(n2294) );
  XOR U2173 ( .A(n2295), .B(n2296), .Z(n2292) );
  AND U2174 ( .A(n359), .B(n2297), .Z(n2296) );
  XNOR U2175 ( .A(p_input[1428]), .B(n2295), .Z(n2297) );
  XOR U2176 ( .A(n2298), .B(n2299), .Z(n2295) );
  AND U2177 ( .A(n363), .B(n2300), .Z(n2299) );
  XNOR U2178 ( .A(p_input[1444]), .B(n2298), .Z(n2300) );
  XOR U2179 ( .A(n2301), .B(n2302), .Z(n2298) );
  AND U2180 ( .A(n367), .B(n2303), .Z(n2302) );
  XNOR U2181 ( .A(p_input[1460]), .B(n2301), .Z(n2303) );
  XOR U2182 ( .A(n2304), .B(n2305), .Z(n2301) );
  AND U2183 ( .A(n371), .B(n2306), .Z(n2305) );
  XNOR U2184 ( .A(p_input[1476]), .B(n2304), .Z(n2306) );
  XOR U2185 ( .A(n2307), .B(n2308), .Z(n2304) );
  AND U2186 ( .A(n375), .B(n2309), .Z(n2308) );
  XNOR U2187 ( .A(p_input[1492]), .B(n2307), .Z(n2309) );
  XOR U2188 ( .A(n2310), .B(n2311), .Z(n2307) );
  AND U2189 ( .A(n379), .B(n2312), .Z(n2311) );
  XNOR U2190 ( .A(p_input[1508]), .B(n2310), .Z(n2312) );
  XOR U2191 ( .A(n2313), .B(n2314), .Z(n2310) );
  AND U2192 ( .A(n383), .B(n2315), .Z(n2314) );
  XNOR U2193 ( .A(p_input[1524]), .B(n2313), .Z(n2315) );
  XOR U2194 ( .A(n2316), .B(n2317), .Z(n2313) );
  AND U2195 ( .A(n387), .B(n2318), .Z(n2317) );
  XNOR U2196 ( .A(p_input[1540]), .B(n2316), .Z(n2318) );
  XOR U2197 ( .A(n2319), .B(n2320), .Z(n2316) );
  AND U2198 ( .A(n391), .B(n2321), .Z(n2320) );
  XNOR U2199 ( .A(p_input[1556]), .B(n2319), .Z(n2321) );
  XOR U2200 ( .A(n2322), .B(n2323), .Z(n2319) );
  AND U2201 ( .A(n395), .B(n2324), .Z(n2323) );
  XNOR U2202 ( .A(p_input[1572]), .B(n2322), .Z(n2324) );
  XOR U2203 ( .A(n2325), .B(n2326), .Z(n2322) );
  AND U2204 ( .A(n399), .B(n2327), .Z(n2326) );
  XNOR U2205 ( .A(p_input[1588]), .B(n2325), .Z(n2327) );
  XOR U2206 ( .A(n2328), .B(n2329), .Z(n2325) );
  AND U2207 ( .A(n403), .B(n2330), .Z(n2329) );
  XNOR U2208 ( .A(p_input[1604]), .B(n2328), .Z(n2330) );
  XOR U2209 ( .A(n2331), .B(n2332), .Z(n2328) );
  AND U2210 ( .A(n407), .B(n2333), .Z(n2332) );
  XNOR U2211 ( .A(p_input[1620]), .B(n2331), .Z(n2333) );
  XOR U2212 ( .A(n2334), .B(n2335), .Z(n2331) );
  AND U2213 ( .A(n411), .B(n2336), .Z(n2335) );
  XNOR U2214 ( .A(p_input[1636]), .B(n2334), .Z(n2336) );
  XOR U2215 ( .A(n2337), .B(n2338), .Z(n2334) );
  AND U2216 ( .A(n415), .B(n2339), .Z(n2338) );
  XNOR U2217 ( .A(p_input[1652]), .B(n2337), .Z(n2339) );
  XOR U2218 ( .A(n2340), .B(n2341), .Z(n2337) );
  AND U2219 ( .A(n419), .B(n2342), .Z(n2341) );
  XNOR U2220 ( .A(p_input[1668]), .B(n2340), .Z(n2342) );
  XOR U2221 ( .A(n2343), .B(n2344), .Z(n2340) );
  AND U2222 ( .A(n423), .B(n2345), .Z(n2344) );
  XNOR U2223 ( .A(p_input[1684]), .B(n2343), .Z(n2345) );
  XOR U2224 ( .A(n2346), .B(n2347), .Z(n2343) );
  AND U2225 ( .A(n427), .B(n2348), .Z(n2347) );
  XNOR U2226 ( .A(p_input[1700]), .B(n2346), .Z(n2348) );
  XOR U2227 ( .A(n2349), .B(n2350), .Z(n2346) );
  AND U2228 ( .A(n431), .B(n2351), .Z(n2350) );
  XNOR U2229 ( .A(p_input[1716]), .B(n2349), .Z(n2351) );
  XOR U2230 ( .A(n2352), .B(n2353), .Z(n2349) );
  AND U2231 ( .A(n435), .B(n2354), .Z(n2353) );
  XNOR U2232 ( .A(p_input[1732]), .B(n2352), .Z(n2354) );
  XOR U2233 ( .A(n2355), .B(n2356), .Z(n2352) );
  AND U2234 ( .A(n439), .B(n2357), .Z(n2356) );
  XNOR U2235 ( .A(p_input[1748]), .B(n2355), .Z(n2357) );
  XOR U2236 ( .A(n2358), .B(n2359), .Z(n2355) );
  AND U2237 ( .A(n443), .B(n2360), .Z(n2359) );
  XNOR U2238 ( .A(p_input[1764]), .B(n2358), .Z(n2360) );
  XOR U2239 ( .A(n2361), .B(n2362), .Z(n2358) );
  AND U2240 ( .A(n447), .B(n2363), .Z(n2362) );
  XNOR U2241 ( .A(p_input[1780]), .B(n2361), .Z(n2363) );
  XOR U2242 ( .A(n2364), .B(n2365), .Z(n2361) );
  AND U2243 ( .A(n451), .B(n2366), .Z(n2365) );
  XNOR U2244 ( .A(p_input[1796]), .B(n2364), .Z(n2366) );
  XOR U2245 ( .A(n2367), .B(n2368), .Z(n2364) );
  AND U2246 ( .A(n455), .B(n2369), .Z(n2368) );
  XNOR U2247 ( .A(p_input[1812]), .B(n2367), .Z(n2369) );
  XOR U2248 ( .A(n2370), .B(n2371), .Z(n2367) );
  AND U2249 ( .A(n459), .B(n2372), .Z(n2371) );
  XNOR U2250 ( .A(p_input[1828]), .B(n2370), .Z(n2372) );
  XOR U2251 ( .A(n2373), .B(n2374), .Z(n2370) );
  AND U2252 ( .A(n463), .B(n2375), .Z(n2374) );
  XNOR U2253 ( .A(p_input[1844]), .B(n2373), .Z(n2375) );
  XOR U2254 ( .A(n2376), .B(n2377), .Z(n2373) );
  AND U2255 ( .A(n467), .B(n2378), .Z(n2377) );
  XNOR U2256 ( .A(p_input[1860]), .B(n2376), .Z(n2378) );
  XOR U2257 ( .A(n2379), .B(n2380), .Z(n2376) );
  AND U2258 ( .A(n471), .B(n2381), .Z(n2380) );
  XNOR U2259 ( .A(p_input[1876]), .B(n2379), .Z(n2381) );
  XOR U2260 ( .A(n2382), .B(n2383), .Z(n2379) );
  AND U2261 ( .A(n475), .B(n2384), .Z(n2383) );
  XNOR U2262 ( .A(p_input[1892]), .B(n2382), .Z(n2384) );
  XOR U2263 ( .A(n2385), .B(n2386), .Z(n2382) );
  AND U2264 ( .A(n479), .B(n2387), .Z(n2386) );
  XNOR U2265 ( .A(p_input[1908]), .B(n2385), .Z(n2387) );
  XOR U2266 ( .A(n2388), .B(n2389), .Z(n2385) );
  AND U2267 ( .A(n483), .B(n2390), .Z(n2389) );
  XNOR U2268 ( .A(p_input[1924]), .B(n2388), .Z(n2390) );
  XOR U2269 ( .A(n2391), .B(n2392), .Z(n2388) );
  AND U2270 ( .A(n487), .B(n2393), .Z(n2392) );
  XNOR U2271 ( .A(p_input[1940]), .B(n2391), .Z(n2393) );
  XOR U2272 ( .A(n2394), .B(n2395), .Z(n2391) );
  AND U2273 ( .A(n491), .B(n2396), .Z(n2395) );
  XNOR U2274 ( .A(p_input[1956]), .B(n2394), .Z(n2396) );
  XOR U2275 ( .A(n2397), .B(n2398), .Z(n2394) );
  AND U2276 ( .A(n495), .B(n2399), .Z(n2398) );
  XNOR U2277 ( .A(p_input[1972]), .B(n2397), .Z(n2399) );
  XOR U2278 ( .A(n2400), .B(n2401), .Z(n2397) );
  AND U2279 ( .A(n499), .B(n2402), .Z(n2401) );
  XNOR U2280 ( .A(p_input[1988]), .B(n2400), .Z(n2402) );
  XNOR U2281 ( .A(n2403), .B(n2404), .Z(n2400) );
  AND U2282 ( .A(n503), .B(n2405), .Z(n2404) );
  XOR U2283 ( .A(p_input[2004]), .B(n2403), .Z(n2405) );
  XOR U2284 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n2406), .Z(n2403) );
  AND U2285 ( .A(n506), .B(n2407), .Z(n2406) );
  XOR U2286 ( .A(p_input[2020]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n2407)
         );
  XNOR U2287 ( .A(n2408), .B(n2409), .Z(o[3]) );
  AND U2288 ( .A(n3), .B(n2410), .Z(n2408) );
  XNOR U2289 ( .A(p_input[3]), .B(n2409), .Z(n2410) );
  XOR U2290 ( .A(n2411), .B(n2412), .Z(n2409) );
  AND U2291 ( .A(n7), .B(n2413), .Z(n2412) );
  XNOR U2292 ( .A(p_input[19]), .B(n2411), .Z(n2413) );
  XOR U2293 ( .A(n2414), .B(n2415), .Z(n2411) );
  AND U2294 ( .A(n11), .B(n2416), .Z(n2415) );
  XNOR U2295 ( .A(p_input[35]), .B(n2414), .Z(n2416) );
  XOR U2296 ( .A(n2417), .B(n2418), .Z(n2414) );
  AND U2297 ( .A(n15), .B(n2419), .Z(n2418) );
  XNOR U2298 ( .A(p_input[51]), .B(n2417), .Z(n2419) );
  XOR U2299 ( .A(n2420), .B(n2421), .Z(n2417) );
  AND U2300 ( .A(n19), .B(n2422), .Z(n2421) );
  XNOR U2301 ( .A(p_input[67]), .B(n2420), .Z(n2422) );
  XOR U2302 ( .A(n2423), .B(n2424), .Z(n2420) );
  AND U2303 ( .A(n23), .B(n2425), .Z(n2424) );
  XNOR U2304 ( .A(p_input[83]), .B(n2423), .Z(n2425) );
  XOR U2305 ( .A(n2426), .B(n2427), .Z(n2423) );
  AND U2306 ( .A(n27), .B(n2428), .Z(n2427) );
  XNOR U2307 ( .A(p_input[99]), .B(n2426), .Z(n2428) );
  XOR U2308 ( .A(n2429), .B(n2430), .Z(n2426) );
  AND U2309 ( .A(n31), .B(n2431), .Z(n2430) );
  XNOR U2310 ( .A(p_input[115]), .B(n2429), .Z(n2431) );
  XOR U2311 ( .A(n2432), .B(n2433), .Z(n2429) );
  AND U2312 ( .A(n35), .B(n2434), .Z(n2433) );
  XNOR U2313 ( .A(p_input[131]), .B(n2432), .Z(n2434) );
  XOR U2314 ( .A(n2435), .B(n2436), .Z(n2432) );
  AND U2315 ( .A(n39), .B(n2437), .Z(n2436) );
  XNOR U2316 ( .A(p_input[147]), .B(n2435), .Z(n2437) );
  XOR U2317 ( .A(n2438), .B(n2439), .Z(n2435) );
  AND U2318 ( .A(n43), .B(n2440), .Z(n2439) );
  XNOR U2319 ( .A(p_input[163]), .B(n2438), .Z(n2440) );
  XOR U2320 ( .A(n2441), .B(n2442), .Z(n2438) );
  AND U2321 ( .A(n47), .B(n2443), .Z(n2442) );
  XNOR U2322 ( .A(p_input[179]), .B(n2441), .Z(n2443) );
  XOR U2323 ( .A(n2444), .B(n2445), .Z(n2441) );
  AND U2324 ( .A(n51), .B(n2446), .Z(n2445) );
  XNOR U2325 ( .A(p_input[195]), .B(n2444), .Z(n2446) );
  XOR U2326 ( .A(n2447), .B(n2448), .Z(n2444) );
  AND U2327 ( .A(n55), .B(n2449), .Z(n2448) );
  XNOR U2328 ( .A(p_input[211]), .B(n2447), .Z(n2449) );
  XOR U2329 ( .A(n2450), .B(n2451), .Z(n2447) );
  AND U2330 ( .A(n59), .B(n2452), .Z(n2451) );
  XNOR U2331 ( .A(p_input[227]), .B(n2450), .Z(n2452) );
  XOR U2332 ( .A(n2453), .B(n2454), .Z(n2450) );
  AND U2333 ( .A(n63), .B(n2455), .Z(n2454) );
  XNOR U2334 ( .A(p_input[243]), .B(n2453), .Z(n2455) );
  XOR U2335 ( .A(n2456), .B(n2457), .Z(n2453) );
  AND U2336 ( .A(n67), .B(n2458), .Z(n2457) );
  XNOR U2337 ( .A(p_input[259]), .B(n2456), .Z(n2458) );
  XOR U2338 ( .A(n2459), .B(n2460), .Z(n2456) );
  AND U2339 ( .A(n71), .B(n2461), .Z(n2460) );
  XNOR U2340 ( .A(p_input[275]), .B(n2459), .Z(n2461) );
  XOR U2341 ( .A(n2462), .B(n2463), .Z(n2459) );
  AND U2342 ( .A(n75), .B(n2464), .Z(n2463) );
  XNOR U2343 ( .A(p_input[291]), .B(n2462), .Z(n2464) );
  XOR U2344 ( .A(n2465), .B(n2466), .Z(n2462) );
  AND U2345 ( .A(n79), .B(n2467), .Z(n2466) );
  XNOR U2346 ( .A(p_input[307]), .B(n2465), .Z(n2467) );
  XOR U2347 ( .A(n2468), .B(n2469), .Z(n2465) );
  AND U2348 ( .A(n83), .B(n2470), .Z(n2469) );
  XNOR U2349 ( .A(p_input[323]), .B(n2468), .Z(n2470) );
  XOR U2350 ( .A(n2471), .B(n2472), .Z(n2468) );
  AND U2351 ( .A(n87), .B(n2473), .Z(n2472) );
  XNOR U2352 ( .A(p_input[339]), .B(n2471), .Z(n2473) );
  XOR U2353 ( .A(n2474), .B(n2475), .Z(n2471) );
  AND U2354 ( .A(n91), .B(n2476), .Z(n2475) );
  XNOR U2355 ( .A(p_input[355]), .B(n2474), .Z(n2476) );
  XOR U2356 ( .A(n2477), .B(n2478), .Z(n2474) );
  AND U2357 ( .A(n95), .B(n2479), .Z(n2478) );
  XNOR U2358 ( .A(p_input[371]), .B(n2477), .Z(n2479) );
  XOR U2359 ( .A(n2480), .B(n2481), .Z(n2477) );
  AND U2360 ( .A(n99), .B(n2482), .Z(n2481) );
  XNOR U2361 ( .A(p_input[387]), .B(n2480), .Z(n2482) );
  XOR U2362 ( .A(n2483), .B(n2484), .Z(n2480) );
  AND U2363 ( .A(n103), .B(n2485), .Z(n2484) );
  XNOR U2364 ( .A(p_input[403]), .B(n2483), .Z(n2485) );
  XOR U2365 ( .A(n2486), .B(n2487), .Z(n2483) );
  AND U2366 ( .A(n107), .B(n2488), .Z(n2487) );
  XNOR U2367 ( .A(p_input[419]), .B(n2486), .Z(n2488) );
  XOR U2368 ( .A(n2489), .B(n2490), .Z(n2486) );
  AND U2369 ( .A(n111), .B(n2491), .Z(n2490) );
  XNOR U2370 ( .A(p_input[435]), .B(n2489), .Z(n2491) );
  XOR U2371 ( .A(n2492), .B(n2493), .Z(n2489) );
  AND U2372 ( .A(n115), .B(n2494), .Z(n2493) );
  XNOR U2373 ( .A(p_input[451]), .B(n2492), .Z(n2494) );
  XOR U2374 ( .A(n2495), .B(n2496), .Z(n2492) );
  AND U2375 ( .A(n119), .B(n2497), .Z(n2496) );
  XNOR U2376 ( .A(p_input[467]), .B(n2495), .Z(n2497) );
  XOR U2377 ( .A(n2498), .B(n2499), .Z(n2495) );
  AND U2378 ( .A(n123), .B(n2500), .Z(n2499) );
  XNOR U2379 ( .A(p_input[483]), .B(n2498), .Z(n2500) );
  XOR U2380 ( .A(n2501), .B(n2502), .Z(n2498) );
  AND U2381 ( .A(n127), .B(n2503), .Z(n2502) );
  XNOR U2382 ( .A(p_input[499]), .B(n2501), .Z(n2503) );
  XOR U2383 ( .A(n2504), .B(n2505), .Z(n2501) );
  AND U2384 ( .A(n131), .B(n2506), .Z(n2505) );
  XNOR U2385 ( .A(p_input[515]), .B(n2504), .Z(n2506) );
  XOR U2386 ( .A(n2507), .B(n2508), .Z(n2504) );
  AND U2387 ( .A(n135), .B(n2509), .Z(n2508) );
  XNOR U2388 ( .A(p_input[531]), .B(n2507), .Z(n2509) );
  XOR U2389 ( .A(n2510), .B(n2511), .Z(n2507) );
  AND U2390 ( .A(n139), .B(n2512), .Z(n2511) );
  XNOR U2391 ( .A(p_input[547]), .B(n2510), .Z(n2512) );
  XOR U2392 ( .A(n2513), .B(n2514), .Z(n2510) );
  AND U2393 ( .A(n143), .B(n2515), .Z(n2514) );
  XNOR U2394 ( .A(p_input[563]), .B(n2513), .Z(n2515) );
  XOR U2395 ( .A(n2516), .B(n2517), .Z(n2513) );
  AND U2396 ( .A(n147), .B(n2518), .Z(n2517) );
  XNOR U2397 ( .A(p_input[579]), .B(n2516), .Z(n2518) );
  XOR U2398 ( .A(n2519), .B(n2520), .Z(n2516) );
  AND U2399 ( .A(n151), .B(n2521), .Z(n2520) );
  XNOR U2400 ( .A(p_input[595]), .B(n2519), .Z(n2521) );
  XOR U2401 ( .A(n2522), .B(n2523), .Z(n2519) );
  AND U2402 ( .A(n155), .B(n2524), .Z(n2523) );
  XNOR U2403 ( .A(p_input[611]), .B(n2522), .Z(n2524) );
  XOR U2404 ( .A(n2525), .B(n2526), .Z(n2522) );
  AND U2405 ( .A(n159), .B(n2527), .Z(n2526) );
  XNOR U2406 ( .A(p_input[627]), .B(n2525), .Z(n2527) );
  XOR U2407 ( .A(n2528), .B(n2529), .Z(n2525) );
  AND U2408 ( .A(n163), .B(n2530), .Z(n2529) );
  XNOR U2409 ( .A(p_input[643]), .B(n2528), .Z(n2530) );
  XOR U2410 ( .A(n2531), .B(n2532), .Z(n2528) );
  AND U2411 ( .A(n167), .B(n2533), .Z(n2532) );
  XNOR U2412 ( .A(p_input[659]), .B(n2531), .Z(n2533) );
  XOR U2413 ( .A(n2534), .B(n2535), .Z(n2531) );
  AND U2414 ( .A(n171), .B(n2536), .Z(n2535) );
  XNOR U2415 ( .A(p_input[675]), .B(n2534), .Z(n2536) );
  XOR U2416 ( .A(n2537), .B(n2538), .Z(n2534) );
  AND U2417 ( .A(n175), .B(n2539), .Z(n2538) );
  XNOR U2418 ( .A(p_input[691]), .B(n2537), .Z(n2539) );
  XOR U2419 ( .A(n2540), .B(n2541), .Z(n2537) );
  AND U2420 ( .A(n179), .B(n2542), .Z(n2541) );
  XNOR U2421 ( .A(p_input[707]), .B(n2540), .Z(n2542) );
  XOR U2422 ( .A(n2543), .B(n2544), .Z(n2540) );
  AND U2423 ( .A(n183), .B(n2545), .Z(n2544) );
  XNOR U2424 ( .A(p_input[723]), .B(n2543), .Z(n2545) );
  XOR U2425 ( .A(n2546), .B(n2547), .Z(n2543) );
  AND U2426 ( .A(n187), .B(n2548), .Z(n2547) );
  XNOR U2427 ( .A(p_input[739]), .B(n2546), .Z(n2548) );
  XOR U2428 ( .A(n2549), .B(n2550), .Z(n2546) );
  AND U2429 ( .A(n191), .B(n2551), .Z(n2550) );
  XNOR U2430 ( .A(p_input[755]), .B(n2549), .Z(n2551) );
  XOR U2431 ( .A(n2552), .B(n2553), .Z(n2549) );
  AND U2432 ( .A(n195), .B(n2554), .Z(n2553) );
  XNOR U2433 ( .A(p_input[771]), .B(n2552), .Z(n2554) );
  XOR U2434 ( .A(n2555), .B(n2556), .Z(n2552) );
  AND U2435 ( .A(n199), .B(n2557), .Z(n2556) );
  XNOR U2436 ( .A(p_input[787]), .B(n2555), .Z(n2557) );
  XOR U2437 ( .A(n2558), .B(n2559), .Z(n2555) );
  AND U2438 ( .A(n203), .B(n2560), .Z(n2559) );
  XNOR U2439 ( .A(p_input[803]), .B(n2558), .Z(n2560) );
  XOR U2440 ( .A(n2561), .B(n2562), .Z(n2558) );
  AND U2441 ( .A(n207), .B(n2563), .Z(n2562) );
  XNOR U2442 ( .A(p_input[819]), .B(n2561), .Z(n2563) );
  XOR U2443 ( .A(n2564), .B(n2565), .Z(n2561) );
  AND U2444 ( .A(n211), .B(n2566), .Z(n2565) );
  XNOR U2445 ( .A(p_input[835]), .B(n2564), .Z(n2566) );
  XOR U2446 ( .A(n2567), .B(n2568), .Z(n2564) );
  AND U2447 ( .A(n215), .B(n2569), .Z(n2568) );
  XNOR U2448 ( .A(p_input[851]), .B(n2567), .Z(n2569) );
  XOR U2449 ( .A(n2570), .B(n2571), .Z(n2567) );
  AND U2450 ( .A(n219), .B(n2572), .Z(n2571) );
  XNOR U2451 ( .A(p_input[867]), .B(n2570), .Z(n2572) );
  XOR U2452 ( .A(n2573), .B(n2574), .Z(n2570) );
  AND U2453 ( .A(n223), .B(n2575), .Z(n2574) );
  XNOR U2454 ( .A(p_input[883]), .B(n2573), .Z(n2575) );
  XOR U2455 ( .A(n2576), .B(n2577), .Z(n2573) );
  AND U2456 ( .A(n227), .B(n2578), .Z(n2577) );
  XNOR U2457 ( .A(p_input[899]), .B(n2576), .Z(n2578) );
  XOR U2458 ( .A(n2579), .B(n2580), .Z(n2576) );
  AND U2459 ( .A(n231), .B(n2581), .Z(n2580) );
  XNOR U2460 ( .A(p_input[915]), .B(n2579), .Z(n2581) );
  XOR U2461 ( .A(n2582), .B(n2583), .Z(n2579) );
  AND U2462 ( .A(n235), .B(n2584), .Z(n2583) );
  XNOR U2463 ( .A(p_input[931]), .B(n2582), .Z(n2584) );
  XOR U2464 ( .A(n2585), .B(n2586), .Z(n2582) );
  AND U2465 ( .A(n239), .B(n2587), .Z(n2586) );
  XNOR U2466 ( .A(p_input[947]), .B(n2585), .Z(n2587) );
  XOR U2467 ( .A(n2588), .B(n2589), .Z(n2585) );
  AND U2468 ( .A(n243), .B(n2590), .Z(n2589) );
  XNOR U2469 ( .A(p_input[963]), .B(n2588), .Z(n2590) );
  XOR U2470 ( .A(n2591), .B(n2592), .Z(n2588) );
  AND U2471 ( .A(n247), .B(n2593), .Z(n2592) );
  XNOR U2472 ( .A(p_input[979]), .B(n2591), .Z(n2593) );
  XOR U2473 ( .A(n2594), .B(n2595), .Z(n2591) );
  AND U2474 ( .A(n251), .B(n2596), .Z(n2595) );
  XNOR U2475 ( .A(p_input[995]), .B(n2594), .Z(n2596) );
  XOR U2476 ( .A(n2597), .B(n2598), .Z(n2594) );
  AND U2477 ( .A(n255), .B(n2599), .Z(n2598) );
  XNOR U2478 ( .A(p_input[1011]), .B(n2597), .Z(n2599) );
  XOR U2479 ( .A(n2600), .B(n2601), .Z(n2597) );
  AND U2480 ( .A(n259), .B(n2602), .Z(n2601) );
  XNOR U2481 ( .A(p_input[1027]), .B(n2600), .Z(n2602) );
  XOR U2482 ( .A(n2603), .B(n2604), .Z(n2600) );
  AND U2483 ( .A(n263), .B(n2605), .Z(n2604) );
  XNOR U2484 ( .A(p_input[1043]), .B(n2603), .Z(n2605) );
  XOR U2485 ( .A(n2606), .B(n2607), .Z(n2603) );
  AND U2486 ( .A(n267), .B(n2608), .Z(n2607) );
  XNOR U2487 ( .A(p_input[1059]), .B(n2606), .Z(n2608) );
  XOR U2488 ( .A(n2609), .B(n2610), .Z(n2606) );
  AND U2489 ( .A(n271), .B(n2611), .Z(n2610) );
  XNOR U2490 ( .A(p_input[1075]), .B(n2609), .Z(n2611) );
  XOR U2491 ( .A(n2612), .B(n2613), .Z(n2609) );
  AND U2492 ( .A(n275), .B(n2614), .Z(n2613) );
  XNOR U2493 ( .A(p_input[1091]), .B(n2612), .Z(n2614) );
  XOR U2494 ( .A(n2615), .B(n2616), .Z(n2612) );
  AND U2495 ( .A(n279), .B(n2617), .Z(n2616) );
  XNOR U2496 ( .A(p_input[1107]), .B(n2615), .Z(n2617) );
  XOR U2497 ( .A(n2618), .B(n2619), .Z(n2615) );
  AND U2498 ( .A(n283), .B(n2620), .Z(n2619) );
  XNOR U2499 ( .A(p_input[1123]), .B(n2618), .Z(n2620) );
  XOR U2500 ( .A(n2621), .B(n2622), .Z(n2618) );
  AND U2501 ( .A(n287), .B(n2623), .Z(n2622) );
  XNOR U2502 ( .A(p_input[1139]), .B(n2621), .Z(n2623) );
  XOR U2503 ( .A(n2624), .B(n2625), .Z(n2621) );
  AND U2504 ( .A(n291), .B(n2626), .Z(n2625) );
  XNOR U2505 ( .A(p_input[1155]), .B(n2624), .Z(n2626) );
  XOR U2506 ( .A(n2627), .B(n2628), .Z(n2624) );
  AND U2507 ( .A(n295), .B(n2629), .Z(n2628) );
  XNOR U2508 ( .A(p_input[1171]), .B(n2627), .Z(n2629) );
  XOR U2509 ( .A(n2630), .B(n2631), .Z(n2627) );
  AND U2510 ( .A(n299), .B(n2632), .Z(n2631) );
  XNOR U2511 ( .A(p_input[1187]), .B(n2630), .Z(n2632) );
  XOR U2512 ( .A(n2633), .B(n2634), .Z(n2630) );
  AND U2513 ( .A(n303), .B(n2635), .Z(n2634) );
  XNOR U2514 ( .A(p_input[1203]), .B(n2633), .Z(n2635) );
  XOR U2515 ( .A(n2636), .B(n2637), .Z(n2633) );
  AND U2516 ( .A(n307), .B(n2638), .Z(n2637) );
  XNOR U2517 ( .A(p_input[1219]), .B(n2636), .Z(n2638) );
  XOR U2518 ( .A(n2639), .B(n2640), .Z(n2636) );
  AND U2519 ( .A(n311), .B(n2641), .Z(n2640) );
  XNOR U2520 ( .A(p_input[1235]), .B(n2639), .Z(n2641) );
  XOR U2521 ( .A(n2642), .B(n2643), .Z(n2639) );
  AND U2522 ( .A(n315), .B(n2644), .Z(n2643) );
  XNOR U2523 ( .A(p_input[1251]), .B(n2642), .Z(n2644) );
  XOR U2524 ( .A(n2645), .B(n2646), .Z(n2642) );
  AND U2525 ( .A(n319), .B(n2647), .Z(n2646) );
  XNOR U2526 ( .A(p_input[1267]), .B(n2645), .Z(n2647) );
  XOR U2527 ( .A(n2648), .B(n2649), .Z(n2645) );
  AND U2528 ( .A(n323), .B(n2650), .Z(n2649) );
  XNOR U2529 ( .A(p_input[1283]), .B(n2648), .Z(n2650) );
  XOR U2530 ( .A(n2651), .B(n2652), .Z(n2648) );
  AND U2531 ( .A(n327), .B(n2653), .Z(n2652) );
  XNOR U2532 ( .A(p_input[1299]), .B(n2651), .Z(n2653) );
  XOR U2533 ( .A(n2654), .B(n2655), .Z(n2651) );
  AND U2534 ( .A(n331), .B(n2656), .Z(n2655) );
  XNOR U2535 ( .A(p_input[1315]), .B(n2654), .Z(n2656) );
  XOR U2536 ( .A(n2657), .B(n2658), .Z(n2654) );
  AND U2537 ( .A(n335), .B(n2659), .Z(n2658) );
  XNOR U2538 ( .A(p_input[1331]), .B(n2657), .Z(n2659) );
  XOR U2539 ( .A(n2660), .B(n2661), .Z(n2657) );
  AND U2540 ( .A(n339), .B(n2662), .Z(n2661) );
  XNOR U2541 ( .A(p_input[1347]), .B(n2660), .Z(n2662) );
  XOR U2542 ( .A(n2663), .B(n2664), .Z(n2660) );
  AND U2543 ( .A(n343), .B(n2665), .Z(n2664) );
  XNOR U2544 ( .A(p_input[1363]), .B(n2663), .Z(n2665) );
  XOR U2545 ( .A(n2666), .B(n2667), .Z(n2663) );
  AND U2546 ( .A(n347), .B(n2668), .Z(n2667) );
  XNOR U2547 ( .A(p_input[1379]), .B(n2666), .Z(n2668) );
  XOR U2548 ( .A(n2669), .B(n2670), .Z(n2666) );
  AND U2549 ( .A(n351), .B(n2671), .Z(n2670) );
  XNOR U2550 ( .A(p_input[1395]), .B(n2669), .Z(n2671) );
  XOR U2551 ( .A(n2672), .B(n2673), .Z(n2669) );
  AND U2552 ( .A(n355), .B(n2674), .Z(n2673) );
  XNOR U2553 ( .A(p_input[1411]), .B(n2672), .Z(n2674) );
  XOR U2554 ( .A(n2675), .B(n2676), .Z(n2672) );
  AND U2555 ( .A(n359), .B(n2677), .Z(n2676) );
  XNOR U2556 ( .A(p_input[1427]), .B(n2675), .Z(n2677) );
  XOR U2557 ( .A(n2678), .B(n2679), .Z(n2675) );
  AND U2558 ( .A(n363), .B(n2680), .Z(n2679) );
  XNOR U2559 ( .A(p_input[1443]), .B(n2678), .Z(n2680) );
  XOR U2560 ( .A(n2681), .B(n2682), .Z(n2678) );
  AND U2561 ( .A(n367), .B(n2683), .Z(n2682) );
  XNOR U2562 ( .A(p_input[1459]), .B(n2681), .Z(n2683) );
  XOR U2563 ( .A(n2684), .B(n2685), .Z(n2681) );
  AND U2564 ( .A(n371), .B(n2686), .Z(n2685) );
  XNOR U2565 ( .A(p_input[1475]), .B(n2684), .Z(n2686) );
  XOR U2566 ( .A(n2687), .B(n2688), .Z(n2684) );
  AND U2567 ( .A(n375), .B(n2689), .Z(n2688) );
  XNOR U2568 ( .A(p_input[1491]), .B(n2687), .Z(n2689) );
  XOR U2569 ( .A(n2690), .B(n2691), .Z(n2687) );
  AND U2570 ( .A(n379), .B(n2692), .Z(n2691) );
  XNOR U2571 ( .A(p_input[1507]), .B(n2690), .Z(n2692) );
  XOR U2572 ( .A(n2693), .B(n2694), .Z(n2690) );
  AND U2573 ( .A(n383), .B(n2695), .Z(n2694) );
  XNOR U2574 ( .A(p_input[1523]), .B(n2693), .Z(n2695) );
  XOR U2575 ( .A(n2696), .B(n2697), .Z(n2693) );
  AND U2576 ( .A(n387), .B(n2698), .Z(n2697) );
  XNOR U2577 ( .A(p_input[1539]), .B(n2696), .Z(n2698) );
  XOR U2578 ( .A(n2699), .B(n2700), .Z(n2696) );
  AND U2579 ( .A(n391), .B(n2701), .Z(n2700) );
  XNOR U2580 ( .A(p_input[1555]), .B(n2699), .Z(n2701) );
  XOR U2581 ( .A(n2702), .B(n2703), .Z(n2699) );
  AND U2582 ( .A(n395), .B(n2704), .Z(n2703) );
  XNOR U2583 ( .A(p_input[1571]), .B(n2702), .Z(n2704) );
  XOR U2584 ( .A(n2705), .B(n2706), .Z(n2702) );
  AND U2585 ( .A(n399), .B(n2707), .Z(n2706) );
  XNOR U2586 ( .A(p_input[1587]), .B(n2705), .Z(n2707) );
  XOR U2587 ( .A(n2708), .B(n2709), .Z(n2705) );
  AND U2588 ( .A(n403), .B(n2710), .Z(n2709) );
  XNOR U2589 ( .A(p_input[1603]), .B(n2708), .Z(n2710) );
  XOR U2590 ( .A(n2711), .B(n2712), .Z(n2708) );
  AND U2591 ( .A(n407), .B(n2713), .Z(n2712) );
  XNOR U2592 ( .A(p_input[1619]), .B(n2711), .Z(n2713) );
  XOR U2593 ( .A(n2714), .B(n2715), .Z(n2711) );
  AND U2594 ( .A(n411), .B(n2716), .Z(n2715) );
  XNOR U2595 ( .A(p_input[1635]), .B(n2714), .Z(n2716) );
  XOR U2596 ( .A(n2717), .B(n2718), .Z(n2714) );
  AND U2597 ( .A(n415), .B(n2719), .Z(n2718) );
  XNOR U2598 ( .A(p_input[1651]), .B(n2717), .Z(n2719) );
  XOR U2599 ( .A(n2720), .B(n2721), .Z(n2717) );
  AND U2600 ( .A(n419), .B(n2722), .Z(n2721) );
  XNOR U2601 ( .A(p_input[1667]), .B(n2720), .Z(n2722) );
  XOR U2602 ( .A(n2723), .B(n2724), .Z(n2720) );
  AND U2603 ( .A(n423), .B(n2725), .Z(n2724) );
  XNOR U2604 ( .A(p_input[1683]), .B(n2723), .Z(n2725) );
  XOR U2605 ( .A(n2726), .B(n2727), .Z(n2723) );
  AND U2606 ( .A(n427), .B(n2728), .Z(n2727) );
  XNOR U2607 ( .A(p_input[1699]), .B(n2726), .Z(n2728) );
  XOR U2608 ( .A(n2729), .B(n2730), .Z(n2726) );
  AND U2609 ( .A(n431), .B(n2731), .Z(n2730) );
  XNOR U2610 ( .A(p_input[1715]), .B(n2729), .Z(n2731) );
  XOR U2611 ( .A(n2732), .B(n2733), .Z(n2729) );
  AND U2612 ( .A(n435), .B(n2734), .Z(n2733) );
  XNOR U2613 ( .A(p_input[1731]), .B(n2732), .Z(n2734) );
  XOR U2614 ( .A(n2735), .B(n2736), .Z(n2732) );
  AND U2615 ( .A(n439), .B(n2737), .Z(n2736) );
  XNOR U2616 ( .A(p_input[1747]), .B(n2735), .Z(n2737) );
  XOR U2617 ( .A(n2738), .B(n2739), .Z(n2735) );
  AND U2618 ( .A(n443), .B(n2740), .Z(n2739) );
  XNOR U2619 ( .A(p_input[1763]), .B(n2738), .Z(n2740) );
  XOR U2620 ( .A(n2741), .B(n2742), .Z(n2738) );
  AND U2621 ( .A(n447), .B(n2743), .Z(n2742) );
  XNOR U2622 ( .A(p_input[1779]), .B(n2741), .Z(n2743) );
  XOR U2623 ( .A(n2744), .B(n2745), .Z(n2741) );
  AND U2624 ( .A(n451), .B(n2746), .Z(n2745) );
  XNOR U2625 ( .A(p_input[1795]), .B(n2744), .Z(n2746) );
  XOR U2626 ( .A(n2747), .B(n2748), .Z(n2744) );
  AND U2627 ( .A(n455), .B(n2749), .Z(n2748) );
  XNOR U2628 ( .A(p_input[1811]), .B(n2747), .Z(n2749) );
  XOR U2629 ( .A(n2750), .B(n2751), .Z(n2747) );
  AND U2630 ( .A(n459), .B(n2752), .Z(n2751) );
  XNOR U2631 ( .A(p_input[1827]), .B(n2750), .Z(n2752) );
  XOR U2632 ( .A(n2753), .B(n2754), .Z(n2750) );
  AND U2633 ( .A(n463), .B(n2755), .Z(n2754) );
  XNOR U2634 ( .A(p_input[1843]), .B(n2753), .Z(n2755) );
  XOR U2635 ( .A(n2756), .B(n2757), .Z(n2753) );
  AND U2636 ( .A(n467), .B(n2758), .Z(n2757) );
  XNOR U2637 ( .A(p_input[1859]), .B(n2756), .Z(n2758) );
  XOR U2638 ( .A(n2759), .B(n2760), .Z(n2756) );
  AND U2639 ( .A(n471), .B(n2761), .Z(n2760) );
  XNOR U2640 ( .A(p_input[1875]), .B(n2759), .Z(n2761) );
  XOR U2641 ( .A(n2762), .B(n2763), .Z(n2759) );
  AND U2642 ( .A(n475), .B(n2764), .Z(n2763) );
  XNOR U2643 ( .A(p_input[1891]), .B(n2762), .Z(n2764) );
  XOR U2644 ( .A(n2765), .B(n2766), .Z(n2762) );
  AND U2645 ( .A(n479), .B(n2767), .Z(n2766) );
  XNOR U2646 ( .A(p_input[1907]), .B(n2765), .Z(n2767) );
  XOR U2647 ( .A(n2768), .B(n2769), .Z(n2765) );
  AND U2648 ( .A(n483), .B(n2770), .Z(n2769) );
  XNOR U2649 ( .A(p_input[1923]), .B(n2768), .Z(n2770) );
  XOR U2650 ( .A(n2771), .B(n2772), .Z(n2768) );
  AND U2651 ( .A(n487), .B(n2773), .Z(n2772) );
  XNOR U2652 ( .A(p_input[1939]), .B(n2771), .Z(n2773) );
  XOR U2653 ( .A(n2774), .B(n2775), .Z(n2771) );
  AND U2654 ( .A(n491), .B(n2776), .Z(n2775) );
  XNOR U2655 ( .A(p_input[1955]), .B(n2774), .Z(n2776) );
  XOR U2656 ( .A(n2777), .B(n2778), .Z(n2774) );
  AND U2657 ( .A(n495), .B(n2779), .Z(n2778) );
  XNOR U2658 ( .A(p_input[1971]), .B(n2777), .Z(n2779) );
  XOR U2659 ( .A(n2780), .B(n2781), .Z(n2777) );
  AND U2660 ( .A(n499), .B(n2782), .Z(n2781) );
  XNOR U2661 ( .A(p_input[1987]), .B(n2780), .Z(n2782) );
  XNOR U2662 ( .A(n2783), .B(n2784), .Z(n2780) );
  AND U2663 ( .A(n503), .B(n2785), .Z(n2784) );
  XOR U2664 ( .A(p_input[2003]), .B(n2783), .Z(n2785) );
  XOR U2665 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n2786), .Z(n2783) );
  AND U2666 ( .A(n506), .B(n2787), .Z(n2786) );
  XOR U2667 ( .A(p_input[2019]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n2787)
         );
  XNOR U2668 ( .A(n2788), .B(n2789), .Z(o[2]) );
  AND U2669 ( .A(n3), .B(n2790), .Z(n2788) );
  XNOR U2670 ( .A(p_input[2]), .B(n2789), .Z(n2790) );
  XOR U2671 ( .A(n2791), .B(n2792), .Z(n2789) );
  AND U2672 ( .A(n7), .B(n2793), .Z(n2792) );
  XNOR U2673 ( .A(p_input[18]), .B(n2791), .Z(n2793) );
  XOR U2674 ( .A(n2794), .B(n2795), .Z(n2791) );
  AND U2675 ( .A(n11), .B(n2796), .Z(n2795) );
  XNOR U2676 ( .A(p_input[34]), .B(n2794), .Z(n2796) );
  XOR U2677 ( .A(n2797), .B(n2798), .Z(n2794) );
  AND U2678 ( .A(n15), .B(n2799), .Z(n2798) );
  XNOR U2679 ( .A(p_input[50]), .B(n2797), .Z(n2799) );
  XOR U2680 ( .A(n2800), .B(n2801), .Z(n2797) );
  AND U2681 ( .A(n19), .B(n2802), .Z(n2801) );
  XNOR U2682 ( .A(p_input[66]), .B(n2800), .Z(n2802) );
  XOR U2683 ( .A(n2803), .B(n2804), .Z(n2800) );
  AND U2684 ( .A(n23), .B(n2805), .Z(n2804) );
  XNOR U2685 ( .A(p_input[82]), .B(n2803), .Z(n2805) );
  XOR U2686 ( .A(n2806), .B(n2807), .Z(n2803) );
  AND U2687 ( .A(n27), .B(n2808), .Z(n2807) );
  XNOR U2688 ( .A(p_input[98]), .B(n2806), .Z(n2808) );
  XOR U2689 ( .A(n2809), .B(n2810), .Z(n2806) );
  AND U2690 ( .A(n31), .B(n2811), .Z(n2810) );
  XNOR U2691 ( .A(p_input[114]), .B(n2809), .Z(n2811) );
  XOR U2692 ( .A(n2812), .B(n2813), .Z(n2809) );
  AND U2693 ( .A(n35), .B(n2814), .Z(n2813) );
  XNOR U2694 ( .A(p_input[130]), .B(n2812), .Z(n2814) );
  XOR U2695 ( .A(n2815), .B(n2816), .Z(n2812) );
  AND U2696 ( .A(n39), .B(n2817), .Z(n2816) );
  XNOR U2697 ( .A(p_input[146]), .B(n2815), .Z(n2817) );
  XOR U2698 ( .A(n2818), .B(n2819), .Z(n2815) );
  AND U2699 ( .A(n43), .B(n2820), .Z(n2819) );
  XNOR U2700 ( .A(p_input[162]), .B(n2818), .Z(n2820) );
  XOR U2701 ( .A(n2821), .B(n2822), .Z(n2818) );
  AND U2702 ( .A(n47), .B(n2823), .Z(n2822) );
  XNOR U2703 ( .A(p_input[178]), .B(n2821), .Z(n2823) );
  XOR U2704 ( .A(n2824), .B(n2825), .Z(n2821) );
  AND U2705 ( .A(n51), .B(n2826), .Z(n2825) );
  XNOR U2706 ( .A(p_input[194]), .B(n2824), .Z(n2826) );
  XOR U2707 ( .A(n2827), .B(n2828), .Z(n2824) );
  AND U2708 ( .A(n55), .B(n2829), .Z(n2828) );
  XNOR U2709 ( .A(p_input[210]), .B(n2827), .Z(n2829) );
  XOR U2710 ( .A(n2830), .B(n2831), .Z(n2827) );
  AND U2711 ( .A(n59), .B(n2832), .Z(n2831) );
  XNOR U2712 ( .A(p_input[226]), .B(n2830), .Z(n2832) );
  XOR U2713 ( .A(n2833), .B(n2834), .Z(n2830) );
  AND U2714 ( .A(n63), .B(n2835), .Z(n2834) );
  XNOR U2715 ( .A(p_input[242]), .B(n2833), .Z(n2835) );
  XOR U2716 ( .A(n2836), .B(n2837), .Z(n2833) );
  AND U2717 ( .A(n67), .B(n2838), .Z(n2837) );
  XNOR U2718 ( .A(p_input[258]), .B(n2836), .Z(n2838) );
  XOR U2719 ( .A(n2839), .B(n2840), .Z(n2836) );
  AND U2720 ( .A(n71), .B(n2841), .Z(n2840) );
  XNOR U2721 ( .A(p_input[274]), .B(n2839), .Z(n2841) );
  XOR U2722 ( .A(n2842), .B(n2843), .Z(n2839) );
  AND U2723 ( .A(n75), .B(n2844), .Z(n2843) );
  XNOR U2724 ( .A(p_input[290]), .B(n2842), .Z(n2844) );
  XOR U2725 ( .A(n2845), .B(n2846), .Z(n2842) );
  AND U2726 ( .A(n79), .B(n2847), .Z(n2846) );
  XNOR U2727 ( .A(p_input[306]), .B(n2845), .Z(n2847) );
  XOR U2728 ( .A(n2848), .B(n2849), .Z(n2845) );
  AND U2729 ( .A(n83), .B(n2850), .Z(n2849) );
  XNOR U2730 ( .A(p_input[322]), .B(n2848), .Z(n2850) );
  XOR U2731 ( .A(n2851), .B(n2852), .Z(n2848) );
  AND U2732 ( .A(n87), .B(n2853), .Z(n2852) );
  XNOR U2733 ( .A(p_input[338]), .B(n2851), .Z(n2853) );
  XOR U2734 ( .A(n2854), .B(n2855), .Z(n2851) );
  AND U2735 ( .A(n91), .B(n2856), .Z(n2855) );
  XNOR U2736 ( .A(p_input[354]), .B(n2854), .Z(n2856) );
  XOR U2737 ( .A(n2857), .B(n2858), .Z(n2854) );
  AND U2738 ( .A(n95), .B(n2859), .Z(n2858) );
  XNOR U2739 ( .A(p_input[370]), .B(n2857), .Z(n2859) );
  XOR U2740 ( .A(n2860), .B(n2861), .Z(n2857) );
  AND U2741 ( .A(n99), .B(n2862), .Z(n2861) );
  XNOR U2742 ( .A(p_input[386]), .B(n2860), .Z(n2862) );
  XOR U2743 ( .A(n2863), .B(n2864), .Z(n2860) );
  AND U2744 ( .A(n103), .B(n2865), .Z(n2864) );
  XNOR U2745 ( .A(p_input[402]), .B(n2863), .Z(n2865) );
  XOR U2746 ( .A(n2866), .B(n2867), .Z(n2863) );
  AND U2747 ( .A(n107), .B(n2868), .Z(n2867) );
  XNOR U2748 ( .A(p_input[418]), .B(n2866), .Z(n2868) );
  XOR U2749 ( .A(n2869), .B(n2870), .Z(n2866) );
  AND U2750 ( .A(n111), .B(n2871), .Z(n2870) );
  XNOR U2751 ( .A(p_input[434]), .B(n2869), .Z(n2871) );
  XOR U2752 ( .A(n2872), .B(n2873), .Z(n2869) );
  AND U2753 ( .A(n115), .B(n2874), .Z(n2873) );
  XNOR U2754 ( .A(p_input[450]), .B(n2872), .Z(n2874) );
  XOR U2755 ( .A(n2875), .B(n2876), .Z(n2872) );
  AND U2756 ( .A(n119), .B(n2877), .Z(n2876) );
  XNOR U2757 ( .A(p_input[466]), .B(n2875), .Z(n2877) );
  XOR U2758 ( .A(n2878), .B(n2879), .Z(n2875) );
  AND U2759 ( .A(n123), .B(n2880), .Z(n2879) );
  XNOR U2760 ( .A(p_input[482]), .B(n2878), .Z(n2880) );
  XOR U2761 ( .A(n2881), .B(n2882), .Z(n2878) );
  AND U2762 ( .A(n127), .B(n2883), .Z(n2882) );
  XNOR U2763 ( .A(p_input[498]), .B(n2881), .Z(n2883) );
  XOR U2764 ( .A(n2884), .B(n2885), .Z(n2881) );
  AND U2765 ( .A(n131), .B(n2886), .Z(n2885) );
  XNOR U2766 ( .A(p_input[514]), .B(n2884), .Z(n2886) );
  XOR U2767 ( .A(n2887), .B(n2888), .Z(n2884) );
  AND U2768 ( .A(n135), .B(n2889), .Z(n2888) );
  XNOR U2769 ( .A(p_input[530]), .B(n2887), .Z(n2889) );
  XOR U2770 ( .A(n2890), .B(n2891), .Z(n2887) );
  AND U2771 ( .A(n139), .B(n2892), .Z(n2891) );
  XNOR U2772 ( .A(p_input[546]), .B(n2890), .Z(n2892) );
  XOR U2773 ( .A(n2893), .B(n2894), .Z(n2890) );
  AND U2774 ( .A(n143), .B(n2895), .Z(n2894) );
  XNOR U2775 ( .A(p_input[562]), .B(n2893), .Z(n2895) );
  XOR U2776 ( .A(n2896), .B(n2897), .Z(n2893) );
  AND U2777 ( .A(n147), .B(n2898), .Z(n2897) );
  XNOR U2778 ( .A(p_input[578]), .B(n2896), .Z(n2898) );
  XOR U2779 ( .A(n2899), .B(n2900), .Z(n2896) );
  AND U2780 ( .A(n151), .B(n2901), .Z(n2900) );
  XNOR U2781 ( .A(p_input[594]), .B(n2899), .Z(n2901) );
  XOR U2782 ( .A(n2902), .B(n2903), .Z(n2899) );
  AND U2783 ( .A(n155), .B(n2904), .Z(n2903) );
  XNOR U2784 ( .A(p_input[610]), .B(n2902), .Z(n2904) );
  XOR U2785 ( .A(n2905), .B(n2906), .Z(n2902) );
  AND U2786 ( .A(n159), .B(n2907), .Z(n2906) );
  XNOR U2787 ( .A(p_input[626]), .B(n2905), .Z(n2907) );
  XOR U2788 ( .A(n2908), .B(n2909), .Z(n2905) );
  AND U2789 ( .A(n163), .B(n2910), .Z(n2909) );
  XNOR U2790 ( .A(p_input[642]), .B(n2908), .Z(n2910) );
  XOR U2791 ( .A(n2911), .B(n2912), .Z(n2908) );
  AND U2792 ( .A(n167), .B(n2913), .Z(n2912) );
  XNOR U2793 ( .A(p_input[658]), .B(n2911), .Z(n2913) );
  XOR U2794 ( .A(n2914), .B(n2915), .Z(n2911) );
  AND U2795 ( .A(n171), .B(n2916), .Z(n2915) );
  XNOR U2796 ( .A(p_input[674]), .B(n2914), .Z(n2916) );
  XOR U2797 ( .A(n2917), .B(n2918), .Z(n2914) );
  AND U2798 ( .A(n175), .B(n2919), .Z(n2918) );
  XNOR U2799 ( .A(p_input[690]), .B(n2917), .Z(n2919) );
  XOR U2800 ( .A(n2920), .B(n2921), .Z(n2917) );
  AND U2801 ( .A(n179), .B(n2922), .Z(n2921) );
  XNOR U2802 ( .A(p_input[706]), .B(n2920), .Z(n2922) );
  XOR U2803 ( .A(n2923), .B(n2924), .Z(n2920) );
  AND U2804 ( .A(n183), .B(n2925), .Z(n2924) );
  XNOR U2805 ( .A(p_input[722]), .B(n2923), .Z(n2925) );
  XOR U2806 ( .A(n2926), .B(n2927), .Z(n2923) );
  AND U2807 ( .A(n187), .B(n2928), .Z(n2927) );
  XNOR U2808 ( .A(p_input[738]), .B(n2926), .Z(n2928) );
  XOR U2809 ( .A(n2929), .B(n2930), .Z(n2926) );
  AND U2810 ( .A(n191), .B(n2931), .Z(n2930) );
  XNOR U2811 ( .A(p_input[754]), .B(n2929), .Z(n2931) );
  XOR U2812 ( .A(n2932), .B(n2933), .Z(n2929) );
  AND U2813 ( .A(n195), .B(n2934), .Z(n2933) );
  XNOR U2814 ( .A(p_input[770]), .B(n2932), .Z(n2934) );
  XOR U2815 ( .A(n2935), .B(n2936), .Z(n2932) );
  AND U2816 ( .A(n199), .B(n2937), .Z(n2936) );
  XNOR U2817 ( .A(p_input[786]), .B(n2935), .Z(n2937) );
  XOR U2818 ( .A(n2938), .B(n2939), .Z(n2935) );
  AND U2819 ( .A(n203), .B(n2940), .Z(n2939) );
  XNOR U2820 ( .A(p_input[802]), .B(n2938), .Z(n2940) );
  XOR U2821 ( .A(n2941), .B(n2942), .Z(n2938) );
  AND U2822 ( .A(n207), .B(n2943), .Z(n2942) );
  XNOR U2823 ( .A(p_input[818]), .B(n2941), .Z(n2943) );
  XOR U2824 ( .A(n2944), .B(n2945), .Z(n2941) );
  AND U2825 ( .A(n211), .B(n2946), .Z(n2945) );
  XNOR U2826 ( .A(p_input[834]), .B(n2944), .Z(n2946) );
  XOR U2827 ( .A(n2947), .B(n2948), .Z(n2944) );
  AND U2828 ( .A(n215), .B(n2949), .Z(n2948) );
  XNOR U2829 ( .A(p_input[850]), .B(n2947), .Z(n2949) );
  XOR U2830 ( .A(n2950), .B(n2951), .Z(n2947) );
  AND U2831 ( .A(n219), .B(n2952), .Z(n2951) );
  XNOR U2832 ( .A(p_input[866]), .B(n2950), .Z(n2952) );
  XOR U2833 ( .A(n2953), .B(n2954), .Z(n2950) );
  AND U2834 ( .A(n223), .B(n2955), .Z(n2954) );
  XNOR U2835 ( .A(p_input[882]), .B(n2953), .Z(n2955) );
  XOR U2836 ( .A(n2956), .B(n2957), .Z(n2953) );
  AND U2837 ( .A(n227), .B(n2958), .Z(n2957) );
  XNOR U2838 ( .A(p_input[898]), .B(n2956), .Z(n2958) );
  XOR U2839 ( .A(n2959), .B(n2960), .Z(n2956) );
  AND U2840 ( .A(n231), .B(n2961), .Z(n2960) );
  XNOR U2841 ( .A(p_input[914]), .B(n2959), .Z(n2961) );
  XOR U2842 ( .A(n2962), .B(n2963), .Z(n2959) );
  AND U2843 ( .A(n235), .B(n2964), .Z(n2963) );
  XNOR U2844 ( .A(p_input[930]), .B(n2962), .Z(n2964) );
  XOR U2845 ( .A(n2965), .B(n2966), .Z(n2962) );
  AND U2846 ( .A(n239), .B(n2967), .Z(n2966) );
  XNOR U2847 ( .A(p_input[946]), .B(n2965), .Z(n2967) );
  XOR U2848 ( .A(n2968), .B(n2969), .Z(n2965) );
  AND U2849 ( .A(n243), .B(n2970), .Z(n2969) );
  XNOR U2850 ( .A(p_input[962]), .B(n2968), .Z(n2970) );
  XOR U2851 ( .A(n2971), .B(n2972), .Z(n2968) );
  AND U2852 ( .A(n247), .B(n2973), .Z(n2972) );
  XNOR U2853 ( .A(p_input[978]), .B(n2971), .Z(n2973) );
  XOR U2854 ( .A(n2974), .B(n2975), .Z(n2971) );
  AND U2855 ( .A(n251), .B(n2976), .Z(n2975) );
  XNOR U2856 ( .A(p_input[994]), .B(n2974), .Z(n2976) );
  XOR U2857 ( .A(n2977), .B(n2978), .Z(n2974) );
  AND U2858 ( .A(n255), .B(n2979), .Z(n2978) );
  XNOR U2859 ( .A(p_input[1010]), .B(n2977), .Z(n2979) );
  XOR U2860 ( .A(n2980), .B(n2981), .Z(n2977) );
  AND U2861 ( .A(n259), .B(n2982), .Z(n2981) );
  XNOR U2862 ( .A(p_input[1026]), .B(n2980), .Z(n2982) );
  XOR U2863 ( .A(n2983), .B(n2984), .Z(n2980) );
  AND U2864 ( .A(n263), .B(n2985), .Z(n2984) );
  XNOR U2865 ( .A(p_input[1042]), .B(n2983), .Z(n2985) );
  XOR U2866 ( .A(n2986), .B(n2987), .Z(n2983) );
  AND U2867 ( .A(n267), .B(n2988), .Z(n2987) );
  XNOR U2868 ( .A(p_input[1058]), .B(n2986), .Z(n2988) );
  XOR U2869 ( .A(n2989), .B(n2990), .Z(n2986) );
  AND U2870 ( .A(n271), .B(n2991), .Z(n2990) );
  XNOR U2871 ( .A(p_input[1074]), .B(n2989), .Z(n2991) );
  XOR U2872 ( .A(n2992), .B(n2993), .Z(n2989) );
  AND U2873 ( .A(n275), .B(n2994), .Z(n2993) );
  XNOR U2874 ( .A(p_input[1090]), .B(n2992), .Z(n2994) );
  XOR U2875 ( .A(n2995), .B(n2996), .Z(n2992) );
  AND U2876 ( .A(n279), .B(n2997), .Z(n2996) );
  XNOR U2877 ( .A(p_input[1106]), .B(n2995), .Z(n2997) );
  XOR U2878 ( .A(n2998), .B(n2999), .Z(n2995) );
  AND U2879 ( .A(n283), .B(n3000), .Z(n2999) );
  XNOR U2880 ( .A(p_input[1122]), .B(n2998), .Z(n3000) );
  XOR U2881 ( .A(n3001), .B(n3002), .Z(n2998) );
  AND U2882 ( .A(n287), .B(n3003), .Z(n3002) );
  XNOR U2883 ( .A(p_input[1138]), .B(n3001), .Z(n3003) );
  XOR U2884 ( .A(n3004), .B(n3005), .Z(n3001) );
  AND U2885 ( .A(n291), .B(n3006), .Z(n3005) );
  XNOR U2886 ( .A(p_input[1154]), .B(n3004), .Z(n3006) );
  XOR U2887 ( .A(n3007), .B(n3008), .Z(n3004) );
  AND U2888 ( .A(n295), .B(n3009), .Z(n3008) );
  XNOR U2889 ( .A(p_input[1170]), .B(n3007), .Z(n3009) );
  XOR U2890 ( .A(n3010), .B(n3011), .Z(n3007) );
  AND U2891 ( .A(n299), .B(n3012), .Z(n3011) );
  XNOR U2892 ( .A(p_input[1186]), .B(n3010), .Z(n3012) );
  XOR U2893 ( .A(n3013), .B(n3014), .Z(n3010) );
  AND U2894 ( .A(n303), .B(n3015), .Z(n3014) );
  XNOR U2895 ( .A(p_input[1202]), .B(n3013), .Z(n3015) );
  XOR U2896 ( .A(n3016), .B(n3017), .Z(n3013) );
  AND U2897 ( .A(n307), .B(n3018), .Z(n3017) );
  XNOR U2898 ( .A(p_input[1218]), .B(n3016), .Z(n3018) );
  XOR U2899 ( .A(n3019), .B(n3020), .Z(n3016) );
  AND U2900 ( .A(n311), .B(n3021), .Z(n3020) );
  XNOR U2901 ( .A(p_input[1234]), .B(n3019), .Z(n3021) );
  XOR U2902 ( .A(n3022), .B(n3023), .Z(n3019) );
  AND U2903 ( .A(n315), .B(n3024), .Z(n3023) );
  XNOR U2904 ( .A(p_input[1250]), .B(n3022), .Z(n3024) );
  XOR U2905 ( .A(n3025), .B(n3026), .Z(n3022) );
  AND U2906 ( .A(n319), .B(n3027), .Z(n3026) );
  XNOR U2907 ( .A(p_input[1266]), .B(n3025), .Z(n3027) );
  XOR U2908 ( .A(n3028), .B(n3029), .Z(n3025) );
  AND U2909 ( .A(n323), .B(n3030), .Z(n3029) );
  XNOR U2910 ( .A(p_input[1282]), .B(n3028), .Z(n3030) );
  XOR U2911 ( .A(n3031), .B(n3032), .Z(n3028) );
  AND U2912 ( .A(n327), .B(n3033), .Z(n3032) );
  XNOR U2913 ( .A(p_input[1298]), .B(n3031), .Z(n3033) );
  XOR U2914 ( .A(n3034), .B(n3035), .Z(n3031) );
  AND U2915 ( .A(n331), .B(n3036), .Z(n3035) );
  XNOR U2916 ( .A(p_input[1314]), .B(n3034), .Z(n3036) );
  XOR U2917 ( .A(n3037), .B(n3038), .Z(n3034) );
  AND U2918 ( .A(n335), .B(n3039), .Z(n3038) );
  XNOR U2919 ( .A(p_input[1330]), .B(n3037), .Z(n3039) );
  XOR U2920 ( .A(n3040), .B(n3041), .Z(n3037) );
  AND U2921 ( .A(n339), .B(n3042), .Z(n3041) );
  XNOR U2922 ( .A(p_input[1346]), .B(n3040), .Z(n3042) );
  XOR U2923 ( .A(n3043), .B(n3044), .Z(n3040) );
  AND U2924 ( .A(n343), .B(n3045), .Z(n3044) );
  XNOR U2925 ( .A(p_input[1362]), .B(n3043), .Z(n3045) );
  XOR U2926 ( .A(n3046), .B(n3047), .Z(n3043) );
  AND U2927 ( .A(n347), .B(n3048), .Z(n3047) );
  XNOR U2928 ( .A(p_input[1378]), .B(n3046), .Z(n3048) );
  XOR U2929 ( .A(n3049), .B(n3050), .Z(n3046) );
  AND U2930 ( .A(n351), .B(n3051), .Z(n3050) );
  XNOR U2931 ( .A(p_input[1394]), .B(n3049), .Z(n3051) );
  XOR U2932 ( .A(n3052), .B(n3053), .Z(n3049) );
  AND U2933 ( .A(n355), .B(n3054), .Z(n3053) );
  XNOR U2934 ( .A(p_input[1410]), .B(n3052), .Z(n3054) );
  XOR U2935 ( .A(n3055), .B(n3056), .Z(n3052) );
  AND U2936 ( .A(n359), .B(n3057), .Z(n3056) );
  XNOR U2937 ( .A(p_input[1426]), .B(n3055), .Z(n3057) );
  XOR U2938 ( .A(n3058), .B(n3059), .Z(n3055) );
  AND U2939 ( .A(n363), .B(n3060), .Z(n3059) );
  XNOR U2940 ( .A(p_input[1442]), .B(n3058), .Z(n3060) );
  XOR U2941 ( .A(n3061), .B(n3062), .Z(n3058) );
  AND U2942 ( .A(n367), .B(n3063), .Z(n3062) );
  XNOR U2943 ( .A(p_input[1458]), .B(n3061), .Z(n3063) );
  XOR U2944 ( .A(n3064), .B(n3065), .Z(n3061) );
  AND U2945 ( .A(n371), .B(n3066), .Z(n3065) );
  XNOR U2946 ( .A(p_input[1474]), .B(n3064), .Z(n3066) );
  XOR U2947 ( .A(n3067), .B(n3068), .Z(n3064) );
  AND U2948 ( .A(n375), .B(n3069), .Z(n3068) );
  XNOR U2949 ( .A(p_input[1490]), .B(n3067), .Z(n3069) );
  XOR U2950 ( .A(n3070), .B(n3071), .Z(n3067) );
  AND U2951 ( .A(n379), .B(n3072), .Z(n3071) );
  XNOR U2952 ( .A(p_input[1506]), .B(n3070), .Z(n3072) );
  XOR U2953 ( .A(n3073), .B(n3074), .Z(n3070) );
  AND U2954 ( .A(n383), .B(n3075), .Z(n3074) );
  XNOR U2955 ( .A(p_input[1522]), .B(n3073), .Z(n3075) );
  XOR U2956 ( .A(n3076), .B(n3077), .Z(n3073) );
  AND U2957 ( .A(n387), .B(n3078), .Z(n3077) );
  XNOR U2958 ( .A(p_input[1538]), .B(n3076), .Z(n3078) );
  XOR U2959 ( .A(n3079), .B(n3080), .Z(n3076) );
  AND U2960 ( .A(n391), .B(n3081), .Z(n3080) );
  XNOR U2961 ( .A(p_input[1554]), .B(n3079), .Z(n3081) );
  XOR U2962 ( .A(n3082), .B(n3083), .Z(n3079) );
  AND U2963 ( .A(n395), .B(n3084), .Z(n3083) );
  XNOR U2964 ( .A(p_input[1570]), .B(n3082), .Z(n3084) );
  XOR U2965 ( .A(n3085), .B(n3086), .Z(n3082) );
  AND U2966 ( .A(n399), .B(n3087), .Z(n3086) );
  XNOR U2967 ( .A(p_input[1586]), .B(n3085), .Z(n3087) );
  XOR U2968 ( .A(n3088), .B(n3089), .Z(n3085) );
  AND U2969 ( .A(n403), .B(n3090), .Z(n3089) );
  XNOR U2970 ( .A(p_input[1602]), .B(n3088), .Z(n3090) );
  XOR U2971 ( .A(n3091), .B(n3092), .Z(n3088) );
  AND U2972 ( .A(n407), .B(n3093), .Z(n3092) );
  XNOR U2973 ( .A(p_input[1618]), .B(n3091), .Z(n3093) );
  XOR U2974 ( .A(n3094), .B(n3095), .Z(n3091) );
  AND U2975 ( .A(n411), .B(n3096), .Z(n3095) );
  XNOR U2976 ( .A(p_input[1634]), .B(n3094), .Z(n3096) );
  XOR U2977 ( .A(n3097), .B(n3098), .Z(n3094) );
  AND U2978 ( .A(n415), .B(n3099), .Z(n3098) );
  XNOR U2979 ( .A(p_input[1650]), .B(n3097), .Z(n3099) );
  XOR U2980 ( .A(n3100), .B(n3101), .Z(n3097) );
  AND U2981 ( .A(n419), .B(n3102), .Z(n3101) );
  XNOR U2982 ( .A(p_input[1666]), .B(n3100), .Z(n3102) );
  XOR U2983 ( .A(n3103), .B(n3104), .Z(n3100) );
  AND U2984 ( .A(n423), .B(n3105), .Z(n3104) );
  XNOR U2985 ( .A(p_input[1682]), .B(n3103), .Z(n3105) );
  XOR U2986 ( .A(n3106), .B(n3107), .Z(n3103) );
  AND U2987 ( .A(n427), .B(n3108), .Z(n3107) );
  XNOR U2988 ( .A(p_input[1698]), .B(n3106), .Z(n3108) );
  XOR U2989 ( .A(n3109), .B(n3110), .Z(n3106) );
  AND U2990 ( .A(n431), .B(n3111), .Z(n3110) );
  XNOR U2991 ( .A(p_input[1714]), .B(n3109), .Z(n3111) );
  XOR U2992 ( .A(n3112), .B(n3113), .Z(n3109) );
  AND U2993 ( .A(n435), .B(n3114), .Z(n3113) );
  XNOR U2994 ( .A(p_input[1730]), .B(n3112), .Z(n3114) );
  XOR U2995 ( .A(n3115), .B(n3116), .Z(n3112) );
  AND U2996 ( .A(n439), .B(n3117), .Z(n3116) );
  XNOR U2997 ( .A(p_input[1746]), .B(n3115), .Z(n3117) );
  XOR U2998 ( .A(n3118), .B(n3119), .Z(n3115) );
  AND U2999 ( .A(n443), .B(n3120), .Z(n3119) );
  XNOR U3000 ( .A(p_input[1762]), .B(n3118), .Z(n3120) );
  XOR U3001 ( .A(n3121), .B(n3122), .Z(n3118) );
  AND U3002 ( .A(n447), .B(n3123), .Z(n3122) );
  XNOR U3003 ( .A(p_input[1778]), .B(n3121), .Z(n3123) );
  XOR U3004 ( .A(n3124), .B(n3125), .Z(n3121) );
  AND U3005 ( .A(n451), .B(n3126), .Z(n3125) );
  XNOR U3006 ( .A(p_input[1794]), .B(n3124), .Z(n3126) );
  XOR U3007 ( .A(n3127), .B(n3128), .Z(n3124) );
  AND U3008 ( .A(n455), .B(n3129), .Z(n3128) );
  XNOR U3009 ( .A(p_input[1810]), .B(n3127), .Z(n3129) );
  XOR U3010 ( .A(n3130), .B(n3131), .Z(n3127) );
  AND U3011 ( .A(n459), .B(n3132), .Z(n3131) );
  XNOR U3012 ( .A(p_input[1826]), .B(n3130), .Z(n3132) );
  XOR U3013 ( .A(n3133), .B(n3134), .Z(n3130) );
  AND U3014 ( .A(n463), .B(n3135), .Z(n3134) );
  XNOR U3015 ( .A(p_input[1842]), .B(n3133), .Z(n3135) );
  XOR U3016 ( .A(n3136), .B(n3137), .Z(n3133) );
  AND U3017 ( .A(n467), .B(n3138), .Z(n3137) );
  XNOR U3018 ( .A(p_input[1858]), .B(n3136), .Z(n3138) );
  XOR U3019 ( .A(n3139), .B(n3140), .Z(n3136) );
  AND U3020 ( .A(n471), .B(n3141), .Z(n3140) );
  XNOR U3021 ( .A(p_input[1874]), .B(n3139), .Z(n3141) );
  XOR U3022 ( .A(n3142), .B(n3143), .Z(n3139) );
  AND U3023 ( .A(n475), .B(n3144), .Z(n3143) );
  XNOR U3024 ( .A(p_input[1890]), .B(n3142), .Z(n3144) );
  XOR U3025 ( .A(n3145), .B(n3146), .Z(n3142) );
  AND U3026 ( .A(n479), .B(n3147), .Z(n3146) );
  XNOR U3027 ( .A(p_input[1906]), .B(n3145), .Z(n3147) );
  XOR U3028 ( .A(n3148), .B(n3149), .Z(n3145) );
  AND U3029 ( .A(n483), .B(n3150), .Z(n3149) );
  XNOR U3030 ( .A(p_input[1922]), .B(n3148), .Z(n3150) );
  XOR U3031 ( .A(n3151), .B(n3152), .Z(n3148) );
  AND U3032 ( .A(n487), .B(n3153), .Z(n3152) );
  XNOR U3033 ( .A(p_input[1938]), .B(n3151), .Z(n3153) );
  XOR U3034 ( .A(n3154), .B(n3155), .Z(n3151) );
  AND U3035 ( .A(n491), .B(n3156), .Z(n3155) );
  XNOR U3036 ( .A(p_input[1954]), .B(n3154), .Z(n3156) );
  XOR U3037 ( .A(n3157), .B(n3158), .Z(n3154) );
  AND U3038 ( .A(n495), .B(n3159), .Z(n3158) );
  XNOR U3039 ( .A(p_input[1970]), .B(n3157), .Z(n3159) );
  XOR U3040 ( .A(n3160), .B(n3161), .Z(n3157) );
  AND U3041 ( .A(n499), .B(n3162), .Z(n3161) );
  XNOR U3042 ( .A(p_input[1986]), .B(n3160), .Z(n3162) );
  XNOR U3043 ( .A(n3163), .B(n3164), .Z(n3160) );
  AND U3044 ( .A(n503), .B(n3165), .Z(n3164) );
  XOR U3045 ( .A(p_input[2002]), .B(n3163), .Z(n3165) );
  XOR U3046 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n3166), .Z(n3163) );
  AND U3047 ( .A(n506), .B(n3167), .Z(n3166) );
  XOR U3048 ( .A(p_input[2018]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n3167)
         );
  XNOR U3049 ( .A(n3168), .B(n3169), .Z(o[1]) );
  AND U3050 ( .A(n3), .B(n3170), .Z(n3168) );
  XNOR U3051 ( .A(p_input[1]), .B(n3169), .Z(n3170) );
  XOR U3052 ( .A(n3171), .B(n3172), .Z(n3169) );
  AND U3053 ( .A(n7), .B(n3173), .Z(n3172) );
  XNOR U3054 ( .A(p_input[17]), .B(n3171), .Z(n3173) );
  XOR U3055 ( .A(n3174), .B(n3175), .Z(n3171) );
  AND U3056 ( .A(n11), .B(n3176), .Z(n3175) );
  XNOR U3057 ( .A(p_input[33]), .B(n3174), .Z(n3176) );
  XOR U3058 ( .A(n3177), .B(n3178), .Z(n3174) );
  AND U3059 ( .A(n15), .B(n3179), .Z(n3178) );
  XNOR U3060 ( .A(p_input[49]), .B(n3177), .Z(n3179) );
  XOR U3061 ( .A(n3180), .B(n3181), .Z(n3177) );
  AND U3062 ( .A(n19), .B(n3182), .Z(n3181) );
  XNOR U3063 ( .A(p_input[65]), .B(n3180), .Z(n3182) );
  XOR U3064 ( .A(n3183), .B(n3184), .Z(n3180) );
  AND U3065 ( .A(n23), .B(n3185), .Z(n3184) );
  XNOR U3066 ( .A(p_input[81]), .B(n3183), .Z(n3185) );
  XOR U3067 ( .A(n3186), .B(n3187), .Z(n3183) );
  AND U3068 ( .A(n27), .B(n3188), .Z(n3187) );
  XNOR U3069 ( .A(p_input[97]), .B(n3186), .Z(n3188) );
  XOR U3070 ( .A(n3189), .B(n3190), .Z(n3186) );
  AND U3071 ( .A(n31), .B(n3191), .Z(n3190) );
  XNOR U3072 ( .A(p_input[113]), .B(n3189), .Z(n3191) );
  XOR U3073 ( .A(n3192), .B(n3193), .Z(n3189) );
  AND U3074 ( .A(n35), .B(n3194), .Z(n3193) );
  XNOR U3075 ( .A(p_input[129]), .B(n3192), .Z(n3194) );
  XOR U3076 ( .A(n3195), .B(n3196), .Z(n3192) );
  AND U3077 ( .A(n39), .B(n3197), .Z(n3196) );
  XNOR U3078 ( .A(p_input[145]), .B(n3195), .Z(n3197) );
  XOR U3079 ( .A(n3198), .B(n3199), .Z(n3195) );
  AND U3080 ( .A(n43), .B(n3200), .Z(n3199) );
  XNOR U3081 ( .A(p_input[161]), .B(n3198), .Z(n3200) );
  XOR U3082 ( .A(n3201), .B(n3202), .Z(n3198) );
  AND U3083 ( .A(n47), .B(n3203), .Z(n3202) );
  XNOR U3084 ( .A(p_input[177]), .B(n3201), .Z(n3203) );
  XOR U3085 ( .A(n3204), .B(n3205), .Z(n3201) );
  AND U3086 ( .A(n51), .B(n3206), .Z(n3205) );
  XNOR U3087 ( .A(p_input[193]), .B(n3204), .Z(n3206) );
  XOR U3088 ( .A(n3207), .B(n3208), .Z(n3204) );
  AND U3089 ( .A(n55), .B(n3209), .Z(n3208) );
  XNOR U3090 ( .A(p_input[209]), .B(n3207), .Z(n3209) );
  XOR U3091 ( .A(n3210), .B(n3211), .Z(n3207) );
  AND U3092 ( .A(n59), .B(n3212), .Z(n3211) );
  XNOR U3093 ( .A(p_input[225]), .B(n3210), .Z(n3212) );
  XOR U3094 ( .A(n3213), .B(n3214), .Z(n3210) );
  AND U3095 ( .A(n63), .B(n3215), .Z(n3214) );
  XNOR U3096 ( .A(p_input[241]), .B(n3213), .Z(n3215) );
  XOR U3097 ( .A(n3216), .B(n3217), .Z(n3213) );
  AND U3098 ( .A(n67), .B(n3218), .Z(n3217) );
  XNOR U3099 ( .A(p_input[257]), .B(n3216), .Z(n3218) );
  XOR U3100 ( .A(n3219), .B(n3220), .Z(n3216) );
  AND U3101 ( .A(n71), .B(n3221), .Z(n3220) );
  XNOR U3102 ( .A(p_input[273]), .B(n3219), .Z(n3221) );
  XOR U3103 ( .A(n3222), .B(n3223), .Z(n3219) );
  AND U3104 ( .A(n75), .B(n3224), .Z(n3223) );
  XNOR U3105 ( .A(p_input[289]), .B(n3222), .Z(n3224) );
  XOR U3106 ( .A(n3225), .B(n3226), .Z(n3222) );
  AND U3107 ( .A(n79), .B(n3227), .Z(n3226) );
  XNOR U3108 ( .A(p_input[305]), .B(n3225), .Z(n3227) );
  XOR U3109 ( .A(n3228), .B(n3229), .Z(n3225) );
  AND U3110 ( .A(n83), .B(n3230), .Z(n3229) );
  XNOR U3111 ( .A(p_input[321]), .B(n3228), .Z(n3230) );
  XOR U3112 ( .A(n3231), .B(n3232), .Z(n3228) );
  AND U3113 ( .A(n87), .B(n3233), .Z(n3232) );
  XNOR U3114 ( .A(p_input[337]), .B(n3231), .Z(n3233) );
  XOR U3115 ( .A(n3234), .B(n3235), .Z(n3231) );
  AND U3116 ( .A(n91), .B(n3236), .Z(n3235) );
  XNOR U3117 ( .A(p_input[353]), .B(n3234), .Z(n3236) );
  XOR U3118 ( .A(n3237), .B(n3238), .Z(n3234) );
  AND U3119 ( .A(n95), .B(n3239), .Z(n3238) );
  XNOR U3120 ( .A(p_input[369]), .B(n3237), .Z(n3239) );
  XOR U3121 ( .A(n3240), .B(n3241), .Z(n3237) );
  AND U3122 ( .A(n99), .B(n3242), .Z(n3241) );
  XNOR U3123 ( .A(p_input[385]), .B(n3240), .Z(n3242) );
  XOR U3124 ( .A(n3243), .B(n3244), .Z(n3240) );
  AND U3125 ( .A(n103), .B(n3245), .Z(n3244) );
  XNOR U3126 ( .A(p_input[401]), .B(n3243), .Z(n3245) );
  XOR U3127 ( .A(n3246), .B(n3247), .Z(n3243) );
  AND U3128 ( .A(n107), .B(n3248), .Z(n3247) );
  XNOR U3129 ( .A(p_input[417]), .B(n3246), .Z(n3248) );
  XOR U3130 ( .A(n3249), .B(n3250), .Z(n3246) );
  AND U3131 ( .A(n111), .B(n3251), .Z(n3250) );
  XNOR U3132 ( .A(p_input[433]), .B(n3249), .Z(n3251) );
  XOR U3133 ( .A(n3252), .B(n3253), .Z(n3249) );
  AND U3134 ( .A(n115), .B(n3254), .Z(n3253) );
  XNOR U3135 ( .A(p_input[449]), .B(n3252), .Z(n3254) );
  XOR U3136 ( .A(n3255), .B(n3256), .Z(n3252) );
  AND U3137 ( .A(n119), .B(n3257), .Z(n3256) );
  XNOR U3138 ( .A(p_input[465]), .B(n3255), .Z(n3257) );
  XOR U3139 ( .A(n3258), .B(n3259), .Z(n3255) );
  AND U3140 ( .A(n123), .B(n3260), .Z(n3259) );
  XNOR U3141 ( .A(p_input[481]), .B(n3258), .Z(n3260) );
  XOR U3142 ( .A(n3261), .B(n3262), .Z(n3258) );
  AND U3143 ( .A(n127), .B(n3263), .Z(n3262) );
  XNOR U3144 ( .A(p_input[497]), .B(n3261), .Z(n3263) );
  XOR U3145 ( .A(n3264), .B(n3265), .Z(n3261) );
  AND U3146 ( .A(n131), .B(n3266), .Z(n3265) );
  XNOR U3147 ( .A(p_input[513]), .B(n3264), .Z(n3266) );
  XOR U3148 ( .A(n3267), .B(n3268), .Z(n3264) );
  AND U3149 ( .A(n135), .B(n3269), .Z(n3268) );
  XNOR U3150 ( .A(p_input[529]), .B(n3267), .Z(n3269) );
  XOR U3151 ( .A(n3270), .B(n3271), .Z(n3267) );
  AND U3152 ( .A(n139), .B(n3272), .Z(n3271) );
  XNOR U3153 ( .A(p_input[545]), .B(n3270), .Z(n3272) );
  XOR U3154 ( .A(n3273), .B(n3274), .Z(n3270) );
  AND U3155 ( .A(n143), .B(n3275), .Z(n3274) );
  XNOR U3156 ( .A(p_input[561]), .B(n3273), .Z(n3275) );
  XOR U3157 ( .A(n3276), .B(n3277), .Z(n3273) );
  AND U3158 ( .A(n147), .B(n3278), .Z(n3277) );
  XNOR U3159 ( .A(p_input[577]), .B(n3276), .Z(n3278) );
  XOR U3160 ( .A(n3279), .B(n3280), .Z(n3276) );
  AND U3161 ( .A(n151), .B(n3281), .Z(n3280) );
  XNOR U3162 ( .A(p_input[593]), .B(n3279), .Z(n3281) );
  XOR U3163 ( .A(n3282), .B(n3283), .Z(n3279) );
  AND U3164 ( .A(n155), .B(n3284), .Z(n3283) );
  XNOR U3165 ( .A(p_input[609]), .B(n3282), .Z(n3284) );
  XOR U3166 ( .A(n3285), .B(n3286), .Z(n3282) );
  AND U3167 ( .A(n159), .B(n3287), .Z(n3286) );
  XNOR U3168 ( .A(p_input[625]), .B(n3285), .Z(n3287) );
  XOR U3169 ( .A(n3288), .B(n3289), .Z(n3285) );
  AND U3170 ( .A(n163), .B(n3290), .Z(n3289) );
  XNOR U3171 ( .A(p_input[641]), .B(n3288), .Z(n3290) );
  XOR U3172 ( .A(n3291), .B(n3292), .Z(n3288) );
  AND U3173 ( .A(n167), .B(n3293), .Z(n3292) );
  XNOR U3174 ( .A(p_input[657]), .B(n3291), .Z(n3293) );
  XOR U3175 ( .A(n3294), .B(n3295), .Z(n3291) );
  AND U3176 ( .A(n171), .B(n3296), .Z(n3295) );
  XNOR U3177 ( .A(p_input[673]), .B(n3294), .Z(n3296) );
  XOR U3178 ( .A(n3297), .B(n3298), .Z(n3294) );
  AND U3179 ( .A(n175), .B(n3299), .Z(n3298) );
  XNOR U3180 ( .A(p_input[689]), .B(n3297), .Z(n3299) );
  XOR U3181 ( .A(n3300), .B(n3301), .Z(n3297) );
  AND U3182 ( .A(n179), .B(n3302), .Z(n3301) );
  XNOR U3183 ( .A(p_input[705]), .B(n3300), .Z(n3302) );
  XOR U3184 ( .A(n3303), .B(n3304), .Z(n3300) );
  AND U3185 ( .A(n183), .B(n3305), .Z(n3304) );
  XNOR U3186 ( .A(p_input[721]), .B(n3303), .Z(n3305) );
  XOR U3187 ( .A(n3306), .B(n3307), .Z(n3303) );
  AND U3188 ( .A(n187), .B(n3308), .Z(n3307) );
  XNOR U3189 ( .A(p_input[737]), .B(n3306), .Z(n3308) );
  XOR U3190 ( .A(n3309), .B(n3310), .Z(n3306) );
  AND U3191 ( .A(n191), .B(n3311), .Z(n3310) );
  XNOR U3192 ( .A(p_input[753]), .B(n3309), .Z(n3311) );
  XOR U3193 ( .A(n3312), .B(n3313), .Z(n3309) );
  AND U3194 ( .A(n195), .B(n3314), .Z(n3313) );
  XNOR U3195 ( .A(p_input[769]), .B(n3312), .Z(n3314) );
  XOR U3196 ( .A(n3315), .B(n3316), .Z(n3312) );
  AND U3197 ( .A(n199), .B(n3317), .Z(n3316) );
  XNOR U3198 ( .A(p_input[785]), .B(n3315), .Z(n3317) );
  XOR U3199 ( .A(n3318), .B(n3319), .Z(n3315) );
  AND U3200 ( .A(n203), .B(n3320), .Z(n3319) );
  XNOR U3201 ( .A(p_input[801]), .B(n3318), .Z(n3320) );
  XOR U3202 ( .A(n3321), .B(n3322), .Z(n3318) );
  AND U3203 ( .A(n207), .B(n3323), .Z(n3322) );
  XNOR U3204 ( .A(p_input[817]), .B(n3321), .Z(n3323) );
  XOR U3205 ( .A(n3324), .B(n3325), .Z(n3321) );
  AND U3206 ( .A(n211), .B(n3326), .Z(n3325) );
  XNOR U3207 ( .A(p_input[833]), .B(n3324), .Z(n3326) );
  XOR U3208 ( .A(n3327), .B(n3328), .Z(n3324) );
  AND U3209 ( .A(n215), .B(n3329), .Z(n3328) );
  XNOR U3210 ( .A(p_input[849]), .B(n3327), .Z(n3329) );
  XOR U3211 ( .A(n3330), .B(n3331), .Z(n3327) );
  AND U3212 ( .A(n219), .B(n3332), .Z(n3331) );
  XNOR U3213 ( .A(p_input[865]), .B(n3330), .Z(n3332) );
  XOR U3214 ( .A(n3333), .B(n3334), .Z(n3330) );
  AND U3215 ( .A(n223), .B(n3335), .Z(n3334) );
  XNOR U3216 ( .A(p_input[881]), .B(n3333), .Z(n3335) );
  XOR U3217 ( .A(n3336), .B(n3337), .Z(n3333) );
  AND U3218 ( .A(n227), .B(n3338), .Z(n3337) );
  XNOR U3219 ( .A(p_input[897]), .B(n3336), .Z(n3338) );
  XOR U3220 ( .A(n3339), .B(n3340), .Z(n3336) );
  AND U3221 ( .A(n231), .B(n3341), .Z(n3340) );
  XNOR U3222 ( .A(p_input[913]), .B(n3339), .Z(n3341) );
  XOR U3223 ( .A(n3342), .B(n3343), .Z(n3339) );
  AND U3224 ( .A(n235), .B(n3344), .Z(n3343) );
  XNOR U3225 ( .A(p_input[929]), .B(n3342), .Z(n3344) );
  XOR U3226 ( .A(n3345), .B(n3346), .Z(n3342) );
  AND U3227 ( .A(n239), .B(n3347), .Z(n3346) );
  XNOR U3228 ( .A(p_input[945]), .B(n3345), .Z(n3347) );
  XOR U3229 ( .A(n3348), .B(n3349), .Z(n3345) );
  AND U3230 ( .A(n243), .B(n3350), .Z(n3349) );
  XNOR U3231 ( .A(p_input[961]), .B(n3348), .Z(n3350) );
  XOR U3232 ( .A(n3351), .B(n3352), .Z(n3348) );
  AND U3233 ( .A(n247), .B(n3353), .Z(n3352) );
  XNOR U3234 ( .A(p_input[977]), .B(n3351), .Z(n3353) );
  XOR U3235 ( .A(n3354), .B(n3355), .Z(n3351) );
  AND U3236 ( .A(n251), .B(n3356), .Z(n3355) );
  XNOR U3237 ( .A(p_input[993]), .B(n3354), .Z(n3356) );
  XOR U3238 ( .A(n3357), .B(n3358), .Z(n3354) );
  AND U3239 ( .A(n255), .B(n3359), .Z(n3358) );
  XNOR U3240 ( .A(p_input[1009]), .B(n3357), .Z(n3359) );
  XOR U3241 ( .A(n3360), .B(n3361), .Z(n3357) );
  AND U3242 ( .A(n259), .B(n3362), .Z(n3361) );
  XNOR U3243 ( .A(p_input[1025]), .B(n3360), .Z(n3362) );
  XOR U3244 ( .A(n3363), .B(n3364), .Z(n3360) );
  AND U3245 ( .A(n263), .B(n3365), .Z(n3364) );
  XNOR U3246 ( .A(p_input[1041]), .B(n3363), .Z(n3365) );
  XOR U3247 ( .A(n3366), .B(n3367), .Z(n3363) );
  AND U3248 ( .A(n267), .B(n3368), .Z(n3367) );
  XNOR U3249 ( .A(p_input[1057]), .B(n3366), .Z(n3368) );
  XOR U3250 ( .A(n3369), .B(n3370), .Z(n3366) );
  AND U3251 ( .A(n271), .B(n3371), .Z(n3370) );
  XNOR U3252 ( .A(p_input[1073]), .B(n3369), .Z(n3371) );
  XOR U3253 ( .A(n3372), .B(n3373), .Z(n3369) );
  AND U3254 ( .A(n275), .B(n3374), .Z(n3373) );
  XNOR U3255 ( .A(p_input[1089]), .B(n3372), .Z(n3374) );
  XOR U3256 ( .A(n3375), .B(n3376), .Z(n3372) );
  AND U3257 ( .A(n279), .B(n3377), .Z(n3376) );
  XNOR U3258 ( .A(p_input[1105]), .B(n3375), .Z(n3377) );
  XOR U3259 ( .A(n3378), .B(n3379), .Z(n3375) );
  AND U3260 ( .A(n283), .B(n3380), .Z(n3379) );
  XNOR U3261 ( .A(p_input[1121]), .B(n3378), .Z(n3380) );
  XOR U3262 ( .A(n3381), .B(n3382), .Z(n3378) );
  AND U3263 ( .A(n287), .B(n3383), .Z(n3382) );
  XNOR U3264 ( .A(p_input[1137]), .B(n3381), .Z(n3383) );
  XOR U3265 ( .A(n3384), .B(n3385), .Z(n3381) );
  AND U3266 ( .A(n291), .B(n3386), .Z(n3385) );
  XNOR U3267 ( .A(p_input[1153]), .B(n3384), .Z(n3386) );
  XOR U3268 ( .A(n3387), .B(n3388), .Z(n3384) );
  AND U3269 ( .A(n295), .B(n3389), .Z(n3388) );
  XNOR U3270 ( .A(p_input[1169]), .B(n3387), .Z(n3389) );
  XOR U3271 ( .A(n3390), .B(n3391), .Z(n3387) );
  AND U3272 ( .A(n299), .B(n3392), .Z(n3391) );
  XNOR U3273 ( .A(p_input[1185]), .B(n3390), .Z(n3392) );
  XOR U3274 ( .A(n3393), .B(n3394), .Z(n3390) );
  AND U3275 ( .A(n303), .B(n3395), .Z(n3394) );
  XNOR U3276 ( .A(p_input[1201]), .B(n3393), .Z(n3395) );
  XOR U3277 ( .A(n3396), .B(n3397), .Z(n3393) );
  AND U3278 ( .A(n307), .B(n3398), .Z(n3397) );
  XNOR U3279 ( .A(p_input[1217]), .B(n3396), .Z(n3398) );
  XOR U3280 ( .A(n3399), .B(n3400), .Z(n3396) );
  AND U3281 ( .A(n311), .B(n3401), .Z(n3400) );
  XNOR U3282 ( .A(p_input[1233]), .B(n3399), .Z(n3401) );
  XOR U3283 ( .A(n3402), .B(n3403), .Z(n3399) );
  AND U3284 ( .A(n315), .B(n3404), .Z(n3403) );
  XNOR U3285 ( .A(p_input[1249]), .B(n3402), .Z(n3404) );
  XOR U3286 ( .A(n3405), .B(n3406), .Z(n3402) );
  AND U3287 ( .A(n319), .B(n3407), .Z(n3406) );
  XNOR U3288 ( .A(p_input[1265]), .B(n3405), .Z(n3407) );
  XOR U3289 ( .A(n3408), .B(n3409), .Z(n3405) );
  AND U3290 ( .A(n323), .B(n3410), .Z(n3409) );
  XNOR U3291 ( .A(p_input[1281]), .B(n3408), .Z(n3410) );
  XOR U3292 ( .A(n3411), .B(n3412), .Z(n3408) );
  AND U3293 ( .A(n327), .B(n3413), .Z(n3412) );
  XNOR U3294 ( .A(p_input[1297]), .B(n3411), .Z(n3413) );
  XOR U3295 ( .A(n3414), .B(n3415), .Z(n3411) );
  AND U3296 ( .A(n331), .B(n3416), .Z(n3415) );
  XNOR U3297 ( .A(p_input[1313]), .B(n3414), .Z(n3416) );
  XOR U3298 ( .A(n3417), .B(n3418), .Z(n3414) );
  AND U3299 ( .A(n335), .B(n3419), .Z(n3418) );
  XNOR U3300 ( .A(p_input[1329]), .B(n3417), .Z(n3419) );
  XOR U3301 ( .A(n3420), .B(n3421), .Z(n3417) );
  AND U3302 ( .A(n339), .B(n3422), .Z(n3421) );
  XNOR U3303 ( .A(p_input[1345]), .B(n3420), .Z(n3422) );
  XOR U3304 ( .A(n3423), .B(n3424), .Z(n3420) );
  AND U3305 ( .A(n343), .B(n3425), .Z(n3424) );
  XNOR U3306 ( .A(p_input[1361]), .B(n3423), .Z(n3425) );
  XOR U3307 ( .A(n3426), .B(n3427), .Z(n3423) );
  AND U3308 ( .A(n347), .B(n3428), .Z(n3427) );
  XNOR U3309 ( .A(p_input[1377]), .B(n3426), .Z(n3428) );
  XOR U3310 ( .A(n3429), .B(n3430), .Z(n3426) );
  AND U3311 ( .A(n351), .B(n3431), .Z(n3430) );
  XNOR U3312 ( .A(p_input[1393]), .B(n3429), .Z(n3431) );
  XOR U3313 ( .A(n3432), .B(n3433), .Z(n3429) );
  AND U3314 ( .A(n355), .B(n3434), .Z(n3433) );
  XNOR U3315 ( .A(p_input[1409]), .B(n3432), .Z(n3434) );
  XOR U3316 ( .A(n3435), .B(n3436), .Z(n3432) );
  AND U3317 ( .A(n359), .B(n3437), .Z(n3436) );
  XNOR U3318 ( .A(p_input[1425]), .B(n3435), .Z(n3437) );
  XOR U3319 ( .A(n3438), .B(n3439), .Z(n3435) );
  AND U3320 ( .A(n363), .B(n3440), .Z(n3439) );
  XNOR U3321 ( .A(p_input[1441]), .B(n3438), .Z(n3440) );
  XOR U3322 ( .A(n3441), .B(n3442), .Z(n3438) );
  AND U3323 ( .A(n367), .B(n3443), .Z(n3442) );
  XNOR U3324 ( .A(p_input[1457]), .B(n3441), .Z(n3443) );
  XOR U3325 ( .A(n3444), .B(n3445), .Z(n3441) );
  AND U3326 ( .A(n371), .B(n3446), .Z(n3445) );
  XNOR U3327 ( .A(p_input[1473]), .B(n3444), .Z(n3446) );
  XOR U3328 ( .A(n3447), .B(n3448), .Z(n3444) );
  AND U3329 ( .A(n375), .B(n3449), .Z(n3448) );
  XNOR U3330 ( .A(p_input[1489]), .B(n3447), .Z(n3449) );
  XOR U3331 ( .A(n3450), .B(n3451), .Z(n3447) );
  AND U3332 ( .A(n379), .B(n3452), .Z(n3451) );
  XNOR U3333 ( .A(p_input[1505]), .B(n3450), .Z(n3452) );
  XOR U3334 ( .A(n3453), .B(n3454), .Z(n3450) );
  AND U3335 ( .A(n383), .B(n3455), .Z(n3454) );
  XNOR U3336 ( .A(p_input[1521]), .B(n3453), .Z(n3455) );
  XOR U3337 ( .A(n3456), .B(n3457), .Z(n3453) );
  AND U3338 ( .A(n387), .B(n3458), .Z(n3457) );
  XNOR U3339 ( .A(p_input[1537]), .B(n3456), .Z(n3458) );
  XOR U3340 ( .A(n3459), .B(n3460), .Z(n3456) );
  AND U3341 ( .A(n391), .B(n3461), .Z(n3460) );
  XNOR U3342 ( .A(p_input[1553]), .B(n3459), .Z(n3461) );
  XOR U3343 ( .A(n3462), .B(n3463), .Z(n3459) );
  AND U3344 ( .A(n395), .B(n3464), .Z(n3463) );
  XNOR U3345 ( .A(p_input[1569]), .B(n3462), .Z(n3464) );
  XOR U3346 ( .A(n3465), .B(n3466), .Z(n3462) );
  AND U3347 ( .A(n399), .B(n3467), .Z(n3466) );
  XNOR U3348 ( .A(p_input[1585]), .B(n3465), .Z(n3467) );
  XOR U3349 ( .A(n3468), .B(n3469), .Z(n3465) );
  AND U3350 ( .A(n403), .B(n3470), .Z(n3469) );
  XNOR U3351 ( .A(p_input[1601]), .B(n3468), .Z(n3470) );
  XOR U3352 ( .A(n3471), .B(n3472), .Z(n3468) );
  AND U3353 ( .A(n407), .B(n3473), .Z(n3472) );
  XNOR U3354 ( .A(p_input[1617]), .B(n3471), .Z(n3473) );
  XOR U3355 ( .A(n3474), .B(n3475), .Z(n3471) );
  AND U3356 ( .A(n411), .B(n3476), .Z(n3475) );
  XNOR U3357 ( .A(p_input[1633]), .B(n3474), .Z(n3476) );
  XOR U3358 ( .A(n3477), .B(n3478), .Z(n3474) );
  AND U3359 ( .A(n415), .B(n3479), .Z(n3478) );
  XNOR U3360 ( .A(p_input[1649]), .B(n3477), .Z(n3479) );
  XOR U3361 ( .A(n3480), .B(n3481), .Z(n3477) );
  AND U3362 ( .A(n419), .B(n3482), .Z(n3481) );
  XNOR U3363 ( .A(p_input[1665]), .B(n3480), .Z(n3482) );
  XOR U3364 ( .A(n3483), .B(n3484), .Z(n3480) );
  AND U3365 ( .A(n423), .B(n3485), .Z(n3484) );
  XNOR U3366 ( .A(p_input[1681]), .B(n3483), .Z(n3485) );
  XOR U3367 ( .A(n3486), .B(n3487), .Z(n3483) );
  AND U3368 ( .A(n427), .B(n3488), .Z(n3487) );
  XNOR U3369 ( .A(p_input[1697]), .B(n3486), .Z(n3488) );
  XOR U3370 ( .A(n3489), .B(n3490), .Z(n3486) );
  AND U3371 ( .A(n431), .B(n3491), .Z(n3490) );
  XNOR U3372 ( .A(p_input[1713]), .B(n3489), .Z(n3491) );
  XOR U3373 ( .A(n3492), .B(n3493), .Z(n3489) );
  AND U3374 ( .A(n435), .B(n3494), .Z(n3493) );
  XNOR U3375 ( .A(p_input[1729]), .B(n3492), .Z(n3494) );
  XOR U3376 ( .A(n3495), .B(n3496), .Z(n3492) );
  AND U3377 ( .A(n439), .B(n3497), .Z(n3496) );
  XNOR U3378 ( .A(p_input[1745]), .B(n3495), .Z(n3497) );
  XOR U3379 ( .A(n3498), .B(n3499), .Z(n3495) );
  AND U3380 ( .A(n443), .B(n3500), .Z(n3499) );
  XNOR U3381 ( .A(p_input[1761]), .B(n3498), .Z(n3500) );
  XOR U3382 ( .A(n3501), .B(n3502), .Z(n3498) );
  AND U3383 ( .A(n447), .B(n3503), .Z(n3502) );
  XNOR U3384 ( .A(p_input[1777]), .B(n3501), .Z(n3503) );
  XOR U3385 ( .A(n3504), .B(n3505), .Z(n3501) );
  AND U3386 ( .A(n451), .B(n3506), .Z(n3505) );
  XNOR U3387 ( .A(p_input[1793]), .B(n3504), .Z(n3506) );
  XOR U3388 ( .A(n3507), .B(n3508), .Z(n3504) );
  AND U3389 ( .A(n455), .B(n3509), .Z(n3508) );
  XNOR U3390 ( .A(p_input[1809]), .B(n3507), .Z(n3509) );
  XOR U3391 ( .A(n3510), .B(n3511), .Z(n3507) );
  AND U3392 ( .A(n459), .B(n3512), .Z(n3511) );
  XNOR U3393 ( .A(p_input[1825]), .B(n3510), .Z(n3512) );
  XOR U3394 ( .A(n3513), .B(n3514), .Z(n3510) );
  AND U3395 ( .A(n463), .B(n3515), .Z(n3514) );
  XNOR U3396 ( .A(p_input[1841]), .B(n3513), .Z(n3515) );
  XOR U3397 ( .A(n3516), .B(n3517), .Z(n3513) );
  AND U3398 ( .A(n467), .B(n3518), .Z(n3517) );
  XNOR U3399 ( .A(p_input[1857]), .B(n3516), .Z(n3518) );
  XOR U3400 ( .A(n3519), .B(n3520), .Z(n3516) );
  AND U3401 ( .A(n471), .B(n3521), .Z(n3520) );
  XNOR U3402 ( .A(p_input[1873]), .B(n3519), .Z(n3521) );
  XOR U3403 ( .A(n3522), .B(n3523), .Z(n3519) );
  AND U3404 ( .A(n475), .B(n3524), .Z(n3523) );
  XNOR U3405 ( .A(p_input[1889]), .B(n3522), .Z(n3524) );
  XOR U3406 ( .A(n3525), .B(n3526), .Z(n3522) );
  AND U3407 ( .A(n479), .B(n3527), .Z(n3526) );
  XNOR U3408 ( .A(p_input[1905]), .B(n3525), .Z(n3527) );
  XOR U3409 ( .A(n3528), .B(n3529), .Z(n3525) );
  AND U3410 ( .A(n483), .B(n3530), .Z(n3529) );
  XNOR U3411 ( .A(p_input[1921]), .B(n3528), .Z(n3530) );
  XOR U3412 ( .A(n3531), .B(n3532), .Z(n3528) );
  AND U3413 ( .A(n487), .B(n3533), .Z(n3532) );
  XNOR U3414 ( .A(p_input[1937]), .B(n3531), .Z(n3533) );
  XOR U3415 ( .A(n3534), .B(n3535), .Z(n3531) );
  AND U3416 ( .A(n491), .B(n3536), .Z(n3535) );
  XNOR U3417 ( .A(p_input[1953]), .B(n3534), .Z(n3536) );
  XOR U3418 ( .A(n3537), .B(n3538), .Z(n3534) );
  AND U3419 ( .A(n495), .B(n3539), .Z(n3538) );
  XNOR U3420 ( .A(p_input[1969]), .B(n3537), .Z(n3539) );
  XOR U3421 ( .A(n3540), .B(n3541), .Z(n3537) );
  AND U3422 ( .A(n499), .B(n3542), .Z(n3541) );
  XNOR U3423 ( .A(p_input[1985]), .B(n3540), .Z(n3542) );
  XNOR U3424 ( .A(n3543), .B(n3544), .Z(n3540) );
  AND U3425 ( .A(n503), .B(n3545), .Z(n3544) );
  XOR U3426 ( .A(p_input[2001]), .B(n3543), .Z(n3545) );
  XOR U3427 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n3546), .Z(n3543) );
  AND U3428 ( .A(n506), .B(n3547), .Z(n3546) );
  XOR U3429 ( .A(p_input[2017]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n3547)
         );
  XNOR U3430 ( .A(n3548), .B(n3549), .Z(o[15]) );
  AND U3431 ( .A(n3), .B(n3550), .Z(n3548) );
  XNOR U3432 ( .A(p_input[15]), .B(n3549), .Z(n3550) );
  XOR U3433 ( .A(n3551), .B(n3552), .Z(n3549) );
  AND U3434 ( .A(n7), .B(n3553), .Z(n3552) );
  XNOR U3435 ( .A(p_input[31]), .B(n3551), .Z(n3553) );
  XOR U3436 ( .A(n3554), .B(n3555), .Z(n3551) );
  AND U3437 ( .A(n11), .B(n3556), .Z(n3555) );
  XNOR U3438 ( .A(p_input[47]), .B(n3554), .Z(n3556) );
  XOR U3439 ( .A(n3557), .B(n3558), .Z(n3554) );
  AND U3440 ( .A(n15), .B(n3559), .Z(n3558) );
  XNOR U3441 ( .A(p_input[63]), .B(n3557), .Z(n3559) );
  XOR U3442 ( .A(n3560), .B(n3561), .Z(n3557) );
  AND U3443 ( .A(n19), .B(n3562), .Z(n3561) );
  XNOR U3444 ( .A(p_input[79]), .B(n3560), .Z(n3562) );
  XOR U3445 ( .A(n3563), .B(n3564), .Z(n3560) );
  AND U3446 ( .A(n23), .B(n3565), .Z(n3564) );
  XNOR U3447 ( .A(p_input[95]), .B(n3563), .Z(n3565) );
  XOR U3448 ( .A(n3566), .B(n3567), .Z(n3563) );
  AND U3449 ( .A(n27), .B(n3568), .Z(n3567) );
  XNOR U3450 ( .A(p_input[111]), .B(n3566), .Z(n3568) );
  XOR U3451 ( .A(n3569), .B(n3570), .Z(n3566) );
  AND U3452 ( .A(n31), .B(n3571), .Z(n3570) );
  XNOR U3453 ( .A(p_input[127]), .B(n3569), .Z(n3571) );
  XOR U3454 ( .A(n3572), .B(n3573), .Z(n3569) );
  AND U3455 ( .A(n35), .B(n3574), .Z(n3573) );
  XNOR U3456 ( .A(p_input[143]), .B(n3572), .Z(n3574) );
  XOR U3457 ( .A(n3575), .B(n3576), .Z(n3572) );
  AND U3458 ( .A(n39), .B(n3577), .Z(n3576) );
  XNOR U3459 ( .A(p_input[159]), .B(n3575), .Z(n3577) );
  XOR U3460 ( .A(n3578), .B(n3579), .Z(n3575) );
  AND U3461 ( .A(n43), .B(n3580), .Z(n3579) );
  XNOR U3462 ( .A(p_input[175]), .B(n3578), .Z(n3580) );
  XOR U3463 ( .A(n3581), .B(n3582), .Z(n3578) );
  AND U3464 ( .A(n47), .B(n3583), .Z(n3582) );
  XNOR U3465 ( .A(p_input[191]), .B(n3581), .Z(n3583) );
  XOR U3466 ( .A(n3584), .B(n3585), .Z(n3581) );
  AND U3467 ( .A(n51), .B(n3586), .Z(n3585) );
  XNOR U3468 ( .A(p_input[207]), .B(n3584), .Z(n3586) );
  XOR U3469 ( .A(n3587), .B(n3588), .Z(n3584) );
  AND U3470 ( .A(n55), .B(n3589), .Z(n3588) );
  XNOR U3471 ( .A(p_input[223]), .B(n3587), .Z(n3589) );
  XOR U3472 ( .A(n3590), .B(n3591), .Z(n3587) );
  AND U3473 ( .A(n59), .B(n3592), .Z(n3591) );
  XNOR U3474 ( .A(p_input[239]), .B(n3590), .Z(n3592) );
  XOR U3475 ( .A(n3593), .B(n3594), .Z(n3590) );
  AND U3476 ( .A(n63), .B(n3595), .Z(n3594) );
  XNOR U3477 ( .A(p_input[255]), .B(n3593), .Z(n3595) );
  XOR U3478 ( .A(n3596), .B(n3597), .Z(n3593) );
  AND U3479 ( .A(n67), .B(n3598), .Z(n3597) );
  XNOR U3480 ( .A(p_input[271]), .B(n3596), .Z(n3598) );
  XOR U3481 ( .A(n3599), .B(n3600), .Z(n3596) );
  AND U3482 ( .A(n71), .B(n3601), .Z(n3600) );
  XNOR U3483 ( .A(p_input[287]), .B(n3599), .Z(n3601) );
  XOR U3484 ( .A(n3602), .B(n3603), .Z(n3599) );
  AND U3485 ( .A(n75), .B(n3604), .Z(n3603) );
  XNOR U3486 ( .A(p_input[303]), .B(n3602), .Z(n3604) );
  XOR U3487 ( .A(n3605), .B(n3606), .Z(n3602) );
  AND U3488 ( .A(n79), .B(n3607), .Z(n3606) );
  XNOR U3489 ( .A(p_input[319]), .B(n3605), .Z(n3607) );
  XOR U3490 ( .A(n3608), .B(n3609), .Z(n3605) );
  AND U3491 ( .A(n83), .B(n3610), .Z(n3609) );
  XNOR U3492 ( .A(p_input[335]), .B(n3608), .Z(n3610) );
  XOR U3493 ( .A(n3611), .B(n3612), .Z(n3608) );
  AND U3494 ( .A(n87), .B(n3613), .Z(n3612) );
  XNOR U3495 ( .A(p_input[351]), .B(n3611), .Z(n3613) );
  XOR U3496 ( .A(n3614), .B(n3615), .Z(n3611) );
  AND U3497 ( .A(n91), .B(n3616), .Z(n3615) );
  XNOR U3498 ( .A(p_input[367]), .B(n3614), .Z(n3616) );
  XOR U3499 ( .A(n3617), .B(n3618), .Z(n3614) );
  AND U3500 ( .A(n95), .B(n3619), .Z(n3618) );
  XNOR U3501 ( .A(p_input[383]), .B(n3617), .Z(n3619) );
  XOR U3502 ( .A(n3620), .B(n3621), .Z(n3617) );
  AND U3503 ( .A(n99), .B(n3622), .Z(n3621) );
  XNOR U3504 ( .A(p_input[399]), .B(n3620), .Z(n3622) );
  XOR U3505 ( .A(n3623), .B(n3624), .Z(n3620) );
  AND U3506 ( .A(n103), .B(n3625), .Z(n3624) );
  XNOR U3507 ( .A(p_input[415]), .B(n3623), .Z(n3625) );
  XOR U3508 ( .A(n3626), .B(n3627), .Z(n3623) );
  AND U3509 ( .A(n107), .B(n3628), .Z(n3627) );
  XNOR U3510 ( .A(p_input[431]), .B(n3626), .Z(n3628) );
  XOR U3511 ( .A(n3629), .B(n3630), .Z(n3626) );
  AND U3512 ( .A(n111), .B(n3631), .Z(n3630) );
  XNOR U3513 ( .A(p_input[447]), .B(n3629), .Z(n3631) );
  XOR U3514 ( .A(n3632), .B(n3633), .Z(n3629) );
  AND U3515 ( .A(n115), .B(n3634), .Z(n3633) );
  XNOR U3516 ( .A(p_input[463]), .B(n3632), .Z(n3634) );
  XOR U3517 ( .A(n3635), .B(n3636), .Z(n3632) );
  AND U3518 ( .A(n119), .B(n3637), .Z(n3636) );
  XNOR U3519 ( .A(p_input[479]), .B(n3635), .Z(n3637) );
  XOR U3520 ( .A(n3638), .B(n3639), .Z(n3635) );
  AND U3521 ( .A(n123), .B(n3640), .Z(n3639) );
  XNOR U3522 ( .A(p_input[495]), .B(n3638), .Z(n3640) );
  XOR U3523 ( .A(n3641), .B(n3642), .Z(n3638) );
  AND U3524 ( .A(n127), .B(n3643), .Z(n3642) );
  XNOR U3525 ( .A(p_input[511]), .B(n3641), .Z(n3643) );
  XOR U3526 ( .A(n3644), .B(n3645), .Z(n3641) );
  AND U3527 ( .A(n131), .B(n3646), .Z(n3645) );
  XNOR U3528 ( .A(p_input[527]), .B(n3644), .Z(n3646) );
  XOR U3529 ( .A(n3647), .B(n3648), .Z(n3644) );
  AND U3530 ( .A(n135), .B(n3649), .Z(n3648) );
  XNOR U3531 ( .A(p_input[543]), .B(n3647), .Z(n3649) );
  XOR U3532 ( .A(n3650), .B(n3651), .Z(n3647) );
  AND U3533 ( .A(n139), .B(n3652), .Z(n3651) );
  XNOR U3534 ( .A(p_input[559]), .B(n3650), .Z(n3652) );
  XOR U3535 ( .A(n3653), .B(n3654), .Z(n3650) );
  AND U3536 ( .A(n143), .B(n3655), .Z(n3654) );
  XNOR U3537 ( .A(p_input[575]), .B(n3653), .Z(n3655) );
  XOR U3538 ( .A(n3656), .B(n3657), .Z(n3653) );
  AND U3539 ( .A(n147), .B(n3658), .Z(n3657) );
  XNOR U3540 ( .A(p_input[591]), .B(n3656), .Z(n3658) );
  XOR U3541 ( .A(n3659), .B(n3660), .Z(n3656) );
  AND U3542 ( .A(n151), .B(n3661), .Z(n3660) );
  XNOR U3543 ( .A(p_input[607]), .B(n3659), .Z(n3661) );
  XOR U3544 ( .A(n3662), .B(n3663), .Z(n3659) );
  AND U3545 ( .A(n155), .B(n3664), .Z(n3663) );
  XNOR U3546 ( .A(p_input[623]), .B(n3662), .Z(n3664) );
  XOR U3547 ( .A(n3665), .B(n3666), .Z(n3662) );
  AND U3548 ( .A(n159), .B(n3667), .Z(n3666) );
  XNOR U3549 ( .A(p_input[639]), .B(n3665), .Z(n3667) );
  XOR U3550 ( .A(n3668), .B(n3669), .Z(n3665) );
  AND U3551 ( .A(n163), .B(n3670), .Z(n3669) );
  XNOR U3552 ( .A(p_input[655]), .B(n3668), .Z(n3670) );
  XOR U3553 ( .A(n3671), .B(n3672), .Z(n3668) );
  AND U3554 ( .A(n167), .B(n3673), .Z(n3672) );
  XNOR U3555 ( .A(p_input[671]), .B(n3671), .Z(n3673) );
  XOR U3556 ( .A(n3674), .B(n3675), .Z(n3671) );
  AND U3557 ( .A(n171), .B(n3676), .Z(n3675) );
  XNOR U3558 ( .A(p_input[687]), .B(n3674), .Z(n3676) );
  XOR U3559 ( .A(n3677), .B(n3678), .Z(n3674) );
  AND U3560 ( .A(n175), .B(n3679), .Z(n3678) );
  XNOR U3561 ( .A(p_input[703]), .B(n3677), .Z(n3679) );
  XOR U3562 ( .A(n3680), .B(n3681), .Z(n3677) );
  AND U3563 ( .A(n179), .B(n3682), .Z(n3681) );
  XNOR U3564 ( .A(p_input[719]), .B(n3680), .Z(n3682) );
  XOR U3565 ( .A(n3683), .B(n3684), .Z(n3680) );
  AND U3566 ( .A(n183), .B(n3685), .Z(n3684) );
  XNOR U3567 ( .A(p_input[735]), .B(n3683), .Z(n3685) );
  XOR U3568 ( .A(n3686), .B(n3687), .Z(n3683) );
  AND U3569 ( .A(n187), .B(n3688), .Z(n3687) );
  XNOR U3570 ( .A(p_input[751]), .B(n3686), .Z(n3688) );
  XOR U3571 ( .A(n3689), .B(n3690), .Z(n3686) );
  AND U3572 ( .A(n191), .B(n3691), .Z(n3690) );
  XNOR U3573 ( .A(p_input[767]), .B(n3689), .Z(n3691) );
  XOR U3574 ( .A(n3692), .B(n3693), .Z(n3689) );
  AND U3575 ( .A(n195), .B(n3694), .Z(n3693) );
  XNOR U3576 ( .A(p_input[783]), .B(n3692), .Z(n3694) );
  XOR U3577 ( .A(n3695), .B(n3696), .Z(n3692) );
  AND U3578 ( .A(n199), .B(n3697), .Z(n3696) );
  XNOR U3579 ( .A(p_input[799]), .B(n3695), .Z(n3697) );
  XOR U3580 ( .A(n3698), .B(n3699), .Z(n3695) );
  AND U3581 ( .A(n203), .B(n3700), .Z(n3699) );
  XNOR U3582 ( .A(p_input[815]), .B(n3698), .Z(n3700) );
  XOR U3583 ( .A(n3701), .B(n3702), .Z(n3698) );
  AND U3584 ( .A(n207), .B(n3703), .Z(n3702) );
  XNOR U3585 ( .A(p_input[831]), .B(n3701), .Z(n3703) );
  XOR U3586 ( .A(n3704), .B(n3705), .Z(n3701) );
  AND U3587 ( .A(n211), .B(n3706), .Z(n3705) );
  XNOR U3588 ( .A(p_input[847]), .B(n3704), .Z(n3706) );
  XOR U3589 ( .A(n3707), .B(n3708), .Z(n3704) );
  AND U3590 ( .A(n215), .B(n3709), .Z(n3708) );
  XNOR U3591 ( .A(p_input[863]), .B(n3707), .Z(n3709) );
  XOR U3592 ( .A(n3710), .B(n3711), .Z(n3707) );
  AND U3593 ( .A(n219), .B(n3712), .Z(n3711) );
  XNOR U3594 ( .A(p_input[879]), .B(n3710), .Z(n3712) );
  XOR U3595 ( .A(n3713), .B(n3714), .Z(n3710) );
  AND U3596 ( .A(n223), .B(n3715), .Z(n3714) );
  XNOR U3597 ( .A(p_input[895]), .B(n3713), .Z(n3715) );
  XOR U3598 ( .A(n3716), .B(n3717), .Z(n3713) );
  AND U3599 ( .A(n227), .B(n3718), .Z(n3717) );
  XNOR U3600 ( .A(p_input[911]), .B(n3716), .Z(n3718) );
  XOR U3601 ( .A(n3719), .B(n3720), .Z(n3716) );
  AND U3602 ( .A(n231), .B(n3721), .Z(n3720) );
  XNOR U3603 ( .A(p_input[927]), .B(n3719), .Z(n3721) );
  XOR U3604 ( .A(n3722), .B(n3723), .Z(n3719) );
  AND U3605 ( .A(n235), .B(n3724), .Z(n3723) );
  XNOR U3606 ( .A(p_input[943]), .B(n3722), .Z(n3724) );
  XOR U3607 ( .A(n3725), .B(n3726), .Z(n3722) );
  AND U3608 ( .A(n239), .B(n3727), .Z(n3726) );
  XNOR U3609 ( .A(p_input[959]), .B(n3725), .Z(n3727) );
  XOR U3610 ( .A(n3728), .B(n3729), .Z(n3725) );
  AND U3611 ( .A(n243), .B(n3730), .Z(n3729) );
  XNOR U3612 ( .A(p_input[975]), .B(n3728), .Z(n3730) );
  XOR U3613 ( .A(n3731), .B(n3732), .Z(n3728) );
  AND U3614 ( .A(n247), .B(n3733), .Z(n3732) );
  XNOR U3615 ( .A(p_input[991]), .B(n3731), .Z(n3733) );
  XOR U3616 ( .A(n3734), .B(n3735), .Z(n3731) );
  AND U3617 ( .A(n251), .B(n3736), .Z(n3735) );
  XNOR U3618 ( .A(p_input[1007]), .B(n3734), .Z(n3736) );
  XOR U3619 ( .A(n3737), .B(n3738), .Z(n3734) );
  AND U3620 ( .A(n255), .B(n3739), .Z(n3738) );
  XNOR U3621 ( .A(p_input[1023]), .B(n3737), .Z(n3739) );
  XOR U3622 ( .A(n3740), .B(n3741), .Z(n3737) );
  AND U3623 ( .A(n259), .B(n3742), .Z(n3741) );
  XNOR U3624 ( .A(p_input[1039]), .B(n3740), .Z(n3742) );
  XOR U3625 ( .A(n3743), .B(n3744), .Z(n3740) );
  AND U3626 ( .A(n263), .B(n3745), .Z(n3744) );
  XNOR U3627 ( .A(p_input[1055]), .B(n3743), .Z(n3745) );
  XOR U3628 ( .A(n3746), .B(n3747), .Z(n3743) );
  AND U3629 ( .A(n267), .B(n3748), .Z(n3747) );
  XNOR U3630 ( .A(p_input[1071]), .B(n3746), .Z(n3748) );
  XOR U3631 ( .A(n3749), .B(n3750), .Z(n3746) );
  AND U3632 ( .A(n271), .B(n3751), .Z(n3750) );
  XNOR U3633 ( .A(p_input[1087]), .B(n3749), .Z(n3751) );
  XOR U3634 ( .A(n3752), .B(n3753), .Z(n3749) );
  AND U3635 ( .A(n275), .B(n3754), .Z(n3753) );
  XNOR U3636 ( .A(p_input[1103]), .B(n3752), .Z(n3754) );
  XOR U3637 ( .A(n3755), .B(n3756), .Z(n3752) );
  AND U3638 ( .A(n279), .B(n3757), .Z(n3756) );
  XNOR U3639 ( .A(p_input[1119]), .B(n3755), .Z(n3757) );
  XOR U3640 ( .A(n3758), .B(n3759), .Z(n3755) );
  AND U3641 ( .A(n283), .B(n3760), .Z(n3759) );
  XNOR U3642 ( .A(p_input[1135]), .B(n3758), .Z(n3760) );
  XOR U3643 ( .A(n3761), .B(n3762), .Z(n3758) );
  AND U3644 ( .A(n287), .B(n3763), .Z(n3762) );
  XNOR U3645 ( .A(p_input[1151]), .B(n3761), .Z(n3763) );
  XOR U3646 ( .A(n3764), .B(n3765), .Z(n3761) );
  AND U3647 ( .A(n291), .B(n3766), .Z(n3765) );
  XNOR U3648 ( .A(p_input[1167]), .B(n3764), .Z(n3766) );
  XOR U3649 ( .A(n3767), .B(n3768), .Z(n3764) );
  AND U3650 ( .A(n295), .B(n3769), .Z(n3768) );
  XNOR U3651 ( .A(p_input[1183]), .B(n3767), .Z(n3769) );
  XOR U3652 ( .A(n3770), .B(n3771), .Z(n3767) );
  AND U3653 ( .A(n299), .B(n3772), .Z(n3771) );
  XNOR U3654 ( .A(p_input[1199]), .B(n3770), .Z(n3772) );
  XOR U3655 ( .A(n3773), .B(n3774), .Z(n3770) );
  AND U3656 ( .A(n303), .B(n3775), .Z(n3774) );
  XNOR U3657 ( .A(p_input[1215]), .B(n3773), .Z(n3775) );
  XOR U3658 ( .A(n3776), .B(n3777), .Z(n3773) );
  AND U3659 ( .A(n307), .B(n3778), .Z(n3777) );
  XNOR U3660 ( .A(p_input[1231]), .B(n3776), .Z(n3778) );
  XOR U3661 ( .A(n3779), .B(n3780), .Z(n3776) );
  AND U3662 ( .A(n311), .B(n3781), .Z(n3780) );
  XNOR U3663 ( .A(p_input[1247]), .B(n3779), .Z(n3781) );
  XOR U3664 ( .A(n3782), .B(n3783), .Z(n3779) );
  AND U3665 ( .A(n315), .B(n3784), .Z(n3783) );
  XNOR U3666 ( .A(p_input[1263]), .B(n3782), .Z(n3784) );
  XOR U3667 ( .A(n3785), .B(n3786), .Z(n3782) );
  AND U3668 ( .A(n319), .B(n3787), .Z(n3786) );
  XNOR U3669 ( .A(p_input[1279]), .B(n3785), .Z(n3787) );
  XOR U3670 ( .A(n3788), .B(n3789), .Z(n3785) );
  AND U3671 ( .A(n323), .B(n3790), .Z(n3789) );
  XNOR U3672 ( .A(p_input[1295]), .B(n3788), .Z(n3790) );
  XOR U3673 ( .A(n3791), .B(n3792), .Z(n3788) );
  AND U3674 ( .A(n327), .B(n3793), .Z(n3792) );
  XNOR U3675 ( .A(p_input[1311]), .B(n3791), .Z(n3793) );
  XOR U3676 ( .A(n3794), .B(n3795), .Z(n3791) );
  AND U3677 ( .A(n331), .B(n3796), .Z(n3795) );
  XNOR U3678 ( .A(p_input[1327]), .B(n3794), .Z(n3796) );
  XOR U3679 ( .A(n3797), .B(n3798), .Z(n3794) );
  AND U3680 ( .A(n335), .B(n3799), .Z(n3798) );
  XNOR U3681 ( .A(p_input[1343]), .B(n3797), .Z(n3799) );
  XOR U3682 ( .A(n3800), .B(n3801), .Z(n3797) );
  AND U3683 ( .A(n339), .B(n3802), .Z(n3801) );
  XNOR U3684 ( .A(p_input[1359]), .B(n3800), .Z(n3802) );
  XOR U3685 ( .A(n3803), .B(n3804), .Z(n3800) );
  AND U3686 ( .A(n343), .B(n3805), .Z(n3804) );
  XNOR U3687 ( .A(p_input[1375]), .B(n3803), .Z(n3805) );
  XOR U3688 ( .A(n3806), .B(n3807), .Z(n3803) );
  AND U3689 ( .A(n347), .B(n3808), .Z(n3807) );
  XNOR U3690 ( .A(p_input[1391]), .B(n3806), .Z(n3808) );
  XOR U3691 ( .A(n3809), .B(n3810), .Z(n3806) );
  AND U3692 ( .A(n351), .B(n3811), .Z(n3810) );
  XNOR U3693 ( .A(p_input[1407]), .B(n3809), .Z(n3811) );
  XOR U3694 ( .A(n3812), .B(n3813), .Z(n3809) );
  AND U3695 ( .A(n355), .B(n3814), .Z(n3813) );
  XNOR U3696 ( .A(p_input[1423]), .B(n3812), .Z(n3814) );
  XOR U3697 ( .A(n3815), .B(n3816), .Z(n3812) );
  AND U3698 ( .A(n359), .B(n3817), .Z(n3816) );
  XNOR U3699 ( .A(p_input[1439]), .B(n3815), .Z(n3817) );
  XOR U3700 ( .A(n3818), .B(n3819), .Z(n3815) );
  AND U3701 ( .A(n363), .B(n3820), .Z(n3819) );
  XNOR U3702 ( .A(p_input[1455]), .B(n3818), .Z(n3820) );
  XOR U3703 ( .A(n3821), .B(n3822), .Z(n3818) );
  AND U3704 ( .A(n367), .B(n3823), .Z(n3822) );
  XNOR U3705 ( .A(p_input[1471]), .B(n3821), .Z(n3823) );
  XOR U3706 ( .A(n3824), .B(n3825), .Z(n3821) );
  AND U3707 ( .A(n371), .B(n3826), .Z(n3825) );
  XNOR U3708 ( .A(p_input[1487]), .B(n3824), .Z(n3826) );
  XOR U3709 ( .A(n3827), .B(n3828), .Z(n3824) );
  AND U3710 ( .A(n375), .B(n3829), .Z(n3828) );
  XNOR U3711 ( .A(p_input[1503]), .B(n3827), .Z(n3829) );
  XOR U3712 ( .A(n3830), .B(n3831), .Z(n3827) );
  AND U3713 ( .A(n379), .B(n3832), .Z(n3831) );
  XNOR U3714 ( .A(p_input[1519]), .B(n3830), .Z(n3832) );
  XOR U3715 ( .A(n3833), .B(n3834), .Z(n3830) );
  AND U3716 ( .A(n383), .B(n3835), .Z(n3834) );
  XNOR U3717 ( .A(p_input[1535]), .B(n3833), .Z(n3835) );
  XOR U3718 ( .A(n3836), .B(n3837), .Z(n3833) );
  AND U3719 ( .A(n387), .B(n3838), .Z(n3837) );
  XNOR U3720 ( .A(p_input[1551]), .B(n3836), .Z(n3838) );
  XOR U3721 ( .A(n3839), .B(n3840), .Z(n3836) );
  AND U3722 ( .A(n391), .B(n3841), .Z(n3840) );
  XNOR U3723 ( .A(p_input[1567]), .B(n3839), .Z(n3841) );
  XOR U3724 ( .A(n3842), .B(n3843), .Z(n3839) );
  AND U3725 ( .A(n395), .B(n3844), .Z(n3843) );
  XNOR U3726 ( .A(p_input[1583]), .B(n3842), .Z(n3844) );
  XOR U3727 ( .A(n3845), .B(n3846), .Z(n3842) );
  AND U3728 ( .A(n399), .B(n3847), .Z(n3846) );
  XNOR U3729 ( .A(p_input[1599]), .B(n3845), .Z(n3847) );
  XOR U3730 ( .A(n3848), .B(n3849), .Z(n3845) );
  AND U3731 ( .A(n403), .B(n3850), .Z(n3849) );
  XNOR U3732 ( .A(p_input[1615]), .B(n3848), .Z(n3850) );
  XOR U3733 ( .A(n3851), .B(n3852), .Z(n3848) );
  AND U3734 ( .A(n407), .B(n3853), .Z(n3852) );
  XNOR U3735 ( .A(p_input[1631]), .B(n3851), .Z(n3853) );
  XOR U3736 ( .A(n3854), .B(n3855), .Z(n3851) );
  AND U3737 ( .A(n411), .B(n3856), .Z(n3855) );
  XNOR U3738 ( .A(p_input[1647]), .B(n3854), .Z(n3856) );
  XOR U3739 ( .A(n3857), .B(n3858), .Z(n3854) );
  AND U3740 ( .A(n415), .B(n3859), .Z(n3858) );
  XNOR U3741 ( .A(p_input[1663]), .B(n3857), .Z(n3859) );
  XOR U3742 ( .A(n3860), .B(n3861), .Z(n3857) );
  AND U3743 ( .A(n419), .B(n3862), .Z(n3861) );
  XNOR U3744 ( .A(p_input[1679]), .B(n3860), .Z(n3862) );
  XOR U3745 ( .A(n3863), .B(n3864), .Z(n3860) );
  AND U3746 ( .A(n423), .B(n3865), .Z(n3864) );
  XNOR U3747 ( .A(p_input[1695]), .B(n3863), .Z(n3865) );
  XOR U3748 ( .A(n3866), .B(n3867), .Z(n3863) );
  AND U3749 ( .A(n427), .B(n3868), .Z(n3867) );
  XNOR U3750 ( .A(p_input[1711]), .B(n3866), .Z(n3868) );
  XOR U3751 ( .A(n3869), .B(n3870), .Z(n3866) );
  AND U3752 ( .A(n431), .B(n3871), .Z(n3870) );
  XNOR U3753 ( .A(p_input[1727]), .B(n3869), .Z(n3871) );
  XOR U3754 ( .A(n3872), .B(n3873), .Z(n3869) );
  AND U3755 ( .A(n435), .B(n3874), .Z(n3873) );
  XNOR U3756 ( .A(p_input[1743]), .B(n3872), .Z(n3874) );
  XOR U3757 ( .A(n3875), .B(n3876), .Z(n3872) );
  AND U3758 ( .A(n439), .B(n3877), .Z(n3876) );
  XNOR U3759 ( .A(p_input[1759]), .B(n3875), .Z(n3877) );
  XOR U3760 ( .A(n3878), .B(n3879), .Z(n3875) );
  AND U3761 ( .A(n443), .B(n3880), .Z(n3879) );
  XNOR U3762 ( .A(p_input[1775]), .B(n3878), .Z(n3880) );
  XOR U3763 ( .A(n3881), .B(n3882), .Z(n3878) );
  AND U3764 ( .A(n447), .B(n3883), .Z(n3882) );
  XNOR U3765 ( .A(p_input[1791]), .B(n3881), .Z(n3883) );
  XOR U3766 ( .A(n3884), .B(n3885), .Z(n3881) );
  AND U3767 ( .A(n451), .B(n3886), .Z(n3885) );
  XNOR U3768 ( .A(p_input[1807]), .B(n3884), .Z(n3886) );
  XOR U3769 ( .A(n3887), .B(n3888), .Z(n3884) );
  AND U3770 ( .A(n455), .B(n3889), .Z(n3888) );
  XNOR U3771 ( .A(p_input[1823]), .B(n3887), .Z(n3889) );
  XOR U3772 ( .A(n3890), .B(n3891), .Z(n3887) );
  AND U3773 ( .A(n459), .B(n3892), .Z(n3891) );
  XNOR U3774 ( .A(p_input[1839]), .B(n3890), .Z(n3892) );
  XOR U3775 ( .A(n3893), .B(n3894), .Z(n3890) );
  AND U3776 ( .A(n463), .B(n3895), .Z(n3894) );
  XNOR U3777 ( .A(p_input[1855]), .B(n3893), .Z(n3895) );
  XOR U3778 ( .A(n3896), .B(n3897), .Z(n3893) );
  AND U3779 ( .A(n467), .B(n3898), .Z(n3897) );
  XNOR U3780 ( .A(p_input[1871]), .B(n3896), .Z(n3898) );
  XOR U3781 ( .A(n3899), .B(n3900), .Z(n3896) );
  AND U3782 ( .A(n471), .B(n3901), .Z(n3900) );
  XNOR U3783 ( .A(p_input[1887]), .B(n3899), .Z(n3901) );
  XOR U3784 ( .A(n3902), .B(n3903), .Z(n3899) );
  AND U3785 ( .A(n475), .B(n3904), .Z(n3903) );
  XNOR U3786 ( .A(p_input[1903]), .B(n3902), .Z(n3904) );
  XOR U3787 ( .A(n3905), .B(n3906), .Z(n3902) );
  AND U3788 ( .A(n479), .B(n3907), .Z(n3906) );
  XNOR U3789 ( .A(p_input[1919]), .B(n3905), .Z(n3907) );
  XOR U3790 ( .A(n3908), .B(n3909), .Z(n3905) );
  AND U3791 ( .A(n483), .B(n3910), .Z(n3909) );
  XNOR U3792 ( .A(p_input[1935]), .B(n3908), .Z(n3910) );
  XOR U3793 ( .A(n3911), .B(n3912), .Z(n3908) );
  AND U3794 ( .A(n487), .B(n3913), .Z(n3912) );
  XNOR U3795 ( .A(p_input[1951]), .B(n3911), .Z(n3913) );
  XOR U3796 ( .A(n3914), .B(n3915), .Z(n3911) );
  AND U3797 ( .A(n491), .B(n3916), .Z(n3915) );
  XNOR U3798 ( .A(p_input[1967]), .B(n3914), .Z(n3916) );
  XOR U3799 ( .A(n3917), .B(n3918), .Z(n3914) );
  AND U3800 ( .A(n495), .B(n3919), .Z(n3918) );
  XNOR U3801 ( .A(p_input[1983]), .B(n3917), .Z(n3919) );
  XOR U3802 ( .A(n3920), .B(n3921), .Z(n3917) );
  AND U3803 ( .A(n499), .B(n3922), .Z(n3921) );
  XNOR U3804 ( .A(p_input[1999]), .B(n3920), .Z(n3922) );
  XNOR U3805 ( .A(n3923), .B(n3924), .Z(n3920) );
  AND U3806 ( .A(n503), .B(n3925), .Z(n3924) );
  XOR U3807 ( .A(p_input[2015]), .B(n3923), .Z(n3925) );
  XOR U3808 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n3926), .Z(n3923) );
  AND U3809 ( .A(n506), .B(n3927), .Z(n3926) );
  XOR U3810 ( .A(p_input[2031]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n3927)
         );
  XNOR U3811 ( .A(n3928), .B(n3929), .Z(o[14]) );
  AND U3812 ( .A(n3), .B(n3930), .Z(n3928) );
  XNOR U3813 ( .A(p_input[14]), .B(n3929), .Z(n3930) );
  XOR U3814 ( .A(n3931), .B(n3932), .Z(n3929) );
  AND U3815 ( .A(n7), .B(n3933), .Z(n3932) );
  XNOR U3816 ( .A(p_input[30]), .B(n3931), .Z(n3933) );
  XOR U3817 ( .A(n3934), .B(n3935), .Z(n3931) );
  AND U3818 ( .A(n11), .B(n3936), .Z(n3935) );
  XNOR U3819 ( .A(p_input[46]), .B(n3934), .Z(n3936) );
  XOR U3820 ( .A(n3937), .B(n3938), .Z(n3934) );
  AND U3821 ( .A(n15), .B(n3939), .Z(n3938) );
  XNOR U3822 ( .A(p_input[62]), .B(n3937), .Z(n3939) );
  XOR U3823 ( .A(n3940), .B(n3941), .Z(n3937) );
  AND U3824 ( .A(n19), .B(n3942), .Z(n3941) );
  XNOR U3825 ( .A(p_input[78]), .B(n3940), .Z(n3942) );
  XOR U3826 ( .A(n3943), .B(n3944), .Z(n3940) );
  AND U3827 ( .A(n23), .B(n3945), .Z(n3944) );
  XNOR U3828 ( .A(p_input[94]), .B(n3943), .Z(n3945) );
  XOR U3829 ( .A(n3946), .B(n3947), .Z(n3943) );
  AND U3830 ( .A(n27), .B(n3948), .Z(n3947) );
  XNOR U3831 ( .A(p_input[110]), .B(n3946), .Z(n3948) );
  XOR U3832 ( .A(n3949), .B(n3950), .Z(n3946) );
  AND U3833 ( .A(n31), .B(n3951), .Z(n3950) );
  XNOR U3834 ( .A(p_input[126]), .B(n3949), .Z(n3951) );
  XOR U3835 ( .A(n3952), .B(n3953), .Z(n3949) );
  AND U3836 ( .A(n35), .B(n3954), .Z(n3953) );
  XNOR U3837 ( .A(p_input[142]), .B(n3952), .Z(n3954) );
  XOR U3838 ( .A(n3955), .B(n3956), .Z(n3952) );
  AND U3839 ( .A(n39), .B(n3957), .Z(n3956) );
  XNOR U3840 ( .A(p_input[158]), .B(n3955), .Z(n3957) );
  XOR U3841 ( .A(n3958), .B(n3959), .Z(n3955) );
  AND U3842 ( .A(n43), .B(n3960), .Z(n3959) );
  XNOR U3843 ( .A(p_input[174]), .B(n3958), .Z(n3960) );
  XOR U3844 ( .A(n3961), .B(n3962), .Z(n3958) );
  AND U3845 ( .A(n47), .B(n3963), .Z(n3962) );
  XNOR U3846 ( .A(p_input[190]), .B(n3961), .Z(n3963) );
  XOR U3847 ( .A(n3964), .B(n3965), .Z(n3961) );
  AND U3848 ( .A(n51), .B(n3966), .Z(n3965) );
  XNOR U3849 ( .A(p_input[206]), .B(n3964), .Z(n3966) );
  XOR U3850 ( .A(n3967), .B(n3968), .Z(n3964) );
  AND U3851 ( .A(n55), .B(n3969), .Z(n3968) );
  XNOR U3852 ( .A(p_input[222]), .B(n3967), .Z(n3969) );
  XOR U3853 ( .A(n3970), .B(n3971), .Z(n3967) );
  AND U3854 ( .A(n59), .B(n3972), .Z(n3971) );
  XNOR U3855 ( .A(p_input[238]), .B(n3970), .Z(n3972) );
  XOR U3856 ( .A(n3973), .B(n3974), .Z(n3970) );
  AND U3857 ( .A(n63), .B(n3975), .Z(n3974) );
  XNOR U3858 ( .A(p_input[254]), .B(n3973), .Z(n3975) );
  XOR U3859 ( .A(n3976), .B(n3977), .Z(n3973) );
  AND U3860 ( .A(n67), .B(n3978), .Z(n3977) );
  XNOR U3861 ( .A(p_input[270]), .B(n3976), .Z(n3978) );
  XOR U3862 ( .A(n3979), .B(n3980), .Z(n3976) );
  AND U3863 ( .A(n71), .B(n3981), .Z(n3980) );
  XNOR U3864 ( .A(p_input[286]), .B(n3979), .Z(n3981) );
  XOR U3865 ( .A(n3982), .B(n3983), .Z(n3979) );
  AND U3866 ( .A(n75), .B(n3984), .Z(n3983) );
  XNOR U3867 ( .A(p_input[302]), .B(n3982), .Z(n3984) );
  XOR U3868 ( .A(n3985), .B(n3986), .Z(n3982) );
  AND U3869 ( .A(n79), .B(n3987), .Z(n3986) );
  XNOR U3870 ( .A(p_input[318]), .B(n3985), .Z(n3987) );
  XOR U3871 ( .A(n3988), .B(n3989), .Z(n3985) );
  AND U3872 ( .A(n83), .B(n3990), .Z(n3989) );
  XNOR U3873 ( .A(p_input[334]), .B(n3988), .Z(n3990) );
  XOR U3874 ( .A(n3991), .B(n3992), .Z(n3988) );
  AND U3875 ( .A(n87), .B(n3993), .Z(n3992) );
  XNOR U3876 ( .A(p_input[350]), .B(n3991), .Z(n3993) );
  XOR U3877 ( .A(n3994), .B(n3995), .Z(n3991) );
  AND U3878 ( .A(n91), .B(n3996), .Z(n3995) );
  XNOR U3879 ( .A(p_input[366]), .B(n3994), .Z(n3996) );
  XOR U3880 ( .A(n3997), .B(n3998), .Z(n3994) );
  AND U3881 ( .A(n95), .B(n3999), .Z(n3998) );
  XNOR U3882 ( .A(p_input[382]), .B(n3997), .Z(n3999) );
  XOR U3883 ( .A(n4000), .B(n4001), .Z(n3997) );
  AND U3884 ( .A(n99), .B(n4002), .Z(n4001) );
  XNOR U3885 ( .A(p_input[398]), .B(n4000), .Z(n4002) );
  XOR U3886 ( .A(n4003), .B(n4004), .Z(n4000) );
  AND U3887 ( .A(n103), .B(n4005), .Z(n4004) );
  XNOR U3888 ( .A(p_input[414]), .B(n4003), .Z(n4005) );
  XOR U3889 ( .A(n4006), .B(n4007), .Z(n4003) );
  AND U3890 ( .A(n107), .B(n4008), .Z(n4007) );
  XNOR U3891 ( .A(p_input[430]), .B(n4006), .Z(n4008) );
  XOR U3892 ( .A(n4009), .B(n4010), .Z(n4006) );
  AND U3893 ( .A(n111), .B(n4011), .Z(n4010) );
  XNOR U3894 ( .A(p_input[446]), .B(n4009), .Z(n4011) );
  XOR U3895 ( .A(n4012), .B(n4013), .Z(n4009) );
  AND U3896 ( .A(n115), .B(n4014), .Z(n4013) );
  XNOR U3897 ( .A(p_input[462]), .B(n4012), .Z(n4014) );
  XOR U3898 ( .A(n4015), .B(n4016), .Z(n4012) );
  AND U3899 ( .A(n119), .B(n4017), .Z(n4016) );
  XNOR U3900 ( .A(p_input[478]), .B(n4015), .Z(n4017) );
  XOR U3901 ( .A(n4018), .B(n4019), .Z(n4015) );
  AND U3902 ( .A(n123), .B(n4020), .Z(n4019) );
  XNOR U3903 ( .A(p_input[494]), .B(n4018), .Z(n4020) );
  XOR U3904 ( .A(n4021), .B(n4022), .Z(n4018) );
  AND U3905 ( .A(n127), .B(n4023), .Z(n4022) );
  XNOR U3906 ( .A(p_input[510]), .B(n4021), .Z(n4023) );
  XOR U3907 ( .A(n4024), .B(n4025), .Z(n4021) );
  AND U3908 ( .A(n131), .B(n4026), .Z(n4025) );
  XNOR U3909 ( .A(p_input[526]), .B(n4024), .Z(n4026) );
  XOR U3910 ( .A(n4027), .B(n4028), .Z(n4024) );
  AND U3911 ( .A(n135), .B(n4029), .Z(n4028) );
  XNOR U3912 ( .A(p_input[542]), .B(n4027), .Z(n4029) );
  XOR U3913 ( .A(n4030), .B(n4031), .Z(n4027) );
  AND U3914 ( .A(n139), .B(n4032), .Z(n4031) );
  XNOR U3915 ( .A(p_input[558]), .B(n4030), .Z(n4032) );
  XOR U3916 ( .A(n4033), .B(n4034), .Z(n4030) );
  AND U3917 ( .A(n143), .B(n4035), .Z(n4034) );
  XNOR U3918 ( .A(p_input[574]), .B(n4033), .Z(n4035) );
  XOR U3919 ( .A(n4036), .B(n4037), .Z(n4033) );
  AND U3920 ( .A(n147), .B(n4038), .Z(n4037) );
  XNOR U3921 ( .A(p_input[590]), .B(n4036), .Z(n4038) );
  XOR U3922 ( .A(n4039), .B(n4040), .Z(n4036) );
  AND U3923 ( .A(n151), .B(n4041), .Z(n4040) );
  XNOR U3924 ( .A(p_input[606]), .B(n4039), .Z(n4041) );
  XOR U3925 ( .A(n4042), .B(n4043), .Z(n4039) );
  AND U3926 ( .A(n155), .B(n4044), .Z(n4043) );
  XNOR U3927 ( .A(p_input[622]), .B(n4042), .Z(n4044) );
  XOR U3928 ( .A(n4045), .B(n4046), .Z(n4042) );
  AND U3929 ( .A(n159), .B(n4047), .Z(n4046) );
  XNOR U3930 ( .A(p_input[638]), .B(n4045), .Z(n4047) );
  XOR U3931 ( .A(n4048), .B(n4049), .Z(n4045) );
  AND U3932 ( .A(n163), .B(n4050), .Z(n4049) );
  XNOR U3933 ( .A(p_input[654]), .B(n4048), .Z(n4050) );
  XOR U3934 ( .A(n4051), .B(n4052), .Z(n4048) );
  AND U3935 ( .A(n167), .B(n4053), .Z(n4052) );
  XNOR U3936 ( .A(p_input[670]), .B(n4051), .Z(n4053) );
  XOR U3937 ( .A(n4054), .B(n4055), .Z(n4051) );
  AND U3938 ( .A(n171), .B(n4056), .Z(n4055) );
  XNOR U3939 ( .A(p_input[686]), .B(n4054), .Z(n4056) );
  XOR U3940 ( .A(n4057), .B(n4058), .Z(n4054) );
  AND U3941 ( .A(n175), .B(n4059), .Z(n4058) );
  XNOR U3942 ( .A(p_input[702]), .B(n4057), .Z(n4059) );
  XOR U3943 ( .A(n4060), .B(n4061), .Z(n4057) );
  AND U3944 ( .A(n179), .B(n4062), .Z(n4061) );
  XNOR U3945 ( .A(p_input[718]), .B(n4060), .Z(n4062) );
  XOR U3946 ( .A(n4063), .B(n4064), .Z(n4060) );
  AND U3947 ( .A(n183), .B(n4065), .Z(n4064) );
  XNOR U3948 ( .A(p_input[734]), .B(n4063), .Z(n4065) );
  XOR U3949 ( .A(n4066), .B(n4067), .Z(n4063) );
  AND U3950 ( .A(n187), .B(n4068), .Z(n4067) );
  XNOR U3951 ( .A(p_input[750]), .B(n4066), .Z(n4068) );
  XOR U3952 ( .A(n4069), .B(n4070), .Z(n4066) );
  AND U3953 ( .A(n191), .B(n4071), .Z(n4070) );
  XNOR U3954 ( .A(p_input[766]), .B(n4069), .Z(n4071) );
  XOR U3955 ( .A(n4072), .B(n4073), .Z(n4069) );
  AND U3956 ( .A(n195), .B(n4074), .Z(n4073) );
  XNOR U3957 ( .A(p_input[782]), .B(n4072), .Z(n4074) );
  XOR U3958 ( .A(n4075), .B(n4076), .Z(n4072) );
  AND U3959 ( .A(n199), .B(n4077), .Z(n4076) );
  XNOR U3960 ( .A(p_input[798]), .B(n4075), .Z(n4077) );
  XOR U3961 ( .A(n4078), .B(n4079), .Z(n4075) );
  AND U3962 ( .A(n203), .B(n4080), .Z(n4079) );
  XNOR U3963 ( .A(p_input[814]), .B(n4078), .Z(n4080) );
  XOR U3964 ( .A(n4081), .B(n4082), .Z(n4078) );
  AND U3965 ( .A(n207), .B(n4083), .Z(n4082) );
  XNOR U3966 ( .A(p_input[830]), .B(n4081), .Z(n4083) );
  XOR U3967 ( .A(n4084), .B(n4085), .Z(n4081) );
  AND U3968 ( .A(n211), .B(n4086), .Z(n4085) );
  XNOR U3969 ( .A(p_input[846]), .B(n4084), .Z(n4086) );
  XOR U3970 ( .A(n4087), .B(n4088), .Z(n4084) );
  AND U3971 ( .A(n215), .B(n4089), .Z(n4088) );
  XNOR U3972 ( .A(p_input[862]), .B(n4087), .Z(n4089) );
  XOR U3973 ( .A(n4090), .B(n4091), .Z(n4087) );
  AND U3974 ( .A(n219), .B(n4092), .Z(n4091) );
  XNOR U3975 ( .A(p_input[878]), .B(n4090), .Z(n4092) );
  XOR U3976 ( .A(n4093), .B(n4094), .Z(n4090) );
  AND U3977 ( .A(n223), .B(n4095), .Z(n4094) );
  XNOR U3978 ( .A(p_input[894]), .B(n4093), .Z(n4095) );
  XOR U3979 ( .A(n4096), .B(n4097), .Z(n4093) );
  AND U3980 ( .A(n227), .B(n4098), .Z(n4097) );
  XNOR U3981 ( .A(p_input[910]), .B(n4096), .Z(n4098) );
  XOR U3982 ( .A(n4099), .B(n4100), .Z(n4096) );
  AND U3983 ( .A(n231), .B(n4101), .Z(n4100) );
  XNOR U3984 ( .A(p_input[926]), .B(n4099), .Z(n4101) );
  XOR U3985 ( .A(n4102), .B(n4103), .Z(n4099) );
  AND U3986 ( .A(n235), .B(n4104), .Z(n4103) );
  XNOR U3987 ( .A(p_input[942]), .B(n4102), .Z(n4104) );
  XOR U3988 ( .A(n4105), .B(n4106), .Z(n4102) );
  AND U3989 ( .A(n239), .B(n4107), .Z(n4106) );
  XNOR U3990 ( .A(p_input[958]), .B(n4105), .Z(n4107) );
  XOR U3991 ( .A(n4108), .B(n4109), .Z(n4105) );
  AND U3992 ( .A(n243), .B(n4110), .Z(n4109) );
  XNOR U3993 ( .A(p_input[974]), .B(n4108), .Z(n4110) );
  XOR U3994 ( .A(n4111), .B(n4112), .Z(n4108) );
  AND U3995 ( .A(n247), .B(n4113), .Z(n4112) );
  XNOR U3996 ( .A(p_input[990]), .B(n4111), .Z(n4113) );
  XOR U3997 ( .A(n4114), .B(n4115), .Z(n4111) );
  AND U3998 ( .A(n251), .B(n4116), .Z(n4115) );
  XNOR U3999 ( .A(p_input[1006]), .B(n4114), .Z(n4116) );
  XOR U4000 ( .A(n4117), .B(n4118), .Z(n4114) );
  AND U4001 ( .A(n255), .B(n4119), .Z(n4118) );
  XNOR U4002 ( .A(p_input[1022]), .B(n4117), .Z(n4119) );
  XOR U4003 ( .A(n4120), .B(n4121), .Z(n4117) );
  AND U4004 ( .A(n259), .B(n4122), .Z(n4121) );
  XNOR U4005 ( .A(p_input[1038]), .B(n4120), .Z(n4122) );
  XOR U4006 ( .A(n4123), .B(n4124), .Z(n4120) );
  AND U4007 ( .A(n263), .B(n4125), .Z(n4124) );
  XNOR U4008 ( .A(p_input[1054]), .B(n4123), .Z(n4125) );
  XOR U4009 ( .A(n4126), .B(n4127), .Z(n4123) );
  AND U4010 ( .A(n267), .B(n4128), .Z(n4127) );
  XNOR U4011 ( .A(p_input[1070]), .B(n4126), .Z(n4128) );
  XOR U4012 ( .A(n4129), .B(n4130), .Z(n4126) );
  AND U4013 ( .A(n271), .B(n4131), .Z(n4130) );
  XNOR U4014 ( .A(p_input[1086]), .B(n4129), .Z(n4131) );
  XOR U4015 ( .A(n4132), .B(n4133), .Z(n4129) );
  AND U4016 ( .A(n275), .B(n4134), .Z(n4133) );
  XNOR U4017 ( .A(p_input[1102]), .B(n4132), .Z(n4134) );
  XOR U4018 ( .A(n4135), .B(n4136), .Z(n4132) );
  AND U4019 ( .A(n279), .B(n4137), .Z(n4136) );
  XNOR U4020 ( .A(p_input[1118]), .B(n4135), .Z(n4137) );
  XOR U4021 ( .A(n4138), .B(n4139), .Z(n4135) );
  AND U4022 ( .A(n283), .B(n4140), .Z(n4139) );
  XNOR U4023 ( .A(p_input[1134]), .B(n4138), .Z(n4140) );
  XOR U4024 ( .A(n4141), .B(n4142), .Z(n4138) );
  AND U4025 ( .A(n287), .B(n4143), .Z(n4142) );
  XNOR U4026 ( .A(p_input[1150]), .B(n4141), .Z(n4143) );
  XOR U4027 ( .A(n4144), .B(n4145), .Z(n4141) );
  AND U4028 ( .A(n291), .B(n4146), .Z(n4145) );
  XNOR U4029 ( .A(p_input[1166]), .B(n4144), .Z(n4146) );
  XOR U4030 ( .A(n4147), .B(n4148), .Z(n4144) );
  AND U4031 ( .A(n295), .B(n4149), .Z(n4148) );
  XNOR U4032 ( .A(p_input[1182]), .B(n4147), .Z(n4149) );
  XOR U4033 ( .A(n4150), .B(n4151), .Z(n4147) );
  AND U4034 ( .A(n299), .B(n4152), .Z(n4151) );
  XNOR U4035 ( .A(p_input[1198]), .B(n4150), .Z(n4152) );
  XOR U4036 ( .A(n4153), .B(n4154), .Z(n4150) );
  AND U4037 ( .A(n303), .B(n4155), .Z(n4154) );
  XNOR U4038 ( .A(p_input[1214]), .B(n4153), .Z(n4155) );
  XOR U4039 ( .A(n4156), .B(n4157), .Z(n4153) );
  AND U4040 ( .A(n307), .B(n4158), .Z(n4157) );
  XNOR U4041 ( .A(p_input[1230]), .B(n4156), .Z(n4158) );
  XOR U4042 ( .A(n4159), .B(n4160), .Z(n4156) );
  AND U4043 ( .A(n311), .B(n4161), .Z(n4160) );
  XNOR U4044 ( .A(p_input[1246]), .B(n4159), .Z(n4161) );
  XOR U4045 ( .A(n4162), .B(n4163), .Z(n4159) );
  AND U4046 ( .A(n315), .B(n4164), .Z(n4163) );
  XNOR U4047 ( .A(p_input[1262]), .B(n4162), .Z(n4164) );
  XOR U4048 ( .A(n4165), .B(n4166), .Z(n4162) );
  AND U4049 ( .A(n319), .B(n4167), .Z(n4166) );
  XNOR U4050 ( .A(p_input[1278]), .B(n4165), .Z(n4167) );
  XOR U4051 ( .A(n4168), .B(n4169), .Z(n4165) );
  AND U4052 ( .A(n323), .B(n4170), .Z(n4169) );
  XNOR U4053 ( .A(p_input[1294]), .B(n4168), .Z(n4170) );
  XOR U4054 ( .A(n4171), .B(n4172), .Z(n4168) );
  AND U4055 ( .A(n327), .B(n4173), .Z(n4172) );
  XNOR U4056 ( .A(p_input[1310]), .B(n4171), .Z(n4173) );
  XOR U4057 ( .A(n4174), .B(n4175), .Z(n4171) );
  AND U4058 ( .A(n331), .B(n4176), .Z(n4175) );
  XNOR U4059 ( .A(p_input[1326]), .B(n4174), .Z(n4176) );
  XOR U4060 ( .A(n4177), .B(n4178), .Z(n4174) );
  AND U4061 ( .A(n335), .B(n4179), .Z(n4178) );
  XNOR U4062 ( .A(p_input[1342]), .B(n4177), .Z(n4179) );
  XOR U4063 ( .A(n4180), .B(n4181), .Z(n4177) );
  AND U4064 ( .A(n339), .B(n4182), .Z(n4181) );
  XNOR U4065 ( .A(p_input[1358]), .B(n4180), .Z(n4182) );
  XOR U4066 ( .A(n4183), .B(n4184), .Z(n4180) );
  AND U4067 ( .A(n343), .B(n4185), .Z(n4184) );
  XNOR U4068 ( .A(p_input[1374]), .B(n4183), .Z(n4185) );
  XOR U4069 ( .A(n4186), .B(n4187), .Z(n4183) );
  AND U4070 ( .A(n347), .B(n4188), .Z(n4187) );
  XNOR U4071 ( .A(p_input[1390]), .B(n4186), .Z(n4188) );
  XOR U4072 ( .A(n4189), .B(n4190), .Z(n4186) );
  AND U4073 ( .A(n351), .B(n4191), .Z(n4190) );
  XNOR U4074 ( .A(p_input[1406]), .B(n4189), .Z(n4191) );
  XOR U4075 ( .A(n4192), .B(n4193), .Z(n4189) );
  AND U4076 ( .A(n355), .B(n4194), .Z(n4193) );
  XNOR U4077 ( .A(p_input[1422]), .B(n4192), .Z(n4194) );
  XOR U4078 ( .A(n4195), .B(n4196), .Z(n4192) );
  AND U4079 ( .A(n359), .B(n4197), .Z(n4196) );
  XNOR U4080 ( .A(p_input[1438]), .B(n4195), .Z(n4197) );
  XOR U4081 ( .A(n4198), .B(n4199), .Z(n4195) );
  AND U4082 ( .A(n363), .B(n4200), .Z(n4199) );
  XNOR U4083 ( .A(p_input[1454]), .B(n4198), .Z(n4200) );
  XOR U4084 ( .A(n4201), .B(n4202), .Z(n4198) );
  AND U4085 ( .A(n367), .B(n4203), .Z(n4202) );
  XNOR U4086 ( .A(p_input[1470]), .B(n4201), .Z(n4203) );
  XOR U4087 ( .A(n4204), .B(n4205), .Z(n4201) );
  AND U4088 ( .A(n371), .B(n4206), .Z(n4205) );
  XNOR U4089 ( .A(p_input[1486]), .B(n4204), .Z(n4206) );
  XOR U4090 ( .A(n4207), .B(n4208), .Z(n4204) );
  AND U4091 ( .A(n375), .B(n4209), .Z(n4208) );
  XNOR U4092 ( .A(p_input[1502]), .B(n4207), .Z(n4209) );
  XOR U4093 ( .A(n4210), .B(n4211), .Z(n4207) );
  AND U4094 ( .A(n379), .B(n4212), .Z(n4211) );
  XNOR U4095 ( .A(p_input[1518]), .B(n4210), .Z(n4212) );
  XOR U4096 ( .A(n4213), .B(n4214), .Z(n4210) );
  AND U4097 ( .A(n383), .B(n4215), .Z(n4214) );
  XNOR U4098 ( .A(p_input[1534]), .B(n4213), .Z(n4215) );
  XOR U4099 ( .A(n4216), .B(n4217), .Z(n4213) );
  AND U4100 ( .A(n387), .B(n4218), .Z(n4217) );
  XNOR U4101 ( .A(p_input[1550]), .B(n4216), .Z(n4218) );
  XOR U4102 ( .A(n4219), .B(n4220), .Z(n4216) );
  AND U4103 ( .A(n391), .B(n4221), .Z(n4220) );
  XNOR U4104 ( .A(p_input[1566]), .B(n4219), .Z(n4221) );
  XOR U4105 ( .A(n4222), .B(n4223), .Z(n4219) );
  AND U4106 ( .A(n395), .B(n4224), .Z(n4223) );
  XNOR U4107 ( .A(p_input[1582]), .B(n4222), .Z(n4224) );
  XOR U4108 ( .A(n4225), .B(n4226), .Z(n4222) );
  AND U4109 ( .A(n399), .B(n4227), .Z(n4226) );
  XNOR U4110 ( .A(p_input[1598]), .B(n4225), .Z(n4227) );
  XOR U4111 ( .A(n4228), .B(n4229), .Z(n4225) );
  AND U4112 ( .A(n403), .B(n4230), .Z(n4229) );
  XNOR U4113 ( .A(p_input[1614]), .B(n4228), .Z(n4230) );
  XOR U4114 ( .A(n4231), .B(n4232), .Z(n4228) );
  AND U4115 ( .A(n407), .B(n4233), .Z(n4232) );
  XNOR U4116 ( .A(p_input[1630]), .B(n4231), .Z(n4233) );
  XOR U4117 ( .A(n4234), .B(n4235), .Z(n4231) );
  AND U4118 ( .A(n411), .B(n4236), .Z(n4235) );
  XNOR U4119 ( .A(p_input[1646]), .B(n4234), .Z(n4236) );
  XOR U4120 ( .A(n4237), .B(n4238), .Z(n4234) );
  AND U4121 ( .A(n415), .B(n4239), .Z(n4238) );
  XNOR U4122 ( .A(p_input[1662]), .B(n4237), .Z(n4239) );
  XOR U4123 ( .A(n4240), .B(n4241), .Z(n4237) );
  AND U4124 ( .A(n419), .B(n4242), .Z(n4241) );
  XNOR U4125 ( .A(p_input[1678]), .B(n4240), .Z(n4242) );
  XOR U4126 ( .A(n4243), .B(n4244), .Z(n4240) );
  AND U4127 ( .A(n423), .B(n4245), .Z(n4244) );
  XNOR U4128 ( .A(p_input[1694]), .B(n4243), .Z(n4245) );
  XOR U4129 ( .A(n4246), .B(n4247), .Z(n4243) );
  AND U4130 ( .A(n427), .B(n4248), .Z(n4247) );
  XNOR U4131 ( .A(p_input[1710]), .B(n4246), .Z(n4248) );
  XOR U4132 ( .A(n4249), .B(n4250), .Z(n4246) );
  AND U4133 ( .A(n431), .B(n4251), .Z(n4250) );
  XNOR U4134 ( .A(p_input[1726]), .B(n4249), .Z(n4251) );
  XOR U4135 ( .A(n4252), .B(n4253), .Z(n4249) );
  AND U4136 ( .A(n435), .B(n4254), .Z(n4253) );
  XNOR U4137 ( .A(p_input[1742]), .B(n4252), .Z(n4254) );
  XOR U4138 ( .A(n4255), .B(n4256), .Z(n4252) );
  AND U4139 ( .A(n439), .B(n4257), .Z(n4256) );
  XNOR U4140 ( .A(p_input[1758]), .B(n4255), .Z(n4257) );
  XOR U4141 ( .A(n4258), .B(n4259), .Z(n4255) );
  AND U4142 ( .A(n443), .B(n4260), .Z(n4259) );
  XNOR U4143 ( .A(p_input[1774]), .B(n4258), .Z(n4260) );
  XOR U4144 ( .A(n4261), .B(n4262), .Z(n4258) );
  AND U4145 ( .A(n447), .B(n4263), .Z(n4262) );
  XNOR U4146 ( .A(p_input[1790]), .B(n4261), .Z(n4263) );
  XOR U4147 ( .A(n4264), .B(n4265), .Z(n4261) );
  AND U4148 ( .A(n451), .B(n4266), .Z(n4265) );
  XNOR U4149 ( .A(p_input[1806]), .B(n4264), .Z(n4266) );
  XOR U4150 ( .A(n4267), .B(n4268), .Z(n4264) );
  AND U4151 ( .A(n455), .B(n4269), .Z(n4268) );
  XNOR U4152 ( .A(p_input[1822]), .B(n4267), .Z(n4269) );
  XOR U4153 ( .A(n4270), .B(n4271), .Z(n4267) );
  AND U4154 ( .A(n459), .B(n4272), .Z(n4271) );
  XNOR U4155 ( .A(p_input[1838]), .B(n4270), .Z(n4272) );
  XOR U4156 ( .A(n4273), .B(n4274), .Z(n4270) );
  AND U4157 ( .A(n463), .B(n4275), .Z(n4274) );
  XNOR U4158 ( .A(p_input[1854]), .B(n4273), .Z(n4275) );
  XOR U4159 ( .A(n4276), .B(n4277), .Z(n4273) );
  AND U4160 ( .A(n467), .B(n4278), .Z(n4277) );
  XNOR U4161 ( .A(p_input[1870]), .B(n4276), .Z(n4278) );
  XOR U4162 ( .A(n4279), .B(n4280), .Z(n4276) );
  AND U4163 ( .A(n471), .B(n4281), .Z(n4280) );
  XNOR U4164 ( .A(p_input[1886]), .B(n4279), .Z(n4281) );
  XOR U4165 ( .A(n4282), .B(n4283), .Z(n4279) );
  AND U4166 ( .A(n475), .B(n4284), .Z(n4283) );
  XNOR U4167 ( .A(p_input[1902]), .B(n4282), .Z(n4284) );
  XOR U4168 ( .A(n4285), .B(n4286), .Z(n4282) );
  AND U4169 ( .A(n479), .B(n4287), .Z(n4286) );
  XNOR U4170 ( .A(p_input[1918]), .B(n4285), .Z(n4287) );
  XOR U4171 ( .A(n4288), .B(n4289), .Z(n4285) );
  AND U4172 ( .A(n483), .B(n4290), .Z(n4289) );
  XNOR U4173 ( .A(p_input[1934]), .B(n4288), .Z(n4290) );
  XOR U4174 ( .A(n4291), .B(n4292), .Z(n4288) );
  AND U4175 ( .A(n487), .B(n4293), .Z(n4292) );
  XNOR U4176 ( .A(p_input[1950]), .B(n4291), .Z(n4293) );
  XOR U4177 ( .A(n4294), .B(n4295), .Z(n4291) );
  AND U4178 ( .A(n491), .B(n4296), .Z(n4295) );
  XNOR U4179 ( .A(p_input[1966]), .B(n4294), .Z(n4296) );
  XOR U4180 ( .A(n4297), .B(n4298), .Z(n4294) );
  AND U4181 ( .A(n495), .B(n4299), .Z(n4298) );
  XNOR U4182 ( .A(p_input[1982]), .B(n4297), .Z(n4299) );
  XOR U4183 ( .A(n4300), .B(n4301), .Z(n4297) );
  AND U4184 ( .A(n499), .B(n4302), .Z(n4301) );
  XNOR U4185 ( .A(p_input[1998]), .B(n4300), .Z(n4302) );
  XNOR U4186 ( .A(n4303), .B(n4304), .Z(n4300) );
  AND U4187 ( .A(n503), .B(n4305), .Z(n4304) );
  XOR U4188 ( .A(p_input[2014]), .B(n4303), .Z(n4305) );
  XOR U4189 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n4306), .Z(n4303) );
  AND U4190 ( .A(n506), .B(n4307), .Z(n4306) );
  XOR U4191 ( .A(p_input[2030]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n4307)
         );
  XNOR U4192 ( .A(n4308), .B(n4309), .Z(o[13]) );
  AND U4193 ( .A(n3), .B(n4310), .Z(n4308) );
  XNOR U4194 ( .A(p_input[13]), .B(n4309), .Z(n4310) );
  XOR U4195 ( .A(n4311), .B(n4312), .Z(n4309) );
  AND U4196 ( .A(n7), .B(n4313), .Z(n4312) );
  XNOR U4197 ( .A(p_input[29]), .B(n4311), .Z(n4313) );
  XOR U4198 ( .A(n4314), .B(n4315), .Z(n4311) );
  AND U4199 ( .A(n11), .B(n4316), .Z(n4315) );
  XNOR U4200 ( .A(p_input[45]), .B(n4314), .Z(n4316) );
  XOR U4201 ( .A(n4317), .B(n4318), .Z(n4314) );
  AND U4202 ( .A(n15), .B(n4319), .Z(n4318) );
  XNOR U4203 ( .A(p_input[61]), .B(n4317), .Z(n4319) );
  XOR U4204 ( .A(n4320), .B(n4321), .Z(n4317) );
  AND U4205 ( .A(n19), .B(n4322), .Z(n4321) );
  XNOR U4206 ( .A(p_input[77]), .B(n4320), .Z(n4322) );
  XOR U4207 ( .A(n4323), .B(n4324), .Z(n4320) );
  AND U4208 ( .A(n23), .B(n4325), .Z(n4324) );
  XNOR U4209 ( .A(p_input[93]), .B(n4323), .Z(n4325) );
  XOR U4210 ( .A(n4326), .B(n4327), .Z(n4323) );
  AND U4211 ( .A(n27), .B(n4328), .Z(n4327) );
  XNOR U4212 ( .A(p_input[109]), .B(n4326), .Z(n4328) );
  XOR U4213 ( .A(n4329), .B(n4330), .Z(n4326) );
  AND U4214 ( .A(n31), .B(n4331), .Z(n4330) );
  XNOR U4215 ( .A(p_input[125]), .B(n4329), .Z(n4331) );
  XOR U4216 ( .A(n4332), .B(n4333), .Z(n4329) );
  AND U4217 ( .A(n35), .B(n4334), .Z(n4333) );
  XNOR U4218 ( .A(p_input[141]), .B(n4332), .Z(n4334) );
  XOR U4219 ( .A(n4335), .B(n4336), .Z(n4332) );
  AND U4220 ( .A(n39), .B(n4337), .Z(n4336) );
  XNOR U4221 ( .A(p_input[157]), .B(n4335), .Z(n4337) );
  XOR U4222 ( .A(n4338), .B(n4339), .Z(n4335) );
  AND U4223 ( .A(n43), .B(n4340), .Z(n4339) );
  XNOR U4224 ( .A(p_input[173]), .B(n4338), .Z(n4340) );
  XOR U4225 ( .A(n4341), .B(n4342), .Z(n4338) );
  AND U4226 ( .A(n47), .B(n4343), .Z(n4342) );
  XNOR U4227 ( .A(p_input[189]), .B(n4341), .Z(n4343) );
  XOR U4228 ( .A(n4344), .B(n4345), .Z(n4341) );
  AND U4229 ( .A(n51), .B(n4346), .Z(n4345) );
  XNOR U4230 ( .A(p_input[205]), .B(n4344), .Z(n4346) );
  XOR U4231 ( .A(n4347), .B(n4348), .Z(n4344) );
  AND U4232 ( .A(n55), .B(n4349), .Z(n4348) );
  XNOR U4233 ( .A(p_input[221]), .B(n4347), .Z(n4349) );
  XOR U4234 ( .A(n4350), .B(n4351), .Z(n4347) );
  AND U4235 ( .A(n59), .B(n4352), .Z(n4351) );
  XNOR U4236 ( .A(p_input[237]), .B(n4350), .Z(n4352) );
  XOR U4237 ( .A(n4353), .B(n4354), .Z(n4350) );
  AND U4238 ( .A(n63), .B(n4355), .Z(n4354) );
  XNOR U4239 ( .A(p_input[253]), .B(n4353), .Z(n4355) );
  XOR U4240 ( .A(n4356), .B(n4357), .Z(n4353) );
  AND U4241 ( .A(n67), .B(n4358), .Z(n4357) );
  XNOR U4242 ( .A(p_input[269]), .B(n4356), .Z(n4358) );
  XOR U4243 ( .A(n4359), .B(n4360), .Z(n4356) );
  AND U4244 ( .A(n71), .B(n4361), .Z(n4360) );
  XNOR U4245 ( .A(p_input[285]), .B(n4359), .Z(n4361) );
  XOR U4246 ( .A(n4362), .B(n4363), .Z(n4359) );
  AND U4247 ( .A(n75), .B(n4364), .Z(n4363) );
  XNOR U4248 ( .A(p_input[301]), .B(n4362), .Z(n4364) );
  XOR U4249 ( .A(n4365), .B(n4366), .Z(n4362) );
  AND U4250 ( .A(n79), .B(n4367), .Z(n4366) );
  XNOR U4251 ( .A(p_input[317]), .B(n4365), .Z(n4367) );
  XOR U4252 ( .A(n4368), .B(n4369), .Z(n4365) );
  AND U4253 ( .A(n83), .B(n4370), .Z(n4369) );
  XNOR U4254 ( .A(p_input[333]), .B(n4368), .Z(n4370) );
  XOR U4255 ( .A(n4371), .B(n4372), .Z(n4368) );
  AND U4256 ( .A(n87), .B(n4373), .Z(n4372) );
  XNOR U4257 ( .A(p_input[349]), .B(n4371), .Z(n4373) );
  XOR U4258 ( .A(n4374), .B(n4375), .Z(n4371) );
  AND U4259 ( .A(n91), .B(n4376), .Z(n4375) );
  XNOR U4260 ( .A(p_input[365]), .B(n4374), .Z(n4376) );
  XOR U4261 ( .A(n4377), .B(n4378), .Z(n4374) );
  AND U4262 ( .A(n95), .B(n4379), .Z(n4378) );
  XNOR U4263 ( .A(p_input[381]), .B(n4377), .Z(n4379) );
  XOR U4264 ( .A(n4380), .B(n4381), .Z(n4377) );
  AND U4265 ( .A(n99), .B(n4382), .Z(n4381) );
  XNOR U4266 ( .A(p_input[397]), .B(n4380), .Z(n4382) );
  XOR U4267 ( .A(n4383), .B(n4384), .Z(n4380) );
  AND U4268 ( .A(n103), .B(n4385), .Z(n4384) );
  XNOR U4269 ( .A(p_input[413]), .B(n4383), .Z(n4385) );
  XOR U4270 ( .A(n4386), .B(n4387), .Z(n4383) );
  AND U4271 ( .A(n107), .B(n4388), .Z(n4387) );
  XNOR U4272 ( .A(p_input[429]), .B(n4386), .Z(n4388) );
  XOR U4273 ( .A(n4389), .B(n4390), .Z(n4386) );
  AND U4274 ( .A(n111), .B(n4391), .Z(n4390) );
  XNOR U4275 ( .A(p_input[445]), .B(n4389), .Z(n4391) );
  XOR U4276 ( .A(n4392), .B(n4393), .Z(n4389) );
  AND U4277 ( .A(n115), .B(n4394), .Z(n4393) );
  XNOR U4278 ( .A(p_input[461]), .B(n4392), .Z(n4394) );
  XOR U4279 ( .A(n4395), .B(n4396), .Z(n4392) );
  AND U4280 ( .A(n119), .B(n4397), .Z(n4396) );
  XNOR U4281 ( .A(p_input[477]), .B(n4395), .Z(n4397) );
  XOR U4282 ( .A(n4398), .B(n4399), .Z(n4395) );
  AND U4283 ( .A(n123), .B(n4400), .Z(n4399) );
  XNOR U4284 ( .A(p_input[493]), .B(n4398), .Z(n4400) );
  XOR U4285 ( .A(n4401), .B(n4402), .Z(n4398) );
  AND U4286 ( .A(n127), .B(n4403), .Z(n4402) );
  XNOR U4287 ( .A(p_input[509]), .B(n4401), .Z(n4403) );
  XOR U4288 ( .A(n4404), .B(n4405), .Z(n4401) );
  AND U4289 ( .A(n131), .B(n4406), .Z(n4405) );
  XNOR U4290 ( .A(p_input[525]), .B(n4404), .Z(n4406) );
  XOR U4291 ( .A(n4407), .B(n4408), .Z(n4404) );
  AND U4292 ( .A(n135), .B(n4409), .Z(n4408) );
  XNOR U4293 ( .A(p_input[541]), .B(n4407), .Z(n4409) );
  XOR U4294 ( .A(n4410), .B(n4411), .Z(n4407) );
  AND U4295 ( .A(n139), .B(n4412), .Z(n4411) );
  XNOR U4296 ( .A(p_input[557]), .B(n4410), .Z(n4412) );
  XOR U4297 ( .A(n4413), .B(n4414), .Z(n4410) );
  AND U4298 ( .A(n143), .B(n4415), .Z(n4414) );
  XNOR U4299 ( .A(p_input[573]), .B(n4413), .Z(n4415) );
  XOR U4300 ( .A(n4416), .B(n4417), .Z(n4413) );
  AND U4301 ( .A(n147), .B(n4418), .Z(n4417) );
  XNOR U4302 ( .A(p_input[589]), .B(n4416), .Z(n4418) );
  XOR U4303 ( .A(n4419), .B(n4420), .Z(n4416) );
  AND U4304 ( .A(n151), .B(n4421), .Z(n4420) );
  XNOR U4305 ( .A(p_input[605]), .B(n4419), .Z(n4421) );
  XOR U4306 ( .A(n4422), .B(n4423), .Z(n4419) );
  AND U4307 ( .A(n155), .B(n4424), .Z(n4423) );
  XNOR U4308 ( .A(p_input[621]), .B(n4422), .Z(n4424) );
  XOR U4309 ( .A(n4425), .B(n4426), .Z(n4422) );
  AND U4310 ( .A(n159), .B(n4427), .Z(n4426) );
  XNOR U4311 ( .A(p_input[637]), .B(n4425), .Z(n4427) );
  XOR U4312 ( .A(n4428), .B(n4429), .Z(n4425) );
  AND U4313 ( .A(n163), .B(n4430), .Z(n4429) );
  XNOR U4314 ( .A(p_input[653]), .B(n4428), .Z(n4430) );
  XOR U4315 ( .A(n4431), .B(n4432), .Z(n4428) );
  AND U4316 ( .A(n167), .B(n4433), .Z(n4432) );
  XNOR U4317 ( .A(p_input[669]), .B(n4431), .Z(n4433) );
  XOR U4318 ( .A(n4434), .B(n4435), .Z(n4431) );
  AND U4319 ( .A(n171), .B(n4436), .Z(n4435) );
  XNOR U4320 ( .A(p_input[685]), .B(n4434), .Z(n4436) );
  XOR U4321 ( .A(n4437), .B(n4438), .Z(n4434) );
  AND U4322 ( .A(n175), .B(n4439), .Z(n4438) );
  XNOR U4323 ( .A(p_input[701]), .B(n4437), .Z(n4439) );
  XOR U4324 ( .A(n4440), .B(n4441), .Z(n4437) );
  AND U4325 ( .A(n179), .B(n4442), .Z(n4441) );
  XNOR U4326 ( .A(p_input[717]), .B(n4440), .Z(n4442) );
  XOR U4327 ( .A(n4443), .B(n4444), .Z(n4440) );
  AND U4328 ( .A(n183), .B(n4445), .Z(n4444) );
  XNOR U4329 ( .A(p_input[733]), .B(n4443), .Z(n4445) );
  XOR U4330 ( .A(n4446), .B(n4447), .Z(n4443) );
  AND U4331 ( .A(n187), .B(n4448), .Z(n4447) );
  XNOR U4332 ( .A(p_input[749]), .B(n4446), .Z(n4448) );
  XOR U4333 ( .A(n4449), .B(n4450), .Z(n4446) );
  AND U4334 ( .A(n191), .B(n4451), .Z(n4450) );
  XNOR U4335 ( .A(p_input[765]), .B(n4449), .Z(n4451) );
  XOR U4336 ( .A(n4452), .B(n4453), .Z(n4449) );
  AND U4337 ( .A(n195), .B(n4454), .Z(n4453) );
  XNOR U4338 ( .A(p_input[781]), .B(n4452), .Z(n4454) );
  XOR U4339 ( .A(n4455), .B(n4456), .Z(n4452) );
  AND U4340 ( .A(n199), .B(n4457), .Z(n4456) );
  XNOR U4341 ( .A(p_input[797]), .B(n4455), .Z(n4457) );
  XOR U4342 ( .A(n4458), .B(n4459), .Z(n4455) );
  AND U4343 ( .A(n203), .B(n4460), .Z(n4459) );
  XNOR U4344 ( .A(p_input[813]), .B(n4458), .Z(n4460) );
  XOR U4345 ( .A(n4461), .B(n4462), .Z(n4458) );
  AND U4346 ( .A(n207), .B(n4463), .Z(n4462) );
  XNOR U4347 ( .A(p_input[829]), .B(n4461), .Z(n4463) );
  XOR U4348 ( .A(n4464), .B(n4465), .Z(n4461) );
  AND U4349 ( .A(n211), .B(n4466), .Z(n4465) );
  XNOR U4350 ( .A(p_input[845]), .B(n4464), .Z(n4466) );
  XOR U4351 ( .A(n4467), .B(n4468), .Z(n4464) );
  AND U4352 ( .A(n215), .B(n4469), .Z(n4468) );
  XNOR U4353 ( .A(p_input[861]), .B(n4467), .Z(n4469) );
  XOR U4354 ( .A(n4470), .B(n4471), .Z(n4467) );
  AND U4355 ( .A(n219), .B(n4472), .Z(n4471) );
  XNOR U4356 ( .A(p_input[877]), .B(n4470), .Z(n4472) );
  XOR U4357 ( .A(n4473), .B(n4474), .Z(n4470) );
  AND U4358 ( .A(n223), .B(n4475), .Z(n4474) );
  XNOR U4359 ( .A(p_input[893]), .B(n4473), .Z(n4475) );
  XOR U4360 ( .A(n4476), .B(n4477), .Z(n4473) );
  AND U4361 ( .A(n227), .B(n4478), .Z(n4477) );
  XNOR U4362 ( .A(p_input[909]), .B(n4476), .Z(n4478) );
  XOR U4363 ( .A(n4479), .B(n4480), .Z(n4476) );
  AND U4364 ( .A(n231), .B(n4481), .Z(n4480) );
  XNOR U4365 ( .A(p_input[925]), .B(n4479), .Z(n4481) );
  XOR U4366 ( .A(n4482), .B(n4483), .Z(n4479) );
  AND U4367 ( .A(n235), .B(n4484), .Z(n4483) );
  XNOR U4368 ( .A(p_input[941]), .B(n4482), .Z(n4484) );
  XOR U4369 ( .A(n4485), .B(n4486), .Z(n4482) );
  AND U4370 ( .A(n239), .B(n4487), .Z(n4486) );
  XNOR U4371 ( .A(p_input[957]), .B(n4485), .Z(n4487) );
  XOR U4372 ( .A(n4488), .B(n4489), .Z(n4485) );
  AND U4373 ( .A(n243), .B(n4490), .Z(n4489) );
  XNOR U4374 ( .A(p_input[973]), .B(n4488), .Z(n4490) );
  XOR U4375 ( .A(n4491), .B(n4492), .Z(n4488) );
  AND U4376 ( .A(n247), .B(n4493), .Z(n4492) );
  XNOR U4377 ( .A(p_input[989]), .B(n4491), .Z(n4493) );
  XOR U4378 ( .A(n4494), .B(n4495), .Z(n4491) );
  AND U4379 ( .A(n251), .B(n4496), .Z(n4495) );
  XNOR U4380 ( .A(p_input[1005]), .B(n4494), .Z(n4496) );
  XOR U4381 ( .A(n4497), .B(n4498), .Z(n4494) );
  AND U4382 ( .A(n255), .B(n4499), .Z(n4498) );
  XNOR U4383 ( .A(p_input[1021]), .B(n4497), .Z(n4499) );
  XOR U4384 ( .A(n4500), .B(n4501), .Z(n4497) );
  AND U4385 ( .A(n259), .B(n4502), .Z(n4501) );
  XNOR U4386 ( .A(p_input[1037]), .B(n4500), .Z(n4502) );
  XOR U4387 ( .A(n4503), .B(n4504), .Z(n4500) );
  AND U4388 ( .A(n263), .B(n4505), .Z(n4504) );
  XNOR U4389 ( .A(p_input[1053]), .B(n4503), .Z(n4505) );
  XOR U4390 ( .A(n4506), .B(n4507), .Z(n4503) );
  AND U4391 ( .A(n267), .B(n4508), .Z(n4507) );
  XNOR U4392 ( .A(p_input[1069]), .B(n4506), .Z(n4508) );
  XOR U4393 ( .A(n4509), .B(n4510), .Z(n4506) );
  AND U4394 ( .A(n271), .B(n4511), .Z(n4510) );
  XNOR U4395 ( .A(p_input[1085]), .B(n4509), .Z(n4511) );
  XOR U4396 ( .A(n4512), .B(n4513), .Z(n4509) );
  AND U4397 ( .A(n275), .B(n4514), .Z(n4513) );
  XNOR U4398 ( .A(p_input[1101]), .B(n4512), .Z(n4514) );
  XOR U4399 ( .A(n4515), .B(n4516), .Z(n4512) );
  AND U4400 ( .A(n279), .B(n4517), .Z(n4516) );
  XNOR U4401 ( .A(p_input[1117]), .B(n4515), .Z(n4517) );
  XOR U4402 ( .A(n4518), .B(n4519), .Z(n4515) );
  AND U4403 ( .A(n283), .B(n4520), .Z(n4519) );
  XNOR U4404 ( .A(p_input[1133]), .B(n4518), .Z(n4520) );
  XOR U4405 ( .A(n4521), .B(n4522), .Z(n4518) );
  AND U4406 ( .A(n287), .B(n4523), .Z(n4522) );
  XNOR U4407 ( .A(p_input[1149]), .B(n4521), .Z(n4523) );
  XOR U4408 ( .A(n4524), .B(n4525), .Z(n4521) );
  AND U4409 ( .A(n291), .B(n4526), .Z(n4525) );
  XNOR U4410 ( .A(p_input[1165]), .B(n4524), .Z(n4526) );
  XOR U4411 ( .A(n4527), .B(n4528), .Z(n4524) );
  AND U4412 ( .A(n295), .B(n4529), .Z(n4528) );
  XNOR U4413 ( .A(p_input[1181]), .B(n4527), .Z(n4529) );
  XOR U4414 ( .A(n4530), .B(n4531), .Z(n4527) );
  AND U4415 ( .A(n299), .B(n4532), .Z(n4531) );
  XNOR U4416 ( .A(p_input[1197]), .B(n4530), .Z(n4532) );
  XOR U4417 ( .A(n4533), .B(n4534), .Z(n4530) );
  AND U4418 ( .A(n303), .B(n4535), .Z(n4534) );
  XNOR U4419 ( .A(p_input[1213]), .B(n4533), .Z(n4535) );
  XOR U4420 ( .A(n4536), .B(n4537), .Z(n4533) );
  AND U4421 ( .A(n307), .B(n4538), .Z(n4537) );
  XNOR U4422 ( .A(p_input[1229]), .B(n4536), .Z(n4538) );
  XOR U4423 ( .A(n4539), .B(n4540), .Z(n4536) );
  AND U4424 ( .A(n311), .B(n4541), .Z(n4540) );
  XNOR U4425 ( .A(p_input[1245]), .B(n4539), .Z(n4541) );
  XOR U4426 ( .A(n4542), .B(n4543), .Z(n4539) );
  AND U4427 ( .A(n315), .B(n4544), .Z(n4543) );
  XNOR U4428 ( .A(p_input[1261]), .B(n4542), .Z(n4544) );
  XOR U4429 ( .A(n4545), .B(n4546), .Z(n4542) );
  AND U4430 ( .A(n319), .B(n4547), .Z(n4546) );
  XNOR U4431 ( .A(p_input[1277]), .B(n4545), .Z(n4547) );
  XOR U4432 ( .A(n4548), .B(n4549), .Z(n4545) );
  AND U4433 ( .A(n323), .B(n4550), .Z(n4549) );
  XNOR U4434 ( .A(p_input[1293]), .B(n4548), .Z(n4550) );
  XOR U4435 ( .A(n4551), .B(n4552), .Z(n4548) );
  AND U4436 ( .A(n327), .B(n4553), .Z(n4552) );
  XNOR U4437 ( .A(p_input[1309]), .B(n4551), .Z(n4553) );
  XOR U4438 ( .A(n4554), .B(n4555), .Z(n4551) );
  AND U4439 ( .A(n331), .B(n4556), .Z(n4555) );
  XNOR U4440 ( .A(p_input[1325]), .B(n4554), .Z(n4556) );
  XOR U4441 ( .A(n4557), .B(n4558), .Z(n4554) );
  AND U4442 ( .A(n335), .B(n4559), .Z(n4558) );
  XNOR U4443 ( .A(p_input[1341]), .B(n4557), .Z(n4559) );
  XOR U4444 ( .A(n4560), .B(n4561), .Z(n4557) );
  AND U4445 ( .A(n339), .B(n4562), .Z(n4561) );
  XNOR U4446 ( .A(p_input[1357]), .B(n4560), .Z(n4562) );
  XOR U4447 ( .A(n4563), .B(n4564), .Z(n4560) );
  AND U4448 ( .A(n343), .B(n4565), .Z(n4564) );
  XNOR U4449 ( .A(p_input[1373]), .B(n4563), .Z(n4565) );
  XOR U4450 ( .A(n4566), .B(n4567), .Z(n4563) );
  AND U4451 ( .A(n347), .B(n4568), .Z(n4567) );
  XNOR U4452 ( .A(p_input[1389]), .B(n4566), .Z(n4568) );
  XOR U4453 ( .A(n4569), .B(n4570), .Z(n4566) );
  AND U4454 ( .A(n351), .B(n4571), .Z(n4570) );
  XNOR U4455 ( .A(p_input[1405]), .B(n4569), .Z(n4571) );
  XOR U4456 ( .A(n4572), .B(n4573), .Z(n4569) );
  AND U4457 ( .A(n355), .B(n4574), .Z(n4573) );
  XNOR U4458 ( .A(p_input[1421]), .B(n4572), .Z(n4574) );
  XOR U4459 ( .A(n4575), .B(n4576), .Z(n4572) );
  AND U4460 ( .A(n359), .B(n4577), .Z(n4576) );
  XNOR U4461 ( .A(p_input[1437]), .B(n4575), .Z(n4577) );
  XOR U4462 ( .A(n4578), .B(n4579), .Z(n4575) );
  AND U4463 ( .A(n363), .B(n4580), .Z(n4579) );
  XNOR U4464 ( .A(p_input[1453]), .B(n4578), .Z(n4580) );
  XOR U4465 ( .A(n4581), .B(n4582), .Z(n4578) );
  AND U4466 ( .A(n367), .B(n4583), .Z(n4582) );
  XNOR U4467 ( .A(p_input[1469]), .B(n4581), .Z(n4583) );
  XOR U4468 ( .A(n4584), .B(n4585), .Z(n4581) );
  AND U4469 ( .A(n371), .B(n4586), .Z(n4585) );
  XNOR U4470 ( .A(p_input[1485]), .B(n4584), .Z(n4586) );
  XOR U4471 ( .A(n4587), .B(n4588), .Z(n4584) );
  AND U4472 ( .A(n375), .B(n4589), .Z(n4588) );
  XNOR U4473 ( .A(p_input[1501]), .B(n4587), .Z(n4589) );
  XOR U4474 ( .A(n4590), .B(n4591), .Z(n4587) );
  AND U4475 ( .A(n379), .B(n4592), .Z(n4591) );
  XNOR U4476 ( .A(p_input[1517]), .B(n4590), .Z(n4592) );
  XOR U4477 ( .A(n4593), .B(n4594), .Z(n4590) );
  AND U4478 ( .A(n383), .B(n4595), .Z(n4594) );
  XNOR U4479 ( .A(p_input[1533]), .B(n4593), .Z(n4595) );
  XOR U4480 ( .A(n4596), .B(n4597), .Z(n4593) );
  AND U4481 ( .A(n387), .B(n4598), .Z(n4597) );
  XNOR U4482 ( .A(p_input[1549]), .B(n4596), .Z(n4598) );
  XOR U4483 ( .A(n4599), .B(n4600), .Z(n4596) );
  AND U4484 ( .A(n391), .B(n4601), .Z(n4600) );
  XNOR U4485 ( .A(p_input[1565]), .B(n4599), .Z(n4601) );
  XOR U4486 ( .A(n4602), .B(n4603), .Z(n4599) );
  AND U4487 ( .A(n395), .B(n4604), .Z(n4603) );
  XNOR U4488 ( .A(p_input[1581]), .B(n4602), .Z(n4604) );
  XOR U4489 ( .A(n4605), .B(n4606), .Z(n4602) );
  AND U4490 ( .A(n399), .B(n4607), .Z(n4606) );
  XNOR U4491 ( .A(p_input[1597]), .B(n4605), .Z(n4607) );
  XOR U4492 ( .A(n4608), .B(n4609), .Z(n4605) );
  AND U4493 ( .A(n403), .B(n4610), .Z(n4609) );
  XNOR U4494 ( .A(p_input[1613]), .B(n4608), .Z(n4610) );
  XOR U4495 ( .A(n4611), .B(n4612), .Z(n4608) );
  AND U4496 ( .A(n407), .B(n4613), .Z(n4612) );
  XNOR U4497 ( .A(p_input[1629]), .B(n4611), .Z(n4613) );
  XOR U4498 ( .A(n4614), .B(n4615), .Z(n4611) );
  AND U4499 ( .A(n411), .B(n4616), .Z(n4615) );
  XNOR U4500 ( .A(p_input[1645]), .B(n4614), .Z(n4616) );
  XOR U4501 ( .A(n4617), .B(n4618), .Z(n4614) );
  AND U4502 ( .A(n415), .B(n4619), .Z(n4618) );
  XNOR U4503 ( .A(p_input[1661]), .B(n4617), .Z(n4619) );
  XOR U4504 ( .A(n4620), .B(n4621), .Z(n4617) );
  AND U4505 ( .A(n419), .B(n4622), .Z(n4621) );
  XNOR U4506 ( .A(p_input[1677]), .B(n4620), .Z(n4622) );
  XOR U4507 ( .A(n4623), .B(n4624), .Z(n4620) );
  AND U4508 ( .A(n423), .B(n4625), .Z(n4624) );
  XNOR U4509 ( .A(p_input[1693]), .B(n4623), .Z(n4625) );
  XOR U4510 ( .A(n4626), .B(n4627), .Z(n4623) );
  AND U4511 ( .A(n427), .B(n4628), .Z(n4627) );
  XNOR U4512 ( .A(p_input[1709]), .B(n4626), .Z(n4628) );
  XOR U4513 ( .A(n4629), .B(n4630), .Z(n4626) );
  AND U4514 ( .A(n431), .B(n4631), .Z(n4630) );
  XNOR U4515 ( .A(p_input[1725]), .B(n4629), .Z(n4631) );
  XOR U4516 ( .A(n4632), .B(n4633), .Z(n4629) );
  AND U4517 ( .A(n435), .B(n4634), .Z(n4633) );
  XNOR U4518 ( .A(p_input[1741]), .B(n4632), .Z(n4634) );
  XOR U4519 ( .A(n4635), .B(n4636), .Z(n4632) );
  AND U4520 ( .A(n439), .B(n4637), .Z(n4636) );
  XNOR U4521 ( .A(p_input[1757]), .B(n4635), .Z(n4637) );
  XOR U4522 ( .A(n4638), .B(n4639), .Z(n4635) );
  AND U4523 ( .A(n443), .B(n4640), .Z(n4639) );
  XNOR U4524 ( .A(p_input[1773]), .B(n4638), .Z(n4640) );
  XOR U4525 ( .A(n4641), .B(n4642), .Z(n4638) );
  AND U4526 ( .A(n447), .B(n4643), .Z(n4642) );
  XNOR U4527 ( .A(p_input[1789]), .B(n4641), .Z(n4643) );
  XOR U4528 ( .A(n4644), .B(n4645), .Z(n4641) );
  AND U4529 ( .A(n451), .B(n4646), .Z(n4645) );
  XNOR U4530 ( .A(p_input[1805]), .B(n4644), .Z(n4646) );
  XOR U4531 ( .A(n4647), .B(n4648), .Z(n4644) );
  AND U4532 ( .A(n455), .B(n4649), .Z(n4648) );
  XNOR U4533 ( .A(p_input[1821]), .B(n4647), .Z(n4649) );
  XOR U4534 ( .A(n4650), .B(n4651), .Z(n4647) );
  AND U4535 ( .A(n459), .B(n4652), .Z(n4651) );
  XNOR U4536 ( .A(p_input[1837]), .B(n4650), .Z(n4652) );
  XOR U4537 ( .A(n4653), .B(n4654), .Z(n4650) );
  AND U4538 ( .A(n463), .B(n4655), .Z(n4654) );
  XNOR U4539 ( .A(p_input[1853]), .B(n4653), .Z(n4655) );
  XOR U4540 ( .A(n4656), .B(n4657), .Z(n4653) );
  AND U4541 ( .A(n467), .B(n4658), .Z(n4657) );
  XNOR U4542 ( .A(p_input[1869]), .B(n4656), .Z(n4658) );
  XOR U4543 ( .A(n4659), .B(n4660), .Z(n4656) );
  AND U4544 ( .A(n471), .B(n4661), .Z(n4660) );
  XNOR U4545 ( .A(p_input[1885]), .B(n4659), .Z(n4661) );
  XOR U4546 ( .A(n4662), .B(n4663), .Z(n4659) );
  AND U4547 ( .A(n475), .B(n4664), .Z(n4663) );
  XNOR U4548 ( .A(p_input[1901]), .B(n4662), .Z(n4664) );
  XOR U4549 ( .A(n4665), .B(n4666), .Z(n4662) );
  AND U4550 ( .A(n479), .B(n4667), .Z(n4666) );
  XNOR U4551 ( .A(p_input[1917]), .B(n4665), .Z(n4667) );
  XOR U4552 ( .A(n4668), .B(n4669), .Z(n4665) );
  AND U4553 ( .A(n483), .B(n4670), .Z(n4669) );
  XNOR U4554 ( .A(p_input[1933]), .B(n4668), .Z(n4670) );
  XOR U4555 ( .A(n4671), .B(n4672), .Z(n4668) );
  AND U4556 ( .A(n487), .B(n4673), .Z(n4672) );
  XNOR U4557 ( .A(p_input[1949]), .B(n4671), .Z(n4673) );
  XOR U4558 ( .A(n4674), .B(n4675), .Z(n4671) );
  AND U4559 ( .A(n491), .B(n4676), .Z(n4675) );
  XNOR U4560 ( .A(p_input[1965]), .B(n4674), .Z(n4676) );
  XOR U4561 ( .A(n4677), .B(n4678), .Z(n4674) );
  AND U4562 ( .A(n495), .B(n4679), .Z(n4678) );
  XNOR U4563 ( .A(p_input[1981]), .B(n4677), .Z(n4679) );
  XOR U4564 ( .A(n4680), .B(n4681), .Z(n4677) );
  AND U4565 ( .A(n499), .B(n4682), .Z(n4681) );
  XNOR U4566 ( .A(p_input[1997]), .B(n4680), .Z(n4682) );
  XNOR U4567 ( .A(n4683), .B(n4684), .Z(n4680) );
  AND U4568 ( .A(n503), .B(n4685), .Z(n4684) );
  XOR U4569 ( .A(p_input[2013]), .B(n4683), .Z(n4685) );
  XOR U4570 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n4686), .Z(n4683) );
  AND U4571 ( .A(n506), .B(n4687), .Z(n4686) );
  XOR U4572 ( .A(p_input[2029]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n4687)
         );
  XNOR U4573 ( .A(n4688), .B(n4689), .Z(o[12]) );
  AND U4574 ( .A(n3), .B(n4690), .Z(n4688) );
  XNOR U4575 ( .A(p_input[12]), .B(n4689), .Z(n4690) );
  XOR U4576 ( .A(n4691), .B(n4692), .Z(n4689) );
  AND U4577 ( .A(n7), .B(n4693), .Z(n4692) );
  XNOR U4578 ( .A(p_input[28]), .B(n4691), .Z(n4693) );
  XOR U4579 ( .A(n4694), .B(n4695), .Z(n4691) );
  AND U4580 ( .A(n11), .B(n4696), .Z(n4695) );
  XNOR U4581 ( .A(p_input[44]), .B(n4694), .Z(n4696) );
  XOR U4582 ( .A(n4697), .B(n4698), .Z(n4694) );
  AND U4583 ( .A(n15), .B(n4699), .Z(n4698) );
  XNOR U4584 ( .A(p_input[60]), .B(n4697), .Z(n4699) );
  XOR U4585 ( .A(n4700), .B(n4701), .Z(n4697) );
  AND U4586 ( .A(n19), .B(n4702), .Z(n4701) );
  XNOR U4587 ( .A(p_input[76]), .B(n4700), .Z(n4702) );
  XOR U4588 ( .A(n4703), .B(n4704), .Z(n4700) );
  AND U4589 ( .A(n23), .B(n4705), .Z(n4704) );
  XNOR U4590 ( .A(p_input[92]), .B(n4703), .Z(n4705) );
  XOR U4591 ( .A(n4706), .B(n4707), .Z(n4703) );
  AND U4592 ( .A(n27), .B(n4708), .Z(n4707) );
  XNOR U4593 ( .A(p_input[108]), .B(n4706), .Z(n4708) );
  XOR U4594 ( .A(n4709), .B(n4710), .Z(n4706) );
  AND U4595 ( .A(n31), .B(n4711), .Z(n4710) );
  XNOR U4596 ( .A(p_input[124]), .B(n4709), .Z(n4711) );
  XOR U4597 ( .A(n4712), .B(n4713), .Z(n4709) );
  AND U4598 ( .A(n35), .B(n4714), .Z(n4713) );
  XNOR U4599 ( .A(p_input[140]), .B(n4712), .Z(n4714) );
  XOR U4600 ( .A(n4715), .B(n4716), .Z(n4712) );
  AND U4601 ( .A(n39), .B(n4717), .Z(n4716) );
  XNOR U4602 ( .A(p_input[156]), .B(n4715), .Z(n4717) );
  XOR U4603 ( .A(n4718), .B(n4719), .Z(n4715) );
  AND U4604 ( .A(n43), .B(n4720), .Z(n4719) );
  XNOR U4605 ( .A(p_input[172]), .B(n4718), .Z(n4720) );
  XOR U4606 ( .A(n4721), .B(n4722), .Z(n4718) );
  AND U4607 ( .A(n47), .B(n4723), .Z(n4722) );
  XNOR U4608 ( .A(p_input[188]), .B(n4721), .Z(n4723) );
  XOR U4609 ( .A(n4724), .B(n4725), .Z(n4721) );
  AND U4610 ( .A(n51), .B(n4726), .Z(n4725) );
  XNOR U4611 ( .A(p_input[204]), .B(n4724), .Z(n4726) );
  XOR U4612 ( .A(n4727), .B(n4728), .Z(n4724) );
  AND U4613 ( .A(n55), .B(n4729), .Z(n4728) );
  XNOR U4614 ( .A(p_input[220]), .B(n4727), .Z(n4729) );
  XOR U4615 ( .A(n4730), .B(n4731), .Z(n4727) );
  AND U4616 ( .A(n59), .B(n4732), .Z(n4731) );
  XNOR U4617 ( .A(p_input[236]), .B(n4730), .Z(n4732) );
  XOR U4618 ( .A(n4733), .B(n4734), .Z(n4730) );
  AND U4619 ( .A(n63), .B(n4735), .Z(n4734) );
  XNOR U4620 ( .A(p_input[252]), .B(n4733), .Z(n4735) );
  XOR U4621 ( .A(n4736), .B(n4737), .Z(n4733) );
  AND U4622 ( .A(n67), .B(n4738), .Z(n4737) );
  XNOR U4623 ( .A(p_input[268]), .B(n4736), .Z(n4738) );
  XOR U4624 ( .A(n4739), .B(n4740), .Z(n4736) );
  AND U4625 ( .A(n71), .B(n4741), .Z(n4740) );
  XNOR U4626 ( .A(p_input[284]), .B(n4739), .Z(n4741) );
  XOR U4627 ( .A(n4742), .B(n4743), .Z(n4739) );
  AND U4628 ( .A(n75), .B(n4744), .Z(n4743) );
  XNOR U4629 ( .A(p_input[300]), .B(n4742), .Z(n4744) );
  XOR U4630 ( .A(n4745), .B(n4746), .Z(n4742) );
  AND U4631 ( .A(n79), .B(n4747), .Z(n4746) );
  XNOR U4632 ( .A(p_input[316]), .B(n4745), .Z(n4747) );
  XOR U4633 ( .A(n4748), .B(n4749), .Z(n4745) );
  AND U4634 ( .A(n83), .B(n4750), .Z(n4749) );
  XNOR U4635 ( .A(p_input[332]), .B(n4748), .Z(n4750) );
  XOR U4636 ( .A(n4751), .B(n4752), .Z(n4748) );
  AND U4637 ( .A(n87), .B(n4753), .Z(n4752) );
  XNOR U4638 ( .A(p_input[348]), .B(n4751), .Z(n4753) );
  XOR U4639 ( .A(n4754), .B(n4755), .Z(n4751) );
  AND U4640 ( .A(n91), .B(n4756), .Z(n4755) );
  XNOR U4641 ( .A(p_input[364]), .B(n4754), .Z(n4756) );
  XOR U4642 ( .A(n4757), .B(n4758), .Z(n4754) );
  AND U4643 ( .A(n95), .B(n4759), .Z(n4758) );
  XNOR U4644 ( .A(p_input[380]), .B(n4757), .Z(n4759) );
  XOR U4645 ( .A(n4760), .B(n4761), .Z(n4757) );
  AND U4646 ( .A(n99), .B(n4762), .Z(n4761) );
  XNOR U4647 ( .A(p_input[396]), .B(n4760), .Z(n4762) );
  XOR U4648 ( .A(n4763), .B(n4764), .Z(n4760) );
  AND U4649 ( .A(n103), .B(n4765), .Z(n4764) );
  XNOR U4650 ( .A(p_input[412]), .B(n4763), .Z(n4765) );
  XOR U4651 ( .A(n4766), .B(n4767), .Z(n4763) );
  AND U4652 ( .A(n107), .B(n4768), .Z(n4767) );
  XNOR U4653 ( .A(p_input[428]), .B(n4766), .Z(n4768) );
  XOR U4654 ( .A(n4769), .B(n4770), .Z(n4766) );
  AND U4655 ( .A(n111), .B(n4771), .Z(n4770) );
  XNOR U4656 ( .A(p_input[444]), .B(n4769), .Z(n4771) );
  XOR U4657 ( .A(n4772), .B(n4773), .Z(n4769) );
  AND U4658 ( .A(n115), .B(n4774), .Z(n4773) );
  XNOR U4659 ( .A(p_input[460]), .B(n4772), .Z(n4774) );
  XOR U4660 ( .A(n4775), .B(n4776), .Z(n4772) );
  AND U4661 ( .A(n119), .B(n4777), .Z(n4776) );
  XNOR U4662 ( .A(p_input[476]), .B(n4775), .Z(n4777) );
  XOR U4663 ( .A(n4778), .B(n4779), .Z(n4775) );
  AND U4664 ( .A(n123), .B(n4780), .Z(n4779) );
  XNOR U4665 ( .A(p_input[492]), .B(n4778), .Z(n4780) );
  XOR U4666 ( .A(n4781), .B(n4782), .Z(n4778) );
  AND U4667 ( .A(n127), .B(n4783), .Z(n4782) );
  XNOR U4668 ( .A(p_input[508]), .B(n4781), .Z(n4783) );
  XOR U4669 ( .A(n4784), .B(n4785), .Z(n4781) );
  AND U4670 ( .A(n131), .B(n4786), .Z(n4785) );
  XNOR U4671 ( .A(p_input[524]), .B(n4784), .Z(n4786) );
  XOR U4672 ( .A(n4787), .B(n4788), .Z(n4784) );
  AND U4673 ( .A(n135), .B(n4789), .Z(n4788) );
  XNOR U4674 ( .A(p_input[540]), .B(n4787), .Z(n4789) );
  XOR U4675 ( .A(n4790), .B(n4791), .Z(n4787) );
  AND U4676 ( .A(n139), .B(n4792), .Z(n4791) );
  XNOR U4677 ( .A(p_input[556]), .B(n4790), .Z(n4792) );
  XOR U4678 ( .A(n4793), .B(n4794), .Z(n4790) );
  AND U4679 ( .A(n143), .B(n4795), .Z(n4794) );
  XNOR U4680 ( .A(p_input[572]), .B(n4793), .Z(n4795) );
  XOR U4681 ( .A(n4796), .B(n4797), .Z(n4793) );
  AND U4682 ( .A(n147), .B(n4798), .Z(n4797) );
  XNOR U4683 ( .A(p_input[588]), .B(n4796), .Z(n4798) );
  XOR U4684 ( .A(n4799), .B(n4800), .Z(n4796) );
  AND U4685 ( .A(n151), .B(n4801), .Z(n4800) );
  XNOR U4686 ( .A(p_input[604]), .B(n4799), .Z(n4801) );
  XOR U4687 ( .A(n4802), .B(n4803), .Z(n4799) );
  AND U4688 ( .A(n155), .B(n4804), .Z(n4803) );
  XNOR U4689 ( .A(p_input[620]), .B(n4802), .Z(n4804) );
  XOR U4690 ( .A(n4805), .B(n4806), .Z(n4802) );
  AND U4691 ( .A(n159), .B(n4807), .Z(n4806) );
  XNOR U4692 ( .A(p_input[636]), .B(n4805), .Z(n4807) );
  XOR U4693 ( .A(n4808), .B(n4809), .Z(n4805) );
  AND U4694 ( .A(n163), .B(n4810), .Z(n4809) );
  XNOR U4695 ( .A(p_input[652]), .B(n4808), .Z(n4810) );
  XOR U4696 ( .A(n4811), .B(n4812), .Z(n4808) );
  AND U4697 ( .A(n167), .B(n4813), .Z(n4812) );
  XNOR U4698 ( .A(p_input[668]), .B(n4811), .Z(n4813) );
  XOR U4699 ( .A(n4814), .B(n4815), .Z(n4811) );
  AND U4700 ( .A(n171), .B(n4816), .Z(n4815) );
  XNOR U4701 ( .A(p_input[684]), .B(n4814), .Z(n4816) );
  XOR U4702 ( .A(n4817), .B(n4818), .Z(n4814) );
  AND U4703 ( .A(n175), .B(n4819), .Z(n4818) );
  XNOR U4704 ( .A(p_input[700]), .B(n4817), .Z(n4819) );
  XOR U4705 ( .A(n4820), .B(n4821), .Z(n4817) );
  AND U4706 ( .A(n179), .B(n4822), .Z(n4821) );
  XNOR U4707 ( .A(p_input[716]), .B(n4820), .Z(n4822) );
  XOR U4708 ( .A(n4823), .B(n4824), .Z(n4820) );
  AND U4709 ( .A(n183), .B(n4825), .Z(n4824) );
  XNOR U4710 ( .A(p_input[732]), .B(n4823), .Z(n4825) );
  XOR U4711 ( .A(n4826), .B(n4827), .Z(n4823) );
  AND U4712 ( .A(n187), .B(n4828), .Z(n4827) );
  XNOR U4713 ( .A(p_input[748]), .B(n4826), .Z(n4828) );
  XOR U4714 ( .A(n4829), .B(n4830), .Z(n4826) );
  AND U4715 ( .A(n191), .B(n4831), .Z(n4830) );
  XNOR U4716 ( .A(p_input[764]), .B(n4829), .Z(n4831) );
  XOR U4717 ( .A(n4832), .B(n4833), .Z(n4829) );
  AND U4718 ( .A(n195), .B(n4834), .Z(n4833) );
  XNOR U4719 ( .A(p_input[780]), .B(n4832), .Z(n4834) );
  XOR U4720 ( .A(n4835), .B(n4836), .Z(n4832) );
  AND U4721 ( .A(n199), .B(n4837), .Z(n4836) );
  XNOR U4722 ( .A(p_input[796]), .B(n4835), .Z(n4837) );
  XOR U4723 ( .A(n4838), .B(n4839), .Z(n4835) );
  AND U4724 ( .A(n203), .B(n4840), .Z(n4839) );
  XNOR U4725 ( .A(p_input[812]), .B(n4838), .Z(n4840) );
  XOR U4726 ( .A(n4841), .B(n4842), .Z(n4838) );
  AND U4727 ( .A(n207), .B(n4843), .Z(n4842) );
  XNOR U4728 ( .A(p_input[828]), .B(n4841), .Z(n4843) );
  XOR U4729 ( .A(n4844), .B(n4845), .Z(n4841) );
  AND U4730 ( .A(n211), .B(n4846), .Z(n4845) );
  XNOR U4731 ( .A(p_input[844]), .B(n4844), .Z(n4846) );
  XOR U4732 ( .A(n4847), .B(n4848), .Z(n4844) );
  AND U4733 ( .A(n215), .B(n4849), .Z(n4848) );
  XNOR U4734 ( .A(p_input[860]), .B(n4847), .Z(n4849) );
  XOR U4735 ( .A(n4850), .B(n4851), .Z(n4847) );
  AND U4736 ( .A(n219), .B(n4852), .Z(n4851) );
  XNOR U4737 ( .A(p_input[876]), .B(n4850), .Z(n4852) );
  XOR U4738 ( .A(n4853), .B(n4854), .Z(n4850) );
  AND U4739 ( .A(n223), .B(n4855), .Z(n4854) );
  XNOR U4740 ( .A(p_input[892]), .B(n4853), .Z(n4855) );
  XOR U4741 ( .A(n4856), .B(n4857), .Z(n4853) );
  AND U4742 ( .A(n227), .B(n4858), .Z(n4857) );
  XNOR U4743 ( .A(p_input[908]), .B(n4856), .Z(n4858) );
  XOR U4744 ( .A(n4859), .B(n4860), .Z(n4856) );
  AND U4745 ( .A(n231), .B(n4861), .Z(n4860) );
  XNOR U4746 ( .A(p_input[924]), .B(n4859), .Z(n4861) );
  XOR U4747 ( .A(n4862), .B(n4863), .Z(n4859) );
  AND U4748 ( .A(n235), .B(n4864), .Z(n4863) );
  XNOR U4749 ( .A(p_input[940]), .B(n4862), .Z(n4864) );
  XOR U4750 ( .A(n4865), .B(n4866), .Z(n4862) );
  AND U4751 ( .A(n239), .B(n4867), .Z(n4866) );
  XNOR U4752 ( .A(p_input[956]), .B(n4865), .Z(n4867) );
  XOR U4753 ( .A(n4868), .B(n4869), .Z(n4865) );
  AND U4754 ( .A(n243), .B(n4870), .Z(n4869) );
  XNOR U4755 ( .A(p_input[972]), .B(n4868), .Z(n4870) );
  XOR U4756 ( .A(n4871), .B(n4872), .Z(n4868) );
  AND U4757 ( .A(n247), .B(n4873), .Z(n4872) );
  XNOR U4758 ( .A(p_input[988]), .B(n4871), .Z(n4873) );
  XOR U4759 ( .A(n4874), .B(n4875), .Z(n4871) );
  AND U4760 ( .A(n251), .B(n4876), .Z(n4875) );
  XNOR U4761 ( .A(p_input[1004]), .B(n4874), .Z(n4876) );
  XOR U4762 ( .A(n4877), .B(n4878), .Z(n4874) );
  AND U4763 ( .A(n255), .B(n4879), .Z(n4878) );
  XNOR U4764 ( .A(p_input[1020]), .B(n4877), .Z(n4879) );
  XOR U4765 ( .A(n4880), .B(n4881), .Z(n4877) );
  AND U4766 ( .A(n259), .B(n4882), .Z(n4881) );
  XNOR U4767 ( .A(p_input[1036]), .B(n4880), .Z(n4882) );
  XOR U4768 ( .A(n4883), .B(n4884), .Z(n4880) );
  AND U4769 ( .A(n263), .B(n4885), .Z(n4884) );
  XNOR U4770 ( .A(p_input[1052]), .B(n4883), .Z(n4885) );
  XOR U4771 ( .A(n4886), .B(n4887), .Z(n4883) );
  AND U4772 ( .A(n267), .B(n4888), .Z(n4887) );
  XNOR U4773 ( .A(p_input[1068]), .B(n4886), .Z(n4888) );
  XOR U4774 ( .A(n4889), .B(n4890), .Z(n4886) );
  AND U4775 ( .A(n271), .B(n4891), .Z(n4890) );
  XNOR U4776 ( .A(p_input[1084]), .B(n4889), .Z(n4891) );
  XOR U4777 ( .A(n4892), .B(n4893), .Z(n4889) );
  AND U4778 ( .A(n275), .B(n4894), .Z(n4893) );
  XNOR U4779 ( .A(p_input[1100]), .B(n4892), .Z(n4894) );
  XOR U4780 ( .A(n4895), .B(n4896), .Z(n4892) );
  AND U4781 ( .A(n279), .B(n4897), .Z(n4896) );
  XNOR U4782 ( .A(p_input[1116]), .B(n4895), .Z(n4897) );
  XOR U4783 ( .A(n4898), .B(n4899), .Z(n4895) );
  AND U4784 ( .A(n283), .B(n4900), .Z(n4899) );
  XNOR U4785 ( .A(p_input[1132]), .B(n4898), .Z(n4900) );
  XOR U4786 ( .A(n4901), .B(n4902), .Z(n4898) );
  AND U4787 ( .A(n287), .B(n4903), .Z(n4902) );
  XNOR U4788 ( .A(p_input[1148]), .B(n4901), .Z(n4903) );
  XOR U4789 ( .A(n4904), .B(n4905), .Z(n4901) );
  AND U4790 ( .A(n291), .B(n4906), .Z(n4905) );
  XNOR U4791 ( .A(p_input[1164]), .B(n4904), .Z(n4906) );
  XOR U4792 ( .A(n4907), .B(n4908), .Z(n4904) );
  AND U4793 ( .A(n295), .B(n4909), .Z(n4908) );
  XNOR U4794 ( .A(p_input[1180]), .B(n4907), .Z(n4909) );
  XOR U4795 ( .A(n4910), .B(n4911), .Z(n4907) );
  AND U4796 ( .A(n299), .B(n4912), .Z(n4911) );
  XNOR U4797 ( .A(p_input[1196]), .B(n4910), .Z(n4912) );
  XOR U4798 ( .A(n4913), .B(n4914), .Z(n4910) );
  AND U4799 ( .A(n303), .B(n4915), .Z(n4914) );
  XNOR U4800 ( .A(p_input[1212]), .B(n4913), .Z(n4915) );
  XOR U4801 ( .A(n4916), .B(n4917), .Z(n4913) );
  AND U4802 ( .A(n307), .B(n4918), .Z(n4917) );
  XNOR U4803 ( .A(p_input[1228]), .B(n4916), .Z(n4918) );
  XOR U4804 ( .A(n4919), .B(n4920), .Z(n4916) );
  AND U4805 ( .A(n311), .B(n4921), .Z(n4920) );
  XNOR U4806 ( .A(p_input[1244]), .B(n4919), .Z(n4921) );
  XOR U4807 ( .A(n4922), .B(n4923), .Z(n4919) );
  AND U4808 ( .A(n315), .B(n4924), .Z(n4923) );
  XNOR U4809 ( .A(p_input[1260]), .B(n4922), .Z(n4924) );
  XOR U4810 ( .A(n4925), .B(n4926), .Z(n4922) );
  AND U4811 ( .A(n319), .B(n4927), .Z(n4926) );
  XNOR U4812 ( .A(p_input[1276]), .B(n4925), .Z(n4927) );
  XOR U4813 ( .A(n4928), .B(n4929), .Z(n4925) );
  AND U4814 ( .A(n323), .B(n4930), .Z(n4929) );
  XNOR U4815 ( .A(p_input[1292]), .B(n4928), .Z(n4930) );
  XOR U4816 ( .A(n4931), .B(n4932), .Z(n4928) );
  AND U4817 ( .A(n327), .B(n4933), .Z(n4932) );
  XNOR U4818 ( .A(p_input[1308]), .B(n4931), .Z(n4933) );
  XOR U4819 ( .A(n4934), .B(n4935), .Z(n4931) );
  AND U4820 ( .A(n331), .B(n4936), .Z(n4935) );
  XNOR U4821 ( .A(p_input[1324]), .B(n4934), .Z(n4936) );
  XOR U4822 ( .A(n4937), .B(n4938), .Z(n4934) );
  AND U4823 ( .A(n335), .B(n4939), .Z(n4938) );
  XNOR U4824 ( .A(p_input[1340]), .B(n4937), .Z(n4939) );
  XOR U4825 ( .A(n4940), .B(n4941), .Z(n4937) );
  AND U4826 ( .A(n339), .B(n4942), .Z(n4941) );
  XNOR U4827 ( .A(p_input[1356]), .B(n4940), .Z(n4942) );
  XOR U4828 ( .A(n4943), .B(n4944), .Z(n4940) );
  AND U4829 ( .A(n343), .B(n4945), .Z(n4944) );
  XNOR U4830 ( .A(p_input[1372]), .B(n4943), .Z(n4945) );
  XOR U4831 ( .A(n4946), .B(n4947), .Z(n4943) );
  AND U4832 ( .A(n347), .B(n4948), .Z(n4947) );
  XNOR U4833 ( .A(p_input[1388]), .B(n4946), .Z(n4948) );
  XOR U4834 ( .A(n4949), .B(n4950), .Z(n4946) );
  AND U4835 ( .A(n351), .B(n4951), .Z(n4950) );
  XNOR U4836 ( .A(p_input[1404]), .B(n4949), .Z(n4951) );
  XOR U4837 ( .A(n4952), .B(n4953), .Z(n4949) );
  AND U4838 ( .A(n355), .B(n4954), .Z(n4953) );
  XNOR U4839 ( .A(p_input[1420]), .B(n4952), .Z(n4954) );
  XOR U4840 ( .A(n4955), .B(n4956), .Z(n4952) );
  AND U4841 ( .A(n359), .B(n4957), .Z(n4956) );
  XNOR U4842 ( .A(p_input[1436]), .B(n4955), .Z(n4957) );
  XOR U4843 ( .A(n4958), .B(n4959), .Z(n4955) );
  AND U4844 ( .A(n363), .B(n4960), .Z(n4959) );
  XNOR U4845 ( .A(p_input[1452]), .B(n4958), .Z(n4960) );
  XOR U4846 ( .A(n4961), .B(n4962), .Z(n4958) );
  AND U4847 ( .A(n367), .B(n4963), .Z(n4962) );
  XNOR U4848 ( .A(p_input[1468]), .B(n4961), .Z(n4963) );
  XOR U4849 ( .A(n4964), .B(n4965), .Z(n4961) );
  AND U4850 ( .A(n371), .B(n4966), .Z(n4965) );
  XNOR U4851 ( .A(p_input[1484]), .B(n4964), .Z(n4966) );
  XOR U4852 ( .A(n4967), .B(n4968), .Z(n4964) );
  AND U4853 ( .A(n375), .B(n4969), .Z(n4968) );
  XNOR U4854 ( .A(p_input[1500]), .B(n4967), .Z(n4969) );
  XOR U4855 ( .A(n4970), .B(n4971), .Z(n4967) );
  AND U4856 ( .A(n379), .B(n4972), .Z(n4971) );
  XNOR U4857 ( .A(p_input[1516]), .B(n4970), .Z(n4972) );
  XOR U4858 ( .A(n4973), .B(n4974), .Z(n4970) );
  AND U4859 ( .A(n383), .B(n4975), .Z(n4974) );
  XNOR U4860 ( .A(p_input[1532]), .B(n4973), .Z(n4975) );
  XOR U4861 ( .A(n4976), .B(n4977), .Z(n4973) );
  AND U4862 ( .A(n387), .B(n4978), .Z(n4977) );
  XNOR U4863 ( .A(p_input[1548]), .B(n4976), .Z(n4978) );
  XOR U4864 ( .A(n4979), .B(n4980), .Z(n4976) );
  AND U4865 ( .A(n391), .B(n4981), .Z(n4980) );
  XNOR U4866 ( .A(p_input[1564]), .B(n4979), .Z(n4981) );
  XOR U4867 ( .A(n4982), .B(n4983), .Z(n4979) );
  AND U4868 ( .A(n395), .B(n4984), .Z(n4983) );
  XNOR U4869 ( .A(p_input[1580]), .B(n4982), .Z(n4984) );
  XOR U4870 ( .A(n4985), .B(n4986), .Z(n4982) );
  AND U4871 ( .A(n399), .B(n4987), .Z(n4986) );
  XNOR U4872 ( .A(p_input[1596]), .B(n4985), .Z(n4987) );
  XOR U4873 ( .A(n4988), .B(n4989), .Z(n4985) );
  AND U4874 ( .A(n403), .B(n4990), .Z(n4989) );
  XNOR U4875 ( .A(p_input[1612]), .B(n4988), .Z(n4990) );
  XOR U4876 ( .A(n4991), .B(n4992), .Z(n4988) );
  AND U4877 ( .A(n407), .B(n4993), .Z(n4992) );
  XNOR U4878 ( .A(p_input[1628]), .B(n4991), .Z(n4993) );
  XOR U4879 ( .A(n4994), .B(n4995), .Z(n4991) );
  AND U4880 ( .A(n411), .B(n4996), .Z(n4995) );
  XNOR U4881 ( .A(p_input[1644]), .B(n4994), .Z(n4996) );
  XOR U4882 ( .A(n4997), .B(n4998), .Z(n4994) );
  AND U4883 ( .A(n415), .B(n4999), .Z(n4998) );
  XNOR U4884 ( .A(p_input[1660]), .B(n4997), .Z(n4999) );
  XOR U4885 ( .A(n5000), .B(n5001), .Z(n4997) );
  AND U4886 ( .A(n419), .B(n5002), .Z(n5001) );
  XNOR U4887 ( .A(p_input[1676]), .B(n5000), .Z(n5002) );
  XOR U4888 ( .A(n5003), .B(n5004), .Z(n5000) );
  AND U4889 ( .A(n423), .B(n5005), .Z(n5004) );
  XNOR U4890 ( .A(p_input[1692]), .B(n5003), .Z(n5005) );
  XOR U4891 ( .A(n5006), .B(n5007), .Z(n5003) );
  AND U4892 ( .A(n427), .B(n5008), .Z(n5007) );
  XNOR U4893 ( .A(p_input[1708]), .B(n5006), .Z(n5008) );
  XOR U4894 ( .A(n5009), .B(n5010), .Z(n5006) );
  AND U4895 ( .A(n431), .B(n5011), .Z(n5010) );
  XNOR U4896 ( .A(p_input[1724]), .B(n5009), .Z(n5011) );
  XOR U4897 ( .A(n5012), .B(n5013), .Z(n5009) );
  AND U4898 ( .A(n435), .B(n5014), .Z(n5013) );
  XNOR U4899 ( .A(p_input[1740]), .B(n5012), .Z(n5014) );
  XOR U4900 ( .A(n5015), .B(n5016), .Z(n5012) );
  AND U4901 ( .A(n439), .B(n5017), .Z(n5016) );
  XNOR U4902 ( .A(p_input[1756]), .B(n5015), .Z(n5017) );
  XOR U4903 ( .A(n5018), .B(n5019), .Z(n5015) );
  AND U4904 ( .A(n443), .B(n5020), .Z(n5019) );
  XNOR U4905 ( .A(p_input[1772]), .B(n5018), .Z(n5020) );
  XOR U4906 ( .A(n5021), .B(n5022), .Z(n5018) );
  AND U4907 ( .A(n447), .B(n5023), .Z(n5022) );
  XNOR U4908 ( .A(p_input[1788]), .B(n5021), .Z(n5023) );
  XOR U4909 ( .A(n5024), .B(n5025), .Z(n5021) );
  AND U4910 ( .A(n451), .B(n5026), .Z(n5025) );
  XNOR U4911 ( .A(p_input[1804]), .B(n5024), .Z(n5026) );
  XOR U4912 ( .A(n5027), .B(n5028), .Z(n5024) );
  AND U4913 ( .A(n455), .B(n5029), .Z(n5028) );
  XNOR U4914 ( .A(p_input[1820]), .B(n5027), .Z(n5029) );
  XOR U4915 ( .A(n5030), .B(n5031), .Z(n5027) );
  AND U4916 ( .A(n459), .B(n5032), .Z(n5031) );
  XNOR U4917 ( .A(p_input[1836]), .B(n5030), .Z(n5032) );
  XOR U4918 ( .A(n5033), .B(n5034), .Z(n5030) );
  AND U4919 ( .A(n463), .B(n5035), .Z(n5034) );
  XNOR U4920 ( .A(p_input[1852]), .B(n5033), .Z(n5035) );
  XOR U4921 ( .A(n5036), .B(n5037), .Z(n5033) );
  AND U4922 ( .A(n467), .B(n5038), .Z(n5037) );
  XNOR U4923 ( .A(p_input[1868]), .B(n5036), .Z(n5038) );
  XOR U4924 ( .A(n5039), .B(n5040), .Z(n5036) );
  AND U4925 ( .A(n471), .B(n5041), .Z(n5040) );
  XNOR U4926 ( .A(p_input[1884]), .B(n5039), .Z(n5041) );
  XOR U4927 ( .A(n5042), .B(n5043), .Z(n5039) );
  AND U4928 ( .A(n475), .B(n5044), .Z(n5043) );
  XNOR U4929 ( .A(p_input[1900]), .B(n5042), .Z(n5044) );
  XOR U4930 ( .A(n5045), .B(n5046), .Z(n5042) );
  AND U4931 ( .A(n479), .B(n5047), .Z(n5046) );
  XNOR U4932 ( .A(p_input[1916]), .B(n5045), .Z(n5047) );
  XOR U4933 ( .A(n5048), .B(n5049), .Z(n5045) );
  AND U4934 ( .A(n483), .B(n5050), .Z(n5049) );
  XNOR U4935 ( .A(p_input[1932]), .B(n5048), .Z(n5050) );
  XOR U4936 ( .A(n5051), .B(n5052), .Z(n5048) );
  AND U4937 ( .A(n487), .B(n5053), .Z(n5052) );
  XNOR U4938 ( .A(p_input[1948]), .B(n5051), .Z(n5053) );
  XOR U4939 ( .A(n5054), .B(n5055), .Z(n5051) );
  AND U4940 ( .A(n491), .B(n5056), .Z(n5055) );
  XNOR U4941 ( .A(p_input[1964]), .B(n5054), .Z(n5056) );
  XOR U4942 ( .A(n5057), .B(n5058), .Z(n5054) );
  AND U4943 ( .A(n495), .B(n5059), .Z(n5058) );
  XNOR U4944 ( .A(p_input[1980]), .B(n5057), .Z(n5059) );
  XOR U4945 ( .A(n5060), .B(n5061), .Z(n5057) );
  AND U4946 ( .A(n499), .B(n5062), .Z(n5061) );
  XNOR U4947 ( .A(p_input[1996]), .B(n5060), .Z(n5062) );
  XNOR U4948 ( .A(n5063), .B(n5064), .Z(n5060) );
  AND U4949 ( .A(n503), .B(n5065), .Z(n5064) );
  XOR U4950 ( .A(p_input[2012]), .B(n5063), .Z(n5065) );
  XOR U4951 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n5066), .Z(n5063) );
  AND U4952 ( .A(n506), .B(n5067), .Z(n5066) );
  XOR U4953 ( .A(p_input[2028]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n5067)
         );
  XNOR U4954 ( .A(n5068), .B(n5069), .Z(o[11]) );
  AND U4955 ( .A(n3), .B(n5070), .Z(n5068) );
  XNOR U4956 ( .A(p_input[11]), .B(n5069), .Z(n5070) );
  XOR U4957 ( .A(n5071), .B(n5072), .Z(n5069) );
  AND U4958 ( .A(n7), .B(n5073), .Z(n5072) );
  XNOR U4959 ( .A(p_input[27]), .B(n5071), .Z(n5073) );
  XOR U4960 ( .A(n5074), .B(n5075), .Z(n5071) );
  AND U4961 ( .A(n11), .B(n5076), .Z(n5075) );
  XNOR U4962 ( .A(p_input[43]), .B(n5074), .Z(n5076) );
  XOR U4963 ( .A(n5077), .B(n5078), .Z(n5074) );
  AND U4964 ( .A(n15), .B(n5079), .Z(n5078) );
  XNOR U4965 ( .A(p_input[59]), .B(n5077), .Z(n5079) );
  XOR U4966 ( .A(n5080), .B(n5081), .Z(n5077) );
  AND U4967 ( .A(n19), .B(n5082), .Z(n5081) );
  XNOR U4968 ( .A(p_input[75]), .B(n5080), .Z(n5082) );
  XOR U4969 ( .A(n5083), .B(n5084), .Z(n5080) );
  AND U4970 ( .A(n23), .B(n5085), .Z(n5084) );
  XNOR U4971 ( .A(p_input[91]), .B(n5083), .Z(n5085) );
  XOR U4972 ( .A(n5086), .B(n5087), .Z(n5083) );
  AND U4973 ( .A(n27), .B(n5088), .Z(n5087) );
  XNOR U4974 ( .A(p_input[107]), .B(n5086), .Z(n5088) );
  XOR U4975 ( .A(n5089), .B(n5090), .Z(n5086) );
  AND U4976 ( .A(n31), .B(n5091), .Z(n5090) );
  XNOR U4977 ( .A(p_input[123]), .B(n5089), .Z(n5091) );
  XOR U4978 ( .A(n5092), .B(n5093), .Z(n5089) );
  AND U4979 ( .A(n35), .B(n5094), .Z(n5093) );
  XNOR U4980 ( .A(p_input[139]), .B(n5092), .Z(n5094) );
  XOR U4981 ( .A(n5095), .B(n5096), .Z(n5092) );
  AND U4982 ( .A(n39), .B(n5097), .Z(n5096) );
  XNOR U4983 ( .A(p_input[155]), .B(n5095), .Z(n5097) );
  XOR U4984 ( .A(n5098), .B(n5099), .Z(n5095) );
  AND U4985 ( .A(n43), .B(n5100), .Z(n5099) );
  XNOR U4986 ( .A(p_input[171]), .B(n5098), .Z(n5100) );
  XOR U4987 ( .A(n5101), .B(n5102), .Z(n5098) );
  AND U4988 ( .A(n47), .B(n5103), .Z(n5102) );
  XNOR U4989 ( .A(p_input[187]), .B(n5101), .Z(n5103) );
  XOR U4990 ( .A(n5104), .B(n5105), .Z(n5101) );
  AND U4991 ( .A(n51), .B(n5106), .Z(n5105) );
  XNOR U4992 ( .A(p_input[203]), .B(n5104), .Z(n5106) );
  XOR U4993 ( .A(n5107), .B(n5108), .Z(n5104) );
  AND U4994 ( .A(n55), .B(n5109), .Z(n5108) );
  XNOR U4995 ( .A(p_input[219]), .B(n5107), .Z(n5109) );
  XOR U4996 ( .A(n5110), .B(n5111), .Z(n5107) );
  AND U4997 ( .A(n59), .B(n5112), .Z(n5111) );
  XNOR U4998 ( .A(p_input[235]), .B(n5110), .Z(n5112) );
  XOR U4999 ( .A(n5113), .B(n5114), .Z(n5110) );
  AND U5000 ( .A(n63), .B(n5115), .Z(n5114) );
  XNOR U5001 ( .A(p_input[251]), .B(n5113), .Z(n5115) );
  XOR U5002 ( .A(n5116), .B(n5117), .Z(n5113) );
  AND U5003 ( .A(n67), .B(n5118), .Z(n5117) );
  XNOR U5004 ( .A(p_input[267]), .B(n5116), .Z(n5118) );
  XOR U5005 ( .A(n5119), .B(n5120), .Z(n5116) );
  AND U5006 ( .A(n71), .B(n5121), .Z(n5120) );
  XNOR U5007 ( .A(p_input[283]), .B(n5119), .Z(n5121) );
  XOR U5008 ( .A(n5122), .B(n5123), .Z(n5119) );
  AND U5009 ( .A(n75), .B(n5124), .Z(n5123) );
  XNOR U5010 ( .A(p_input[299]), .B(n5122), .Z(n5124) );
  XOR U5011 ( .A(n5125), .B(n5126), .Z(n5122) );
  AND U5012 ( .A(n79), .B(n5127), .Z(n5126) );
  XNOR U5013 ( .A(p_input[315]), .B(n5125), .Z(n5127) );
  XOR U5014 ( .A(n5128), .B(n5129), .Z(n5125) );
  AND U5015 ( .A(n83), .B(n5130), .Z(n5129) );
  XNOR U5016 ( .A(p_input[331]), .B(n5128), .Z(n5130) );
  XOR U5017 ( .A(n5131), .B(n5132), .Z(n5128) );
  AND U5018 ( .A(n87), .B(n5133), .Z(n5132) );
  XNOR U5019 ( .A(p_input[347]), .B(n5131), .Z(n5133) );
  XOR U5020 ( .A(n5134), .B(n5135), .Z(n5131) );
  AND U5021 ( .A(n91), .B(n5136), .Z(n5135) );
  XNOR U5022 ( .A(p_input[363]), .B(n5134), .Z(n5136) );
  XOR U5023 ( .A(n5137), .B(n5138), .Z(n5134) );
  AND U5024 ( .A(n95), .B(n5139), .Z(n5138) );
  XNOR U5025 ( .A(p_input[379]), .B(n5137), .Z(n5139) );
  XOR U5026 ( .A(n5140), .B(n5141), .Z(n5137) );
  AND U5027 ( .A(n99), .B(n5142), .Z(n5141) );
  XNOR U5028 ( .A(p_input[395]), .B(n5140), .Z(n5142) );
  XOR U5029 ( .A(n5143), .B(n5144), .Z(n5140) );
  AND U5030 ( .A(n103), .B(n5145), .Z(n5144) );
  XNOR U5031 ( .A(p_input[411]), .B(n5143), .Z(n5145) );
  XOR U5032 ( .A(n5146), .B(n5147), .Z(n5143) );
  AND U5033 ( .A(n107), .B(n5148), .Z(n5147) );
  XNOR U5034 ( .A(p_input[427]), .B(n5146), .Z(n5148) );
  XOR U5035 ( .A(n5149), .B(n5150), .Z(n5146) );
  AND U5036 ( .A(n111), .B(n5151), .Z(n5150) );
  XNOR U5037 ( .A(p_input[443]), .B(n5149), .Z(n5151) );
  XOR U5038 ( .A(n5152), .B(n5153), .Z(n5149) );
  AND U5039 ( .A(n115), .B(n5154), .Z(n5153) );
  XNOR U5040 ( .A(p_input[459]), .B(n5152), .Z(n5154) );
  XOR U5041 ( .A(n5155), .B(n5156), .Z(n5152) );
  AND U5042 ( .A(n119), .B(n5157), .Z(n5156) );
  XNOR U5043 ( .A(p_input[475]), .B(n5155), .Z(n5157) );
  XOR U5044 ( .A(n5158), .B(n5159), .Z(n5155) );
  AND U5045 ( .A(n123), .B(n5160), .Z(n5159) );
  XNOR U5046 ( .A(p_input[491]), .B(n5158), .Z(n5160) );
  XOR U5047 ( .A(n5161), .B(n5162), .Z(n5158) );
  AND U5048 ( .A(n127), .B(n5163), .Z(n5162) );
  XNOR U5049 ( .A(p_input[507]), .B(n5161), .Z(n5163) );
  XOR U5050 ( .A(n5164), .B(n5165), .Z(n5161) );
  AND U5051 ( .A(n131), .B(n5166), .Z(n5165) );
  XNOR U5052 ( .A(p_input[523]), .B(n5164), .Z(n5166) );
  XOR U5053 ( .A(n5167), .B(n5168), .Z(n5164) );
  AND U5054 ( .A(n135), .B(n5169), .Z(n5168) );
  XNOR U5055 ( .A(p_input[539]), .B(n5167), .Z(n5169) );
  XOR U5056 ( .A(n5170), .B(n5171), .Z(n5167) );
  AND U5057 ( .A(n139), .B(n5172), .Z(n5171) );
  XNOR U5058 ( .A(p_input[555]), .B(n5170), .Z(n5172) );
  XOR U5059 ( .A(n5173), .B(n5174), .Z(n5170) );
  AND U5060 ( .A(n143), .B(n5175), .Z(n5174) );
  XNOR U5061 ( .A(p_input[571]), .B(n5173), .Z(n5175) );
  XOR U5062 ( .A(n5176), .B(n5177), .Z(n5173) );
  AND U5063 ( .A(n147), .B(n5178), .Z(n5177) );
  XNOR U5064 ( .A(p_input[587]), .B(n5176), .Z(n5178) );
  XOR U5065 ( .A(n5179), .B(n5180), .Z(n5176) );
  AND U5066 ( .A(n151), .B(n5181), .Z(n5180) );
  XNOR U5067 ( .A(p_input[603]), .B(n5179), .Z(n5181) );
  XOR U5068 ( .A(n5182), .B(n5183), .Z(n5179) );
  AND U5069 ( .A(n155), .B(n5184), .Z(n5183) );
  XNOR U5070 ( .A(p_input[619]), .B(n5182), .Z(n5184) );
  XOR U5071 ( .A(n5185), .B(n5186), .Z(n5182) );
  AND U5072 ( .A(n159), .B(n5187), .Z(n5186) );
  XNOR U5073 ( .A(p_input[635]), .B(n5185), .Z(n5187) );
  XOR U5074 ( .A(n5188), .B(n5189), .Z(n5185) );
  AND U5075 ( .A(n163), .B(n5190), .Z(n5189) );
  XNOR U5076 ( .A(p_input[651]), .B(n5188), .Z(n5190) );
  XOR U5077 ( .A(n5191), .B(n5192), .Z(n5188) );
  AND U5078 ( .A(n167), .B(n5193), .Z(n5192) );
  XNOR U5079 ( .A(p_input[667]), .B(n5191), .Z(n5193) );
  XOR U5080 ( .A(n5194), .B(n5195), .Z(n5191) );
  AND U5081 ( .A(n171), .B(n5196), .Z(n5195) );
  XNOR U5082 ( .A(p_input[683]), .B(n5194), .Z(n5196) );
  XOR U5083 ( .A(n5197), .B(n5198), .Z(n5194) );
  AND U5084 ( .A(n175), .B(n5199), .Z(n5198) );
  XNOR U5085 ( .A(p_input[699]), .B(n5197), .Z(n5199) );
  XOR U5086 ( .A(n5200), .B(n5201), .Z(n5197) );
  AND U5087 ( .A(n179), .B(n5202), .Z(n5201) );
  XNOR U5088 ( .A(p_input[715]), .B(n5200), .Z(n5202) );
  XOR U5089 ( .A(n5203), .B(n5204), .Z(n5200) );
  AND U5090 ( .A(n183), .B(n5205), .Z(n5204) );
  XNOR U5091 ( .A(p_input[731]), .B(n5203), .Z(n5205) );
  XOR U5092 ( .A(n5206), .B(n5207), .Z(n5203) );
  AND U5093 ( .A(n187), .B(n5208), .Z(n5207) );
  XNOR U5094 ( .A(p_input[747]), .B(n5206), .Z(n5208) );
  XOR U5095 ( .A(n5209), .B(n5210), .Z(n5206) );
  AND U5096 ( .A(n191), .B(n5211), .Z(n5210) );
  XNOR U5097 ( .A(p_input[763]), .B(n5209), .Z(n5211) );
  XOR U5098 ( .A(n5212), .B(n5213), .Z(n5209) );
  AND U5099 ( .A(n195), .B(n5214), .Z(n5213) );
  XNOR U5100 ( .A(p_input[779]), .B(n5212), .Z(n5214) );
  XOR U5101 ( .A(n5215), .B(n5216), .Z(n5212) );
  AND U5102 ( .A(n199), .B(n5217), .Z(n5216) );
  XNOR U5103 ( .A(p_input[795]), .B(n5215), .Z(n5217) );
  XOR U5104 ( .A(n5218), .B(n5219), .Z(n5215) );
  AND U5105 ( .A(n203), .B(n5220), .Z(n5219) );
  XNOR U5106 ( .A(p_input[811]), .B(n5218), .Z(n5220) );
  XOR U5107 ( .A(n5221), .B(n5222), .Z(n5218) );
  AND U5108 ( .A(n207), .B(n5223), .Z(n5222) );
  XNOR U5109 ( .A(p_input[827]), .B(n5221), .Z(n5223) );
  XOR U5110 ( .A(n5224), .B(n5225), .Z(n5221) );
  AND U5111 ( .A(n211), .B(n5226), .Z(n5225) );
  XNOR U5112 ( .A(p_input[843]), .B(n5224), .Z(n5226) );
  XOR U5113 ( .A(n5227), .B(n5228), .Z(n5224) );
  AND U5114 ( .A(n215), .B(n5229), .Z(n5228) );
  XNOR U5115 ( .A(p_input[859]), .B(n5227), .Z(n5229) );
  XOR U5116 ( .A(n5230), .B(n5231), .Z(n5227) );
  AND U5117 ( .A(n219), .B(n5232), .Z(n5231) );
  XNOR U5118 ( .A(p_input[875]), .B(n5230), .Z(n5232) );
  XOR U5119 ( .A(n5233), .B(n5234), .Z(n5230) );
  AND U5120 ( .A(n223), .B(n5235), .Z(n5234) );
  XNOR U5121 ( .A(p_input[891]), .B(n5233), .Z(n5235) );
  XOR U5122 ( .A(n5236), .B(n5237), .Z(n5233) );
  AND U5123 ( .A(n227), .B(n5238), .Z(n5237) );
  XNOR U5124 ( .A(p_input[907]), .B(n5236), .Z(n5238) );
  XOR U5125 ( .A(n5239), .B(n5240), .Z(n5236) );
  AND U5126 ( .A(n231), .B(n5241), .Z(n5240) );
  XNOR U5127 ( .A(p_input[923]), .B(n5239), .Z(n5241) );
  XOR U5128 ( .A(n5242), .B(n5243), .Z(n5239) );
  AND U5129 ( .A(n235), .B(n5244), .Z(n5243) );
  XNOR U5130 ( .A(p_input[939]), .B(n5242), .Z(n5244) );
  XOR U5131 ( .A(n5245), .B(n5246), .Z(n5242) );
  AND U5132 ( .A(n239), .B(n5247), .Z(n5246) );
  XNOR U5133 ( .A(p_input[955]), .B(n5245), .Z(n5247) );
  XOR U5134 ( .A(n5248), .B(n5249), .Z(n5245) );
  AND U5135 ( .A(n243), .B(n5250), .Z(n5249) );
  XNOR U5136 ( .A(p_input[971]), .B(n5248), .Z(n5250) );
  XOR U5137 ( .A(n5251), .B(n5252), .Z(n5248) );
  AND U5138 ( .A(n247), .B(n5253), .Z(n5252) );
  XNOR U5139 ( .A(p_input[987]), .B(n5251), .Z(n5253) );
  XOR U5140 ( .A(n5254), .B(n5255), .Z(n5251) );
  AND U5141 ( .A(n251), .B(n5256), .Z(n5255) );
  XNOR U5142 ( .A(p_input[1003]), .B(n5254), .Z(n5256) );
  XOR U5143 ( .A(n5257), .B(n5258), .Z(n5254) );
  AND U5144 ( .A(n255), .B(n5259), .Z(n5258) );
  XNOR U5145 ( .A(p_input[1019]), .B(n5257), .Z(n5259) );
  XOR U5146 ( .A(n5260), .B(n5261), .Z(n5257) );
  AND U5147 ( .A(n259), .B(n5262), .Z(n5261) );
  XNOR U5148 ( .A(p_input[1035]), .B(n5260), .Z(n5262) );
  XOR U5149 ( .A(n5263), .B(n5264), .Z(n5260) );
  AND U5150 ( .A(n263), .B(n5265), .Z(n5264) );
  XNOR U5151 ( .A(p_input[1051]), .B(n5263), .Z(n5265) );
  XOR U5152 ( .A(n5266), .B(n5267), .Z(n5263) );
  AND U5153 ( .A(n267), .B(n5268), .Z(n5267) );
  XNOR U5154 ( .A(p_input[1067]), .B(n5266), .Z(n5268) );
  XOR U5155 ( .A(n5269), .B(n5270), .Z(n5266) );
  AND U5156 ( .A(n271), .B(n5271), .Z(n5270) );
  XNOR U5157 ( .A(p_input[1083]), .B(n5269), .Z(n5271) );
  XOR U5158 ( .A(n5272), .B(n5273), .Z(n5269) );
  AND U5159 ( .A(n275), .B(n5274), .Z(n5273) );
  XNOR U5160 ( .A(p_input[1099]), .B(n5272), .Z(n5274) );
  XOR U5161 ( .A(n5275), .B(n5276), .Z(n5272) );
  AND U5162 ( .A(n279), .B(n5277), .Z(n5276) );
  XNOR U5163 ( .A(p_input[1115]), .B(n5275), .Z(n5277) );
  XOR U5164 ( .A(n5278), .B(n5279), .Z(n5275) );
  AND U5165 ( .A(n283), .B(n5280), .Z(n5279) );
  XNOR U5166 ( .A(p_input[1131]), .B(n5278), .Z(n5280) );
  XOR U5167 ( .A(n5281), .B(n5282), .Z(n5278) );
  AND U5168 ( .A(n287), .B(n5283), .Z(n5282) );
  XNOR U5169 ( .A(p_input[1147]), .B(n5281), .Z(n5283) );
  XOR U5170 ( .A(n5284), .B(n5285), .Z(n5281) );
  AND U5171 ( .A(n291), .B(n5286), .Z(n5285) );
  XNOR U5172 ( .A(p_input[1163]), .B(n5284), .Z(n5286) );
  XOR U5173 ( .A(n5287), .B(n5288), .Z(n5284) );
  AND U5174 ( .A(n295), .B(n5289), .Z(n5288) );
  XNOR U5175 ( .A(p_input[1179]), .B(n5287), .Z(n5289) );
  XOR U5176 ( .A(n5290), .B(n5291), .Z(n5287) );
  AND U5177 ( .A(n299), .B(n5292), .Z(n5291) );
  XNOR U5178 ( .A(p_input[1195]), .B(n5290), .Z(n5292) );
  XOR U5179 ( .A(n5293), .B(n5294), .Z(n5290) );
  AND U5180 ( .A(n303), .B(n5295), .Z(n5294) );
  XNOR U5181 ( .A(p_input[1211]), .B(n5293), .Z(n5295) );
  XOR U5182 ( .A(n5296), .B(n5297), .Z(n5293) );
  AND U5183 ( .A(n307), .B(n5298), .Z(n5297) );
  XNOR U5184 ( .A(p_input[1227]), .B(n5296), .Z(n5298) );
  XOR U5185 ( .A(n5299), .B(n5300), .Z(n5296) );
  AND U5186 ( .A(n311), .B(n5301), .Z(n5300) );
  XNOR U5187 ( .A(p_input[1243]), .B(n5299), .Z(n5301) );
  XOR U5188 ( .A(n5302), .B(n5303), .Z(n5299) );
  AND U5189 ( .A(n315), .B(n5304), .Z(n5303) );
  XNOR U5190 ( .A(p_input[1259]), .B(n5302), .Z(n5304) );
  XOR U5191 ( .A(n5305), .B(n5306), .Z(n5302) );
  AND U5192 ( .A(n319), .B(n5307), .Z(n5306) );
  XNOR U5193 ( .A(p_input[1275]), .B(n5305), .Z(n5307) );
  XOR U5194 ( .A(n5308), .B(n5309), .Z(n5305) );
  AND U5195 ( .A(n323), .B(n5310), .Z(n5309) );
  XNOR U5196 ( .A(p_input[1291]), .B(n5308), .Z(n5310) );
  XOR U5197 ( .A(n5311), .B(n5312), .Z(n5308) );
  AND U5198 ( .A(n327), .B(n5313), .Z(n5312) );
  XNOR U5199 ( .A(p_input[1307]), .B(n5311), .Z(n5313) );
  XOR U5200 ( .A(n5314), .B(n5315), .Z(n5311) );
  AND U5201 ( .A(n331), .B(n5316), .Z(n5315) );
  XNOR U5202 ( .A(p_input[1323]), .B(n5314), .Z(n5316) );
  XOR U5203 ( .A(n5317), .B(n5318), .Z(n5314) );
  AND U5204 ( .A(n335), .B(n5319), .Z(n5318) );
  XNOR U5205 ( .A(p_input[1339]), .B(n5317), .Z(n5319) );
  XOR U5206 ( .A(n5320), .B(n5321), .Z(n5317) );
  AND U5207 ( .A(n339), .B(n5322), .Z(n5321) );
  XNOR U5208 ( .A(p_input[1355]), .B(n5320), .Z(n5322) );
  XOR U5209 ( .A(n5323), .B(n5324), .Z(n5320) );
  AND U5210 ( .A(n343), .B(n5325), .Z(n5324) );
  XNOR U5211 ( .A(p_input[1371]), .B(n5323), .Z(n5325) );
  XOR U5212 ( .A(n5326), .B(n5327), .Z(n5323) );
  AND U5213 ( .A(n347), .B(n5328), .Z(n5327) );
  XNOR U5214 ( .A(p_input[1387]), .B(n5326), .Z(n5328) );
  XOR U5215 ( .A(n5329), .B(n5330), .Z(n5326) );
  AND U5216 ( .A(n351), .B(n5331), .Z(n5330) );
  XNOR U5217 ( .A(p_input[1403]), .B(n5329), .Z(n5331) );
  XOR U5218 ( .A(n5332), .B(n5333), .Z(n5329) );
  AND U5219 ( .A(n355), .B(n5334), .Z(n5333) );
  XNOR U5220 ( .A(p_input[1419]), .B(n5332), .Z(n5334) );
  XOR U5221 ( .A(n5335), .B(n5336), .Z(n5332) );
  AND U5222 ( .A(n359), .B(n5337), .Z(n5336) );
  XNOR U5223 ( .A(p_input[1435]), .B(n5335), .Z(n5337) );
  XOR U5224 ( .A(n5338), .B(n5339), .Z(n5335) );
  AND U5225 ( .A(n363), .B(n5340), .Z(n5339) );
  XNOR U5226 ( .A(p_input[1451]), .B(n5338), .Z(n5340) );
  XOR U5227 ( .A(n5341), .B(n5342), .Z(n5338) );
  AND U5228 ( .A(n367), .B(n5343), .Z(n5342) );
  XNOR U5229 ( .A(p_input[1467]), .B(n5341), .Z(n5343) );
  XOR U5230 ( .A(n5344), .B(n5345), .Z(n5341) );
  AND U5231 ( .A(n371), .B(n5346), .Z(n5345) );
  XNOR U5232 ( .A(p_input[1483]), .B(n5344), .Z(n5346) );
  XOR U5233 ( .A(n5347), .B(n5348), .Z(n5344) );
  AND U5234 ( .A(n375), .B(n5349), .Z(n5348) );
  XNOR U5235 ( .A(p_input[1499]), .B(n5347), .Z(n5349) );
  XOR U5236 ( .A(n5350), .B(n5351), .Z(n5347) );
  AND U5237 ( .A(n379), .B(n5352), .Z(n5351) );
  XNOR U5238 ( .A(p_input[1515]), .B(n5350), .Z(n5352) );
  XOR U5239 ( .A(n5353), .B(n5354), .Z(n5350) );
  AND U5240 ( .A(n383), .B(n5355), .Z(n5354) );
  XNOR U5241 ( .A(p_input[1531]), .B(n5353), .Z(n5355) );
  XOR U5242 ( .A(n5356), .B(n5357), .Z(n5353) );
  AND U5243 ( .A(n387), .B(n5358), .Z(n5357) );
  XNOR U5244 ( .A(p_input[1547]), .B(n5356), .Z(n5358) );
  XOR U5245 ( .A(n5359), .B(n5360), .Z(n5356) );
  AND U5246 ( .A(n391), .B(n5361), .Z(n5360) );
  XNOR U5247 ( .A(p_input[1563]), .B(n5359), .Z(n5361) );
  XOR U5248 ( .A(n5362), .B(n5363), .Z(n5359) );
  AND U5249 ( .A(n395), .B(n5364), .Z(n5363) );
  XNOR U5250 ( .A(p_input[1579]), .B(n5362), .Z(n5364) );
  XOR U5251 ( .A(n5365), .B(n5366), .Z(n5362) );
  AND U5252 ( .A(n399), .B(n5367), .Z(n5366) );
  XNOR U5253 ( .A(p_input[1595]), .B(n5365), .Z(n5367) );
  XOR U5254 ( .A(n5368), .B(n5369), .Z(n5365) );
  AND U5255 ( .A(n403), .B(n5370), .Z(n5369) );
  XNOR U5256 ( .A(p_input[1611]), .B(n5368), .Z(n5370) );
  XOR U5257 ( .A(n5371), .B(n5372), .Z(n5368) );
  AND U5258 ( .A(n407), .B(n5373), .Z(n5372) );
  XNOR U5259 ( .A(p_input[1627]), .B(n5371), .Z(n5373) );
  XOR U5260 ( .A(n5374), .B(n5375), .Z(n5371) );
  AND U5261 ( .A(n411), .B(n5376), .Z(n5375) );
  XNOR U5262 ( .A(p_input[1643]), .B(n5374), .Z(n5376) );
  XOR U5263 ( .A(n5377), .B(n5378), .Z(n5374) );
  AND U5264 ( .A(n415), .B(n5379), .Z(n5378) );
  XNOR U5265 ( .A(p_input[1659]), .B(n5377), .Z(n5379) );
  XOR U5266 ( .A(n5380), .B(n5381), .Z(n5377) );
  AND U5267 ( .A(n419), .B(n5382), .Z(n5381) );
  XNOR U5268 ( .A(p_input[1675]), .B(n5380), .Z(n5382) );
  XOR U5269 ( .A(n5383), .B(n5384), .Z(n5380) );
  AND U5270 ( .A(n423), .B(n5385), .Z(n5384) );
  XNOR U5271 ( .A(p_input[1691]), .B(n5383), .Z(n5385) );
  XOR U5272 ( .A(n5386), .B(n5387), .Z(n5383) );
  AND U5273 ( .A(n427), .B(n5388), .Z(n5387) );
  XNOR U5274 ( .A(p_input[1707]), .B(n5386), .Z(n5388) );
  XOR U5275 ( .A(n5389), .B(n5390), .Z(n5386) );
  AND U5276 ( .A(n431), .B(n5391), .Z(n5390) );
  XNOR U5277 ( .A(p_input[1723]), .B(n5389), .Z(n5391) );
  XOR U5278 ( .A(n5392), .B(n5393), .Z(n5389) );
  AND U5279 ( .A(n435), .B(n5394), .Z(n5393) );
  XNOR U5280 ( .A(p_input[1739]), .B(n5392), .Z(n5394) );
  XOR U5281 ( .A(n5395), .B(n5396), .Z(n5392) );
  AND U5282 ( .A(n439), .B(n5397), .Z(n5396) );
  XNOR U5283 ( .A(p_input[1755]), .B(n5395), .Z(n5397) );
  XOR U5284 ( .A(n5398), .B(n5399), .Z(n5395) );
  AND U5285 ( .A(n443), .B(n5400), .Z(n5399) );
  XNOR U5286 ( .A(p_input[1771]), .B(n5398), .Z(n5400) );
  XOR U5287 ( .A(n5401), .B(n5402), .Z(n5398) );
  AND U5288 ( .A(n447), .B(n5403), .Z(n5402) );
  XNOR U5289 ( .A(p_input[1787]), .B(n5401), .Z(n5403) );
  XOR U5290 ( .A(n5404), .B(n5405), .Z(n5401) );
  AND U5291 ( .A(n451), .B(n5406), .Z(n5405) );
  XNOR U5292 ( .A(p_input[1803]), .B(n5404), .Z(n5406) );
  XOR U5293 ( .A(n5407), .B(n5408), .Z(n5404) );
  AND U5294 ( .A(n455), .B(n5409), .Z(n5408) );
  XNOR U5295 ( .A(p_input[1819]), .B(n5407), .Z(n5409) );
  XOR U5296 ( .A(n5410), .B(n5411), .Z(n5407) );
  AND U5297 ( .A(n459), .B(n5412), .Z(n5411) );
  XNOR U5298 ( .A(p_input[1835]), .B(n5410), .Z(n5412) );
  XOR U5299 ( .A(n5413), .B(n5414), .Z(n5410) );
  AND U5300 ( .A(n463), .B(n5415), .Z(n5414) );
  XNOR U5301 ( .A(p_input[1851]), .B(n5413), .Z(n5415) );
  XOR U5302 ( .A(n5416), .B(n5417), .Z(n5413) );
  AND U5303 ( .A(n467), .B(n5418), .Z(n5417) );
  XNOR U5304 ( .A(p_input[1867]), .B(n5416), .Z(n5418) );
  XOR U5305 ( .A(n5419), .B(n5420), .Z(n5416) );
  AND U5306 ( .A(n471), .B(n5421), .Z(n5420) );
  XNOR U5307 ( .A(p_input[1883]), .B(n5419), .Z(n5421) );
  XOR U5308 ( .A(n5422), .B(n5423), .Z(n5419) );
  AND U5309 ( .A(n475), .B(n5424), .Z(n5423) );
  XNOR U5310 ( .A(p_input[1899]), .B(n5422), .Z(n5424) );
  XOR U5311 ( .A(n5425), .B(n5426), .Z(n5422) );
  AND U5312 ( .A(n479), .B(n5427), .Z(n5426) );
  XNOR U5313 ( .A(p_input[1915]), .B(n5425), .Z(n5427) );
  XOR U5314 ( .A(n5428), .B(n5429), .Z(n5425) );
  AND U5315 ( .A(n483), .B(n5430), .Z(n5429) );
  XNOR U5316 ( .A(p_input[1931]), .B(n5428), .Z(n5430) );
  XOR U5317 ( .A(n5431), .B(n5432), .Z(n5428) );
  AND U5318 ( .A(n487), .B(n5433), .Z(n5432) );
  XNOR U5319 ( .A(p_input[1947]), .B(n5431), .Z(n5433) );
  XOR U5320 ( .A(n5434), .B(n5435), .Z(n5431) );
  AND U5321 ( .A(n491), .B(n5436), .Z(n5435) );
  XNOR U5322 ( .A(p_input[1963]), .B(n5434), .Z(n5436) );
  XOR U5323 ( .A(n5437), .B(n5438), .Z(n5434) );
  AND U5324 ( .A(n495), .B(n5439), .Z(n5438) );
  XNOR U5325 ( .A(p_input[1979]), .B(n5437), .Z(n5439) );
  XOR U5326 ( .A(n5440), .B(n5441), .Z(n5437) );
  AND U5327 ( .A(n499), .B(n5442), .Z(n5441) );
  XNOR U5328 ( .A(p_input[1995]), .B(n5440), .Z(n5442) );
  XNOR U5329 ( .A(n5443), .B(n5444), .Z(n5440) );
  AND U5330 ( .A(n503), .B(n5445), .Z(n5444) );
  XOR U5331 ( .A(p_input[2011]), .B(n5443), .Z(n5445) );
  XOR U5332 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n5446), .Z(n5443) );
  AND U5333 ( .A(n506), .B(n5447), .Z(n5446) );
  XOR U5334 ( .A(p_input[2027]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n5447)
         );
  XNOR U5335 ( .A(n5448), .B(n5449), .Z(o[10]) );
  AND U5336 ( .A(n3), .B(n5450), .Z(n5448) );
  XNOR U5337 ( .A(p_input[10]), .B(n5449), .Z(n5450) );
  XOR U5338 ( .A(n5451), .B(n5452), .Z(n5449) );
  AND U5339 ( .A(n7), .B(n5453), .Z(n5452) );
  XNOR U5340 ( .A(p_input[26]), .B(n5451), .Z(n5453) );
  XOR U5341 ( .A(n5454), .B(n5455), .Z(n5451) );
  AND U5342 ( .A(n11), .B(n5456), .Z(n5455) );
  XNOR U5343 ( .A(p_input[42]), .B(n5454), .Z(n5456) );
  XOR U5344 ( .A(n5457), .B(n5458), .Z(n5454) );
  AND U5345 ( .A(n15), .B(n5459), .Z(n5458) );
  XNOR U5346 ( .A(p_input[58]), .B(n5457), .Z(n5459) );
  XOR U5347 ( .A(n5460), .B(n5461), .Z(n5457) );
  AND U5348 ( .A(n19), .B(n5462), .Z(n5461) );
  XNOR U5349 ( .A(p_input[74]), .B(n5460), .Z(n5462) );
  XOR U5350 ( .A(n5463), .B(n5464), .Z(n5460) );
  AND U5351 ( .A(n23), .B(n5465), .Z(n5464) );
  XNOR U5352 ( .A(p_input[90]), .B(n5463), .Z(n5465) );
  XOR U5353 ( .A(n5466), .B(n5467), .Z(n5463) );
  AND U5354 ( .A(n27), .B(n5468), .Z(n5467) );
  XNOR U5355 ( .A(p_input[106]), .B(n5466), .Z(n5468) );
  XOR U5356 ( .A(n5469), .B(n5470), .Z(n5466) );
  AND U5357 ( .A(n31), .B(n5471), .Z(n5470) );
  XNOR U5358 ( .A(p_input[122]), .B(n5469), .Z(n5471) );
  XOR U5359 ( .A(n5472), .B(n5473), .Z(n5469) );
  AND U5360 ( .A(n35), .B(n5474), .Z(n5473) );
  XNOR U5361 ( .A(p_input[138]), .B(n5472), .Z(n5474) );
  XOR U5362 ( .A(n5475), .B(n5476), .Z(n5472) );
  AND U5363 ( .A(n39), .B(n5477), .Z(n5476) );
  XNOR U5364 ( .A(p_input[154]), .B(n5475), .Z(n5477) );
  XOR U5365 ( .A(n5478), .B(n5479), .Z(n5475) );
  AND U5366 ( .A(n43), .B(n5480), .Z(n5479) );
  XNOR U5367 ( .A(p_input[170]), .B(n5478), .Z(n5480) );
  XOR U5368 ( .A(n5481), .B(n5482), .Z(n5478) );
  AND U5369 ( .A(n47), .B(n5483), .Z(n5482) );
  XNOR U5370 ( .A(p_input[186]), .B(n5481), .Z(n5483) );
  XOR U5371 ( .A(n5484), .B(n5485), .Z(n5481) );
  AND U5372 ( .A(n51), .B(n5486), .Z(n5485) );
  XNOR U5373 ( .A(p_input[202]), .B(n5484), .Z(n5486) );
  XOR U5374 ( .A(n5487), .B(n5488), .Z(n5484) );
  AND U5375 ( .A(n55), .B(n5489), .Z(n5488) );
  XNOR U5376 ( .A(p_input[218]), .B(n5487), .Z(n5489) );
  XOR U5377 ( .A(n5490), .B(n5491), .Z(n5487) );
  AND U5378 ( .A(n59), .B(n5492), .Z(n5491) );
  XNOR U5379 ( .A(p_input[234]), .B(n5490), .Z(n5492) );
  XOR U5380 ( .A(n5493), .B(n5494), .Z(n5490) );
  AND U5381 ( .A(n63), .B(n5495), .Z(n5494) );
  XNOR U5382 ( .A(p_input[250]), .B(n5493), .Z(n5495) );
  XOR U5383 ( .A(n5496), .B(n5497), .Z(n5493) );
  AND U5384 ( .A(n67), .B(n5498), .Z(n5497) );
  XNOR U5385 ( .A(p_input[266]), .B(n5496), .Z(n5498) );
  XOR U5386 ( .A(n5499), .B(n5500), .Z(n5496) );
  AND U5387 ( .A(n71), .B(n5501), .Z(n5500) );
  XNOR U5388 ( .A(p_input[282]), .B(n5499), .Z(n5501) );
  XOR U5389 ( .A(n5502), .B(n5503), .Z(n5499) );
  AND U5390 ( .A(n75), .B(n5504), .Z(n5503) );
  XNOR U5391 ( .A(p_input[298]), .B(n5502), .Z(n5504) );
  XOR U5392 ( .A(n5505), .B(n5506), .Z(n5502) );
  AND U5393 ( .A(n79), .B(n5507), .Z(n5506) );
  XNOR U5394 ( .A(p_input[314]), .B(n5505), .Z(n5507) );
  XOR U5395 ( .A(n5508), .B(n5509), .Z(n5505) );
  AND U5396 ( .A(n83), .B(n5510), .Z(n5509) );
  XNOR U5397 ( .A(p_input[330]), .B(n5508), .Z(n5510) );
  XOR U5398 ( .A(n5511), .B(n5512), .Z(n5508) );
  AND U5399 ( .A(n87), .B(n5513), .Z(n5512) );
  XNOR U5400 ( .A(p_input[346]), .B(n5511), .Z(n5513) );
  XOR U5401 ( .A(n5514), .B(n5515), .Z(n5511) );
  AND U5402 ( .A(n91), .B(n5516), .Z(n5515) );
  XNOR U5403 ( .A(p_input[362]), .B(n5514), .Z(n5516) );
  XOR U5404 ( .A(n5517), .B(n5518), .Z(n5514) );
  AND U5405 ( .A(n95), .B(n5519), .Z(n5518) );
  XNOR U5406 ( .A(p_input[378]), .B(n5517), .Z(n5519) );
  XOR U5407 ( .A(n5520), .B(n5521), .Z(n5517) );
  AND U5408 ( .A(n99), .B(n5522), .Z(n5521) );
  XNOR U5409 ( .A(p_input[394]), .B(n5520), .Z(n5522) );
  XOR U5410 ( .A(n5523), .B(n5524), .Z(n5520) );
  AND U5411 ( .A(n103), .B(n5525), .Z(n5524) );
  XNOR U5412 ( .A(p_input[410]), .B(n5523), .Z(n5525) );
  XOR U5413 ( .A(n5526), .B(n5527), .Z(n5523) );
  AND U5414 ( .A(n107), .B(n5528), .Z(n5527) );
  XNOR U5415 ( .A(p_input[426]), .B(n5526), .Z(n5528) );
  XOR U5416 ( .A(n5529), .B(n5530), .Z(n5526) );
  AND U5417 ( .A(n111), .B(n5531), .Z(n5530) );
  XNOR U5418 ( .A(p_input[442]), .B(n5529), .Z(n5531) );
  XOR U5419 ( .A(n5532), .B(n5533), .Z(n5529) );
  AND U5420 ( .A(n115), .B(n5534), .Z(n5533) );
  XNOR U5421 ( .A(p_input[458]), .B(n5532), .Z(n5534) );
  XOR U5422 ( .A(n5535), .B(n5536), .Z(n5532) );
  AND U5423 ( .A(n119), .B(n5537), .Z(n5536) );
  XNOR U5424 ( .A(p_input[474]), .B(n5535), .Z(n5537) );
  XOR U5425 ( .A(n5538), .B(n5539), .Z(n5535) );
  AND U5426 ( .A(n123), .B(n5540), .Z(n5539) );
  XNOR U5427 ( .A(p_input[490]), .B(n5538), .Z(n5540) );
  XOR U5428 ( .A(n5541), .B(n5542), .Z(n5538) );
  AND U5429 ( .A(n127), .B(n5543), .Z(n5542) );
  XNOR U5430 ( .A(p_input[506]), .B(n5541), .Z(n5543) );
  XOR U5431 ( .A(n5544), .B(n5545), .Z(n5541) );
  AND U5432 ( .A(n131), .B(n5546), .Z(n5545) );
  XNOR U5433 ( .A(p_input[522]), .B(n5544), .Z(n5546) );
  XOR U5434 ( .A(n5547), .B(n5548), .Z(n5544) );
  AND U5435 ( .A(n135), .B(n5549), .Z(n5548) );
  XNOR U5436 ( .A(p_input[538]), .B(n5547), .Z(n5549) );
  XOR U5437 ( .A(n5550), .B(n5551), .Z(n5547) );
  AND U5438 ( .A(n139), .B(n5552), .Z(n5551) );
  XNOR U5439 ( .A(p_input[554]), .B(n5550), .Z(n5552) );
  XOR U5440 ( .A(n5553), .B(n5554), .Z(n5550) );
  AND U5441 ( .A(n143), .B(n5555), .Z(n5554) );
  XNOR U5442 ( .A(p_input[570]), .B(n5553), .Z(n5555) );
  XOR U5443 ( .A(n5556), .B(n5557), .Z(n5553) );
  AND U5444 ( .A(n147), .B(n5558), .Z(n5557) );
  XNOR U5445 ( .A(p_input[586]), .B(n5556), .Z(n5558) );
  XOR U5446 ( .A(n5559), .B(n5560), .Z(n5556) );
  AND U5447 ( .A(n151), .B(n5561), .Z(n5560) );
  XNOR U5448 ( .A(p_input[602]), .B(n5559), .Z(n5561) );
  XOR U5449 ( .A(n5562), .B(n5563), .Z(n5559) );
  AND U5450 ( .A(n155), .B(n5564), .Z(n5563) );
  XNOR U5451 ( .A(p_input[618]), .B(n5562), .Z(n5564) );
  XOR U5452 ( .A(n5565), .B(n5566), .Z(n5562) );
  AND U5453 ( .A(n159), .B(n5567), .Z(n5566) );
  XNOR U5454 ( .A(p_input[634]), .B(n5565), .Z(n5567) );
  XOR U5455 ( .A(n5568), .B(n5569), .Z(n5565) );
  AND U5456 ( .A(n163), .B(n5570), .Z(n5569) );
  XNOR U5457 ( .A(p_input[650]), .B(n5568), .Z(n5570) );
  XOR U5458 ( .A(n5571), .B(n5572), .Z(n5568) );
  AND U5459 ( .A(n167), .B(n5573), .Z(n5572) );
  XNOR U5460 ( .A(p_input[666]), .B(n5571), .Z(n5573) );
  XOR U5461 ( .A(n5574), .B(n5575), .Z(n5571) );
  AND U5462 ( .A(n171), .B(n5576), .Z(n5575) );
  XNOR U5463 ( .A(p_input[682]), .B(n5574), .Z(n5576) );
  XOR U5464 ( .A(n5577), .B(n5578), .Z(n5574) );
  AND U5465 ( .A(n175), .B(n5579), .Z(n5578) );
  XNOR U5466 ( .A(p_input[698]), .B(n5577), .Z(n5579) );
  XOR U5467 ( .A(n5580), .B(n5581), .Z(n5577) );
  AND U5468 ( .A(n179), .B(n5582), .Z(n5581) );
  XNOR U5469 ( .A(p_input[714]), .B(n5580), .Z(n5582) );
  XOR U5470 ( .A(n5583), .B(n5584), .Z(n5580) );
  AND U5471 ( .A(n183), .B(n5585), .Z(n5584) );
  XNOR U5472 ( .A(p_input[730]), .B(n5583), .Z(n5585) );
  XOR U5473 ( .A(n5586), .B(n5587), .Z(n5583) );
  AND U5474 ( .A(n187), .B(n5588), .Z(n5587) );
  XNOR U5475 ( .A(p_input[746]), .B(n5586), .Z(n5588) );
  XOR U5476 ( .A(n5589), .B(n5590), .Z(n5586) );
  AND U5477 ( .A(n191), .B(n5591), .Z(n5590) );
  XNOR U5478 ( .A(p_input[762]), .B(n5589), .Z(n5591) );
  XOR U5479 ( .A(n5592), .B(n5593), .Z(n5589) );
  AND U5480 ( .A(n195), .B(n5594), .Z(n5593) );
  XNOR U5481 ( .A(p_input[778]), .B(n5592), .Z(n5594) );
  XOR U5482 ( .A(n5595), .B(n5596), .Z(n5592) );
  AND U5483 ( .A(n199), .B(n5597), .Z(n5596) );
  XNOR U5484 ( .A(p_input[794]), .B(n5595), .Z(n5597) );
  XOR U5485 ( .A(n5598), .B(n5599), .Z(n5595) );
  AND U5486 ( .A(n203), .B(n5600), .Z(n5599) );
  XNOR U5487 ( .A(p_input[810]), .B(n5598), .Z(n5600) );
  XOR U5488 ( .A(n5601), .B(n5602), .Z(n5598) );
  AND U5489 ( .A(n207), .B(n5603), .Z(n5602) );
  XNOR U5490 ( .A(p_input[826]), .B(n5601), .Z(n5603) );
  XOR U5491 ( .A(n5604), .B(n5605), .Z(n5601) );
  AND U5492 ( .A(n211), .B(n5606), .Z(n5605) );
  XNOR U5493 ( .A(p_input[842]), .B(n5604), .Z(n5606) );
  XOR U5494 ( .A(n5607), .B(n5608), .Z(n5604) );
  AND U5495 ( .A(n215), .B(n5609), .Z(n5608) );
  XNOR U5496 ( .A(p_input[858]), .B(n5607), .Z(n5609) );
  XOR U5497 ( .A(n5610), .B(n5611), .Z(n5607) );
  AND U5498 ( .A(n219), .B(n5612), .Z(n5611) );
  XNOR U5499 ( .A(p_input[874]), .B(n5610), .Z(n5612) );
  XOR U5500 ( .A(n5613), .B(n5614), .Z(n5610) );
  AND U5501 ( .A(n223), .B(n5615), .Z(n5614) );
  XNOR U5502 ( .A(p_input[890]), .B(n5613), .Z(n5615) );
  XOR U5503 ( .A(n5616), .B(n5617), .Z(n5613) );
  AND U5504 ( .A(n227), .B(n5618), .Z(n5617) );
  XNOR U5505 ( .A(p_input[906]), .B(n5616), .Z(n5618) );
  XOR U5506 ( .A(n5619), .B(n5620), .Z(n5616) );
  AND U5507 ( .A(n231), .B(n5621), .Z(n5620) );
  XNOR U5508 ( .A(p_input[922]), .B(n5619), .Z(n5621) );
  XOR U5509 ( .A(n5622), .B(n5623), .Z(n5619) );
  AND U5510 ( .A(n235), .B(n5624), .Z(n5623) );
  XNOR U5511 ( .A(p_input[938]), .B(n5622), .Z(n5624) );
  XOR U5512 ( .A(n5625), .B(n5626), .Z(n5622) );
  AND U5513 ( .A(n239), .B(n5627), .Z(n5626) );
  XNOR U5514 ( .A(p_input[954]), .B(n5625), .Z(n5627) );
  XOR U5515 ( .A(n5628), .B(n5629), .Z(n5625) );
  AND U5516 ( .A(n243), .B(n5630), .Z(n5629) );
  XNOR U5517 ( .A(p_input[970]), .B(n5628), .Z(n5630) );
  XOR U5518 ( .A(n5631), .B(n5632), .Z(n5628) );
  AND U5519 ( .A(n247), .B(n5633), .Z(n5632) );
  XNOR U5520 ( .A(p_input[986]), .B(n5631), .Z(n5633) );
  XOR U5521 ( .A(n5634), .B(n5635), .Z(n5631) );
  AND U5522 ( .A(n251), .B(n5636), .Z(n5635) );
  XNOR U5523 ( .A(p_input[1002]), .B(n5634), .Z(n5636) );
  XOR U5524 ( .A(n5637), .B(n5638), .Z(n5634) );
  AND U5525 ( .A(n255), .B(n5639), .Z(n5638) );
  XNOR U5526 ( .A(p_input[1018]), .B(n5637), .Z(n5639) );
  XOR U5527 ( .A(n5640), .B(n5641), .Z(n5637) );
  AND U5528 ( .A(n259), .B(n5642), .Z(n5641) );
  XNOR U5529 ( .A(p_input[1034]), .B(n5640), .Z(n5642) );
  XOR U5530 ( .A(n5643), .B(n5644), .Z(n5640) );
  AND U5531 ( .A(n263), .B(n5645), .Z(n5644) );
  XNOR U5532 ( .A(p_input[1050]), .B(n5643), .Z(n5645) );
  XOR U5533 ( .A(n5646), .B(n5647), .Z(n5643) );
  AND U5534 ( .A(n267), .B(n5648), .Z(n5647) );
  XNOR U5535 ( .A(p_input[1066]), .B(n5646), .Z(n5648) );
  XOR U5536 ( .A(n5649), .B(n5650), .Z(n5646) );
  AND U5537 ( .A(n271), .B(n5651), .Z(n5650) );
  XNOR U5538 ( .A(p_input[1082]), .B(n5649), .Z(n5651) );
  XOR U5539 ( .A(n5652), .B(n5653), .Z(n5649) );
  AND U5540 ( .A(n275), .B(n5654), .Z(n5653) );
  XNOR U5541 ( .A(p_input[1098]), .B(n5652), .Z(n5654) );
  XOR U5542 ( .A(n5655), .B(n5656), .Z(n5652) );
  AND U5543 ( .A(n279), .B(n5657), .Z(n5656) );
  XNOR U5544 ( .A(p_input[1114]), .B(n5655), .Z(n5657) );
  XOR U5545 ( .A(n5658), .B(n5659), .Z(n5655) );
  AND U5546 ( .A(n283), .B(n5660), .Z(n5659) );
  XNOR U5547 ( .A(p_input[1130]), .B(n5658), .Z(n5660) );
  XOR U5548 ( .A(n5661), .B(n5662), .Z(n5658) );
  AND U5549 ( .A(n287), .B(n5663), .Z(n5662) );
  XNOR U5550 ( .A(p_input[1146]), .B(n5661), .Z(n5663) );
  XOR U5551 ( .A(n5664), .B(n5665), .Z(n5661) );
  AND U5552 ( .A(n291), .B(n5666), .Z(n5665) );
  XNOR U5553 ( .A(p_input[1162]), .B(n5664), .Z(n5666) );
  XOR U5554 ( .A(n5667), .B(n5668), .Z(n5664) );
  AND U5555 ( .A(n295), .B(n5669), .Z(n5668) );
  XNOR U5556 ( .A(p_input[1178]), .B(n5667), .Z(n5669) );
  XOR U5557 ( .A(n5670), .B(n5671), .Z(n5667) );
  AND U5558 ( .A(n299), .B(n5672), .Z(n5671) );
  XNOR U5559 ( .A(p_input[1194]), .B(n5670), .Z(n5672) );
  XOR U5560 ( .A(n5673), .B(n5674), .Z(n5670) );
  AND U5561 ( .A(n303), .B(n5675), .Z(n5674) );
  XNOR U5562 ( .A(p_input[1210]), .B(n5673), .Z(n5675) );
  XOR U5563 ( .A(n5676), .B(n5677), .Z(n5673) );
  AND U5564 ( .A(n307), .B(n5678), .Z(n5677) );
  XNOR U5565 ( .A(p_input[1226]), .B(n5676), .Z(n5678) );
  XOR U5566 ( .A(n5679), .B(n5680), .Z(n5676) );
  AND U5567 ( .A(n311), .B(n5681), .Z(n5680) );
  XNOR U5568 ( .A(p_input[1242]), .B(n5679), .Z(n5681) );
  XOR U5569 ( .A(n5682), .B(n5683), .Z(n5679) );
  AND U5570 ( .A(n315), .B(n5684), .Z(n5683) );
  XNOR U5571 ( .A(p_input[1258]), .B(n5682), .Z(n5684) );
  XOR U5572 ( .A(n5685), .B(n5686), .Z(n5682) );
  AND U5573 ( .A(n319), .B(n5687), .Z(n5686) );
  XNOR U5574 ( .A(p_input[1274]), .B(n5685), .Z(n5687) );
  XOR U5575 ( .A(n5688), .B(n5689), .Z(n5685) );
  AND U5576 ( .A(n323), .B(n5690), .Z(n5689) );
  XNOR U5577 ( .A(p_input[1290]), .B(n5688), .Z(n5690) );
  XOR U5578 ( .A(n5691), .B(n5692), .Z(n5688) );
  AND U5579 ( .A(n327), .B(n5693), .Z(n5692) );
  XNOR U5580 ( .A(p_input[1306]), .B(n5691), .Z(n5693) );
  XOR U5581 ( .A(n5694), .B(n5695), .Z(n5691) );
  AND U5582 ( .A(n331), .B(n5696), .Z(n5695) );
  XNOR U5583 ( .A(p_input[1322]), .B(n5694), .Z(n5696) );
  XOR U5584 ( .A(n5697), .B(n5698), .Z(n5694) );
  AND U5585 ( .A(n335), .B(n5699), .Z(n5698) );
  XNOR U5586 ( .A(p_input[1338]), .B(n5697), .Z(n5699) );
  XOR U5587 ( .A(n5700), .B(n5701), .Z(n5697) );
  AND U5588 ( .A(n339), .B(n5702), .Z(n5701) );
  XNOR U5589 ( .A(p_input[1354]), .B(n5700), .Z(n5702) );
  XOR U5590 ( .A(n5703), .B(n5704), .Z(n5700) );
  AND U5591 ( .A(n343), .B(n5705), .Z(n5704) );
  XNOR U5592 ( .A(p_input[1370]), .B(n5703), .Z(n5705) );
  XOR U5593 ( .A(n5706), .B(n5707), .Z(n5703) );
  AND U5594 ( .A(n347), .B(n5708), .Z(n5707) );
  XNOR U5595 ( .A(p_input[1386]), .B(n5706), .Z(n5708) );
  XOR U5596 ( .A(n5709), .B(n5710), .Z(n5706) );
  AND U5597 ( .A(n351), .B(n5711), .Z(n5710) );
  XNOR U5598 ( .A(p_input[1402]), .B(n5709), .Z(n5711) );
  XOR U5599 ( .A(n5712), .B(n5713), .Z(n5709) );
  AND U5600 ( .A(n355), .B(n5714), .Z(n5713) );
  XNOR U5601 ( .A(p_input[1418]), .B(n5712), .Z(n5714) );
  XOR U5602 ( .A(n5715), .B(n5716), .Z(n5712) );
  AND U5603 ( .A(n359), .B(n5717), .Z(n5716) );
  XNOR U5604 ( .A(p_input[1434]), .B(n5715), .Z(n5717) );
  XOR U5605 ( .A(n5718), .B(n5719), .Z(n5715) );
  AND U5606 ( .A(n363), .B(n5720), .Z(n5719) );
  XNOR U5607 ( .A(p_input[1450]), .B(n5718), .Z(n5720) );
  XOR U5608 ( .A(n5721), .B(n5722), .Z(n5718) );
  AND U5609 ( .A(n367), .B(n5723), .Z(n5722) );
  XNOR U5610 ( .A(p_input[1466]), .B(n5721), .Z(n5723) );
  XOR U5611 ( .A(n5724), .B(n5725), .Z(n5721) );
  AND U5612 ( .A(n371), .B(n5726), .Z(n5725) );
  XNOR U5613 ( .A(p_input[1482]), .B(n5724), .Z(n5726) );
  XOR U5614 ( .A(n5727), .B(n5728), .Z(n5724) );
  AND U5615 ( .A(n375), .B(n5729), .Z(n5728) );
  XNOR U5616 ( .A(p_input[1498]), .B(n5727), .Z(n5729) );
  XOR U5617 ( .A(n5730), .B(n5731), .Z(n5727) );
  AND U5618 ( .A(n379), .B(n5732), .Z(n5731) );
  XNOR U5619 ( .A(p_input[1514]), .B(n5730), .Z(n5732) );
  XOR U5620 ( .A(n5733), .B(n5734), .Z(n5730) );
  AND U5621 ( .A(n383), .B(n5735), .Z(n5734) );
  XNOR U5622 ( .A(p_input[1530]), .B(n5733), .Z(n5735) );
  XOR U5623 ( .A(n5736), .B(n5737), .Z(n5733) );
  AND U5624 ( .A(n387), .B(n5738), .Z(n5737) );
  XNOR U5625 ( .A(p_input[1546]), .B(n5736), .Z(n5738) );
  XOR U5626 ( .A(n5739), .B(n5740), .Z(n5736) );
  AND U5627 ( .A(n391), .B(n5741), .Z(n5740) );
  XNOR U5628 ( .A(p_input[1562]), .B(n5739), .Z(n5741) );
  XOR U5629 ( .A(n5742), .B(n5743), .Z(n5739) );
  AND U5630 ( .A(n395), .B(n5744), .Z(n5743) );
  XNOR U5631 ( .A(p_input[1578]), .B(n5742), .Z(n5744) );
  XOR U5632 ( .A(n5745), .B(n5746), .Z(n5742) );
  AND U5633 ( .A(n399), .B(n5747), .Z(n5746) );
  XNOR U5634 ( .A(p_input[1594]), .B(n5745), .Z(n5747) );
  XOR U5635 ( .A(n5748), .B(n5749), .Z(n5745) );
  AND U5636 ( .A(n403), .B(n5750), .Z(n5749) );
  XNOR U5637 ( .A(p_input[1610]), .B(n5748), .Z(n5750) );
  XOR U5638 ( .A(n5751), .B(n5752), .Z(n5748) );
  AND U5639 ( .A(n407), .B(n5753), .Z(n5752) );
  XNOR U5640 ( .A(p_input[1626]), .B(n5751), .Z(n5753) );
  XOR U5641 ( .A(n5754), .B(n5755), .Z(n5751) );
  AND U5642 ( .A(n411), .B(n5756), .Z(n5755) );
  XNOR U5643 ( .A(p_input[1642]), .B(n5754), .Z(n5756) );
  XOR U5644 ( .A(n5757), .B(n5758), .Z(n5754) );
  AND U5645 ( .A(n415), .B(n5759), .Z(n5758) );
  XNOR U5646 ( .A(p_input[1658]), .B(n5757), .Z(n5759) );
  XOR U5647 ( .A(n5760), .B(n5761), .Z(n5757) );
  AND U5648 ( .A(n419), .B(n5762), .Z(n5761) );
  XNOR U5649 ( .A(p_input[1674]), .B(n5760), .Z(n5762) );
  XOR U5650 ( .A(n5763), .B(n5764), .Z(n5760) );
  AND U5651 ( .A(n423), .B(n5765), .Z(n5764) );
  XNOR U5652 ( .A(p_input[1690]), .B(n5763), .Z(n5765) );
  XOR U5653 ( .A(n5766), .B(n5767), .Z(n5763) );
  AND U5654 ( .A(n427), .B(n5768), .Z(n5767) );
  XNOR U5655 ( .A(p_input[1706]), .B(n5766), .Z(n5768) );
  XOR U5656 ( .A(n5769), .B(n5770), .Z(n5766) );
  AND U5657 ( .A(n431), .B(n5771), .Z(n5770) );
  XNOR U5658 ( .A(p_input[1722]), .B(n5769), .Z(n5771) );
  XOR U5659 ( .A(n5772), .B(n5773), .Z(n5769) );
  AND U5660 ( .A(n435), .B(n5774), .Z(n5773) );
  XNOR U5661 ( .A(p_input[1738]), .B(n5772), .Z(n5774) );
  XOR U5662 ( .A(n5775), .B(n5776), .Z(n5772) );
  AND U5663 ( .A(n439), .B(n5777), .Z(n5776) );
  XNOR U5664 ( .A(p_input[1754]), .B(n5775), .Z(n5777) );
  XOR U5665 ( .A(n5778), .B(n5779), .Z(n5775) );
  AND U5666 ( .A(n443), .B(n5780), .Z(n5779) );
  XNOR U5667 ( .A(p_input[1770]), .B(n5778), .Z(n5780) );
  XOR U5668 ( .A(n5781), .B(n5782), .Z(n5778) );
  AND U5669 ( .A(n447), .B(n5783), .Z(n5782) );
  XNOR U5670 ( .A(p_input[1786]), .B(n5781), .Z(n5783) );
  XOR U5671 ( .A(n5784), .B(n5785), .Z(n5781) );
  AND U5672 ( .A(n451), .B(n5786), .Z(n5785) );
  XNOR U5673 ( .A(p_input[1802]), .B(n5784), .Z(n5786) );
  XOR U5674 ( .A(n5787), .B(n5788), .Z(n5784) );
  AND U5675 ( .A(n455), .B(n5789), .Z(n5788) );
  XNOR U5676 ( .A(p_input[1818]), .B(n5787), .Z(n5789) );
  XOR U5677 ( .A(n5790), .B(n5791), .Z(n5787) );
  AND U5678 ( .A(n459), .B(n5792), .Z(n5791) );
  XNOR U5679 ( .A(p_input[1834]), .B(n5790), .Z(n5792) );
  XOR U5680 ( .A(n5793), .B(n5794), .Z(n5790) );
  AND U5681 ( .A(n463), .B(n5795), .Z(n5794) );
  XNOR U5682 ( .A(p_input[1850]), .B(n5793), .Z(n5795) );
  XOR U5683 ( .A(n5796), .B(n5797), .Z(n5793) );
  AND U5684 ( .A(n467), .B(n5798), .Z(n5797) );
  XNOR U5685 ( .A(p_input[1866]), .B(n5796), .Z(n5798) );
  XOR U5686 ( .A(n5799), .B(n5800), .Z(n5796) );
  AND U5687 ( .A(n471), .B(n5801), .Z(n5800) );
  XNOR U5688 ( .A(p_input[1882]), .B(n5799), .Z(n5801) );
  XOR U5689 ( .A(n5802), .B(n5803), .Z(n5799) );
  AND U5690 ( .A(n475), .B(n5804), .Z(n5803) );
  XNOR U5691 ( .A(p_input[1898]), .B(n5802), .Z(n5804) );
  XOR U5692 ( .A(n5805), .B(n5806), .Z(n5802) );
  AND U5693 ( .A(n479), .B(n5807), .Z(n5806) );
  XNOR U5694 ( .A(p_input[1914]), .B(n5805), .Z(n5807) );
  XOR U5695 ( .A(n5808), .B(n5809), .Z(n5805) );
  AND U5696 ( .A(n483), .B(n5810), .Z(n5809) );
  XNOR U5697 ( .A(p_input[1930]), .B(n5808), .Z(n5810) );
  XOR U5698 ( .A(n5811), .B(n5812), .Z(n5808) );
  AND U5699 ( .A(n487), .B(n5813), .Z(n5812) );
  XNOR U5700 ( .A(p_input[1946]), .B(n5811), .Z(n5813) );
  XOR U5701 ( .A(n5814), .B(n5815), .Z(n5811) );
  AND U5702 ( .A(n491), .B(n5816), .Z(n5815) );
  XNOR U5703 ( .A(p_input[1962]), .B(n5814), .Z(n5816) );
  XOR U5704 ( .A(n5817), .B(n5818), .Z(n5814) );
  AND U5705 ( .A(n495), .B(n5819), .Z(n5818) );
  XNOR U5706 ( .A(p_input[1978]), .B(n5817), .Z(n5819) );
  XOR U5707 ( .A(n5820), .B(n5821), .Z(n5817) );
  AND U5708 ( .A(n499), .B(n5822), .Z(n5821) );
  XNOR U5709 ( .A(p_input[1994]), .B(n5820), .Z(n5822) );
  XNOR U5710 ( .A(n5823), .B(n5824), .Z(n5820) );
  AND U5711 ( .A(n503), .B(n5825), .Z(n5824) );
  XOR U5712 ( .A(p_input[2010]), .B(n5823), .Z(n5825) );
  XOR U5713 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n5826), .Z(n5823) );
  AND U5714 ( .A(n506), .B(n5827), .Z(n5826) );
  XOR U5715 ( .A(p_input[2026]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n5827)
         );
  XNOR U5716 ( .A(n5828), .B(n5829), .Z(o[0]) );
  AND U5717 ( .A(n3), .B(n5830), .Z(n5828) );
  XNOR U5718 ( .A(p_input[0]), .B(n5829), .Z(n5830) );
  XOR U5719 ( .A(n5831), .B(n5832), .Z(n5829) );
  AND U5720 ( .A(n7), .B(n5833), .Z(n5832) );
  XNOR U5721 ( .A(p_input[16]), .B(n5831), .Z(n5833) );
  XOR U5722 ( .A(n5834), .B(n5835), .Z(n5831) );
  AND U5723 ( .A(n11), .B(n5836), .Z(n5835) );
  XNOR U5724 ( .A(p_input[32]), .B(n5834), .Z(n5836) );
  XOR U5725 ( .A(n5837), .B(n5838), .Z(n5834) );
  AND U5726 ( .A(n15), .B(n5839), .Z(n5838) );
  XNOR U5727 ( .A(p_input[48]), .B(n5837), .Z(n5839) );
  XOR U5728 ( .A(n5840), .B(n5841), .Z(n5837) );
  AND U5729 ( .A(n19), .B(n5842), .Z(n5841) );
  XNOR U5730 ( .A(p_input[64]), .B(n5840), .Z(n5842) );
  XOR U5731 ( .A(n5843), .B(n5844), .Z(n5840) );
  AND U5732 ( .A(n23), .B(n5845), .Z(n5844) );
  XNOR U5733 ( .A(p_input[80]), .B(n5843), .Z(n5845) );
  XOR U5734 ( .A(n5846), .B(n5847), .Z(n5843) );
  AND U5735 ( .A(n27), .B(n5848), .Z(n5847) );
  XNOR U5736 ( .A(p_input[96]), .B(n5846), .Z(n5848) );
  XOR U5737 ( .A(n5849), .B(n5850), .Z(n5846) );
  AND U5738 ( .A(n31), .B(n5851), .Z(n5850) );
  XNOR U5739 ( .A(p_input[112]), .B(n5849), .Z(n5851) );
  XOR U5740 ( .A(n5852), .B(n5853), .Z(n5849) );
  AND U5741 ( .A(n35), .B(n5854), .Z(n5853) );
  XNOR U5742 ( .A(p_input[128]), .B(n5852), .Z(n5854) );
  XOR U5743 ( .A(n5855), .B(n5856), .Z(n5852) );
  AND U5744 ( .A(n39), .B(n5857), .Z(n5856) );
  XNOR U5745 ( .A(p_input[144]), .B(n5855), .Z(n5857) );
  XOR U5746 ( .A(n5858), .B(n5859), .Z(n5855) );
  AND U5747 ( .A(n43), .B(n5860), .Z(n5859) );
  XNOR U5748 ( .A(p_input[160]), .B(n5858), .Z(n5860) );
  XOR U5749 ( .A(n5861), .B(n5862), .Z(n5858) );
  AND U5750 ( .A(n47), .B(n5863), .Z(n5862) );
  XNOR U5751 ( .A(p_input[176]), .B(n5861), .Z(n5863) );
  XOR U5752 ( .A(n5864), .B(n5865), .Z(n5861) );
  AND U5753 ( .A(n51), .B(n5866), .Z(n5865) );
  XNOR U5754 ( .A(p_input[192]), .B(n5864), .Z(n5866) );
  XOR U5755 ( .A(n5867), .B(n5868), .Z(n5864) );
  AND U5756 ( .A(n55), .B(n5869), .Z(n5868) );
  XNOR U5757 ( .A(p_input[208]), .B(n5867), .Z(n5869) );
  XOR U5758 ( .A(n5870), .B(n5871), .Z(n5867) );
  AND U5759 ( .A(n59), .B(n5872), .Z(n5871) );
  XNOR U5760 ( .A(p_input[224]), .B(n5870), .Z(n5872) );
  XOR U5761 ( .A(n5873), .B(n5874), .Z(n5870) );
  AND U5762 ( .A(n63), .B(n5875), .Z(n5874) );
  XNOR U5763 ( .A(p_input[240]), .B(n5873), .Z(n5875) );
  XOR U5764 ( .A(n5876), .B(n5877), .Z(n5873) );
  AND U5765 ( .A(n67), .B(n5878), .Z(n5877) );
  XNOR U5766 ( .A(p_input[256]), .B(n5876), .Z(n5878) );
  XOR U5767 ( .A(n5879), .B(n5880), .Z(n5876) );
  AND U5768 ( .A(n71), .B(n5881), .Z(n5880) );
  XNOR U5769 ( .A(p_input[272]), .B(n5879), .Z(n5881) );
  XOR U5770 ( .A(n5882), .B(n5883), .Z(n5879) );
  AND U5771 ( .A(n75), .B(n5884), .Z(n5883) );
  XNOR U5772 ( .A(p_input[288]), .B(n5882), .Z(n5884) );
  XOR U5773 ( .A(n5885), .B(n5886), .Z(n5882) );
  AND U5774 ( .A(n79), .B(n5887), .Z(n5886) );
  XNOR U5775 ( .A(p_input[304]), .B(n5885), .Z(n5887) );
  XOR U5776 ( .A(n5888), .B(n5889), .Z(n5885) );
  AND U5777 ( .A(n83), .B(n5890), .Z(n5889) );
  XNOR U5778 ( .A(p_input[320]), .B(n5888), .Z(n5890) );
  XOR U5779 ( .A(n5891), .B(n5892), .Z(n5888) );
  AND U5780 ( .A(n87), .B(n5893), .Z(n5892) );
  XNOR U5781 ( .A(p_input[336]), .B(n5891), .Z(n5893) );
  XOR U5782 ( .A(n5894), .B(n5895), .Z(n5891) );
  AND U5783 ( .A(n91), .B(n5896), .Z(n5895) );
  XNOR U5784 ( .A(p_input[352]), .B(n5894), .Z(n5896) );
  XOR U5785 ( .A(n5897), .B(n5898), .Z(n5894) );
  AND U5786 ( .A(n95), .B(n5899), .Z(n5898) );
  XNOR U5787 ( .A(p_input[368]), .B(n5897), .Z(n5899) );
  XOR U5788 ( .A(n5900), .B(n5901), .Z(n5897) );
  AND U5789 ( .A(n99), .B(n5902), .Z(n5901) );
  XNOR U5790 ( .A(p_input[384]), .B(n5900), .Z(n5902) );
  XOR U5791 ( .A(n5903), .B(n5904), .Z(n5900) );
  AND U5792 ( .A(n103), .B(n5905), .Z(n5904) );
  XNOR U5793 ( .A(p_input[400]), .B(n5903), .Z(n5905) );
  XOR U5794 ( .A(n5906), .B(n5907), .Z(n5903) );
  AND U5795 ( .A(n107), .B(n5908), .Z(n5907) );
  XNOR U5796 ( .A(p_input[416]), .B(n5906), .Z(n5908) );
  XOR U5797 ( .A(n5909), .B(n5910), .Z(n5906) );
  AND U5798 ( .A(n111), .B(n5911), .Z(n5910) );
  XNOR U5799 ( .A(p_input[432]), .B(n5909), .Z(n5911) );
  XOR U5800 ( .A(n5912), .B(n5913), .Z(n5909) );
  AND U5801 ( .A(n115), .B(n5914), .Z(n5913) );
  XNOR U5802 ( .A(p_input[448]), .B(n5912), .Z(n5914) );
  XOR U5803 ( .A(n5915), .B(n5916), .Z(n5912) );
  AND U5804 ( .A(n119), .B(n5917), .Z(n5916) );
  XNOR U5805 ( .A(p_input[464]), .B(n5915), .Z(n5917) );
  XOR U5806 ( .A(n5918), .B(n5919), .Z(n5915) );
  AND U5807 ( .A(n123), .B(n5920), .Z(n5919) );
  XNOR U5808 ( .A(p_input[480]), .B(n5918), .Z(n5920) );
  XOR U5809 ( .A(n5921), .B(n5922), .Z(n5918) );
  AND U5810 ( .A(n127), .B(n5923), .Z(n5922) );
  XNOR U5811 ( .A(p_input[496]), .B(n5921), .Z(n5923) );
  XOR U5812 ( .A(n5924), .B(n5925), .Z(n5921) );
  AND U5813 ( .A(n131), .B(n5926), .Z(n5925) );
  XNOR U5814 ( .A(p_input[512]), .B(n5924), .Z(n5926) );
  XOR U5815 ( .A(n5927), .B(n5928), .Z(n5924) );
  AND U5816 ( .A(n135), .B(n5929), .Z(n5928) );
  XNOR U5817 ( .A(p_input[528]), .B(n5927), .Z(n5929) );
  XOR U5818 ( .A(n5930), .B(n5931), .Z(n5927) );
  AND U5819 ( .A(n139), .B(n5932), .Z(n5931) );
  XNOR U5820 ( .A(p_input[544]), .B(n5930), .Z(n5932) );
  XOR U5821 ( .A(n5933), .B(n5934), .Z(n5930) );
  AND U5822 ( .A(n143), .B(n5935), .Z(n5934) );
  XNOR U5823 ( .A(p_input[560]), .B(n5933), .Z(n5935) );
  XOR U5824 ( .A(n5936), .B(n5937), .Z(n5933) );
  AND U5825 ( .A(n147), .B(n5938), .Z(n5937) );
  XNOR U5826 ( .A(p_input[576]), .B(n5936), .Z(n5938) );
  XOR U5827 ( .A(n5939), .B(n5940), .Z(n5936) );
  AND U5828 ( .A(n151), .B(n5941), .Z(n5940) );
  XNOR U5829 ( .A(p_input[592]), .B(n5939), .Z(n5941) );
  XOR U5830 ( .A(n5942), .B(n5943), .Z(n5939) );
  AND U5831 ( .A(n155), .B(n5944), .Z(n5943) );
  XNOR U5832 ( .A(p_input[608]), .B(n5942), .Z(n5944) );
  XOR U5833 ( .A(n5945), .B(n5946), .Z(n5942) );
  AND U5834 ( .A(n159), .B(n5947), .Z(n5946) );
  XNOR U5835 ( .A(p_input[624]), .B(n5945), .Z(n5947) );
  XOR U5836 ( .A(n5948), .B(n5949), .Z(n5945) );
  AND U5837 ( .A(n163), .B(n5950), .Z(n5949) );
  XNOR U5838 ( .A(p_input[640]), .B(n5948), .Z(n5950) );
  XOR U5839 ( .A(n5951), .B(n5952), .Z(n5948) );
  AND U5840 ( .A(n167), .B(n5953), .Z(n5952) );
  XNOR U5841 ( .A(p_input[656]), .B(n5951), .Z(n5953) );
  XOR U5842 ( .A(n5954), .B(n5955), .Z(n5951) );
  AND U5843 ( .A(n171), .B(n5956), .Z(n5955) );
  XNOR U5844 ( .A(p_input[672]), .B(n5954), .Z(n5956) );
  XOR U5845 ( .A(n5957), .B(n5958), .Z(n5954) );
  AND U5846 ( .A(n175), .B(n5959), .Z(n5958) );
  XNOR U5847 ( .A(p_input[688]), .B(n5957), .Z(n5959) );
  XOR U5848 ( .A(n5960), .B(n5961), .Z(n5957) );
  AND U5849 ( .A(n179), .B(n5962), .Z(n5961) );
  XNOR U5850 ( .A(p_input[704]), .B(n5960), .Z(n5962) );
  XOR U5851 ( .A(n5963), .B(n5964), .Z(n5960) );
  AND U5852 ( .A(n183), .B(n5965), .Z(n5964) );
  XNOR U5853 ( .A(p_input[720]), .B(n5963), .Z(n5965) );
  XOR U5854 ( .A(n5966), .B(n5967), .Z(n5963) );
  AND U5855 ( .A(n187), .B(n5968), .Z(n5967) );
  XNOR U5856 ( .A(p_input[736]), .B(n5966), .Z(n5968) );
  XOR U5857 ( .A(n5969), .B(n5970), .Z(n5966) );
  AND U5858 ( .A(n191), .B(n5971), .Z(n5970) );
  XNOR U5859 ( .A(p_input[752]), .B(n5969), .Z(n5971) );
  XOR U5860 ( .A(n5972), .B(n5973), .Z(n5969) );
  AND U5861 ( .A(n195), .B(n5974), .Z(n5973) );
  XNOR U5862 ( .A(p_input[768]), .B(n5972), .Z(n5974) );
  XOR U5863 ( .A(n5975), .B(n5976), .Z(n5972) );
  AND U5864 ( .A(n199), .B(n5977), .Z(n5976) );
  XNOR U5865 ( .A(p_input[784]), .B(n5975), .Z(n5977) );
  XOR U5866 ( .A(n5978), .B(n5979), .Z(n5975) );
  AND U5867 ( .A(n203), .B(n5980), .Z(n5979) );
  XNOR U5868 ( .A(p_input[800]), .B(n5978), .Z(n5980) );
  XOR U5869 ( .A(n5981), .B(n5982), .Z(n5978) );
  AND U5870 ( .A(n207), .B(n5983), .Z(n5982) );
  XNOR U5871 ( .A(p_input[816]), .B(n5981), .Z(n5983) );
  XOR U5872 ( .A(n5984), .B(n5985), .Z(n5981) );
  AND U5873 ( .A(n211), .B(n5986), .Z(n5985) );
  XNOR U5874 ( .A(p_input[832]), .B(n5984), .Z(n5986) );
  XOR U5875 ( .A(n5987), .B(n5988), .Z(n5984) );
  AND U5876 ( .A(n215), .B(n5989), .Z(n5988) );
  XNOR U5877 ( .A(p_input[848]), .B(n5987), .Z(n5989) );
  XOR U5878 ( .A(n5990), .B(n5991), .Z(n5987) );
  AND U5879 ( .A(n219), .B(n5992), .Z(n5991) );
  XNOR U5880 ( .A(p_input[864]), .B(n5990), .Z(n5992) );
  XOR U5881 ( .A(n5993), .B(n5994), .Z(n5990) );
  AND U5882 ( .A(n223), .B(n5995), .Z(n5994) );
  XNOR U5883 ( .A(p_input[880]), .B(n5993), .Z(n5995) );
  XOR U5884 ( .A(n5996), .B(n5997), .Z(n5993) );
  AND U5885 ( .A(n227), .B(n5998), .Z(n5997) );
  XNOR U5886 ( .A(p_input[896]), .B(n5996), .Z(n5998) );
  XOR U5887 ( .A(n5999), .B(n6000), .Z(n5996) );
  AND U5888 ( .A(n231), .B(n6001), .Z(n6000) );
  XNOR U5889 ( .A(p_input[912]), .B(n5999), .Z(n6001) );
  XOR U5890 ( .A(n6002), .B(n6003), .Z(n5999) );
  AND U5891 ( .A(n235), .B(n6004), .Z(n6003) );
  XNOR U5892 ( .A(p_input[928]), .B(n6002), .Z(n6004) );
  XOR U5893 ( .A(n6005), .B(n6006), .Z(n6002) );
  AND U5894 ( .A(n239), .B(n6007), .Z(n6006) );
  XNOR U5895 ( .A(p_input[944]), .B(n6005), .Z(n6007) );
  XOR U5896 ( .A(n6008), .B(n6009), .Z(n6005) );
  AND U5897 ( .A(n243), .B(n6010), .Z(n6009) );
  XNOR U5898 ( .A(p_input[960]), .B(n6008), .Z(n6010) );
  XOR U5899 ( .A(n6011), .B(n6012), .Z(n6008) );
  AND U5900 ( .A(n247), .B(n6013), .Z(n6012) );
  XNOR U5901 ( .A(p_input[976]), .B(n6011), .Z(n6013) );
  XOR U5902 ( .A(n6014), .B(n6015), .Z(n6011) );
  AND U5903 ( .A(n251), .B(n6016), .Z(n6015) );
  XNOR U5904 ( .A(p_input[992]), .B(n6014), .Z(n6016) );
  XOR U5905 ( .A(n6017), .B(n6018), .Z(n6014) );
  AND U5906 ( .A(n255), .B(n6019), .Z(n6018) );
  XNOR U5907 ( .A(p_input[1008]), .B(n6017), .Z(n6019) );
  XOR U5908 ( .A(n6020), .B(n6021), .Z(n6017) );
  AND U5909 ( .A(n259), .B(n6022), .Z(n6021) );
  XNOR U5910 ( .A(p_input[1024]), .B(n6020), .Z(n6022) );
  XOR U5911 ( .A(n6023), .B(n6024), .Z(n6020) );
  AND U5912 ( .A(n263), .B(n6025), .Z(n6024) );
  XNOR U5913 ( .A(p_input[1040]), .B(n6023), .Z(n6025) );
  XOR U5914 ( .A(n6026), .B(n6027), .Z(n6023) );
  AND U5915 ( .A(n267), .B(n6028), .Z(n6027) );
  XNOR U5916 ( .A(p_input[1056]), .B(n6026), .Z(n6028) );
  XOR U5917 ( .A(n6029), .B(n6030), .Z(n6026) );
  AND U5918 ( .A(n271), .B(n6031), .Z(n6030) );
  XNOR U5919 ( .A(p_input[1072]), .B(n6029), .Z(n6031) );
  XOR U5920 ( .A(n6032), .B(n6033), .Z(n6029) );
  AND U5921 ( .A(n275), .B(n6034), .Z(n6033) );
  XNOR U5922 ( .A(p_input[1088]), .B(n6032), .Z(n6034) );
  XOR U5923 ( .A(n6035), .B(n6036), .Z(n6032) );
  AND U5924 ( .A(n279), .B(n6037), .Z(n6036) );
  XNOR U5925 ( .A(p_input[1104]), .B(n6035), .Z(n6037) );
  XOR U5926 ( .A(n6038), .B(n6039), .Z(n6035) );
  AND U5927 ( .A(n283), .B(n6040), .Z(n6039) );
  XNOR U5928 ( .A(p_input[1120]), .B(n6038), .Z(n6040) );
  XOR U5929 ( .A(n6041), .B(n6042), .Z(n6038) );
  AND U5930 ( .A(n287), .B(n6043), .Z(n6042) );
  XNOR U5931 ( .A(p_input[1136]), .B(n6041), .Z(n6043) );
  XOR U5932 ( .A(n6044), .B(n6045), .Z(n6041) );
  AND U5933 ( .A(n291), .B(n6046), .Z(n6045) );
  XNOR U5934 ( .A(p_input[1152]), .B(n6044), .Z(n6046) );
  XOR U5935 ( .A(n6047), .B(n6048), .Z(n6044) );
  AND U5936 ( .A(n295), .B(n6049), .Z(n6048) );
  XNOR U5937 ( .A(p_input[1168]), .B(n6047), .Z(n6049) );
  XOR U5938 ( .A(n6050), .B(n6051), .Z(n6047) );
  AND U5939 ( .A(n299), .B(n6052), .Z(n6051) );
  XNOR U5940 ( .A(p_input[1184]), .B(n6050), .Z(n6052) );
  XOR U5941 ( .A(n6053), .B(n6054), .Z(n6050) );
  AND U5942 ( .A(n303), .B(n6055), .Z(n6054) );
  XNOR U5943 ( .A(p_input[1200]), .B(n6053), .Z(n6055) );
  XOR U5944 ( .A(n6056), .B(n6057), .Z(n6053) );
  AND U5945 ( .A(n307), .B(n6058), .Z(n6057) );
  XNOR U5946 ( .A(p_input[1216]), .B(n6056), .Z(n6058) );
  XOR U5947 ( .A(n6059), .B(n6060), .Z(n6056) );
  AND U5948 ( .A(n311), .B(n6061), .Z(n6060) );
  XNOR U5949 ( .A(p_input[1232]), .B(n6059), .Z(n6061) );
  XOR U5950 ( .A(n6062), .B(n6063), .Z(n6059) );
  AND U5951 ( .A(n315), .B(n6064), .Z(n6063) );
  XNOR U5952 ( .A(p_input[1248]), .B(n6062), .Z(n6064) );
  XOR U5953 ( .A(n6065), .B(n6066), .Z(n6062) );
  AND U5954 ( .A(n319), .B(n6067), .Z(n6066) );
  XNOR U5955 ( .A(p_input[1264]), .B(n6065), .Z(n6067) );
  XOR U5956 ( .A(n6068), .B(n6069), .Z(n6065) );
  AND U5957 ( .A(n323), .B(n6070), .Z(n6069) );
  XNOR U5958 ( .A(p_input[1280]), .B(n6068), .Z(n6070) );
  XOR U5959 ( .A(n6071), .B(n6072), .Z(n6068) );
  AND U5960 ( .A(n327), .B(n6073), .Z(n6072) );
  XNOR U5961 ( .A(p_input[1296]), .B(n6071), .Z(n6073) );
  XOR U5962 ( .A(n6074), .B(n6075), .Z(n6071) );
  AND U5963 ( .A(n331), .B(n6076), .Z(n6075) );
  XNOR U5964 ( .A(p_input[1312]), .B(n6074), .Z(n6076) );
  XOR U5965 ( .A(n6077), .B(n6078), .Z(n6074) );
  AND U5966 ( .A(n335), .B(n6079), .Z(n6078) );
  XNOR U5967 ( .A(p_input[1328]), .B(n6077), .Z(n6079) );
  XOR U5968 ( .A(n6080), .B(n6081), .Z(n6077) );
  AND U5969 ( .A(n339), .B(n6082), .Z(n6081) );
  XNOR U5970 ( .A(p_input[1344]), .B(n6080), .Z(n6082) );
  XOR U5971 ( .A(n6083), .B(n6084), .Z(n6080) );
  AND U5972 ( .A(n343), .B(n6085), .Z(n6084) );
  XNOR U5973 ( .A(p_input[1360]), .B(n6083), .Z(n6085) );
  XOR U5974 ( .A(n6086), .B(n6087), .Z(n6083) );
  AND U5975 ( .A(n347), .B(n6088), .Z(n6087) );
  XNOR U5976 ( .A(p_input[1376]), .B(n6086), .Z(n6088) );
  XOR U5977 ( .A(n6089), .B(n6090), .Z(n6086) );
  AND U5978 ( .A(n351), .B(n6091), .Z(n6090) );
  XNOR U5979 ( .A(p_input[1392]), .B(n6089), .Z(n6091) );
  XOR U5980 ( .A(n6092), .B(n6093), .Z(n6089) );
  AND U5981 ( .A(n355), .B(n6094), .Z(n6093) );
  XNOR U5982 ( .A(p_input[1408]), .B(n6092), .Z(n6094) );
  XOR U5983 ( .A(n6095), .B(n6096), .Z(n6092) );
  AND U5984 ( .A(n359), .B(n6097), .Z(n6096) );
  XNOR U5985 ( .A(p_input[1424]), .B(n6095), .Z(n6097) );
  XOR U5986 ( .A(n6098), .B(n6099), .Z(n6095) );
  AND U5987 ( .A(n363), .B(n6100), .Z(n6099) );
  XNOR U5988 ( .A(p_input[1440]), .B(n6098), .Z(n6100) );
  XOR U5989 ( .A(n6101), .B(n6102), .Z(n6098) );
  AND U5990 ( .A(n367), .B(n6103), .Z(n6102) );
  XNOR U5991 ( .A(p_input[1456]), .B(n6101), .Z(n6103) );
  XOR U5992 ( .A(n6104), .B(n6105), .Z(n6101) );
  AND U5993 ( .A(n371), .B(n6106), .Z(n6105) );
  XNOR U5994 ( .A(p_input[1472]), .B(n6104), .Z(n6106) );
  XOR U5995 ( .A(n6107), .B(n6108), .Z(n6104) );
  AND U5996 ( .A(n375), .B(n6109), .Z(n6108) );
  XNOR U5997 ( .A(p_input[1488]), .B(n6107), .Z(n6109) );
  XOR U5998 ( .A(n6110), .B(n6111), .Z(n6107) );
  AND U5999 ( .A(n379), .B(n6112), .Z(n6111) );
  XNOR U6000 ( .A(p_input[1504]), .B(n6110), .Z(n6112) );
  XOR U6001 ( .A(n6113), .B(n6114), .Z(n6110) );
  AND U6002 ( .A(n383), .B(n6115), .Z(n6114) );
  XNOR U6003 ( .A(p_input[1520]), .B(n6113), .Z(n6115) );
  XOR U6004 ( .A(n6116), .B(n6117), .Z(n6113) );
  AND U6005 ( .A(n387), .B(n6118), .Z(n6117) );
  XNOR U6006 ( .A(p_input[1536]), .B(n6116), .Z(n6118) );
  XOR U6007 ( .A(n6119), .B(n6120), .Z(n6116) );
  AND U6008 ( .A(n391), .B(n6121), .Z(n6120) );
  XNOR U6009 ( .A(p_input[1552]), .B(n6119), .Z(n6121) );
  XOR U6010 ( .A(n6122), .B(n6123), .Z(n6119) );
  AND U6011 ( .A(n395), .B(n6124), .Z(n6123) );
  XNOR U6012 ( .A(p_input[1568]), .B(n6122), .Z(n6124) );
  XOR U6013 ( .A(n6125), .B(n6126), .Z(n6122) );
  AND U6014 ( .A(n399), .B(n6127), .Z(n6126) );
  XNOR U6015 ( .A(p_input[1584]), .B(n6125), .Z(n6127) );
  XOR U6016 ( .A(n6128), .B(n6129), .Z(n6125) );
  AND U6017 ( .A(n403), .B(n6130), .Z(n6129) );
  XNOR U6018 ( .A(p_input[1600]), .B(n6128), .Z(n6130) );
  XOR U6019 ( .A(n6131), .B(n6132), .Z(n6128) );
  AND U6020 ( .A(n407), .B(n6133), .Z(n6132) );
  XNOR U6021 ( .A(p_input[1616]), .B(n6131), .Z(n6133) );
  XOR U6022 ( .A(n6134), .B(n6135), .Z(n6131) );
  AND U6023 ( .A(n411), .B(n6136), .Z(n6135) );
  XNOR U6024 ( .A(p_input[1632]), .B(n6134), .Z(n6136) );
  XOR U6025 ( .A(n6137), .B(n6138), .Z(n6134) );
  AND U6026 ( .A(n415), .B(n6139), .Z(n6138) );
  XNOR U6027 ( .A(p_input[1648]), .B(n6137), .Z(n6139) );
  XOR U6028 ( .A(n6140), .B(n6141), .Z(n6137) );
  AND U6029 ( .A(n419), .B(n6142), .Z(n6141) );
  XNOR U6030 ( .A(p_input[1664]), .B(n6140), .Z(n6142) );
  XOR U6031 ( .A(n6143), .B(n6144), .Z(n6140) );
  AND U6032 ( .A(n423), .B(n6145), .Z(n6144) );
  XNOR U6033 ( .A(p_input[1680]), .B(n6143), .Z(n6145) );
  XOR U6034 ( .A(n6146), .B(n6147), .Z(n6143) );
  AND U6035 ( .A(n427), .B(n6148), .Z(n6147) );
  XNOR U6036 ( .A(p_input[1696]), .B(n6146), .Z(n6148) );
  XOR U6037 ( .A(n6149), .B(n6150), .Z(n6146) );
  AND U6038 ( .A(n431), .B(n6151), .Z(n6150) );
  XNOR U6039 ( .A(p_input[1712]), .B(n6149), .Z(n6151) );
  XOR U6040 ( .A(n6152), .B(n6153), .Z(n6149) );
  AND U6041 ( .A(n435), .B(n6154), .Z(n6153) );
  XNOR U6042 ( .A(p_input[1728]), .B(n6152), .Z(n6154) );
  XOR U6043 ( .A(n6155), .B(n6156), .Z(n6152) );
  AND U6044 ( .A(n439), .B(n6157), .Z(n6156) );
  XNOR U6045 ( .A(p_input[1744]), .B(n6155), .Z(n6157) );
  XOR U6046 ( .A(n6158), .B(n6159), .Z(n6155) );
  AND U6047 ( .A(n443), .B(n6160), .Z(n6159) );
  XNOR U6048 ( .A(p_input[1760]), .B(n6158), .Z(n6160) );
  XOR U6049 ( .A(n6161), .B(n6162), .Z(n6158) );
  AND U6050 ( .A(n447), .B(n6163), .Z(n6162) );
  XNOR U6051 ( .A(p_input[1776]), .B(n6161), .Z(n6163) );
  XOR U6052 ( .A(n6164), .B(n6165), .Z(n6161) );
  AND U6053 ( .A(n451), .B(n6166), .Z(n6165) );
  XNOR U6054 ( .A(p_input[1792]), .B(n6164), .Z(n6166) );
  XOR U6055 ( .A(n6167), .B(n6168), .Z(n6164) );
  AND U6056 ( .A(n455), .B(n6169), .Z(n6168) );
  XNOR U6057 ( .A(p_input[1808]), .B(n6167), .Z(n6169) );
  XOR U6058 ( .A(n6170), .B(n6171), .Z(n6167) );
  AND U6059 ( .A(n459), .B(n6172), .Z(n6171) );
  XNOR U6060 ( .A(p_input[1824]), .B(n6170), .Z(n6172) );
  XOR U6061 ( .A(n6173), .B(n6174), .Z(n6170) );
  AND U6062 ( .A(n463), .B(n6175), .Z(n6174) );
  XNOR U6063 ( .A(p_input[1840]), .B(n6173), .Z(n6175) );
  XOR U6064 ( .A(n6176), .B(n6177), .Z(n6173) );
  AND U6065 ( .A(n467), .B(n6178), .Z(n6177) );
  XNOR U6066 ( .A(p_input[1856]), .B(n6176), .Z(n6178) );
  XOR U6067 ( .A(n6179), .B(n6180), .Z(n6176) );
  AND U6068 ( .A(n471), .B(n6181), .Z(n6180) );
  XNOR U6069 ( .A(p_input[1872]), .B(n6179), .Z(n6181) );
  XOR U6070 ( .A(n6182), .B(n6183), .Z(n6179) );
  AND U6071 ( .A(n475), .B(n6184), .Z(n6183) );
  XNOR U6072 ( .A(p_input[1888]), .B(n6182), .Z(n6184) );
  XOR U6073 ( .A(n6185), .B(n6186), .Z(n6182) );
  AND U6074 ( .A(n479), .B(n6187), .Z(n6186) );
  XNOR U6075 ( .A(p_input[1904]), .B(n6185), .Z(n6187) );
  XOR U6076 ( .A(n6188), .B(n6189), .Z(n6185) );
  AND U6077 ( .A(n483), .B(n6190), .Z(n6189) );
  XNOR U6078 ( .A(p_input[1920]), .B(n6188), .Z(n6190) );
  XOR U6079 ( .A(n6191), .B(n6192), .Z(n6188) );
  AND U6080 ( .A(n487), .B(n6193), .Z(n6192) );
  XNOR U6081 ( .A(p_input[1936]), .B(n6191), .Z(n6193) );
  XOR U6082 ( .A(n6194), .B(n6195), .Z(n6191) );
  AND U6083 ( .A(n491), .B(n6196), .Z(n6195) );
  XNOR U6084 ( .A(p_input[1952]), .B(n6194), .Z(n6196) );
  XOR U6085 ( .A(n6197), .B(n6198), .Z(n6194) );
  AND U6086 ( .A(n495), .B(n6199), .Z(n6198) );
  XNOR U6087 ( .A(p_input[1968]), .B(n6197), .Z(n6199) );
  XOR U6088 ( .A(n6200), .B(n6201), .Z(n6197) );
  AND U6089 ( .A(n499), .B(n6202), .Z(n6201) );
  XNOR U6090 ( .A(p_input[1984]), .B(n6200), .Z(n6202) );
  XNOR U6091 ( .A(n6203), .B(n6204), .Z(n6200) );
  AND U6092 ( .A(n503), .B(n6205), .Z(n6204) );
  XOR U6093 ( .A(p_input[2000]), .B(n6203), .Z(n6205) );
  XOR U6094 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n6206), .Z(n6203) );
  AND U6095 ( .A(n506), .B(n6207), .Z(n6206) );
  XOR U6096 ( .A(p_input[2016]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n6207)
         );
  XNOR U6097 ( .A(n6208), .B(n6209), .Z(n3) );
  AND U6098 ( .A(n6210), .B(n6211), .Z(n6209) );
  XOR U6099 ( .A(n6212), .B(n6208), .Z(n6211) );
  AND U6100 ( .A(n6213), .B(n6214), .Z(n6212) );
  XOR U6101 ( .A(n6215), .B(n6208), .Z(n6210) );
  XNOR U6102 ( .A(n6216), .B(n6217), .Z(n6215) );
  AND U6103 ( .A(n7), .B(n6218), .Z(n6217) );
  XOR U6104 ( .A(n6219), .B(n6216), .Z(n6218) );
  XOR U6105 ( .A(n6220), .B(n6221), .Z(n6208) );
  AND U6106 ( .A(n6222), .B(n6223), .Z(n6221) );
  XNOR U6107 ( .A(n6220), .B(n6213), .Z(n6223) );
  XNOR U6108 ( .A(n6224), .B(n6225), .Z(n6213) );
  XOR U6109 ( .A(n6226), .B(n6214), .Z(n6225) );
  AND U6110 ( .A(n6227), .B(n6228), .Z(n6214) );
  AND U6111 ( .A(n6229), .B(n6230), .Z(n6226) );
  XOR U6112 ( .A(n6231), .B(n6224), .Z(n6229) );
  XOR U6113 ( .A(n6232), .B(n6220), .Z(n6222) );
  XNOR U6114 ( .A(n6233), .B(n6234), .Z(n6232) );
  AND U6115 ( .A(n7), .B(n6235), .Z(n6234) );
  XOR U6116 ( .A(n6236), .B(n6233), .Z(n6235) );
  XOR U6117 ( .A(n6237), .B(n6238), .Z(n6220) );
  AND U6118 ( .A(n6239), .B(n6240), .Z(n6238) );
  XNOR U6119 ( .A(n6237), .B(n6227), .Z(n6240) );
  XOR U6120 ( .A(n6241), .B(n6230), .Z(n6227) );
  XNOR U6121 ( .A(n6242), .B(n6224), .Z(n6230) );
  XOR U6122 ( .A(n6243), .B(n6244), .Z(n6224) );
  AND U6123 ( .A(n6245), .B(n6246), .Z(n6244) );
  XOR U6124 ( .A(n6247), .B(n6243), .Z(n6245) );
  XNOR U6125 ( .A(n6248), .B(n6249), .Z(n6242) );
  AND U6126 ( .A(n6250), .B(n6251), .Z(n6249) );
  XOR U6127 ( .A(n6248), .B(n6252), .Z(n6250) );
  XNOR U6128 ( .A(n6231), .B(n6228), .Z(n6241) );
  AND U6129 ( .A(n6253), .B(n6254), .Z(n6228) );
  XOR U6130 ( .A(n6255), .B(n6256), .Z(n6231) );
  AND U6131 ( .A(n6257), .B(n6258), .Z(n6256) );
  XOR U6132 ( .A(n6255), .B(n6259), .Z(n6257) );
  XOR U6133 ( .A(n6260), .B(n6237), .Z(n6239) );
  XNOR U6134 ( .A(n6261), .B(n6262), .Z(n6260) );
  AND U6135 ( .A(n7), .B(n6263), .Z(n6262) );
  XNOR U6136 ( .A(n6264), .B(n6261), .Z(n6263) );
  XOR U6137 ( .A(n6265), .B(n6266), .Z(n6237) );
  AND U6138 ( .A(n6267), .B(n6268), .Z(n6266) );
  XNOR U6139 ( .A(n6265), .B(n6253), .Z(n6268) );
  XOR U6140 ( .A(n6269), .B(n6246), .Z(n6253) );
  XNOR U6141 ( .A(n6270), .B(n6252), .Z(n6246) );
  XNOR U6142 ( .A(n6271), .B(n6272), .Z(n6252) );
  NOR U6143 ( .A(n6273), .B(n6274), .Z(n6272) );
  XOR U6144 ( .A(n6271), .B(n6275), .Z(n6273) );
  XNOR U6145 ( .A(n6251), .B(n6243), .Z(n6270) );
  XOR U6146 ( .A(n6276), .B(n6277), .Z(n6243) );
  AND U6147 ( .A(n6278), .B(n6279), .Z(n6277) );
  XNOR U6148 ( .A(n6276), .B(n6280), .Z(n6278) );
  XNOR U6149 ( .A(n6281), .B(n6248), .Z(n6251) );
  XOR U6150 ( .A(n6282), .B(n6283), .Z(n6248) );
  AND U6151 ( .A(n6284), .B(n6285), .Z(n6283) );
  XOR U6152 ( .A(n6282), .B(n6286), .Z(n6284) );
  XNOR U6153 ( .A(n6287), .B(n6288), .Z(n6281) );
  NOR U6154 ( .A(n6289), .B(n6290), .Z(n6288) );
  XNOR U6155 ( .A(n6287), .B(n6291), .Z(n6289) );
  XNOR U6156 ( .A(n6247), .B(n6254), .Z(n6269) );
  NOR U6157 ( .A(n6292), .B(n6293), .Z(n6254) );
  XOR U6158 ( .A(n6259), .B(n6258), .Z(n6247) );
  XNOR U6159 ( .A(n6294), .B(n6255), .Z(n6258) );
  XOR U6160 ( .A(n6295), .B(n6296), .Z(n6255) );
  AND U6161 ( .A(n6297), .B(n6298), .Z(n6296) );
  XOR U6162 ( .A(n6295), .B(n6299), .Z(n6297) );
  XNOR U6163 ( .A(n6300), .B(n6301), .Z(n6294) );
  NOR U6164 ( .A(n6302), .B(n6303), .Z(n6301) );
  XNOR U6165 ( .A(n6300), .B(n6304), .Z(n6302) );
  XOR U6166 ( .A(n6305), .B(n6306), .Z(n6259) );
  NOR U6167 ( .A(n6307), .B(n6308), .Z(n6306) );
  XNOR U6168 ( .A(n6305), .B(n6309), .Z(n6307) );
  XNOR U6169 ( .A(n6310), .B(n6311), .Z(n6267) );
  XOR U6170 ( .A(n6265), .B(n6312), .Z(n6311) );
  AND U6171 ( .A(n7), .B(n6313), .Z(n6312) );
  XOR U6172 ( .A(n6314), .B(n6310), .Z(n6313) );
  AND U6173 ( .A(n6315), .B(n6292), .Z(n6265) );
  XOR U6174 ( .A(n6316), .B(n6293), .Z(n6292) );
  XNOR U6175 ( .A(p_input[0]), .B(p_input[2048]), .Z(n6293) );
  XOR U6176 ( .A(n6280), .B(n6279), .Z(n6316) );
  XNOR U6177 ( .A(n6317), .B(n6286), .Z(n6279) );
  XNOR U6178 ( .A(n6275), .B(n6274), .Z(n6286) );
  XNOR U6179 ( .A(n6318), .B(n6271), .Z(n6274) );
  XNOR U6180 ( .A(p_input[10]), .B(p_input[2058]), .Z(n6271) );
  XOR U6181 ( .A(p_input[11]), .B(n6319), .Z(n6318) );
  XOR U6182 ( .A(p_input[12]), .B(p_input[2060]), .Z(n6275) );
  XOR U6183 ( .A(n6285), .B(n6320), .Z(n6317) );
  IV U6184 ( .A(n6276), .Z(n6320) );
  XOR U6185 ( .A(p_input[1]), .B(p_input[2049]), .Z(n6276) );
  XNOR U6186 ( .A(n6321), .B(n6291), .Z(n6285) );
  XNOR U6187 ( .A(p_input[15]), .B(n6322), .Z(n6291) );
  XOR U6188 ( .A(n6282), .B(n6290), .Z(n6321) );
  XOR U6189 ( .A(n6323), .B(n6287), .Z(n6290) );
  XOR U6190 ( .A(p_input[13]), .B(p_input[2061]), .Z(n6287) );
  XOR U6191 ( .A(p_input[14]), .B(n6324), .Z(n6323) );
  XNOR U6192 ( .A(n6325), .B(p_input[9]), .Z(n6282) );
  XNOR U6193 ( .A(n6299), .B(n6298), .Z(n6280) );
  XNOR U6194 ( .A(n6326), .B(n6304), .Z(n6298) );
  XOR U6195 ( .A(p_input[2056]), .B(p_input[8]), .Z(n6304) );
  XOR U6196 ( .A(n6295), .B(n6303), .Z(n6326) );
  XOR U6197 ( .A(n6327), .B(n6300), .Z(n6303) );
  XOR U6198 ( .A(p_input[2054]), .B(p_input[6]), .Z(n6300) );
  XNOR U6199 ( .A(p_input[2055]), .B(p_input[7]), .Z(n6327) );
  XNOR U6200 ( .A(n6328), .B(p_input[2]), .Z(n6295) );
  XNOR U6201 ( .A(n6309), .B(n6308), .Z(n6299) );
  XOR U6202 ( .A(n6329), .B(n6305), .Z(n6308) );
  XOR U6203 ( .A(p_input[2051]), .B(p_input[3]), .Z(n6305) );
  XNOR U6204 ( .A(p_input[2052]), .B(p_input[4]), .Z(n6329) );
  XOR U6205 ( .A(p_input[2053]), .B(p_input[5]), .Z(n6309) );
  XNOR U6206 ( .A(n6330), .B(n6331), .Z(n6315) );
  AND U6207 ( .A(n7), .B(n6332), .Z(n6331) );
  XNOR U6208 ( .A(n6333), .B(n6334), .Z(n6332) );
  XNOR U6209 ( .A(n6335), .B(n6336), .Z(n7) );
  AND U6210 ( .A(n6337), .B(n6338), .Z(n6336) );
  XOR U6211 ( .A(n6219), .B(n6335), .Z(n6338) );
  AND U6212 ( .A(n6339), .B(n6340), .Z(n6219) );
  XNOR U6213 ( .A(n6216), .B(n6335), .Z(n6337) );
  XOR U6214 ( .A(n6341), .B(n6342), .Z(n6216) );
  AND U6215 ( .A(n11), .B(n6343), .Z(n6342) );
  XOR U6216 ( .A(n6344), .B(n6341), .Z(n6343) );
  XOR U6217 ( .A(n6345), .B(n6346), .Z(n6335) );
  AND U6218 ( .A(n6347), .B(n6348), .Z(n6346) );
  XNOR U6219 ( .A(n6345), .B(n6339), .Z(n6348) );
  IV U6220 ( .A(n6236), .Z(n6339) );
  XOR U6221 ( .A(n6349), .B(n6350), .Z(n6236) );
  XOR U6222 ( .A(n6351), .B(n6340), .Z(n6350) );
  AND U6223 ( .A(n6264), .B(n6352), .Z(n6340) );
  AND U6224 ( .A(n6353), .B(n6354), .Z(n6351) );
  XOR U6225 ( .A(n6355), .B(n6349), .Z(n6353) );
  XNOR U6226 ( .A(n6233), .B(n6345), .Z(n6347) );
  XOR U6227 ( .A(n6356), .B(n6357), .Z(n6233) );
  AND U6228 ( .A(n11), .B(n6358), .Z(n6357) );
  XOR U6229 ( .A(n6359), .B(n6356), .Z(n6358) );
  XOR U6230 ( .A(n6360), .B(n6361), .Z(n6345) );
  AND U6231 ( .A(n6362), .B(n6363), .Z(n6361) );
  XNOR U6232 ( .A(n6360), .B(n6264), .Z(n6363) );
  XOR U6233 ( .A(n6364), .B(n6354), .Z(n6264) );
  XNOR U6234 ( .A(n6365), .B(n6349), .Z(n6354) );
  XOR U6235 ( .A(n6366), .B(n6367), .Z(n6349) );
  AND U6236 ( .A(n6368), .B(n6369), .Z(n6367) );
  XOR U6237 ( .A(n6370), .B(n6366), .Z(n6368) );
  XNOR U6238 ( .A(n6371), .B(n6372), .Z(n6365) );
  AND U6239 ( .A(n6373), .B(n6374), .Z(n6372) );
  XOR U6240 ( .A(n6371), .B(n6375), .Z(n6373) );
  XNOR U6241 ( .A(n6355), .B(n6352), .Z(n6364) );
  AND U6242 ( .A(n6376), .B(n6377), .Z(n6352) );
  XOR U6243 ( .A(n6378), .B(n6379), .Z(n6355) );
  AND U6244 ( .A(n6380), .B(n6381), .Z(n6379) );
  XOR U6245 ( .A(n6378), .B(n6382), .Z(n6380) );
  XNOR U6246 ( .A(n6261), .B(n6360), .Z(n6362) );
  XOR U6247 ( .A(n6383), .B(n6384), .Z(n6261) );
  AND U6248 ( .A(n11), .B(n6385), .Z(n6384) );
  XNOR U6249 ( .A(n6386), .B(n6383), .Z(n6385) );
  XOR U6250 ( .A(n6387), .B(n6388), .Z(n6360) );
  AND U6251 ( .A(n6389), .B(n6390), .Z(n6388) );
  XNOR U6252 ( .A(n6387), .B(n6376), .Z(n6390) );
  IV U6253 ( .A(n6314), .Z(n6376) );
  XNOR U6254 ( .A(n6391), .B(n6369), .Z(n6314) );
  XNOR U6255 ( .A(n6392), .B(n6375), .Z(n6369) );
  XOR U6256 ( .A(n6393), .B(n6394), .Z(n6375) );
  NOR U6257 ( .A(n6395), .B(n6396), .Z(n6394) );
  XNOR U6258 ( .A(n6393), .B(n6397), .Z(n6395) );
  XNOR U6259 ( .A(n6374), .B(n6366), .Z(n6392) );
  XOR U6260 ( .A(n6398), .B(n6399), .Z(n6366) );
  AND U6261 ( .A(n6400), .B(n6401), .Z(n6399) );
  XNOR U6262 ( .A(n6398), .B(n6402), .Z(n6400) );
  XNOR U6263 ( .A(n6403), .B(n6371), .Z(n6374) );
  XOR U6264 ( .A(n6404), .B(n6405), .Z(n6371) );
  AND U6265 ( .A(n6406), .B(n6407), .Z(n6405) );
  XOR U6266 ( .A(n6404), .B(n6408), .Z(n6406) );
  XNOR U6267 ( .A(n6409), .B(n6410), .Z(n6403) );
  NOR U6268 ( .A(n6411), .B(n6412), .Z(n6410) );
  XOR U6269 ( .A(n6409), .B(n6413), .Z(n6411) );
  XNOR U6270 ( .A(n6370), .B(n6377), .Z(n6391) );
  NOR U6271 ( .A(n6333), .B(n6414), .Z(n6377) );
  XOR U6272 ( .A(n6382), .B(n6381), .Z(n6370) );
  XNOR U6273 ( .A(n6415), .B(n6378), .Z(n6381) );
  XOR U6274 ( .A(n6416), .B(n6417), .Z(n6378) );
  AND U6275 ( .A(n6418), .B(n6419), .Z(n6417) );
  XNOR U6276 ( .A(n6420), .B(n6421), .Z(n6418) );
  IV U6277 ( .A(n6416), .Z(n6420) );
  XNOR U6278 ( .A(n6422), .B(n6423), .Z(n6415) );
  NOR U6279 ( .A(n6424), .B(n6425), .Z(n6423) );
  XNOR U6280 ( .A(n6422), .B(n6426), .Z(n6424) );
  XOR U6281 ( .A(n6427), .B(n6428), .Z(n6382) );
  NOR U6282 ( .A(n6429), .B(n6430), .Z(n6428) );
  XNOR U6283 ( .A(n6427), .B(n6431), .Z(n6429) );
  XNOR U6284 ( .A(n6310), .B(n6387), .Z(n6389) );
  XOR U6285 ( .A(n6432), .B(n6433), .Z(n6310) );
  AND U6286 ( .A(n11), .B(n6434), .Z(n6433) );
  XOR U6287 ( .A(n6435), .B(n6432), .Z(n6434) );
  AND U6288 ( .A(n6334), .B(n6333), .Z(n6387) );
  XOR U6289 ( .A(n6436), .B(n6414), .Z(n6333) );
  XNOR U6290 ( .A(p_input[16]), .B(p_input[2048]), .Z(n6414) );
  XOR U6291 ( .A(n6402), .B(n6401), .Z(n6436) );
  XNOR U6292 ( .A(n6437), .B(n6408), .Z(n6401) );
  XNOR U6293 ( .A(n6397), .B(n6396), .Z(n6408) );
  XOR U6294 ( .A(n6438), .B(n6393), .Z(n6396) );
  XNOR U6295 ( .A(n6439), .B(p_input[26]), .Z(n6393) );
  XNOR U6296 ( .A(p_input[2059]), .B(p_input[27]), .Z(n6438) );
  XOR U6297 ( .A(p_input[2060]), .B(p_input[28]), .Z(n6397) );
  XOR U6298 ( .A(n6407), .B(n6440), .Z(n6437) );
  IV U6299 ( .A(n6398), .Z(n6440) );
  XOR U6300 ( .A(p_input[17]), .B(p_input[2049]), .Z(n6398) );
  XOR U6301 ( .A(n6441), .B(n6413), .Z(n6407) );
  XNOR U6302 ( .A(p_input[2063]), .B(p_input[31]), .Z(n6413) );
  XOR U6303 ( .A(n6404), .B(n6412), .Z(n6441) );
  XOR U6304 ( .A(n6442), .B(n6409), .Z(n6412) );
  XOR U6305 ( .A(p_input[2061]), .B(p_input[29]), .Z(n6409) );
  XNOR U6306 ( .A(p_input[2062]), .B(p_input[30]), .Z(n6442) );
  XNOR U6307 ( .A(n6325), .B(p_input[25]), .Z(n6404) );
  XNOR U6308 ( .A(n6421), .B(n6419), .Z(n6402) );
  XNOR U6309 ( .A(n6443), .B(n6426), .Z(n6419) );
  XOR U6310 ( .A(p_input[2056]), .B(p_input[24]), .Z(n6426) );
  XOR U6311 ( .A(n6416), .B(n6425), .Z(n6443) );
  XOR U6312 ( .A(n6444), .B(n6422), .Z(n6425) );
  XOR U6313 ( .A(p_input[2054]), .B(p_input[22]), .Z(n6422) );
  XNOR U6314 ( .A(p_input[2055]), .B(p_input[23]), .Z(n6444) );
  XOR U6315 ( .A(p_input[18]), .B(p_input[2050]), .Z(n6416) );
  XNOR U6316 ( .A(n6431), .B(n6430), .Z(n6421) );
  XOR U6317 ( .A(n6445), .B(n6427), .Z(n6430) );
  XOR U6318 ( .A(p_input[19]), .B(p_input[2051]), .Z(n6427) );
  XNOR U6319 ( .A(p_input[2052]), .B(p_input[20]), .Z(n6445) );
  XOR U6320 ( .A(p_input[2053]), .B(p_input[21]), .Z(n6431) );
  IV U6321 ( .A(n6330), .Z(n6334) );
  XNOR U6322 ( .A(n6446), .B(n6447), .Z(n6330) );
  AND U6323 ( .A(n11), .B(n6448), .Z(n6447) );
  XNOR U6324 ( .A(n6449), .B(n6446), .Z(n6448) );
  XNOR U6325 ( .A(n6450), .B(n6451), .Z(n11) );
  AND U6326 ( .A(n6452), .B(n6453), .Z(n6451) );
  XOR U6327 ( .A(n6344), .B(n6450), .Z(n6453) );
  AND U6328 ( .A(n6454), .B(n6455), .Z(n6344) );
  XNOR U6329 ( .A(n6341), .B(n6450), .Z(n6452) );
  XOR U6330 ( .A(n6456), .B(n6457), .Z(n6341) );
  AND U6331 ( .A(n15), .B(n6458), .Z(n6457) );
  XOR U6332 ( .A(n6459), .B(n6456), .Z(n6458) );
  XOR U6333 ( .A(n6460), .B(n6461), .Z(n6450) );
  AND U6334 ( .A(n6462), .B(n6463), .Z(n6461) );
  XNOR U6335 ( .A(n6460), .B(n6454), .Z(n6463) );
  IV U6336 ( .A(n6359), .Z(n6454) );
  XOR U6337 ( .A(n6464), .B(n6465), .Z(n6359) );
  XOR U6338 ( .A(n6466), .B(n6455), .Z(n6465) );
  AND U6339 ( .A(n6386), .B(n6467), .Z(n6455) );
  AND U6340 ( .A(n6468), .B(n6469), .Z(n6466) );
  XOR U6341 ( .A(n6470), .B(n6464), .Z(n6468) );
  XNOR U6342 ( .A(n6356), .B(n6460), .Z(n6462) );
  XOR U6343 ( .A(n6471), .B(n6472), .Z(n6356) );
  AND U6344 ( .A(n15), .B(n6473), .Z(n6472) );
  XOR U6345 ( .A(n6474), .B(n6471), .Z(n6473) );
  XOR U6346 ( .A(n6475), .B(n6476), .Z(n6460) );
  AND U6347 ( .A(n6477), .B(n6478), .Z(n6476) );
  XNOR U6348 ( .A(n6475), .B(n6386), .Z(n6478) );
  XOR U6349 ( .A(n6479), .B(n6469), .Z(n6386) );
  XNOR U6350 ( .A(n6480), .B(n6464), .Z(n6469) );
  XOR U6351 ( .A(n6481), .B(n6482), .Z(n6464) );
  AND U6352 ( .A(n6483), .B(n6484), .Z(n6482) );
  XOR U6353 ( .A(n6485), .B(n6481), .Z(n6483) );
  XNOR U6354 ( .A(n6486), .B(n6487), .Z(n6480) );
  AND U6355 ( .A(n6488), .B(n6489), .Z(n6487) );
  XOR U6356 ( .A(n6486), .B(n6490), .Z(n6488) );
  XNOR U6357 ( .A(n6470), .B(n6467), .Z(n6479) );
  AND U6358 ( .A(n6491), .B(n6492), .Z(n6467) );
  XOR U6359 ( .A(n6493), .B(n6494), .Z(n6470) );
  AND U6360 ( .A(n6495), .B(n6496), .Z(n6494) );
  XOR U6361 ( .A(n6493), .B(n6497), .Z(n6495) );
  XNOR U6362 ( .A(n6383), .B(n6475), .Z(n6477) );
  XOR U6363 ( .A(n6498), .B(n6499), .Z(n6383) );
  AND U6364 ( .A(n15), .B(n6500), .Z(n6499) );
  XNOR U6365 ( .A(n6501), .B(n6498), .Z(n6500) );
  XOR U6366 ( .A(n6502), .B(n6503), .Z(n6475) );
  AND U6367 ( .A(n6504), .B(n6505), .Z(n6503) );
  XNOR U6368 ( .A(n6502), .B(n6491), .Z(n6505) );
  IV U6369 ( .A(n6435), .Z(n6491) );
  XNOR U6370 ( .A(n6506), .B(n6484), .Z(n6435) );
  XNOR U6371 ( .A(n6507), .B(n6490), .Z(n6484) );
  XOR U6372 ( .A(n6508), .B(n6509), .Z(n6490) );
  NOR U6373 ( .A(n6510), .B(n6511), .Z(n6509) );
  XNOR U6374 ( .A(n6508), .B(n6512), .Z(n6510) );
  XNOR U6375 ( .A(n6489), .B(n6481), .Z(n6507) );
  XOR U6376 ( .A(n6513), .B(n6514), .Z(n6481) );
  AND U6377 ( .A(n6515), .B(n6516), .Z(n6514) );
  XNOR U6378 ( .A(n6513), .B(n6517), .Z(n6515) );
  XNOR U6379 ( .A(n6518), .B(n6486), .Z(n6489) );
  XOR U6380 ( .A(n6519), .B(n6520), .Z(n6486) );
  AND U6381 ( .A(n6521), .B(n6522), .Z(n6520) );
  XOR U6382 ( .A(n6519), .B(n6523), .Z(n6521) );
  XNOR U6383 ( .A(n6524), .B(n6525), .Z(n6518) );
  NOR U6384 ( .A(n6526), .B(n6527), .Z(n6525) );
  XOR U6385 ( .A(n6524), .B(n6528), .Z(n6526) );
  XNOR U6386 ( .A(n6485), .B(n6492), .Z(n6506) );
  NOR U6387 ( .A(n6449), .B(n6529), .Z(n6492) );
  XOR U6388 ( .A(n6497), .B(n6496), .Z(n6485) );
  XNOR U6389 ( .A(n6530), .B(n6493), .Z(n6496) );
  XOR U6390 ( .A(n6531), .B(n6532), .Z(n6493) );
  AND U6391 ( .A(n6533), .B(n6534), .Z(n6532) );
  XOR U6392 ( .A(n6531), .B(n6535), .Z(n6533) );
  XNOR U6393 ( .A(n6536), .B(n6537), .Z(n6530) );
  NOR U6394 ( .A(n6538), .B(n6539), .Z(n6537) );
  XNOR U6395 ( .A(n6536), .B(n6540), .Z(n6538) );
  XOR U6396 ( .A(n6541), .B(n6542), .Z(n6497) );
  NOR U6397 ( .A(n6543), .B(n6544), .Z(n6542) );
  XNOR U6398 ( .A(n6541), .B(n6545), .Z(n6543) );
  XNOR U6399 ( .A(n6432), .B(n6502), .Z(n6504) );
  XOR U6400 ( .A(n6546), .B(n6547), .Z(n6432) );
  AND U6401 ( .A(n15), .B(n6548), .Z(n6547) );
  XOR U6402 ( .A(n6549), .B(n6546), .Z(n6548) );
  AND U6403 ( .A(n6446), .B(n6449), .Z(n6502) );
  XOR U6404 ( .A(n6550), .B(n6529), .Z(n6449) );
  XNOR U6405 ( .A(p_input[2048]), .B(p_input[32]), .Z(n6529) );
  XOR U6406 ( .A(n6517), .B(n6516), .Z(n6550) );
  XNOR U6407 ( .A(n6551), .B(n6523), .Z(n6516) );
  XNOR U6408 ( .A(n6512), .B(n6511), .Z(n6523) );
  XOR U6409 ( .A(n6552), .B(n6508), .Z(n6511) );
  XNOR U6410 ( .A(n6439), .B(p_input[42]), .Z(n6508) );
  XNOR U6411 ( .A(p_input[2059]), .B(p_input[43]), .Z(n6552) );
  XOR U6412 ( .A(p_input[2060]), .B(p_input[44]), .Z(n6512) );
  XNOR U6413 ( .A(n6522), .B(n6513), .Z(n6551) );
  XNOR U6414 ( .A(n6553), .B(p_input[33]), .Z(n6513) );
  XOR U6415 ( .A(n6554), .B(n6528), .Z(n6522) );
  XNOR U6416 ( .A(p_input[2063]), .B(p_input[47]), .Z(n6528) );
  XOR U6417 ( .A(n6519), .B(n6527), .Z(n6554) );
  XOR U6418 ( .A(n6555), .B(n6524), .Z(n6527) );
  XOR U6419 ( .A(p_input[2061]), .B(p_input[45]), .Z(n6524) );
  XNOR U6420 ( .A(p_input[2062]), .B(p_input[46]), .Z(n6555) );
  XNOR U6421 ( .A(n6325), .B(p_input[41]), .Z(n6519) );
  XNOR U6422 ( .A(n6535), .B(n6534), .Z(n6517) );
  XNOR U6423 ( .A(n6556), .B(n6540), .Z(n6534) );
  XOR U6424 ( .A(p_input[2056]), .B(p_input[40]), .Z(n6540) );
  XOR U6425 ( .A(n6531), .B(n6539), .Z(n6556) );
  XOR U6426 ( .A(n6557), .B(n6536), .Z(n6539) );
  XOR U6427 ( .A(p_input[2054]), .B(p_input[38]), .Z(n6536) );
  XNOR U6428 ( .A(p_input[2055]), .B(p_input[39]), .Z(n6557) );
  XNOR U6429 ( .A(n6328), .B(p_input[34]), .Z(n6531) );
  XNOR U6430 ( .A(n6545), .B(n6544), .Z(n6535) );
  XOR U6431 ( .A(n6558), .B(n6541), .Z(n6544) );
  XOR U6432 ( .A(p_input[2051]), .B(p_input[35]), .Z(n6541) );
  XNOR U6433 ( .A(p_input[2052]), .B(p_input[36]), .Z(n6558) );
  XOR U6434 ( .A(p_input[2053]), .B(p_input[37]), .Z(n6545) );
  XOR U6435 ( .A(n6559), .B(n6560), .Z(n6446) );
  AND U6436 ( .A(n15), .B(n6561), .Z(n6560) );
  XNOR U6437 ( .A(n6562), .B(n6559), .Z(n6561) );
  XNOR U6438 ( .A(n6563), .B(n6564), .Z(n15) );
  AND U6439 ( .A(n6565), .B(n6566), .Z(n6564) );
  XOR U6440 ( .A(n6459), .B(n6563), .Z(n6566) );
  AND U6441 ( .A(n6567), .B(n6568), .Z(n6459) );
  XNOR U6442 ( .A(n6456), .B(n6563), .Z(n6565) );
  XOR U6443 ( .A(n6569), .B(n6570), .Z(n6456) );
  AND U6444 ( .A(n19), .B(n6571), .Z(n6570) );
  XOR U6445 ( .A(n6572), .B(n6569), .Z(n6571) );
  XOR U6446 ( .A(n6573), .B(n6574), .Z(n6563) );
  AND U6447 ( .A(n6575), .B(n6576), .Z(n6574) );
  XNOR U6448 ( .A(n6573), .B(n6567), .Z(n6576) );
  IV U6449 ( .A(n6474), .Z(n6567) );
  XOR U6450 ( .A(n6577), .B(n6578), .Z(n6474) );
  XOR U6451 ( .A(n6579), .B(n6568), .Z(n6578) );
  AND U6452 ( .A(n6501), .B(n6580), .Z(n6568) );
  AND U6453 ( .A(n6581), .B(n6582), .Z(n6579) );
  XOR U6454 ( .A(n6583), .B(n6577), .Z(n6581) );
  XNOR U6455 ( .A(n6471), .B(n6573), .Z(n6575) );
  XOR U6456 ( .A(n6584), .B(n6585), .Z(n6471) );
  AND U6457 ( .A(n19), .B(n6586), .Z(n6585) );
  XOR U6458 ( .A(n6587), .B(n6584), .Z(n6586) );
  XOR U6459 ( .A(n6588), .B(n6589), .Z(n6573) );
  AND U6460 ( .A(n6590), .B(n6591), .Z(n6589) );
  XNOR U6461 ( .A(n6588), .B(n6501), .Z(n6591) );
  XOR U6462 ( .A(n6592), .B(n6582), .Z(n6501) );
  XNOR U6463 ( .A(n6593), .B(n6577), .Z(n6582) );
  XOR U6464 ( .A(n6594), .B(n6595), .Z(n6577) );
  AND U6465 ( .A(n6596), .B(n6597), .Z(n6595) );
  XOR U6466 ( .A(n6598), .B(n6594), .Z(n6596) );
  XNOR U6467 ( .A(n6599), .B(n6600), .Z(n6593) );
  AND U6468 ( .A(n6601), .B(n6602), .Z(n6600) );
  XOR U6469 ( .A(n6599), .B(n6603), .Z(n6601) );
  XNOR U6470 ( .A(n6583), .B(n6580), .Z(n6592) );
  AND U6471 ( .A(n6604), .B(n6605), .Z(n6580) );
  XOR U6472 ( .A(n6606), .B(n6607), .Z(n6583) );
  AND U6473 ( .A(n6608), .B(n6609), .Z(n6607) );
  XOR U6474 ( .A(n6606), .B(n6610), .Z(n6608) );
  XNOR U6475 ( .A(n6498), .B(n6588), .Z(n6590) );
  XOR U6476 ( .A(n6611), .B(n6612), .Z(n6498) );
  AND U6477 ( .A(n19), .B(n6613), .Z(n6612) );
  XNOR U6478 ( .A(n6614), .B(n6611), .Z(n6613) );
  XOR U6479 ( .A(n6615), .B(n6616), .Z(n6588) );
  AND U6480 ( .A(n6617), .B(n6618), .Z(n6616) );
  XNOR U6481 ( .A(n6615), .B(n6604), .Z(n6618) );
  IV U6482 ( .A(n6549), .Z(n6604) );
  XNOR U6483 ( .A(n6619), .B(n6597), .Z(n6549) );
  XNOR U6484 ( .A(n6620), .B(n6603), .Z(n6597) );
  XOR U6485 ( .A(n6621), .B(n6622), .Z(n6603) );
  NOR U6486 ( .A(n6623), .B(n6624), .Z(n6622) );
  XNOR U6487 ( .A(n6621), .B(n6625), .Z(n6623) );
  XNOR U6488 ( .A(n6602), .B(n6594), .Z(n6620) );
  XOR U6489 ( .A(n6626), .B(n6627), .Z(n6594) );
  AND U6490 ( .A(n6628), .B(n6629), .Z(n6627) );
  XNOR U6491 ( .A(n6626), .B(n6630), .Z(n6628) );
  XNOR U6492 ( .A(n6631), .B(n6599), .Z(n6602) );
  XOR U6493 ( .A(n6632), .B(n6633), .Z(n6599) );
  AND U6494 ( .A(n6634), .B(n6635), .Z(n6633) );
  XOR U6495 ( .A(n6632), .B(n6636), .Z(n6634) );
  XNOR U6496 ( .A(n6637), .B(n6638), .Z(n6631) );
  NOR U6497 ( .A(n6639), .B(n6640), .Z(n6638) );
  XOR U6498 ( .A(n6637), .B(n6641), .Z(n6639) );
  XNOR U6499 ( .A(n6598), .B(n6605), .Z(n6619) );
  NOR U6500 ( .A(n6562), .B(n6642), .Z(n6605) );
  XOR U6501 ( .A(n6610), .B(n6609), .Z(n6598) );
  XNOR U6502 ( .A(n6643), .B(n6606), .Z(n6609) );
  XOR U6503 ( .A(n6644), .B(n6645), .Z(n6606) );
  AND U6504 ( .A(n6646), .B(n6647), .Z(n6645) );
  XOR U6505 ( .A(n6644), .B(n6648), .Z(n6646) );
  XNOR U6506 ( .A(n6649), .B(n6650), .Z(n6643) );
  NOR U6507 ( .A(n6651), .B(n6652), .Z(n6650) );
  XNOR U6508 ( .A(n6649), .B(n6653), .Z(n6651) );
  XOR U6509 ( .A(n6654), .B(n6655), .Z(n6610) );
  NOR U6510 ( .A(n6656), .B(n6657), .Z(n6655) );
  XNOR U6511 ( .A(n6654), .B(n6658), .Z(n6656) );
  XNOR U6512 ( .A(n6546), .B(n6615), .Z(n6617) );
  XOR U6513 ( .A(n6659), .B(n6660), .Z(n6546) );
  AND U6514 ( .A(n19), .B(n6661), .Z(n6660) );
  XOR U6515 ( .A(n6662), .B(n6659), .Z(n6661) );
  AND U6516 ( .A(n6559), .B(n6562), .Z(n6615) );
  XOR U6517 ( .A(n6663), .B(n6642), .Z(n6562) );
  XNOR U6518 ( .A(p_input[2048]), .B(p_input[48]), .Z(n6642) );
  XOR U6519 ( .A(n6630), .B(n6629), .Z(n6663) );
  XNOR U6520 ( .A(n6664), .B(n6636), .Z(n6629) );
  XNOR U6521 ( .A(n6625), .B(n6624), .Z(n6636) );
  XOR U6522 ( .A(n6665), .B(n6621), .Z(n6624) );
  XNOR U6523 ( .A(n6439), .B(p_input[58]), .Z(n6621) );
  XNOR U6524 ( .A(p_input[2059]), .B(p_input[59]), .Z(n6665) );
  XOR U6525 ( .A(p_input[2060]), .B(p_input[60]), .Z(n6625) );
  XNOR U6526 ( .A(n6635), .B(n6626), .Z(n6664) );
  XNOR U6527 ( .A(n6553), .B(p_input[49]), .Z(n6626) );
  XOR U6528 ( .A(n6666), .B(n6641), .Z(n6635) );
  XNOR U6529 ( .A(p_input[2063]), .B(p_input[63]), .Z(n6641) );
  XOR U6530 ( .A(n6632), .B(n6640), .Z(n6666) );
  XOR U6531 ( .A(n6667), .B(n6637), .Z(n6640) );
  XOR U6532 ( .A(p_input[2061]), .B(p_input[61]), .Z(n6637) );
  XNOR U6533 ( .A(p_input[2062]), .B(p_input[62]), .Z(n6667) );
  XNOR U6534 ( .A(n6325), .B(p_input[57]), .Z(n6632) );
  XNOR U6535 ( .A(n6648), .B(n6647), .Z(n6630) );
  XNOR U6536 ( .A(n6668), .B(n6653), .Z(n6647) );
  XOR U6537 ( .A(p_input[2056]), .B(p_input[56]), .Z(n6653) );
  XOR U6538 ( .A(n6644), .B(n6652), .Z(n6668) );
  XOR U6539 ( .A(n6669), .B(n6649), .Z(n6652) );
  XOR U6540 ( .A(p_input[2054]), .B(p_input[54]), .Z(n6649) );
  XNOR U6541 ( .A(p_input[2055]), .B(p_input[55]), .Z(n6669) );
  XNOR U6542 ( .A(n6328), .B(p_input[50]), .Z(n6644) );
  XNOR U6543 ( .A(n6658), .B(n6657), .Z(n6648) );
  XOR U6544 ( .A(n6670), .B(n6654), .Z(n6657) );
  XOR U6545 ( .A(p_input[2051]), .B(p_input[51]), .Z(n6654) );
  XNOR U6546 ( .A(p_input[2052]), .B(p_input[52]), .Z(n6670) );
  XOR U6547 ( .A(p_input[2053]), .B(p_input[53]), .Z(n6658) );
  XOR U6548 ( .A(n6671), .B(n6672), .Z(n6559) );
  AND U6549 ( .A(n19), .B(n6673), .Z(n6672) );
  XNOR U6550 ( .A(n6674), .B(n6671), .Z(n6673) );
  XNOR U6551 ( .A(n6675), .B(n6676), .Z(n19) );
  AND U6552 ( .A(n6677), .B(n6678), .Z(n6676) );
  XOR U6553 ( .A(n6572), .B(n6675), .Z(n6678) );
  AND U6554 ( .A(n6679), .B(n6680), .Z(n6572) );
  XNOR U6555 ( .A(n6569), .B(n6675), .Z(n6677) );
  XOR U6556 ( .A(n6681), .B(n6682), .Z(n6569) );
  AND U6557 ( .A(n23), .B(n6683), .Z(n6682) );
  XOR U6558 ( .A(n6684), .B(n6681), .Z(n6683) );
  XOR U6559 ( .A(n6685), .B(n6686), .Z(n6675) );
  AND U6560 ( .A(n6687), .B(n6688), .Z(n6686) );
  XNOR U6561 ( .A(n6685), .B(n6679), .Z(n6688) );
  IV U6562 ( .A(n6587), .Z(n6679) );
  XOR U6563 ( .A(n6689), .B(n6690), .Z(n6587) );
  XOR U6564 ( .A(n6691), .B(n6680), .Z(n6690) );
  AND U6565 ( .A(n6614), .B(n6692), .Z(n6680) );
  AND U6566 ( .A(n6693), .B(n6694), .Z(n6691) );
  XOR U6567 ( .A(n6695), .B(n6689), .Z(n6693) );
  XNOR U6568 ( .A(n6584), .B(n6685), .Z(n6687) );
  XOR U6569 ( .A(n6696), .B(n6697), .Z(n6584) );
  AND U6570 ( .A(n23), .B(n6698), .Z(n6697) );
  XOR U6571 ( .A(n6699), .B(n6696), .Z(n6698) );
  XOR U6572 ( .A(n6700), .B(n6701), .Z(n6685) );
  AND U6573 ( .A(n6702), .B(n6703), .Z(n6701) );
  XNOR U6574 ( .A(n6700), .B(n6614), .Z(n6703) );
  XOR U6575 ( .A(n6704), .B(n6694), .Z(n6614) );
  XNOR U6576 ( .A(n6705), .B(n6689), .Z(n6694) );
  XOR U6577 ( .A(n6706), .B(n6707), .Z(n6689) );
  AND U6578 ( .A(n6708), .B(n6709), .Z(n6707) );
  XOR U6579 ( .A(n6710), .B(n6706), .Z(n6708) );
  XNOR U6580 ( .A(n6711), .B(n6712), .Z(n6705) );
  AND U6581 ( .A(n6713), .B(n6714), .Z(n6712) );
  XOR U6582 ( .A(n6711), .B(n6715), .Z(n6713) );
  XNOR U6583 ( .A(n6695), .B(n6692), .Z(n6704) );
  AND U6584 ( .A(n6716), .B(n6717), .Z(n6692) );
  XOR U6585 ( .A(n6718), .B(n6719), .Z(n6695) );
  AND U6586 ( .A(n6720), .B(n6721), .Z(n6719) );
  XOR U6587 ( .A(n6718), .B(n6722), .Z(n6720) );
  XNOR U6588 ( .A(n6611), .B(n6700), .Z(n6702) );
  XOR U6589 ( .A(n6723), .B(n6724), .Z(n6611) );
  AND U6590 ( .A(n23), .B(n6725), .Z(n6724) );
  XNOR U6591 ( .A(n6726), .B(n6723), .Z(n6725) );
  XOR U6592 ( .A(n6727), .B(n6728), .Z(n6700) );
  AND U6593 ( .A(n6729), .B(n6730), .Z(n6728) );
  XNOR U6594 ( .A(n6727), .B(n6716), .Z(n6730) );
  IV U6595 ( .A(n6662), .Z(n6716) );
  XNOR U6596 ( .A(n6731), .B(n6709), .Z(n6662) );
  XNOR U6597 ( .A(n6732), .B(n6715), .Z(n6709) );
  XOR U6598 ( .A(n6733), .B(n6734), .Z(n6715) );
  NOR U6599 ( .A(n6735), .B(n6736), .Z(n6734) );
  XNOR U6600 ( .A(n6733), .B(n6737), .Z(n6735) );
  XNOR U6601 ( .A(n6714), .B(n6706), .Z(n6732) );
  XOR U6602 ( .A(n6738), .B(n6739), .Z(n6706) );
  AND U6603 ( .A(n6740), .B(n6741), .Z(n6739) );
  XNOR U6604 ( .A(n6738), .B(n6742), .Z(n6740) );
  XNOR U6605 ( .A(n6743), .B(n6711), .Z(n6714) );
  XOR U6606 ( .A(n6744), .B(n6745), .Z(n6711) );
  AND U6607 ( .A(n6746), .B(n6747), .Z(n6745) );
  XOR U6608 ( .A(n6744), .B(n6748), .Z(n6746) );
  XNOR U6609 ( .A(n6749), .B(n6750), .Z(n6743) );
  NOR U6610 ( .A(n6751), .B(n6752), .Z(n6750) );
  XOR U6611 ( .A(n6749), .B(n6753), .Z(n6751) );
  XNOR U6612 ( .A(n6710), .B(n6717), .Z(n6731) );
  NOR U6613 ( .A(n6674), .B(n6754), .Z(n6717) );
  XOR U6614 ( .A(n6722), .B(n6721), .Z(n6710) );
  XNOR U6615 ( .A(n6755), .B(n6718), .Z(n6721) );
  XOR U6616 ( .A(n6756), .B(n6757), .Z(n6718) );
  AND U6617 ( .A(n6758), .B(n6759), .Z(n6757) );
  XOR U6618 ( .A(n6756), .B(n6760), .Z(n6758) );
  XNOR U6619 ( .A(n6761), .B(n6762), .Z(n6755) );
  NOR U6620 ( .A(n6763), .B(n6764), .Z(n6762) );
  XNOR U6621 ( .A(n6761), .B(n6765), .Z(n6763) );
  XOR U6622 ( .A(n6766), .B(n6767), .Z(n6722) );
  NOR U6623 ( .A(n6768), .B(n6769), .Z(n6767) );
  XNOR U6624 ( .A(n6766), .B(n6770), .Z(n6768) );
  XNOR U6625 ( .A(n6659), .B(n6727), .Z(n6729) );
  XOR U6626 ( .A(n6771), .B(n6772), .Z(n6659) );
  AND U6627 ( .A(n23), .B(n6773), .Z(n6772) );
  XOR U6628 ( .A(n6774), .B(n6771), .Z(n6773) );
  AND U6629 ( .A(n6671), .B(n6674), .Z(n6727) );
  XOR U6630 ( .A(n6775), .B(n6754), .Z(n6674) );
  XNOR U6631 ( .A(p_input[2048]), .B(p_input[64]), .Z(n6754) );
  XOR U6632 ( .A(n6742), .B(n6741), .Z(n6775) );
  XNOR U6633 ( .A(n6776), .B(n6748), .Z(n6741) );
  XNOR U6634 ( .A(n6737), .B(n6736), .Z(n6748) );
  XOR U6635 ( .A(n6777), .B(n6733), .Z(n6736) );
  XNOR U6636 ( .A(n6439), .B(p_input[74]), .Z(n6733) );
  XNOR U6637 ( .A(p_input[2059]), .B(p_input[75]), .Z(n6777) );
  XOR U6638 ( .A(p_input[2060]), .B(p_input[76]), .Z(n6737) );
  XNOR U6639 ( .A(n6747), .B(n6738), .Z(n6776) );
  XNOR U6640 ( .A(n6553), .B(p_input[65]), .Z(n6738) );
  XOR U6641 ( .A(n6778), .B(n6753), .Z(n6747) );
  XNOR U6642 ( .A(p_input[2063]), .B(p_input[79]), .Z(n6753) );
  XOR U6643 ( .A(n6744), .B(n6752), .Z(n6778) );
  XOR U6644 ( .A(n6779), .B(n6749), .Z(n6752) );
  XOR U6645 ( .A(p_input[2061]), .B(p_input[77]), .Z(n6749) );
  XNOR U6646 ( .A(p_input[2062]), .B(p_input[78]), .Z(n6779) );
  XNOR U6647 ( .A(n6325), .B(p_input[73]), .Z(n6744) );
  XNOR U6648 ( .A(n6760), .B(n6759), .Z(n6742) );
  XNOR U6649 ( .A(n6780), .B(n6765), .Z(n6759) );
  XOR U6650 ( .A(p_input[2056]), .B(p_input[72]), .Z(n6765) );
  XOR U6651 ( .A(n6756), .B(n6764), .Z(n6780) );
  XOR U6652 ( .A(n6781), .B(n6761), .Z(n6764) );
  XOR U6653 ( .A(p_input[2054]), .B(p_input[70]), .Z(n6761) );
  XNOR U6654 ( .A(p_input[2055]), .B(p_input[71]), .Z(n6781) );
  XNOR U6655 ( .A(n6328), .B(p_input[66]), .Z(n6756) );
  XNOR U6656 ( .A(n6770), .B(n6769), .Z(n6760) );
  XOR U6657 ( .A(n6782), .B(n6766), .Z(n6769) );
  XOR U6658 ( .A(p_input[2051]), .B(p_input[67]), .Z(n6766) );
  XNOR U6659 ( .A(p_input[2052]), .B(p_input[68]), .Z(n6782) );
  XOR U6660 ( .A(p_input[2053]), .B(p_input[69]), .Z(n6770) );
  XOR U6661 ( .A(n6783), .B(n6784), .Z(n6671) );
  AND U6662 ( .A(n23), .B(n6785), .Z(n6784) );
  XNOR U6663 ( .A(n6786), .B(n6783), .Z(n6785) );
  XNOR U6664 ( .A(n6787), .B(n6788), .Z(n23) );
  AND U6665 ( .A(n6789), .B(n6790), .Z(n6788) );
  XOR U6666 ( .A(n6684), .B(n6787), .Z(n6790) );
  AND U6667 ( .A(n6791), .B(n6792), .Z(n6684) );
  XNOR U6668 ( .A(n6681), .B(n6787), .Z(n6789) );
  XOR U6669 ( .A(n6793), .B(n6794), .Z(n6681) );
  AND U6670 ( .A(n27), .B(n6795), .Z(n6794) );
  XOR U6671 ( .A(n6796), .B(n6793), .Z(n6795) );
  XOR U6672 ( .A(n6797), .B(n6798), .Z(n6787) );
  AND U6673 ( .A(n6799), .B(n6800), .Z(n6798) );
  XNOR U6674 ( .A(n6797), .B(n6791), .Z(n6800) );
  IV U6675 ( .A(n6699), .Z(n6791) );
  XOR U6676 ( .A(n6801), .B(n6802), .Z(n6699) );
  XOR U6677 ( .A(n6803), .B(n6792), .Z(n6802) );
  AND U6678 ( .A(n6726), .B(n6804), .Z(n6792) );
  AND U6679 ( .A(n6805), .B(n6806), .Z(n6803) );
  XOR U6680 ( .A(n6807), .B(n6801), .Z(n6805) );
  XNOR U6681 ( .A(n6696), .B(n6797), .Z(n6799) );
  XOR U6682 ( .A(n6808), .B(n6809), .Z(n6696) );
  AND U6683 ( .A(n27), .B(n6810), .Z(n6809) );
  XOR U6684 ( .A(n6811), .B(n6808), .Z(n6810) );
  XOR U6685 ( .A(n6812), .B(n6813), .Z(n6797) );
  AND U6686 ( .A(n6814), .B(n6815), .Z(n6813) );
  XNOR U6687 ( .A(n6812), .B(n6726), .Z(n6815) );
  XOR U6688 ( .A(n6816), .B(n6806), .Z(n6726) );
  XNOR U6689 ( .A(n6817), .B(n6801), .Z(n6806) );
  XOR U6690 ( .A(n6818), .B(n6819), .Z(n6801) );
  AND U6691 ( .A(n6820), .B(n6821), .Z(n6819) );
  XOR U6692 ( .A(n6822), .B(n6818), .Z(n6820) );
  XNOR U6693 ( .A(n6823), .B(n6824), .Z(n6817) );
  AND U6694 ( .A(n6825), .B(n6826), .Z(n6824) );
  XOR U6695 ( .A(n6823), .B(n6827), .Z(n6825) );
  XNOR U6696 ( .A(n6807), .B(n6804), .Z(n6816) );
  AND U6697 ( .A(n6828), .B(n6829), .Z(n6804) );
  XOR U6698 ( .A(n6830), .B(n6831), .Z(n6807) );
  AND U6699 ( .A(n6832), .B(n6833), .Z(n6831) );
  XOR U6700 ( .A(n6830), .B(n6834), .Z(n6832) );
  XNOR U6701 ( .A(n6723), .B(n6812), .Z(n6814) );
  XOR U6702 ( .A(n6835), .B(n6836), .Z(n6723) );
  AND U6703 ( .A(n27), .B(n6837), .Z(n6836) );
  XNOR U6704 ( .A(n6838), .B(n6835), .Z(n6837) );
  XOR U6705 ( .A(n6839), .B(n6840), .Z(n6812) );
  AND U6706 ( .A(n6841), .B(n6842), .Z(n6840) );
  XNOR U6707 ( .A(n6839), .B(n6828), .Z(n6842) );
  IV U6708 ( .A(n6774), .Z(n6828) );
  XNOR U6709 ( .A(n6843), .B(n6821), .Z(n6774) );
  XNOR U6710 ( .A(n6844), .B(n6827), .Z(n6821) );
  XOR U6711 ( .A(n6845), .B(n6846), .Z(n6827) );
  NOR U6712 ( .A(n6847), .B(n6848), .Z(n6846) );
  XNOR U6713 ( .A(n6845), .B(n6849), .Z(n6847) );
  XNOR U6714 ( .A(n6826), .B(n6818), .Z(n6844) );
  XOR U6715 ( .A(n6850), .B(n6851), .Z(n6818) );
  AND U6716 ( .A(n6852), .B(n6853), .Z(n6851) );
  XNOR U6717 ( .A(n6850), .B(n6854), .Z(n6852) );
  XNOR U6718 ( .A(n6855), .B(n6823), .Z(n6826) );
  XOR U6719 ( .A(n6856), .B(n6857), .Z(n6823) );
  AND U6720 ( .A(n6858), .B(n6859), .Z(n6857) );
  XOR U6721 ( .A(n6856), .B(n6860), .Z(n6858) );
  XNOR U6722 ( .A(n6861), .B(n6862), .Z(n6855) );
  NOR U6723 ( .A(n6863), .B(n6864), .Z(n6862) );
  XOR U6724 ( .A(n6861), .B(n6865), .Z(n6863) );
  XNOR U6725 ( .A(n6822), .B(n6829), .Z(n6843) );
  NOR U6726 ( .A(n6786), .B(n6866), .Z(n6829) );
  XOR U6727 ( .A(n6834), .B(n6833), .Z(n6822) );
  XNOR U6728 ( .A(n6867), .B(n6830), .Z(n6833) );
  XOR U6729 ( .A(n6868), .B(n6869), .Z(n6830) );
  AND U6730 ( .A(n6870), .B(n6871), .Z(n6869) );
  XOR U6731 ( .A(n6868), .B(n6872), .Z(n6870) );
  XNOR U6732 ( .A(n6873), .B(n6874), .Z(n6867) );
  NOR U6733 ( .A(n6875), .B(n6876), .Z(n6874) );
  XNOR U6734 ( .A(n6873), .B(n6877), .Z(n6875) );
  XOR U6735 ( .A(n6878), .B(n6879), .Z(n6834) );
  NOR U6736 ( .A(n6880), .B(n6881), .Z(n6879) );
  XNOR U6737 ( .A(n6878), .B(n6882), .Z(n6880) );
  XNOR U6738 ( .A(n6771), .B(n6839), .Z(n6841) );
  XOR U6739 ( .A(n6883), .B(n6884), .Z(n6771) );
  AND U6740 ( .A(n27), .B(n6885), .Z(n6884) );
  XOR U6741 ( .A(n6886), .B(n6883), .Z(n6885) );
  AND U6742 ( .A(n6783), .B(n6786), .Z(n6839) );
  XOR U6743 ( .A(n6887), .B(n6866), .Z(n6786) );
  XNOR U6744 ( .A(p_input[2048]), .B(p_input[80]), .Z(n6866) );
  XOR U6745 ( .A(n6854), .B(n6853), .Z(n6887) );
  XNOR U6746 ( .A(n6888), .B(n6860), .Z(n6853) );
  XNOR U6747 ( .A(n6849), .B(n6848), .Z(n6860) );
  XOR U6748 ( .A(n6889), .B(n6845), .Z(n6848) );
  XNOR U6749 ( .A(n6439), .B(p_input[90]), .Z(n6845) );
  XNOR U6750 ( .A(p_input[2059]), .B(p_input[91]), .Z(n6889) );
  XOR U6751 ( .A(p_input[2060]), .B(p_input[92]), .Z(n6849) );
  XNOR U6752 ( .A(n6859), .B(n6850), .Z(n6888) );
  XNOR U6753 ( .A(n6553), .B(p_input[81]), .Z(n6850) );
  XOR U6754 ( .A(n6890), .B(n6865), .Z(n6859) );
  XNOR U6755 ( .A(p_input[2063]), .B(p_input[95]), .Z(n6865) );
  XOR U6756 ( .A(n6856), .B(n6864), .Z(n6890) );
  XOR U6757 ( .A(n6891), .B(n6861), .Z(n6864) );
  XOR U6758 ( .A(p_input[2061]), .B(p_input[93]), .Z(n6861) );
  XNOR U6759 ( .A(p_input[2062]), .B(p_input[94]), .Z(n6891) );
  XNOR U6760 ( .A(n6325), .B(p_input[89]), .Z(n6856) );
  XNOR U6761 ( .A(n6872), .B(n6871), .Z(n6854) );
  XNOR U6762 ( .A(n6892), .B(n6877), .Z(n6871) );
  XOR U6763 ( .A(p_input[2056]), .B(p_input[88]), .Z(n6877) );
  XOR U6764 ( .A(n6868), .B(n6876), .Z(n6892) );
  XOR U6765 ( .A(n6893), .B(n6873), .Z(n6876) );
  XOR U6766 ( .A(p_input[2054]), .B(p_input[86]), .Z(n6873) );
  XNOR U6767 ( .A(p_input[2055]), .B(p_input[87]), .Z(n6893) );
  XNOR U6768 ( .A(n6328), .B(p_input[82]), .Z(n6868) );
  XNOR U6769 ( .A(n6882), .B(n6881), .Z(n6872) );
  XOR U6770 ( .A(n6894), .B(n6878), .Z(n6881) );
  XOR U6771 ( .A(p_input[2051]), .B(p_input[83]), .Z(n6878) );
  XNOR U6772 ( .A(p_input[2052]), .B(p_input[84]), .Z(n6894) );
  XOR U6773 ( .A(p_input[2053]), .B(p_input[85]), .Z(n6882) );
  XOR U6774 ( .A(n6895), .B(n6896), .Z(n6783) );
  AND U6775 ( .A(n27), .B(n6897), .Z(n6896) );
  XNOR U6776 ( .A(n6898), .B(n6895), .Z(n6897) );
  XNOR U6777 ( .A(n6899), .B(n6900), .Z(n27) );
  AND U6778 ( .A(n6901), .B(n6902), .Z(n6900) );
  XOR U6779 ( .A(n6796), .B(n6899), .Z(n6902) );
  AND U6780 ( .A(n6903), .B(n6904), .Z(n6796) );
  XNOR U6781 ( .A(n6793), .B(n6899), .Z(n6901) );
  XOR U6782 ( .A(n6905), .B(n6906), .Z(n6793) );
  AND U6783 ( .A(n31), .B(n6907), .Z(n6906) );
  XOR U6784 ( .A(n6908), .B(n6905), .Z(n6907) );
  XOR U6785 ( .A(n6909), .B(n6910), .Z(n6899) );
  AND U6786 ( .A(n6911), .B(n6912), .Z(n6910) );
  XNOR U6787 ( .A(n6909), .B(n6903), .Z(n6912) );
  IV U6788 ( .A(n6811), .Z(n6903) );
  XOR U6789 ( .A(n6913), .B(n6914), .Z(n6811) );
  XOR U6790 ( .A(n6915), .B(n6904), .Z(n6914) );
  AND U6791 ( .A(n6838), .B(n6916), .Z(n6904) );
  AND U6792 ( .A(n6917), .B(n6918), .Z(n6915) );
  XOR U6793 ( .A(n6919), .B(n6913), .Z(n6917) );
  XNOR U6794 ( .A(n6808), .B(n6909), .Z(n6911) );
  XOR U6795 ( .A(n6920), .B(n6921), .Z(n6808) );
  AND U6796 ( .A(n31), .B(n6922), .Z(n6921) );
  XOR U6797 ( .A(n6923), .B(n6920), .Z(n6922) );
  XOR U6798 ( .A(n6924), .B(n6925), .Z(n6909) );
  AND U6799 ( .A(n6926), .B(n6927), .Z(n6925) );
  XNOR U6800 ( .A(n6924), .B(n6838), .Z(n6927) );
  XOR U6801 ( .A(n6928), .B(n6918), .Z(n6838) );
  XNOR U6802 ( .A(n6929), .B(n6913), .Z(n6918) );
  XOR U6803 ( .A(n6930), .B(n6931), .Z(n6913) );
  AND U6804 ( .A(n6932), .B(n6933), .Z(n6931) );
  XOR U6805 ( .A(n6934), .B(n6930), .Z(n6932) );
  XNOR U6806 ( .A(n6935), .B(n6936), .Z(n6929) );
  AND U6807 ( .A(n6937), .B(n6938), .Z(n6936) );
  XOR U6808 ( .A(n6935), .B(n6939), .Z(n6937) );
  XNOR U6809 ( .A(n6919), .B(n6916), .Z(n6928) );
  AND U6810 ( .A(n6940), .B(n6941), .Z(n6916) );
  XOR U6811 ( .A(n6942), .B(n6943), .Z(n6919) );
  AND U6812 ( .A(n6944), .B(n6945), .Z(n6943) );
  XOR U6813 ( .A(n6942), .B(n6946), .Z(n6944) );
  XNOR U6814 ( .A(n6835), .B(n6924), .Z(n6926) );
  XOR U6815 ( .A(n6947), .B(n6948), .Z(n6835) );
  AND U6816 ( .A(n31), .B(n6949), .Z(n6948) );
  XNOR U6817 ( .A(n6950), .B(n6947), .Z(n6949) );
  XOR U6818 ( .A(n6951), .B(n6952), .Z(n6924) );
  AND U6819 ( .A(n6953), .B(n6954), .Z(n6952) );
  XNOR U6820 ( .A(n6951), .B(n6940), .Z(n6954) );
  IV U6821 ( .A(n6886), .Z(n6940) );
  XNOR U6822 ( .A(n6955), .B(n6933), .Z(n6886) );
  XNOR U6823 ( .A(n6956), .B(n6939), .Z(n6933) );
  XNOR U6824 ( .A(n6957), .B(n6958), .Z(n6939) );
  NOR U6825 ( .A(n6959), .B(n6960), .Z(n6958) );
  XOR U6826 ( .A(n6957), .B(n6961), .Z(n6959) );
  XNOR U6827 ( .A(n6938), .B(n6930), .Z(n6956) );
  XOR U6828 ( .A(n6962), .B(n6963), .Z(n6930) );
  AND U6829 ( .A(n6964), .B(n6965), .Z(n6963) );
  XOR U6830 ( .A(n6962), .B(n6966), .Z(n6964) );
  XNOR U6831 ( .A(n6967), .B(n6935), .Z(n6938) );
  XOR U6832 ( .A(n6968), .B(n6969), .Z(n6935) );
  AND U6833 ( .A(n6970), .B(n6971), .Z(n6969) );
  XNOR U6834 ( .A(n6972), .B(n6973), .Z(n6970) );
  IV U6835 ( .A(n6968), .Z(n6972) );
  XNOR U6836 ( .A(n6974), .B(n6975), .Z(n6967) );
  NOR U6837 ( .A(n6976), .B(n6977), .Z(n6975) );
  XNOR U6838 ( .A(n6974), .B(n6978), .Z(n6976) );
  XNOR U6839 ( .A(n6934), .B(n6941), .Z(n6955) );
  NOR U6840 ( .A(n6898), .B(n6979), .Z(n6941) );
  XOR U6841 ( .A(n6946), .B(n6945), .Z(n6934) );
  XNOR U6842 ( .A(n6980), .B(n6942), .Z(n6945) );
  XOR U6843 ( .A(n6981), .B(n6982), .Z(n6942) );
  AND U6844 ( .A(n6983), .B(n6984), .Z(n6982) );
  XOR U6845 ( .A(n6981), .B(n6985), .Z(n6983) );
  XNOR U6846 ( .A(n6986), .B(n6987), .Z(n6980) );
  NOR U6847 ( .A(n6988), .B(n6989), .Z(n6987) );
  XNOR U6848 ( .A(n6986), .B(n6990), .Z(n6988) );
  XOR U6849 ( .A(n6991), .B(n6992), .Z(n6946) );
  NOR U6850 ( .A(n6993), .B(n6994), .Z(n6992) );
  XNOR U6851 ( .A(n6991), .B(n6995), .Z(n6993) );
  XNOR U6852 ( .A(n6883), .B(n6951), .Z(n6953) );
  XOR U6853 ( .A(n6996), .B(n6997), .Z(n6883) );
  AND U6854 ( .A(n31), .B(n6998), .Z(n6997) );
  XOR U6855 ( .A(n6999), .B(n6996), .Z(n6998) );
  AND U6856 ( .A(n6895), .B(n6898), .Z(n6951) );
  XOR U6857 ( .A(n7000), .B(n6979), .Z(n6898) );
  XNOR U6858 ( .A(p_input[2048]), .B(p_input[96]), .Z(n6979) );
  XNOR U6859 ( .A(n6966), .B(n6965), .Z(n7000) );
  XNOR U6860 ( .A(n7001), .B(n6973), .Z(n6965) );
  XNOR U6861 ( .A(n6961), .B(n6960), .Z(n6973) );
  XNOR U6862 ( .A(n7002), .B(n6957), .Z(n6960) );
  XNOR U6863 ( .A(p_input[106]), .B(p_input[2058]), .Z(n6957) );
  XOR U6864 ( .A(p_input[107]), .B(n6319), .Z(n7002) );
  XOR U6865 ( .A(p_input[108]), .B(p_input[2060]), .Z(n6961) );
  XNOR U6866 ( .A(n6971), .B(n6962), .Z(n7001) );
  XNOR U6867 ( .A(n6553), .B(p_input[97]), .Z(n6962) );
  XNOR U6868 ( .A(n7003), .B(n6978), .Z(n6971) );
  XNOR U6869 ( .A(p_input[111]), .B(n6322), .Z(n6978) );
  XOR U6870 ( .A(n6968), .B(n6977), .Z(n7003) );
  XOR U6871 ( .A(n7004), .B(n6974), .Z(n6977) );
  XOR U6872 ( .A(p_input[109]), .B(p_input[2061]), .Z(n6974) );
  XOR U6873 ( .A(p_input[110]), .B(n6324), .Z(n7004) );
  XOR U6874 ( .A(p_input[105]), .B(p_input[2057]), .Z(n6968) );
  XOR U6875 ( .A(n6985), .B(n6984), .Z(n6966) );
  XNOR U6876 ( .A(n7005), .B(n6990), .Z(n6984) );
  XOR U6877 ( .A(p_input[104]), .B(p_input[2056]), .Z(n6990) );
  XOR U6878 ( .A(n6981), .B(n6989), .Z(n7005) );
  XOR U6879 ( .A(n7006), .B(n6986), .Z(n6989) );
  XOR U6880 ( .A(p_input[102]), .B(p_input[2054]), .Z(n6986) );
  XOR U6881 ( .A(p_input[103]), .B(n7007), .Z(n7006) );
  XNOR U6882 ( .A(n6328), .B(p_input[98]), .Z(n6981) );
  XNOR U6883 ( .A(n6995), .B(n6994), .Z(n6985) );
  XOR U6884 ( .A(n7008), .B(n6991), .Z(n6994) );
  XOR U6885 ( .A(p_input[2051]), .B(p_input[99]), .Z(n6991) );
  XOR U6886 ( .A(p_input[100]), .B(n7009), .Z(n7008) );
  XOR U6887 ( .A(p_input[101]), .B(p_input[2053]), .Z(n6995) );
  XOR U6888 ( .A(n7010), .B(n7011), .Z(n6895) );
  AND U6889 ( .A(n31), .B(n7012), .Z(n7011) );
  XNOR U6890 ( .A(n7013), .B(n7010), .Z(n7012) );
  XNOR U6891 ( .A(n7014), .B(n7015), .Z(n31) );
  AND U6892 ( .A(n7016), .B(n7017), .Z(n7015) );
  XOR U6893 ( .A(n6908), .B(n7014), .Z(n7017) );
  AND U6894 ( .A(n7018), .B(n7019), .Z(n6908) );
  XNOR U6895 ( .A(n6905), .B(n7014), .Z(n7016) );
  XOR U6896 ( .A(n7020), .B(n7021), .Z(n6905) );
  AND U6897 ( .A(n35), .B(n7022), .Z(n7021) );
  XOR U6898 ( .A(n7023), .B(n7020), .Z(n7022) );
  XOR U6899 ( .A(n7024), .B(n7025), .Z(n7014) );
  AND U6900 ( .A(n7026), .B(n7027), .Z(n7025) );
  XNOR U6901 ( .A(n7024), .B(n7018), .Z(n7027) );
  IV U6902 ( .A(n6923), .Z(n7018) );
  XOR U6903 ( .A(n7028), .B(n7029), .Z(n6923) );
  XOR U6904 ( .A(n7030), .B(n7019), .Z(n7029) );
  AND U6905 ( .A(n6950), .B(n7031), .Z(n7019) );
  AND U6906 ( .A(n7032), .B(n7033), .Z(n7030) );
  XOR U6907 ( .A(n7034), .B(n7028), .Z(n7032) );
  XNOR U6908 ( .A(n6920), .B(n7024), .Z(n7026) );
  XOR U6909 ( .A(n7035), .B(n7036), .Z(n6920) );
  AND U6910 ( .A(n35), .B(n7037), .Z(n7036) );
  XOR U6911 ( .A(n7038), .B(n7035), .Z(n7037) );
  XOR U6912 ( .A(n7039), .B(n7040), .Z(n7024) );
  AND U6913 ( .A(n7041), .B(n7042), .Z(n7040) );
  XNOR U6914 ( .A(n7039), .B(n6950), .Z(n7042) );
  XOR U6915 ( .A(n7043), .B(n7033), .Z(n6950) );
  XNOR U6916 ( .A(n7044), .B(n7028), .Z(n7033) );
  XOR U6917 ( .A(n7045), .B(n7046), .Z(n7028) );
  AND U6918 ( .A(n7047), .B(n7048), .Z(n7046) );
  XOR U6919 ( .A(n7049), .B(n7045), .Z(n7047) );
  XNOR U6920 ( .A(n7050), .B(n7051), .Z(n7044) );
  AND U6921 ( .A(n7052), .B(n7053), .Z(n7051) );
  XOR U6922 ( .A(n7050), .B(n7054), .Z(n7052) );
  XNOR U6923 ( .A(n7034), .B(n7031), .Z(n7043) );
  AND U6924 ( .A(n7055), .B(n7056), .Z(n7031) );
  XOR U6925 ( .A(n7057), .B(n7058), .Z(n7034) );
  AND U6926 ( .A(n7059), .B(n7060), .Z(n7058) );
  XOR U6927 ( .A(n7057), .B(n7061), .Z(n7059) );
  XNOR U6928 ( .A(n6947), .B(n7039), .Z(n7041) );
  XOR U6929 ( .A(n7062), .B(n7063), .Z(n6947) );
  AND U6930 ( .A(n35), .B(n7064), .Z(n7063) );
  XNOR U6931 ( .A(n7065), .B(n7062), .Z(n7064) );
  XOR U6932 ( .A(n7066), .B(n7067), .Z(n7039) );
  AND U6933 ( .A(n7068), .B(n7069), .Z(n7067) );
  XNOR U6934 ( .A(n7066), .B(n7055), .Z(n7069) );
  IV U6935 ( .A(n6999), .Z(n7055) );
  XNOR U6936 ( .A(n7070), .B(n7048), .Z(n6999) );
  XNOR U6937 ( .A(n7071), .B(n7054), .Z(n7048) );
  XNOR U6938 ( .A(n7072), .B(n7073), .Z(n7054) );
  NOR U6939 ( .A(n7074), .B(n7075), .Z(n7073) );
  XOR U6940 ( .A(n7072), .B(n7076), .Z(n7074) );
  XNOR U6941 ( .A(n7053), .B(n7045), .Z(n7071) );
  XOR U6942 ( .A(n7077), .B(n7078), .Z(n7045) );
  AND U6943 ( .A(n7079), .B(n7080), .Z(n7078) );
  XOR U6944 ( .A(n7077), .B(n7081), .Z(n7079) );
  XNOR U6945 ( .A(n7082), .B(n7050), .Z(n7053) );
  XOR U6946 ( .A(n7083), .B(n7084), .Z(n7050) );
  AND U6947 ( .A(n7085), .B(n7086), .Z(n7084) );
  XNOR U6948 ( .A(n7087), .B(n7088), .Z(n7085) );
  IV U6949 ( .A(n7083), .Z(n7087) );
  XNOR U6950 ( .A(n7089), .B(n7090), .Z(n7082) );
  NOR U6951 ( .A(n7091), .B(n7092), .Z(n7090) );
  XNOR U6952 ( .A(n7089), .B(n7093), .Z(n7091) );
  XNOR U6953 ( .A(n7049), .B(n7056), .Z(n7070) );
  NOR U6954 ( .A(n7013), .B(n7094), .Z(n7056) );
  XOR U6955 ( .A(n7061), .B(n7060), .Z(n7049) );
  XNOR U6956 ( .A(n7095), .B(n7057), .Z(n7060) );
  XOR U6957 ( .A(n7096), .B(n7097), .Z(n7057) );
  AND U6958 ( .A(n7098), .B(n7099), .Z(n7097) );
  XNOR U6959 ( .A(n7100), .B(n7101), .Z(n7098) );
  IV U6960 ( .A(n7096), .Z(n7100) );
  XNOR U6961 ( .A(n7102), .B(n7103), .Z(n7095) );
  NOR U6962 ( .A(n7104), .B(n7105), .Z(n7103) );
  XNOR U6963 ( .A(n7102), .B(n7106), .Z(n7104) );
  XOR U6964 ( .A(n7107), .B(n7108), .Z(n7061) );
  NOR U6965 ( .A(n7109), .B(n7110), .Z(n7108) );
  XNOR U6966 ( .A(n7107), .B(n7111), .Z(n7109) );
  XNOR U6967 ( .A(n6996), .B(n7066), .Z(n7068) );
  XOR U6968 ( .A(n7112), .B(n7113), .Z(n6996) );
  AND U6969 ( .A(n35), .B(n7114), .Z(n7113) );
  XOR U6970 ( .A(n7115), .B(n7112), .Z(n7114) );
  AND U6971 ( .A(n7010), .B(n7013), .Z(n7066) );
  XOR U6972 ( .A(n7116), .B(n7094), .Z(n7013) );
  XNOR U6973 ( .A(p_input[112]), .B(p_input[2048]), .Z(n7094) );
  XNOR U6974 ( .A(n7081), .B(n7080), .Z(n7116) );
  XNOR U6975 ( .A(n7117), .B(n7088), .Z(n7080) );
  XNOR U6976 ( .A(n7076), .B(n7075), .Z(n7088) );
  XNOR U6977 ( .A(n7118), .B(n7072), .Z(n7075) );
  XNOR U6978 ( .A(p_input[122]), .B(p_input[2058]), .Z(n7072) );
  XOR U6979 ( .A(p_input[123]), .B(n6319), .Z(n7118) );
  XOR U6980 ( .A(p_input[124]), .B(p_input[2060]), .Z(n7076) );
  XOR U6981 ( .A(n7086), .B(n7119), .Z(n7117) );
  IV U6982 ( .A(n7077), .Z(n7119) );
  XOR U6983 ( .A(p_input[113]), .B(p_input[2049]), .Z(n7077) );
  XNOR U6984 ( .A(n7120), .B(n7093), .Z(n7086) );
  XNOR U6985 ( .A(p_input[127]), .B(n6322), .Z(n7093) );
  XOR U6986 ( .A(n7083), .B(n7092), .Z(n7120) );
  XOR U6987 ( .A(n7121), .B(n7089), .Z(n7092) );
  XOR U6988 ( .A(p_input[125]), .B(p_input[2061]), .Z(n7089) );
  XOR U6989 ( .A(p_input[126]), .B(n6324), .Z(n7121) );
  XOR U6990 ( .A(p_input[121]), .B(p_input[2057]), .Z(n7083) );
  XOR U6991 ( .A(n7101), .B(n7099), .Z(n7081) );
  XNOR U6992 ( .A(n7122), .B(n7106), .Z(n7099) );
  XOR U6993 ( .A(p_input[120]), .B(p_input[2056]), .Z(n7106) );
  XOR U6994 ( .A(n7096), .B(n7105), .Z(n7122) );
  XOR U6995 ( .A(n7123), .B(n7102), .Z(n7105) );
  XOR U6996 ( .A(p_input[118]), .B(p_input[2054]), .Z(n7102) );
  XOR U6997 ( .A(p_input[119]), .B(n7007), .Z(n7123) );
  XOR U6998 ( .A(p_input[114]), .B(p_input[2050]), .Z(n7096) );
  XNOR U6999 ( .A(n7111), .B(n7110), .Z(n7101) );
  XOR U7000 ( .A(n7124), .B(n7107), .Z(n7110) );
  XOR U7001 ( .A(p_input[115]), .B(p_input[2051]), .Z(n7107) );
  XOR U7002 ( .A(p_input[116]), .B(n7009), .Z(n7124) );
  XOR U7003 ( .A(p_input[117]), .B(p_input[2053]), .Z(n7111) );
  XOR U7004 ( .A(n7125), .B(n7126), .Z(n7010) );
  AND U7005 ( .A(n35), .B(n7127), .Z(n7126) );
  XNOR U7006 ( .A(n7128), .B(n7125), .Z(n7127) );
  XNOR U7007 ( .A(n7129), .B(n7130), .Z(n35) );
  AND U7008 ( .A(n7131), .B(n7132), .Z(n7130) );
  XOR U7009 ( .A(n7023), .B(n7129), .Z(n7132) );
  AND U7010 ( .A(n7133), .B(n7134), .Z(n7023) );
  XNOR U7011 ( .A(n7020), .B(n7129), .Z(n7131) );
  XOR U7012 ( .A(n7135), .B(n7136), .Z(n7020) );
  AND U7013 ( .A(n39), .B(n7137), .Z(n7136) );
  XOR U7014 ( .A(n7138), .B(n7135), .Z(n7137) );
  XOR U7015 ( .A(n7139), .B(n7140), .Z(n7129) );
  AND U7016 ( .A(n7141), .B(n7142), .Z(n7140) );
  XNOR U7017 ( .A(n7139), .B(n7133), .Z(n7142) );
  IV U7018 ( .A(n7038), .Z(n7133) );
  XOR U7019 ( .A(n7143), .B(n7144), .Z(n7038) );
  XOR U7020 ( .A(n7145), .B(n7134), .Z(n7144) );
  AND U7021 ( .A(n7065), .B(n7146), .Z(n7134) );
  AND U7022 ( .A(n7147), .B(n7148), .Z(n7145) );
  XOR U7023 ( .A(n7149), .B(n7143), .Z(n7147) );
  XNOR U7024 ( .A(n7035), .B(n7139), .Z(n7141) );
  XOR U7025 ( .A(n7150), .B(n7151), .Z(n7035) );
  AND U7026 ( .A(n39), .B(n7152), .Z(n7151) );
  XOR U7027 ( .A(n7153), .B(n7150), .Z(n7152) );
  XOR U7028 ( .A(n7154), .B(n7155), .Z(n7139) );
  AND U7029 ( .A(n7156), .B(n7157), .Z(n7155) );
  XNOR U7030 ( .A(n7154), .B(n7065), .Z(n7157) );
  XOR U7031 ( .A(n7158), .B(n7148), .Z(n7065) );
  XNOR U7032 ( .A(n7159), .B(n7143), .Z(n7148) );
  XOR U7033 ( .A(n7160), .B(n7161), .Z(n7143) );
  AND U7034 ( .A(n7162), .B(n7163), .Z(n7161) );
  XOR U7035 ( .A(n7164), .B(n7160), .Z(n7162) );
  XNOR U7036 ( .A(n7165), .B(n7166), .Z(n7159) );
  AND U7037 ( .A(n7167), .B(n7168), .Z(n7166) );
  XOR U7038 ( .A(n7165), .B(n7169), .Z(n7167) );
  XNOR U7039 ( .A(n7149), .B(n7146), .Z(n7158) );
  AND U7040 ( .A(n7170), .B(n7171), .Z(n7146) );
  XOR U7041 ( .A(n7172), .B(n7173), .Z(n7149) );
  AND U7042 ( .A(n7174), .B(n7175), .Z(n7173) );
  XOR U7043 ( .A(n7172), .B(n7176), .Z(n7174) );
  XNOR U7044 ( .A(n7062), .B(n7154), .Z(n7156) );
  XOR U7045 ( .A(n7177), .B(n7178), .Z(n7062) );
  AND U7046 ( .A(n39), .B(n7179), .Z(n7178) );
  XNOR U7047 ( .A(n7180), .B(n7177), .Z(n7179) );
  XOR U7048 ( .A(n7181), .B(n7182), .Z(n7154) );
  AND U7049 ( .A(n7183), .B(n7184), .Z(n7182) );
  XNOR U7050 ( .A(n7181), .B(n7170), .Z(n7184) );
  IV U7051 ( .A(n7115), .Z(n7170) );
  XNOR U7052 ( .A(n7185), .B(n7163), .Z(n7115) );
  XNOR U7053 ( .A(n7186), .B(n7169), .Z(n7163) );
  XNOR U7054 ( .A(n7187), .B(n7188), .Z(n7169) );
  NOR U7055 ( .A(n7189), .B(n7190), .Z(n7188) );
  XOR U7056 ( .A(n7187), .B(n7191), .Z(n7189) );
  XNOR U7057 ( .A(n7168), .B(n7160), .Z(n7186) );
  XOR U7058 ( .A(n7192), .B(n7193), .Z(n7160) );
  AND U7059 ( .A(n7194), .B(n7195), .Z(n7193) );
  XOR U7060 ( .A(n7192), .B(n7196), .Z(n7194) );
  XNOR U7061 ( .A(n7197), .B(n7165), .Z(n7168) );
  XOR U7062 ( .A(n7198), .B(n7199), .Z(n7165) );
  AND U7063 ( .A(n7200), .B(n7201), .Z(n7199) );
  XNOR U7064 ( .A(n7202), .B(n7203), .Z(n7200) );
  IV U7065 ( .A(n7198), .Z(n7202) );
  XNOR U7066 ( .A(n7204), .B(n7205), .Z(n7197) );
  NOR U7067 ( .A(n7206), .B(n7207), .Z(n7205) );
  XNOR U7068 ( .A(n7204), .B(n7208), .Z(n7206) );
  XNOR U7069 ( .A(n7164), .B(n7171), .Z(n7185) );
  NOR U7070 ( .A(n7128), .B(n7209), .Z(n7171) );
  XOR U7071 ( .A(n7176), .B(n7175), .Z(n7164) );
  XNOR U7072 ( .A(n7210), .B(n7172), .Z(n7175) );
  XOR U7073 ( .A(n7211), .B(n7212), .Z(n7172) );
  AND U7074 ( .A(n7213), .B(n7214), .Z(n7212) );
  XNOR U7075 ( .A(n7215), .B(n7216), .Z(n7213) );
  IV U7076 ( .A(n7211), .Z(n7215) );
  XNOR U7077 ( .A(n7217), .B(n7218), .Z(n7210) );
  NOR U7078 ( .A(n7219), .B(n7220), .Z(n7218) );
  XNOR U7079 ( .A(n7217), .B(n7221), .Z(n7219) );
  XOR U7080 ( .A(n7222), .B(n7223), .Z(n7176) );
  NOR U7081 ( .A(n7224), .B(n7225), .Z(n7223) );
  XNOR U7082 ( .A(n7222), .B(n7226), .Z(n7224) );
  XNOR U7083 ( .A(n7112), .B(n7181), .Z(n7183) );
  XOR U7084 ( .A(n7227), .B(n7228), .Z(n7112) );
  AND U7085 ( .A(n39), .B(n7229), .Z(n7228) );
  XOR U7086 ( .A(n7230), .B(n7227), .Z(n7229) );
  AND U7087 ( .A(n7125), .B(n7128), .Z(n7181) );
  XOR U7088 ( .A(n7231), .B(n7209), .Z(n7128) );
  XNOR U7089 ( .A(p_input[128]), .B(p_input[2048]), .Z(n7209) );
  XNOR U7090 ( .A(n7196), .B(n7195), .Z(n7231) );
  XNOR U7091 ( .A(n7232), .B(n7203), .Z(n7195) );
  XNOR U7092 ( .A(n7191), .B(n7190), .Z(n7203) );
  XNOR U7093 ( .A(n7233), .B(n7187), .Z(n7190) );
  XNOR U7094 ( .A(p_input[138]), .B(p_input[2058]), .Z(n7187) );
  XOR U7095 ( .A(p_input[139]), .B(n6319), .Z(n7233) );
  XOR U7096 ( .A(p_input[140]), .B(p_input[2060]), .Z(n7191) );
  XOR U7097 ( .A(n7201), .B(n7234), .Z(n7232) );
  IV U7098 ( .A(n7192), .Z(n7234) );
  XOR U7099 ( .A(p_input[129]), .B(p_input[2049]), .Z(n7192) );
  XNOR U7100 ( .A(n7235), .B(n7208), .Z(n7201) );
  XNOR U7101 ( .A(p_input[143]), .B(n6322), .Z(n7208) );
  XOR U7102 ( .A(n7198), .B(n7207), .Z(n7235) );
  XOR U7103 ( .A(n7236), .B(n7204), .Z(n7207) );
  XOR U7104 ( .A(p_input[141]), .B(p_input[2061]), .Z(n7204) );
  XOR U7105 ( .A(p_input[142]), .B(n6324), .Z(n7236) );
  XOR U7106 ( .A(p_input[137]), .B(p_input[2057]), .Z(n7198) );
  XOR U7107 ( .A(n7216), .B(n7214), .Z(n7196) );
  XNOR U7108 ( .A(n7237), .B(n7221), .Z(n7214) );
  XOR U7109 ( .A(p_input[136]), .B(p_input[2056]), .Z(n7221) );
  XOR U7110 ( .A(n7211), .B(n7220), .Z(n7237) );
  XOR U7111 ( .A(n7238), .B(n7217), .Z(n7220) );
  XOR U7112 ( .A(p_input[134]), .B(p_input[2054]), .Z(n7217) );
  XOR U7113 ( .A(p_input[135]), .B(n7007), .Z(n7238) );
  XOR U7114 ( .A(p_input[130]), .B(p_input[2050]), .Z(n7211) );
  XNOR U7115 ( .A(n7226), .B(n7225), .Z(n7216) );
  XOR U7116 ( .A(n7239), .B(n7222), .Z(n7225) );
  XOR U7117 ( .A(p_input[131]), .B(p_input[2051]), .Z(n7222) );
  XOR U7118 ( .A(p_input[132]), .B(n7009), .Z(n7239) );
  XOR U7119 ( .A(p_input[133]), .B(p_input[2053]), .Z(n7226) );
  XOR U7120 ( .A(n7240), .B(n7241), .Z(n7125) );
  AND U7121 ( .A(n39), .B(n7242), .Z(n7241) );
  XNOR U7122 ( .A(n7243), .B(n7240), .Z(n7242) );
  XNOR U7123 ( .A(n7244), .B(n7245), .Z(n39) );
  AND U7124 ( .A(n7246), .B(n7247), .Z(n7245) );
  XOR U7125 ( .A(n7138), .B(n7244), .Z(n7247) );
  AND U7126 ( .A(n7248), .B(n7249), .Z(n7138) );
  XNOR U7127 ( .A(n7135), .B(n7244), .Z(n7246) );
  XOR U7128 ( .A(n7250), .B(n7251), .Z(n7135) );
  AND U7129 ( .A(n43), .B(n7252), .Z(n7251) );
  XOR U7130 ( .A(n7253), .B(n7250), .Z(n7252) );
  XOR U7131 ( .A(n7254), .B(n7255), .Z(n7244) );
  AND U7132 ( .A(n7256), .B(n7257), .Z(n7255) );
  XNOR U7133 ( .A(n7254), .B(n7248), .Z(n7257) );
  IV U7134 ( .A(n7153), .Z(n7248) );
  XOR U7135 ( .A(n7258), .B(n7259), .Z(n7153) );
  XOR U7136 ( .A(n7260), .B(n7249), .Z(n7259) );
  AND U7137 ( .A(n7180), .B(n7261), .Z(n7249) );
  AND U7138 ( .A(n7262), .B(n7263), .Z(n7260) );
  XOR U7139 ( .A(n7264), .B(n7258), .Z(n7262) );
  XNOR U7140 ( .A(n7150), .B(n7254), .Z(n7256) );
  XOR U7141 ( .A(n7265), .B(n7266), .Z(n7150) );
  AND U7142 ( .A(n43), .B(n7267), .Z(n7266) );
  XOR U7143 ( .A(n7268), .B(n7265), .Z(n7267) );
  XOR U7144 ( .A(n7269), .B(n7270), .Z(n7254) );
  AND U7145 ( .A(n7271), .B(n7272), .Z(n7270) );
  XNOR U7146 ( .A(n7269), .B(n7180), .Z(n7272) );
  XOR U7147 ( .A(n7273), .B(n7263), .Z(n7180) );
  XNOR U7148 ( .A(n7274), .B(n7258), .Z(n7263) );
  XOR U7149 ( .A(n7275), .B(n7276), .Z(n7258) );
  AND U7150 ( .A(n7277), .B(n7278), .Z(n7276) );
  XOR U7151 ( .A(n7279), .B(n7275), .Z(n7277) );
  XNOR U7152 ( .A(n7280), .B(n7281), .Z(n7274) );
  AND U7153 ( .A(n7282), .B(n7283), .Z(n7281) );
  XOR U7154 ( .A(n7280), .B(n7284), .Z(n7282) );
  XNOR U7155 ( .A(n7264), .B(n7261), .Z(n7273) );
  AND U7156 ( .A(n7285), .B(n7286), .Z(n7261) );
  XOR U7157 ( .A(n7287), .B(n7288), .Z(n7264) );
  AND U7158 ( .A(n7289), .B(n7290), .Z(n7288) );
  XOR U7159 ( .A(n7287), .B(n7291), .Z(n7289) );
  XNOR U7160 ( .A(n7177), .B(n7269), .Z(n7271) );
  XOR U7161 ( .A(n7292), .B(n7293), .Z(n7177) );
  AND U7162 ( .A(n43), .B(n7294), .Z(n7293) );
  XNOR U7163 ( .A(n7295), .B(n7292), .Z(n7294) );
  XOR U7164 ( .A(n7296), .B(n7297), .Z(n7269) );
  AND U7165 ( .A(n7298), .B(n7299), .Z(n7297) );
  XNOR U7166 ( .A(n7296), .B(n7285), .Z(n7299) );
  IV U7167 ( .A(n7230), .Z(n7285) );
  XNOR U7168 ( .A(n7300), .B(n7278), .Z(n7230) );
  XNOR U7169 ( .A(n7301), .B(n7284), .Z(n7278) );
  XNOR U7170 ( .A(n7302), .B(n7303), .Z(n7284) );
  NOR U7171 ( .A(n7304), .B(n7305), .Z(n7303) );
  XOR U7172 ( .A(n7302), .B(n7306), .Z(n7304) );
  XNOR U7173 ( .A(n7283), .B(n7275), .Z(n7301) );
  XOR U7174 ( .A(n7307), .B(n7308), .Z(n7275) );
  AND U7175 ( .A(n7309), .B(n7310), .Z(n7308) );
  XOR U7176 ( .A(n7307), .B(n7311), .Z(n7309) );
  XNOR U7177 ( .A(n7312), .B(n7280), .Z(n7283) );
  XOR U7178 ( .A(n7313), .B(n7314), .Z(n7280) );
  AND U7179 ( .A(n7315), .B(n7316), .Z(n7314) );
  XNOR U7180 ( .A(n7317), .B(n7318), .Z(n7315) );
  IV U7181 ( .A(n7313), .Z(n7317) );
  XNOR U7182 ( .A(n7319), .B(n7320), .Z(n7312) );
  NOR U7183 ( .A(n7321), .B(n7322), .Z(n7320) );
  XNOR U7184 ( .A(n7319), .B(n7323), .Z(n7321) );
  XNOR U7185 ( .A(n7279), .B(n7286), .Z(n7300) );
  NOR U7186 ( .A(n7243), .B(n7324), .Z(n7286) );
  XOR U7187 ( .A(n7291), .B(n7290), .Z(n7279) );
  XNOR U7188 ( .A(n7325), .B(n7287), .Z(n7290) );
  XOR U7189 ( .A(n7326), .B(n7327), .Z(n7287) );
  AND U7190 ( .A(n7328), .B(n7329), .Z(n7327) );
  XNOR U7191 ( .A(n7330), .B(n7331), .Z(n7328) );
  IV U7192 ( .A(n7326), .Z(n7330) );
  XNOR U7193 ( .A(n7332), .B(n7333), .Z(n7325) );
  NOR U7194 ( .A(n7334), .B(n7335), .Z(n7333) );
  XNOR U7195 ( .A(n7332), .B(n7336), .Z(n7334) );
  XOR U7196 ( .A(n7337), .B(n7338), .Z(n7291) );
  NOR U7197 ( .A(n7339), .B(n7340), .Z(n7338) );
  XNOR U7198 ( .A(n7337), .B(n7341), .Z(n7339) );
  XNOR U7199 ( .A(n7227), .B(n7296), .Z(n7298) );
  XOR U7200 ( .A(n7342), .B(n7343), .Z(n7227) );
  AND U7201 ( .A(n43), .B(n7344), .Z(n7343) );
  XOR U7202 ( .A(n7345), .B(n7342), .Z(n7344) );
  AND U7203 ( .A(n7240), .B(n7243), .Z(n7296) );
  XOR U7204 ( .A(n7346), .B(n7324), .Z(n7243) );
  XNOR U7205 ( .A(p_input[144]), .B(p_input[2048]), .Z(n7324) );
  XNOR U7206 ( .A(n7311), .B(n7310), .Z(n7346) );
  XNOR U7207 ( .A(n7347), .B(n7318), .Z(n7310) );
  XNOR U7208 ( .A(n7306), .B(n7305), .Z(n7318) );
  XNOR U7209 ( .A(n7348), .B(n7302), .Z(n7305) );
  XNOR U7210 ( .A(p_input[154]), .B(p_input[2058]), .Z(n7302) );
  XOR U7211 ( .A(p_input[155]), .B(n6319), .Z(n7348) );
  XOR U7212 ( .A(p_input[156]), .B(p_input[2060]), .Z(n7306) );
  XOR U7213 ( .A(n7316), .B(n7349), .Z(n7347) );
  IV U7214 ( .A(n7307), .Z(n7349) );
  XOR U7215 ( .A(p_input[145]), .B(p_input[2049]), .Z(n7307) );
  XNOR U7216 ( .A(n7350), .B(n7323), .Z(n7316) );
  XNOR U7217 ( .A(p_input[159]), .B(n6322), .Z(n7323) );
  XOR U7218 ( .A(n7313), .B(n7322), .Z(n7350) );
  XOR U7219 ( .A(n7351), .B(n7319), .Z(n7322) );
  XOR U7220 ( .A(p_input[157]), .B(p_input[2061]), .Z(n7319) );
  XOR U7221 ( .A(p_input[158]), .B(n6324), .Z(n7351) );
  XOR U7222 ( .A(p_input[153]), .B(p_input[2057]), .Z(n7313) );
  XOR U7223 ( .A(n7331), .B(n7329), .Z(n7311) );
  XNOR U7224 ( .A(n7352), .B(n7336), .Z(n7329) );
  XOR U7225 ( .A(p_input[152]), .B(p_input[2056]), .Z(n7336) );
  XOR U7226 ( .A(n7326), .B(n7335), .Z(n7352) );
  XOR U7227 ( .A(n7353), .B(n7332), .Z(n7335) );
  XOR U7228 ( .A(p_input[150]), .B(p_input[2054]), .Z(n7332) );
  XOR U7229 ( .A(p_input[151]), .B(n7007), .Z(n7353) );
  XOR U7230 ( .A(p_input[146]), .B(p_input[2050]), .Z(n7326) );
  XNOR U7231 ( .A(n7341), .B(n7340), .Z(n7331) );
  XOR U7232 ( .A(n7354), .B(n7337), .Z(n7340) );
  XOR U7233 ( .A(p_input[147]), .B(p_input[2051]), .Z(n7337) );
  XOR U7234 ( .A(p_input[148]), .B(n7009), .Z(n7354) );
  XOR U7235 ( .A(p_input[149]), .B(p_input[2053]), .Z(n7341) );
  XOR U7236 ( .A(n7355), .B(n7356), .Z(n7240) );
  AND U7237 ( .A(n43), .B(n7357), .Z(n7356) );
  XNOR U7238 ( .A(n7358), .B(n7355), .Z(n7357) );
  XNOR U7239 ( .A(n7359), .B(n7360), .Z(n43) );
  AND U7240 ( .A(n7361), .B(n7362), .Z(n7360) );
  XOR U7241 ( .A(n7253), .B(n7359), .Z(n7362) );
  AND U7242 ( .A(n7363), .B(n7364), .Z(n7253) );
  XNOR U7243 ( .A(n7250), .B(n7359), .Z(n7361) );
  XOR U7244 ( .A(n7365), .B(n7366), .Z(n7250) );
  AND U7245 ( .A(n47), .B(n7367), .Z(n7366) );
  XOR U7246 ( .A(n7368), .B(n7365), .Z(n7367) );
  XOR U7247 ( .A(n7369), .B(n7370), .Z(n7359) );
  AND U7248 ( .A(n7371), .B(n7372), .Z(n7370) );
  XNOR U7249 ( .A(n7369), .B(n7363), .Z(n7372) );
  IV U7250 ( .A(n7268), .Z(n7363) );
  XOR U7251 ( .A(n7373), .B(n7374), .Z(n7268) );
  XOR U7252 ( .A(n7375), .B(n7364), .Z(n7374) );
  AND U7253 ( .A(n7295), .B(n7376), .Z(n7364) );
  AND U7254 ( .A(n7377), .B(n7378), .Z(n7375) );
  XOR U7255 ( .A(n7379), .B(n7373), .Z(n7377) );
  XNOR U7256 ( .A(n7265), .B(n7369), .Z(n7371) );
  XOR U7257 ( .A(n7380), .B(n7381), .Z(n7265) );
  AND U7258 ( .A(n47), .B(n7382), .Z(n7381) );
  XOR U7259 ( .A(n7383), .B(n7380), .Z(n7382) );
  XOR U7260 ( .A(n7384), .B(n7385), .Z(n7369) );
  AND U7261 ( .A(n7386), .B(n7387), .Z(n7385) );
  XNOR U7262 ( .A(n7384), .B(n7295), .Z(n7387) );
  XOR U7263 ( .A(n7388), .B(n7378), .Z(n7295) );
  XNOR U7264 ( .A(n7389), .B(n7373), .Z(n7378) );
  XOR U7265 ( .A(n7390), .B(n7391), .Z(n7373) );
  AND U7266 ( .A(n7392), .B(n7393), .Z(n7391) );
  XOR U7267 ( .A(n7394), .B(n7390), .Z(n7392) );
  XNOR U7268 ( .A(n7395), .B(n7396), .Z(n7389) );
  AND U7269 ( .A(n7397), .B(n7398), .Z(n7396) );
  XOR U7270 ( .A(n7395), .B(n7399), .Z(n7397) );
  XNOR U7271 ( .A(n7379), .B(n7376), .Z(n7388) );
  AND U7272 ( .A(n7400), .B(n7401), .Z(n7376) );
  XOR U7273 ( .A(n7402), .B(n7403), .Z(n7379) );
  AND U7274 ( .A(n7404), .B(n7405), .Z(n7403) );
  XOR U7275 ( .A(n7402), .B(n7406), .Z(n7404) );
  XNOR U7276 ( .A(n7292), .B(n7384), .Z(n7386) );
  XOR U7277 ( .A(n7407), .B(n7408), .Z(n7292) );
  AND U7278 ( .A(n47), .B(n7409), .Z(n7408) );
  XNOR U7279 ( .A(n7410), .B(n7407), .Z(n7409) );
  XOR U7280 ( .A(n7411), .B(n7412), .Z(n7384) );
  AND U7281 ( .A(n7413), .B(n7414), .Z(n7412) );
  XNOR U7282 ( .A(n7411), .B(n7400), .Z(n7414) );
  IV U7283 ( .A(n7345), .Z(n7400) );
  XNOR U7284 ( .A(n7415), .B(n7393), .Z(n7345) );
  XNOR U7285 ( .A(n7416), .B(n7399), .Z(n7393) );
  XNOR U7286 ( .A(n7417), .B(n7418), .Z(n7399) );
  NOR U7287 ( .A(n7419), .B(n7420), .Z(n7418) );
  XOR U7288 ( .A(n7417), .B(n7421), .Z(n7419) );
  XNOR U7289 ( .A(n7398), .B(n7390), .Z(n7416) );
  XOR U7290 ( .A(n7422), .B(n7423), .Z(n7390) );
  AND U7291 ( .A(n7424), .B(n7425), .Z(n7423) );
  XOR U7292 ( .A(n7422), .B(n7426), .Z(n7424) );
  XNOR U7293 ( .A(n7427), .B(n7395), .Z(n7398) );
  XOR U7294 ( .A(n7428), .B(n7429), .Z(n7395) );
  AND U7295 ( .A(n7430), .B(n7431), .Z(n7429) );
  XNOR U7296 ( .A(n7432), .B(n7433), .Z(n7430) );
  IV U7297 ( .A(n7428), .Z(n7432) );
  XNOR U7298 ( .A(n7434), .B(n7435), .Z(n7427) );
  NOR U7299 ( .A(n7436), .B(n7437), .Z(n7435) );
  XNOR U7300 ( .A(n7434), .B(n7438), .Z(n7436) );
  XNOR U7301 ( .A(n7394), .B(n7401), .Z(n7415) );
  NOR U7302 ( .A(n7358), .B(n7439), .Z(n7401) );
  XOR U7303 ( .A(n7406), .B(n7405), .Z(n7394) );
  XNOR U7304 ( .A(n7440), .B(n7402), .Z(n7405) );
  XOR U7305 ( .A(n7441), .B(n7442), .Z(n7402) );
  AND U7306 ( .A(n7443), .B(n7444), .Z(n7442) );
  XNOR U7307 ( .A(n7445), .B(n7446), .Z(n7443) );
  IV U7308 ( .A(n7441), .Z(n7445) );
  XNOR U7309 ( .A(n7447), .B(n7448), .Z(n7440) );
  NOR U7310 ( .A(n7449), .B(n7450), .Z(n7448) );
  XNOR U7311 ( .A(n7447), .B(n7451), .Z(n7449) );
  XOR U7312 ( .A(n7452), .B(n7453), .Z(n7406) );
  NOR U7313 ( .A(n7454), .B(n7455), .Z(n7453) );
  XNOR U7314 ( .A(n7452), .B(n7456), .Z(n7454) );
  XNOR U7315 ( .A(n7342), .B(n7411), .Z(n7413) );
  XOR U7316 ( .A(n7457), .B(n7458), .Z(n7342) );
  AND U7317 ( .A(n47), .B(n7459), .Z(n7458) );
  XOR U7318 ( .A(n7460), .B(n7457), .Z(n7459) );
  AND U7319 ( .A(n7355), .B(n7358), .Z(n7411) );
  XOR U7320 ( .A(n7461), .B(n7439), .Z(n7358) );
  XNOR U7321 ( .A(p_input[160]), .B(p_input[2048]), .Z(n7439) );
  XNOR U7322 ( .A(n7426), .B(n7425), .Z(n7461) );
  XNOR U7323 ( .A(n7462), .B(n7433), .Z(n7425) );
  XNOR U7324 ( .A(n7421), .B(n7420), .Z(n7433) );
  XNOR U7325 ( .A(n7463), .B(n7417), .Z(n7420) );
  XNOR U7326 ( .A(p_input[170]), .B(p_input[2058]), .Z(n7417) );
  XOR U7327 ( .A(p_input[171]), .B(n6319), .Z(n7463) );
  XOR U7328 ( .A(p_input[172]), .B(p_input[2060]), .Z(n7421) );
  XOR U7329 ( .A(n7431), .B(n7464), .Z(n7462) );
  IV U7330 ( .A(n7422), .Z(n7464) );
  XOR U7331 ( .A(p_input[161]), .B(p_input[2049]), .Z(n7422) );
  XNOR U7332 ( .A(n7465), .B(n7438), .Z(n7431) );
  XNOR U7333 ( .A(p_input[175]), .B(n6322), .Z(n7438) );
  XOR U7334 ( .A(n7428), .B(n7437), .Z(n7465) );
  XOR U7335 ( .A(n7466), .B(n7434), .Z(n7437) );
  XOR U7336 ( .A(p_input[173]), .B(p_input[2061]), .Z(n7434) );
  XOR U7337 ( .A(p_input[174]), .B(n6324), .Z(n7466) );
  XOR U7338 ( .A(p_input[169]), .B(p_input[2057]), .Z(n7428) );
  XOR U7339 ( .A(n7446), .B(n7444), .Z(n7426) );
  XNOR U7340 ( .A(n7467), .B(n7451), .Z(n7444) );
  XOR U7341 ( .A(p_input[168]), .B(p_input[2056]), .Z(n7451) );
  XOR U7342 ( .A(n7441), .B(n7450), .Z(n7467) );
  XOR U7343 ( .A(n7468), .B(n7447), .Z(n7450) );
  XOR U7344 ( .A(p_input[166]), .B(p_input[2054]), .Z(n7447) );
  XOR U7345 ( .A(p_input[167]), .B(n7007), .Z(n7468) );
  XOR U7346 ( .A(p_input[162]), .B(p_input[2050]), .Z(n7441) );
  XNOR U7347 ( .A(n7456), .B(n7455), .Z(n7446) );
  XOR U7348 ( .A(n7469), .B(n7452), .Z(n7455) );
  XOR U7349 ( .A(p_input[163]), .B(p_input[2051]), .Z(n7452) );
  XOR U7350 ( .A(p_input[164]), .B(n7009), .Z(n7469) );
  XOR U7351 ( .A(p_input[165]), .B(p_input[2053]), .Z(n7456) );
  XOR U7352 ( .A(n7470), .B(n7471), .Z(n7355) );
  AND U7353 ( .A(n47), .B(n7472), .Z(n7471) );
  XNOR U7354 ( .A(n7473), .B(n7470), .Z(n7472) );
  XNOR U7355 ( .A(n7474), .B(n7475), .Z(n47) );
  AND U7356 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR U7357 ( .A(n7368), .B(n7474), .Z(n7477) );
  AND U7358 ( .A(n7478), .B(n7479), .Z(n7368) );
  XNOR U7359 ( .A(n7365), .B(n7474), .Z(n7476) );
  XOR U7360 ( .A(n7480), .B(n7481), .Z(n7365) );
  AND U7361 ( .A(n51), .B(n7482), .Z(n7481) );
  XOR U7362 ( .A(n7483), .B(n7480), .Z(n7482) );
  XOR U7363 ( .A(n7484), .B(n7485), .Z(n7474) );
  AND U7364 ( .A(n7486), .B(n7487), .Z(n7485) );
  XNOR U7365 ( .A(n7484), .B(n7478), .Z(n7487) );
  IV U7366 ( .A(n7383), .Z(n7478) );
  XOR U7367 ( .A(n7488), .B(n7489), .Z(n7383) );
  XOR U7368 ( .A(n7490), .B(n7479), .Z(n7489) );
  AND U7369 ( .A(n7410), .B(n7491), .Z(n7479) );
  AND U7370 ( .A(n7492), .B(n7493), .Z(n7490) );
  XOR U7371 ( .A(n7494), .B(n7488), .Z(n7492) );
  XNOR U7372 ( .A(n7380), .B(n7484), .Z(n7486) );
  XOR U7373 ( .A(n7495), .B(n7496), .Z(n7380) );
  AND U7374 ( .A(n51), .B(n7497), .Z(n7496) );
  XOR U7375 ( .A(n7498), .B(n7495), .Z(n7497) );
  XOR U7376 ( .A(n7499), .B(n7500), .Z(n7484) );
  AND U7377 ( .A(n7501), .B(n7502), .Z(n7500) );
  XNOR U7378 ( .A(n7499), .B(n7410), .Z(n7502) );
  XOR U7379 ( .A(n7503), .B(n7493), .Z(n7410) );
  XNOR U7380 ( .A(n7504), .B(n7488), .Z(n7493) );
  XOR U7381 ( .A(n7505), .B(n7506), .Z(n7488) );
  AND U7382 ( .A(n7507), .B(n7508), .Z(n7506) );
  XOR U7383 ( .A(n7509), .B(n7505), .Z(n7507) );
  XNOR U7384 ( .A(n7510), .B(n7511), .Z(n7504) );
  AND U7385 ( .A(n7512), .B(n7513), .Z(n7511) );
  XOR U7386 ( .A(n7510), .B(n7514), .Z(n7512) );
  XNOR U7387 ( .A(n7494), .B(n7491), .Z(n7503) );
  AND U7388 ( .A(n7515), .B(n7516), .Z(n7491) );
  XOR U7389 ( .A(n7517), .B(n7518), .Z(n7494) );
  AND U7390 ( .A(n7519), .B(n7520), .Z(n7518) );
  XOR U7391 ( .A(n7517), .B(n7521), .Z(n7519) );
  XNOR U7392 ( .A(n7407), .B(n7499), .Z(n7501) );
  XOR U7393 ( .A(n7522), .B(n7523), .Z(n7407) );
  AND U7394 ( .A(n51), .B(n7524), .Z(n7523) );
  XNOR U7395 ( .A(n7525), .B(n7522), .Z(n7524) );
  XOR U7396 ( .A(n7526), .B(n7527), .Z(n7499) );
  AND U7397 ( .A(n7528), .B(n7529), .Z(n7527) );
  XNOR U7398 ( .A(n7526), .B(n7515), .Z(n7529) );
  IV U7399 ( .A(n7460), .Z(n7515) );
  XNOR U7400 ( .A(n7530), .B(n7508), .Z(n7460) );
  XNOR U7401 ( .A(n7531), .B(n7514), .Z(n7508) );
  XNOR U7402 ( .A(n7532), .B(n7533), .Z(n7514) );
  NOR U7403 ( .A(n7534), .B(n7535), .Z(n7533) );
  XOR U7404 ( .A(n7532), .B(n7536), .Z(n7534) );
  XNOR U7405 ( .A(n7513), .B(n7505), .Z(n7531) );
  XOR U7406 ( .A(n7537), .B(n7538), .Z(n7505) );
  AND U7407 ( .A(n7539), .B(n7540), .Z(n7538) );
  XOR U7408 ( .A(n7537), .B(n7541), .Z(n7539) );
  XNOR U7409 ( .A(n7542), .B(n7510), .Z(n7513) );
  XOR U7410 ( .A(n7543), .B(n7544), .Z(n7510) );
  AND U7411 ( .A(n7545), .B(n7546), .Z(n7544) );
  XNOR U7412 ( .A(n7547), .B(n7548), .Z(n7545) );
  IV U7413 ( .A(n7543), .Z(n7547) );
  XNOR U7414 ( .A(n7549), .B(n7550), .Z(n7542) );
  NOR U7415 ( .A(n7551), .B(n7552), .Z(n7550) );
  XNOR U7416 ( .A(n7549), .B(n7553), .Z(n7551) );
  XNOR U7417 ( .A(n7509), .B(n7516), .Z(n7530) );
  NOR U7418 ( .A(n7473), .B(n7554), .Z(n7516) );
  XOR U7419 ( .A(n7521), .B(n7520), .Z(n7509) );
  XNOR U7420 ( .A(n7555), .B(n7517), .Z(n7520) );
  XOR U7421 ( .A(n7556), .B(n7557), .Z(n7517) );
  AND U7422 ( .A(n7558), .B(n7559), .Z(n7557) );
  XNOR U7423 ( .A(n7560), .B(n7561), .Z(n7558) );
  IV U7424 ( .A(n7556), .Z(n7560) );
  XNOR U7425 ( .A(n7562), .B(n7563), .Z(n7555) );
  NOR U7426 ( .A(n7564), .B(n7565), .Z(n7563) );
  XNOR U7427 ( .A(n7562), .B(n7566), .Z(n7564) );
  XOR U7428 ( .A(n7567), .B(n7568), .Z(n7521) );
  NOR U7429 ( .A(n7569), .B(n7570), .Z(n7568) );
  XNOR U7430 ( .A(n7567), .B(n7571), .Z(n7569) );
  XNOR U7431 ( .A(n7457), .B(n7526), .Z(n7528) );
  XOR U7432 ( .A(n7572), .B(n7573), .Z(n7457) );
  AND U7433 ( .A(n51), .B(n7574), .Z(n7573) );
  XOR U7434 ( .A(n7575), .B(n7572), .Z(n7574) );
  AND U7435 ( .A(n7470), .B(n7473), .Z(n7526) );
  XOR U7436 ( .A(n7576), .B(n7554), .Z(n7473) );
  XNOR U7437 ( .A(p_input[176]), .B(p_input[2048]), .Z(n7554) );
  XNOR U7438 ( .A(n7541), .B(n7540), .Z(n7576) );
  XNOR U7439 ( .A(n7577), .B(n7548), .Z(n7540) );
  XNOR U7440 ( .A(n7536), .B(n7535), .Z(n7548) );
  XNOR U7441 ( .A(n7578), .B(n7532), .Z(n7535) );
  XNOR U7442 ( .A(p_input[186]), .B(p_input[2058]), .Z(n7532) );
  XOR U7443 ( .A(p_input[187]), .B(n6319), .Z(n7578) );
  XOR U7444 ( .A(p_input[188]), .B(p_input[2060]), .Z(n7536) );
  XOR U7445 ( .A(n7546), .B(n7579), .Z(n7577) );
  IV U7446 ( .A(n7537), .Z(n7579) );
  XOR U7447 ( .A(p_input[177]), .B(p_input[2049]), .Z(n7537) );
  XNOR U7448 ( .A(n7580), .B(n7553), .Z(n7546) );
  XNOR U7449 ( .A(p_input[191]), .B(n6322), .Z(n7553) );
  XOR U7450 ( .A(n7543), .B(n7552), .Z(n7580) );
  XOR U7451 ( .A(n7581), .B(n7549), .Z(n7552) );
  XOR U7452 ( .A(p_input[189]), .B(p_input[2061]), .Z(n7549) );
  XOR U7453 ( .A(p_input[190]), .B(n6324), .Z(n7581) );
  XOR U7454 ( .A(p_input[185]), .B(p_input[2057]), .Z(n7543) );
  XOR U7455 ( .A(n7561), .B(n7559), .Z(n7541) );
  XNOR U7456 ( .A(n7582), .B(n7566), .Z(n7559) );
  XOR U7457 ( .A(p_input[184]), .B(p_input[2056]), .Z(n7566) );
  XOR U7458 ( .A(n7556), .B(n7565), .Z(n7582) );
  XOR U7459 ( .A(n7583), .B(n7562), .Z(n7565) );
  XOR U7460 ( .A(p_input[182]), .B(p_input[2054]), .Z(n7562) );
  XOR U7461 ( .A(p_input[183]), .B(n7007), .Z(n7583) );
  XOR U7462 ( .A(p_input[178]), .B(p_input[2050]), .Z(n7556) );
  XNOR U7463 ( .A(n7571), .B(n7570), .Z(n7561) );
  XOR U7464 ( .A(n7584), .B(n7567), .Z(n7570) );
  XOR U7465 ( .A(p_input[179]), .B(p_input[2051]), .Z(n7567) );
  XOR U7466 ( .A(p_input[180]), .B(n7009), .Z(n7584) );
  XOR U7467 ( .A(p_input[181]), .B(p_input[2053]), .Z(n7571) );
  XOR U7468 ( .A(n7585), .B(n7586), .Z(n7470) );
  AND U7469 ( .A(n51), .B(n7587), .Z(n7586) );
  XNOR U7470 ( .A(n7588), .B(n7585), .Z(n7587) );
  XNOR U7471 ( .A(n7589), .B(n7590), .Z(n51) );
  AND U7472 ( .A(n7591), .B(n7592), .Z(n7590) );
  XOR U7473 ( .A(n7483), .B(n7589), .Z(n7592) );
  AND U7474 ( .A(n7593), .B(n7594), .Z(n7483) );
  XNOR U7475 ( .A(n7480), .B(n7589), .Z(n7591) );
  XOR U7476 ( .A(n7595), .B(n7596), .Z(n7480) );
  AND U7477 ( .A(n55), .B(n7597), .Z(n7596) );
  XOR U7478 ( .A(n7598), .B(n7595), .Z(n7597) );
  XOR U7479 ( .A(n7599), .B(n7600), .Z(n7589) );
  AND U7480 ( .A(n7601), .B(n7602), .Z(n7600) );
  XNOR U7481 ( .A(n7599), .B(n7593), .Z(n7602) );
  IV U7482 ( .A(n7498), .Z(n7593) );
  XOR U7483 ( .A(n7603), .B(n7604), .Z(n7498) );
  XOR U7484 ( .A(n7605), .B(n7594), .Z(n7604) );
  AND U7485 ( .A(n7525), .B(n7606), .Z(n7594) );
  AND U7486 ( .A(n7607), .B(n7608), .Z(n7605) );
  XOR U7487 ( .A(n7609), .B(n7603), .Z(n7607) );
  XNOR U7488 ( .A(n7495), .B(n7599), .Z(n7601) );
  XOR U7489 ( .A(n7610), .B(n7611), .Z(n7495) );
  AND U7490 ( .A(n55), .B(n7612), .Z(n7611) );
  XOR U7491 ( .A(n7613), .B(n7610), .Z(n7612) );
  XOR U7492 ( .A(n7614), .B(n7615), .Z(n7599) );
  AND U7493 ( .A(n7616), .B(n7617), .Z(n7615) );
  XNOR U7494 ( .A(n7614), .B(n7525), .Z(n7617) );
  XOR U7495 ( .A(n7618), .B(n7608), .Z(n7525) );
  XNOR U7496 ( .A(n7619), .B(n7603), .Z(n7608) );
  XOR U7497 ( .A(n7620), .B(n7621), .Z(n7603) );
  AND U7498 ( .A(n7622), .B(n7623), .Z(n7621) );
  XOR U7499 ( .A(n7624), .B(n7620), .Z(n7622) );
  XNOR U7500 ( .A(n7625), .B(n7626), .Z(n7619) );
  AND U7501 ( .A(n7627), .B(n7628), .Z(n7626) );
  XOR U7502 ( .A(n7625), .B(n7629), .Z(n7627) );
  XNOR U7503 ( .A(n7609), .B(n7606), .Z(n7618) );
  AND U7504 ( .A(n7630), .B(n7631), .Z(n7606) );
  XOR U7505 ( .A(n7632), .B(n7633), .Z(n7609) );
  AND U7506 ( .A(n7634), .B(n7635), .Z(n7633) );
  XOR U7507 ( .A(n7632), .B(n7636), .Z(n7634) );
  XNOR U7508 ( .A(n7522), .B(n7614), .Z(n7616) );
  XOR U7509 ( .A(n7637), .B(n7638), .Z(n7522) );
  AND U7510 ( .A(n55), .B(n7639), .Z(n7638) );
  XNOR U7511 ( .A(n7640), .B(n7637), .Z(n7639) );
  XOR U7512 ( .A(n7641), .B(n7642), .Z(n7614) );
  AND U7513 ( .A(n7643), .B(n7644), .Z(n7642) );
  XNOR U7514 ( .A(n7641), .B(n7630), .Z(n7644) );
  IV U7515 ( .A(n7575), .Z(n7630) );
  XNOR U7516 ( .A(n7645), .B(n7623), .Z(n7575) );
  XNOR U7517 ( .A(n7646), .B(n7629), .Z(n7623) );
  XNOR U7518 ( .A(n7647), .B(n7648), .Z(n7629) );
  NOR U7519 ( .A(n7649), .B(n7650), .Z(n7648) );
  XOR U7520 ( .A(n7647), .B(n7651), .Z(n7649) );
  XNOR U7521 ( .A(n7628), .B(n7620), .Z(n7646) );
  XOR U7522 ( .A(n7652), .B(n7653), .Z(n7620) );
  AND U7523 ( .A(n7654), .B(n7655), .Z(n7653) );
  XOR U7524 ( .A(n7652), .B(n7656), .Z(n7654) );
  XNOR U7525 ( .A(n7657), .B(n7625), .Z(n7628) );
  XOR U7526 ( .A(n7658), .B(n7659), .Z(n7625) );
  AND U7527 ( .A(n7660), .B(n7661), .Z(n7659) );
  XNOR U7528 ( .A(n7662), .B(n7663), .Z(n7660) );
  IV U7529 ( .A(n7658), .Z(n7662) );
  XNOR U7530 ( .A(n7664), .B(n7665), .Z(n7657) );
  NOR U7531 ( .A(n7666), .B(n7667), .Z(n7665) );
  XOR U7532 ( .A(n7664), .B(n7668), .Z(n7666) );
  XNOR U7533 ( .A(n7624), .B(n7631), .Z(n7645) );
  NOR U7534 ( .A(n7588), .B(n7669), .Z(n7631) );
  XOR U7535 ( .A(n7636), .B(n7635), .Z(n7624) );
  XNOR U7536 ( .A(n7670), .B(n7632), .Z(n7635) );
  XOR U7537 ( .A(n7671), .B(n7672), .Z(n7632) );
  AND U7538 ( .A(n7673), .B(n7674), .Z(n7672) );
  XNOR U7539 ( .A(n7675), .B(n7676), .Z(n7673) );
  IV U7540 ( .A(n7671), .Z(n7675) );
  XNOR U7541 ( .A(n7677), .B(n7678), .Z(n7670) );
  NOR U7542 ( .A(n7679), .B(n7680), .Z(n7678) );
  XNOR U7543 ( .A(n7677), .B(n7681), .Z(n7679) );
  XOR U7544 ( .A(n7682), .B(n7683), .Z(n7636) );
  NOR U7545 ( .A(n7684), .B(n7685), .Z(n7683) );
  XNOR U7546 ( .A(n7682), .B(n7686), .Z(n7684) );
  XNOR U7547 ( .A(n7572), .B(n7641), .Z(n7643) );
  XOR U7548 ( .A(n7687), .B(n7688), .Z(n7572) );
  AND U7549 ( .A(n55), .B(n7689), .Z(n7688) );
  XOR U7550 ( .A(n7690), .B(n7687), .Z(n7689) );
  AND U7551 ( .A(n7585), .B(n7588), .Z(n7641) );
  XOR U7552 ( .A(n7691), .B(n7669), .Z(n7588) );
  XNOR U7553 ( .A(p_input[192]), .B(p_input[2048]), .Z(n7669) );
  XNOR U7554 ( .A(n7656), .B(n7655), .Z(n7691) );
  XNOR U7555 ( .A(n7692), .B(n7663), .Z(n7655) );
  XNOR U7556 ( .A(n7651), .B(n7650), .Z(n7663) );
  XNOR U7557 ( .A(n7693), .B(n7647), .Z(n7650) );
  XNOR U7558 ( .A(p_input[202]), .B(p_input[2058]), .Z(n7647) );
  XOR U7559 ( .A(p_input[203]), .B(n6319), .Z(n7693) );
  XOR U7560 ( .A(p_input[204]), .B(p_input[2060]), .Z(n7651) );
  XOR U7561 ( .A(n7661), .B(n7694), .Z(n7692) );
  IV U7562 ( .A(n7652), .Z(n7694) );
  XOR U7563 ( .A(p_input[193]), .B(p_input[2049]), .Z(n7652) );
  XOR U7564 ( .A(n7695), .B(n7668), .Z(n7661) );
  XNOR U7565 ( .A(p_input[2063]), .B(p_input[207]), .Z(n7668) );
  XOR U7566 ( .A(n7658), .B(n7667), .Z(n7695) );
  XOR U7567 ( .A(n7696), .B(n7664), .Z(n7667) );
  XOR U7568 ( .A(p_input[205]), .B(p_input[2061]), .Z(n7664) );
  XNOR U7569 ( .A(p_input[2062]), .B(p_input[206]), .Z(n7696) );
  XOR U7570 ( .A(p_input[201]), .B(p_input[2057]), .Z(n7658) );
  XOR U7571 ( .A(n7676), .B(n7674), .Z(n7656) );
  XNOR U7572 ( .A(n7697), .B(n7681), .Z(n7674) );
  XOR U7573 ( .A(p_input[200]), .B(p_input[2056]), .Z(n7681) );
  XOR U7574 ( .A(n7671), .B(n7680), .Z(n7697) );
  XOR U7575 ( .A(n7698), .B(n7677), .Z(n7680) );
  XOR U7576 ( .A(p_input[198]), .B(p_input[2054]), .Z(n7677) );
  XOR U7577 ( .A(p_input[199]), .B(n7007), .Z(n7698) );
  XOR U7578 ( .A(p_input[194]), .B(p_input[2050]), .Z(n7671) );
  XNOR U7579 ( .A(n7686), .B(n7685), .Z(n7676) );
  XOR U7580 ( .A(n7699), .B(n7682), .Z(n7685) );
  XOR U7581 ( .A(p_input[195]), .B(p_input[2051]), .Z(n7682) );
  XOR U7582 ( .A(p_input[196]), .B(n7009), .Z(n7699) );
  XOR U7583 ( .A(p_input[197]), .B(p_input[2053]), .Z(n7686) );
  XOR U7584 ( .A(n7700), .B(n7701), .Z(n7585) );
  AND U7585 ( .A(n55), .B(n7702), .Z(n7701) );
  XNOR U7586 ( .A(n7703), .B(n7700), .Z(n7702) );
  XNOR U7587 ( .A(n7704), .B(n7705), .Z(n55) );
  AND U7588 ( .A(n7706), .B(n7707), .Z(n7705) );
  XOR U7589 ( .A(n7598), .B(n7704), .Z(n7707) );
  AND U7590 ( .A(n7708), .B(n7709), .Z(n7598) );
  XNOR U7591 ( .A(n7595), .B(n7704), .Z(n7706) );
  XOR U7592 ( .A(n7710), .B(n7711), .Z(n7595) );
  AND U7593 ( .A(n59), .B(n7712), .Z(n7711) );
  XOR U7594 ( .A(n7713), .B(n7710), .Z(n7712) );
  XOR U7595 ( .A(n7714), .B(n7715), .Z(n7704) );
  AND U7596 ( .A(n7716), .B(n7717), .Z(n7715) );
  XNOR U7597 ( .A(n7714), .B(n7708), .Z(n7717) );
  IV U7598 ( .A(n7613), .Z(n7708) );
  XOR U7599 ( .A(n7718), .B(n7719), .Z(n7613) );
  XOR U7600 ( .A(n7720), .B(n7709), .Z(n7719) );
  AND U7601 ( .A(n7640), .B(n7721), .Z(n7709) );
  AND U7602 ( .A(n7722), .B(n7723), .Z(n7720) );
  XOR U7603 ( .A(n7724), .B(n7718), .Z(n7722) );
  XNOR U7604 ( .A(n7610), .B(n7714), .Z(n7716) );
  XOR U7605 ( .A(n7725), .B(n7726), .Z(n7610) );
  AND U7606 ( .A(n59), .B(n7727), .Z(n7726) );
  XOR U7607 ( .A(n7728), .B(n7725), .Z(n7727) );
  XOR U7608 ( .A(n7729), .B(n7730), .Z(n7714) );
  AND U7609 ( .A(n7731), .B(n7732), .Z(n7730) );
  XNOR U7610 ( .A(n7729), .B(n7640), .Z(n7732) );
  XOR U7611 ( .A(n7733), .B(n7723), .Z(n7640) );
  XNOR U7612 ( .A(n7734), .B(n7718), .Z(n7723) );
  XOR U7613 ( .A(n7735), .B(n7736), .Z(n7718) );
  AND U7614 ( .A(n7737), .B(n7738), .Z(n7736) );
  XOR U7615 ( .A(n7739), .B(n7735), .Z(n7737) );
  XNOR U7616 ( .A(n7740), .B(n7741), .Z(n7734) );
  AND U7617 ( .A(n7742), .B(n7743), .Z(n7741) );
  XOR U7618 ( .A(n7740), .B(n7744), .Z(n7742) );
  XNOR U7619 ( .A(n7724), .B(n7721), .Z(n7733) );
  AND U7620 ( .A(n7745), .B(n7746), .Z(n7721) );
  XOR U7621 ( .A(n7747), .B(n7748), .Z(n7724) );
  AND U7622 ( .A(n7749), .B(n7750), .Z(n7748) );
  XOR U7623 ( .A(n7747), .B(n7751), .Z(n7749) );
  XNOR U7624 ( .A(n7637), .B(n7729), .Z(n7731) );
  XOR U7625 ( .A(n7752), .B(n7753), .Z(n7637) );
  AND U7626 ( .A(n59), .B(n7754), .Z(n7753) );
  XNOR U7627 ( .A(n7755), .B(n7752), .Z(n7754) );
  XOR U7628 ( .A(n7756), .B(n7757), .Z(n7729) );
  AND U7629 ( .A(n7758), .B(n7759), .Z(n7757) );
  XNOR U7630 ( .A(n7756), .B(n7745), .Z(n7759) );
  IV U7631 ( .A(n7690), .Z(n7745) );
  XNOR U7632 ( .A(n7760), .B(n7738), .Z(n7690) );
  XNOR U7633 ( .A(n7761), .B(n7744), .Z(n7738) );
  XOR U7634 ( .A(n7762), .B(n7763), .Z(n7744) );
  NOR U7635 ( .A(n7764), .B(n7765), .Z(n7763) );
  XNOR U7636 ( .A(n7762), .B(n7766), .Z(n7764) );
  XNOR U7637 ( .A(n7743), .B(n7735), .Z(n7761) );
  XOR U7638 ( .A(n7767), .B(n7768), .Z(n7735) );
  AND U7639 ( .A(n7769), .B(n7770), .Z(n7768) );
  XNOR U7640 ( .A(n7767), .B(n7771), .Z(n7769) );
  XNOR U7641 ( .A(n7772), .B(n7740), .Z(n7743) );
  XOR U7642 ( .A(n7773), .B(n7774), .Z(n7740) );
  AND U7643 ( .A(n7775), .B(n7776), .Z(n7774) );
  XOR U7644 ( .A(n7773), .B(n7777), .Z(n7775) );
  XNOR U7645 ( .A(n7778), .B(n7779), .Z(n7772) );
  NOR U7646 ( .A(n7780), .B(n7781), .Z(n7779) );
  XOR U7647 ( .A(n7778), .B(n7782), .Z(n7780) );
  XNOR U7648 ( .A(n7739), .B(n7746), .Z(n7760) );
  NOR U7649 ( .A(n7703), .B(n7783), .Z(n7746) );
  XOR U7650 ( .A(n7751), .B(n7750), .Z(n7739) );
  XNOR U7651 ( .A(n7784), .B(n7747), .Z(n7750) );
  XOR U7652 ( .A(n7785), .B(n7786), .Z(n7747) );
  AND U7653 ( .A(n7787), .B(n7788), .Z(n7786) );
  XOR U7654 ( .A(n7785), .B(n7789), .Z(n7787) );
  XNOR U7655 ( .A(n7790), .B(n7791), .Z(n7784) );
  NOR U7656 ( .A(n7792), .B(n7793), .Z(n7791) );
  XNOR U7657 ( .A(n7790), .B(n7794), .Z(n7792) );
  XOR U7658 ( .A(n7795), .B(n7796), .Z(n7751) );
  NOR U7659 ( .A(n7797), .B(n7798), .Z(n7796) );
  XNOR U7660 ( .A(n7795), .B(n7799), .Z(n7797) );
  XNOR U7661 ( .A(n7687), .B(n7756), .Z(n7758) );
  XOR U7662 ( .A(n7800), .B(n7801), .Z(n7687) );
  AND U7663 ( .A(n59), .B(n7802), .Z(n7801) );
  XOR U7664 ( .A(n7803), .B(n7800), .Z(n7802) );
  AND U7665 ( .A(n7700), .B(n7703), .Z(n7756) );
  XOR U7666 ( .A(n7804), .B(n7783), .Z(n7703) );
  XNOR U7667 ( .A(p_input[2048]), .B(p_input[208]), .Z(n7783) );
  XOR U7668 ( .A(n7771), .B(n7770), .Z(n7804) );
  XNOR U7669 ( .A(n7805), .B(n7777), .Z(n7770) );
  XNOR U7670 ( .A(n7766), .B(n7765), .Z(n7777) );
  XOR U7671 ( .A(n7806), .B(n7762), .Z(n7765) );
  XNOR U7672 ( .A(n6439), .B(p_input[218]), .Z(n7762) );
  XNOR U7673 ( .A(p_input[2059]), .B(p_input[219]), .Z(n7806) );
  XOR U7674 ( .A(p_input[2060]), .B(p_input[220]), .Z(n7766) );
  XNOR U7675 ( .A(n7776), .B(n7767), .Z(n7805) );
  XNOR U7676 ( .A(n6553), .B(p_input[209]), .Z(n7767) );
  XOR U7677 ( .A(n7807), .B(n7782), .Z(n7776) );
  XNOR U7678 ( .A(p_input[2063]), .B(p_input[223]), .Z(n7782) );
  XOR U7679 ( .A(n7773), .B(n7781), .Z(n7807) );
  XOR U7680 ( .A(n7808), .B(n7778), .Z(n7781) );
  XOR U7681 ( .A(p_input[2061]), .B(p_input[221]), .Z(n7778) );
  XNOR U7682 ( .A(p_input[2062]), .B(p_input[222]), .Z(n7808) );
  XNOR U7683 ( .A(n6325), .B(p_input[217]), .Z(n7773) );
  XNOR U7684 ( .A(n7789), .B(n7788), .Z(n7771) );
  XNOR U7685 ( .A(n7809), .B(n7794), .Z(n7788) );
  XOR U7686 ( .A(p_input[2056]), .B(p_input[216]), .Z(n7794) );
  XOR U7687 ( .A(n7785), .B(n7793), .Z(n7809) );
  XOR U7688 ( .A(n7810), .B(n7790), .Z(n7793) );
  XOR U7689 ( .A(p_input[2054]), .B(p_input[214]), .Z(n7790) );
  XNOR U7690 ( .A(p_input[2055]), .B(p_input[215]), .Z(n7810) );
  XNOR U7691 ( .A(n6328), .B(p_input[210]), .Z(n7785) );
  XNOR U7692 ( .A(n7799), .B(n7798), .Z(n7789) );
  XOR U7693 ( .A(n7811), .B(n7795), .Z(n7798) );
  XOR U7694 ( .A(p_input[2051]), .B(p_input[211]), .Z(n7795) );
  XNOR U7695 ( .A(p_input[2052]), .B(p_input[212]), .Z(n7811) );
  XOR U7696 ( .A(p_input[2053]), .B(p_input[213]), .Z(n7799) );
  XOR U7697 ( .A(n7812), .B(n7813), .Z(n7700) );
  AND U7698 ( .A(n59), .B(n7814), .Z(n7813) );
  XNOR U7699 ( .A(n7815), .B(n7812), .Z(n7814) );
  XNOR U7700 ( .A(n7816), .B(n7817), .Z(n59) );
  AND U7701 ( .A(n7818), .B(n7819), .Z(n7817) );
  XOR U7702 ( .A(n7713), .B(n7816), .Z(n7819) );
  AND U7703 ( .A(n7820), .B(n7821), .Z(n7713) );
  XNOR U7704 ( .A(n7710), .B(n7816), .Z(n7818) );
  XOR U7705 ( .A(n7822), .B(n7823), .Z(n7710) );
  AND U7706 ( .A(n63), .B(n7824), .Z(n7823) );
  XOR U7707 ( .A(n7825), .B(n7822), .Z(n7824) );
  XOR U7708 ( .A(n7826), .B(n7827), .Z(n7816) );
  AND U7709 ( .A(n7828), .B(n7829), .Z(n7827) );
  XNOR U7710 ( .A(n7826), .B(n7820), .Z(n7829) );
  IV U7711 ( .A(n7728), .Z(n7820) );
  XOR U7712 ( .A(n7830), .B(n7831), .Z(n7728) );
  XOR U7713 ( .A(n7832), .B(n7821), .Z(n7831) );
  AND U7714 ( .A(n7755), .B(n7833), .Z(n7821) );
  AND U7715 ( .A(n7834), .B(n7835), .Z(n7832) );
  XOR U7716 ( .A(n7836), .B(n7830), .Z(n7834) );
  XNOR U7717 ( .A(n7725), .B(n7826), .Z(n7828) );
  XOR U7718 ( .A(n7837), .B(n7838), .Z(n7725) );
  AND U7719 ( .A(n63), .B(n7839), .Z(n7838) );
  XOR U7720 ( .A(n7840), .B(n7837), .Z(n7839) );
  XOR U7721 ( .A(n7841), .B(n7842), .Z(n7826) );
  AND U7722 ( .A(n7843), .B(n7844), .Z(n7842) );
  XNOR U7723 ( .A(n7841), .B(n7755), .Z(n7844) );
  XOR U7724 ( .A(n7845), .B(n7835), .Z(n7755) );
  XNOR U7725 ( .A(n7846), .B(n7830), .Z(n7835) );
  XOR U7726 ( .A(n7847), .B(n7848), .Z(n7830) );
  AND U7727 ( .A(n7849), .B(n7850), .Z(n7848) );
  XOR U7728 ( .A(n7851), .B(n7847), .Z(n7849) );
  XNOR U7729 ( .A(n7852), .B(n7853), .Z(n7846) );
  AND U7730 ( .A(n7854), .B(n7855), .Z(n7853) );
  XOR U7731 ( .A(n7852), .B(n7856), .Z(n7854) );
  XNOR U7732 ( .A(n7836), .B(n7833), .Z(n7845) );
  AND U7733 ( .A(n7857), .B(n7858), .Z(n7833) );
  XOR U7734 ( .A(n7859), .B(n7860), .Z(n7836) );
  AND U7735 ( .A(n7861), .B(n7862), .Z(n7860) );
  XOR U7736 ( .A(n7859), .B(n7863), .Z(n7861) );
  XNOR U7737 ( .A(n7752), .B(n7841), .Z(n7843) );
  XOR U7738 ( .A(n7864), .B(n7865), .Z(n7752) );
  AND U7739 ( .A(n63), .B(n7866), .Z(n7865) );
  XNOR U7740 ( .A(n7867), .B(n7864), .Z(n7866) );
  XOR U7741 ( .A(n7868), .B(n7869), .Z(n7841) );
  AND U7742 ( .A(n7870), .B(n7871), .Z(n7869) );
  XNOR U7743 ( .A(n7868), .B(n7857), .Z(n7871) );
  IV U7744 ( .A(n7803), .Z(n7857) );
  XNOR U7745 ( .A(n7872), .B(n7850), .Z(n7803) );
  XNOR U7746 ( .A(n7873), .B(n7856), .Z(n7850) );
  XOR U7747 ( .A(n7874), .B(n7875), .Z(n7856) );
  NOR U7748 ( .A(n7876), .B(n7877), .Z(n7875) );
  XNOR U7749 ( .A(n7874), .B(n7878), .Z(n7876) );
  XNOR U7750 ( .A(n7855), .B(n7847), .Z(n7873) );
  XOR U7751 ( .A(n7879), .B(n7880), .Z(n7847) );
  AND U7752 ( .A(n7881), .B(n7882), .Z(n7880) );
  XNOR U7753 ( .A(n7879), .B(n7883), .Z(n7881) );
  XNOR U7754 ( .A(n7884), .B(n7852), .Z(n7855) );
  XOR U7755 ( .A(n7885), .B(n7886), .Z(n7852) );
  AND U7756 ( .A(n7887), .B(n7888), .Z(n7886) );
  XOR U7757 ( .A(n7885), .B(n7889), .Z(n7887) );
  XNOR U7758 ( .A(n7890), .B(n7891), .Z(n7884) );
  NOR U7759 ( .A(n7892), .B(n7893), .Z(n7891) );
  XOR U7760 ( .A(n7890), .B(n7894), .Z(n7892) );
  XNOR U7761 ( .A(n7851), .B(n7858), .Z(n7872) );
  NOR U7762 ( .A(n7815), .B(n7895), .Z(n7858) );
  XOR U7763 ( .A(n7863), .B(n7862), .Z(n7851) );
  XNOR U7764 ( .A(n7896), .B(n7859), .Z(n7862) );
  XOR U7765 ( .A(n7897), .B(n7898), .Z(n7859) );
  AND U7766 ( .A(n7899), .B(n7900), .Z(n7898) );
  XOR U7767 ( .A(n7897), .B(n7901), .Z(n7899) );
  XNOR U7768 ( .A(n7902), .B(n7903), .Z(n7896) );
  NOR U7769 ( .A(n7904), .B(n7905), .Z(n7903) );
  XNOR U7770 ( .A(n7902), .B(n7906), .Z(n7904) );
  XOR U7771 ( .A(n7907), .B(n7908), .Z(n7863) );
  NOR U7772 ( .A(n7909), .B(n7910), .Z(n7908) );
  XNOR U7773 ( .A(n7907), .B(n7911), .Z(n7909) );
  XNOR U7774 ( .A(n7800), .B(n7868), .Z(n7870) );
  XOR U7775 ( .A(n7912), .B(n7913), .Z(n7800) );
  AND U7776 ( .A(n63), .B(n7914), .Z(n7913) );
  XOR U7777 ( .A(n7915), .B(n7912), .Z(n7914) );
  AND U7778 ( .A(n7812), .B(n7815), .Z(n7868) );
  XOR U7779 ( .A(n7916), .B(n7895), .Z(n7815) );
  XNOR U7780 ( .A(p_input[2048]), .B(p_input[224]), .Z(n7895) );
  XOR U7781 ( .A(n7883), .B(n7882), .Z(n7916) );
  XNOR U7782 ( .A(n7917), .B(n7889), .Z(n7882) );
  XNOR U7783 ( .A(n7878), .B(n7877), .Z(n7889) );
  XOR U7784 ( .A(n7918), .B(n7874), .Z(n7877) );
  XNOR U7785 ( .A(n6439), .B(p_input[234]), .Z(n7874) );
  XNOR U7786 ( .A(p_input[2059]), .B(p_input[235]), .Z(n7918) );
  XOR U7787 ( .A(p_input[2060]), .B(p_input[236]), .Z(n7878) );
  XNOR U7788 ( .A(n7888), .B(n7879), .Z(n7917) );
  XNOR U7789 ( .A(n6553), .B(p_input[225]), .Z(n7879) );
  XOR U7790 ( .A(n7919), .B(n7894), .Z(n7888) );
  XNOR U7791 ( .A(p_input[2063]), .B(p_input[239]), .Z(n7894) );
  XOR U7792 ( .A(n7885), .B(n7893), .Z(n7919) );
  XOR U7793 ( .A(n7920), .B(n7890), .Z(n7893) );
  XOR U7794 ( .A(p_input[2061]), .B(p_input[237]), .Z(n7890) );
  XNOR U7795 ( .A(p_input[2062]), .B(p_input[238]), .Z(n7920) );
  XNOR U7796 ( .A(n6325), .B(p_input[233]), .Z(n7885) );
  XNOR U7797 ( .A(n7901), .B(n7900), .Z(n7883) );
  XNOR U7798 ( .A(n7921), .B(n7906), .Z(n7900) );
  XOR U7799 ( .A(p_input[2056]), .B(p_input[232]), .Z(n7906) );
  XOR U7800 ( .A(n7897), .B(n7905), .Z(n7921) );
  XOR U7801 ( .A(n7922), .B(n7902), .Z(n7905) );
  XOR U7802 ( .A(p_input[2054]), .B(p_input[230]), .Z(n7902) );
  XNOR U7803 ( .A(p_input[2055]), .B(p_input[231]), .Z(n7922) );
  XNOR U7804 ( .A(n6328), .B(p_input[226]), .Z(n7897) );
  XNOR U7805 ( .A(n7911), .B(n7910), .Z(n7901) );
  XOR U7806 ( .A(n7923), .B(n7907), .Z(n7910) );
  XOR U7807 ( .A(p_input[2051]), .B(p_input[227]), .Z(n7907) );
  XNOR U7808 ( .A(p_input[2052]), .B(p_input[228]), .Z(n7923) );
  XOR U7809 ( .A(p_input[2053]), .B(p_input[229]), .Z(n7911) );
  XOR U7810 ( .A(n7924), .B(n7925), .Z(n7812) );
  AND U7811 ( .A(n63), .B(n7926), .Z(n7925) );
  XNOR U7812 ( .A(n7927), .B(n7924), .Z(n7926) );
  XNOR U7813 ( .A(n7928), .B(n7929), .Z(n63) );
  AND U7814 ( .A(n7930), .B(n7931), .Z(n7929) );
  XOR U7815 ( .A(n7825), .B(n7928), .Z(n7931) );
  AND U7816 ( .A(n7932), .B(n7933), .Z(n7825) );
  XNOR U7817 ( .A(n7822), .B(n7928), .Z(n7930) );
  XOR U7818 ( .A(n7934), .B(n7935), .Z(n7822) );
  AND U7819 ( .A(n67), .B(n7936), .Z(n7935) );
  XOR U7820 ( .A(n7937), .B(n7934), .Z(n7936) );
  XOR U7821 ( .A(n7938), .B(n7939), .Z(n7928) );
  AND U7822 ( .A(n7940), .B(n7941), .Z(n7939) );
  XNOR U7823 ( .A(n7938), .B(n7932), .Z(n7941) );
  IV U7824 ( .A(n7840), .Z(n7932) );
  XOR U7825 ( .A(n7942), .B(n7943), .Z(n7840) );
  XOR U7826 ( .A(n7944), .B(n7933), .Z(n7943) );
  AND U7827 ( .A(n7867), .B(n7945), .Z(n7933) );
  AND U7828 ( .A(n7946), .B(n7947), .Z(n7944) );
  XOR U7829 ( .A(n7948), .B(n7942), .Z(n7946) );
  XNOR U7830 ( .A(n7837), .B(n7938), .Z(n7940) );
  XOR U7831 ( .A(n7949), .B(n7950), .Z(n7837) );
  AND U7832 ( .A(n67), .B(n7951), .Z(n7950) );
  XOR U7833 ( .A(n7952), .B(n7949), .Z(n7951) );
  XOR U7834 ( .A(n7953), .B(n7954), .Z(n7938) );
  AND U7835 ( .A(n7955), .B(n7956), .Z(n7954) );
  XNOR U7836 ( .A(n7953), .B(n7867), .Z(n7956) );
  XOR U7837 ( .A(n7957), .B(n7947), .Z(n7867) );
  XNOR U7838 ( .A(n7958), .B(n7942), .Z(n7947) );
  XOR U7839 ( .A(n7959), .B(n7960), .Z(n7942) );
  AND U7840 ( .A(n7961), .B(n7962), .Z(n7960) );
  XOR U7841 ( .A(n7963), .B(n7959), .Z(n7961) );
  XNOR U7842 ( .A(n7964), .B(n7965), .Z(n7958) );
  AND U7843 ( .A(n7966), .B(n7967), .Z(n7965) );
  XOR U7844 ( .A(n7964), .B(n7968), .Z(n7966) );
  XNOR U7845 ( .A(n7948), .B(n7945), .Z(n7957) );
  AND U7846 ( .A(n7969), .B(n7970), .Z(n7945) );
  XOR U7847 ( .A(n7971), .B(n7972), .Z(n7948) );
  AND U7848 ( .A(n7973), .B(n7974), .Z(n7972) );
  XOR U7849 ( .A(n7971), .B(n7975), .Z(n7973) );
  XNOR U7850 ( .A(n7864), .B(n7953), .Z(n7955) );
  XOR U7851 ( .A(n7976), .B(n7977), .Z(n7864) );
  AND U7852 ( .A(n67), .B(n7978), .Z(n7977) );
  XNOR U7853 ( .A(n7979), .B(n7976), .Z(n7978) );
  XOR U7854 ( .A(n7980), .B(n7981), .Z(n7953) );
  AND U7855 ( .A(n7982), .B(n7983), .Z(n7981) );
  XNOR U7856 ( .A(n7980), .B(n7969), .Z(n7983) );
  IV U7857 ( .A(n7915), .Z(n7969) );
  XNOR U7858 ( .A(n7984), .B(n7962), .Z(n7915) );
  XNOR U7859 ( .A(n7985), .B(n7968), .Z(n7962) );
  XOR U7860 ( .A(n7986), .B(n7987), .Z(n7968) );
  NOR U7861 ( .A(n7988), .B(n7989), .Z(n7987) );
  XNOR U7862 ( .A(n7986), .B(n7990), .Z(n7988) );
  XNOR U7863 ( .A(n7967), .B(n7959), .Z(n7985) );
  XOR U7864 ( .A(n7991), .B(n7992), .Z(n7959) );
  AND U7865 ( .A(n7993), .B(n7994), .Z(n7992) );
  XNOR U7866 ( .A(n7991), .B(n7995), .Z(n7993) );
  XNOR U7867 ( .A(n7996), .B(n7964), .Z(n7967) );
  XOR U7868 ( .A(n7997), .B(n7998), .Z(n7964) );
  AND U7869 ( .A(n7999), .B(n8000), .Z(n7998) );
  XOR U7870 ( .A(n7997), .B(n8001), .Z(n7999) );
  XNOR U7871 ( .A(n8002), .B(n8003), .Z(n7996) );
  NOR U7872 ( .A(n8004), .B(n8005), .Z(n8003) );
  XOR U7873 ( .A(n8002), .B(n8006), .Z(n8004) );
  XNOR U7874 ( .A(n7963), .B(n7970), .Z(n7984) );
  NOR U7875 ( .A(n7927), .B(n8007), .Z(n7970) );
  XOR U7876 ( .A(n7975), .B(n7974), .Z(n7963) );
  XNOR U7877 ( .A(n8008), .B(n7971), .Z(n7974) );
  XOR U7878 ( .A(n8009), .B(n8010), .Z(n7971) );
  AND U7879 ( .A(n8011), .B(n8012), .Z(n8010) );
  XOR U7880 ( .A(n8009), .B(n8013), .Z(n8011) );
  XNOR U7881 ( .A(n8014), .B(n8015), .Z(n8008) );
  NOR U7882 ( .A(n8016), .B(n8017), .Z(n8015) );
  XNOR U7883 ( .A(n8014), .B(n8018), .Z(n8016) );
  XOR U7884 ( .A(n8019), .B(n8020), .Z(n7975) );
  NOR U7885 ( .A(n8021), .B(n8022), .Z(n8020) );
  XNOR U7886 ( .A(n8019), .B(n8023), .Z(n8021) );
  XNOR U7887 ( .A(n7912), .B(n7980), .Z(n7982) );
  XOR U7888 ( .A(n8024), .B(n8025), .Z(n7912) );
  AND U7889 ( .A(n67), .B(n8026), .Z(n8025) );
  XOR U7890 ( .A(n8027), .B(n8024), .Z(n8026) );
  AND U7891 ( .A(n7924), .B(n7927), .Z(n7980) );
  XOR U7892 ( .A(n8028), .B(n8007), .Z(n7927) );
  XNOR U7893 ( .A(p_input[2048]), .B(p_input[240]), .Z(n8007) );
  XOR U7894 ( .A(n7995), .B(n7994), .Z(n8028) );
  XNOR U7895 ( .A(n8029), .B(n8001), .Z(n7994) );
  XNOR U7896 ( .A(n7990), .B(n7989), .Z(n8001) );
  XOR U7897 ( .A(n8030), .B(n7986), .Z(n7989) );
  XNOR U7898 ( .A(n6439), .B(p_input[250]), .Z(n7986) );
  XNOR U7899 ( .A(p_input[2059]), .B(p_input[251]), .Z(n8030) );
  XOR U7900 ( .A(p_input[2060]), .B(p_input[252]), .Z(n7990) );
  XNOR U7901 ( .A(n8000), .B(n7991), .Z(n8029) );
  XNOR U7902 ( .A(n6553), .B(p_input[241]), .Z(n7991) );
  XOR U7903 ( .A(n8031), .B(n8006), .Z(n8000) );
  XNOR U7904 ( .A(p_input[2063]), .B(p_input[255]), .Z(n8006) );
  XOR U7905 ( .A(n7997), .B(n8005), .Z(n8031) );
  XOR U7906 ( .A(n8032), .B(n8002), .Z(n8005) );
  XOR U7907 ( .A(p_input[2061]), .B(p_input[253]), .Z(n8002) );
  XNOR U7908 ( .A(p_input[2062]), .B(p_input[254]), .Z(n8032) );
  XNOR U7909 ( .A(n6325), .B(p_input[249]), .Z(n7997) );
  XNOR U7910 ( .A(n8013), .B(n8012), .Z(n7995) );
  XNOR U7911 ( .A(n8033), .B(n8018), .Z(n8012) );
  XOR U7912 ( .A(p_input[2056]), .B(p_input[248]), .Z(n8018) );
  XOR U7913 ( .A(n8009), .B(n8017), .Z(n8033) );
  XOR U7914 ( .A(n8034), .B(n8014), .Z(n8017) );
  XOR U7915 ( .A(p_input[2054]), .B(p_input[246]), .Z(n8014) );
  XNOR U7916 ( .A(p_input[2055]), .B(p_input[247]), .Z(n8034) );
  XNOR U7917 ( .A(n6328), .B(p_input[242]), .Z(n8009) );
  XNOR U7918 ( .A(n8023), .B(n8022), .Z(n8013) );
  XOR U7919 ( .A(n8035), .B(n8019), .Z(n8022) );
  XOR U7920 ( .A(p_input[2051]), .B(p_input[243]), .Z(n8019) );
  XNOR U7921 ( .A(p_input[2052]), .B(p_input[244]), .Z(n8035) );
  XOR U7922 ( .A(p_input[2053]), .B(p_input[245]), .Z(n8023) );
  XOR U7923 ( .A(n8036), .B(n8037), .Z(n7924) );
  AND U7924 ( .A(n67), .B(n8038), .Z(n8037) );
  XNOR U7925 ( .A(n8039), .B(n8036), .Z(n8038) );
  XNOR U7926 ( .A(n8040), .B(n8041), .Z(n67) );
  AND U7927 ( .A(n8042), .B(n8043), .Z(n8041) );
  XOR U7928 ( .A(n7937), .B(n8040), .Z(n8043) );
  AND U7929 ( .A(n8044), .B(n8045), .Z(n7937) );
  XNOR U7930 ( .A(n7934), .B(n8040), .Z(n8042) );
  XOR U7931 ( .A(n8046), .B(n8047), .Z(n7934) );
  AND U7932 ( .A(n71), .B(n8048), .Z(n8047) );
  XOR U7933 ( .A(n8049), .B(n8046), .Z(n8048) );
  XOR U7934 ( .A(n8050), .B(n8051), .Z(n8040) );
  AND U7935 ( .A(n8052), .B(n8053), .Z(n8051) );
  XNOR U7936 ( .A(n8050), .B(n8044), .Z(n8053) );
  IV U7937 ( .A(n7952), .Z(n8044) );
  XOR U7938 ( .A(n8054), .B(n8055), .Z(n7952) );
  XOR U7939 ( .A(n8056), .B(n8045), .Z(n8055) );
  AND U7940 ( .A(n7979), .B(n8057), .Z(n8045) );
  AND U7941 ( .A(n8058), .B(n8059), .Z(n8056) );
  XOR U7942 ( .A(n8060), .B(n8054), .Z(n8058) );
  XNOR U7943 ( .A(n7949), .B(n8050), .Z(n8052) );
  XOR U7944 ( .A(n8061), .B(n8062), .Z(n7949) );
  AND U7945 ( .A(n71), .B(n8063), .Z(n8062) );
  XOR U7946 ( .A(n8064), .B(n8061), .Z(n8063) );
  XOR U7947 ( .A(n8065), .B(n8066), .Z(n8050) );
  AND U7948 ( .A(n8067), .B(n8068), .Z(n8066) );
  XNOR U7949 ( .A(n8065), .B(n7979), .Z(n8068) );
  XOR U7950 ( .A(n8069), .B(n8059), .Z(n7979) );
  XNOR U7951 ( .A(n8070), .B(n8054), .Z(n8059) );
  XOR U7952 ( .A(n8071), .B(n8072), .Z(n8054) );
  AND U7953 ( .A(n8073), .B(n8074), .Z(n8072) );
  XOR U7954 ( .A(n8075), .B(n8071), .Z(n8073) );
  XNOR U7955 ( .A(n8076), .B(n8077), .Z(n8070) );
  AND U7956 ( .A(n8078), .B(n8079), .Z(n8077) );
  XOR U7957 ( .A(n8076), .B(n8080), .Z(n8078) );
  XNOR U7958 ( .A(n8060), .B(n8057), .Z(n8069) );
  AND U7959 ( .A(n8081), .B(n8082), .Z(n8057) );
  XOR U7960 ( .A(n8083), .B(n8084), .Z(n8060) );
  AND U7961 ( .A(n8085), .B(n8086), .Z(n8084) );
  XOR U7962 ( .A(n8083), .B(n8087), .Z(n8085) );
  XNOR U7963 ( .A(n7976), .B(n8065), .Z(n8067) );
  XOR U7964 ( .A(n8088), .B(n8089), .Z(n7976) );
  AND U7965 ( .A(n71), .B(n8090), .Z(n8089) );
  XNOR U7966 ( .A(n8091), .B(n8088), .Z(n8090) );
  XOR U7967 ( .A(n8092), .B(n8093), .Z(n8065) );
  AND U7968 ( .A(n8094), .B(n8095), .Z(n8093) );
  XNOR U7969 ( .A(n8092), .B(n8081), .Z(n8095) );
  IV U7970 ( .A(n8027), .Z(n8081) );
  XNOR U7971 ( .A(n8096), .B(n8074), .Z(n8027) );
  XNOR U7972 ( .A(n8097), .B(n8080), .Z(n8074) );
  XOR U7973 ( .A(n8098), .B(n8099), .Z(n8080) );
  NOR U7974 ( .A(n8100), .B(n8101), .Z(n8099) );
  XNOR U7975 ( .A(n8098), .B(n8102), .Z(n8100) );
  XNOR U7976 ( .A(n8079), .B(n8071), .Z(n8097) );
  XOR U7977 ( .A(n8103), .B(n8104), .Z(n8071) );
  AND U7978 ( .A(n8105), .B(n8106), .Z(n8104) );
  XNOR U7979 ( .A(n8103), .B(n8107), .Z(n8105) );
  XNOR U7980 ( .A(n8108), .B(n8076), .Z(n8079) );
  XOR U7981 ( .A(n8109), .B(n8110), .Z(n8076) );
  AND U7982 ( .A(n8111), .B(n8112), .Z(n8110) );
  XOR U7983 ( .A(n8109), .B(n8113), .Z(n8111) );
  XNOR U7984 ( .A(n8114), .B(n8115), .Z(n8108) );
  NOR U7985 ( .A(n8116), .B(n8117), .Z(n8115) );
  XOR U7986 ( .A(n8114), .B(n8118), .Z(n8116) );
  XNOR U7987 ( .A(n8075), .B(n8082), .Z(n8096) );
  NOR U7988 ( .A(n8039), .B(n8119), .Z(n8082) );
  XOR U7989 ( .A(n8087), .B(n8086), .Z(n8075) );
  XNOR U7990 ( .A(n8120), .B(n8083), .Z(n8086) );
  XOR U7991 ( .A(n8121), .B(n8122), .Z(n8083) );
  AND U7992 ( .A(n8123), .B(n8124), .Z(n8122) );
  XOR U7993 ( .A(n8121), .B(n8125), .Z(n8123) );
  XNOR U7994 ( .A(n8126), .B(n8127), .Z(n8120) );
  NOR U7995 ( .A(n8128), .B(n8129), .Z(n8127) );
  XNOR U7996 ( .A(n8126), .B(n8130), .Z(n8128) );
  XOR U7997 ( .A(n8131), .B(n8132), .Z(n8087) );
  NOR U7998 ( .A(n8133), .B(n8134), .Z(n8132) );
  XNOR U7999 ( .A(n8131), .B(n8135), .Z(n8133) );
  XNOR U8000 ( .A(n8024), .B(n8092), .Z(n8094) );
  XOR U8001 ( .A(n8136), .B(n8137), .Z(n8024) );
  AND U8002 ( .A(n71), .B(n8138), .Z(n8137) );
  XOR U8003 ( .A(n8139), .B(n8136), .Z(n8138) );
  AND U8004 ( .A(n8036), .B(n8039), .Z(n8092) );
  XOR U8005 ( .A(n8140), .B(n8119), .Z(n8039) );
  XNOR U8006 ( .A(p_input[2048]), .B(p_input[256]), .Z(n8119) );
  XOR U8007 ( .A(n8107), .B(n8106), .Z(n8140) );
  XNOR U8008 ( .A(n8141), .B(n8113), .Z(n8106) );
  XNOR U8009 ( .A(n8102), .B(n8101), .Z(n8113) );
  XOR U8010 ( .A(n8142), .B(n8098), .Z(n8101) );
  XNOR U8011 ( .A(n6439), .B(p_input[266]), .Z(n8098) );
  XNOR U8012 ( .A(p_input[2059]), .B(p_input[267]), .Z(n8142) );
  XOR U8013 ( .A(p_input[2060]), .B(p_input[268]), .Z(n8102) );
  XNOR U8014 ( .A(n8112), .B(n8103), .Z(n8141) );
  XNOR U8015 ( .A(n6553), .B(p_input[257]), .Z(n8103) );
  XOR U8016 ( .A(n8143), .B(n8118), .Z(n8112) );
  XNOR U8017 ( .A(p_input[2063]), .B(p_input[271]), .Z(n8118) );
  XOR U8018 ( .A(n8109), .B(n8117), .Z(n8143) );
  XOR U8019 ( .A(n8144), .B(n8114), .Z(n8117) );
  XOR U8020 ( .A(p_input[2061]), .B(p_input[269]), .Z(n8114) );
  XNOR U8021 ( .A(p_input[2062]), .B(p_input[270]), .Z(n8144) );
  XNOR U8022 ( .A(n6325), .B(p_input[265]), .Z(n8109) );
  XNOR U8023 ( .A(n8125), .B(n8124), .Z(n8107) );
  XNOR U8024 ( .A(n8145), .B(n8130), .Z(n8124) );
  XOR U8025 ( .A(p_input[2056]), .B(p_input[264]), .Z(n8130) );
  XOR U8026 ( .A(n8121), .B(n8129), .Z(n8145) );
  XOR U8027 ( .A(n8146), .B(n8126), .Z(n8129) );
  XOR U8028 ( .A(p_input[2054]), .B(p_input[262]), .Z(n8126) );
  XNOR U8029 ( .A(p_input[2055]), .B(p_input[263]), .Z(n8146) );
  XNOR U8030 ( .A(n6328), .B(p_input[258]), .Z(n8121) );
  XNOR U8031 ( .A(n8135), .B(n8134), .Z(n8125) );
  XOR U8032 ( .A(n8147), .B(n8131), .Z(n8134) );
  XOR U8033 ( .A(p_input[2051]), .B(p_input[259]), .Z(n8131) );
  XNOR U8034 ( .A(p_input[2052]), .B(p_input[260]), .Z(n8147) );
  XOR U8035 ( .A(p_input[2053]), .B(p_input[261]), .Z(n8135) );
  XOR U8036 ( .A(n8148), .B(n8149), .Z(n8036) );
  AND U8037 ( .A(n71), .B(n8150), .Z(n8149) );
  XNOR U8038 ( .A(n8151), .B(n8148), .Z(n8150) );
  XNOR U8039 ( .A(n8152), .B(n8153), .Z(n71) );
  AND U8040 ( .A(n8154), .B(n8155), .Z(n8153) );
  XOR U8041 ( .A(n8049), .B(n8152), .Z(n8155) );
  AND U8042 ( .A(n8156), .B(n8157), .Z(n8049) );
  XNOR U8043 ( .A(n8046), .B(n8152), .Z(n8154) );
  XOR U8044 ( .A(n8158), .B(n8159), .Z(n8046) );
  AND U8045 ( .A(n75), .B(n8160), .Z(n8159) );
  XOR U8046 ( .A(n8161), .B(n8158), .Z(n8160) );
  XOR U8047 ( .A(n8162), .B(n8163), .Z(n8152) );
  AND U8048 ( .A(n8164), .B(n8165), .Z(n8163) );
  XNOR U8049 ( .A(n8162), .B(n8156), .Z(n8165) );
  IV U8050 ( .A(n8064), .Z(n8156) );
  XOR U8051 ( .A(n8166), .B(n8167), .Z(n8064) );
  XOR U8052 ( .A(n8168), .B(n8157), .Z(n8167) );
  AND U8053 ( .A(n8091), .B(n8169), .Z(n8157) );
  AND U8054 ( .A(n8170), .B(n8171), .Z(n8168) );
  XOR U8055 ( .A(n8172), .B(n8166), .Z(n8170) );
  XNOR U8056 ( .A(n8061), .B(n8162), .Z(n8164) );
  XOR U8057 ( .A(n8173), .B(n8174), .Z(n8061) );
  AND U8058 ( .A(n75), .B(n8175), .Z(n8174) );
  XOR U8059 ( .A(n8176), .B(n8173), .Z(n8175) );
  XOR U8060 ( .A(n8177), .B(n8178), .Z(n8162) );
  AND U8061 ( .A(n8179), .B(n8180), .Z(n8178) );
  XNOR U8062 ( .A(n8177), .B(n8091), .Z(n8180) );
  XOR U8063 ( .A(n8181), .B(n8171), .Z(n8091) );
  XNOR U8064 ( .A(n8182), .B(n8166), .Z(n8171) );
  XOR U8065 ( .A(n8183), .B(n8184), .Z(n8166) );
  AND U8066 ( .A(n8185), .B(n8186), .Z(n8184) );
  XOR U8067 ( .A(n8187), .B(n8183), .Z(n8185) );
  XNOR U8068 ( .A(n8188), .B(n8189), .Z(n8182) );
  AND U8069 ( .A(n8190), .B(n8191), .Z(n8189) );
  XOR U8070 ( .A(n8188), .B(n8192), .Z(n8190) );
  XNOR U8071 ( .A(n8172), .B(n8169), .Z(n8181) );
  AND U8072 ( .A(n8193), .B(n8194), .Z(n8169) );
  XOR U8073 ( .A(n8195), .B(n8196), .Z(n8172) );
  AND U8074 ( .A(n8197), .B(n8198), .Z(n8196) );
  XOR U8075 ( .A(n8195), .B(n8199), .Z(n8197) );
  XNOR U8076 ( .A(n8088), .B(n8177), .Z(n8179) );
  XOR U8077 ( .A(n8200), .B(n8201), .Z(n8088) );
  AND U8078 ( .A(n75), .B(n8202), .Z(n8201) );
  XNOR U8079 ( .A(n8203), .B(n8200), .Z(n8202) );
  XOR U8080 ( .A(n8204), .B(n8205), .Z(n8177) );
  AND U8081 ( .A(n8206), .B(n8207), .Z(n8205) );
  XNOR U8082 ( .A(n8204), .B(n8193), .Z(n8207) );
  IV U8083 ( .A(n8139), .Z(n8193) );
  XNOR U8084 ( .A(n8208), .B(n8186), .Z(n8139) );
  XNOR U8085 ( .A(n8209), .B(n8192), .Z(n8186) );
  XOR U8086 ( .A(n8210), .B(n8211), .Z(n8192) );
  NOR U8087 ( .A(n8212), .B(n8213), .Z(n8211) );
  XNOR U8088 ( .A(n8210), .B(n8214), .Z(n8212) );
  XNOR U8089 ( .A(n8191), .B(n8183), .Z(n8209) );
  XOR U8090 ( .A(n8215), .B(n8216), .Z(n8183) );
  AND U8091 ( .A(n8217), .B(n8218), .Z(n8216) );
  XNOR U8092 ( .A(n8215), .B(n8219), .Z(n8217) );
  XNOR U8093 ( .A(n8220), .B(n8188), .Z(n8191) );
  XOR U8094 ( .A(n8221), .B(n8222), .Z(n8188) );
  AND U8095 ( .A(n8223), .B(n8224), .Z(n8222) );
  XOR U8096 ( .A(n8221), .B(n8225), .Z(n8223) );
  XNOR U8097 ( .A(n8226), .B(n8227), .Z(n8220) );
  NOR U8098 ( .A(n8228), .B(n8229), .Z(n8227) );
  XOR U8099 ( .A(n8226), .B(n8230), .Z(n8228) );
  XNOR U8100 ( .A(n8187), .B(n8194), .Z(n8208) );
  NOR U8101 ( .A(n8151), .B(n8231), .Z(n8194) );
  XOR U8102 ( .A(n8199), .B(n8198), .Z(n8187) );
  XNOR U8103 ( .A(n8232), .B(n8195), .Z(n8198) );
  XOR U8104 ( .A(n8233), .B(n8234), .Z(n8195) );
  AND U8105 ( .A(n8235), .B(n8236), .Z(n8234) );
  XOR U8106 ( .A(n8233), .B(n8237), .Z(n8235) );
  XNOR U8107 ( .A(n8238), .B(n8239), .Z(n8232) );
  NOR U8108 ( .A(n8240), .B(n8241), .Z(n8239) );
  XNOR U8109 ( .A(n8238), .B(n8242), .Z(n8240) );
  XOR U8110 ( .A(n8243), .B(n8244), .Z(n8199) );
  NOR U8111 ( .A(n8245), .B(n8246), .Z(n8244) );
  XNOR U8112 ( .A(n8243), .B(n8247), .Z(n8245) );
  XNOR U8113 ( .A(n8136), .B(n8204), .Z(n8206) );
  XOR U8114 ( .A(n8248), .B(n8249), .Z(n8136) );
  AND U8115 ( .A(n75), .B(n8250), .Z(n8249) );
  XOR U8116 ( .A(n8251), .B(n8248), .Z(n8250) );
  AND U8117 ( .A(n8148), .B(n8151), .Z(n8204) );
  XOR U8118 ( .A(n8252), .B(n8231), .Z(n8151) );
  XNOR U8119 ( .A(p_input[2048]), .B(p_input[272]), .Z(n8231) );
  XOR U8120 ( .A(n8219), .B(n8218), .Z(n8252) );
  XNOR U8121 ( .A(n8253), .B(n8225), .Z(n8218) );
  XNOR U8122 ( .A(n8214), .B(n8213), .Z(n8225) );
  XOR U8123 ( .A(n8254), .B(n8210), .Z(n8213) );
  XNOR U8124 ( .A(n6439), .B(p_input[282]), .Z(n8210) );
  XNOR U8125 ( .A(p_input[2059]), .B(p_input[283]), .Z(n8254) );
  XOR U8126 ( .A(p_input[2060]), .B(p_input[284]), .Z(n8214) );
  XNOR U8127 ( .A(n8224), .B(n8215), .Z(n8253) );
  XNOR U8128 ( .A(n6553), .B(p_input[273]), .Z(n8215) );
  XOR U8129 ( .A(n8255), .B(n8230), .Z(n8224) );
  XNOR U8130 ( .A(p_input[2063]), .B(p_input[287]), .Z(n8230) );
  XOR U8131 ( .A(n8221), .B(n8229), .Z(n8255) );
  XOR U8132 ( .A(n8256), .B(n8226), .Z(n8229) );
  XOR U8133 ( .A(p_input[2061]), .B(p_input[285]), .Z(n8226) );
  XNOR U8134 ( .A(p_input[2062]), .B(p_input[286]), .Z(n8256) );
  XNOR U8135 ( .A(n6325), .B(p_input[281]), .Z(n8221) );
  XNOR U8136 ( .A(n8237), .B(n8236), .Z(n8219) );
  XNOR U8137 ( .A(n8257), .B(n8242), .Z(n8236) );
  XOR U8138 ( .A(p_input[2056]), .B(p_input[280]), .Z(n8242) );
  XOR U8139 ( .A(n8233), .B(n8241), .Z(n8257) );
  XOR U8140 ( .A(n8258), .B(n8238), .Z(n8241) );
  XOR U8141 ( .A(p_input[2054]), .B(p_input[278]), .Z(n8238) );
  XNOR U8142 ( .A(p_input[2055]), .B(p_input[279]), .Z(n8258) );
  XNOR U8143 ( .A(n6328), .B(p_input[274]), .Z(n8233) );
  XNOR U8144 ( .A(n8247), .B(n8246), .Z(n8237) );
  XOR U8145 ( .A(n8259), .B(n8243), .Z(n8246) );
  XOR U8146 ( .A(p_input[2051]), .B(p_input[275]), .Z(n8243) );
  XNOR U8147 ( .A(p_input[2052]), .B(p_input[276]), .Z(n8259) );
  XOR U8148 ( .A(p_input[2053]), .B(p_input[277]), .Z(n8247) );
  XOR U8149 ( .A(n8260), .B(n8261), .Z(n8148) );
  AND U8150 ( .A(n75), .B(n8262), .Z(n8261) );
  XNOR U8151 ( .A(n8263), .B(n8260), .Z(n8262) );
  XNOR U8152 ( .A(n8264), .B(n8265), .Z(n75) );
  AND U8153 ( .A(n8266), .B(n8267), .Z(n8265) );
  XOR U8154 ( .A(n8161), .B(n8264), .Z(n8267) );
  AND U8155 ( .A(n8268), .B(n8269), .Z(n8161) );
  XNOR U8156 ( .A(n8158), .B(n8264), .Z(n8266) );
  XOR U8157 ( .A(n8270), .B(n8271), .Z(n8158) );
  AND U8158 ( .A(n79), .B(n8272), .Z(n8271) );
  XOR U8159 ( .A(n8273), .B(n8270), .Z(n8272) );
  XOR U8160 ( .A(n8274), .B(n8275), .Z(n8264) );
  AND U8161 ( .A(n8276), .B(n8277), .Z(n8275) );
  XNOR U8162 ( .A(n8274), .B(n8268), .Z(n8277) );
  IV U8163 ( .A(n8176), .Z(n8268) );
  XOR U8164 ( .A(n8278), .B(n8279), .Z(n8176) );
  XOR U8165 ( .A(n8280), .B(n8269), .Z(n8279) );
  AND U8166 ( .A(n8203), .B(n8281), .Z(n8269) );
  AND U8167 ( .A(n8282), .B(n8283), .Z(n8280) );
  XOR U8168 ( .A(n8284), .B(n8278), .Z(n8282) );
  XNOR U8169 ( .A(n8173), .B(n8274), .Z(n8276) );
  XOR U8170 ( .A(n8285), .B(n8286), .Z(n8173) );
  AND U8171 ( .A(n79), .B(n8287), .Z(n8286) );
  XOR U8172 ( .A(n8288), .B(n8285), .Z(n8287) );
  XOR U8173 ( .A(n8289), .B(n8290), .Z(n8274) );
  AND U8174 ( .A(n8291), .B(n8292), .Z(n8290) );
  XNOR U8175 ( .A(n8289), .B(n8203), .Z(n8292) );
  XOR U8176 ( .A(n8293), .B(n8283), .Z(n8203) );
  XNOR U8177 ( .A(n8294), .B(n8278), .Z(n8283) );
  XOR U8178 ( .A(n8295), .B(n8296), .Z(n8278) );
  AND U8179 ( .A(n8297), .B(n8298), .Z(n8296) );
  XOR U8180 ( .A(n8299), .B(n8295), .Z(n8297) );
  XNOR U8181 ( .A(n8300), .B(n8301), .Z(n8294) );
  AND U8182 ( .A(n8302), .B(n8303), .Z(n8301) );
  XOR U8183 ( .A(n8300), .B(n8304), .Z(n8302) );
  XNOR U8184 ( .A(n8284), .B(n8281), .Z(n8293) );
  AND U8185 ( .A(n8305), .B(n8306), .Z(n8281) );
  XOR U8186 ( .A(n8307), .B(n8308), .Z(n8284) );
  AND U8187 ( .A(n8309), .B(n8310), .Z(n8308) );
  XOR U8188 ( .A(n8307), .B(n8311), .Z(n8309) );
  XNOR U8189 ( .A(n8200), .B(n8289), .Z(n8291) );
  XOR U8190 ( .A(n8312), .B(n8313), .Z(n8200) );
  AND U8191 ( .A(n79), .B(n8314), .Z(n8313) );
  XNOR U8192 ( .A(n8315), .B(n8312), .Z(n8314) );
  XOR U8193 ( .A(n8316), .B(n8317), .Z(n8289) );
  AND U8194 ( .A(n8318), .B(n8319), .Z(n8317) );
  XNOR U8195 ( .A(n8316), .B(n8305), .Z(n8319) );
  IV U8196 ( .A(n8251), .Z(n8305) );
  XNOR U8197 ( .A(n8320), .B(n8298), .Z(n8251) );
  XNOR U8198 ( .A(n8321), .B(n8304), .Z(n8298) );
  XOR U8199 ( .A(n8322), .B(n8323), .Z(n8304) );
  NOR U8200 ( .A(n8324), .B(n8325), .Z(n8323) );
  XNOR U8201 ( .A(n8322), .B(n8326), .Z(n8324) );
  XNOR U8202 ( .A(n8303), .B(n8295), .Z(n8321) );
  XOR U8203 ( .A(n8327), .B(n8328), .Z(n8295) );
  AND U8204 ( .A(n8329), .B(n8330), .Z(n8328) );
  XNOR U8205 ( .A(n8327), .B(n8331), .Z(n8329) );
  XNOR U8206 ( .A(n8332), .B(n8300), .Z(n8303) );
  XOR U8207 ( .A(n8333), .B(n8334), .Z(n8300) );
  AND U8208 ( .A(n8335), .B(n8336), .Z(n8334) );
  XOR U8209 ( .A(n8333), .B(n8337), .Z(n8335) );
  XNOR U8210 ( .A(n8338), .B(n8339), .Z(n8332) );
  NOR U8211 ( .A(n8340), .B(n8341), .Z(n8339) );
  XOR U8212 ( .A(n8338), .B(n8342), .Z(n8340) );
  XNOR U8213 ( .A(n8299), .B(n8306), .Z(n8320) );
  NOR U8214 ( .A(n8263), .B(n8343), .Z(n8306) );
  XOR U8215 ( .A(n8311), .B(n8310), .Z(n8299) );
  XNOR U8216 ( .A(n8344), .B(n8307), .Z(n8310) );
  XOR U8217 ( .A(n8345), .B(n8346), .Z(n8307) );
  AND U8218 ( .A(n8347), .B(n8348), .Z(n8346) );
  XOR U8219 ( .A(n8345), .B(n8349), .Z(n8347) );
  XNOR U8220 ( .A(n8350), .B(n8351), .Z(n8344) );
  NOR U8221 ( .A(n8352), .B(n8353), .Z(n8351) );
  XNOR U8222 ( .A(n8350), .B(n8354), .Z(n8352) );
  XOR U8223 ( .A(n8355), .B(n8356), .Z(n8311) );
  NOR U8224 ( .A(n8357), .B(n8358), .Z(n8356) );
  XNOR U8225 ( .A(n8355), .B(n8359), .Z(n8357) );
  XNOR U8226 ( .A(n8248), .B(n8316), .Z(n8318) );
  XOR U8227 ( .A(n8360), .B(n8361), .Z(n8248) );
  AND U8228 ( .A(n79), .B(n8362), .Z(n8361) );
  XOR U8229 ( .A(n8363), .B(n8360), .Z(n8362) );
  AND U8230 ( .A(n8260), .B(n8263), .Z(n8316) );
  XOR U8231 ( .A(n8364), .B(n8343), .Z(n8263) );
  XNOR U8232 ( .A(p_input[2048]), .B(p_input[288]), .Z(n8343) );
  XOR U8233 ( .A(n8331), .B(n8330), .Z(n8364) );
  XNOR U8234 ( .A(n8365), .B(n8337), .Z(n8330) );
  XNOR U8235 ( .A(n8326), .B(n8325), .Z(n8337) );
  XOR U8236 ( .A(n8366), .B(n8322), .Z(n8325) );
  XNOR U8237 ( .A(n6439), .B(p_input[298]), .Z(n8322) );
  XNOR U8238 ( .A(p_input[2059]), .B(p_input[299]), .Z(n8366) );
  XOR U8239 ( .A(p_input[2060]), .B(p_input[300]), .Z(n8326) );
  XNOR U8240 ( .A(n8336), .B(n8327), .Z(n8365) );
  XNOR U8241 ( .A(n6553), .B(p_input[289]), .Z(n8327) );
  XOR U8242 ( .A(n8367), .B(n8342), .Z(n8336) );
  XNOR U8243 ( .A(p_input[2063]), .B(p_input[303]), .Z(n8342) );
  XOR U8244 ( .A(n8333), .B(n8341), .Z(n8367) );
  XOR U8245 ( .A(n8368), .B(n8338), .Z(n8341) );
  XOR U8246 ( .A(p_input[2061]), .B(p_input[301]), .Z(n8338) );
  XNOR U8247 ( .A(p_input[2062]), .B(p_input[302]), .Z(n8368) );
  XNOR U8248 ( .A(n6325), .B(p_input[297]), .Z(n8333) );
  XNOR U8249 ( .A(n8349), .B(n8348), .Z(n8331) );
  XNOR U8250 ( .A(n8369), .B(n8354), .Z(n8348) );
  XOR U8251 ( .A(p_input[2056]), .B(p_input[296]), .Z(n8354) );
  XOR U8252 ( .A(n8345), .B(n8353), .Z(n8369) );
  XOR U8253 ( .A(n8370), .B(n8350), .Z(n8353) );
  XOR U8254 ( .A(p_input[2054]), .B(p_input[294]), .Z(n8350) );
  XNOR U8255 ( .A(p_input[2055]), .B(p_input[295]), .Z(n8370) );
  XNOR U8256 ( .A(n6328), .B(p_input[290]), .Z(n8345) );
  XNOR U8257 ( .A(n8359), .B(n8358), .Z(n8349) );
  XOR U8258 ( .A(n8371), .B(n8355), .Z(n8358) );
  XOR U8259 ( .A(p_input[2051]), .B(p_input[291]), .Z(n8355) );
  XNOR U8260 ( .A(p_input[2052]), .B(p_input[292]), .Z(n8371) );
  XOR U8261 ( .A(p_input[2053]), .B(p_input[293]), .Z(n8359) );
  XOR U8262 ( .A(n8372), .B(n8373), .Z(n8260) );
  AND U8263 ( .A(n79), .B(n8374), .Z(n8373) );
  XNOR U8264 ( .A(n8375), .B(n8372), .Z(n8374) );
  XNOR U8265 ( .A(n8376), .B(n8377), .Z(n79) );
  AND U8266 ( .A(n8378), .B(n8379), .Z(n8377) );
  XOR U8267 ( .A(n8273), .B(n8376), .Z(n8379) );
  AND U8268 ( .A(n8380), .B(n8381), .Z(n8273) );
  XNOR U8269 ( .A(n8270), .B(n8376), .Z(n8378) );
  XOR U8270 ( .A(n8382), .B(n8383), .Z(n8270) );
  AND U8271 ( .A(n83), .B(n8384), .Z(n8383) );
  XOR U8272 ( .A(n8385), .B(n8382), .Z(n8384) );
  XOR U8273 ( .A(n8386), .B(n8387), .Z(n8376) );
  AND U8274 ( .A(n8388), .B(n8389), .Z(n8387) );
  XNOR U8275 ( .A(n8386), .B(n8380), .Z(n8389) );
  IV U8276 ( .A(n8288), .Z(n8380) );
  XOR U8277 ( .A(n8390), .B(n8391), .Z(n8288) );
  XOR U8278 ( .A(n8392), .B(n8381), .Z(n8391) );
  AND U8279 ( .A(n8315), .B(n8393), .Z(n8381) );
  AND U8280 ( .A(n8394), .B(n8395), .Z(n8392) );
  XOR U8281 ( .A(n8396), .B(n8390), .Z(n8394) );
  XNOR U8282 ( .A(n8285), .B(n8386), .Z(n8388) );
  XOR U8283 ( .A(n8397), .B(n8398), .Z(n8285) );
  AND U8284 ( .A(n83), .B(n8399), .Z(n8398) );
  XOR U8285 ( .A(n8400), .B(n8397), .Z(n8399) );
  XOR U8286 ( .A(n8401), .B(n8402), .Z(n8386) );
  AND U8287 ( .A(n8403), .B(n8404), .Z(n8402) );
  XNOR U8288 ( .A(n8401), .B(n8315), .Z(n8404) );
  XOR U8289 ( .A(n8405), .B(n8395), .Z(n8315) );
  XNOR U8290 ( .A(n8406), .B(n8390), .Z(n8395) );
  XOR U8291 ( .A(n8407), .B(n8408), .Z(n8390) );
  AND U8292 ( .A(n8409), .B(n8410), .Z(n8408) );
  XOR U8293 ( .A(n8411), .B(n8407), .Z(n8409) );
  XNOR U8294 ( .A(n8412), .B(n8413), .Z(n8406) );
  AND U8295 ( .A(n8414), .B(n8415), .Z(n8413) );
  XOR U8296 ( .A(n8412), .B(n8416), .Z(n8414) );
  XNOR U8297 ( .A(n8396), .B(n8393), .Z(n8405) );
  AND U8298 ( .A(n8417), .B(n8418), .Z(n8393) );
  XOR U8299 ( .A(n8419), .B(n8420), .Z(n8396) );
  AND U8300 ( .A(n8421), .B(n8422), .Z(n8420) );
  XOR U8301 ( .A(n8419), .B(n8423), .Z(n8421) );
  XNOR U8302 ( .A(n8312), .B(n8401), .Z(n8403) );
  XOR U8303 ( .A(n8424), .B(n8425), .Z(n8312) );
  AND U8304 ( .A(n83), .B(n8426), .Z(n8425) );
  XNOR U8305 ( .A(n8427), .B(n8424), .Z(n8426) );
  XOR U8306 ( .A(n8428), .B(n8429), .Z(n8401) );
  AND U8307 ( .A(n8430), .B(n8431), .Z(n8429) );
  XNOR U8308 ( .A(n8428), .B(n8417), .Z(n8431) );
  IV U8309 ( .A(n8363), .Z(n8417) );
  XNOR U8310 ( .A(n8432), .B(n8410), .Z(n8363) );
  XNOR U8311 ( .A(n8433), .B(n8416), .Z(n8410) );
  XOR U8312 ( .A(n8434), .B(n8435), .Z(n8416) );
  NOR U8313 ( .A(n8436), .B(n8437), .Z(n8435) );
  XNOR U8314 ( .A(n8434), .B(n8438), .Z(n8436) );
  XNOR U8315 ( .A(n8415), .B(n8407), .Z(n8433) );
  XOR U8316 ( .A(n8439), .B(n8440), .Z(n8407) );
  AND U8317 ( .A(n8441), .B(n8442), .Z(n8440) );
  XNOR U8318 ( .A(n8439), .B(n8443), .Z(n8441) );
  XNOR U8319 ( .A(n8444), .B(n8412), .Z(n8415) );
  XOR U8320 ( .A(n8445), .B(n8446), .Z(n8412) );
  AND U8321 ( .A(n8447), .B(n8448), .Z(n8446) );
  XOR U8322 ( .A(n8445), .B(n8449), .Z(n8447) );
  XNOR U8323 ( .A(n8450), .B(n8451), .Z(n8444) );
  NOR U8324 ( .A(n8452), .B(n8453), .Z(n8451) );
  XOR U8325 ( .A(n8450), .B(n8454), .Z(n8452) );
  XNOR U8326 ( .A(n8411), .B(n8418), .Z(n8432) );
  NOR U8327 ( .A(n8375), .B(n8455), .Z(n8418) );
  XOR U8328 ( .A(n8423), .B(n8422), .Z(n8411) );
  XNOR U8329 ( .A(n8456), .B(n8419), .Z(n8422) );
  XOR U8330 ( .A(n8457), .B(n8458), .Z(n8419) );
  AND U8331 ( .A(n8459), .B(n8460), .Z(n8458) );
  XOR U8332 ( .A(n8457), .B(n8461), .Z(n8459) );
  XNOR U8333 ( .A(n8462), .B(n8463), .Z(n8456) );
  NOR U8334 ( .A(n8464), .B(n8465), .Z(n8463) );
  XNOR U8335 ( .A(n8462), .B(n8466), .Z(n8464) );
  XOR U8336 ( .A(n8467), .B(n8468), .Z(n8423) );
  NOR U8337 ( .A(n8469), .B(n8470), .Z(n8468) );
  XNOR U8338 ( .A(n8467), .B(n8471), .Z(n8469) );
  XNOR U8339 ( .A(n8360), .B(n8428), .Z(n8430) );
  XOR U8340 ( .A(n8472), .B(n8473), .Z(n8360) );
  AND U8341 ( .A(n83), .B(n8474), .Z(n8473) );
  XOR U8342 ( .A(n8475), .B(n8472), .Z(n8474) );
  AND U8343 ( .A(n8372), .B(n8375), .Z(n8428) );
  XOR U8344 ( .A(n8476), .B(n8455), .Z(n8375) );
  XNOR U8345 ( .A(p_input[2048]), .B(p_input[304]), .Z(n8455) );
  XOR U8346 ( .A(n8443), .B(n8442), .Z(n8476) );
  XNOR U8347 ( .A(n8477), .B(n8449), .Z(n8442) );
  XNOR U8348 ( .A(n8438), .B(n8437), .Z(n8449) );
  XOR U8349 ( .A(n8478), .B(n8434), .Z(n8437) );
  XNOR U8350 ( .A(n6439), .B(p_input[314]), .Z(n8434) );
  XNOR U8351 ( .A(p_input[2059]), .B(p_input[315]), .Z(n8478) );
  XOR U8352 ( .A(p_input[2060]), .B(p_input[316]), .Z(n8438) );
  XNOR U8353 ( .A(n8448), .B(n8439), .Z(n8477) );
  XNOR U8354 ( .A(n6553), .B(p_input[305]), .Z(n8439) );
  XOR U8355 ( .A(n8479), .B(n8454), .Z(n8448) );
  XNOR U8356 ( .A(p_input[2063]), .B(p_input[319]), .Z(n8454) );
  XOR U8357 ( .A(n8445), .B(n8453), .Z(n8479) );
  XOR U8358 ( .A(n8480), .B(n8450), .Z(n8453) );
  XOR U8359 ( .A(p_input[2061]), .B(p_input[317]), .Z(n8450) );
  XNOR U8360 ( .A(p_input[2062]), .B(p_input[318]), .Z(n8480) );
  XNOR U8361 ( .A(n6325), .B(p_input[313]), .Z(n8445) );
  XNOR U8362 ( .A(n8461), .B(n8460), .Z(n8443) );
  XNOR U8363 ( .A(n8481), .B(n8466), .Z(n8460) );
  XOR U8364 ( .A(p_input[2056]), .B(p_input[312]), .Z(n8466) );
  XOR U8365 ( .A(n8457), .B(n8465), .Z(n8481) );
  XOR U8366 ( .A(n8482), .B(n8462), .Z(n8465) );
  XOR U8367 ( .A(p_input[2054]), .B(p_input[310]), .Z(n8462) );
  XNOR U8368 ( .A(p_input[2055]), .B(p_input[311]), .Z(n8482) );
  XNOR U8369 ( .A(n6328), .B(p_input[306]), .Z(n8457) );
  XNOR U8370 ( .A(n8471), .B(n8470), .Z(n8461) );
  XOR U8371 ( .A(n8483), .B(n8467), .Z(n8470) );
  XOR U8372 ( .A(p_input[2051]), .B(p_input[307]), .Z(n8467) );
  XNOR U8373 ( .A(p_input[2052]), .B(p_input[308]), .Z(n8483) );
  XOR U8374 ( .A(p_input[2053]), .B(p_input[309]), .Z(n8471) );
  XOR U8375 ( .A(n8484), .B(n8485), .Z(n8372) );
  AND U8376 ( .A(n83), .B(n8486), .Z(n8485) );
  XNOR U8377 ( .A(n8487), .B(n8484), .Z(n8486) );
  XNOR U8378 ( .A(n8488), .B(n8489), .Z(n83) );
  AND U8379 ( .A(n8490), .B(n8491), .Z(n8489) );
  XOR U8380 ( .A(n8385), .B(n8488), .Z(n8491) );
  AND U8381 ( .A(n8492), .B(n8493), .Z(n8385) );
  XNOR U8382 ( .A(n8382), .B(n8488), .Z(n8490) );
  XOR U8383 ( .A(n8494), .B(n8495), .Z(n8382) );
  AND U8384 ( .A(n87), .B(n8496), .Z(n8495) );
  XOR U8385 ( .A(n8497), .B(n8494), .Z(n8496) );
  XOR U8386 ( .A(n8498), .B(n8499), .Z(n8488) );
  AND U8387 ( .A(n8500), .B(n8501), .Z(n8499) );
  XNOR U8388 ( .A(n8498), .B(n8492), .Z(n8501) );
  IV U8389 ( .A(n8400), .Z(n8492) );
  XOR U8390 ( .A(n8502), .B(n8503), .Z(n8400) );
  XOR U8391 ( .A(n8504), .B(n8493), .Z(n8503) );
  AND U8392 ( .A(n8427), .B(n8505), .Z(n8493) );
  AND U8393 ( .A(n8506), .B(n8507), .Z(n8504) );
  XOR U8394 ( .A(n8508), .B(n8502), .Z(n8506) );
  XNOR U8395 ( .A(n8397), .B(n8498), .Z(n8500) );
  XOR U8396 ( .A(n8509), .B(n8510), .Z(n8397) );
  AND U8397 ( .A(n87), .B(n8511), .Z(n8510) );
  XOR U8398 ( .A(n8512), .B(n8509), .Z(n8511) );
  XOR U8399 ( .A(n8513), .B(n8514), .Z(n8498) );
  AND U8400 ( .A(n8515), .B(n8516), .Z(n8514) );
  XNOR U8401 ( .A(n8513), .B(n8427), .Z(n8516) );
  XOR U8402 ( .A(n8517), .B(n8507), .Z(n8427) );
  XNOR U8403 ( .A(n8518), .B(n8502), .Z(n8507) );
  XOR U8404 ( .A(n8519), .B(n8520), .Z(n8502) );
  AND U8405 ( .A(n8521), .B(n8522), .Z(n8520) );
  XOR U8406 ( .A(n8523), .B(n8519), .Z(n8521) );
  XNOR U8407 ( .A(n8524), .B(n8525), .Z(n8518) );
  AND U8408 ( .A(n8526), .B(n8527), .Z(n8525) );
  XOR U8409 ( .A(n8524), .B(n8528), .Z(n8526) );
  XNOR U8410 ( .A(n8508), .B(n8505), .Z(n8517) );
  AND U8411 ( .A(n8529), .B(n8530), .Z(n8505) );
  XOR U8412 ( .A(n8531), .B(n8532), .Z(n8508) );
  AND U8413 ( .A(n8533), .B(n8534), .Z(n8532) );
  XOR U8414 ( .A(n8531), .B(n8535), .Z(n8533) );
  XNOR U8415 ( .A(n8424), .B(n8513), .Z(n8515) );
  XOR U8416 ( .A(n8536), .B(n8537), .Z(n8424) );
  AND U8417 ( .A(n87), .B(n8538), .Z(n8537) );
  XNOR U8418 ( .A(n8539), .B(n8536), .Z(n8538) );
  XOR U8419 ( .A(n8540), .B(n8541), .Z(n8513) );
  AND U8420 ( .A(n8542), .B(n8543), .Z(n8541) );
  XNOR U8421 ( .A(n8540), .B(n8529), .Z(n8543) );
  IV U8422 ( .A(n8475), .Z(n8529) );
  XNOR U8423 ( .A(n8544), .B(n8522), .Z(n8475) );
  XNOR U8424 ( .A(n8545), .B(n8528), .Z(n8522) );
  XOR U8425 ( .A(n8546), .B(n8547), .Z(n8528) );
  NOR U8426 ( .A(n8548), .B(n8549), .Z(n8547) );
  XNOR U8427 ( .A(n8546), .B(n8550), .Z(n8548) );
  XNOR U8428 ( .A(n8527), .B(n8519), .Z(n8545) );
  XOR U8429 ( .A(n8551), .B(n8552), .Z(n8519) );
  AND U8430 ( .A(n8553), .B(n8554), .Z(n8552) );
  XNOR U8431 ( .A(n8551), .B(n8555), .Z(n8553) );
  XNOR U8432 ( .A(n8556), .B(n8524), .Z(n8527) );
  XOR U8433 ( .A(n8557), .B(n8558), .Z(n8524) );
  AND U8434 ( .A(n8559), .B(n8560), .Z(n8558) );
  XOR U8435 ( .A(n8557), .B(n8561), .Z(n8559) );
  XNOR U8436 ( .A(n8562), .B(n8563), .Z(n8556) );
  NOR U8437 ( .A(n8564), .B(n8565), .Z(n8563) );
  XOR U8438 ( .A(n8562), .B(n8566), .Z(n8564) );
  XNOR U8439 ( .A(n8523), .B(n8530), .Z(n8544) );
  NOR U8440 ( .A(n8487), .B(n8567), .Z(n8530) );
  XOR U8441 ( .A(n8535), .B(n8534), .Z(n8523) );
  XNOR U8442 ( .A(n8568), .B(n8531), .Z(n8534) );
  XOR U8443 ( .A(n8569), .B(n8570), .Z(n8531) );
  AND U8444 ( .A(n8571), .B(n8572), .Z(n8570) );
  XOR U8445 ( .A(n8569), .B(n8573), .Z(n8571) );
  XNOR U8446 ( .A(n8574), .B(n8575), .Z(n8568) );
  NOR U8447 ( .A(n8576), .B(n8577), .Z(n8575) );
  XNOR U8448 ( .A(n8574), .B(n8578), .Z(n8576) );
  XOR U8449 ( .A(n8579), .B(n8580), .Z(n8535) );
  NOR U8450 ( .A(n8581), .B(n8582), .Z(n8580) );
  XNOR U8451 ( .A(n8579), .B(n8583), .Z(n8581) );
  XNOR U8452 ( .A(n8472), .B(n8540), .Z(n8542) );
  XOR U8453 ( .A(n8584), .B(n8585), .Z(n8472) );
  AND U8454 ( .A(n87), .B(n8586), .Z(n8585) );
  XOR U8455 ( .A(n8587), .B(n8584), .Z(n8586) );
  AND U8456 ( .A(n8484), .B(n8487), .Z(n8540) );
  XOR U8457 ( .A(n8588), .B(n8567), .Z(n8487) );
  XNOR U8458 ( .A(p_input[2048]), .B(p_input[320]), .Z(n8567) );
  XOR U8459 ( .A(n8555), .B(n8554), .Z(n8588) );
  XNOR U8460 ( .A(n8589), .B(n8561), .Z(n8554) );
  XNOR U8461 ( .A(n8550), .B(n8549), .Z(n8561) );
  XOR U8462 ( .A(n8590), .B(n8546), .Z(n8549) );
  XNOR U8463 ( .A(n6439), .B(p_input[330]), .Z(n8546) );
  XNOR U8464 ( .A(p_input[2059]), .B(p_input[331]), .Z(n8590) );
  XOR U8465 ( .A(p_input[2060]), .B(p_input[332]), .Z(n8550) );
  XNOR U8466 ( .A(n8560), .B(n8551), .Z(n8589) );
  XNOR U8467 ( .A(n6553), .B(p_input[321]), .Z(n8551) );
  XOR U8468 ( .A(n8591), .B(n8566), .Z(n8560) );
  XNOR U8469 ( .A(p_input[2063]), .B(p_input[335]), .Z(n8566) );
  XOR U8470 ( .A(n8557), .B(n8565), .Z(n8591) );
  XOR U8471 ( .A(n8592), .B(n8562), .Z(n8565) );
  XOR U8472 ( .A(p_input[2061]), .B(p_input[333]), .Z(n8562) );
  XNOR U8473 ( .A(p_input[2062]), .B(p_input[334]), .Z(n8592) );
  XNOR U8474 ( .A(n6325), .B(p_input[329]), .Z(n8557) );
  XNOR U8475 ( .A(n8573), .B(n8572), .Z(n8555) );
  XNOR U8476 ( .A(n8593), .B(n8578), .Z(n8572) );
  XOR U8477 ( .A(p_input[2056]), .B(p_input[328]), .Z(n8578) );
  XOR U8478 ( .A(n8569), .B(n8577), .Z(n8593) );
  XOR U8479 ( .A(n8594), .B(n8574), .Z(n8577) );
  XOR U8480 ( .A(p_input[2054]), .B(p_input[326]), .Z(n8574) );
  XNOR U8481 ( .A(p_input[2055]), .B(p_input[327]), .Z(n8594) );
  XNOR U8482 ( .A(n6328), .B(p_input[322]), .Z(n8569) );
  XNOR U8483 ( .A(n8583), .B(n8582), .Z(n8573) );
  XOR U8484 ( .A(n8595), .B(n8579), .Z(n8582) );
  XOR U8485 ( .A(p_input[2051]), .B(p_input[323]), .Z(n8579) );
  XNOR U8486 ( .A(p_input[2052]), .B(p_input[324]), .Z(n8595) );
  XOR U8487 ( .A(p_input[2053]), .B(p_input[325]), .Z(n8583) );
  XOR U8488 ( .A(n8596), .B(n8597), .Z(n8484) );
  AND U8489 ( .A(n87), .B(n8598), .Z(n8597) );
  XNOR U8490 ( .A(n8599), .B(n8596), .Z(n8598) );
  XNOR U8491 ( .A(n8600), .B(n8601), .Z(n87) );
  AND U8492 ( .A(n8602), .B(n8603), .Z(n8601) );
  XOR U8493 ( .A(n8497), .B(n8600), .Z(n8603) );
  AND U8494 ( .A(n8604), .B(n8605), .Z(n8497) );
  XNOR U8495 ( .A(n8494), .B(n8600), .Z(n8602) );
  XOR U8496 ( .A(n8606), .B(n8607), .Z(n8494) );
  AND U8497 ( .A(n91), .B(n8608), .Z(n8607) );
  XOR U8498 ( .A(n8609), .B(n8606), .Z(n8608) );
  XOR U8499 ( .A(n8610), .B(n8611), .Z(n8600) );
  AND U8500 ( .A(n8612), .B(n8613), .Z(n8611) );
  XNOR U8501 ( .A(n8610), .B(n8604), .Z(n8613) );
  IV U8502 ( .A(n8512), .Z(n8604) );
  XOR U8503 ( .A(n8614), .B(n8615), .Z(n8512) );
  XOR U8504 ( .A(n8616), .B(n8605), .Z(n8615) );
  AND U8505 ( .A(n8539), .B(n8617), .Z(n8605) );
  AND U8506 ( .A(n8618), .B(n8619), .Z(n8616) );
  XOR U8507 ( .A(n8620), .B(n8614), .Z(n8618) );
  XNOR U8508 ( .A(n8509), .B(n8610), .Z(n8612) );
  XOR U8509 ( .A(n8621), .B(n8622), .Z(n8509) );
  AND U8510 ( .A(n91), .B(n8623), .Z(n8622) );
  XOR U8511 ( .A(n8624), .B(n8621), .Z(n8623) );
  XOR U8512 ( .A(n8625), .B(n8626), .Z(n8610) );
  AND U8513 ( .A(n8627), .B(n8628), .Z(n8626) );
  XNOR U8514 ( .A(n8625), .B(n8539), .Z(n8628) );
  XOR U8515 ( .A(n8629), .B(n8619), .Z(n8539) );
  XNOR U8516 ( .A(n8630), .B(n8614), .Z(n8619) );
  XOR U8517 ( .A(n8631), .B(n8632), .Z(n8614) );
  AND U8518 ( .A(n8633), .B(n8634), .Z(n8632) );
  XOR U8519 ( .A(n8635), .B(n8631), .Z(n8633) );
  XNOR U8520 ( .A(n8636), .B(n8637), .Z(n8630) );
  AND U8521 ( .A(n8638), .B(n8639), .Z(n8637) );
  XOR U8522 ( .A(n8636), .B(n8640), .Z(n8638) );
  XNOR U8523 ( .A(n8620), .B(n8617), .Z(n8629) );
  AND U8524 ( .A(n8641), .B(n8642), .Z(n8617) );
  XOR U8525 ( .A(n8643), .B(n8644), .Z(n8620) );
  AND U8526 ( .A(n8645), .B(n8646), .Z(n8644) );
  XOR U8527 ( .A(n8643), .B(n8647), .Z(n8645) );
  XNOR U8528 ( .A(n8536), .B(n8625), .Z(n8627) );
  XOR U8529 ( .A(n8648), .B(n8649), .Z(n8536) );
  AND U8530 ( .A(n91), .B(n8650), .Z(n8649) );
  XNOR U8531 ( .A(n8651), .B(n8648), .Z(n8650) );
  XOR U8532 ( .A(n8652), .B(n8653), .Z(n8625) );
  AND U8533 ( .A(n8654), .B(n8655), .Z(n8653) );
  XNOR U8534 ( .A(n8652), .B(n8641), .Z(n8655) );
  IV U8535 ( .A(n8587), .Z(n8641) );
  XNOR U8536 ( .A(n8656), .B(n8634), .Z(n8587) );
  XNOR U8537 ( .A(n8657), .B(n8640), .Z(n8634) );
  XOR U8538 ( .A(n8658), .B(n8659), .Z(n8640) );
  NOR U8539 ( .A(n8660), .B(n8661), .Z(n8659) );
  XNOR U8540 ( .A(n8658), .B(n8662), .Z(n8660) );
  XNOR U8541 ( .A(n8639), .B(n8631), .Z(n8657) );
  XOR U8542 ( .A(n8663), .B(n8664), .Z(n8631) );
  AND U8543 ( .A(n8665), .B(n8666), .Z(n8664) );
  XNOR U8544 ( .A(n8663), .B(n8667), .Z(n8665) );
  XNOR U8545 ( .A(n8668), .B(n8636), .Z(n8639) );
  XOR U8546 ( .A(n8669), .B(n8670), .Z(n8636) );
  AND U8547 ( .A(n8671), .B(n8672), .Z(n8670) );
  XOR U8548 ( .A(n8669), .B(n8673), .Z(n8671) );
  XNOR U8549 ( .A(n8674), .B(n8675), .Z(n8668) );
  NOR U8550 ( .A(n8676), .B(n8677), .Z(n8675) );
  XOR U8551 ( .A(n8674), .B(n8678), .Z(n8676) );
  XNOR U8552 ( .A(n8635), .B(n8642), .Z(n8656) );
  NOR U8553 ( .A(n8599), .B(n8679), .Z(n8642) );
  XOR U8554 ( .A(n8647), .B(n8646), .Z(n8635) );
  XNOR U8555 ( .A(n8680), .B(n8643), .Z(n8646) );
  XOR U8556 ( .A(n8681), .B(n8682), .Z(n8643) );
  AND U8557 ( .A(n8683), .B(n8684), .Z(n8682) );
  XOR U8558 ( .A(n8681), .B(n8685), .Z(n8683) );
  XNOR U8559 ( .A(n8686), .B(n8687), .Z(n8680) );
  NOR U8560 ( .A(n8688), .B(n8689), .Z(n8687) );
  XNOR U8561 ( .A(n8686), .B(n8690), .Z(n8688) );
  XOR U8562 ( .A(n8691), .B(n8692), .Z(n8647) );
  NOR U8563 ( .A(n8693), .B(n8694), .Z(n8692) );
  XNOR U8564 ( .A(n8691), .B(n8695), .Z(n8693) );
  XNOR U8565 ( .A(n8584), .B(n8652), .Z(n8654) );
  XOR U8566 ( .A(n8696), .B(n8697), .Z(n8584) );
  AND U8567 ( .A(n91), .B(n8698), .Z(n8697) );
  XOR U8568 ( .A(n8699), .B(n8696), .Z(n8698) );
  AND U8569 ( .A(n8596), .B(n8599), .Z(n8652) );
  XOR U8570 ( .A(n8700), .B(n8679), .Z(n8599) );
  XNOR U8571 ( .A(p_input[2048]), .B(p_input[336]), .Z(n8679) );
  XOR U8572 ( .A(n8667), .B(n8666), .Z(n8700) );
  XNOR U8573 ( .A(n8701), .B(n8673), .Z(n8666) );
  XNOR U8574 ( .A(n8662), .B(n8661), .Z(n8673) );
  XOR U8575 ( .A(n8702), .B(n8658), .Z(n8661) );
  XNOR U8576 ( .A(n6439), .B(p_input[346]), .Z(n8658) );
  XNOR U8577 ( .A(p_input[2059]), .B(p_input[347]), .Z(n8702) );
  XOR U8578 ( .A(p_input[2060]), .B(p_input[348]), .Z(n8662) );
  XNOR U8579 ( .A(n8672), .B(n8663), .Z(n8701) );
  XNOR U8580 ( .A(n6553), .B(p_input[337]), .Z(n8663) );
  XOR U8581 ( .A(n8703), .B(n8678), .Z(n8672) );
  XNOR U8582 ( .A(p_input[2063]), .B(p_input[351]), .Z(n8678) );
  XOR U8583 ( .A(n8669), .B(n8677), .Z(n8703) );
  XOR U8584 ( .A(n8704), .B(n8674), .Z(n8677) );
  XOR U8585 ( .A(p_input[2061]), .B(p_input[349]), .Z(n8674) );
  XNOR U8586 ( .A(p_input[2062]), .B(p_input[350]), .Z(n8704) );
  XNOR U8587 ( .A(n6325), .B(p_input[345]), .Z(n8669) );
  XNOR U8588 ( .A(n8685), .B(n8684), .Z(n8667) );
  XNOR U8589 ( .A(n8705), .B(n8690), .Z(n8684) );
  XOR U8590 ( .A(p_input[2056]), .B(p_input[344]), .Z(n8690) );
  XOR U8591 ( .A(n8681), .B(n8689), .Z(n8705) );
  XOR U8592 ( .A(n8706), .B(n8686), .Z(n8689) );
  XOR U8593 ( .A(p_input[2054]), .B(p_input[342]), .Z(n8686) );
  XNOR U8594 ( .A(p_input[2055]), .B(p_input[343]), .Z(n8706) );
  XNOR U8595 ( .A(n6328), .B(p_input[338]), .Z(n8681) );
  XNOR U8596 ( .A(n8695), .B(n8694), .Z(n8685) );
  XOR U8597 ( .A(n8707), .B(n8691), .Z(n8694) );
  XOR U8598 ( .A(p_input[2051]), .B(p_input[339]), .Z(n8691) );
  XNOR U8599 ( .A(p_input[2052]), .B(p_input[340]), .Z(n8707) );
  XOR U8600 ( .A(p_input[2053]), .B(p_input[341]), .Z(n8695) );
  XOR U8601 ( .A(n8708), .B(n8709), .Z(n8596) );
  AND U8602 ( .A(n91), .B(n8710), .Z(n8709) );
  XNOR U8603 ( .A(n8711), .B(n8708), .Z(n8710) );
  XNOR U8604 ( .A(n8712), .B(n8713), .Z(n91) );
  AND U8605 ( .A(n8714), .B(n8715), .Z(n8713) );
  XOR U8606 ( .A(n8609), .B(n8712), .Z(n8715) );
  AND U8607 ( .A(n8716), .B(n8717), .Z(n8609) );
  XNOR U8608 ( .A(n8606), .B(n8712), .Z(n8714) );
  XOR U8609 ( .A(n8718), .B(n8719), .Z(n8606) );
  AND U8610 ( .A(n95), .B(n8720), .Z(n8719) );
  XOR U8611 ( .A(n8721), .B(n8718), .Z(n8720) );
  XOR U8612 ( .A(n8722), .B(n8723), .Z(n8712) );
  AND U8613 ( .A(n8724), .B(n8725), .Z(n8723) );
  XNOR U8614 ( .A(n8722), .B(n8716), .Z(n8725) );
  IV U8615 ( .A(n8624), .Z(n8716) );
  XOR U8616 ( .A(n8726), .B(n8727), .Z(n8624) );
  XOR U8617 ( .A(n8728), .B(n8717), .Z(n8727) );
  AND U8618 ( .A(n8651), .B(n8729), .Z(n8717) );
  AND U8619 ( .A(n8730), .B(n8731), .Z(n8728) );
  XOR U8620 ( .A(n8732), .B(n8726), .Z(n8730) );
  XNOR U8621 ( .A(n8621), .B(n8722), .Z(n8724) );
  XOR U8622 ( .A(n8733), .B(n8734), .Z(n8621) );
  AND U8623 ( .A(n95), .B(n8735), .Z(n8734) );
  XOR U8624 ( .A(n8736), .B(n8733), .Z(n8735) );
  XOR U8625 ( .A(n8737), .B(n8738), .Z(n8722) );
  AND U8626 ( .A(n8739), .B(n8740), .Z(n8738) );
  XNOR U8627 ( .A(n8737), .B(n8651), .Z(n8740) );
  XOR U8628 ( .A(n8741), .B(n8731), .Z(n8651) );
  XNOR U8629 ( .A(n8742), .B(n8726), .Z(n8731) );
  XOR U8630 ( .A(n8743), .B(n8744), .Z(n8726) );
  AND U8631 ( .A(n8745), .B(n8746), .Z(n8744) );
  XOR U8632 ( .A(n8747), .B(n8743), .Z(n8745) );
  XNOR U8633 ( .A(n8748), .B(n8749), .Z(n8742) );
  AND U8634 ( .A(n8750), .B(n8751), .Z(n8749) );
  XOR U8635 ( .A(n8748), .B(n8752), .Z(n8750) );
  XNOR U8636 ( .A(n8732), .B(n8729), .Z(n8741) );
  AND U8637 ( .A(n8753), .B(n8754), .Z(n8729) );
  XOR U8638 ( .A(n8755), .B(n8756), .Z(n8732) );
  AND U8639 ( .A(n8757), .B(n8758), .Z(n8756) );
  XOR U8640 ( .A(n8755), .B(n8759), .Z(n8757) );
  XNOR U8641 ( .A(n8648), .B(n8737), .Z(n8739) );
  XOR U8642 ( .A(n8760), .B(n8761), .Z(n8648) );
  AND U8643 ( .A(n95), .B(n8762), .Z(n8761) );
  XNOR U8644 ( .A(n8763), .B(n8760), .Z(n8762) );
  XOR U8645 ( .A(n8764), .B(n8765), .Z(n8737) );
  AND U8646 ( .A(n8766), .B(n8767), .Z(n8765) );
  XNOR U8647 ( .A(n8764), .B(n8753), .Z(n8767) );
  IV U8648 ( .A(n8699), .Z(n8753) );
  XNOR U8649 ( .A(n8768), .B(n8746), .Z(n8699) );
  XNOR U8650 ( .A(n8769), .B(n8752), .Z(n8746) );
  XOR U8651 ( .A(n8770), .B(n8771), .Z(n8752) );
  NOR U8652 ( .A(n8772), .B(n8773), .Z(n8771) );
  XNOR U8653 ( .A(n8770), .B(n8774), .Z(n8772) );
  XNOR U8654 ( .A(n8751), .B(n8743), .Z(n8769) );
  XOR U8655 ( .A(n8775), .B(n8776), .Z(n8743) );
  AND U8656 ( .A(n8777), .B(n8778), .Z(n8776) );
  XNOR U8657 ( .A(n8775), .B(n8779), .Z(n8777) );
  XNOR U8658 ( .A(n8780), .B(n8748), .Z(n8751) );
  XOR U8659 ( .A(n8781), .B(n8782), .Z(n8748) );
  AND U8660 ( .A(n8783), .B(n8784), .Z(n8782) );
  XOR U8661 ( .A(n8781), .B(n8785), .Z(n8783) );
  XNOR U8662 ( .A(n8786), .B(n8787), .Z(n8780) );
  NOR U8663 ( .A(n8788), .B(n8789), .Z(n8787) );
  XOR U8664 ( .A(n8786), .B(n8790), .Z(n8788) );
  XNOR U8665 ( .A(n8747), .B(n8754), .Z(n8768) );
  NOR U8666 ( .A(n8711), .B(n8791), .Z(n8754) );
  XOR U8667 ( .A(n8759), .B(n8758), .Z(n8747) );
  XNOR U8668 ( .A(n8792), .B(n8755), .Z(n8758) );
  XOR U8669 ( .A(n8793), .B(n8794), .Z(n8755) );
  AND U8670 ( .A(n8795), .B(n8796), .Z(n8794) );
  XOR U8671 ( .A(n8793), .B(n8797), .Z(n8795) );
  XNOR U8672 ( .A(n8798), .B(n8799), .Z(n8792) );
  NOR U8673 ( .A(n8800), .B(n8801), .Z(n8799) );
  XNOR U8674 ( .A(n8798), .B(n8802), .Z(n8800) );
  XOR U8675 ( .A(n8803), .B(n8804), .Z(n8759) );
  NOR U8676 ( .A(n8805), .B(n8806), .Z(n8804) );
  XNOR U8677 ( .A(n8803), .B(n8807), .Z(n8805) );
  XNOR U8678 ( .A(n8696), .B(n8764), .Z(n8766) );
  XOR U8679 ( .A(n8808), .B(n8809), .Z(n8696) );
  AND U8680 ( .A(n95), .B(n8810), .Z(n8809) );
  XOR U8681 ( .A(n8811), .B(n8808), .Z(n8810) );
  AND U8682 ( .A(n8708), .B(n8711), .Z(n8764) );
  XOR U8683 ( .A(n8812), .B(n8791), .Z(n8711) );
  XNOR U8684 ( .A(p_input[2048]), .B(p_input[352]), .Z(n8791) );
  XOR U8685 ( .A(n8779), .B(n8778), .Z(n8812) );
  XNOR U8686 ( .A(n8813), .B(n8785), .Z(n8778) );
  XNOR U8687 ( .A(n8774), .B(n8773), .Z(n8785) );
  XOR U8688 ( .A(n8814), .B(n8770), .Z(n8773) );
  XNOR U8689 ( .A(n6439), .B(p_input[362]), .Z(n8770) );
  XNOR U8690 ( .A(p_input[2059]), .B(p_input[363]), .Z(n8814) );
  XOR U8691 ( .A(p_input[2060]), .B(p_input[364]), .Z(n8774) );
  XNOR U8692 ( .A(n8784), .B(n8775), .Z(n8813) );
  XNOR U8693 ( .A(n6553), .B(p_input[353]), .Z(n8775) );
  XOR U8694 ( .A(n8815), .B(n8790), .Z(n8784) );
  XNOR U8695 ( .A(p_input[2063]), .B(p_input[367]), .Z(n8790) );
  XOR U8696 ( .A(n8781), .B(n8789), .Z(n8815) );
  XOR U8697 ( .A(n8816), .B(n8786), .Z(n8789) );
  XOR U8698 ( .A(p_input[2061]), .B(p_input[365]), .Z(n8786) );
  XNOR U8699 ( .A(p_input[2062]), .B(p_input[366]), .Z(n8816) );
  XNOR U8700 ( .A(n6325), .B(p_input[361]), .Z(n8781) );
  XNOR U8701 ( .A(n8797), .B(n8796), .Z(n8779) );
  XNOR U8702 ( .A(n8817), .B(n8802), .Z(n8796) );
  XOR U8703 ( .A(p_input[2056]), .B(p_input[360]), .Z(n8802) );
  XOR U8704 ( .A(n8793), .B(n8801), .Z(n8817) );
  XOR U8705 ( .A(n8818), .B(n8798), .Z(n8801) );
  XOR U8706 ( .A(p_input[2054]), .B(p_input[358]), .Z(n8798) );
  XNOR U8707 ( .A(p_input[2055]), .B(p_input[359]), .Z(n8818) );
  XNOR U8708 ( .A(n6328), .B(p_input[354]), .Z(n8793) );
  XNOR U8709 ( .A(n8807), .B(n8806), .Z(n8797) );
  XOR U8710 ( .A(n8819), .B(n8803), .Z(n8806) );
  XOR U8711 ( .A(p_input[2051]), .B(p_input[355]), .Z(n8803) );
  XNOR U8712 ( .A(p_input[2052]), .B(p_input[356]), .Z(n8819) );
  XOR U8713 ( .A(p_input[2053]), .B(p_input[357]), .Z(n8807) );
  XOR U8714 ( .A(n8820), .B(n8821), .Z(n8708) );
  AND U8715 ( .A(n95), .B(n8822), .Z(n8821) );
  XNOR U8716 ( .A(n8823), .B(n8820), .Z(n8822) );
  XNOR U8717 ( .A(n8824), .B(n8825), .Z(n95) );
  AND U8718 ( .A(n8826), .B(n8827), .Z(n8825) );
  XOR U8719 ( .A(n8721), .B(n8824), .Z(n8827) );
  AND U8720 ( .A(n8828), .B(n8829), .Z(n8721) );
  XNOR U8721 ( .A(n8718), .B(n8824), .Z(n8826) );
  XOR U8722 ( .A(n8830), .B(n8831), .Z(n8718) );
  AND U8723 ( .A(n99), .B(n8832), .Z(n8831) );
  XOR U8724 ( .A(n8833), .B(n8830), .Z(n8832) );
  XOR U8725 ( .A(n8834), .B(n8835), .Z(n8824) );
  AND U8726 ( .A(n8836), .B(n8837), .Z(n8835) );
  XNOR U8727 ( .A(n8834), .B(n8828), .Z(n8837) );
  IV U8728 ( .A(n8736), .Z(n8828) );
  XOR U8729 ( .A(n8838), .B(n8839), .Z(n8736) );
  XOR U8730 ( .A(n8840), .B(n8829), .Z(n8839) );
  AND U8731 ( .A(n8763), .B(n8841), .Z(n8829) );
  AND U8732 ( .A(n8842), .B(n8843), .Z(n8840) );
  XOR U8733 ( .A(n8844), .B(n8838), .Z(n8842) );
  XNOR U8734 ( .A(n8733), .B(n8834), .Z(n8836) );
  XOR U8735 ( .A(n8845), .B(n8846), .Z(n8733) );
  AND U8736 ( .A(n99), .B(n8847), .Z(n8846) );
  XOR U8737 ( .A(n8848), .B(n8845), .Z(n8847) );
  XOR U8738 ( .A(n8849), .B(n8850), .Z(n8834) );
  AND U8739 ( .A(n8851), .B(n8852), .Z(n8850) );
  XNOR U8740 ( .A(n8849), .B(n8763), .Z(n8852) );
  XOR U8741 ( .A(n8853), .B(n8843), .Z(n8763) );
  XNOR U8742 ( .A(n8854), .B(n8838), .Z(n8843) );
  XOR U8743 ( .A(n8855), .B(n8856), .Z(n8838) );
  AND U8744 ( .A(n8857), .B(n8858), .Z(n8856) );
  XOR U8745 ( .A(n8859), .B(n8855), .Z(n8857) );
  XNOR U8746 ( .A(n8860), .B(n8861), .Z(n8854) );
  AND U8747 ( .A(n8862), .B(n8863), .Z(n8861) );
  XOR U8748 ( .A(n8860), .B(n8864), .Z(n8862) );
  XNOR U8749 ( .A(n8844), .B(n8841), .Z(n8853) );
  AND U8750 ( .A(n8865), .B(n8866), .Z(n8841) );
  XOR U8751 ( .A(n8867), .B(n8868), .Z(n8844) );
  AND U8752 ( .A(n8869), .B(n8870), .Z(n8868) );
  XOR U8753 ( .A(n8867), .B(n8871), .Z(n8869) );
  XNOR U8754 ( .A(n8760), .B(n8849), .Z(n8851) );
  XOR U8755 ( .A(n8872), .B(n8873), .Z(n8760) );
  AND U8756 ( .A(n99), .B(n8874), .Z(n8873) );
  XNOR U8757 ( .A(n8875), .B(n8872), .Z(n8874) );
  XOR U8758 ( .A(n8876), .B(n8877), .Z(n8849) );
  AND U8759 ( .A(n8878), .B(n8879), .Z(n8877) );
  XNOR U8760 ( .A(n8876), .B(n8865), .Z(n8879) );
  IV U8761 ( .A(n8811), .Z(n8865) );
  XNOR U8762 ( .A(n8880), .B(n8858), .Z(n8811) );
  XNOR U8763 ( .A(n8881), .B(n8864), .Z(n8858) );
  XOR U8764 ( .A(n8882), .B(n8883), .Z(n8864) );
  NOR U8765 ( .A(n8884), .B(n8885), .Z(n8883) );
  XNOR U8766 ( .A(n8882), .B(n8886), .Z(n8884) );
  XNOR U8767 ( .A(n8863), .B(n8855), .Z(n8881) );
  XOR U8768 ( .A(n8887), .B(n8888), .Z(n8855) );
  AND U8769 ( .A(n8889), .B(n8890), .Z(n8888) );
  XNOR U8770 ( .A(n8887), .B(n8891), .Z(n8889) );
  XNOR U8771 ( .A(n8892), .B(n8860), .Z(n8863) );
  XOR U8772 ( .A(n8893), .B(n8894), .Z(n8860) );
  AND U8773 ( .A(n8895), .B(n8896), .Z(n8894) );
  XOR U8774 ( .A(n8893), .B(n8897), .Z(n8895) );
  XNOR U8775 ( .A(n8898), .B(n8899), .Z(n8892) );
  NOR U8776 ( .A(n8900), .B(n8901), .Z(n8899) );
  XOR U8777 ( .A(n8898), .B(n8902), .Z(n8900) );
  XNOR U8778 ( .A(n8859), .B(n8866), .Z(n8880) );
  NOR U8779 ( .A(n8823), .B(n8903), .Z(n8866) );
  XOR U8780 ( .A(n8871), .B(n8870), .Z(n8859) );
  XNOR U8781 ( .A(n8904), .B(n8867), .Z(n8870) );
  XOR U8782 ( .A(n8905), .B(n8906), .Z(n8867) );
  AND U8783 ( .A(n8907), .B(n8908), .Z(n8906) );
  XOR U8784 ( .A(n8905), .B(n8909), .Z(n8907) );
  XNOR U8785 ( .A(n8910), .B(n8911), .Z(n8904) );
  NOR U8786 ( .A(n8912), .B(n8913), .Z(n8911) );
  XNOR U8787 ( .A(n8910), .B(n8914), .Z(n8912) );
  XOR U8788 ( .A(n8915), .B(n8916), .Z(n8871) );
  NOR U8789 ( .A(n8917), .B(n8918), .Z(n8916) );
  XNOR U8790 ( .A(n8915), .B(n8919), .Z(n8917) );
  XNOR U8791 ( .A(n8808), .B(n8876), .Z(n8878) );
  XOR U8792 ( .A(n8920), .B(n8921), .Z(n8808) );
  AND U8793 ( .A(n99), .B(n8922), .Z(n8921) );
  XOR U8794 ( .A(n8923), .B(n8920), .Z(n8922) );
  AND U8795 ( .A(n8820), .B(n8823), .Z(n8876) );
  XOR U8796 ( .A(n8924), .B(n8903), .Z(n8823) );
  XNOR U8797 ( .A(p_input[2048]), .B(p_input[368]), .Z(n8903) );
  XOR U8798 ( .A(n8891), .B(n8890), .Z(n8924) );
  XNOR U8799 ( .A(n8925), .B(n8897), .Z(n8890) );
  XNOR U8800 ( .A(n8886), .B(n8885), .Z(n8897) );
  XOR U8801 ( .A(n8926), .B(n8882), .Z(n8885) );
  XNOR U8802 ( .A(n6439), .B(p_input[378]), .Z(n8882) );
  XNOR U8803 ( .A(p_input[2059]), .B(p_input[379]), .Z(n8926) );
  XOR U8804 ( .A(p_input[2060]), .B(p_input[380]), .Z(n8886) );
  XNOR U8805 ( .A(n8896), .B(n8887), .Z(n8925) );
  XNOR U8806 ( .A(n6553), .B(p_input[369]), .Z(n8887) );
  XOR U8807 ( .A(n8927), .B(n8902), .Z(n8896) );
  XNOR U8808 ( .A(p_input[2063]), .B(p_input[383]), .Z(n8902) );
  XOR U8809 ( .A(n8893), .B(n8901), .Z(n8927) );
  XOR U8810 ( .A(n8928), .B(n8898), .Z(n8901) );
  XOR U8811 ( .A(p_input[2061]), .B(p_input[381]), .Z(n8898) );
  XNOR U8812 ( .A(p_input[2062]), .B(p_input[382]), .Z(n8928) );
  XNOR U8813 ( .A(n6325), .B(p_input[377]), .Z(n8893) );
  XNOR U8814 ( .A(n8909), .B(n8908), .Z(n8891) );
  XNOR U8815 ( .A(n8929), .B(n8914), .Z(n8908) );
  XOR U8816 ( .A(p_input[2056]), .B(p_input[376]), .Z(n8914) );
  XOR U8817 ( .A(n8905), .B(n8913), .Z(n8929) );
  XOR U8818 ( .A(n8930), .B(n8910), .Z(n8913) );
  XOR U8819 ( .A(p_input[2054]), .B(p_input[374]), .Z(n8910) );
  XNOR U8820 ( .A(p_input[2055]), .B(p_input[375]), .Z(n8930) );
  XNOR U8821 ( .A(n6328), .B(p_input[370]), .Z(n8905) );
  XNOR U8822 ( .A(n8919), .B(n8918), .Z(n8909) );
  XOR U8823 ( .A(n8931), .B(n8915), .Z(n8918) );
  XOR U8824 ( .A(p_input[2051]), .B(p_input[371]), .Z(n8915) );
  XNOR U8825 ( .A(p_input[2052]), .B(p_input[372]), .Z(n8931) );
  XOR U8826 ( .A(p_input[2053]), .B(p_input[373]), .Z(n8919) );
  XOR U8827 ( .A(n8932), .B(n8933), .Z(n8820) );
  AND U8828 ( .A(n99), .B(n8934), .Z(n8933) );
  XNOR U8829 ( .A(n8935), .B(n8932), .Z(n8934) );
  XNOR U8830 ( .A(n8936), .B(n8937), .Z(n99) );
  AND U8831 ( .A(n8938), .B(n8939), .Z(n8937) );
  XOR U8832 ( .A(n8833), .B(n8936), .Z(n8939) );
  AND U8833 ( .A(n8940), .B(n8941), .Z(n8833) );
  XNOR U8834 ( .A(n8830), .B(n8936), .Z(n8938) );
  XOR U8835 ( .A(n8942), .B(n8943), .Z(n8830) );
  AND U8836 ( .A(n103), .B(n8944), .Z(n8943) );
  XOR U8837 ( .A(n8945), .B(n8942), .Z(n8944) );
  XOR U8838 ( .A(n8946), .B(n8947), .Z(n8936) );
  AND U8839 ( .A(n8948), .B(n8949), .Z(n8947) );
  XNOR U8840 ( .A(n8946), .B(n8940), .Z(n8949) );
  IV U8841 ( .A(n8848), .Z(n8940) );
  XOR U8842 ( .A(n8950), .B(n8951), .Z(n8848) );
  XOR U8843 ( .A(n8952), .B(n8941), .Z(n8951) );
  AND U8844 ( .A(n8875), .B(n8953), .Z(n8941) );
  AND U8845 ( .A(n8954), .B(n8955), .Z(n8952) );
  XOR U8846 ( .A(n8956), .B(n8950), .Z(n8954) );
  XNOR U8847 ( .A(n8845), .B(n8946), .Z(n8948) );
  XOR U8848 ( .A(n8957), .B(n8958), .Z(n8845) );
  AND U8849 ( .A(n103), .B(n8959), .Z(n8958) );
  XOR U8850 ( .A(n8960), .B(n8957), .Z(n8959) );
  XOR U8851 ( .A(n8961), .B(n8962), .Z(n8946) );
  AND U8852 ( .A(n8963), .B(n8964), .Z(n8962) );
  XNOR U8853 ( .A(n8961), .B(n8875), .Z(n8964) );
  XOR U8854 ( .A(n8965), .B(n8955), .Z(n8875) );
  XNOR U8855 ( .A(n8966), .B(n8950), .Z(n8955) );
  XOR U8856 ( .A(n8967), .B(n8968), .Z(n8950) );
  AND U8857 ( .A(n8969), .B(n8970), .Z(n8968) );
  XOR U8858 ( .A(n8971), .B(n8967), .Z(n8969) );
  XNOR U8859 ( .A(n8972), .B(n8973), .Z(n8966) );
  AND U8860 ( .A(n8974), .B(n8975), .Z(n8973) );
  XOR U8861 ( .A(n8972), .B(n8976), .Z(n8974) );
  XNOR U8862 ( .A(n8956), .B(n8953), .Z(n8965) );
  AND U8863 ( .A(n8977), .B(n8978), .Z(n8953) );
  XOR U8864 ( .A(n8979), .B(n8980), .Z(n8956) );
  AND U8865 ( .A(n8981), .B(n8982), .Z(n8980) );
  XOR U8866 ( .A(n8979), .B(n8983), .Z(n8981) );
  XNOR U8867 ( .A(n8872), .B(n8961), .Z(n8963) );
  XOR U8868 ( .A(n8984), .B(n8985), .Z(n8872) );
  AND U8869 ( .A(n103), .B(n8986), .Z(n8985) );
  XNOR U8870 ( .A(n8987), .B(n8984), .Z(n8986) );
  XOR U8871 ( .A(n8988), .B(n8989), .Z(n8961) );
  AND U8872 ( .A(n8990), .B(n8991), .Z(n8989) );
  XNOR U8873 ( .A(n8988), .B(n8977), .Z(n8991) );
  IV U8874 ( .A(n8923), .Z(n8977) );
  XNOR U8875 ( .A(n8992), .B(n8970), .Z(n8923) );
  XNOR U8876 ( .A(n8993), .B(n8976), .Z(n8970) );
  XOR U8877 ( .A(n8994), .B(n8995), .Z(n8976) );
  NOR U8878 ( .A(n8996), .B(n8997), .Z(n8995) );
  XNOR U8879 ( .A(n8994), .B(n8998), .Z(n8996) );
  XNOR U8880 ( .A(n8975), .B(n8967), .Z(n8993) );
  XOR U8881 ( .A(n8999), .B(n9000), .Z(n8967) );
  AND U8882 ( .A(n9001), .B(n9002), .Z(n9000) );
  XNOR U8883 ( .A(n8999), .B(n9003), .Z(n9001) );
  XNOR U8884 ( .A(n9004), .B(n8972), .Z(n8975) );
  XOR U8885 ( .A(n9005), .B(n9006), .Z(n8972) );
  AND U8886 ( .A(n9007), .B(n9008), .Z(n9006) );
  XOR U8887 ( .A(n9005), .B(n9009), .Z(n9007) );
  XNOR U8888 ( .A(n9010), .B(n9011), .Z(n9004) );
  NOR U8889 ( .A(n9012), .B(n9013), .Z(n9011) );
  XOR U8890 ( .A(n9010), .B(n9014), .Z(n9012) );
  XNOR U8891 ( .A(n8971), .B(n8978), .Z(n8992) );
  NOR U8892 ( .A(n8935), .B(n9015), .Z(n8978) );
  XOR U8893 ( .A(n8983), .B(n8982), .Z(n8971) );
  XNOR U8894 ( .A(n9016), .B(n8979), .Z(n8982) );
  XOR U8895 ( .A(n9017), .B(n9018), .Z(n8979) );
  AND U8896 ( .A(n9019), .B(n9020), .Z(n9018) );
  XOR U8897 ( .A(n9017), .B(n9021), .Z(n9019) );
  XNOR U8898 ( .A(n9022), .B(n9023), .Z(n9016) );
  NOR U8899 ( .A(n9024), .B(n9025), .Z(n9023) );
  XNOR U8900 ( .A(n9022), .B(n9026), .Z(n9024) );
  XOR U8901 ( .A(n9027), .B(n9028), .Z(n8983) );
  NOR U8902 ( .A(n9029), .B(n9030), .Z(n9028) );
  XNOR U8903 ( .A(n9027), .B(n9031), .Z(n9029) );
  XNOR U8904 ( .A(n8920), .B(n8988), .Z(n8990) );
  XOR U8905 ( .A(n9032), .B(n9033), .Z(n8920) );
  AND U8906 ( .A(n103), .B(n9034), .Z(n9033) );
  XOR U8907 ( .A(n9035), .B(n9032), .Z(n9034) );
  AND U8908 ( .A(n8932), .B(n8935), .Z(n8988) );
  XOR U8909 ( .A(n9036), .B(n9015), .Z(n8935) );
  XNOR U8910 ( .A(p_input[2048]), .B(p_input[384]), .Z(n9015) );
  XOR U8911 ( .A(n9003), .B(n9002), .Z(n9036) );
  XNOR U8912 ( .A(n9037), .B(n9009), .Z(n9002) );
  XNOR U8913 ( .A(n8998), .B(n8997), .Z(n9009) );
  XOR U8914 ( .A(n9038), .B(n8994), .Z(n8997) );
  XNOR U8915 ( .A(n6439), .B(p_input[394]), .Z(n8994) );
  XNOR U8916 ( .A(p_input[2059]), .B(p_input[395]), .Z(n9038) );
  XOR U8917 ( .A(p_input[2060]), .B(p_input[396]), .Z(n8998) );
  XNOR U8918 ( .A(n9008), .B(n8999), .Z(n9037) );
  XNOR U8919 ( .A(n6553), .B(p_input[385]), .Z(n8999) );
  XOR U8920 ( .A(n9039), .B(n9014), .Z(n9008) );
  XNOR U8921 ( .A(p_input[2063]), .B(p_input[399]), .Z(n9014) );
  XOR U8922 ( .A(n9005), .B(n9013), .Z(n9039) );
  XOR U8923 ( .A(n9040), .B(n9010), .Z(n9013) );
  XOR U8924 ( .A(p_input[2061]), .B(p_input[397]), .Z(n9010) );
  XNOR U8925 ( .A(p_input[2062]), .B(p_input[398]), .Z(n9040) );
  XNOR U8926 ( .A(n6325), .B(p_input[393]), .Z(n9005) );
  XNOR U8927 ( .A(n9021), .B(n9020), .Z(n9003) );
  XNOR U8928 ( .A(n9041), .B(n9026), .Z(n9020) );
  XOR U8929 ( .A(p_input[2056]), .B(p_input[392]), .Z(n9026) );
  XOR U8930 ( .A(n9017), .B(n9025), .Z(n9041) );
  XOR U8931 ( .A(n9042), .B(n9022), .Z(n9025) );
  XOR U8932 ( .A(p_input[2054]), .B(p_input[390]), .Z(n9022) );
  XNOR U8933 ( .A(p_input[2055]), .B(p_input[391]), .Z(n9042) );
  XNOR U8934 ( .A(n6328), .B(p_input[386]), .Z(n9017) );
  XNOR U8935 ( .A(n9031), .B(n9030), .Z(n9021) );
  XOR U8936 ( .A(n9043), .B(n9027), .Z(n9030) );
  XOR U8937 ( .A(p_input[2051]), .B(p_input[387]), .Z(n9027) );
  XNOR U8938 ( .A(p_input[2052]), .B(p_input[388]), .Z(n9043) );
  XOR U8939 ( .A(p_input[2053]), .B(p_input[389]), .Z(n9031) );
  XOR U8940 ( .A(n9044), .B(n9045), .Z(n8932) );
  AND U8941 ( .A(n103), .B(n9046), .Z(n9045) );
  XNOR U8942 ( .A(n9047), .B(n9044), .Z(n9046) );
  XNOR U8943 ( .A(n9048), .B(n9049), .Z(n103) );
  AND U8944 ( .A(n9050), .B(n9051), .Z(n9049) );
  XOR U8945 ( .A(n8945), .B(n9048), .Z(n9051) );
  AND U8946 ( .A(n9052), .B(n9053), .Z(n8945) );
  XNOR U8947 ( .A(n8942), .B(n9048), .Z(n9050) );
  XOR U8948 ( .A(n9054), .B(n9055), .Z(n8942) );
  AND U8949 ( .A(n107), .B(n9056), .Z(n9055) );
  XOR U8950 ( .A(n9057), .B(n9054), .Z(n9056) );
  XOR U8951 ( .A(n9058), .B(n9059), .Z(n9048) );
  AND U8952 ( .A(n9060), .B(n9061), .Z(n9059) );
  XNOR U8953 ( .A(n9058), .B(n9052), .Z(n9061) );
  IV U8954 ( .A(n8960), .Z(n9052) );
  XOR U8955 ( .A(n9062), .B(n9063), .Z(n8960) );
  XOR U8956 ( .A(n9064), .B(n9053), .Z(n9063) );
  AND U8957 ( .A(n8987), .B(n9065), .Z(n9053) );
  AND U8958 ( .A(n9066), .B(n9067), .Z(n9064) );
  XOR U8959 ( .A(n9068), .B(n9062), .Z(n9066) );
  XNOR U8960 ( .A(n8957), .B(n9058), .Z(n9060) );
  XOR U8961 ( .A(n9069), .B(n9070), .Z(n8957) );
  AND U8962 ( .A(n107), .B(n9071), .Z(n9070) );
  XOR U8963 ( .A(n9072), .B(n9069), .Z(n9071) );
  XOR U8964 ( .A(n9073), .B(n9074), .Z(n9058) );
  AND U8965 ( .A(n9075), .B(n9076), .Z(n9074) );
  XNOR U8966 ( .A(n9073), .B(n8987), .Z(n9076) );
  XOR U8967 ( .A(n9077), .B(n9067), .Z(n8987) );
  XNOR U8968 ( .A(n9078), .B(n9062), .Z(n9067) );
  XOR U8969 ( .A(n9079), .B(n9080), .Z(n9062) );
  AND U8970 ( .A(n9081), .B(n9082), .Z(n9080) );
  XOR U8971 ( .A(n9083), .B(n9079), .Z(n9081) );
  XNOR U8972 ( .A(n9084), .B(n9085), .Z(n9078) );
  AND U8973 ( .A(n9086), .B(n9087), .Z(n9085) );
  XOR U8974 ( .A(n9084), .B(n9088), .Z(n9086) );
  XNOR U8975 ( .A(n9068), .B(n9065), .Z(n9077) );
  AND U8976 ( .A(n9089), .B(n9090), .Z(n9065) );
  XOR U8977 ( .A(n9091), .B(n9092), .Z(n9068) );
  AND U8978 ( .A(n9093), .B(n9094), .Z(n9092) );
  XOR U8979 ( .A(n9091), .B(n9095), .Z(n9093) );
  XNOR U8980 ( .A(n8984), .B(n9073), .Z(n9075) );
  XOR U8981 ( .A(n9096), .B(n9097), .Z(n8984) );
  AND U8982 ( .A(n107), .B(n9098), .Z(n9097) );
  XNOR U8983 ( .A(n9099), .B(n9096), .Z(n9098) );
  XOR U8984 ( .A(n9100), .B(n9101), .Z(n9073) );
  AND U8985 ( .A(n9102), .B(n9103), .Z(n9101) );
  XNOR U8986 ( .A(n9100), .B(n9089), .Z(n9103) );
  IV U8987 ( .A(n9035), .Z(n9089) );
  XNOR U8988 ( .A(n9104), .B(n9082), .Z(n9035) );
  XNOR U8989 ( .A(n9105), .B(n9088), .Z(n9082) );
  XOR U8990 ( .A(n9106), .B(n9107), .Z(n9088) );
  NOR U8991 ( .A(n9108), .B(n9109), .Z(n9107) );
  XNOR U8992 ( .A(n9106), .B(n9110), .Z(n9108) );
  XNOR U8993 ( .A(n9087), .B(n9079), .Z(n9105) );
  XOR U8994 ( .A(n9111), .B(n9112), .Z(n9079) );
  AND U8995 ( .A(n9113), .B(n9114), .Z(n9112) );
  XNOR U8996 ( .A(n9111), .B(n9115), .Z(n9113) );
  XNOR U8997 ( .A(n9116), .B(n9084), .Z(n9087) );
  XOR U8998 ( .A(n9117), .B(n9118), .Z(n9084) );
  AND U8999 ( .A(n9119), .B(n9120), .Z(n9118) );
  XOR U9000 ( .A(n9117), .B(n9121), .Z(n9119) );
  XNOR U9001 ( .A(n9122), .B(n9123), .Z(n9116) );
  NOR U9002 ( .A(n9124), .B(n9125), .Z(n9123) );
  XOR U9003 ( .A(n9122), .B(n9126), .Z(n9124) );
  XNOR U9004 ( .A(n9083), .B(n9090), .Z(n9104) );
  NOR U9005 ( .A(n9047), .B(n9127), .Z(n9090) );
  XOR U9006 ( .A(n9095), .B(n9094), .Z(n9083) );
  XNOR U9007 ( .A(n9128), .B(n9091), .Z(n9094) );
  XOR U9008 ( .A(n9129), .B(n9130), .Z(n9091) );
  AND U9009 ( .A(n9131), .B(n9132), .Z(n9130) );
  XOR U9010 ( .A(n9129), .B(n9133), .Z(n9131) );
  XNOR U9011 ( .A(n9134), .B(n9135), .Z(n9128) );
  NOR U9012 ( .A(n9136), .B(n9137), .Z(n9135) );
  XNOR U9013 ( .A(n9134), .B(n9138), .Z(n9136) );
  XOR U9014 ( .A(n9139), .B(n9140), .Z(n9095) );
  NOR U9015 ( .A(n9141), .B(n9142), .Z(n9140) );
  XNOR U9016 ( .A(n9139), .B(n9143), .Z(n9141) );
  XNOR U9017 ( .A(n9032), .B(n9100), .Z(n9102) );
  XOR U9018 ( .A(n9144), .B(n9145), .Z(n9032) );
  AND U9019 ( .A(n107), .B(n9146), .Z(n9145) );
  XOR U9020 ( .A(n9147), .B(n9144), .Z(n9146) );
  AND U9021 ( .A(n9044), .B(n9047), .Z(n9100) );
  XOR U9022 ( .A(n9148), .B(n9127), .Z(n9047) );
  XNOR U9023 ( .A(p_input[2048]), .B(p_input[400]), .Z(n9127) );
  XOR U9024 ( .A(n9115), .B(n9114), .Z(n9148) );
  XNOR U9025 ( .A(n9149), .B(n9121), .Z(n9114) );
  XNOR U9026 ( .A(n9110), .B(n9109), .Z(n9121) );
  XOR U9027 ( .A(n9150), .B(n9106), .Z(n9109) );
  XNOR U9028 ( .A(n6439), .B(p_input[410]), .Z(n9106) );
  XNOR U9029 ( .A(p_input[2059]), .B(p_input[411]), .Z(n9150) );
  XOR U9030 ( .A(p_input[2060]), .B(p_input[412]), .Z(n9110) );
  XNOR U9031 ( .A(n9120), .B(n9111), .Z(n9149) );
  XNOR U9032 ( .A(n6553), .B(p_input[401]), .Z(n9111) );
  XOR U9033 ( .A(n9151), .B(n9126), .Z(n9120) );
  XNOR U9034 ( .A(p_input[2063]), .B(p_input[415]), .Z(n9126) );
  XOR U9035 ( .A(n9117), .B(n9125), .Z(n9151) );
  XOR U9036 ( .A(n9152), .B(n9122), .Z(n9125) );
  XOR U9037 ( .A(p_input[2061]), .B(p_input[413]), .Z(n9122) );
  XNOR U9038 ( .A(p_input[2062]), .B(p_input[414]), .Z(n9152) );
  XNOR U9039 ( .A(n6325), .B(p_input[409]), .Z(n9117) );
  XNOR U9040 ( .A(n9133), .B(n9132), .Z(n9115) );
  XNOR U9041 ( .A(n9153), .B(n9138), .Z(n9132) );
  XOR U9042 ( .A(p_input[2056]), .B(p_input[408]), .Z(n9138) );
  XOR U9043 ( .A(n9129), .B(n9137), .Z(n9153) );
  XOR U9044 ( .A(n9154), .B(n9134), .Z(n9137) );
  XOR U9045 ( .A(p_input[2054]), .B(p_input[406]), .Z(n9134) );
  XNOR U9046 ( .A(p_input[2055]), .B(p_input[407]), .Z(n9154) );
  XNOR U9047 ( .A(n6328), .B(p_input[402]), .Z(n9129) );
  XNOR U9048 ( .A(n9143), .B(n9142), .Z(n9133) );
  XOR U9049 ( .A(n9155), .B(n9139), .Z(n9142) );
  XOR U9050 ( .A(p_input[2051]), .B(p_input[403]), .Z(n9139) );
  XNOR U9051 ( .A(p_input[2052]), .B(p_input[404]), .Z(n9155) );
  XOR U9052 ( .A(p_input[2053]), .B(p_input[405]), .Z(n9143) );
  XOR U9053 ( .A(n9156), .B(n9157), .Z(n9044) );
  AND U9054 ( .A(n107), .B(n9158), .Z(n9157) );
  XNOR U9055 ( .A(n9159), .B(n9156), .Z(n9158) );
  XNOR U9056 ( .A(n9160), .B(n9161), .Z(n107) );
  AND U9057 ( .A(n9162), .B(n9163), .Z(n9161) );
  XOR U9058 ( .A(n9057), .B(n9160), .Z(n9163) );
  AND U9059 ( .A(n9164), .B(n9165), .Z(n9057) );
  XNOR U9060 ( .A(n9054), .B(n9160), .Z(n9162) );
  XOR U9061 ( .A(n9166), .B(n9167), .Z(n9054) );
  AND U9062 ( .A(n111), .B(n9168), .Z(n9167) );
  XOR U9063 ( .A(n9169), .B(n9166), .Z(n9168) );
  XOR U9064 ( .A(n9170), .B(n9171), .Z(n9160) );
  AND U9065 ( .A(n9172), .B(n9173), .Z(n9171) );
  XNOR U9066 ( .A(n9170), .B(n9164), .Z(n9173) );
  IV U9067 ( .A(n9072), .Z(n9164) );
  XOR U9068 ( .A(n9174), .B(n9175), .Z(n9072) );
  XOR U9069 ( .A(n9176), .B(n9165), .Z(n9175) );
  AND U9070 ( .A(n9099), .B(n9177), .Z(n9165) );
  AND U9071 ( .A(n9178), .B(n9179), .Z(n9176) );
  XOR U9072 ( .A(n9180), .B(n9174), .Z(n9178) );
  XNOR U9073 ( .A(n9069), .B(n9170), .Z(n9172) );
  XOR U9074 ( .A(n9181), .B(n9182), .Z(n9069) );
  AND U9075 ( .A(n111), .B(n9183), .Z(n9182) );
  XOR U9076 ( .A(n9184), .B(n9181), .Z(n9183) );
  XOR U9077 ( .A(n9185), .B(n9186), .Z(n9170) );
  AND U9078 ( .A(n9187), .B(n9188), .Z(n9186) );
  XNOR U9079 ( .A(n9185), .B(n9099), .Z(n9188) );
  XOR U9080 ( .A(n9189), .B(n9179), .Z(n9099) );
  XNOR U9081 ( .A(n9190), .B(n9174), .Z(n9179) );
  XOR U9082 ( .A(n9191), .B(n9192), .Z(n9174) );
  AND U9083 ( .A(n9193), .B(n9194), .Z(n9192) );
  XOR U9084 ( .A(n9195), .B(n9191), .Z(n9193) );
  XNOR U9085 ( .A(n9196), .B(n9197), .Z(n9190) );
  AND U9086 ( .A(n9198), .B(n9199), .Z(n9197) );
  XOR U9087 ( .A(n9196), .B(n9200), .Z(n9198) );
  XNOR U9088 ( .A(n9180), .B(n9177), .Z(n9189) );
  AND U9089 ( .A(n9201), .B(n9202), .Z(n9177) );
  XOR U9090 ( .A(n9203), .B(n9204), .Z(n9180) );
  AND U9091 ( .A(n9205), .B(n9206), .Z(n9204) );
  XOR U9092 ( .A(n9203), .B(n9207), .Z(n9205) );
  XNOR U9093 ( .A(n9096), .B(n9185), .Z(n9187) );
  XOR U9094 ( .A(n9208), .B(n9209), .Z(n9096) );
  AND U9095 ( .A(n111), .B(n9210), .Z(n9209) );
  XNOR U9096 ( .A(n9211), .B(n9208), .Z(n9210) );
  XOR U9097 ( .A(n9212), .B(n9213), .Z(n9185) );
  AND U9098 ( .A(n9214), .B(n9215), .Z(n9213) );
  XNOR U9099 ( .A(n9212), .B(n9201), .Z(n9215) );
  IV U9100 ( .A(n9147), .Z(n9201) );
  XNOR U9101 ( .A(n9216), .B(n9194), .Z(n9147) );
  XNOR U9102 ( .A(n9217), .B(n9200), .Z(n9194) );
  XOR U9103 ( .A(n9218), .B(n9219), .Z(n9200) );
  NOR U9104 ( .A(n9220), .B(n9221), .Z(n9219) );
  XNOR U9105 ( .A(n9218), .B(n9222), .Z(n9220) );
  XNOR U9106 ( .A(n9199), .B(n9191), .Z(n9217) );
  XOR U9107 ( .A(n9223), .B(n9224), .Z(n9191) );
  AND U9108 ( .A(n9225), .B(n9226), .Z(n9224) );
  XNOR U9109 ( .A(n9223), .B(n9227), .Z(n9225) );
  XNOR U9110 ( .A(n9228), .B(n9196), .Z(n9199) );
  XOR U9111 ( .A(n9229), .B(n9230), .Z(n9196) );
  AND U9112 ( .A(n9231), .B(n9232), .Z(n9230) );
  XOR U9113 ( .A(n9229), .B(n9233), .Z(n9231) );
  XNOR U9114 ( .A(n9234), .B(n9235), .Z(n9228) );
  NOR U9115 ( .A(n9236), .B(n9237), .Z(n9235) );
  XOR U9116 ( .A(n9234), .B(n9238), .Z(n9236) );
  XNOR U9117 ( .A(n9195), .B(n9202), .Z(n9216) );
  NOR U9118 ( .A(n9159), .B(n9239), .Z(n9202) );
  XOR U9119 ( .A(n9207), .B(n9206), .Z(n9195) );
  XNOR U9120 ( .A(n9240), .B(n9203), .Z(n9206) );
  XOR U9121 ( .A(n9241), .B(n9242), .Z(n9203) );
  AND U9122 ( .A(n9243), .B(n9244), .Z(n9242) );
  XOR U9123 ( .A(n9241), .B(n9245), .Z(n9243) );
  XNOR U9124 ( .A(n9246), .B(n9247), .Z(n9240) );
  NOR U9125 ( .A(n9248), .B(n9249), .Z(n9247) );
  XNOR U9126 ( .A(n9246), .B(n9250), .Z(n9248) );
  XOR U9127 ( .A(n9251), .B(n9252), .Z(n9207) );
  NOR U9128 ( .A(n9253), .B(n9254), .Z(n9252) );
  XNOR U9129 ( .A(n9251), .B(n9255), .Z(n9253) );
  XNOR U9130 ( .A(n9144), .B(n9212), .Z(n9214) );
  XOR U9131 ( .A(n9256), .B(n9257), .Z(n9144) );
  AND U9132 ( .A(n111), .B(n9258), .Z(n9257) );
  XOR U9133 ( .A(n9259), .B(n9256), .Z(n9258) );
  AND U9134 ( .A(n9156), .B(n9159), .Z(n9212) );
  XOR U9135 ( .A(n9260), .B(n9239), .Z(n9159) );
  XNOR U9136 ( .A(p_input[2048]), .B(p_input[416]), .Z(n9239) );
  XOR U9137 ( .A(n9227), .B(n9226), .Z(n9260) );
  XNOR U9138 ( .A(n9261), .B(n9233), .Z(n9226) );
  XNOR U9139 ( .A(n9222), .B(n9221), .Z(n9233) );
  XOR U9140 ( .A(n9262), .B(n9218), .Z(n9221) );
  XNOR U9141 ( .A(n6439), .B(p_input[426]), .Z(n9218) );
  XNOR U9142 ( .A(p_input[2059]), .B(p_input[427]), .Z(n9262) );
  XOR U9143 ( .A(p_input[2060]), .B(p_input[428]), .Z(n9222) );
  XNOR U9144 ( .A(n9232), .B(n9223), .Z(n9261) );
  XNOR U9145 ( .A(n6553), .B(p_input[417]), .Z(n9223) );
  XOR U9146 ( .A(n9263), .B(n9238), .Z(n9232) );
  XNOR U9147 ( .A(p_input[2063]), .B(p_input[431]), .Z(n9238) );
  XOR U9148 ( .A(n9229), .B(n9237), .Z(n9263) );
  XOR U9149 ( .A(n9264), .B(n9234), .Z(n9237) );
  XOR U9150 ( .A(p_input[2061]), .B(p_input[429]), .Z(n9234) );
  XNOR U9151 ( .A(p_input[2062]), .B(p_input[430]), .Z(n9264) );
  XNOR U9152 ( .A(n6325), .B(p_input[425]), .Z(n9229) );
  XNOR U9153 ( .A(n9245), .B(n9244), .Z(n9227) );
  XNOR U9154 ( .A(n9265), .B(n9250), .Z(n9244) );
  XOR U9155 ( .A(p_input[2056]), .B(p_input[424]), .Z(n9250) );
  XOR U9156 ( .A(n9241), .B(n9249), .Z(n9265) );
  XOR U9157 ( .A(n9266), .B(n9246), .Z(n9249) );
  XOR U9158 ( .A(p_input[2054]), .B(p_input[422]), .Z(n9246) );
  XNOR U9159 ( .A(p_input[2055]), .B(p_input[423]), .Z(n9266) );
  XNOR U9160 ( .A(n6328), .B(p_input[418]), .Z(n9241) );
  XNOR U9161 ( .A(n9255), .B(n9254), .Z(n9245) );
  XOR U9162 ( .A(n9267), .B(n9251), .Z(n9254) );
  XOR U9163 ( .A(p_input[2051]), .B(p_input[419]), .Z(n9251) );
  XNOR U9164 ( .A(p_input[2052]), .B(p_input[420]), .Z(n9267) );
  XOR U9165 ( .A(p_input[2053]), .B(p_input[421]), .Z(n9255) );
  XOR U9166 ( .A(n9268), .B(n9269), .Z(n9156) );
  AND U9167 ( .A(n111), .B(n9270), .Z(n9269) );
  XNOR U9168 ( .A(n9271), .B(n9268), .Z(n9270) );
  XNOR U9169 ( .A(n9272), .B(n9273), .Z(n111) );
  AND U9170 ( .A(n9274), .B(n9275), .Z(n9273) );
  XOR U9171 ( .A(n9169), .B(n9272), .Z(n9275) );
  AND U9172 ( .A(n9276), .B(n9277), .Z(n9169) );
  XNOR U9173 ( .A(n9166), .B(n9272), .Z(n9274) );
  XOR U9174 ( .A(n9278), .B(n9279), .Z(n9166) );
  AND U9175 ( .A(n115), .B(n9280), .Z(n9279) );
  XOR U9176 ( .A(n9281), .B(n9278), .Z(n9280) );
  XOR U9177 ( .A(n9282), .B(n9283), .Z(n9272) );
  AND U9178 ( .A(n9284), .B(n9285), .Z(n9283) );
  XNOR U9179 ( .A(n9282), .B(n9276), .Z(n9285) );
  IV U9180 ( .A(n9184), .Z(n9276) );
  XOR U9181 ( .A(n9286), .B(n9287), .Z(n9184) );
  XOR U9182 ( .A(n9288), .B(n9277), .Z(n9287) );
  AND U9183 ( .A(n9211), .B(n9289), .Z(n9277) );
  AND U9184 ( .A(n9290), .B(n9291), .Z(n9288) );
  XOR U9185 ( .A(n9292), .B(n9286), .Z(n9290) );
  XNOR U9186 ( .A(n9181), .B(n9282), .Z(n9284) );
  XOR U9187 ( .A(n9293), .B(n9294), .Z(n9181) );
  AND U9188 ( .A(n115), .B(n9295), .Z(n9294) );
  XOR U9189 ( .A(n9296), .B(n9293), .Z(n9295) );
  XOR U9190 ( .A(n9297), .B(n9298), .Z(n9282) );
  AND U9191 ( .A(n9299), .B(n9300), .Z(n9298) );
  XNOR U9192 ( .A(n9297), .B(n9211), .Z(n9300) );
  XOR U9193 ( .A(n9301), .B(n9291), .Z(n9211) );
  XNOR U9194 ( .A(n9302), .B(n9286), .Z(n9291) );
  XOR U9195 ( .A(n9303), .B(n9304), .Z(n9286) );
  AND U9196 ( .A(n9305), .B(n9306), .Z(n9304) );
  XOR U9197 ( .A(n9307), .B(n9303), .Z(n9305) );
  XNOR U9198 ( .A(n9308), .B(n9309), .Z(n9302) );
  AND U9199 ( .A(n9310), .B(n9311), .Z(n9309) );
  XOR U9200 ( .A(n9308), .B(n9312), .Z(n9310) );
  XNOR U9201 ( .A(n9292), .B(n9289), .Z(n9301) );
  AND U9202 ( .A(n9313), .B(n9314), .Z(n9289) );
  XOR U9203 ( .A(n9315), .B(n9316), .Z(n9292) );
  AND U9204 ( .A(n9317), .B(n9318), .Z(n9316) );
  XOR U9205 ( .A(n9315), .B(n9319), .Z(n9317) );
  XNOR U9206 ( .A(n9208), .B(n9297), .Z(n9299) );
  XOR U9207 ( .A(n9320), .B(n9321), .Z(n9208) );
  AND U9208 ( .A(n115), .B(n9322), .Z(n9321) );
  XNOR U9209 ( .A(n9323), .B(n9320), .Z(n9322) );
  XOR U9210 ( .A(n9324), .B(n9325), .Z(n9297) );
  AND U9211 ( .A(n9326), .B(n9327), .Z(n9325) );
  XNOR U9212 ( .A(n9324), .B(n9313), .Z(n9327) );
  IV U9213 ( .A(n9259), .Z(n9313) );
  XNOR U9214 ( .A(n9328), .B(n9306), .Z(n9259) );
  XNOR U9215 ( .A(n9329), .B(n9312), .Z(n9306) );
  XOR U9216 ( .A(n9330), .B(n9331), .Z(n9312) );
  NOR U9217 ( .A(n9332), .B(n9333), .Z(n9331) );
  XNOR U9218 ( .A(n9330), .B(n9334), .Z(n9332) );
  XNOR U9219 ( .A(n9311), .B(n9303), .Z(n9329) );
  XOR U9220 ( .A(n9335), .B(n9336), .Z(n9303) );
  AND U9221 ( .A(n9337), .B(n9338), .Z(n9336) );
  XNOR U9222 ( .A(n9335), .B(n9339), .Z(n9337) );
  XNOR U9223 ( .A(n9340), .B(n9308), .Z(n9311) );
  XOR U9224 ( .A(n9341), .B(n9342), .Z(n9308) );
  AND U9225 ( .A(n9343), .B(n9344), .Z(n9342) );
  XOR U9226 ( .A(n9341), .B(n9345), .Z(n9343) );
  XNOR U9227 ( .A(n9346), .B(n9347), .Z(n9340) );
  NOR U9228 ( .A(n9348), .B(n9349), .Z(n9347) );
  XOR U9229 ( .A(n9346), .B(n9350), .Z(n9348) );
  XNOR U9230 ( .A(n9307), .B(n9314), .Z(n9328) );
  NOR U9231 ( .A(n9271), .B(n9351), .Z(n9314) );
  XOR U9232 ( .A(n9319), .B(n9318), .Z(n9307) );
  XNOR U9233 ( .A(n9352), .B(n9315), .Z(n9318) );
  XOR U9234 ( .A(n9353), .B(n9354), .Z(n9315) );
  AND U9235 ( .A(n9355), .B(n9356), .Z(n9354) );
  XOR U9236 ( .A(n9353), .B(n9357), .Z(n9355) );
  XNOR U9237 ( .A(n9358), .B(n9359), .Z(n9352) );
  NOR U9238 ( .A(n9360), .B(n9361), .Z(n9359) );
  XNOR U9239 ( .A(n9358), .B(n9362), .Z(n9360) );
  XOR U9240 ( .A(n9363), .B(n9364), .Z(n9319) );
  NOR U9241 ( .A(n9365), .B(n9366), .Z(n9364) );
  XNOR U9242 ( .A(n9363), .B(n9367), .Z(n9365) );
  XNOR U9243 ( .A(n9256), .B(n9324), .Z(n9326) );
  XOR U9244 ( .A(n9368), .B(n9369), .Z(n9256) );
  AND U9245 ( .A(n115), .B(n9370), .Z(n9369) );
  XOR U9246 ( .A(n9371), .B(n9368), .Z(n9370) );
  AND U9247 ( .A(n9268), .B(n9271), .Z(n9324) );
  XOR U9248 ( .A(n9372), .B(n9351), .Z(n9271) );
  XNOR U9249 ( .A(p_input[2048]), .B(p_input[432]), .Z(n9351) );
  XOR U9250 ( .A(n9339), .B(n9338), .Z(n9372) );
  XNOR U9251 ( .A(n9373), .B(n9345), .Z(n9338) );
  XNOR U9252 ( .A(n9334), .B(n9333), .Z(n9345) );
  XOR U9253 ( .A(n9374), .B(n9330), .Z(n9333) );
  XNOR U9254 ( .A(n6439), .B(p_input[442]), .Z(n9330) );
  XNOR U9255 ( .A(p_input[2059]), .B(p_input[443]), .Z(n9374) );
  XOR U9256 ( .A(p_input[2060]), .B(p_input[444]), .Z(n9334) );
  XNOR U9257 ( .A(n9344), .B(n9335), .Z(n9373) );
  XNOR U9258 ( .A(n6553), .B(p_input[433]), .Z(n9335) );
  XOR U9259 ( .A(n9375), .B(n9350), .Z(n9344) );
  XNOR U9260 ( .A(p_input[2063]), .B(p_input[447]), .Z(n9350) );
  XOR U9261 ( .A(n9341), .B(n9349), .Z(n9375) );
  XOR U9262 ( .A(n9376), .B(n9346), .Z(n9349) );
  XOR U9263 ( .A(p_input[2061]), .B(p_input[445]), .Z(n9346) );
  XNOR U9264 ( .A(p_input[2062]), .B(p_input[446]), .Z(n9376) );
  XNOR U9265 ( .A(n6325), .B(p_input[441]), .Z(n9341) );
  XNOR U9266 ( .A(n9357), .B(n9356), .Z(n9339) );
  XNOR U9267 ( .A(n9377), .B(n9362), .Z(n9356) );
  XOR U9268 ( .A(p_input[2056]), .B(p_input[440]), .Z(n9362) );
  XOR U9269 ( .A(n9353), .B(n9361), .Z(n9377) );
  XOR U9270 ( .A(n9378), .B(n9358), .Z(n9361) );
  XOR U9271 ( .A(p_input[2054]), .B(p_input[438]), .Z(n9358) );
  XNOR U9272 ( .A(p_input[2055]), .B(p_input[439]), .Z(n9378) );
  XNOR U9273 ( .A(n6328), .B(p_input[434]), .Z(n9353) );
  XNOR U9274 ( .A(n9367), .B(n9366), .Z(n9357) );
  XOR U9275 ( .A(n9379), .B(n9363), .Z(n9366) );
  XOR U9276 ( .A(p_input[2051]), .B(p_input[435]), .Z(n9363) );
  XNOR U9277 ( .A(p_input[2052]), .B(p_input[436]), .Z(n9379) );
  XOR U9278 ( .A(p_input[2053]), .B(p_input[437]), .Z(n9367) );
  XOR U9279 ( .A(n9380), .B(n9381), .Z(n9268) );
  AND U9280 ( .A(n115), .B(n9382), .Z(n9381) );
  XNOR U9281 ( .A(n9383), .B(n9380), .Z(n9382) );
  XNOR U9282 ( .A(n9384), .B(n9385), .Z(n115) );
  AND U9283 ( .A(n9386), .B(n9387), .Z(n9385) );
  XOR U9284 ( .A(n9281), .B(n9384), .Z(n9387) );
  AND U9285 ( .A(n9388), .B(n9389), .Z(n9281) );
  XNOR U9286 ( .A(n9278), .B(n9384), .Z(n9386) );
  XOR U9287 ( .A(n9390), .B(n9391), .Z(n9278) );
  AND U9288 ( .A(n119), .B(n9392), .Z(n9391) );
  XOR U9289 ( .A(n9393), .B(n9390), .Z(n9392) );
  XOR U9290 ( .A(n9394), .B(n9395), .Z(n9384) );
  AND U9291 ( .A(n9396), .B(n9397), .Z(n9395) );
  XNOR U9292 ( .A(n9394), .B(n9388), .Z(n9397) );
  IV U9293 ( .A(n9296), .Z(n9388) );
  XOR U9294 ( .A(n9398), .B(n9399), .Z(n9296) );
  XOR U9295 ( .A(n9400), .B(n9389), .Z(n9399) );
  AND U9296 ( .A(n9323), .B(n9401), .Z(n9389) );
  AND U9297 ( .A(n9402), .B(n9403), .Z(n9400) );
  XOR U9298 ( .A(n9404), .B(n9398), .Z(n9402) );
  XNOR U9299 ( .A(n9293), .B(n9394), .Z(n9396) );
  XOR U9300 ( .A(n9405), .B(n9406), .Z(n9293) );
  AND U9301 ( .A(n119), .B(n9407), .Z(n9406) );
  XOR U9302 ( .A(n9408), .B(n9405), .Z(n9407) );
  XOR U9303 ( .A(n9409), .B(n9410), .Z(n9394) );
  AND U9304 ( .A(n9411), .B(n9412), .Z(n9410) );
  XNOR U9305 ( .A(n9409), .B(n9323), .Z(n9412) );
  XOR U9306 ( .A(n9413), .B(n9403), .Z(n9323) );
  XNOR U9307 ( .A(n9414), .B(n9398), .Z(n9403) );
  XOR U9308 ( .A(n9415), .B(n9416), .Z(n9398) );
  AND U9309 ( .A(n9417), .B(n9418), .Z(n9416) );
  XOR U9310 ( .A(n9419), .B(n9415), .Z(n9417) );
  XNOR U9311 ( .A(n9420), .B(n9421), .Z(n9414) );
  AND U9312 ( .A(n9422), .B(n9423), .Z(n9421) );
  XOR U9313 ( .A(n9420), .B(n9424), .Z(n9422) );
  XNOR U9314 ( .A(n9404), .B(n9401), .Z(n9413) );
  AND U9315 ( .A(n9425), .B(n9426), .Z(n9401) );
  XOR U9316 ( .A(n9427), .B(n9428), .Z(n9404) );
  AND U9317 ( .A(n9429), .B(n9430), .Z(n9428) );
  XOR U9318 ( .A(n9427), .B(n9431), .Z(n9429) );
  XNOR U9319 ( .A(n9320), .B(n9409), .Z(n9411) );
  XOR U9320 ( .A(n9432), .B(n9433), .Z(n9320) );
  AND U9321 ( .A(n119), .B(n9434), .Z(n9433) );
  XNOR U9322 ( .A(n9435), .B(n9432), .Z(n9434) );
  XOR U9323 ( .A(n9436), .B(n9437), .Z(n9409) );
  AND U9324 ( .A(n9438), .B(n9439), .Z(n9437) );
  XNOR U9325 ( .A(n9436), .B(n9425), .Z(n9439) );
  IV U9326 ( .A(n9371), .Z(n9425) );
  XNOR U9327 ( .A(n9440), .B(n9418), .Z(n9371) );
  XNOR U9328 ( .A(n9441), .B(n9424), .Z(n9418) );
  XOR U9329 ( .A(n9442), .B(n9443), .Z(n9424) );
  NOR U9330 ( .A(n9444), .B(n9445), .Z(n9443) );
  XNOR U9331 ( .A(n9442), .B(n9446), .Z(n9444) );
  XNOR U9332 ( .A(n9423), .B(n9415), .Z(n9441) );
  XOR U9333 ( .A(n9447), .B(n9448), .Z(n9415) );
  AND U9334 ( .A(n9449), .B(n9450), .Z(n9448) );
  XNOR U9335 ( .A(n9447), .B(n9451), .Z(n9449) );
  XNOR U9336 ( .A(n9452), .B(n9420), .Z(n9423) );
  XOR U9337 ( .A(n9453), .B(n9454), .Z(n9420) );
  AND U9338 ( .A(n9455), .B(n9456), .Z(n9454) );
  XOR U9339 ( .A(n9453), .B(n9457), .Z(n9455) );
  XNOR U9340 ( .A(n9458), .B(n9459), .Z(n9452) );
  NOR U9341 ( .A(n9460), .B(n9461), .Z(n9459) );
  XOR U9342 ( .A(n9458), .B(n9462), .Z(n9460) );
  XNOR U9343 ( .A(n9419), .B(n9426), .Z(n9440) );
  NOR U9344 ( .A(n9383), .B(n9463), .Z(n9426) );
  XOR U9345 ( .A(n9431), .B(n9430), .Z(n9419) );
  XNOR U9346 ( .A(n9464), .B(n9427), .Z(n9430) );
  XOR U9347 ( .A(n9465), .B(n9466), .Z(n9427) );
  AND U9348 ( .A(n9467), .B(n9468), .Z(n9466) );
  XOR U9349 ( .A(n9465), .B(n9469), .Z(n9467) );
  XNOR U9350 ( .A(n9470), .B(n9471), .Z(n9464) );
  NOR U9351 ( .A(n9472), .B(n9473), .Z(n9471) );
  XNOR U9352 ( .A(n9470), .B(n9474), .Z(n9472) );
  XOR U9353 ( .A(n9475), .B(n9476), .Z(n9431) );
  NOR U9354 ( .A(n9477), .B(n9478), .Z(n9476) );
  XNOR U9355 ( .A(n9475), .B(n9479), .Z(n9477) );
  XNOR U9356 ( .A(n9368), .B(n9436), .Z(n9438) );
  XOR U9357 ( .A(n9480), .B(n9481), .Z(n9368) );
  AND U9358 ( .A(n119), .B(n9482), .Z(n9481) );
  XOR U9359 ( .A(n9483), .B(n9480), .Z(n9482) );
  AND U9360 ( .A(n9380), .B(n9383), .Z(n9436) );
  XOR U9361 ( .A(n9484), .B(n9463), .Z(n9383) );
  XNOR U9362 ( .A(p_input[2048]), .B(p_input[448]), .Z(n9463) );
  XOR U9363 ( .A(n9451), .B(n9450), .Z(n9484) );
  XNOR U9364 ( .A(n9485), .B(n9457), .Z(n9450) );
  XNOR U9365 ( .A(n9446), .B(n9445), .Z(n9457) );
  XOR U9366 ( .A(n9486), .B(n9442), .Z(n9445) );
  XNOR U9367 ( .A(n6439), .B(p_input[458]), .Z(n9442) );
  XNOR U9368 ( .A(p_input[2059]), .B(p_input[459]), .Z(n9486) );
  XOR U9369 ( .A(p_input[2060]), .B(p_input[460]), .Z(n9446) );
  XNOR U9370 ( .A(n9456), .B(n9447), .Z(n9485) );
  XNOR U9371 ( .A(n6553), .B(p_input[449]), .Z(n9447) );
  XOR U9372 ( .A(n9487), .B(n9462), .Z(n9456) );
  XNOR U9373 ( .A(p_input[2063]), .B(p_input[463]), .Z(n9462) );
  XOR U9374 ( .A(n9453), .B(n9461), .Z(n9487) );
  XOR U9375 ( .A(n9488), .B(n9458), .Z(n9461) );
  XOR U9376 ( .A(p_input[2061]), .B(p_input[461]), .Z(n9458) );
  XNOR U9377 ( .A(p_input[2062]), .B(p_input[462]), .Z(n9488) );
  XNOR U9378 ( .A(n6325), .B(p_input[457]), .Z(n9453) );
  XNOR U9379 ( .A(n9469), .B(n9468), .Z(n9451) );
  XNOR U9380 ( .A(n9489), .B(n9474), .Z(n9468) );
  XOR U9381 ( .A(p_input[2056]), .B(p_input[456]), .Z(n9474) );
  XOR U9382 ( .A(n9465), .B(n9473), .Z(n9489) );
  XOR U9383 ( .A(n9490), .B(n9470), .Z(n9473) );
  XOR U9384 ( .A(p_input[2054]), .B(p_input[454]), .Z(n9470) );
  XNOR U9385 ( .A(p_input[2055]), .B(p_input[455]), .Z(n9490) );
  XNOR U9386 ( .A(n6328), .B(p_input[450]), .Z(n9465) );
  XNOR U9387 ( .A(n9479), .B(n9478), .Z(n9469) );
  XOR U9388 ( .A(n9491), .B(n9475), .Z(n9478) );
  XOR U9389 ( .A(p_input[2051]), .B(p_input[451]), .Z(n9475) );
  XNOR U9390 ( .A(p_input[2052]), .B(p_input[452]), .Z(n9491) );
  XOR U9391 ( .A(p_input[2053]), .B(p_input[453]), .Z(n9479) );
  XOR U9392 ( .A(n9492), .B(n9493), .Z(n9380) );
  AND U9393 ( .A(n119), .B(n9494), .Z(n9493) );
  XNOR U9394 ( .A(n9495), .B(n9492), .Z(n9494) );
  XNOR U9395 ( .A(n9496), .B(n9497), .Z(n119) );
  AND U9396 ( .A(n9498), .B(n9499), .Z(n9497) );
  XOR U9397 ( .A(n9393), .B(n9496), .Z(n9499) );
  AND U9398 ( .A(n9500), .B(n9501), .Z(n9393) );
  XNOR U9399 ( .A(n9390), .B(n9496), .Z(n9498) );
  XOR U9400 ( .A(n9502), .B(n9503), .Z(n9390) );
  AND U9401 ( .A(n123), .B(n9504), .Z(n9503) );
  XOR U9402 ( .A(n9505), .B(n9502), .Z(n9504) );
  XOR U9403 ( .A(n9506), .B(n9507), .Z(n9496) );
  AND U9404 ( .A(n9508), .B(n9509), .Z(n9507) );
  XNOR U9405 ( .A(n9506), .B(n9500), .Z(n9509) );
  IV U9406 ( .A(n9408), .Z(n9500) );
  XOR U9407 ( .A(n9510), .B(n9511), .Z(n9408) );
  XOR U9408 ( .A(n9512), .B(n9501), .Z(n9511) );
  AND U9409 ( .A(n9435), .B(n9513), .Z(n9501) );
  AND U9410 ( .A(n9514), .B(n9515), .Z(n9512) );
  XOR U9411 ( .A(n9516), .B(n9510), .Z(n9514) );
  XNOR U9412 ( .A(n9405), .B(n9506), .Z(n9508) );
  XOR U9413 ( .A(n9517), .B(n9518), .Z(n9405) );
  AND U9414 ( .A(n123), .B(n9519), .Z(n9518) );
  XOR U9415 ( .A(n9520), .B(n9517), .Z(n9519) );
  XOR U9416 ( .A(n9521), .B(n9522), .Z(n9506) );
  AND U9417 ( .A(n9523), .B(n9524), .Z(n9522) );
  XNOR U9418 ( .A(n9521), .B(n9435), .Z(n9524) );
  XOR U9419 ( .A(n9525), .B(n9515), .Z(n9435) );
  XNOR U9420 ( .A(n9526), .B(n9510), .Z(n9515) );
  XOR U9421 ( .A(n9527), .B(n9528), .Z(n9510) );
  AND U9422 ( .A(n9529), .B(n9530), .Z(n9528) );
  XOR U9423 ( .A(n9531), .B(n9527), .Z(n9529) );
  XNOR U9424 ( .A(n9532), .B(n9533), .Z(n9526) );
  AND U9425 ( .A(n9534), .B(n9535), .Z(n9533) );
  XOR U9426 ( .A(n9532), .B(n9536), .Z(n9534) );
  XNOR U9427 ( .A(n9516), .B(n9513), .Z(n9525) );
  AND U9428 ( .A(n9537), .B(n9538), .Z(n9513) );
  XOR U9429 ( .A(n9539), .B(n9540), .Z(n9516) );
  AND U9430 ( .A(n9541), .B(n9542), .Z(n9540) );
  XOR U9431 ( .A(n9539), .B(n9543), .Z(n9541) );
  XNOR U9432 ( .A(n9432), .B(n9521), .Z(n9523) );
  XOR U9433 ( .A(n9544), .B(n9545), .Z(n9432) );
  AND U9434 ( .A(n123), .B(n9546), .Z(n9545) );
  XNOR U9435 ( .A(n9547), .B(n9544), .Z(n9546) );
  XOR U9436 ( .A(n9548), .B(n9549), .Z(n9521) );
  AND U9437 ( .A(n9550), .B(n9551), .Z(n9549) );
  XNOR U9438 ( .A(n9548), .B(n9537), .Z(n9551) );
  IV U9439 ( .A(n9483), .Z(n9537) );
  XNOR U9440 ( .A(n9552), .B(n9530), .Z(n9483) );
  XNOR U9441 ( .A(n9553), .B(n9536), .Z(n9530) );
  XOR U9442 ( .A(n9554), .B(n9555), .Z(n9536) );
  NOR U9443 ( .A(n9556), .B(n9557), .Z(n9555) );
  XNOR U9444 ( .A(n9554), .B(n9558), .Z(n9556) );
  XNOR U9445 ( .A(n9535), .B(n9527), .Z(n9553) );
  XOR U9446 ( .A(n9559), .B(n9560), .Z(n9527) );
  AND U9447 ( .A(n9561), .B(n9562), .Z(n9560) );
  XNOR U9448 ( .A(n9559), .B(n9563), .Z(n9561) );
  XNOR U9449 ( .A(n9564), .B(n9532), .Z(n9535) );
  XOR U9450 ( .A(n9565), .B(n9566), .Z(n9532) );
  AND U9451 ( .A(n9567), .B(n9568), .Z(n9566) );
  XOR U9452 ( .A(n9565), .B(n9569), .Z(n9567) );
  XNOR U9453 ( .A(n9570), .B(n9571), .Z(n9564) );
  NOR U9454 ( .A(n9572), .B(n9573), .Z(n9571) );
  XOR U9455 ( .A(n9570), .B(n9574), .Z(n9572) );
  XNOR U9456 ( .A(n9531), .B(n9538), .Z(n9552) );
  NOR U9457 ( .A(n9495), .B(n9575), .Z(n9538) );
  XOR U9458 ( .A(n9543), .B(n9542), .Z(n9531) );
  XNOR U9459 ( .A(n9576), .B(n9539), .Z(n9542) );
  XOR U9460 ( .A(n9577), .B(n9578), .Z(n9539) );
  AND U9461 ( .A(n9579), .B(n9580), .Z(n9578) );
  XOR U9462 ( .A(n9577), .B(n9581), .Z(n9579) );
  XNOR U9463 ( .A(n9582), .B(n9583), .Z(n9576) );
  NOR U9464 ( .A(n9584), .B(n9585), .Z(n9583) );
  XNOR U9465 ( .A(n9582), .B(n9586), .Z(n9584) );
  XOR U9466 ( .A(n9587), .B(n9588), .Z(n9543) );
  NOR U9467 ( .A(n9589), .B(n9590), .Z(n9588) );
  XNOR U9468 ( .A(n9587), .B(n9591), .Z(n9589) );
  XNOR U9469 ( .A(n9480), .B(n9548), .Z(n9550) );
  XOR U9470 ( .A(n9592), .B(n9593), .Z(n9480) );
  AND U9471 ( .A(n123), .B(n9594), .Z(n9593) );
  XOR U9472 ( .A(n9595), .B(n9592), .Z(n9594) );
  AND U9473 ( .A(n9492), .B(n9495), .Z(n9548) );
  XOR U9474 ( .A(n9596), .B(n9575), .Z(n9495) );
  XNOR U9475 ( .A(p_input[2048]), .B(p_input[464]), .Z(n9575) );
  XOR U9476 ( .A(n9563), .B(n9562), .Z(n9596) );
  XNOR U9477 ( .A(n9597), .B(n9569), .Z(n9562) );
  XNOR U9478 ( .A(n9558), .B(n9557), .Z(n9569) );
  XOR U9479 ( .A(n9598), .B(n9554), .Z(n9557) );
  XNOR U9480 ( .A(n6439), .B(p_input[474]), .Z(n9554) );
  XNOR U9481 ( .A(p_input[2059]), .B(p_input[475]), .Z(n9598) );
  XOR U9482 ( .A(p_input[2060]), .B(p_input[476]), .Z(n9558) );
  XNOR U9483 ( .A(n9568), .B(n9559), .Z(n9597) );
  XNOR U9484 ( .A(n6553), .B(p_input[465]), .Z(n9559) );
  XOR U9485 ( .A(n9599), .B(n9574), .Z(n9568) );
  XNOR U9486 ( .A(p_input[2063]), .B(p_input[479]), .Z(n9574) );
  XOR U9487 ( .A(n9565), .B(n9573), .Z(n9599) );
  XOR U9488 ( .A(n9600), .B(n9570), .Z(n9573) );
  XOR U9489 ( .A(p_input[2061]), .B(p_input[477]), .Z(n9570) );
  XNOR U9490 ( .A(p_input[2062]), .B(p_input[478]), .Z(n9600) );
  XNOR U9491 ( .A(n6325), .B(p_input[473]), .Z(n9565) );
  XNOR U9492 ( .A(n9581), .B(n9580), .Z(n9563) );
  XNOR U9493 ( .A(n9601), .B(n9586), .Z(n9580) );
  XOR U9494 ( .A(p_input[2056]), .B(p_input[472]), .Z(n9586) );
  XOR U9495 ( .A(n9577), .B(n9585), .Z(n9601) );
  XOR U9496 ( .A(n9602), .B(n9582), .Z(n9585) );
  XOR U9497 ( .A(p_input[2054]), .B(p_input[470]), .Z(n9582) );
  XNOR U9498 ( .A(p_input[2055]), .B(p_input[471]), .Z(n9602) );
  XNOR U9499 ( .A(n6328), .B(p_input[466]), .Z(n9577) );
  XNOR U9500 ( .A(n9591), .B(n9590), .Z(n9581) );
  XOR U9501 ( .A(n9603), .B(n9587), .Z(n9590) );
  XOR U9502 ( .A(p_input[2051]), .B(p_input[467]), .Z(n9587) );
  XNOR U9503 ( .A(p_input[2052]), .B(p_input[468]), .Z(n9603) );
  XOR U9504 ( .A(p_input[2053]), .B(p_input[469]), .Z(n9591) );
  XOR U9505 ( .A(n9604), .B(n9605), .Z(n9492) );
  AND U9506 ( .A(n123), .B(n9606), .Z(n9605) );
  XNOR U9507 ( .A(n9607), .B(n9604), .Z(n9606) );
  XNOR U9508 ( .A(n9608), .B(n9609), .Z(n123) );
  AND U9509 ( .A(n9610), .B(n9611), .Z(n9609) );
  XOR U9510 ( .A(n9505), .B(n9608), .Z(n9611) );
  AND U9511 ( .A(n9612), .B(n9613), .Z(n9505) );
  XNOR U9512 ( .A(n9502), .B(n9608), .Z(n9610) );
  XOR U9513 ( .A(n9614), .B(n9615), .Z(n9502) );
  AND U9514 ( .A(n127), .B(n9616), .Z(n9615) );
  XOR U9515 ( .A(n9617), .B(n9614), .Z(n9616) );
  XOR U9516 ( .A(n9618), .B(n9619), .Z(n9608) );
  AND U9517 ( .A(n9620), .B(n9621), .Z(n9619) );
  XNOR U9518 ( .A(n9618), .B(n9612), .Z(n9621) );
  IV U9519 ( .A(n9520), .Z(n9612) );
  XOR U9520 ( .A(n9622), .B(n9623), .Z(n9520) );
  XOR U9521 ( .A(n9624), .B(n9613), .Z(n9623) );
  AND U9522 ( .A(n9547), .B(n9625), .Z(n9613) );
  AND U9523 ( .A(n9626), .B(n9627), .Z(n9624) );
  XOR U9524 ( .A(n9628), .B(n9622), .Z(n9626) );
  XNOR U9525 ( .A(n9517), .B(n9618), .Z(n9620) );
  XOR U9526 ( .A(n9629), .B(n9630), .Z(n9517) );
  AND U9527 ( .A(n127), .B(n9631), .Z(n9630) );
  XOR U9528 ( .A(n9632), .B(n9629), .Z(n9631) );
  XOR U9529 ( .A(n9633), .B(n9634), .Z(n9618) );
  AND U9530 ( .A(n9635), .B(n9636), .Z(n9634) );
  XNOR U9531 ( .A(n9633), .B(n9547), .Z(n9636) );
  XOR U9532 ( .A(n9637), .B(n9627), .Z(n9547) );
  XNOR U9533 ( .A(n9638), .B(n9622), .Z(n9627) );
  XOR U9534 ( .A(n9639), .B(n9640), .Z(n9622) );
  AND U9535 ( .A(n9641), .B(n9642), .Z(n9640) );
  XOR U9536 ( .A(n9643), .B(n9639), .Z(n9641) );
  XNOR U9537 ( .A(n9644), .B(n9645), .Z(n9638) );
  AND U9538 ( .A(n9646), .B(n9647), .Z(n9645) );
  XOR U9539 ( .A(n9644), .B(n9648), .Z(n9646) );
  XNOR U9540 ( .A(n9628), .B(n9625), .Z(n9637) );
  AND U9541 ( .A(n9649), .B(n9650), .Z(n9625) );
  XOR U9542 ( .A(n9651), .B(n9652), .Z(n9628) );
  AND U9543 ( .A(n9653), .B(n9654), .Z(n9652) );
  XOR U9544 ( .A(n9651), .B(n9655), .Z(n9653) );
  XNOR U9545 ( .A(n9544), .B(n9633), .Z(n9635) );
  XOR U9546 ( .A(n9656), .B(n9657), .Z(n9544) );
  AND U9547 ( .A(n127), .B(n9658), .Z(n9657) );
  XNOR U9548 ( .A(n9659), .B(n9656), .Z(n9658) );
  XOR U9549 ( .A(n9660), .B(n9661), .Z(n9633) );
  AND U9550 ( .A(n9662), .B(n9663), .Z(n9661) );
  XNOR U9551 ( .A(n9660), .B(n9649), .Z(n9663) );
  IV U9552 ( .A(n9595), .Z(n9649) );
  XNOR U9553 ( .A(n9664), .B(n9642), .Z(n9595) );
  XNOR U9554 ( .A(n9665), .B(n9648), .Z(n9642) );
  XOR U9555 ( .A(n9666), .B(n9667), .Z(n9648) );
  NOR U9556 ( .A(n9668), .B(n9669), .Z(n9667) );
  XNOR U9557 ( .A(n9666), .B(n9670), .Z(n9668) );
  XNOR U9558 ( .A(n9647), .B(n9639), .Z(n9665) );
  XOR U9559 ( .A(n9671), .B(n9672), .Z(n9639) );
  AND U9560 ( .A(n9673), .B(n9674), .Z(n9672) );
  XNOR U9561 ( .A(n9671), .B(n9675), .Z(n9673) );
  XNOR U9562 ( .A(n9676), .B(n9644), .Z(n9647) );
  XOR U9563 ( .A(n9677), .B(n9678), .Z(n9644) );
  AND U9564 ( .A(n9679), .B(n9680), .Z(n9678) );
  XOR U9565 ( .A(n9677), .B(n9681), .Z(n9679) );
  XNOR U9566 ( .A(n9682), .B(n9683), .Z(n9676) );
  NOR U9567 ( .A(n9684), .B(n9685), .Z(n9683) );
  XOR U9568 ( .A(n9682), .B(n9686), .Z(n9684) );
  XNOR U9569 ( .A(n9643), .B(n9650), .Z(n9664) );
  NOR U9570 ( .A(n9607), .B(n9687), .Z(n9650) );
  XOR U9571 ( .A(n9655), .B(n9654), .Z(n9643) );
  XNOR U9572 ( .A(n9688), .B(n9651), .Z(n9654) );
  XOR U9573 ( .A(n9689), .B(n9690), .Z(n9651) );
  AND U9574 ( .A(n9691), .B(n9692), .Z(n9690) );
  XOR U9575 ( .A(n9689), .B(n9693), .Z(n9691) );
  XNOR U9576 ( .A(n9694), .B(n9695), .Z(n9688) );
  NOR U9577 ( .A(n9696), .B(n9697), .Z(n9695) );
  XNOR U9578 ( .A(n9694), .B(n9698), .Z(n9696) );
  XOR U9579 ( .A(n9699), .B(n9700), .Z(n9655) );
  NOR U9580 ( .A(n9701), .B(n9702), .Z(n9700) );
  XNOR U9581 ( .A(n9699), .B(n9703), .Z(n9701) );
  XNOR U9582 ( .A(n9592), .B(n9660), .Z(n9662) );
  XOR U9583 ( .A(n9704), .B(n9705), .Z(n9592) );
  AND U9584 ( .A(n127), .B(n9706), .Z(n9705) );
  XOR U9585 ( .A(n9707), .B(n9704), .Z(n9706) );
  AND U9586 ( .A(n9604), .B(n9607), .Z(n9660) );
  XOR U9587 ( .A(n9708), .B(n9687), .Z(n9607) );
  XNOR U9588 ( .A(p_input[2048]), .B(p_input[480]), .Z(n9687) );
  XOR U9589 ( .A(n9675), .B(n9674), .Z(n9708) );
  XNOR U9590 ( .A(n9709), .B(n9681), .Z(n9674) );
  XNOR U9591 ( .A(n9670), .B(n9669), .Z(n9681) );
  XOR U9592 ( .A(n9710), .B(n9666), .Z(n9669) );
  XNOR U9593 ( .A(n6439), .B(p_input[490]), .Z(n9666) );
  XNOR U9594 ( .A(p_input[2059]), .B(p_input[491]), .Z(n9710) );
  XOR U9595 ( .A(p_input[2060]), .B(p_input[492]), .Z(n9670) );
  XNOR U9596 ( .A(n9680), .B(n9671), .Z(n9709) );
  XNOR U9597 ( .A(n6553), .B(p_input[481]), .Z(n9671) );
  XOR U9598 ( .A(n9711), .B(n9686), .Z(n9680) );
  XNOR U9599 ( .A(p_input[2063]), .B(p_input[495]), .Z(n9686) );
  XOR U9600 ( .A(n9677), .B(n9685), .Z(n9711) );
  XOR U9601 ( .A(n9712), .B(n9682), .Z(n9685) );
  XOR U9602 ( .A(p_input[2061]), .B(p_input[493]), .Z(n9682) );
  XNOR U9603 ( .A(p_input[2062]), .B(p_input[494]), .Z(n9712) );
  XNOR U9604 ( .A(n6325), .B(p_input[489]), .Z(n9677) );
  XNOR U9605 ( .A(n9693), .B(n9692), .Z(n9675) );
  XNOR U9606 ( .A(n9713), .B(n9698), .Z(n9692) );
  XOR U9607 ( .A(p_input[2056]), .B(p_input[488]), .Z(n9698) );
  XOR U9608 ( .A(n9689), .B(n9697), .Z(n9713) );
  XOR U9609 ( .A(n9714), .B(n9694), .Z(n9697) );
  XOR U9610 ( .A(p_input[2054]), .B(p_input[486]), .Z(n9694) );
  XNOR U9611 ( .A(p_input[2055]), .B(p_input[487]), .Z(n9714) );
  XNOR U9612 ( .A(n6328), .B(p_input[482]), .Z(n9689) );
  XNOR U9613 ( .A(n9703), .B(n9702), .Z(n9693) );
  XOR U9614 ( .A(n9715), .B(n9699), .Z(n9702) );
  XOR U9615 ( .A(p_input[2051]), .B(p_input[483]), .Z(n9699) );
  XNOR U9616 ( .A(p_input[2052]), .B(p_input[484]), .Z(n9715) );
  XOR U9617 ( .A(p_input[2053]), .B(p_input[485]), .Z(n9703) );
  XOR U9618 ( .A(n9716), .B(n9717), .Z(n9604) );
  AND U9619 ( .A(n127), .B(n9718), .Z(n9717) );
  XNOR U9620 ( .A(n9719), .B(n9716), .Z(n9718) );
  XNOR U9621 ( .A(n9720), .B(n9721), .Z(n127) );
  AND U9622 ( .A(n9722), .B(n9723), .Z(n9721) );
  XOR U9623 ( .A(n9617), .B(n9720), .Z(n9723) );
  AND U9624 ( .A(n9724), .B(n9725), .Z(n9617) );
  XNOR U9625 ( .A(n9614), .B(n9720), .Z(n9722) );
  XOR U9626 ( .A(n9726), .B(n9727), .Z(n9614) );
  AND U9627 ( .A(n131), .B(n9728), .Z(n9727) );
  XOR U9628 ( .A(n9729), .B(n9726), .Z(n9728) );
  XOR U9629 ( .A(n9730), .B(n9731), .Z(n9720) );
  AND U9630 ( .A(n9732), .B(n9733), .Z(n9731) );
  XNOR U9631 ( .A(n9730), .B(n9724), .Z(n9733) );
  IV U9632 ( .A(n9632), .Z(n9724) );
  XOR U9633 ( .A(n9734), .B(n9735), .Z(n9632) );
  XOR U9634 ( .A(n9736), .B(n9725), .Z(n9735) );
  AND U9635 ( .A(n9659), .B(n9737), .Z(n9725) );
  AND U9636 ( .A(n9738), .B(n9739), .Z(n9736) );
  XOR U9637 ( .A(n9740), .B(n9734), .Z(n9738) );
  XNOR U9638 ( .A(n9629), .B(n9730), .Z(n9732) );
  XOR U9639 ( .A(n9741), .B(n9742), .Z(n9629) );
  AND U9640 ( .A(n131), .B(n9743), .Z(n9742) );
  XOR U9641 ( .A(n9744), .B(n9741), .Z(n9743) );
  XOR U9642 ( .A(n9745), .B(n9746), .Z(n9730) );
  AND U9643 ( .A(n9747), .B(n9748), .Z(n9746) );
  XNOR U9644 ( .A(n9745), .B(n9659), .Z(n9748) );
  XOR U9645 ( .A(n9749), .B(n9739), .Z(n9659) );
  XNOR U9646 ( .A(n9750), .B(n9734), .Z(n9739) );
  XOR U9647 ( .A(n9751), .B(n9752), .Z(n9734) );
  AND U9648 ( .A(n9753), .B(n9754), .Z(n9752) );
  XOR U9649 ( .A(n9755), .B(n9751), .Z(n9753) );
  XNOR U9650 ( .A(n9756), .B(n9757), .Z(n9750) );
  AND U9651 ( .A(n9758), .B(n9759), .Z(n9757) );
  XOR U9652 ( .A(n9756), .B(n9760), .Z(n9758) );
  XNOR U9653 ( .A(n9740), .B(n9737), .Z(n9749) );
  AND U9654 ( .A(n9761), .B(n9762), .Z(n9737) );
  XOR U9655 ( .A(n9763), .B(n9764), .Z(n9740) );
  AND U9656 ( .A(n9765), .B(n9766), .Z(n9764) );
  XOR U9657 ( .A(n9763), .B(n9767), .Z(n9765) );
  XNOR U9658 ( .A(n9656), .B(n9745), .Z(n9747) );
  XOR U9659 ( .A(n9768), .B(n9769), .Z(n9656) );
  AND U9660 ( .A(n131), .B(n9770), .Z(n9769) );
  XNOR U9661 ( .A(n9771), .B(n9768), .Z(n9770) );
  XOR U9662 ( .A(n9772), .B(n9773), .Z(n9745) );
  AND U9663 ( .A(n9774), .B(n9775), .Z(n9773) );
  XNOR U9664 ( .A(n9772), .B(n9761), .Z(n9775) );
  IV U9665 ( .A(n9707), .Z(n9761) );
  XNOR U9666 ( .A(n9776), .B(n9754), .Z(n9707) );
  XNOR U9667 ( .A(n9777), .B(n9760), .Z(n9754) );
  XOR U9668 ( .A(n9778), .B(n9779), .Z(n9760) );
  NOR U9669 ( .A(n9780), .B(n9781), .Z(n9779) );
  XNOR U9670 ( .A(n9778), .B(n9782), .Z(n9780) );
  XNOR U9671 ( .A(n9759), .B(n9751), .Z(n9777) );
  XOR U9672 ( .A(n9783), .B(n9784), .Z(n9751) );
  AND U9673 ( .A(n9785), .B(n9786), .Z(n9784) );
  XNOR U9674 ( .A(n9783), .B(n9787), .Z(n9785) );
  XNOR U9675 ( .A(n9788), .B(n9756), .Z(n9759) );
  XOR U9676 ( .A(n9789), .B(n9790), .Z(n9756) );
  AND U9677 ( .A(n9791), .B(n9792), .Z(n9790) );
  XOR U9678 ( .A(n9789), .B(n9793), .Z(n9791) );
  XNOR U9679 ( .A(n9794), .B(n9795), .Z(n9788) );
  NOR U9680 ( .A(n9796), .B(n9797), .Z(n9795) );
  XOR U9681 ( .A(n9794), .B(n9798), .Z(n9796) );
  XNOR U9682 ( .A(n9755), .B(n9762), .Z(n9776) );
  NOR U9683 ( .A(n9719), .B(n9799), .Z(n9762) );
  XOR U9684 ( .A(n9767), .B(n9766), .Z(n9755) );
  XNOR U9685 ( .A(n9800), .B(n9763), .Z(n9766) );
  XOR U9686 ( .A(n9801), .B(n9802), .Z(n9763) );
  AND U9687 ( .A(n9803), .B(n9804), .Z(n9802) );
  XOR U9688 ( .A(n9801), .B(n9805), .Z(n9803) );
  XNOR U9689 ( .A(n9806), .B(n9807), .Z(n9800) );
  NOR U9690 ( .A(n9808), .B(n9809), .Z(n9807) );
  XNOR U9691 ( .A(n9806), .B(n9810), .Z(n9808) );
  XOR U9692 ( .A(n9811), .B(n9812), .Z(n9767) );
  NOR U9693 ( .A(n9813), .B(n9814), .Z(n9812) );
  XNOR U9694 ( .A(n9811), .B(n9815), .Z(n9813) );
  XNOR U9695 ( .A(n9704), .B(n9772), .Z(n9774) );
  XOR U9696 ( .A(n9816), .B(n9817), .Z(n9704) );
  AND U9697 ( .A(n131), .B(n9818), .Z(n9817) );
  XOR U9698 ( .A(n9819), .B(n9816), .Z(n9818) );
  AND U9699 ( .A(n9716), .B(n9719), .Z(n9772) );
  XOR U9700 ( .A(n9820), .B(n9799), .Z(n9719) );
  XNOR U9701 ( .A(p_input[2048]), .B(p_input[496]), .Z(n9799) );
  XOR U9702 ( .A(n9787), .B(n9786), .Z(n9820) );
  XNOR U9703 ( .A(n9821), .B(n9793), .Z(n9786) );
  XNOR U9704 ( .A(n9782), .B(n9781), .Z(n9793) );
  XOR U9705 ( .A(n9822), .B(n9778), .Z(n9781) );
  XNOR U9706 ( .A(n6439), .B(p_input[506]), .Z(n9778) );
  XNOR U9707 ( .A(p_input[2059]), .B(p_input[507]), .Z(n9822) );
  XOR U9708 ( .A(p_input[2060]), .B(p_input[508]), .Z(n9782) );
  XNOR U9709 ( .A(n9792), .B(n9783), .Z(n9821) );
  XNOR U9710 ( .A(n6553), .B(p_input[497]), .Z(n9783) );
  XOR U9711 ( .A(n9823), .B(n9798), .Z(n9792) );
  XNOR U9712 ( .A(p_input[2063]), .B(p_input[511]), .Z(n9798) );
  XOR U9713 ( .A(n9789), .B(n9797), .Z(n9823) );
  XOR U9714 ( .A(n9824), .B(n9794), .Z(n9797) );
  XOR U9715 ( .A(p_input[2061]), .B(p_input[509]), .Z(n9794) );
  XNOR U9716 ( .A(p_input[2062]), .B(p_input[510]), .Z(n9824) );
  XNOR U9717 ( .A(n6325), .B(p_input[505]), .Z(n9789) );
  XNOR U9718 ( .A(n9805), .B(n9804), .Z(n9787) );
  XNOR U9719 ( .A(n9825), .B(n9810), .Z(n9804) );
  XOR U9720 ( .A(p_input[2056]), .B(p_input[504]), .Z(n9810) );
  XOR U9721 ( .A(n9801), .B(n9809), .Z(n9825) );
  XOR U9722 ( .A(n9826), .B(n9806), .Z(n9809) );
  XOR U9723 ( .A(p_input[2054]), .B(p_input[502]), .Z(n9806) );
  XNOR U9724 ( .A(p_input[2055]), .B(p_input[503]), .Z(n9826) );
  XNOR U9725 ( .A(n6328), .B(p_input[498]), .Z(n9801) );
  XNOR U9726 ( .A(n9815), .B(n9814), .Z(n9805) );
  XOR U9727 ( .A(n9827), .B(n9811), .Z(n9814) );
  XOR U9728 ( .A(p_input[2051]), .B(p_input[499]), .Z(n9811) );
  XNOR U9729 ( .A(p_input[2052]), .B(p_input[500]), .Z(n9827) );
  XOR U9730 ( .A(p_input[2053]), .B(p_input[501]), .Z(n9815) );
  XOR U9731 ( .A(n9828), .B(n9829), .Z(n9716) );
  AND U9732 ( .A(n131), .B(n9830), .Z(n9829) );
  XNOR U9733 ( .A(n9831), .B(n9828), .Z(n9830) );
  XNOR U9734 ( .A(n9832), .B(n9833), .Z(n131) );
  AND U9735 ( .A(n9834), .B(n9835), .Z(n9833) );
  XOR U9736 ( .A(n9729), .B(n9832), .Z(n9835) );
  AND U9737 ( .A(n9836), .B(n9837), .Z(n9729) );
  XNOR U9738 ( .A(n9726), .B(n9832), .Z(n9834) );
  XOR U9739 ( .A(n9838), .B(n9839), .Z(n9726) );
  AND U9740 ( .A(n135), .B(n9840), .Z(n9839) );
  XOR U9741 ( .A(n9841), .B(n9838), .Z(n9840) );
  XOR U9742 ( .A(n9842), .B(n9843), .Z(n9832) );
  AND U9743 ( .A(n9844), .B(n9845), .Z(n9843) );
  XNOR U9744 ( .A(n9842), .B(n9836), .Z(n9845) );
  IV U9745 ( .A(n9744), .Z(n9836) );
  XOR U9746 ( .A(n9846), .B(n9847), .Z(n9744) );
  XOR U9747 ( .A(n9848), .B(n9837), .Z(n9847) );
  AND U9748 ( .A(n9771), .B(n9849), .Z(n9837) );
  AND U9749 ( .A(n9850), .B(n9851), .Z(n9848) );
  XOR U9750 ( .A(n9852), .B(n9846), .Z(n9850) );
  XNOR U9751 ( .A(n9741), .B(n9842), .Z(n9844) );
  XOR U9752 ( .A(n9853), .B(n9854), .Z(n9741) );
  AND U9753 ( .A(n135), .B(n9855), .Z(n9854) );
  XOR U9754 ( .A(n9856), .B(n9853), .Z(n9855) );
  XOR U9755 ( .A(n9857), .B(n9858), .Z(n9842) );
  AND U9756 ( .A(n9859), .B(n9860), .Z(n9858) );
  XNOR U9757 ( .A(n9857), .B(n9771), .Z(n9860) );
  XOR U9758 ( .A(n9861), .B(n9851), .Z(n9771) );
  XNOR U9759 ( .A(n9862), .B(n9846), .Z(n9851) );
  XOR U9760 ( .A(n9863), .B(n9864), .Z(n9846) );
  AND U9761 ( .A(n9865), .B(n9866), .Z(n9864) );
  XOR U9762 ( .A(n9867), .B(n9863), .Z(n9865) );
  XNOR U9763 ( .A(n9868), .B(n9869), .Z(n9862) );
  AND U9764 ( .A(n9870), .B(n9871), .Z(n9869) );
  XOR U9765 ( .A(n9868), .B(n9872), .Z(n9870) );
  XNOR U9766 ( .A(n9852), .B(n9849), .Z(n9861) );
  AND U9767 ( .A(n9873), .B(n9874), .Z(n9849) );
  XOR U9768 ( .A(n9875), .B(n9876), .Z(n9852) );
  AND U9769 ( .A(n9877), .B(n9878), .Z(n9876) );
  XOR U9770 ( .A(n9875), .B(n9879), .Z(n9877) );
  XNOR U9771 ( .A(n9768), .B(n9857), .Z(n9859) );
  XOR U9772 ( .A(n9880), .B(n9881), .Z(n9768) );
  AND U9773 ( .A(n135), .B(n9882), .Z(n9881) );
  XNOR U9774 ( .A(n9883), .B(n9880), .Z(n9882) );
  XOR U9775 ( .A(n9884), .B(n9885), .Z(n9857) );
  AND U9776 ( .A(n9886), .B(n9887), .Z(n9885) );
  XNOR U9777 ( .A(n9884), .B(n9873), .Z(n9887) );
  IV U9778 ( .A(n9819), .Z(n9873) );
  XNOR U9779 ( .A(n9888), .B(n9866), .Z(n9819) );
  XNOR U9780 ( .A(n9889), .B(n9872), .Z(n9866) );
  XOR U9781 ( .A(n9890), .B(n9891), .Z(n9872) );
  NOR U9782 ( .A(n9892), .B(n9893), .Z(n9891) );
  XNOR U9783 ( .A(n9890), .B(n9894), .Z(n9892) );
  XNOR U9784 ( .A(n9871), .B(n9863), .Z(n9889) );
  XOR U9785 ( .A(n9895), .B(n9896), .Z(n9863) );
  AND U9786 ( .A(n9897), .B(n9898), .Z(n9896) );
  XNOR U9787 ( .A(n9895), .B(n9899), .Z(n9897) );
  XNOR U9788 ( .A(n9900), .B(n9868), .Z(n9871) );
  XOR U9789 ( .A(n9901), .B(n9902), .Z(n9868) );
  AND U9790 ( .A(n9903), .B(n9904), .Z(n9902) );
  XOR U9791 ( .A(n9901), .B(n9905), .Z(n9903) );
  XNOR U9792 ( .A(n9906), .B(n9907), .Z(n9900) );
  NOR U9793 ( .A(n9908), .B(n9909), .Z(n9907) );
  XOR U9794 ( .A(n9906), .B(n9910), .Z(n9908) );
  XNOR U9795 ( .A(n9867), .B(n9874), .Z(n9888) );
  NOR U9796 ( .A(n9831), .B(n9911), .Z(n9874) );
  XOR U9797 ( .A(n9879), .B(n9878), .Z(n9867) );
  XNOR U9798 ( .A(n9912), .B(n9875), .Z(n9878) );
  XOR U9799 ( .A(n9913), .B(n9914), .Z(n9875) );
  AND U9800 ( .A(n9915), .B(n9916), .Z(n9914) );
  XOR U9801 ( .A(n9913), .B(n9917), .Z(n9915) );
  XNOR U9802 ( .A(n9918), .B(n9919), .Z(n9912) );
  NOR U9803 ( .A(n9920), .B(n9921), .Z(n9919) );
  XNOR U9804 ( .A(n9918), .B(n9922), .Z(n9920) );
  XOR U9805 ( .A(n9923), .B(n9924), .Z(n9879) );
  NOR U9806 ( .A(n9925), .B(n9926), .Z(n9924) );
  XNOR U9807 ( .A(n9923), .B(n9927), .Z(n9925) );
  XNOR U9808 ( .A(n9816), .B(n9884), .Z(n9886) );
  XOR U9809 ( .A(n9928), .B(n9929), .Z(n9816) );
  AND U9810 ( .A(n135), .B(n9930), .Z(n9929) );
  XOR U9811 ( .A(n9931), .B(n9928), .Z(n9930) );
  AND U9812 ( .A(n9828), .B(n9831), .Z(n9884) );
  XOR U9813 ( .A(n9932), .B(n9911), .Z(n9831) );
  XNOR U9814 ( .A(p_input[2048]), .B(p_input[512]), .Z(n9911) );
  XOR U9815 ( .A(n9899), .B(n9898), .Z(n9932) );
  XNOR U9816 ( .A(n9933), .B(n9905), .Z(n9898) );
  XNOR U9817 ( .A(n9894), .B(n9893), .Z(n9905) );
  XOR U9818 ( .A(n9934), .B(n9890), .Z(n9893) );
  XNOR U9819 ( .A(n6439), .B(p_input[522]), .Z(n9890) );
  XNOR U9820 ( .A(p_input[2059]), .B(p_input[523]), .Z(n9934) );
  XOR U9821 ( .A(p_input[2060]), .B(p_input[524]), .Z(n9894) );
  XNOR U9822 ( .A(n9904), .B(n9895), .Z(n9933) );
  XNOR U9823 ( .A(n6553), .B(p_input[513]), .Z(n9895) );
  XOR U9824 ( .A(n9935), .B(n9910), .Z(n9904) );
  XNOR U9825 ( .A(p_input[2063]), .B(p_input[527]), .Z(n9910) );
  XOR U9826 ( .A(n9901), .B(n9909), .Z(n9935) );
  XOR U9827 ( .A(n9936), .B(n9906), .Z(n9909) );
  XOR U9828 ( .A(p_input[2061]), .B(p_input[525]), .Z(n9906) );
  XNOR U9829 ( .A(p_input[2062]), .B(p_input[526]), .Z(n9936) );
  XNOR U9830 ( .A(n6325), .B(p_input[521]), .Z(n9901) );
  XNOR U9831 ( .A(n9917), .B(n9916), .Z(n9899) );
  XNOR U9832 ( .A(n9937), .B(n9922), .Z(n9916) );
  XOR U9833 ( .A(p_input[2056]), .B(p_input[520]), .Z(n9922) );
  XOR U9834 ( .A(n9913), .B(n9921), .Z(n9937) );
  XOR U9835 ( .A(n9938), .B(n9918), .Z(n9921) );
  XOR U9836 ( .A(p_input[2054]), .B(p_input[518]), .Z(n9918) );
  XNOR U9837 ( .A(p_input[2055]), .B(p_input[519]), .Z(n9938) );
  XNOR U9838 ( .A(n6328), .B(p_input[514]), .Z(n9913) );
  XNOR U9839 ( .A(n9927), .B(n9926), .Z(n9917) );
  XOR U9840 ( .A(n9939), .B(n9923), .Z(n9926) );
  XOR U9841 ( .A(p_input[2051]), .B(p_input[515]), .Z(n9923) );
  XNOR U9842 ( .A(p_input[2052]), .B(p_input[516]), .Z(n9939) );
  XOR U9843 ( .A(p_input[2053]), .B(p_input[517]), .Z(n9927) );
  XOR U9844 ( .A(n9940), .B(n9941), .Z(n9828) );
  AND U9845 ( .A(n135), .B(n9942), .Z(n9941) );
  XNOR U9846 ( .A(n9943), .B(n9940), .Z(n9942) );
  XNOR U9847 ( .A(n9944), .B(n9945), .Z(n135) );
  AND U9848 ( .A(n9946), .B(n9947), .Z(n9945) );
  XOR U9849 ( .A(n9841), .B(n9944), .Z(n9947) );
  AND U9850 ( .A(n9948), .B(n9949), .Z(n9841) );
  XNOR U9851 ( .A(n9838), .B(n9944), .Z(n9946) );
  XOR U9852 ( .A(n9950), .B(n9951), .Z(n9838) );
  AND U9853 ( .A(n139), .B(n9952), .Z(n9951) );
  XOR U9854 ( .A(n9953), .B(n9950), .Z(n9952) );
  XOR U9855 ( .A(n9954), .B(n9955), .Z(n9944) );
  AND U9856 ( .A(n9956), .B(n9957), .Z(n9955) );
  XNOR U9857 ( .A(n9954), .B(n9948), .Z(n9957) );
  IV U9858 ( .A(n9856), .Z(n9948) );
  XOR U9859 ( .A(n9958), .B(n9959), .Z(n9856) );
  XOR U9860 ( .A(n9960), .B(n9949), .Z(n9959) );
  AND U9861 ( .A(n9883), .B(n9961), .Z(n9949) );
  AND U9862 ( .A(n9962), .B(n9963), .Z(n9960) );
  XOR U9863 ( .A(n9964), .B(n9958), .Z(n9962) );
  XNOR U9864 ( .A(n9853), .B(n9954), .Z(n9956) );
  XOR U9865 ( .A(n9965), .B(n9966), .Z(n9853) );
  AND U9866 ( .A(n139), .B(n9967), .Z(n9966) );
  XOR U9867 ( .A(n9968), .B(n9965), .Z(n9967) );
  XOR U9868 ( .A(n9969), .B(n9970), .Z(n9954) );
  AND U9869 ( .A(n9971), .B(n9972), .Z(n9970) );
  XNOR U9870 ( .A(n9969), .B(n9883), .Z(n9972) );
  XOR U9871 ( .A(n9973), .B(n9963), .Z(n9883) );
  XNOR U9872 ( .A(n9974), .B(n9958), .Z(n9963) );
  XOR U9873 ( .A(n9975), .B(n9976), .Z(n9958) );
  AND U9874 ( .A(n9977), .B(n9978), .Z(n9976) );
  XOR U9875 ( .A(n9979), .B(n9975), .Z(n9977) );
  XNOR U9876 ( .A(n9980), .B(n9981), .Z(n9974) );
  AND U9877 ( .A(n9982), .B(n9983), .Z(n9981) );
  XOR U9878 ( .A(n9980), .B(n9984), .Z(n9982) );
  XNOR U9879 ( .A(n9964), .B(n9961), .Z(n9973) );
  AND U9880 ( .A(n9985), .B(n9986), .Z(n9961) );
  XOR U9881 ( .A(n9987), .B(n9988), .Z(n9964) );
  AND U9882 ( .A(n9989), .B(n9990), .Z(n9988) );
  XOR U9883 ( .A(n9987), .B(n9991), .Z(n9989) );
  XNOR U9884 ( .A(n9880), .B(n9969), .Z(n9971) );
  XOR U9885 ( .A(n9992), .B(n9993), .Z(n9880) );
  AND U9886 ( .A(n139), .B(n9994), .Z(n9993) );
  XNOR U9887 ( .A(n9995), .B(n9992), .Z(n9994) );
  XOR U9888 ( .A(n9996), .B(n9997), .Z(n9969) );
  AND U9889 ( .A(n9998), .B(n9999), .Z(n9997) );
  XNOR U9890 ( .A(n9996), .B(n9985), .Z(n9999) );
  IV U9891 ( .A(n9931), .Z(n9985) );
  XNOR U9892 ( .A(n10000), .B(n9978), .Z(n9931) );
  XNOR U9893 ( .A(n10001), .B(n9984), .Z(n9978) );
  XOR U9894 ( .A(n10002), .B(n10003), .Z(n9984) );
  NOR U9895 ( .A(n10004), .B(n10005), .Z(n10003) );
  XNOR U9896 ( .A(n10002), .B(n10006), .Z(n10004) );
  XNOR U9897 ( .A(n9983), .B(n9975), .Z(n10001) );
  XOR U9898 ( .A(n10007), .B(n10008), .Z(n9975) );
  AND U9899 ( .A(n10009), .B(n10010), .Z(n10008) );
  XNOR U9900 ( .A(n10007), .B(n10011), .Z(n10009) );
  XNOR U9901 ( .A(n10012), .B(n9980), .Z(n9983) );
  XOR U9902 ( .A(n10013), .B(n10014), .Z(n9980) );
  AND U9903 ( .A(n10015), .B(n10016), .Z(n10014) );
  XOR U9904 ( .A(n10013), .B(n10017), .Z(n10015) );
  XNOR U9905 ( .A(n10018), .B(n10019), .Z(n10012) );
  NOR U9906 ( .A(n10020), .B(n10021), .Z(n10019) );
  XOR U9907 ( .A(n10018), .B(n10022), .Z(n10020) );
  XNOR U9908 ( .A(n9979), .B(n9986), .Z(n10000) );
  NOR U9909 ( .A(n9943), .B(n10023), .Z(n9986) );
  XOR U9910 ( .A(n9991), .B(n9990), .Z(n9979) );
  XNOR U9911 ( .A(n10024), .B(n9987), .Z(n9990) );
  XOR U9912 ( .A(n10025), .B(n10026), .Z(n9987) );
  AND U9913 ( .A(n10027), .B(n10028), .Z(n10026) );
  XOR U9914 ( .A(n10025), .B(n10029), .Z(n10027) );
  XNOR U9915 ( .A(n10030), .B(n10031), .Z(n10024) );
  NOR U9916 ( .A(n10032), .B(n10033), .Z(n10031) );
  XNOR U9917 ( .A(n10030), .B(n10034), .Z(n10032) );
  XOR U9918 ( .A(n10035), .B(n10036), .Z(n9991) );
  NOR U9919 ( .A(n10037), .B(n10038), .Z(n10036) );
  XNOR U9920 ( .A(n10035), .B(n10039), .Z(n10037) );
  XNOR U9921 ( .A(n9928), .B(n9996), .Z(n9998) );
  XOR U9922 ( .A(n10040), .B(n10041), .Z(n9928) );
  AND U9923 ( .A(n139), .B(n10042), .Z(n10041) );
  XOR U9924 ( .A(n10043), .B(n10040), .Z(n10042) );
  AND U9925 ( .A(n9940), .B(n9943), .Z(n9996) );
  XOR U9926 ( .A(n10044), .B(n10023), .Z(n9943) );
  XNOR U9927 ( .A(p_input[2048]), .B(p_input[528]), .Z(n10023) );
  XOR U9928 ( .A(n10011), .B(n10010), .Z(n10044) );
  XNOR U9929 ( .A(n10045), .B(n10017), .Z(n10010) );
  XNOR U9930 ( .A(n10006), .B(n10005), .Z(n10017) );
  XOR U9931 ( .A(n10046), .B(n10002), .Z(n10005) );
  XNOR U9932 ( .A(n6439), .B(p_input[538]), .Z(n10002) );
  XNOR U9933 ( .A(p_input[2059]), .B(p_input[539]), .Z(n10046) );
  XOR U9934 ( .A(p_input[2060]), .B(p_input[540]), .Z(n10006) );
  XNOR U9935 ( .A(n10016), .B(n10007), .Z(n10045) );
  XNOR U9936 ( .A(n6553), .B(p_input[529]), .Z(n10007) );
  XOR U9937 ( .A(n10047), .B(n10022), .Z(n10016) );
  XNOR U9938 ( .A(p_input[2063]), .B(p_input[543]), .Z(n10022) );
  XOR U9939 ( .A(n10013), .B(n10021), .Z(n10047) );
  XOR U9940 ( .A(n10048), .B(n10018), .Z(n10021) );
  XOR U9941 ( .A(p_input[2061]), .B(p_input[541]), .Z(n10018) );
  XNOR U9942 ( .A(p_input[2062]), .B(p_input[542]), .Z(n10048) );
  XNOR U9943 ( .A(n6325), .B(p_input[537]), .Z(n10013) );
  XNOR U9944 ( .A(n10029), .B(n10028), .Z(n10011) );
  XNOR U9945 ( .A(n10049), .B(n10034), .Z(n10028) );
  XOR U9946 ( .A(p_input[2056]), .B(p_input[536]), .Z(n10034) );
  XOR U9947 ( .A(n10025), .B(n10033), .Z(n10049) );
  XOR U9948 ( .A(n10050), .B(n10030), .Z(n10033) );
  XOR U9949 ( .A(p_input[2054]), .B(p_input[534]), .Z(n10030) );
  XNOR U9950 ( .A(p_input[2055]), .B(p_input[535]), .Z(n10050) );
  XNOR U9951 ( .A(n6328), .B(p_input[530]), .Z(n10025) );
  XNOR U9952 ( .A(n10039), .B(n10038), .Z(n10029) );
  XOR U9953 ( .A(n10051), .B(n10035), .Z(n10038) );
  XOR U9954 ( .A(p_input[2051]), .B(p_input[531]), .Z(n10035) );
  XNOR U9955 ( .A(p_input[2052]), .B(p_input[532]), .Z(n10051) );
  XOR U9956 ( .A(p_input[2053]), .B(p_input[533]), .Z(n10039) );
  XOR U9957 ( .A(n10052), .B(n10053), .Z(n9940) );
  AND U9958 ( .A(n139), .B(n10054), .Z(n10053) );
  XNOR U9959 ( .A(n10055), .B(n10052), .Z(n10054) );
  XNOR U9960 ( .A(n10056), .B(n10057), .Z(n139) );
  AND U9961 ( .A(n10058), .B(n10059), .Z(n10057) );
  XOR U9962 ( .A(n9953), .B(n10056), .Z(n10059) );
  AND U9963 ( .A(n10060), .B(n10061), .Z(n9953) );
  XNOR U9964 ( .A(n9950), .B(n10056), .Z(n10058) );
  XOR U9965 ( .A(n10062), .B(n10063), .Z(n9950) );
  AND U9966 ( .A(n143), .B(n10064), .Z(n10063) );
  XOR U9967 ( .A(n10065), .B(n10062), .Z(n10064) );
  XOR U9968 ( .A(n10066), .B(n10067), .Z(n10056) );
  AND U9969 ( .A(n10068), .B(n10069), .Z(n10067) );
  XNOR U9970 ( .A(n10066), .B(n10060), .Z(n10069) );
  IV U9971 ( .A(n9968), .Z(n10060) );
  XOR U9972 ( .A(n10070), .B(n10071), .Z(n9968) );
  XOR U9973 ( .A(n10072), .B(n10061), .Z(n10071) );
  AND U9974 ( .A(n9995), .B(n10073), .Z(n10061) );
  AND U9975 ( .A(n10074), .B(n10075), .Z(n10072) );
  XOR U9976 ( .A(n10076), .B(n10070), .Z(n10074) );
  XNOR U9977 ( .A(n9965), .B(n10066), .Z(n10068) );
  XOR U9978 ( .A(n10077), .B(n10078), .Z(n9965) );
  AND U9979 ( .A(n143), .B(n10079), .Z(n10078) );
  XOR U9980 ( .A(n10080), .B(n10077), .Z(n10079) );
  XOR U9981 ( .A(n10081), .B(n10082), .Z(n10066) );
  AND U9982 ( .A(n10083), .B(n10084), .Z(n10082) );
  XNOR U9983 ( .A(n10081), .B(n9995), .Z(n10084) );
  XOR U9984 ( .A(n10085), .B(n10075), .Z(n9995) );
  XNOR U9985 ( .A(n10086), .B(n10070), .Z(n10075) );
  XOR U9986 ( .A(n10087), .B(n10088), .Z(n10070) );
  AND U9987 ( .A(n10089), .B(n10090), .Z(n10088) );
  XOR U9988 ( .A(n10091), .B(n10087), .Z(n10089) );
  XNOR U9989 ( .A(n10092), .B(n10093), .Z(n10086) );
  AND U9990 ( .A(n10094), .B(n10095), .Z(n10093) );
  XOR U9991 ( .A(n10092), .B(n10096), .Z(n10094) );
  XNOR U9992 ( .A(n10076), .B(n10073), .Z(n10085) );
  AND U9993 ( .A(n10097), .B(n10098), .Z(n10073) );
  XOR U9994 ( .A(n10099), .B(n10100), .Z(n10076) );
  AND U9995 ( .A(n10101), .B(n10102), .Z(n10100) );
  XOR U9996 ( .A(n10099), .B(n10103), .Z(n10101) );
  XNOR U9997 ( .A(n9992), .B(n10081), .Z(n10083) );
  XOR U9998 ( .A(n10104), .B(n10105), .Z(n9992) );
  AND U9999 ( .A(n143), .B(n10106), .Z(n10105) );
  XNOR U10000 ( .A(n10107), .B(n10104), .Z(n10106) );
  XOR U10001 ( .A(n10108), .B(n10109), .Z(n10081) );
  AND U10002 ( .A(n10110), .B(n10111), .Z(n10109) );
  XNOR U10003 ( .A(n10108), .B(n10097), .Z(n10111) );
  IV U10004 ( .A(n10043), .Z(n10097) );
  XNOR U10005 ( .A(n10112), .B(n10090), .Z(n10043) );
  XNOR U10006 ( .A(n10113), .B(n10096), .Z(n10090) );
  XOR U10007 ( .A(n10114), .B(n10115), .Z(n10096) );
  NOR U10008 ( .A(n10116), .B(n10117), .Z(n10115) );
  XNOR U10009 ( .A(n10114), .B(n10118), .Z(n10116) );
  XNOR U10010 ( .A(n10095), .B(n10087), .Z(n10113) );
  XOR U10011 ( .A(n10119), .B(n10120), .Z(n10087) );
  AND U10012 ( .A(n10121), .B(n10122), .Z(n10120) );
  XNOR U10013 ( .A(n10119), .B(n10123), .Z(n10121) );
  XNOR U10014 ( .A(n10124), .B(n10092), .Z(n10095) );
  XOR U10015 ( .A(n10125), .B(n10126), .Z(n10092) );
  AND U10016 ( .A(n10127), .B(n10128), .Z(n10126) );
  XOR U10017 ( .A(n10125), .B(n10129), .Z(n10127) );
  XNOR U10018 ( .A(n10130), .B(n10131), .Z(n10124) );
  NOR U10019 ( .A(n10132), .B(n10133), .Z(n10131) );
  XOR U10020 ( .A(n10130), .B(n10134), .Z(n10132) );
  XNOR U10021 ( .A(n10091), .B(n10098), .Z(n10112) );
  NOR U10022 ( .A(n10055), .B(n10135), .Z(n10098) );
  XOR U10023 ( .A(n10103), .B(n10102), .Z(n10091) );
  XNOR U10024 ( .A(n10136), .B(n10099), .Z(n10102) );
  XOR U10025 ( .A(n10137), .B(n10138), .Z(n10099) );
  AND U10026 ( .A(n10139), .B(n10140), .Z(n10138) );
  XOR U10027 ( .A(n10137), .B(n10141), .Z(n10139) );
  XNOR U10028 ( .A(n10142), .B(n10143), .Z(n10136) );
  NOR U10029 ( .A(n10144), .B(n10145), .Z(n10143) );
  XNOR U10030 ( .A(n10142), .B(n10146), .Z(n10144) );
  XOR U10031 ( .A(n10147), .B(n10148), .Z(n10103) );
  NOR U10032 ( .A(n10149), .B(n10150), .Z(n10148) );
  XNOR U10033 ( .A(n10147), .B(n10151), .Z(n10149) );
  XNOR U10034 ( .A(n10040), .B(n10108), .Z(n10110) );
  XOR U10035 ( .A(n10152), .B(n10153), .Z(n10040) );
  AND U10036 ( .A(n143), .B(n10154), .Z(n10153) );
  XOR U10037 ( .A(n10155), .B(n10152), .Z(n10154) );
  AND U10038 ( .A(n10052), .B(n10055), .Z(n10108) );
  XOR U10039 ( .A(n10156), .B(n10135), .Z(n10055) );
  XNOR U10040 ( .A(p_input[2048]), .B(p_input[544]), .Z(n10135) );
  XOR U10041 ( .A(n10123), .B(n10122), .Z(n10156) );
  XNOR U10042 ( .A(n10157), .B(n10129), .Z(n10122) );
  XNOR U10043 ( .A(n10118), .B(n10117), .Z(n10129) );
  XOR U10044 ( .A(n10158), .B(n10114), .Z(n10117) );
  XNOR U10045 ( .A(n6439), .B(p_input[554]), .Z(n10114) );
  XNOR U10046 ( .A(p_input[2059]), .B(p_input[555]), .Z(n10158) );
  XOR U10047 ( .A(p_input[2060]), .B(p_input[556]), .Z(n10118) );
  XNOR U10048 ( .A(n10128), .B(n10119), .Z(n10157) );
  XNOR U10049 ( .A(n6553), .B(p_input[545]), .Z(n10119) );
  XOR U10050 ( .A(n10159), .B(n10134), .Z(n10128) );
  XNOR U10051 ( .A(p_input[2063]), .B(p_input[559]), .Z(n10134) );
  XOR U10052 ( .A(n10125), .B(n10133), .Z(n10159) );
  XOR U10053 ( .A(n10160), .B(n10130), .Z(n10133) );
  XOR U10054 ( .A(p_input[2061]), .B(p_input[557]), .Z(n10130) );
  XNOR U10055 ( .A(p_input[2062]), .B(p_input[558]), .Z(n10160) );
  XNOR U10056 ( .A(n6325), .B(p_input[553]), .Z(n10125) );
  XNOR U10057 ( .A(n10141), .B(n10140), .Z(n10123) );
  XNOR U10058 ( .A(n10161), .B(n10146), .Z(n10140) );
  XOR U10059 ( .A(p_input[2056]), .B(p_input[552]), .Z(n10146) );
  XOR U10060 ( .A(n10137), .B(n10145), .Z(n10161) );
  XOR U10061 ( .A(n10162), .B(n10142), .Z(n10145) );
  XOR U10062 ( .A(p_input[2054]), .B(p_input[550]), .Z(n10142) );
  XNOR U10063 ( .A(p_input[2055]), .B(p_input[551]), .Z(n10162) );
  XNOR U10064 ( .A(n6328), .B(p_input[546]), .Z(n10137) );
  XNOR U10065 ( .A(n10151), .B(n10150), .Z(n10141) );
  XOR U10066 ( .A(n10163), .B(n10147), .Z(n10150) );
  XOR U10067 ( .A(p_input[2051]), .B(p_input[547]), .Z(n10147) );
  XNOR U10068 ( .A(p_input[2052]), .B(p_input[548]), .Z(n10163) );
  XOR U10069 ( .A(p_input[2053]), .B(p_input[549]), .Z(n10151) );
  XOR U10070 ( .A(n10164), .B(n10165), .Z(n10052) );
  AND U10071 ( .A(n143), .B(n10166), .Z(n10165) );
  XNOR U10072 ( .A(n10167), .B(n10164), .Z(n10166) );
  XNOR U10073 ( .A(n10168), .B(n10169), .Z(n143) );
  AND U10074 ( .A(n10170), .B(n10171), .Z(n10169) );
  XOR U10075 ( .A(n10065), .B(n10168), .Z(n10171) );
  AND U10076 ( .A(n10172), .B(n10173), .Z(n10065) );
  XNOR U10077 ( .A(n10062), .B(n10168), .Z(n10170) );
  XOR U10078 ( .A(n10174), .B(n10175), .Z(n10062) );
  AND U10079 ( .A(n147), .B(n10176), .Z(n10175) );
  XOR U10080 ( .A(n10177), .B(n10174), .Z(n10176) );
  XOR U10081 ( .A(n10178), .B(n10179), .Z(n10168) );
  AND U10082 ( .A(n10180), .B(n10181), .Z(n10179) );
  XNOR U10083 ( .A(n10178), .B(n10172), .Z(n10181) );
  IV U10084 ( .A(n10080), .Z(n10172) );
  XOR U10085 ( .A(n10182), .B(n10183), .Z(n10080) );
  XOR U10086 ( .A(n10184), .B(n10173), .Z(n10183) );
  AND U10087 ( .A(n10107), .B(n10185), .Z(n10173) );
  AND U10088 ( .A(n10186), .B(n10187), .Z(n10184) );
  XOR U10089 ( .A(n10188), .B(n10182), .Z(n10186) );
  XNOR U10090 ( .A(n10077), .B(n10178), .Z(n10180) );
  XOR U10091 ( .A(n10189), .B(n10190), .Z(n10077) );
  AND U10092 ( .A(n147), .B(n10191), .Z(n10190) );
  XOR U10093 ( .A(n10192), .B(n10189), .Z(n10191) );
  XOR U10094 ( .A(n10193), .B(n10194), .Z(n10178) );
  AND U10095 ( .A(n10195), .B(n10196), .Z(n10194) );
  XNOR U10096 ( .A(n10193), .B(n10107), .Z(n10196) );
  XOR U10097 ( .A(n10197), .B(n10187), .Z(n10107) );
  XNOR U10098 ( .A(n10198), .B(n10182), .Z(n10187) );
  XOR U10099 ( .A(n10199), .B(n10200), .Z(n10182) );
  AND U10100 ( .A(n10201), .B(n10202), .Z(n10200) );
  XOR U10101 ( .A(n10203), .B(n10199), .Z(n10201) );
  XNOR U10102 ( .A(n10204), .B(n10205), .Z(n10198) );
  AND U10103 ( .A(n10206), .B(n10207), .Z(n10205) );
  XOR U10104 ( .A(n10204), .B(n10208), .Z(n10206) );
  XNOR U10105 ( .A(n10188), .B(n10185), .Z(n10197) );
  AND U10106 ( .A(n10209), .B(n10210), .Z(n10185) );
  XOR U10107 ( .A(n10211), .B(n10212), .Z(n10188) );
  AND U10108 ( .A(n10213), .B(n10214), .Z(n10212) );
  XOR U10109 ( .A(n10211), .B(n10215), .Z(n10213) );
  XNOR U10110 ( .A(n10104), .B(n10193), .Z(n10195) );
  XOR U10111 ( .A(n10216), .B(n10217), .Z(n10104) );
  AND U10112 ( .A(n147), .B(n10218), .Z(n10217) );
  XNOR U10113 ( .A(n10219), .B(n10216), .Z(n10218) );
  XOR U10114 ( .A(n10220), .B(n10221), .Z(n10193) );
  AND U10115 ( .A(n10222), .B(n10223), .Z(n10221) );
  XNOR U10116 ( .A(n10220), .B(n10209), .Z(n10223) );
  IV U10117 ( .A(n10155), .Z(n10209) );
  XNOR U10118 ( .A(n10224), .B(n10202), .Z(n10155) );
  XNOR U10119 ( .A(n10225), .B(n10208), .Z(n10202) );
  XOR U10120 ( .A(n10226), .B(n10227), .Z(n10208) );
  NOR U10121 ( .A(n10228), .B(n10229), .Z(n10227) );
  XNOR U10122 ( .A(n10226), .B(n10230), .Z(n10228) );
  XNOR U10123 ( .A(n10207), .B(n10199), .Z(n10225) );
  XOR U10124 ( .A(n10231), .B(n10232), .Z(n10199) );
  AND U10125 ( .A(n10233), .B(n10234), .Z(n10232) );
  XNOR U10126 ( .A(n10231), .B(n10235), .Z(n10233) );
  XNOR U10127 ( .A(n10236), .B(n10204), .Z(n10207) );
  XOR U10128 ( .A(n10237), .B(n10238), .Z(n10204) );
  AND U10129 ( .A(n10239), .B(n10240), .Z(n10238) );
  XOR U10130 ( .A(n10237), .B(n10241), .Z(n10239) );
  XNOR U10131 ( .A(n10242), .B(n10243), .Z(n10236) );
  NOR U10132 ( .A(n10244), .B(n10245), .Z(n10243) );
  XOR U10133 ( .A(n10242), .B(n10246), .Z(n10244) );
  XNOR U10134 ( .A(n10203), .B(n10210), .Z(n10224) );
  NOR U10135 ( .A(n10167), .B(n10247), .Z(n10210) );
  XOR U10136 ( .A(n10215), .B(n10214), .Z(n10203) );
  XNOR U10137 ( .A(n10248), .B(n10211), .Z(n10214) );
  XOR U10138 ( .A(n10249), .B(n10250), .Z(n10211) );
  AND U10139 ( .A(n10251), .B(n10252), .Z(n10250) );
  XOR U10140 ( .A(n10249), .B(n10253), .Z(n10251) );
  XNOR U10141 ( .A(n10254), .B(n10255), .Z(n10248) );
  NOR U10142 ( .A(n10256), .B(n10257), .Z(n10255) );
  XNOR U10143 ( .A(n10254), .B(n10258), .Z(n10256) );
  XOR U10144 ( .A(n10259), .B(n10260), .Z(n10215) );
  NOR U10145 ( .A(n10261), .B(n10262), .Z(n10260) );
  XNOR U10146 ( .A(n10259), .B(n10263), .Z(n10261) );
  XNOR U10147 ( .A(n10152), .B(n10220), .Z(n10222) );
  XOR U10148 ( .A(n10264), .B(n10265), .Z(n10152) );
  AND U10149 ( .A(n147), .B(n10266), .Z(n10265) );
  XOR U10150 ( .A(n10267), .B(n10264), .Z(n10266) );
  AND U10151 ( .A(n10164), .B(n10167), .Z(n10220) );
  XOR U10152 ( .A(n10268), .B(n10247), .Z(n10167) );
  XNOR U10153 ( .A(p_input[2048]), .B(p_input[560]), .Z(n10247) );
  XOR U10154 ( .A(n10235), .B(n10234), .Z(n10268) );
  XNOR U10155 ( .A(n10269), .B(n10241), .Z(n10234) );
  XNOR U10156 ( .A(n10230), .B(n10229), .Z(n10241) );
  XOR U10157 ( .A(n10270), .B(n10226), .Z(n10229) );
  XNOR U10158 ( .A(n6439), .B(p_input[570]), .Z(n10226) );
  XNOR U10159 ( .A(p_input[2059]), .B(p_input[571]), .Z(n10270) );
  XOR U10160 ( .A(p_input[2060]), .B(p_input[572]), .Z(n10230) );
  XNOR U10161 ( .A(n10240), .B(n10231), .Z(n10269) );
  XNOR U10162 ( .A(n6553), .B(p_input[561]), .Z(n10231) );
  XOR U10163 ( .A(n10271), .B(n10246), .Z(n10240) );
  XNOR U10164 ( .A(p_input[2063]), .B(p_input[575]), .Z(n10246) );
  XOR U10165 ( .A(n10237), .B(n10245), .Z(n10271) );
  XOR U10166 ( .A(n10272), .B(n10242), .Z(n10245) );
  XOR U10167 ( .A(p_input[2061]), .B(p_input[573]), .Z(n10242) );
  XNOR U10168 ( .A(p_input[2062]), .B(p_input[574]), .Z(n10272) );
  XNOR U10169 ( .A(n6325), .B(p_input[569]), .Z(n10237) );
  XNOR U10170 ( .A(n10253), .B(n10252), .Z(n10235) );
  XNOR U10171 ( .A(n10273), .B(n10258), .Z(n10252) );
  XOR U10172 ( .A(p_input[2056]), .B(p_input[568]), .Z(n10258) );
  XOR U10173 ( .A(n10249), .B(n10257), .Z(n10273) );
  XOR U10174 ( .A(n10274), .B(n10254), .Z(n10257) );
  XOR U10175 ( .A(p_input[2054]), .B(p_input[566]), .Z(n10254) );
  XNOR U10176 ( .A(p_input[2055]), .B(p_input[567]), .Z(n10274) );
  XNOR U10177 ( .A(n6328), .B(p_input[562]), .Z(n10249) );
  XNOR U10178 ( .A(n10263), .B(n10262), .Z(n10253) );
  XOR U10179 ( .A(n10275), .B(n10259), .Z(n10262) );
  XOR U10180 ( .A(p_input[2051]), .B(p_input[563]), .Z(n10259) );
  XNOR U10181 ( .A(p_input[2052]), .B(p_input[564]), .Z(n10275) );
  XOR U10182 ( .A(p_input[2053]), .B(p_input[565]), .Z(n10263) );
  XOR U10183 ( .A(n10276), .B(n10277), .Z(n10164) );
  AND U10184 ( .A(n147), .B(n10278), .Z(n10277) );
  XNOR U10185 ( .A(n10279), .B(n10276), .Z(n10278) );
  XNOR U10186 ( .A(n10280), .B(n10281), .Z(n147) );
  AND U10187 ( .A(n10282), .B(n10283), .Z(n10281) );
  XOR U10188 ( .A(n10177), .B(n10280), .Z(n10283) );
  AND U10189 ( .A(n10284), .B(n10285), .Z(n10177) );
  XNOR U10190 ( .A(n10174), .B(n10280), .Z(n10282) );
  XOR U10191 ( .A(n10286), .B(n10287), .Z(n10174) );
  AND U10192 ( .A(n151), .B(n10288), .Z(n10287) );
  XOR U10193 ( .A(n10289), .B(n10286), .Z(n10288) );
  XOR U10194 ( .A(n10290), .B(n10291), .Z(n10280) );
  AND U10195 ( .A(n10292), .B(n10293), .Z(n10291) );
  XNOR U10196 ( .A(n10290), .B(n10284), .Z(n10293) );
  IV U10197 ( .A(n10192), .Z(n10284) );
  XOR U10198 ( .A(n10294), .B(n10295), .Z(n10192) );
  XOR U10199 ( .A(n10296), .B(n10285), .Z(n10295) );
  AND U10200 ( .A(n10219), .B(n10297), .Z(n10285) );
  AND U10201 ( .A(n10298), .B(n10299), .Z(n10296) );
  XOR U10202 ( .A(n10300), .B(n10294), .Z(n10298) );
  XNOR U10203 ( .A(n10189), .B(n10290), .Z(n10292) );
  XOR U10204 ( .A(n10301), .B(n10302), .Z(n10189) );
  AND U10205 ( .A(n151), .B(n10303), .Z(n10302) );
  XOR U10206 ( .A(n10304), .B(n10301), .Z(n10303) );
  XOR U10207 ( .A(n10305), .B(n10306), .Z(n10290) );
  AND U10208 ( .A(n10307), .B(n10308), .Z(n10306) );
  XNOR U10209 ( .A(n10305), .B(n10219), .Z(n10308) );
  XOR U10210 ( .A(n10309), .B(n10299), .Z(n10219) );
  XNOR U10211 ( .A(n10310), .B(n10294), .Z(n10299) );
  XOR U10212 ( .A(n10311), .B(n10312), .Z(n10294) );
  AND U10213 ( .A(n10313), .B(n10314), .Z(n10312) );
  XOR U10214 ( .A(n10315), .B(n10311), .Z(n10313) );
  XNOR U10215 ( .A(n10316), .B(n10317), .Z(n10310) );
  AND U10216 ( .A(n10318), .B(n10319), .Z(n10317) );
  XOR U10217 ( .A(n10316), .B(n10320), .Z(n10318) );
  XNOR U10218 ( .A(n10300), .B(n10297), .Z(n10309) );
  AND U10219 ( .A(n10321), .B(n10322), .Z(n10297) );
  XOR U10220 ( .A(n10323), .B(n10324), .Z(n10300) );
  AND U10221 ( .A(n10325), .B(n10326), .Z(n10324) );
  XOR U10222 ( .A(n10323), .B(n10327), .Z(n10325) );
  XNOR U10223 ( .A(n10216), .B(n10305), .Z(n10307) );
  XOR U10224 ( .A(n10328), .B(n10329), .Z(n10216) );
  AND U10225 ( .A(n151), .B(n10330), .Z(n10329) );
  XNOR U10226 ( .A(n10331), .B(n10328), .Z(n10330) );
  XOR U10227 ( .A(n10332), .B(n10333), .Z(n10305) );
  AND U10228 ( .A(n10334), .B(n10335), .Z(n10333) );
  XNOR U10229 ( .A(n10332), .B(n10321), .Z(n10335) );
  IV U10230 ( .A(n10267), .Z(n10321) );
  XNOR U10231 ( .A(n10336), .B(n10314), .Z(n10267) );
  XNOR U10232 ( .A(n10337), .B(n10320), .Z(n10314) );
  XOR U10233 ( .A(n10338), .B(n10339), .Z(n10320) );
  NOR U10234 ( .A(n10340), .B(n10341), .Z(n10339) );
  XNOR U10235 ( .A(n10338), .B(n10342), .Z(n10340) );
  XNOR U10236 ( .A(n10319), .B(n10311), .Z(n10337) );
  XOR U10237 ( .A(n10343), .B(n10344), .Z(n10311) );
  AND U10238 ( .A(n10345), .B(n10346), .Z(n10344) );
  XNOR U10239 ( .A(n10343), .B(n10347), .Z(n10345) );
  XNOR U10240 ( .A(n10348), .B(n10316), .Z(n10319) );
  XOR U10241 ( .A(n10349), .B(n10350), .Z(n10316) );
  AND U10242 ( .A(n10351), .B(n10352), .Z(n10350) );
  XOR U10243 ( .A(n10349), .B(n10353), .Z(n10351) );
  XNOR U10244 ( .A(n10354), .B(n10355), .Z(n10348) );
  NOR U10245 ( .A(n10356), .B(n10357), .Z(n10355) );
  XOR U10246 ( .A(n10354), .B(n10358), .Z(n10356) );
  XNOR U10247 ( .A(n10315), .B(n10322), .Z(n10336) );
  NOR U10248 ( .A(n10279), .B(n10359), .Z(n10322) );
  XOR U10249 ( .A(n10327), .B(n10326), .Z(n10315) );
  XNOR U10250 ( .A(n10360), .B(n10323), .Z(n10326) );
  XOR U10251 ( .A(n10361), .B(n10362), .Z(n10323) );
  AND U10252 ( .A(n10363), .B(n10364), .Z(n10362) );
  XOR U10253 ( .A(n10361), .B(n10365), .Z(n10363) );
  XNOR U10254 ( .A(n10366), .B(n10367), .Z(n10360) );
  NOR U10255 ( .A(n10368), .B(n10369), .Z(n10367) );
  XNOR U10256 ( .A(n10366), .B(n10370), .Z(n10368) );
  XOR U10257 ( .A(n10371), .B(n10372), .Z(n10327) );
  NOR U10258 ( .A(n10373), .B(n10374), .Z(n10372) );
  XNOR U10259 ( .A(n10371), .B(n10375), .Z(n10373) );
  XNOR U10260 ( .A(n10264), .B(n10332), .Z(n10334) );
  XOR U10261 ( .A(n10376), .B(n10377), .Z(n10264) );
  AND U10262 ( .A(n151), .B(n10378), .Z(n10377) );
  XOR U10263 ( .A(n10379), .B(n10376), .Z(n10378) );
  AND U10264 ( .A(n10276), .B(n10279), .Z(n10332) );
  XOR U10265 ( .A(n10380), .B(n10359), .Z(n10279) );
  XNOR U10266 ( .A(p_input[2048]), .B(p_input[576]), .Z(n10359) );
  XOR U10267 ( .A(n10347), .B(n10346), .Z(n10380) );
  XNOR U10268 ( .A(n10381), .B(n10353), .Z(n10346) );
  XNOR U10269 ( .A(n10342), .B(n10341), .Z(n10353) );
  XOR U10270 ( .A(n10382), .B(n10338), .Z(n10341) );
  XNOR U10271 ( .A(n6439), .B(p_input[586]), .Z(n10338) );
  XNOR U10272 ( .A(p_input[2059]), .B(p_input[587]), .Z(n10382) );
  XOR U10273 ( .A(p_input[2060]), .B(p_input[588]), .Z(n10342) );
  XNOR U10274 ( .A(n10352), .B(n10343), .Z(n10381) );
  XNOR U10275 ( .A(n6553), .B(p_input[577]), .Z(n10343) );
  XOR U10276 ( .A(n10383), .B(n10358), .Z(n10352) );
  XNOR U10277 ( .A(p_input[2063]), .B(p_input[591]), .Z(n10358) );
  XOR U10278 ( .A(n10349), .B(n10357), .Z(n10383) );
  XOR U10279 ( .A(n10384), .B(n10354), .Z(n10357) );
  XOR U10280 ( .A(p_input[2061]), .B(p_input[589]), .Z(n10354) );
  XNOR U10281 ( .A(p_input[2062]), .B(p_input[590]), .Z(n10384) );
  XNOR U10282 ( .A(n6325), .B(p_input[585]), .Z(n10349) );
  XNOR U10283 ( .A(n10365), .B(n10364), .Z(n10347) );
  XNOR U10284 ( .A(n10385), .B(n10370), .Z(n10364) );
  XOR U10285 ( .A(p_input[2056]), .B(p_input[584]), .Z(n10370) );
  XOR U10286 ( .A(n10361), .B(n10369), .Z(n10385) );
  XOR U10287 ( .A(n10386), .B(n10366), .Z(n10369) );
  XOR U10288 ( .A(p_input[2054]), .B(p_input[582]), .Z(n10366) );
  XNOR U10289 ( .A(p_input[2055]), .B(p_input[583]), .Z(n10386) );
  XNOR U10290 ( .A(n6328), .B(p_input[578]), .Z(n10361) );
  XNOR U10291 ( .A(n10375), .B(n10374), .Z(n10365) );
  XOR U10292 ( .A(n10387), .B(n10371), .Z(n10374) );
  XOR U10293 ( .A(p_input[2051]), .B(p_input[579]), .Z(n10371) );
  XNOR U10294 ( .A(p_input[2052]), .B(p_input[580]), .Z(n10387) );
  XOR U10295 ( .A(p_input[2053]), .B(p_input[581]), .Z(n10375) );
  XOR U10296 ( .A(n10388), .B(n10389), .Z(n10276) );
  AND U10297 ( .A(n151), .B(n10390), .Z(n10389) );
  XNOR U10298 ( .A(n10391), .B(n10388), .Z(n10390) );
  XNOR U10299 ( .A(n10392), .B(n10393), .Z(n151) );
  AND U10300 ( .A(n10394), .B(n10395), .Z(n10393) );
  XOR U10301 ( .A(n10289), .B(n10392), .Z(n10395) );
  AND U10302 ( .A(n10396), .B(n10397), .Z(n10289) );
  XNOR U10303 ( .A(n10286), .B(n10392), .Z(n10394) );
  XOR U10304 ( .A(n10398), .B(n10399), .Z(n10286) );
  AND U10305 ( .A(n155), .B(n10400), .Z(n10399) );
  XOR U10306 ( .A(n10401), .B(n10398), .Z(n10400) );
  XOR U10307 ( .A(n10402), .B(n10403), .Z(n10392) );
  AND U10308 ( .A(n10404), .B(n10405), .Z(n10403) );
  XNOR U10309 ( .A(n10402), .B(n10396), .Z(n10405) );
  IV U10310 ( .A(n10304), .Z(n10396) );
  XOR U10311 ( .A(n10406), .B(n10407), .Z(n10304) );
  XOR U10312 ( .A(n10408), .B(n10397), .Z(n10407) );
  AND U10313 ( .A(n10331), .B(n10409), .Z(n10397) );
  AND U10314 ( .A(n10410), .B(n10411), .Z(n10408) );
  XOR U10315 ( .A(n10412), .B(n10406), .Z(n10410) );
  XNOR U10316 ( .A(n10301), .B(n10402), .Z(n10404) );
  XOR U10317 ( .A(n10413), .B(n10414), .Z(n10301) );
  AND U10318 ( .A(n155), .B(n10415), .Z(n10414) );
  XOR U10319 ( .A(n10416), .B(n10413), .Z(n10415) );
  XOR U10320 ( .A(n10417), .B(n10418), .Z(n10402) );
  AND U10321 ( .A(n10419), .B(n10420), .Z(n10418) );
  XNOR U10322 ( .A(n10417), .B(n10331), .Z(n10420) );
  XOR U10323 ( .A(n10421), .B(n10411), .Z(n10331) );
  XNOR U10324 ( .A(n10422), .B(n10406), .Z(n10411) );
  XOR U10325 ( .A(n10423), .B(n10424), .Z(n10406) );
  AND U10326 ( .A(n10425), .B(n10426), .Z(n10424) );
  XOR U10327 ( .A(n10427), .B(n10423), .Z(n10425) );
  XNOR U10328 ( .A(n10428), .B(n10429), .Z(n10422) );
  AND U10329 ( .A(n10430), .B(n10431), .Z(n10429) );
  XOR U10330 ( .A(n10428), .B(n10432), .Z(n10430) );
  XNOR U10331 ( .A(n10412), .B(n10409), .Z(n10421) );
  AND U10332 ( .A(n10433), .B(n10434), .Z(n10409) );
  XOR U10333 ( .A(n10435), .B(n10436), .Z(n10412) );
  AND U10334 ( .A(n10437), .B(n10438), .Z(n10436) );
  XOR U10335 ( .A(n10435), .B(n10439), .Z(n10437) );
  XNOR U10336 ( .A(n10328), .B(n10417), .Z(n10419) );
  XOR U10337 ( .A(n10440), .B(n10441), .Z(n10328) );
  AND U10338 ( .A(n155), .B(n10442), .Z(n10441) );
  XNOR U10339 ( .A(n10443), .B(n10440), .Z(n10442) );
  XOR U10340 ( .A(n10444), .B(n10445), .Z(n10417) );
  AND U10341 ( .A(n10446), .B(n10447), .Z(n10445) );
  XNOR U10342 ( .A(n10444), .B(n10433), .Z(n10447) );
  IV U10343 ( .A(n10379), .Z(n10433) );
  XNOR U10344 ( .A(n10448), .B(n10426), .Z(n10379) );
  XNOR U10345 ( .A(n10449), .B(n10432), .Z(n10426) );
  XOR U10346 ( .A(n10450), .B(n10451), .Z(n10432) );
  NOR U10347 ( .A(n10452), .B(n10453), .Z(n10451) );
  XNOR U10348 ( .A(n10450), .B(n10454), .Z(n10452) );
  XNOR U10349 ( .A(n10431), .B(n10423), .Z(n10449) );
  XOR U10350 ( .A(n10455), .B(n10456), .Z(n10423) );
  AND U10351 ( .A(n10457), .B(n10458), .Z(n10456) );
  XNOR U10352 ( .A(n10455), .B(n10459), .Z(n10457) );
  XNOR U10353 ( .A(n10460), .B(n10428), .Z(n10431) );
  XOR U10354 ( .A(n10461), .B(n10462), .Z(n10428) );
  AND U10355 ( .A(n10463), .B(n10464), .Z(n10462) );
  XOR U10356 ( .A(n10461), .B(n10465), .Z(n10463) );
  XNOR U10357 ( .A(n10466), .B(n10467), .Z(n10460) );
  NOR U10358 ( .A(n10468), .B(n10469), .Z(n10467) );
  XOR U10359 ( .A(n10466), .B(n10470), .Z(n10468) );
  XNOR U10360 ( .A(n10427), .B(n10434), .Z(n10448) );
  NOR U10361 ( .A(n10391), .B(n10471), .Z(n10434) );
  XOR U10362 ( .A(n10439), .B(n10438), .Z(n10427) );
  XNOR U10363 ( .A(n10472), .B(n10435), .Z(n10438) );
  XOR U10364 ( .A(n10473), .B(n10474), .Z(n10435) );
  AND U10365 ( .A(n10475), .B(n10476), .Z(n10474) );
  XOR U10366 ( .A(n10473), .B(n10477), .Z(n10475) );
  XNOR U10367 ( .A(n10478), .B(n10479), .Z(n10472) );
  NOR U10368 ( .A(n10480), .B(n10481), .Z(n10479) );
  XNOR U10369 ( .A(n10478), .B(n10482), .Z(n10480) );
  XOR U10370 ( .A(n10483), .B(n10484), .Z(n10439) );
  NOR U10371 ( .A(n10485), .B(n10486), .Z(n10484) );
  XNOR U10372 ( .A(n10483), .B(n10487), .Z(n10485) );
  XNOR U10373 ( .A(n10376), .B(n10444), .Z(n10446) );
  XOR U10374 ( .A(n10488), .B(n10489), .Z(n10376) );
  AND U10375 ( .A(n155), .B(n10490), .Z(n10489) );
  XOR U10376 ( .A(n10491), .B(n10488), .Z(n10490) );
  AND U10377 ( .A(n10388), .B(n10391), .Z(n10444) );
  XOR U10378 ( .A(n10492), .B(n10471), .Z(n10391) );
  XNOR U10379 ( .A(p_input[2048]), .B(p_input[592]), .Z(n10471) );
  XOR U10380 ( .A(n10459), .B(n10458), .Z(n10492) );
  XNOR U10381 ( .A(n10493), .B(n10465), .Z(n10458) );
  XNOR U10382 ( .A(n10454), .B(n10453), .Z(n10465) );
  XOR U10383 ( .A(n10494), .B(n10450), .Z(n10453) );
  XNOR U10384 ( .A(n6439), .B(p_input[602]), .Z(n10450) );
  XNOR U10385 ( .A(p_input[2059]), .B(p_input[603]), .Z(n10494) );
  XOR U10386 ( .A(p_input[2060]), .B(p_input[604]), .Z(n10454) );
  XNOR U10387 ( .A(n10464), .B(n10455), .Z(n10493) );
  XNOR U10388 ( .A(n6553), .B(p_input[593]), .Z(n10455) );
  XOR U10389 ( .A(n10495), .B(n10470), .Z(n10464) );
  XNOR U10390 ( .A(p_input[2063]), .B(p_input[607]), .Z(n10470) );
  XOR U10391 ( .A(n10461), .B(n10469), .Z(n10495) );
  XOR U10392 ( .A(n10496), .B(n10466), .Z(n10469) );
  XOR U10393 ( .A(p_input[2061]), .B(p_input[605]), .Z(n10466) );
  XNOR U10394 ( .A(p_input[2062]), .B(p_input[606]), .Z(n10496) );
  XNOR U10395 ( .A(n6325), .B(p_input[601]), .Z(n10461) );
  XNOR U10396 ( .A(n10477), .B(n10476), .Z(n10459) );
  XNOR U10397 ( .A(n10497), .B(n10482), .Z(n10476) );
  XOR U10398 ( .A(p_input[2056]), .B(p_input[600]), .Z(n10482) );
  XOR U10399 ( .A(n10473), .B(n10481), .Z(n10497) );
  XOR U10400 ( .A(n10498), .B(n10478), .Z(n10481) );
  XOR U10401 ( .A(p_input[2054]), .B(p_input[598]), .Z(n10478) );
  XNOR U10402 ( .A(p_input[2055]), .B(p_input[599]), .Z(n10498) );
  XNOR U10403 ( .A(n6328), .B(p_input[594]), .Z(n10473) );
  XNOR U10404 ( .A(n10487), .B(n10486), .Z(n10477) );
  XOR U10405 ( .A(n10499), .B(n10483), .Z(n10486) );
  XOR U10406 ( .A(p_input[2051]), .B(p_input[595]), .Z(n10483) );
  XNOR U10407 ( .A(p_input[2052]), .B(p_input[596]), .Z(n10499) );
  XOR U10408 ( .A(p_input[2053]), .B(p_input[597]), .Z(n10487) );
  XOR U10409 ( .A(n10500), .B(n10501), .Z(n10388) );
  AND U10410 ( .A(n155), .B(n10502), .Z(n10501) );
  XNOR U10411 ( .A(n10503), .B(n10500), .Z(n10502) );
  XNOR U10412 ( .A(n10504), .B(n10505), .Z(n155) );
  AND U10413 ( .A(n10506), .B(n10507), .Z(n10505) );
  XOR U10414 ( .A(n10401), .B(n10504), .Z(n10507) );
  AND U10415 ( .A(n10508), .B(n10509), .Z(n10401) );
  XNOR U10416 ( .A(n10398), .B(n10504), .Z(n10506) );
  XOR U10417 ( .A(n10510), .B(n10511), .Z(n10398) );
  AND U10418 ( .A(n159), .B(n10512), .Z(n10511) );
  XOR U10419 ( .A(n10513), .B(n10510), .Z(n10512) );
  XOR U10420 ( .A(n10514), .B(n10515), .Z(n10504) );
  AND U10421 ( .A(n10516), .B(n10517), .Z(n10515) );
  XNOR U10422 ( .A(n10514), .B(n10508), .Z(n10517) );
  IV U10423 ( .A(n10416), .Z(n10508) );
  XOR U10424 ( .A(n10518), .B(n10519), .Z(n10416) );
  XOR U10425 ( .A(n10520), .B(n10509), .Z(n10519) );
  AND U10426 ( .A(n10443), .B(n10521), .Z(n10509) );
  AND U10427 ( .A(n10522), .B(n10523), .Z(n10520) );
  XOR U10428 ( .A(n10524), .B(n10518), .Z(n10522) );
  XNOR U10429 ( .A(n10413), .B(n10514), .Z(n10516) );
  XOR U10430 ( .A(n10525), .B(n10526), .Z(n10413) );
  AND U10431 ( .A(n159), .B(n10527), .Z(n10526) );
  XOR U10432 ( .A(n10528), .B(n10525), .Z(n10527) );
  XOR U10433 ( .A(n10529), .B(n10530), .Z(n10514) );
  AND U10434 ( .A(n10531), .B(n10532), .Z(n10530) );
  XNOR U10435 ( .A(n10529), .B(n10443), .Z(n10532) );
  XOR U10436 ( .A(n10533), .B(n10523), .Z(n10443) );
  XNOR U10437 ( .A(n10534), .B(n10518), .Z(n10523) );
  XOR U10438 ( .A(n10535), .B(n10536), .Z(n10518) );
  AND U10439 ( .A(n10537), .B(n10538), .Z(n10536) );
  XOR U10440 ( .A(n10539), .B(n10535), .Z(n10537) );
  XNOR U10441 ( .A(n10540), .B(n10541), .Z(n10534) );
  AND U10442 ( .A(n10542), .B(n10543), .Z(n10541) );
  XOR U10443 ( .A(n10540), .B(n10544), .Z(n10542) );
  XNOR U10444 ( .A(n10524), .B(n10521), .Z(n10533) );
  AND U10445 ( .A(n10545), .B(n10546), .Z(n10521) );
  XOR U10446 ( .A(n10547), .B(n10548), .Z(n10524) );
  AND U10447 ( .A(n10549), .B(n10550), .Z(n10548) );
  XOR U10448 ( .A(n10547), .B(n10551), .Z(n10549) );
  XNOR U10449 ( .A(n10440), .B(n10529), .Z(n10531) );
  XOR U10450 ( .A(n10552), .B(n10553), .Z(n10440) );
  AND U10451 ( .A(n159), .B(n10554), .Z(n10553) );
  XNOR U10452 ( .A(n10555), .B(n10552), .Z(n10554) );
  XOR U10453 ( .A(n10556), .B(n10557), .Z(n10529) );
  AND U10454 ( .A(n10558), .B(n10559), .Z(n10557) );
  XNOR U10455 ( .A(n10556), .B(n10545), .Z(n10559) );
  IV U10456 ( .A(n10491), .Z(n10545) );
  XNOR U10457 ( .A(n10560), .B(n10538), .Z(n10491) );
  XNOR U10458 ( .A(n10561), .B(n10544), .Z(n10538) );
  XOR U10459 ( .A(n10562), .B(n10563), .Z(n10544) );
  NOR U10460 ( .A(n10564), .B(n10565), .Z(n10563) );
  XNOR U10461 ( .A(n10562), .B(n10566), .Z(n10564) );
  XNOR U10462 ( .A(n10543), .B(n10535), .Z(n10561) );
  XOR U10463 ( .A(n10567), .B(n10568), .Z(n10535) );
  AND U10464 ( .A(n10569), .B(n10570), .Z(n10568) );
  XNOR U10465 ( .A(n10567), .B(n10571), .Z(n10569) );
  XNOR U10466 ( .A(n10572), .B(n10540), .Z(n10543) );
  XOR U10467 ( .A(n10573), .B(n10574), .Z(n10540) );
  AND U10468 ( .A(n10575), .B(n10576), .Z(n10574) );
  XOR U10469 ( .A(n10573), .B(n10577), .Z(n10575) );
  XNOR U10470 ( .A(n10578), .B(n10579), .Z(n10572) );
  NOR U10471 ( .A(n10580), .B(n10581), .Z(n10579) );
  XOR U10472 ( .A(n10578), .B(n10582), .Z(n10580) );
  XNOR U10473 ( .A(n10539), .B(n10546), .Z(n10560) );
  NOR U10474 ( .A(n10503), .B(n10583), .Z(n10546) );
  XOR U10475 ( .A(n10551), .B(n10550), .Z(n10539) );
  XNOR U10476 ( .A(n10584), .B(n10547), .Z(n10550) );
  XOR U10477 ( .A(n10585), .B(n10586), .Z(n10547) );
  AND U10478 ( .A(n10587), .B(n10588), .Z(n10586) );
  XOR U10479 ( .A(n10585), .B(n10589), .Z(n10587) );
  XNOR U10480 ( .A(n10590), .B(n10591), .Z(n10584) );
  NOR U10481 ( .A(n10592), .B(n10593), .Z(n10591) );
  XNOR U10482 ( .A(n10590), .B(n10594), .Z(n10592) );
  XOR U10483 ( .A(n10595), .B(n10596), .Z(n10551) );
  NOR U10484 ( .A(n10597), .B(n10598), .Z(n10596) );
  XNOR U10485 ( .A(n10595), .B(n10599), .Z(n10597) );
  XNOR U10486 ( .A(n10488), .B(n10556), .Z(n10558) );
  XOR U10487 ( .A(n10600), .B(n10601), .Z(n10488) );
  AND U10488 ( .A(n159), .B(n10602), .Z(n10601) );
  XOR U10489 ( .A(n10603), .B(n10600), .Z(n10602) );
  AND U10490 ( .A(n10500), .B(n10503), .Z(n10556) );
  XOR U10491 ( .A(n10604), .B(n10583), .Z(n10503) );
  XNOR U10492 ( .A(p_input[2048]), .B(p_input[608]), .Z(n10583) );
  XOR U10493 ( .A(n10571), .B(n10570), .Z(n10604) );
  XNOR U10494 ( .A(n10605), .B(n10577), .Z(n10570) );
  XNOR U10495 ( .A(n10566), .B(n10565), .Z(n10577) );
  XOR U10496 ( .A(n10606), .B(n10562), .Z(n10565) );
  XNOR U10497 ( .A(n6439), .B(p_input[618]), .Z(n10562) );
  XNOR U10498 ( .A(p_input[2059]), .B(p_input[619]), .Z(n10606) );
  XOR U10499 ( .A(p_input[2060]), .B(p_input[620]), .Z(n10566) );
  XNOR U10500 ( .A(n10576), .B(n10567), .Z(n10605) );
  XNOR U10501 ( .A(n6553), .B(p_input[609]), .Z(n10567) );
  XOR U10502 ( .A(n10607), .B(n10582), .Z(n10576) );
  XNOR U10503 ( .A(p_input[2063]), .B(p_input[623]), .Z(n10582) );
  XOR U10504 ( .A(n10573), .B(n10581), .Z(n10607) );
  XOR U10505 ( .A(n10608), .B(n10578), .Z(n10581) );
  XOR U10506 ( .A(p_input[2061]), .B(p_input[621]), .Z(n10578) );
  XNOR U10507 ( .A(p_input[2062]), .B(p_input[622]), .Z(n10608) );
  XNOR U10508 ( .A(n6325), .B(p_input[617]), .Z(n10573) );
  XNOR U10509 ( .A(n10589), .B(n10588), .Z(n10571) );
  XNOR U10510 ( .A(n10609), .B(n10594), .Z(n10588) );
  XOR U10511 ( .A(p_input[2056]), .B(p_input[616]), .Z(n10594) );
  XOR U10512 ( .A(n10585), .B(n10593), .Z(n10609) );
  XOR U10513 ( .A(n10610), .B(n10590), .Z(n10593) );
  XOR U10514 ( .A(p_input[2054]), .B(p_input[614]), .Z(n10590) );
  XNOR U10515 ( .A(p_input[2055]), .B(p_input[615]), .Z(n10610) );
  XNOR U10516 ( .A(n6328), .B(p_input[610]), .Z(n10585) );
  XNOR U10517 ( .A(n10599), .B(n10598), .Z(n10589) );
  XOR U10518 ( .A(n10611), .B(n10595), .Z(n10598) );
  XOR U10519 ( .A(p_input[2051]), .B(p_input[611]), .Z(n10595) );
  XNOR U10520 ( .A(p_input[2052]), .B(p_input[612]), .Z(n10611) );
  XOR U10521 ( .A(p_input[2053]), .B(p_input[613]), .Z(n10599) );
  XOR U10522 ( .A(n10612), .B(n10613), .Z(n10500) );
  AND U10523 ( .A(n159), .B(n10614), .Z(n10613) );
  XNOR U10524 ( .A(n10615), .B(n10612), .Z(n10614) );
  XNOR U10525 ( .A(n10616), .B(n10617), .Z(n159) );
  AND U10526 ( .A(n10618), .B(n10619), .Z(n10617) );
  XOR U10527 ( .A(n10513), .B(n10616), .Z(n10619) );
  AND U10528 ( .A(n10620), .B(n10621), .Z(n10513) );
  XNOR U10529 ( .A(n10510), .B(n10616), .Z(n10618) );
  XOR U10530 ( .A(n10622), .B(n10623), .Z(n10510) );
  AND U10531 ( .A(n163), .B(n10624), .Z(n10623) );
  XOR U10532 ( .A(n10625), .B(n10622), .Z(n10624) );
  XOR U10533 ( .A(n10626), .B(n10627), .Z(n10616) );
  AND U10534 ( .A(n10628), .B(n10629), .Z(n10627) );
  XNOR U10535 ( .A(n10626), .B(n10620), .Z(n10629) );
  IV U10536 ( .A(n10528), .Z(n10620) );
  XOR U10537 ( .A(n10630), .B(n10631), .Z(n10528) );
  XOR U10538 ( .A(n10632), .B(n10621), .Z(n10631) );
  AND U10539 ( .A(n10555), .B(n10633), .Z(n10621) );
  AND U10540 ( .A(n10634), .B(n10635), .Z(n10632) );
  XOR U10541 ( .A(n10636), .B(n10630), .Z(n10634) );
  XNOR U10542 ( .A(n10525), .B(n10626), .Z(n10628) );
  XOR U10543 ( .A(n10637), .B(n10638), .Z(n10525) );
  AND U10544 ( .A(n163), .B(n10639), .Z(n10638) );
  XOR U10545 ( .A(n10640), .B(n10637), .Z(n10639) );
  XOR U10546 ( .A(n10641), .B(n10642), .Z(n10626) );
  AND U10547 ( .A(n10643), .B(n10644), .Z(n10642) );
  XNOR U10548 ( .A(n10641), .B(n10555), .Z(n10644) );
  XOR U10549 ( .A(n10645), .B(n10635), .Z(n10555) );
  XNOR U10550 ( .A(n10646), .B(n10630), .Z(n10635) );
  XOR U10551 ( .A(n10647), .B(n10648), .Z(n10630) );
  AND U10552 ( .A(n10649), .B(n10650), .Z(n10648) );
  XOR U10553 ( .A(n10651), .B(n10647), .Z(n10649) );
  XNOR U10554 ( .A(n10652), .B(n10653), .Z(n10646) );
  AND U10555 ( .A(n10654), .B(n10655), .Z(n10653) );
  XOR U10556 ( .A(n10652), .B(n10656), .Z(n10654) );
  XNOR U10557 ( .A(n10636), .B(n10633), .Z(n10645) );
  AND U10558 ( .A(n10657), .B(n10658), .Z(n10633) );
  XOR U10559 ( .A(n10659), .B(n10660), .Z(n10636) );
  AND U10560 ( .A(n10661), .B(n10662), .Z(n10660) );
  XOR U10561 ( .A(n10659), .B(n10663), .Z(n10661) );
  XNOR U10562 ( .A(n10552), .B(n10641), .Z(n10643) );
  XOR U10563 ( .A(n10664), .B(n10665), .Z(n10552) );
  AND U10564 ( .A(n163), .B(n10666), .Z(n10665) );
  XNOR U10565 ( .A(n10667), .B(n10664), .Z(n10666) );
  XOR U10566 ( .A(n10668), .B(n10669), .Z(n10641) );
  AND U10567 ( .A(n10670), .B(n10671), .Z(n10669) );
  XNOR U10568 ( .A(n10668), .B(n10657), .Z(n10671) );
  IV U10569 ( .A(n10603), .Z(n10657) );
  XNOR U10570 ( .A(n10672), .B(n10650), .Z(n10603) );
  XNOR U10571 ( .A(n10673), .B(n10656), .Z(n10650) );
  XOR U10572 ( .A(n10674), .B(n10675), .Z(n10656) );
  NOR U10573 ( .A(n10676), .B(n10677), .Z(n10675) );
  XNOR U10574 ( .A(n10674), .B(n10678), .Z(n10676) );
  XNOR U10575 ( .A(n10655), .B(n10647), .Z(n10673) );
  XOR U10576 ( .A(n10679), .B(n10680), .Z(n10647) );
  AND U10577 ( .A(n10681), .B(n10682), .Z(n10680) );
  XNOR U10578 ( .A(n10679), .B(n10683), .Z(n10681) );
  XNOR U10579 ( .A(n10684), .B(n10652), .Z(n10655) );
  XOR U10580 ( .A(n10685), .B(n10686), .Z(n10652) );
  AND U10581 ( .A(n10687), .B(n10688), .Z(n10686) );
  XOR U10582 ( .A(n10685), .B(n10689), .Z(n10687) );
  XNOR U10583 ( .A(n10690), .B(n10691), .Z(n10684) );
  NOR U10584 ( .A(n10692), .B(n10693), .Z(n10691) );
  XOR U10585 ( .A(n10690), .B(n10694), .Z(n10692) );
  XNOR U10586 ( .A(n10651), .B(n10658), .Z(n10672) );
  NOR U10587 ( .A(n10615), .B(n10695), .Z(n10658) );
  XOR U10588 ( .A(n10663), .B(n10662), .Z(n10651) );
  XNOR U10589 ( .A(n10696), .B(n10659), .Z(n10662) );
  XOR U10590 ( .A(n10697), .B(n10698), .Z(n10659) );
  AND U10591 ( .A(n10699), .B(n10700), .Z(n10698) );
  XOR U10592 ( .A(n10697), .B(n10701), .Z(n10699) );
  XNOR U10593 ( .A(n10702), .B(n10703), .Z(n10696) );
  NOR U10594 ( .A(n10704), .B(n10705), .Z(n10703) );
  XNOR U10595 ( .A(n10702), .B(n10706), .Z(n10704) );
  XOR U10596 ( .A(n10707), .B(n10708), .Z(n10663) );
  NOR U10597 ( .A(n10709), .B(n10710), .Z(n10708) );
  XNOR U10598 ( .A(n10707), .B(n10711), .Z(n10709) );
  XNOR U10599 ( .A(n10600), .B(n10668), .Z(n10670) );
  XOR U10600 ( .A(n10712), .B(n10713), .Z(n10600) );
  AND U10601 ( .A(n163), .B(n10714), .Z(n10713) );
  XOR U10602 ( .A(n10715), .B(n10712), .Z(n10714) );
  AND U10603 ( .A(n10612), .B(n10615), .Z(n10668) );
  XOR U10604 ( .A(n10716), .B(n10695), .Z(n10615) );
  XNOR U10605 ( .A(p_input[2048]), .B(p_input[624]), .Z(n10695) );
  XOR U10606 ( .A(n10683), .B(n10682), .Z(n10716) );
  XNOR U10607 ( .A(n10717), .B(n10689), .Z(n10682) );
  XNOR U10608 ( .A(n10678), .B(n10677), .Z(n10689) );
  XOR U10609 ( .A(n10718), .B(n10674), .Z(n10677) );
  XNOR U10610 ( .A(n6439), .B(p_input[634]), .Z(n10674) );
  XNOR U10611 ( .A(p_input[2059]), .B(p_input[635]), .Z(n10718) );
  XOR U10612 ( .A(p_input[2060]), .B(p_input[636]), .Z(n10678) );
  XNOR U10613 ( .A(n10688), .B(n10679), .Z(n10717) );
  XNOR U10614 ( .A(n6553), .B(p_input[625]), .Z(n10679) );
  XOR U10615 ( .A(n10719), .B(n10694), .Z(n10688) );
  XNOR U10616 ( .A(p_input[2063]), .B(p_input[639]), .Z(n10694) );
  XOR U10617 ( .A(n10685), .B(n10693), .Z(n10719) );
  XOR U10618 ( .A(n10720), .B(n10690), .Z(n10693) );
  XOR U10619 ( .A(p_input[2061]), .B(p_input[637]), .Z(n10690) );
  XNOR U10620 ( .A(p_input[2062]), .B(p_input[638]), .Z(n10720) );
  XNOR U10621 ( .A(n6325), .B(p_input[633]), .Z(n10685) );
  XNOR U10622 ( .A(n10701), .B(n10700), .Z(n10683) );
  XNOR U10623 ( .A(n10721), .B(n10706), .Z(n10700) );
  XOR U10624 ( .A(p_input[2056]), .B(p_input[632]), .Z(n10706) );
  XOR U10625 ( .A(n10697), .B(n10705), .Z(n10721) );
  XOR U10626 ( .A(n10722), .B(n10702), .Z(n10705) );
  XOR U10627 ( .A(p_input[2054]), .B(p_input[630]), .Z(n10702) );
  XNOR U10628 ( .A(p_input[2055]), .B(p_input[631]), .Z(n10722) );
  XNOR U10629 ( .A(n6328), .B(p_input[626]), .Z(n10697) );
  XNOR U10630 ( .A(n10711), .B(n10710), .Z(n10701) );
  XOR U10631 ( .A(n10723), .B(n10707), .Z(n10710) );
  XOR U10632 ( .A(p_input[2051]), .B(p_input[627]), .Z(n10707) );
  XNOR U10633 ( .A(p_input[2052]), .B(p_input[628]), .Z(n10723) );
  XOR U10634 ( .A(p_input[2053]), .B(p_input[629]), .Z(n10711) );
  XOR U10635 ( .A(n10724), .B(n10725), .Z(n10612) );
  AND U10636 ( .A(n163), .B(n10726), .Z(n10725) );
  XNOR U10637 ( .A(n10727), .B(n10724), .Z(n10726) );
  XNOR U10638 ( .A(n10728), .B(n10729), .Z(n163) );
  AND U10639 ( .A(n10730), .B(n10731), .Z(n10729) );
  XOR U10640 ( .A(n10625), .B(n10728), .Z(n10731) );
  AND U10641 ( .A(n10732), .B(n10733), .Z(n10625) );
  XNOR U10642 ( .A(n10622), .B(n10728), .Z(n10730) );
  XOR U10643 ( .A(n10734), .B(n10735), .Z(n10622) );
  AND U10644 ( .A(n167), .B(n10736), .Z(n10735) );
  XOR U10645 ( .A(n10737), .B(n10734), .Z(n10736) );
  XOR U10646 ( .A(n10738), .B(n10739), .Z(n10728) );
  AND U10647 ( .A(n10740), .B(n10741), .Z(n10739) );
  XNOR U10648 ( .A(n10738), .B(n10732), .Z(n10741) );
  IV U10649 ( .A(n10640), .Z(n10732) );
  XOR U10650 ( .A(n10742), .B(n10743), .Z(n10640) );
  XOR U10651 ( .A(n10744), .B(n10733), .Z(n10743) );
  AND U10652 ( .A(n10667), .B(n10745), .Z(n10733) );
  AND U10653 ( .A(n10746), .B(n10747), .Z(n10744) );
  XOR U10654 ( .A(n10748), .B(n10742), .Z(n10746) );
  XNOR U10655 ( .A(n10637), .B(n10738), .Z(n10740) );
  XOR U10656 ( .A(n10749), .B(n10750), .Z(n10637) );
  AND U10657 ( .A(n167), .B(n10751), .Z(n10750) );
  XOR U10658 ( .A(n10752), .B(n10749), .Z(n10751) );
  XOR U10659 ( .A(n10753), .B(n10754), .Z(n10738) );
  AND U10660 ( .A(n10755), .B(n10756), .Z(n10754) );
  XNOR U10661 ( .A(n10753), .B(n10667), .Z(n10756) );
  XOR U10662 ( .A(n10757), .B(n10747), .Z(n10667) );
  XNOR U10663 ( .A(n10758), .B(n10742), .Z(n10747) );
  XOR U10664 ( .A(n10759), .B(n10760), .Z(n10742) );
  AND U10665 ( .A(n10761), .B(n10762), .Z(n10760) );
  XOR U10666 ( .A(n10763), .B(n10759), .Z(n10761) );
  XNOR U10667 ( .A(n10764), .B(n10765), .Z(n10758) );
  AND U10668 ( .A(n10766), .B(n10767), .Z(n10765) );
  XOR U10669 ( .A(n10764), .B(n10768), .Z(n10766) );
  XNOR U10670 ( .A(n10748), .B(n10745), .Z(n10757) );
  AND U10671 ( .A(n10769), .B(n10770), .Z(n10745) );
  XOR U10672 ( .A(n10771), .B(n10772), .Z(n10748) );
  AND U10673 ( .A(n10773), .B(n10774), .Z(n10772) );
  XOR U10674 ( .A(n10771), .B(n10775), .Z(n10773) );
  XNOR U10675 ( .A(n10664), .B(n10753), .Z(n10755) );
  XOR U10676 ( .A(n10776), .B(n10777), .Z(n10664) );
  AND U10677 ( .A(n167), .B(n10778), .Z(n10777) );
  XNOR U10678 ( .A(n10779), .B(n10776), .Z(n10778) );
  XOR U10679 ( .A(n10780), .B(n10781), .Z(n10753) );
  AND U10680 ( .A(n10782), .B(n10783), .Z(n10781) );
  XNOR U10681 ( .A(n10780), .B(n10769), .Z(n10783) );
  IV U10682 ( .A(n10715), .Z(n10769) );
  XNOR U10683 ( .A(n10784), .B(n10762), .Z(n10715) );
  XNOR U10684 ( .A(n10785), .B(n10768), .Z(n10762) );
  XOR U10685 ( .A(n10786), .B(n10787), .Z(n10768) );
  NOR U10686 ( .A(n10788), .B(n10789), .Z(n10787) );
  XNOR U10687 ( .A(n10786), .B(n10790), .Z(n10788) );
  XNOR U10688 ( .A(n10767), .B(n10759), .Z(n10785) );
  XOR U10689 ( .A(n10791), .B(n10792), .Z(n10759) );
  AND U10690 ( .A(n10793), .B(n10794), .Z(n10792) );
  XNOR U10691 ( .A(n10791), .B(n10795), .Z(n10793) );
  XNOR U10692 ( .A(n10796), .B(n10764), .Z(n10767) );
  XOR U10693 ( .A(n10797), .B(n10798), .Z(n10764) );
  AND U10694 ( .A(n10799), .B(n10800), .Z(n10798) );
  XOR U10695 ( .A(n10797), .B(n10801), .Z(n10799) );
  XNOR U10696 ( .A(n10802), .B(n10803), .Z(n10796) );
  NOR U10697 ( .A(n10804), .B(n10805), .Z(n10803) );
  XOR U10698 ( .A(n10802), .B(n10806), .Z(n10804) );
  XNOR U10699 ( .A(n10763), .B(n10770), .Z(n10784) );
  NOR U10700 ( .A(n10727), .B(n10807), .Z(n10770) );
  XOR U10701 ( .A(n10775), .B(n10774), .Z(n10763) );
  XNOR U10702 ( .A(n10808), .B(n10771), .Z(n10774) );
  XOR U10703 ( .A(n10809), .B(n10810), .Z(n10771) );
  AND U10704 ( .A(n10811), .B(n10812), .Z(n10810) );
  XOR U10705 ( .A(n10809), .B(n10813), .Z(n10811) );
  XNOR U10706 ( .A(n10814), .B(n10815), .Z(n10808) );
  NOR U10707 ( .A(n10816), .B(n10817), .Z(n10815) );
  XNOR U10708 ( .A(n10814), .B(n10818), .Z(n10816) );
  XOR U10709 ( .A(n10819), .B(n10820), .Z(n10775) );
  NOR U10710 ( .A(n10821), .B(n10822), .Z(n10820) );
  XNOR U10711 ( .A(n10819), .B(n10823), .Z(n10821) );
  XNOR U10712 ( .A(n10712), .B(n10780), .Z(n10782) );
  XOR U10713 ( .A(n10824), .B(n10825), .Z(n10712) );
  AND U10714 ( .A(n167), .B(n10826), .Z(n10825) );
  XOR U10715 ( .A(n10827), .B(n10824), .Z(n10826) );
  AND U10716 ( .A(n10724), .B(n10727), .Z(n10780) );
  XOR U10717 ( .A(n10828), .B(n10807), .Z(n10727) );
  XNOR U10718 ( .A(p_input[2048]), .B(p_input[640]), .Z(n10807) );
  XOR U10719 ( .A(n10795), .B(n10794), .Z(n10828) );
  XNOR U10720 ( .A(n10829), .B(n10801), .Z(n10794) );
  XNOR U10721 ( .A(n10790), .B(n10789), .Z(n10801) );
  XOR U10722 ( .A(n10830), .B(n10786), .Z(n10789) );
  XNOR U10723 ( .A(n6439), .B(p_input[650]), .Z(n10786) );
  XNOR U10724 ( .A(p_input[2059]), .B(p_input[651]), .Z(n10830) );
  XOR U10725 ( .A(p_input[2060]), .B(p_input[652]), .Z(n10790) );
  XNOR U10726 ( .A(n10800), .B(n10791), .Z(n10829) );
  XNOR U10727 ( .A(n6553), .B(p_input[641]), .Z(n10791) );
  XOR U10728 ( .A(n10831), .B(n10806), .Z(n10800) );
  XNOR U10729 ( .A(p_input[2063]), .B(p_input[655]), .Z(n10806) );
  XOR U10730 ( .A(n10797), .B(n10805), .Z(n10831) );
  XOR U10731 ( .A(n10832), .B(n10802), .Z(n10805) );
  XOR U10732 ( .A(p_input[2061]), .B(p_input[653]), .Z(n10802) );
  XNOR U10733 ( .A(p_input[2062]), .B(p_input[654]), .Z(n10832) );
  XNOR U10734 ( .A(n6325), .B(p_input[649]), .Z(n10797) );
  XNOR U10735 ( .A(n10813), .B(n10812), .Z(n10795) );
  XNOR U10736 ( .A(n10833), .B(n10818), .Z(n10812) );
  XOR U10737 ( .A(p_input[2056]), .B(p_input[648]), .Z(n10818) );
  XOR U10738 ( .A(n10809), .B(n10817), .Z(n10833) );
  XOR U10739 ( .A(n10834), .B(n10814), .Z(n10817) );
  XOR U10740 ( .A(p_input[2054]), .B(p_input[646]), .Z(n10814) );
  XNOR U10741 ( .A(p_input[2055]), .B(p_input[647]), .Z(n10834) );
  XNOR U10742 ( .A(n6328), .B(p_input[642]), .Z(n10809) );
  XNOR U10743 ( .A(n10823), .B(n10822), .Z(n10813) );
  XOR U10744 ( .A(n10835), .B(n10819), .Z(n10822) );
  XOR U10745 ( .A(p_input[2051]), .B(p_input[643]), .Z(n10819) );
  XNOR U10746 ( .A(p_input[2052]), .B(p_input[644]), .Z(n10835) );
  XOR U10747 ( .A(p_input[2053]), .B(p_input[645]), .Z(n10823) );
  XOR U10748 ( .A(n10836), .B(n10837), .Z(n10724) );
  AND U10749 ( .A(n167), .B(n10838), .Z(n10837) );
  XNOR U10750 ( .A(n10839), .B(n10836), .Z(n10838) );
  XNOR U10751 ( .A(n10840), .B(n10841), .Z(n167) );
  AND U10752 ( .A(n10842), .B(n10843), .Z(n10841) );
  XOR U10753 ( .A(n10737), .B(n10840), .Z(n10843) );
  AND U10754 ( .A(n10844), .B(n10845), .Z(n10737) );
  XNOR U10755 ( .A(n10734), .B(n10840), .Z(n10842) );
  XOR U10756 ( .A(n10846), .B(n10847), .Z(n10734) );
  AND U10757 ( .A(n171), .B(n10848), .Z(n10847) );
  XOR U10758 ( .A(n10849), .B(n10846), .Z(n10848) );
  XOR U10759 ( .A(n10850), .B(n10851), .Z(n10840) );
  AND U10760 ( .A(n10852), .B(n10853), .Z(n10851) );
  XNOR U10761 ( .A(n10850), .B(n10844), .Z(n10853) );
  IV U10762 ( .A(n10752), .Z(n10844) );
  XOR U10763 ( .A(n10854), .B(n10855), .Z(n10752) );
  XOR U10764 ( .A(n10856), .B(n10845), .Z(n10855) );
  AND U10765 ( .A(n10779), .B(n10857), .Z(n10845) );
  AND U10766 ( .A(n10858), .B(n10859), .Z(n10856) );
  XOR U10767 ( .A(n10860), .B(n10854), .Z(n10858) );
  XNOR U10768 ( .A(n10749), .B(n10850), .Z(n10852) );
  XOR U10769 ( .A(n10861), .B(n10862), .Z(n10749) );
  AND U10770 ( .A(n171), .B(n10863), .Z(n10862) );
  XOR U10771 ( .A(n10864), .B(n10861), .Z(n10863) );
  XOR U10772 ( .A(n10865), .B(n10866), .Z(n10850) );
  AND U10773 ( .A(n10867), .B(n10868), .Z(n10866) );
  XNOR U10774 ( .A(n10865), .B(n10779), .Z(n10868) );
  XOR U10775 ( .A(n10869), .B(n10859), .Z(n10779) );
  XNOR U10776 ( .A(n10870), .B(n10854), .Z(n10859) );
  XOR U10777 ( .A(n10871), .B(n10872), .Z(n10854) );
  AND U10778 ( .A(n10873), .B(n10874), .Z(n10872) );
  XOR U10779 ( .A(n10875), .B(n10871), .Z(n10873) );
  XNOR U10780 ( .A(n10876), .B(n10877), .Z(n10870) );
  AND U10781 ( .A(n10878), .B(n10879), .Z(n10877) );
  XOR U10782 ( .A(n10876), .B(n10880), .Z(n10878) );
  XNOR U10783 ( .A(n10860), .B(n10857), .Z(n10869) );
  AND U10784 ( .A(n10881), .B(n10882), .Z(n10857) );
  XOR U10785 ( .A(n10883), .B(n10884), .Z(n10860) );
  AND U10786 ( .A(n10885), .B(n10886), .Z(n10884) );
  XOR U10787 ( .A(n10883), .B(n10887), .Z(n10885) );
  XNOR U10788 ( .A(n10776), .B(n10865), .Z(n10867) );
  XOR U10789 ( .A(n10888), .B(n10889), .Z(n10776) );
  AND U10790 ( .A(n171), .B(n10890), .Z(n10889) );
  XNOR U10791 ( .A(n10891), .B(n10888), .Z(n10890) );
  XOR U10792 ( .A(n10892), .B(n10893), .Z(n10865) );
  AND U10793 ( .A(n10894), .B(n10895), .Z(n10893) );
  XNOR U10794 ( .A(n10892), .B(n10881), .Z(n10895) );
  IV U10795 ( .A(n10827), .Z(n10881) );
  XNOR U10796 ( .A(n10896), .B(n10874), .Z(n10827) );
  XNOR U10797 ( .A(n10897), .B(n10880), .Z(n10874) );
  XOR U10798 ( .A(n10898), .B(n10899), .Z(n10880) );
  NOR U10799 ( .A(n10900), .B(n10901), .Z(n10899) );
  XNOR U10800 ( .A(n10898), .B(n10902), .Z(n10900) );
  XNOR U10801 ( .A(n10879), .B(n10871), .Z(n10897) );
  XOR U10802 ( .A(n10903), .B(n10904), .Z(n10871) );
  AND U10803 ( .A(n10905), .B(n10906), .Z(n10904) );
  XNOR U10804 ( .A(n10903), .B(n10907), .Z(n10905) );
  XNOR U10805 ( .A(n10908), .B(n10876), .Z(n10879) );
  XOR U10806 ( .A(n10909), .B(n10910), .Z(n10876) );
  AND U10807 ( .A(n10911), .B(n10912), .Z(n10910) );
  XOR U10808 ( .A(n10909), .B(n10913), .Z(n10911) );
  XNOR U10809 ( .A(n10914), .B(n10915), .Z(n10908) );
  NOR U10810 ( .A(n10916), .B(n10917), .Z(n10915) );
  XOR U10811 ( .A(n10914), .B(n10918), .Z(n10916) );
  XNOR U10812 ( .A(n10875), .B(n10882), .Z(n10896) );
  NOR U10813 ( .A(n10839), .B(n10919), .Z(n10882) );
  XOR U10814 ( .A(n10887), .B(n10886), .Z(n10875) );
  XNOR U10815 ( .A(n10920), .B(n10883), .Z(n10886) );
  XOR U10816 ( .A(n10921), .B(n10922), .Z(n10883) );
  AND U10817 ( .A(n10923), .B(n10924), .Z(n10922) );
  XOR U10818 ( .A(n10921), .B(n10925), .Z(n10923) );
  XNOR U10819 ( .A(n10926), .B(n10927), .Z(n10920) );
  NOR U10820 ( .A(n10928), .B(n10929), .Z(n10927) );
  XNOR U10821 ( .A(n10926), .B(n10930), .Z(n10928) );
  XOR U10822 ( .A(n10931), .B(n10932), .Z(n10887) );
  NOR U10823 ( .A(n10933), .B(n10934), .Z(n10932) );
  XNOR U10824 ( .A(n10931), .B(n10935), .Z(n10933) );
  XNOR U10825 ( .A(n10824), .B(n10892), .Z(n10894) );
  XOR U10826 ( .A(n10936), .B(n10937), .Z(n10824) );
  AND U10827 ( .A(n171), .B(n10938), .Z(n10937) );
  XOR U10828 ( .A(n10939), .B(n10936), .Z(n10938) );
  AND U10829 ( .A(n10836), .B(n10839), .Z(n10892) );
  XOR U10830 ( .A(n10940), .B(n10919), .Z(n10839) );
  XNOR U10831 ( .A(p_input[2048]), .B(p_input[656]), .Z(n10919) );
  XOR U10832 ( .A(n10907), .B(n10906), .Z(n10940) );
  XNOR U10833 ( .A(n10941), .B(n10913), .Z(n10906) );
  XNOR U10834 ( .A(n10902), .B(n10901), .Z(n10913) );
  XOR U10835 ( .A(n10942), .B(n10898), .Z(n10901) );
  XNOR U10836 ( .A(n6439), .B(p_input[666]), .Z(n10898) );
  XNOR U10837 ( .A(p_input[2059]), .B(p_input[667]), .Z(n10942) );
  XOR U10838 ( .A(p_input[2060]), .B(p_input[668]), .Z(n10902) );
  XNOR U10839 ( .A(n10912), .B(n10903), .Z(n10941) );
  XNOR U10840 ( .A(n6553), .B(p_input[657]), .Z(n10903) );
  XOR U10841 ( .A(n10943), .B(n10918), .Z(n10912) );
  XNOR U10842 ( .A(p_input[2063]), .B(p_input[671]), .Z(n10918) );
  XOR U10843 ( .A(n10909), .B(n10917), .Z(n10943) );
  XOR U10844 ( .A(n10944), .B(n10914), .Z(n10917) );
  XOR U10845 ( .A(p_input[2061]), .B(p_input[669]), .Z(n10914) );
  XNOR U10846 ( .A(p_input[2062]), .B(p_input[670]), .Z(n10944) );
  XNOR U10847 ( .A(n6325), .B(p_input[665]), .Z(n10909) );
  XNOR U10848 ( .A(n10925), .B(n10924), .Z(n10907) );
  XNOR U10849 ( .A(n10945), .B(n10930), .Z(n10924) );
  XOR U10850 ( .A(p_input[2056]), .B(p_input[664]), .Z(n10930) );
  XOR U10851 ( .A(n10921), .B(n10929), .Z(n10945) );
  XOR U10852 ( .A(n10946), .B(n10926), .Z(n10929) );
  XOR U10853 ( .A(p_input[2054]), .B(p_input[662]), .Z(n10926) );
  XNOR U10854 ( .A(p_input[2055]), .B(p_input[663]), .Z(n10946) );
  XNOR U10855 ( .A(n6328), .B(p_input[658]), .Z(n10921) );
  XNOR U10856 ( .A(n10935), .B(n10934), .Z(n10925) );
  XOR U10857 ( .A(n10947), .B(n10931), .Z(n10934) );
  XOR U10858 ( .A(p_input[2051]), .B(p_input[659]), .Z(n10931) );
  XNOR U10859 ( .A(p_input[2052]), .B(p_input[660]), .Z(n10947) );
  XOR U10860 ( .A(p_input[2053]), .B(p_input[661]), .Z(n10935) );
  XOR U10861 ( .A(n10948), .B(n10949), .Z(n10836) );
  AND U10862 ( .A(n171), .B(n10950), .Z(n10949) );
  XNOR U10863 ( .A(n10951), .B(n10948), .Z(n10950) );
  XNOR U10864 ( .A(n10952), .B(n10953), .Z(n171) );
  AND U10865 ( .A(n10954), .B(n10955), .Z(n10953) );
  XOR U10866 ( .A(n10849), .B(n10952), .Z(n10955) );
  AND U10867 ( .A(n10956), .B(n10957), .Z(n10849) );
  XNOR U10868 ( .A(n10846), .B(n10952), .Z(n10954) );
  XOR U10869 ( .A(n10958), .B(n10959), .Z(n10846) );
  AND U10870 ( .A(n175), .B(n10960), .Z(n10959) );
  XOR U10871 ( .A(n10961), .B(n10958), .Z(n10960) );
  XOR U10872 ( .A(n10962), .B(n10963), .Z(n10952) );
  AND U10873 ( .A(n10964), .B(n10965), .Z(n10963) );
  XNOR U10874 ( .A(n10962), .B(n10956), .Z(n10965) );
  IV U10875 ( .A(n10864), .Z(n10956) );
  XOR U10876 ( .A(n10966), .B(n10967), .Z(n10864) );
  XOR U10877 ( .A(n10968), .B(n10957), .Z(n10967) );
  AND U10878 ( .A(n10891), .B(n10969), .Z(n10957) );
  AND U10879 ( .A(n10970), .B(n10971), .Z(n10968) );
  XOR U10880 ( .A(n10972), .B(n10966), .Z(n10970) );
  XNOR U10881 ( .A(n10861), .B(n10962), .Z(n10964) );
  XOR U10882 ( .A(n10973), .B(n10974), .Z(n10861) );
  AND U10883 ( .A(n175), .B(n10975), .Z(n10974) );
  XOR U10884 ( .A(n10976), .B(n10973), .Z(n10975) );
  XOR U10885 ( .A(n10977), .B(n10978), .Z(n10962) );
  AND U10886 ( .A(n10979), .B(n10980), .Z(n10978) );
  XNOR U10887 ( .A(n10977), .B(n10891), .Z(n10980) );
  XOR U10888 ( .A(n10981), .B(n10971), .Z(n10891) );
  XNOR U10889 ( .A(n10982), .B(n10966), .Z(n10971) );
  XOR U10890 ( .A(n10983), .B(n10984), .Z(n10966) );
  AND U10891 ( .A(n10985), .B(n10986), .Z(n10984) );
  XOR U10892 ( .A(n10987), .B(n10983), .Z(n10985) );
  XNOR U10893 ( .A(n10988), .B(n10989), .Z(n10982) );
  AND U10894 ( .A(n10990), .B(n10991), .Z(n10989) );
  XOR U10895 ( .A(n10988), .B(n10992), .Z(n10990) );
  XNOR U10896 ( .A(n10972), .B(n10969), .Z(n10981) );
  AND U10897 ( .A(n10993), .B(n10994), .Z(n10969) );
  XOR U10898 ( .A(n10995), .B(n10996), .Z(n10972) );
  AND U10899 ( .A(n10997), .B(n10998), .Z(n10996) );
  XOR U10900 ( .A(n10995), .B(n10999), .Z(n10997) );
  XNOR U10901 ( .A(n10888), .B(n10977), .Z(n10979) );
  XOR U10902 ( .A(n11000), .B(n11001), .Z(n10888) );
  AND U10903 ( .A(n175), .B(n11002), .Z(n11001) );
  XNOR U10904 ( .A(n11003), .B(n11000), .Z(n11002) );
  XOR U10905 ( .A(n11004), .B(n11005), .Z(n10977) );
  AND U10906 ( .A(n11006), .B(n11007), .Z(n11005) );
  XNOR U10907 ( .A(n11004), .B(n10993), .Z(n11007) );
  IV U10908 ( .A(n10939), .Z(n10993) );
  XNOR U10909 ( .A(n11008), .B(n10986), .Z(n10939) );
  XNOR U10910 ( .A(n11009), .B(n10992), .Z(n10986) );
  XOR U10911 ( .A(n11010), .B(n11011), .Z(n10992) );
  NOR U10912 ( .A(n11012), .B(n11013), .Z(n11011) );
  XNOR U10913 ( .A(n11010), .B(n11014), .Z(n11012) );
  XNOR U10914 ( .A(n10991), .B(n10983), .Z(n11009) );
  XOR U10915 ( .A(n11015), .B(n11016), .Z(n10983) );
  AND U10916 ( .A(n11017), .B(n11018), .Z(n11016) );
  XNOR U10917 ( .A(n11015), .B(n11019), .Z(n11017) );
  XNOR U10918 ( .A(n11020), .B(n10988), .Z(n10991) );
  XOR U10919 ( .A(n11021), .B(n11022), .Z(n10988) );
  AND U10920 ( .A(n11023), .B(n11024), .Z(n11022) );
  XOR U10921 ( .A(n11021), .B(n11025), .Z(n11023) );
  XNOR U10922 ( .A(n11026), .B(n11027), .Z(n11020) );
  NOR U10923 ( .A(n11028), .B(n11029), .Z(n11027) );
  XOR U10924 ( .A(n11026), .B(n11030), .Z(n11028) );
  XNOR U10925 ( .A(n10987), .B(n10994), .Z(n11008) );
  NOR U10926 ( .A(n10951), .B(n11031), .Z(n10994) );
  XOR U10927 ( .A(n10999), .B(n10998), .Z(n10987) );
  XNOR U10928 ( .A(n11032), .B(n10995), .Z(n10998) );
  XOR U10929 ( .A(n11033), .B(n11034), .Z(n10995) );
  AND U10930 ( .A(n11035), .B(n11036), .Z(n11034) );
  XOR U10931 ( .A(n11033), .B(n11037), .Z(n11035) );
  XNOR U10932 ( .A(n11038), .B(n11039), .Z(n11032) );
  NOR U10933 ( .A(n11040), .B(n11041), .Z(n11039) );
  XNOR U10934 ( .A(n11038), .B(n11042), .Z(n11040) );
  XOR U10935 ( .A(n11043), .B(n11044), .Z(n10999) );
  NOR U10936 ( .A(n11045), .B(n11046), .Z(n11044) );
  XNOR U10937 ( .A(n11043), .B(n11047), .Z(n11045) );
  XNOR U10938 ( .A(n10936), .B(n11004), .Z(n11006) );
  XOR U10939 ( .A(n11048), .B(n11049), .Z(n10936) );
  AND U10940 ( .A(n175), .B(n11050), .Z(n11049) );
  XOR U10941 ( .A(n11051), .B(n11048), .Z(n11050) );
  AND U10942 ( .A(n10948), .B(n10951), .Z(n11004) );
  XOR U10943 ( .A(n11052), .B(n11031), .Z(n10951) );
  XNOR U10944 ( .A(p_input[2048]), .B(p_input[672]), .Z(n11031) );
  XOR U10945 ( .A(n11019), .B(n11018), .Z(n11052) );
  XNOR U10946 ( .A(n11053), .B(n11025), .Z(n11018) );
  XNOR U10947 ( .A(n11014), .B(n11013), .Z(n11025) );
  XOR U10948 ( .A(n11054), .B(n11010), .Z(n11013) );
  XNOR U10949 ( .A(n6439), .B(p_input[682]), .Z(n11010) );
  XNOR U10950 ( .A(p_input[2059]), .B(p_input[683]), .Z(n11054) );
  XOR U10951 ( .A(p_input[2060]), .B(p_input[684]), .Z(n11014) );
  XNOR U10952 ( .A(n11024), .B(n11015), .Z(n11053) );
  XNOR U10953 ( .A(n6553), .B(p_input[673]), .Z(n11015) );
  XOR U10954 ( .A(n11055), .B(n11030), .Z(n11024) );
  XNOR U10955 ( .A(p_input[2063]), .B(p_input[687]), .Z(n11030) );
  XOR U10956 ( .A(n11021), .B(n11029), .Z(n11055) );
  XOR U10957 ( .A(n11056), .B(n11026), .Z(n11029) );
  XOR U10958 ( .A(p_input[2061]), .B(p_input[685]), .Z(n11026) );
  XNOR U10959 ( .A(p_input[2062]), .B(p_input[686]), .Z(n11056) );
  XNOR U10960 ( .A(n6325), .B(p_input[681]), .Z(n11021) );
  XNOR U10961 ( .A(n11037), .B(n11036), .Z(n11019) );
  XNOR U10962 ( .A(n11057), .B(n11042), .Z(n11036) );
  XOR U10963 ( .A(p_input[2056]), .B(p_input[680]), .Z(n11042) );
  XOR U10964 ( .A(n11033), .B(n11041), .Z(n11057) );
  XOR U10965 ( .A(n11058), .B(n11038), .Z(n11041) );
  XOR U10966 ( .A(p_input[2054]), .B(p_input[678]), .Z(n11038) );
  XNOR U10967 ( .A(p_input[2055]), .B(p_input[679]), .Z(n11058) );
  XNOR U10968 ( .A(n6328), .B(p_input[674]), .Z(n11033) );
  XNOR U10969 ( .A(n11047), .B(n11046), .Z(n11037) );
  XOR U10970 ( .A(n11059), .B(n11043), .Z(n11046) );
  XOR U10971 ( .A(p_input[2051]), .B(p_input[675]), .Z(n11043) );
  XNOR U10972 ( .A(p_input[2052]), .B(p_input[676]), .Z(n11059) );
  XOR U10973 ( .A(p_input[2053]), .B(p_input[677]), .Z(n11047) );
  XOR U10974 ( .A(n11060), .B(n11061), .Z(n10948) );
  AND U10975 ( .A(n175), .B(n11062), .Z(n11061) );
  XNOR U10976 ( .A(n11063), .B(n11060), .Z(n11062) );
  XNOR U10977 ( .A(n11064), .B(n11065), .Z(n175) );
  AND U10978 ( .A(n11066), .B(n11067), .Z(n11065) );
  XOR U10979 ( .A(n10961), .B(n11064), .Z(n11067) );
  AND U10980 ( .A(n11068), .B(n11069), .Z(n10961) );
  XNOR U10981 ( .A(n10958), .B(n11064), .Z(n11066) );
  XOR U10982 ( .A(n11070), .B(n11071), .Z(n10958) );
  AND U10983 ( .A(n179), .B(n11072), .Z(n11071) );
  XOR U10984 ( .A(n11073), .B(n11070), .Z(n11072) );
  XOR U10985 ( .A(n11074), .B(n11075), .Z(n11064) );
  AND U10986 ( .A(n11076), .B(n11077), .Z(n11075) );
  XNOR U10987 ( .A(n11074), .B(n11068), .Z(n11077) );
  IV U10988 ( .A(n10976), .Z(n11068) );
  XOR U10989 ( .A(n11078), .B(n11079), .Z(n10976) );
  XOR U10990 ( .A(n11080), .B(n11069), .Z(n11079) );
  AND U10991 ( .A(n11003), .B(n11081), .Z(n11069) );
  AND U10992 ( .A(n11082), .B(n11083), .Z(n11080) );
  XOR U10993 ( .A(n11084), .B(n11078), .Z(n11082) );
  XNOR U10994 ( .A(n10973), .B(n11074), .Z(n11076) );
  XOR U10995 ( .A(n11085), .B(n11086), .Z(n10973) );
  AND U10996 ( .A(n179), .B(n11087), .Z(n11086) );
  XOR U10997 ( .A(n11088), .B(n11085), .Z(n11087) );
  XOR U10998 ( .A(n11089), .B(n11090), .Z(n11074) );
  AND U10999 ( .A(n11091), .B(n11092), .Z(n11090) );
  XNOR U11000 ( .A(n11089), .B(n11003), .Z(n11092) );
  XOR U11001 ( .A(n11093), .B(n11083), .Z(n11003) );
  XNOR U11002 ( .A(n11094), .B(n11078), .Z(n11083) );
  XOR U11003 ( .A(n11095), .B(n11096), .Z(n11078) );
  AND U11004 ( .A(n11097), .B(n11098), .Z(n11096) );
  XOR U11005 ( .A(n11099), .B(n11095), .Z(n11097) );
  XNOR U11006 ( .A(n11100), .B(n11101), .Z(n11094) );
  AND U11007 ( .A(n11102), .B(n11103), .Z(n11101) );
  XOR U11008 ( .A(n11100), .B(n11104), .Z(n11102) );
  XNOR U11009 ( .A(n11084), .B(n11081), .Z(n11093) );
  AND U11010 ( .A(n11105), .B(n11106), .Z(n11081) );
  XOR U11011 ( .A(n11107), .B(n11108), .Z(n11084) );
  AND U11012 ( .A(n11109), .B(n11110), .Z(n11108) );
  XOR U11013 ( .A(n11107), .B(n11111), .Z(n11109) );
  XNOR U11014 ( .A(n11000), .B(n11089), .Z(n11091) );
  XOR U11015 ( .A(n11112), .B(n11113), .Z(n11000) );
  AND U11016 ( .A(n179), .B(n11114), .Z(n11113) );
  XNOR U11017 ( .A(n11115), .B(n11112), .Z(n11114) );
  XOR U11018 ( .A(n11116), .B(n11117), .Z(n11089) );
  AND U11019 ( .A(n11118), .B(n11119), .Z(n11117) );
  XNOR U11020 ( .A(n11116), .B(n11105), .Z(n11119) );
  IV U11021 ( .A(n11051), .Z(n11105) );
  XNOR U11022 ( .A(n11120), .B(n11098), .Z(n11051) );
  XNOR U11023 ( .A(n11121), .B(n11104), .Z(n11098) );
  XOR U11024 ( .A(n11122), .B(n11123), .Z(n11104) );
  NOR U11025 ( .A(n11124), .B(n11125), .Z(n11123) );
  XNOR U11026 ( .A(n11122), .B(n11126), .Z(n11124) );
  XNOR U11027 ( .A(n11103), .B(n11095), .Z(n11121) );
  XOR U11028 ( .A(n11127), .B(n11128), .Z(n11095) );
  AND U11029 ( .A(n11129), .B(n11130), .Z(n11128) );
  XNOR U11030 ( .A(n11127), .B(n11131), .Z(n11129) );
  XNOR U11031 ( .A(n11132), .B(n11100), .Z(n11103) );
  XOR U11032 ( .A(n11133), .B(n11134), .Z(n11100) );
  AND U11033 ( .A(n11135), .B(n11136), .Z(n11134) );
  XOR U11034 ( .A(n11133), .B(n11137), .Z(n11135) );
  XNOR U11035 ( .A(n11138), .B(n11139), .Z(n11132) );
  NOR U11036 ( .A(n11140), .B(n11141), .Z(n11139) );
  XOR U11037 ( .A(n11138), .B(n11142), .Z(n11140) );
  XNOR U11038 ( .A(n11099), .B(n11106), .Z(n11120) );
  NOR U11039 ( .A(n11063), .B(n11143), .Z(n11106) );
  XOR U11040 ( .A(n11111), .B(n11110), .Z(n11099) );
  XNOR U11041 ( .A(n11144), .B(n11107), .Z(n11110) );
  XOR U11042 ( .A(n11145), .B(n11146), .Z(n11107) );
  AND U11043 ( .A(n11147), .B(n11148), .Z(n11146) );
  XOR U11044 ( .A(n11145), .B(n11149), .Z(n11147) );
  XNOR U11045 ( .A(n11150), .B(n11151), .Z(n11144) );
  NOR U11046 ( .A(n11152), .B(n11153), .Z(n11151) );
  XNOR U11047 ( .A(n11150), .B(n11154), .Z(n11152) );
  XOR U11048 ( .A(n11155), .B(n11156), .Z(n11111) );
  NOR U11049 ( .A(n11157), .B(n11158), .Z(n11156) );
  XNOR U11050 ( .A(n11155), .B(n11159), .Z(n11157) );
  XNOR U11051 ( .A(n11048), .B(n11116), .Z(n11118) );
  XOR U11052 ( .A(n11160), .B(n11161), .Z(n11048) );
  AND U11053 ( .A(n179), .B(n11162), .Z(n11161) );
  XOR U11054 ( .A(n11163), .B(n11160), .Z(n11162) );
  AND U11055 ( .A(n11060), .B(n11063), .Z(n11116) );
  XOR U11056 ( .A(n11164), .B(n11143), .Z(n11063) );
  XNOR U11057 ( .A(p_input[2048]), .B(p_input[688]), .Z(n11143) );
  XOR U11058 ( .A(n11131), .B(n11130), .Z(n11164) );
  XNOR U11059 ( .A(n11165), .B(n11137), .Z(n11130) );
  XNOR U11060 ( .A(n11126), .B(n11125), .Z(n11137) );
  XOR U11061 ( .A(n11166), .B(n11122), .Z(n11125) );
  XNOR U11062 ( .A(n6439), .B(p_input[698]), .Z(n11122) );
  XNOR U11063 ( .A(p_input[2059]), .B(p_input[699]), .Z(n11166) );
  XOR U11064 ( .A(p_input[2060]), .B(p_input[700]), .Z(n11126) );
  XNOR U11065 ( .A(n11136), .B(n11127), .Z(n11165) );
  XNOR U11066 ( .A(n6553), .B(p_input[689]), .Z(n11127) );
  XOR U11067 ( .A(n11167), .B(n11142), .Z(n11136) );
  XNOR U11068 ( .A(p_input[2063]), .B(p_input[703]), .Z(n11142) );
  XOR U11069 ( .A(n11133), .B(n11141), .Z(n11167) );
  XOR U11070 ( .A(n11168), .B(n11138), .Z(n11141) );
  XOR U11071 ( .A(p_input[2061]), .B(p_input[701]), .Z(n11138) );
  XNOR U11072 ( .A(p_input[2062]), .B(p_input[702]), .Z(n11168) );
  XNOR U11073 ( .A(n6325), .B(p_input[697]), .Z(n11133) );
  XNOR U11074 ( .A(n11149), .B(n11148), .Z(n11131) );
  XNOR U11075 ( .A(n11169), .B(n11154), .Z(n11148) );
  XOR U11076 ( .A(p_input[2056]), .B(p_input[696]), .Z(n11154) );
  XOR U11077 ( .A(n11145), .B(n11153), .Z(n11169) );
  XOR U11078 ( .A(n11170), .B(n11150), .Z(n11153) );
  XOR U11079 ( .A(p_input[2054]), .B(p_input[694]), .Z(n11150) );
  XNOR U11080 ( .A(p_input[2055]), .B(p_input[695]), .Z(n11170) );
  XNOR U11081 ( .A(n6328), .B(p_input[690]), .Z(n11145) );
  XNOR U11082 ( .A(n11159), .B(n11158), .Z(n11149) );
  XOR U11083 ( .A(n11171), .B(n11155), .Z(n11158) );
  XOR U11084 ( .A(p_input[2051]), .B(p_input[691]), .Z(n11155) );
  XNOR U11085 ( .A(p_input[2052]), .B(p_input[692]), .Z(n11171) );
  XOR U11086 ( .A(p_input[2053]), .B(p_input[693]), .Z(n11159) );
  XOR U11087 ( .A(n11172), .B(n11173), .Z(n11060) );
  AND U11088 ( .A(n179), .B(n11174), .Z(n11173) );
  XNOR U11089 ( .A(n11175), .B(n11172), .Z(n11174) );
  XNOR U11090 ( .A(n11176), .B(n11177), .Z(n179) );
  AND U11091 ( .A(n11178), .B(n11179), .Z(n11177) );
  XOR U11092 ( .A(n11073), .B(n11176), .Z(n11179) );
  AND U11093 ( .A(n11180), .B(n11181), .Z(n11073) );
  XNOR U11094 ( .A(n11070), .B(n11176), .Z(n11178) );
  XOR U11095 ( .A(n11182), .B(n11183), .Z(n11070) );
  AND U11096 ( .A(n183), .B(n11184), .Z(n11183) );
  XOR U11097 ( .A(n11185), .B(n11182), .Z(n11184) );
  XOR U11098 ( .A(n11186), .B(n11187), .Z(n11176) );
  AND U11099 ( .A(n11188), .B(n11189), .Z(n11187) );
  XNOR U11100 ( .A(n11186), .B(n11180), .Z(n11189) );
  IV U11101 ( .A(n11088), .Z(n11180) );
  XOR U11102 ( .A(n11190), .B(n11191), .Z(n11088) );
  XOR U11103 ( .A(n11192), .B(n11181), .Z(n11191) );
  AND U11104 ( .A(n11115), .B(n11193), .Z(n11181) );
  AND U11105 ( .A(n11194), .B(n11195), .Z(n11192) );
  XOR U11106 ( .A(n11196), .B(n11190), .Z(n11194) );
  XNOR U11107 ( .A(n11085), .B(n11186), .Z(n11188) );
  XOR U11108 ( .A(n11197), .B(n11198), .Z(n11085) );
  AND U11109 ( .A(n183), .B(n11199), .Z(n11198) );
  XOR U11110 ( .A(n11200), .B(n11197), .Z(n11199) );
  XOR U11111 ( .A(n11201), .B(n11202), .Z(n11186) );
  AND U11112 ( .A(n11203), .B(n11204), .Z(n11202) );
  XNOR U11113 ( .A(n11201), .B(n11115), .Z(n11204) );
  XOR U11114 ( .A(n11205), .B(n11195), .Z(n11115) );
  XNOR U11115 ( .A(n11206), .B(n11190), .Z(n11195) );
  XOR U11116 ( .A(n11207), .B(n11208), .Z(n11190) );
  AND U11117 ( .A(n11209), .B(n11210), .Z(n11208) );
  XOR U11118 ( .A(n11211), .B(n11207), .Z(n11209) );
  XNOR U11119 ( .A(n11212), .B(n11213), .Z(n11206) );
  AND U11120 ( .A(n11214), .B(n11215), .Z(n11213) );
  XOR U11121 ( .A(n11212), .B(n11216), .Z(n11214) );
  XNOR U11122 ( .A(n11196), .B(n11193), .Z(n11205) );
  AND U11123 ( .A(n11217), .B(n11218), .Z(n11193) );
  XOR U11124 ( .A(n11219), .B(n11220), .Z(n11196) );
  AND U11125 ( .A(n11221), .B(n11222), .Z(n11220) );
  XOR U11126 ( .A(n11219), .B(n11223), .Z(n11221) );
  XNOR U11127 ( .A(n11112), .B(n11201), .Z(n11203) );
  XOR U11128 ( .A(n11224), .B(n11225), .Z(n11112) );
  AND U11129 ( .A(n183), .B(n11226), .Z(n11225) );
  XNOR U11130 ( .A(n11227), .B(n11224), .Z(n11226) );
  XOR U11131 ( .A(n11228), .B(n11229), .Z(n11201) );
  AND U11132 ( .A(n11230), .B(n11231), .Z(n11229) );
  XNOR U11133 ( .A(n11228), .B(n11217), .Z(n11231) );
  IV U11134 ( .A(n11163), .Z(n11217) );
  XNOR U11135 ( .A(n11232), .B(n11210), .Z(n11163) );
  XNOR U11136 ( .A(n11233), .B(n11216), .Z(n11210) );
  XOR U11137 ( .A(n11234), .B(n11235), .Z(n11216) );
  NOR U11138 ( .A(n11236), .B(n11237), .Z(n11235) );
  XNOR U11139 ( .A(n11234), .B(n11238), .Z(n11236) );
  XNOR U11140 ( .A(n11215), .B(n11207), .Z(n11233) );
  XOR U11141 ( .A(n11239), .B(n11240), .Z(n11207) );
  AND U11142 ( .A(n11241), .B(n11242), .Z(n11240) );
  XNOR U11143 ( .A(n11239), .B(n11243), .Z(n11241) );
  XNOR U11144 ( .A(n11244), .B(n11212), .Z(n11215) );
  XOR U11145 ( .A(n11245), .B(n11246), .Z(n11212) );
  AND U11146 ( .A(n11247), .B(n11248), .Z(n11246) );
  XOR U11147 ( .A(n11245), .B(n11249), .Z(n11247) );
  XNOR U11148 ( .A(n11250), .B(n11251), .Z(n11244) );
  NOR U11149 ( .A(n11252), .B(n11253), .Z(n11251) );
  XOR U11150 ( .A(n11250), .B(n11254), .Z(n11252) );
  XNOR U11151 ( .A(n11211), .B(n11218), .Z(n11232) );
  NOR U11152 ( .A(n11175), .B(n11255), .Z(n11218) );
  XOR U11153 ( .A(n11223), .B(n11222), .Z(n11211) );
  XNOR U11154 ( .A(n11256), .B(n11219), .Z(n11222) );
  XOR U11155 ( .A(n11257), .B(n11258), .Z(n11219) );
  AND U11156 ( .A(n11259), .B(n11260), .Z(n11258) );
  XOR U11157 ( .A(n11257), .B(n11261), .Z(n11259) );
  XNOR U11158 ( .A(n11262), .B(n11263), .Z(n11256) );
  NOR U11159 ( .A(n11264), .B(n11265), .Z(n11263) );
  XNOR U11160 ( .A(n11262), .B(n11266), .Z(n11264) );
  XOR U11161 ( .A(n11267), .B(n11268), .Z(n11223) );
  NOR U11162 ( .A(n11269), .B(n11270), .Z(n11268) );
  XNOR U11163 ( .A(n11267), .B(n11271), .Z(n11269) );
  XNOR U11164 ( .A(n11160), .B(n11228), .Z(n11230) );
  XOR U11165 ( .A(n11272), .B(n11273), .Z(n11160) );
  AND U11166 ( .A(n183), .B(n11274), .Z(n11273) );
  XOR U11167 ( .A(n11275), .B(n11272), .Z(n11274) );
  AND U11168 ( .A(n11172), .B(n11175), .Z(n11228) );
  XOR U11169 ( .A(n11276), .B(n11255), .Z(n11175) );
  XNOR U11170 ( .A(p_input[2048]), .B(p_input[704]), .Z(n11255) );
  XOR U11171 ( .A(n11243), .B(n11242), .Z(n11276) );
  XNOR U11172 ( .A(n11277), .B(n11249), .Z(n11242) );
  XNOR U11173 ( .A(n11238), .B(n11237), .Z(n11249) );
  XOR U11174 ( .A(n11278), .B(n11234), .Z(n11237) );
  XNOR U11175 ( .A(n6439), .B(p_input[714]), .Z(n11234) );
  XNOR U11176 ( .A(p_input[2059]), .B(p_input[715]), .Z(n11278) );
  XOR U11177 ( .A(p_input[2060]), .B(p_input[716]), .Z(n11238) );
  XNOR U11178 ( .A(n11248), .B(n11239), .Z(n11277) );
  XNOR U11179 ( .A(n6553), .B(p_input[705]), .Z(n11239) );
  XOR U11180 ( .A(n11279), .B(n11254), .Z(n11248) );
  XNOR U11181 ( .A(p_input[2063]), .B(p_input[719]), .Z(n11254) );
  XOR U11182 ( .A(n11245), .B(n11253), .Z(n11279) );
  XOR U11183 ( .A(n11280), .B(n11250), .Z(n11253) );
  XOR U11184 ( .A(p_input[2061]), .B(p_input[717]), .Z(n11250) );
  XNOR U11185 ( .A(p_input[2062]), .B(p_input[718]), .Z(n11280) );
  XNOR U11186 ( .A(n6325), .B(p_input[713]), .Z(n11245) );
  XNOR U11187 ( .A(n11261), .B(n11260), .Z(n11243) );
  XNOR U11188 ( .A(n11281), .B(n11266), .Z(n11260) );
  XOR U11189 ( .A(p_input[2056]), .B(p_input[712]), .Z(n11266) );
  XOR U11190 ( .A(n11257), .B(n11265), .Z(n11281) );
  XOR U11191 ( .A(n11282), .B(n11262), .Z(n11265) );
  XOR U11192 ( .A(p_input[2054]), .B(p_input[710]), .Z(n11262) );
  XNOR U11193 ( .A(p_input[2055]), .B(p_input[711]), .Z(n11282) );
  XNOR U11194 ( .A(n6328), .B(p_input[706]), .Z(n11257) );
  XNOR U11195 ( .A(n11271), .B(n11270), .Z(n11261) );
  XOR U11196 ( .A(n11283), .B(n11267), .Z(n11270) );
  XOR U11197 ( .A(p_input[2051]), .B(p_input[707]), .Z(n11267) );
  XNOR U11198 ( .A(p_input[2052]), .B(p_input[708]), .Z(n11283) );
  XOR U11199 ( .A(p_input[2053]), .B(p_input[709]), .Z(n11271) );
  XOR U11200 ( .A(n11284), .B(n11285), .Z(n11172) );
  AND U11201 ( .A(n183), .B(n11286), .Z(n11285) );
  XNOR U11202 ( .A(n11287), .B(n11284), .Z(n11286) );
  XNOR U11203 ( .A(n11288), .B(n11289), .Z(n183) );
  AND U11204 ( .A(n11290), .B(n11291), .Z(n11289) );
  XOR U11205 ( .A(n11185), .B(n11288), .Z(n11291) );
  AND U11206 ( .A(n11292), .B(n11293), .Z(n11185) );
  XNOR U11207 ( .A(n11182), .B(n11288), .Z(n11290) );
  XOR U11208 ( .A(n11294), .B(n11295), .Z(n11182) );
  AND U11209 ( .A(n187), .B(n11296), .Z(n11295) );
  XOR U11210 ( .A(n11297), .B(n11294), .Z(n11296) );
  XOR U11211 ( .A(n11298), .B(n11299), .Z(n11288) );
  AND U11212 ( .A(n11300), .B(n11301), .Z(n11299) );
  XNOR U11213 ( .A(n11298), .B(n11292), .Z(n11301) );
  IV U11214 ( .A(n11200), .Z(n11292) );
  XOR U11215 ( .A(n11302), .B(n11303), .Z(n11200) );
  XOR U11216 ( .A(n11304), .B(n11293), .Z(n11303) );
  AND U11217 ( .A(n11227), .B(n11305), .Z(n11293) );
  AND U11218 ( .A(n11306), .B(n11307), .Z(n11304) );
  XOR U11219 ( .A(n11308), .B(n11302), .Z(n11306) );
  XNOR U11220 ( .A(n11197), .B(n11298), .Z(n11300) );
  XOR U11221 ( .A(n11309), .B(n11310), .Z(n11197) );
  AND U11222 ( .A(n187), .B(n11311), .Z(n11310) );
  XOR U11223 ( .A(n11312), .B(n11309), .Z(n11311) );
  XOR U11224 ( .A(n11313), .B(n11314), .Z(n11298) );
  AND U11225 ( .A(n11315), .B(n11316), .Z(n11314) );
  XNOR U11226 ( .A(n11313), .B(n11227), .Z(n11316) );
  XOR U11227 ( .A(n11317), .B(n11307), .Z(n11227) );
  XNOR U11228 ( .A(n11318), .B(n11302), .Z(n11307) );
  XOR U11229 ( .A(n11319), .B(n11320), .Z(n11302) );
  AND U11230 ( .A(n11321), .B(n11322), .Z(n11320) );
  XOR U11231 ( .A(n11323), .B(n11319), .Z(n11321) );
  XNOR U11232 ( .A(n11324), .B(n11325), .Z(n11318) );
  AND U11233 ( .A(n11326), .B(n11327), .Z(n11325) );
  XOR U11234 ( .A(n11324), .B(n11328), .Z(n11326) );
  XNOR U11235 ( .A(n11308), .B(n11305), .Z(n11317) );
  AND U11236 ( .A(n11329), .B(n11330), .Z(n11305) );
  XOR U11237 ( .A(n11331), .B(n11332), .Z(n11308) );
  AND U11238 ( .A(n11333), .B(n11334), .Z(n11332) );
  XOR U11239 ( .A(n11331), .B(n11335), .Z(n11333) );
  XNOR U11240 ( .A(n11224), .B(n11313), .Z(n11315) );
  XOR U11241 ( .A(n11336), .B(n11337), .Z(n11224) );
  AND U11242 ( .A(n187), .B(n11338), .Z(n11337) );
  XNOR U11243 ( .A(n11339), .B(n11336), .Z(n11338) );
  XOR U11244 ( .A(n11340), .B(n11341), .Z(n11313) );
  AND U11245 ( .A(n11342), .B(n11343), .Z(n11341) );
  XNOR U11246 ( .A(n11340), .B(n11329), .Z(n11343) );
  IV U11247 ( .A(n11275), .Z(n11329) );
  XNOR U11248 ( .A(n11344), .B(n11322), .Z(n11275) );
  XNOR U11249 ( .A(n11345), .B(n11328), .Z(n11322) );
  XOR U11250 ( .A(n11346), .B(n11347), .Z(n11328) );
  NOR U11251 ( .A(n11348), .B(n11349), .Z(n11347) );
  XNOR U11252 ( .A(n11346), .B(n11350), .Z(n11348) );
  XNOR U11253 ( .A(n11327), .B(n11319), .Z(n11345) );
  XOR U11254 ( .A(n11351), .B(n11352), .Z(n11319) );
  AND U11255 ( .A(n11353), .B(n11354), .Z(n11352) );
  XNOR U11256 ( .A(n11351), .B(n11355), .Z(n11353) );
  XNOR U11257 ( .A(n11356), .B(n11324), .Z(n11327) );
  XOR U11258 ( .A(n11357), .B(n11358), .Z(n11324) );
  AND U11259 ( .A(n11359), .B(n11360), .Z(n11358) );
  XOR U11260 ( .A(n11357), .B(n11361), .Z(n11359) );
  XNOR U11261 ( .A(n11362), .B(n11363), .Z(n11356) );
  NOR U11262 ( .A(n11364), .B(n11365), .Z(n11363) );
  XOR U11263 ( .A(n11362), .B(n11366), .Z(n11364) );
  XNOR U11264 ( .A(n11323), .B(n11330), .Z(n11344) );
  NOR U11265 ( .A(n11287), .B(n11367), .Z(n11330) );
  XOR U11266 ( .A(n11335), .B(n11334), .Z(n11323) );
  XNOR U11267 ( .A(n11368), .B(n11331), .Z(n11334) );
  XOR U11268 ( .A(n11369), .B(n11370), .Z(n11331) );
  AND U11269 ( .A(n11371), .B(n11372), .Z(n11370) );
  XOR U11270 ( .A(n11369), .B(n11373), .Z(n11371) );
  XNOR U11271 ( .A(n11374), .B(n11375), .Z(n11368) );
  NOR U11272 ( .A(n11376), .B(n11377), .Z(n11375) );
  XNOR U11273 ( .A(n11374), .B(n11378), .Z(n11376) );
  XOR U11274 ( .A(n11379), .B(n11380), .Z(n11335) );
  NOR U11275 ( .A(n11381), .B(n11382), .Z(n11380) );
  XNOR U11276 ( .A(n11379), .B(n11383), .Z(n11381) );
  XNOR U11277 ( .A(n11272), .B(n11340), .Z(n11342) );
  XOR U11278 ( .A(n11384), .B(n11385), .Z(n11272) );
  AND U11279 ( .A(n187), .B(n11386), .Z(n11385) );
  XOR U11280 ( .A(n11387), .B(n11384), .Z(n11386) );
  AND U11281 ( .A(n11284), .B(n11287), .Z(n11340) );
  XOR U11282 ( .A(n11388), .B(n11367), .Z(n11287) );
  XNOR U11283 ( .A(p_input[2048]), .B(p_input[720]), .Z(n11367) );
  XOR U11284 ( .A(n11355), .B(n11354), .Z(n11388) );
  XNOR U11285 ( .A(n11389), .B(n11361), .Z(n11354) );
  XNOR U11286 ( .A(n11350), .B(n11349), .Z(n11361) );
  XOR U11287 ( .A(n11390), .B(n11346), .Z(n11349) );
  XNOR U11288 ( .A(n6439), .B(p_input[730]), .Z(n11346) );
  XNOR U11289 ( .A(p_input[2059]), .B(p_input[731]), .Z(n11390) );
  XOR U11290 ( .A(p_input[2060]), .B(p_input[732]), .Z(n11350) );
  XNOR U11291 ( .A(n11360), .B(n11351), .Z(n11389) );
  XNOR U11292 ( .A(n6553), .B(p_input[721]), .Z(n11351) );
  XOR U11293 ( .A(n11391), .B(n11366), .Z(n11360) );
  XNOR U11294 ( .A(p_input[2063]), .B(p_input[735]), .Z(n11366) );
  XOR U11295 ( .A(n11357), .B(n11365), .Z(n11391) );
  XOR U11296 ( .A(n11392), .B(n11362), .Z(n11365) );
  XOR U11297 ( .A(p_input[2061]), .B(p_input[733]), .Z(n11362) );
  XNOR U11298 ( .A(p_input[2062]), .B(p_input[734]), .Z(n11392) );
  XNOR U11299 ( .A(n6325), .B(p_input[729]), .Z(n11357) );
  XNOR U11300 ( .A(n11373), .B(n11372), .Z(n11355) );
  XNOR U11301 ( .A(n11393), .B(n11378), .Z(n11372) );
  XOR U11302 ( .A(p_input[2056]), .B(p_input[728]), .Z(n11378) );
  XOR U11303 ( .A(n11369), .B(n11377), .Z(n11393) );
  XOR U11304 ( .A(n11394), .B(n11374), .Z(n11377) );
  XOR U11305 ( .A(p_input[2054]), .B(p_input[726]), .Z(n11374) );
  XNOR U11306 ( .A(p_input[2055]), .B(p_input[727]), .Z(n11394) );
  XNOR U11307 ( .A(n6328), .B(p_input[722]), .Z(n11369) );
  XNOR U11308 ( .A(n11383), .B(n11382), .Z(n11373) );
  XOR U11309 ( .A(n11395), .B(n11379), .Z(n11382) );
  XOR U11310 ( .A(p_input[2051]), .B(p_input[723]), .Z(n11379) );
  XNOR U11311 ( .A(p_input[2052]), .B(p_input[724]), .Z(n11395) );
  XOR U11312 ( .A(p_input[2053]), .B(p_input[725]), .Z(n11383) );
  XOR U11313 ( .A(n11396), .B(n11397), .Z(n11284) );
  AND U11314 ( .A(n187), .B(n11398), .Z(n11397) );
  XNOR U11315 ( .A(n11399), .B(n11396), .Z(n11398) );
  XNOR U11316 ( .A(n11400), .B(n11401), .Z(n187) );
  AND U11317 ( .A(n11402), .B(n11403), .Z(n11401) );
  XOR U11318 ( .A(n11297), .B(n11400), .Z(n11403) );
  AND U11319 ( .A(n11404), .B(n11405), .Z(n11297) );
  XNOR U11320 ( .A(n11294), .B(n11400), .Z(n11402) );
  XOR U11321 ( .A(n11406), .B(n11407), .Z(n11294) );
  AND U11322 ( .A(n191), .B(n11408), .Z(n11407) );
  XOR U11323 ( .A(n11409), .B(n11406), .Z(n11408) );
  XOR U11324 ( .A(n11410), .B(n11411), .Z(n11400) );
  AND U11325 ( .A(n11412), .B(n11413), .Z(n11411) );
  XNOR U11326 ( .A(n11410), .B(n11404), .Z(n11413) );
  IV U11327 ( .A(n11312), .Z(n11404) );
  XOR U11328 ( .A(n11414), .B(n11415), .Z(n11312) );
  XOR U11329 ( .A(n11416), .B(n11405), .Z(n11415) );
  AND U11330 ( .A(n11339), .B(n11417), .Z(n11405) );
  AND U11331 ( .A(n11418), .B(n11419), .Z(n11416) );
  XOR U11332 ( .A(n11420), .B(n11414), .Z(n11418) );
  XNOR U11333 ( .A(n11309), .B(n11410), .Z(n11412) );
  XOR U11334 ( .A(n11421), .B(n11422), .Z(n11309) );
  AND U11335 ( .A(n191), .B(n11423), .Z(n11422) );
  XOR U11336 ( .A(n11424), .B(n11421), .Z(n11423) );
  XOR U11337 ( .A(n11425), .B(n11426), .Z(n11410) );
  AND U11338 ( .A(n11427), .B(n11428), .Z(n11426) );
  XNOR U11339 ( .A(n11425), .B(n11339), .Z(n11428) );
  XOR U11340 ( .A(n11429), .B(n11419), .Z(n11339) );
  XNOR U11341 ( .A(n11430), .B(n11414), .Z(n11419) );
  XOR U11342 ( .A(n11431), .B(n11432), .Z(n11414) );
  AND U11343 ( .A(n11433), .B(n11434), .Z(n11432) );
  XOR U11344 ( .A(n11435), .B(n11431), .Z(n11433) );
  XNOR U11345 ( .A(n11436), .B(n11437), .Z(n11430) );
  AND U11346 ( .A(n11438), .B(n11439), .Z(n11437) );
  XOR U11347 ( .A(n11436), .B(n11440), .Z(n11438) );
  XNOR U11348 ( .A(n11420), .B(n11417), .Z(n11429) );
  AND U11349 ( .A(n11441), .B(n11442), .Z(n11417) );
  XOR U11350 ( .A(n11443), .B(n11444), .Z(n11420) );
  AND U11351 ( .A(n11445), .B(n11446), .Z(n11444) );
  XOR U11352 ( .A(n11443), .B(n11447), .Z(n11445) );
  XNOR U11353 ( .A(n11336), .B(n11425), .Z(n11427) );
  XOR U11354 ( .A(n11448), .B(n11449), .Z(n11336) );
  AND U11355 ( .A(n191), .B(n11450), .Z(n11449) );
  XNOR U11356 ( .A(n11451), .B(n11448), .Z(n11450) );
  XOR U11357 ( .A(n11452), .B(n11453), .Z(n11425) );
  AND U11358 ( .A(n11454), .B(n11455), .Z(n11453) );
  XNOR U11359 ( .A(n11452), .B(n11441), .Z(n11455) );
  IV U11360 ( .A(n11387), .Z(n11441) );
  XNOR U11361 ( .A(n11456), .B(n11434), .Z(n11387) );
  XNOR U11362 ( .A(n11457), .B(n11440), .Z(n11434) );
  XOR U11363 ( .A(n11458), .B(n11459), .Z(n11440) );
  NOR U11364 ( .A(n11460), .B(n11461), .Z(n11459) );
  XNOR U11365 ( .A(n11458), .B(n11462), .Z(n11460) );
  XNOR U11366 ( .A(n11439), .B(n11431), .Z(n11457) );
  XOR U11367 ( .A(n11463), .B(n11464), .Z(n11431) );
  AND U11368 ( .A(n11465), .B(n11466), .Z(n11464) );
  XNOR U11369 ( .A(n11463), .B(n11467), .Z(n11465) );
  XNOR U11370 ( .A(n11468), .B(n11436), .Z(n11439) );
  XOR U11371 ( .A(n11469), .B(n11470), .Z(n11436) );
  AND U11372 ( .A(n11471), .B(n11472), .Z(n11470) );
  XOR U11373 ( .A(n11469), .B(n11473), .Z(n11471) );
  XNOR U11374 ( .A(n11474), .B(n11475), .Z(n11468) );
  NOR U11375 ( .A(n11476), .B(n11477), .Z(n11475) );
  XOR U11376 ( .A(n11474), .B(n11478), .Z(n11476) );
  XNOR U11377 ( .A(n11435), .B(n11442), .Z(n11456) );
  NOR U11378 ( .A(n11399), .B(n11479), .Z(n11442) );
  XOR U11379 ( .A(n11447), .B(n11446), .Z(n11435) );
  XNOR U11380 ( .A(n11480), .B(n11443), .Z(n11446) );
  XOR U11381 ( .A(n11481), .B(n11482), .Z(n11443) );
  AND U11382 ( .A(n11483), .B(n11484), .Z(n11482) );
  XOR U11383 ( .A(n11481), .B(n11485), .Z(n11483) );
  XNOR U11384 ( .A(n11486), .B(n11487), .Z(n11480) );
  NOR U11385 ( .A(n11488), .B(n11489), .Z(n11487) );
  XNOR U11386 ( .A(n11486), .B(n11490), .Z(n11488) );
  XOR U11387 ( .A(n11491), .B(n11492), .Z(n11447) );
  NOR U11388 ( .A(n11493), .B(n11494), .Z(n11492) );
  XNOR U11389 ( .A(n11491), .B(n11495), .Z(n11493) );
  XNOR U11390 ( .A(n11384), .B(n11452), .Z(n11454) );
  XOR U11391 ( .A(n11496), .B(n11497), .Z(n11384) );
  AND U11392 ( .A(n191), .B(n11498), .Z(n11497) );
  XOR U11393 ( .A(n11499), .B(n11496), .Z(n11498) );
  AND U11394 ( .A(n11396), .B(n11399), .Z(n11452) );
  XOR U11395 ( .A(n11500), .B(n11479), .Z(n11399) );
  XNOR U11396 ( .A(p_input[2048]), .B(p_input[736]), .Z(n11479) );
  XOR U11397 ( .A(n11467), .B(n11466), .Z(n11500) );
  XNOR U11398 ( .A(n11501), .B(n11473), .Z(n11466) );
  XNOR U11399 ( .A(n11462), .B(n11461), .Z(n11473) );
  XOR U11400 ( .A(n11502), .B(n11458), .Z(n11461) );
  XNOR U11401 ( .A(n6439), .B(p_input[746]), .Z(n11458) );
  XNOR U11402 ( .A(p_input[2059]), .B(p_input[747]), .Z(n11502) );
  XOR U11403 ( .A(p_input[2060]), .B(p_input[748]), .Z(n11462) );
  XNOR U11404 ( .A(n11472), .B(n11463), .Z(n11501) );
  XNOR U11405 ( .A(n6553), .B(p_input[737]), .Z(n11463) );
  XOR U11406 ( .A(n11503), .B(n11478), .Z(n11472) );
  XNOR U11407 ( .A(p_input[2063]), .B(p_input[751]), .Z(n11478) );
  XOR U11408 ( .A(n11469), .B(n11477), .Z(n11503) );
  XOR U11409 ( .A(n11504), .B(n11474), .Z(n11477) );
  XOR U11410 ( .A(p_input[2061]), .B(p_input[749]), .Z(n11474) );
  XNOR U11411 ( .A(p_input[2062]), .B(p_input[750]), .Z(n11504) );
  XNOR U11412 ( .A(n6325), .B(p_input[745]), .Z(n11469) );
  XNOR U11413 ( .A(n11485), .B(n11484), .Z(n11467) );
  XNOR U11414 ( .A(n11505), .B(n11490), .Z(n11484) );
  XOR U11415 ( .A(p_input[2056]), .B(p_input[744]), .Z(n11490) );
  XOR U11416 ( .A(n11481), .B(n11489), .Z(n11505) );
  XOR U11417 ( .A(n11506), .B(n11486), .Z(n11489) );
  XOR U11418 ( .A(p_input[2054]), .B(p_input[742]), .Z(n11486) );
  XNOR U11419 ( .A(p_input[2055]), .B(p_input[743]), .Z(n11506) );
  XNOR U11420 ( .A(n6328), .B(p_input[738]), .Z(n11481) );
  XNOR U11421 ( .A(n11495), .B(n11494), .Z(n11485) );
  XOR U11422 ( .A(n11507), .B(n11491), .Z(n11494) );
  XOR U11423 ( .A(p_input[2051]), .B(p_input[739]), .Z(n11491) );
  XNOR U11424 ( .A(p_input[2052]), .B(p_input[740]), .Z(n11507) );
  XOR U11425 ( .A(p_input[2053]), .B(p_input[741]), .Z(n11495) );
  XOR U11426 ( .A(n11508), .B(n11509), .Z(n11396) );
  AND U11427 ( .A(n191), .B(n11510), .Z(n11509) );
  XNOR U11428 ( .A(n11511), .B(n11508), .Z(n11510) );
  XNOR U11429 ( .A(n11512), .B(n11513), .Z(n191) );
  AND U11430 ( .A(n11514), .B(n11515), .Z(n11513) );
  XOR U11431 ( .A(n11409), .B(n11512), .Z(n11515) );
  AND U11432 ( .A(n11516), .B(n11517), .Z(n11409) );
  XNOR U11433 ( .A(n11406), .B(n11512), .Z(n11514) );
  XOR U11434 ( .A(n11518), .B(n11519), .Z(n11406) );
  AND U11435 ( .A(n195), .B(n11520), .Z(n11519) );
  XOR U11436 ( .A(n11521), .B(n11518), .Z(n11520) );
  XOR U11437 ( .A(n11522), .B(n11523), .Z(n11512) );
  AND U11438 ( .A(n11524), .B(n11525), .Z(n11523) );
  XNOR U11439 ( .A(n11522), .B(n11516), .Z(n11525) );
  IV U11440 ( .A(n11424), .Z(n11516) );
  XOR U11441 ( .A(n11526), .B(n11527), .Z(n11424) );
  XOR U11442 ( .A(n11528), .B(n11517), .Z(n11527) );
  AND U11443 ( .A(n11451), .B(n11529), .Z(n11517) );
  AND U11444 ( .A(n11530), .B(n11531), .Z(n11528) );
  XOR U11445 ( .A(n11532), .B(n11526), .Z(n11530) );
  XNOR U11446 ( .A(n11421), .B(n11522), .Z(n11524) );
  XOR U11447 ( .A(n11533), .B(n11534), .Z(n11421) );
  AND U11448 ( .A(n195), .B(n11535), .Z(n11534) );
  XOR U11449 ( .A(n11536), .B(n11533), .Z(n11535) );
  XOR U11450 ( .A(n11537), .B(n11538), .Z(n11522) );
  AND U11451 ( .A(n11539), .B(n11540), .Z(n11538) );
  XNOR U11452 ( .A(n11537), .B(n11451), .Z(n11540) );
  XOR U11453 ( .A(n11541), .B(n11531), .Z(n11451) );
  XNOR U11454 ( .A(n11542), .B(n11526), .Z(n11531) );
  XOR U11455 ( .A(n11543), .B(n11544), .Z(n11526) );
  AND U11456 ( .A(n11545), .B(n11546), .Z(n11544) );
  XOR U11457 ( .A(n11547), .B(n11543), .Z(n11545) );
  XNOR U11458 ( .A(n11548), .B(n11549), .Z(n11542) );
  AND U11459 ( .A(n11550), .B(n11551), .Z(n11549) );
  XOR U11460 ( .A(n11548), .B(n11552), .Z(n11550) );
  XNOR U11461 ( .A(n11532), .B(n11529), .Z(n11541) );
  AND U11462 ( .A(n11553), .B(n11554), .Z(n11529) );
  XOR U11463 ( .A(n11555), .B(n11556), .Z(n11532) );
  AND U11464 ( .A(n11557), .B(n11558), .Z(n11556) );
  XOR U11465 ( .A(n11555), .B(n11559), .Z(n11557) );
  XNOR U11466 ( .A(n11448), .B(n11537), .Z(n11539) );
  XOR U11467 ( .A(n11560), .B(n11561), .Z(n11448) );
  AND U11468 ( .A(n195), .B(n11562), .Z(n11561) );
  XNOR U11469 ( .A(n11563), .B(n11560), .Z(n11562) );
  XOR U11470 ( .A(n11564), .B(n11565), .Z(n11537) );
  AND U11471 ( .A(n11566), .B(n11567), .Z(n11565) );
  XNOR U11472 ( .A(n11564), .B(n11553), .Z(n11567) );
  IV U11473 ( .A(n11499), .Z(n11553) );
  XNOR U11474 ( .A(n11568), .B(n11546), .Z(n11499) );
  XNOR U11475 ( .A(n11569), .B(n11552), .Z(n11546) );
  XOR U11476 ( .A(n11570), .B(n11571), .Z(n11552) );
  NOR U11477 ( .A(n11572), .B(n11573), .Z(n11571) );
  XNOR U11478 ( .A(n11570), .B(n11574), .Z(n11572) );
  XNOR U11479 ( .A(n11551), .B(n11543), .Z(n11569) );
  XOR U11480 ( .A(n11575), .B(n11576), .Z(n11543) );
  AND U11481 ( .A(n11577), .B(n11578), .Z(n11576) );
  XNOR U11482 ( .A(n11575), .B(n11579), .Z(n11577) );
  XNOR U11483 ( .A(n11580), .B(n11548), .Z(n11551) );
  XOR U11484 ( .A(n11581), .B(n11582), .Z(n11548) );
  AND U11485 ( .A(n11583), .B(n11584), .Z(n11582) );
  XOR U11486 ( .A(n11581), .B(n11585), .Z(n11583) );
  XNOR U11487 ( .A(n11586), .B(n11587), .Z(n11580) );
  NOR U11488 ( .A(n11588), .B(n11589), .Z(n11587) );
  XOR U11489 ( .A(n11586), .B(n11590), .Z(n11588) );
  XNOR U11490 ( .A(n11547), .B(n11554), .Z(n11568) );
  NOR U11491 ( .A(n11511), .B(n11591), .Z(n11554) );
  XOR U11492 ( .A(n11559), .B(n11558), .Z(n11547) );
  XNOR U11493 ( .A(n11592), .B(n11555), .Z(n11558) );
  XOR U11494 ( .A(n11593), .B(n11594), .Z(n11555) );
  AND U11495 ( .A(n11595), .B(n11596), .Z(n11594) );
  XOR U11496 ( .A(n11593), .B(n11597), .Z(n11595) );
  XNOR U11497 ( .A(n11598), .B(n11599), .Z(n11592) );
  NOR U11498 ( .A(n11600), .B(n11601), .Z(n11599) );
  XNOR U11499 ( .A(n11598), .B(n11602), .Z(n11600) );
  XOR U11500 ( .A(n11603), .B(n11604), .Z(n11559) );
  NOR U11501 ( .A(n11605), .B(n11606), .Z(n11604) );
  XNOR U11502 ( .A(n11603), .B(n11607), .Z(n11605) );
  XNOR U11503 ( .A(n11496), .B(n11564), .Z(n11566) );
  XOR U11504 ( .A(n11608), .B(n11609), .Z(n11496) );
  AND U11505 ( .A(n195), .B(n11610), .Z(n11609) );
  XOR U11506 ( .A(n11611), .B(n11608), .Z(n11610) );
  AND U11507 ( .A(n11508), .B(n11511), .Z(n11564) );
  XOR U11508 ( .A(n11612), .B(n11591), .Z(n11511) );
  XNOR U11509 ( .A(p_input[2048]), .B(p_input[752]), .Z(n11591) );
  XOR U11510 ( .A(n11579), .B(n11578), .Z(n11612) );
  XNOR U11511 ( .A(n11613), .B(n11585), .Z(n11578) );
  XNOR U11512 ( .A(n11574), .B(n11573), .Z(n11585) );
  XOR U11513 ( .A(n11614), .B(n11570), .Z(n11573) );
  XNOR U11514 ( .A(n6439), .B(p_input[762]), .Z(n11570) );
  XNOR U11515 ( .A(p_input[2059]), .B(p_input[763]), .Z(n11614) );
  XOR U11516 ( .A(p_input[2060]), .B(p_input[764]), .Z(n11574) );
  XNOR U11517 ( .A(n11584), .B(n11575), .Z(n11613) );
  XNOR U11518 ( .A(n6553), .B(p_input[753]), .Z(n11575) );
  XOR U11519 ( .A(n11615), .B(n11590), .Z(n11584) );
  XNOR U11520 ( .A(p_input[2063]), .B(p_input[767]), .Z(n11590) );
  XOR U11521 ( .A(n11581), .B(n11589), .Z(n11615) );
  XOR U11522 ( .A(n11616), .B(n11586), .Z(n11589) );
  XOR U11523 ( .A(p_input[2061]), .B(p_input[765]), .Z(n11586) );
  XNOR U11524 ( .A(p_input[2062]), .B(p_input[766]), .Z(n11616) );
  XNOR U11525 ( .A(n6325), .B(p_input[761]), .Z(n11581) );
  XNOR U11526 ( .A(n11597), .B(n11596), .Z(n11579) );
  XNOR U11527 ( .A(n11617), .B(n11602), .Z(n11596) );
  XOR U11528 ( .A(p_input[2056]), .B(p_input[760]), .Z(n11602) );
  XOR U11529 ( .A(n11593), .B(n11601), .Z(n11617) );
  XOR U11530 ( .A(n11618), .B(n11598), .Z(n11601) );
  XOR U11531 ( .A(p_input[2054]), .B(p_input[758]), .Z(n11598) );
  XNOR U11532 ( .A(p_input[2055]), .B(p_input[759]), .Z(n11618) );
  XNOR U11533 ( .A(n6328), .B(p_input[754]), .Z(n11593) );
  XNOR U11534 ( .A(n11607), .B(n11606), .Z(n11597) );
  XOR U11535 ( .A(n11619), .B(n11603), .Z(n11606) );
  XOR U11536 ( .A(p_input[2051]), .B(p_input[755]), .Z(n11603) );
  XNOR U11537 ( .A(p_input[2052]), .B(p_input[756]), .Z(n11619) );
  XOR U11538 ( .A(p_input[2053]), .B(p_input[757]), .Z(n11607) );
  XOR U11539 ( .A(n11620), .B(n11621), .Z(n11508) );
  AND U11540 ( .A(n195), .B(n11622), .Z(n11621) );
  XNOR U11541 ( .A(n11623), .B(n11620), .Z(n11622) );
  XNOR U11542 ( .A(n11624), .B(n11625), .Z(n195) );
  AND U11543 ( .A(n11626), .B(n11627), .Z(n11625) );
  XOR U11544 ( .A(n11521), .B(n11624), .Z(n11627) );
  AND U11545 ( .A(n11628), .B(n11629), .Z(n11521) );
  XNOR U11546 ( .A(n11518), .B(n11624), .Z(n11626) );
  XOR U11547 ( .A(n11630), .B(n11631), .Z(n11518) );
  AND U11548 ( .A(n199), .B(n11632), .Z(n11631) );
  XOR U11549 ( .A(n11633), .B(n11630), .Z(n11632) );
  XOR U11550 ( .A(n11634), .B(n11635), .Z(n11624) );
  AND U11551 ( .A(n11636), .B(n11637), .Z(n11635) );
  XNOR U11552 ( .A(n11634), .B(n11628), .Z(n11637) );
  IV U11553 ( .A(n11536), .Z(n11628) );
  XOR U11554 ( .A(n11638), .B(n11639), .Z(n11536) );
  XOR U11555 ( .A(n11640), .B(n11629), .Z(n11639) );
  AND U11556 ( .A(n11563), .B(n11641), .Z(n11629) );
  AND U11557 ( .A(n11642), .B(n11643), .Z(n11640) );
  XOR U11558 ( .A(n11644), .B(n11638), .Z(n11642) );
  XNOR U11559 ( .A(n11533), .B(n11634), .Z(n11636) );
  XOR U11560 ( .A(n11645), .B(n11646), .Z(n11533) );
  AND U11561 ( .A(n199), .B(n11647), .Z(n11646) );
  XOR U11562 ( .A(n11648), .B(n11645), .Z(n11647) );
  XOR U11563 ( .A(n11649), .B(n11650), .Z(n11634) );
  AND U11564 ( .A(n11651), .B(n11652), .Z(n11650) );
  XNOR U11565 ( .A(n11649), .B(n11563), .Z(n11652) );
  XOR U11566 ( .A(n11653), .B(n11643), .Z(n11563) );
  XNOR U11567 ( .A(n11654), .B(n11638), .Z(n11643) );
  XOR U11568 ( .A(n11655), .B(n11656), .Z(n11638) );
  AND U11569 ( .A(n11657), .B(n11658), .Z(n11656) );
  XOR U11570 ( .A(n11659), .B(n11655), .Z(n11657) );
  XNOR U11571 ( .A(n11660), .B(n11661), .Z(n11654) );
  AND U11572 ( .A(n11662), .B(n11663), .Z(n11661) );
  XOR U11573 ( .A(n11660), .B(n11664), .Z(n11662) );
  XNOR U11574 ( .A(n11644), .B(n11641), .Z(n11653) );
  AND U11575 ( .A(n11665), .B(n11666), .Z(n11641) );
  XOR U11576 ( .A(n11667), .B(n11668), .Z(n11644) );
  AND U11577 ( .A(n11669), .B(n11670), .Z(n11668) );
  XOR U11578 ( .A(n11667), .B(n11671), .Z(n11669) );
  XNOR U11579 ( .A(n11560), .B(n11649), .Z(n11651) );
  XOR U11580 ( .A(n11672), .B(n11673), .Z(n11560) );
  AND U11581 ( .A(n199), .B(n11674), .Z(n11673) );
  XNOR U11582 ( .A(n11675), .B(n11672), .Z(n11674) );
  XOR U11583 ( .A(n11676), .B(n11677), .Z(n11649) );
  AND U11584 ( .A(n11678), .B(n11679), .Z(n11677) );
  XNOR U11585 ( .A(n11676), .B(n11665), .Z(n11679) );
  IV U11586 ( .A(n11611), .Z(n11665) );
  XNOR U11587 ( .A(n11680), .B(n11658), .Z(n11611) );
  XNOR U11588 ( .A(n11681), .B(n11664), .Z(n11658) );
  XOR U11589 ( .A(n11682), .B(n11683), .Z(n11664) );
  NOR U11590 ( .A(n11684), .B(n11685), .Z(n11683) );
  XNOR U11591 ( .A(n11682), .B(n11686), .Z(n11684) );
  XNOR U11592 ( .A(n11663), .B(n11655), .Z(n11681) );
  XOR U11593 ( .A(n11687), .B(n11688), .Z(n11655) );
  AND U11594 ( .A(n11689), .B(n11690), .Z(n11688) );
  XNOR U11595 ( .A(n11687), .B(n11691), .Z(n11689) );
  XNOR U11596 ( .A(n11692), .B(n11660), .Z(n11663) );
  XOR U11597 ( .A(n11693), .B(n11694), .Z(n11660) );
  AND U11598 ( .A(n11695), .B(n11696), .Z(n11694) );
  XOR U11599 ( .A(n11693), .B(n11697), .Z(n11695) );
  XNOR U11600 ( .A(n11698), .B(n11699), .Z(n11692) );
  NOR U11601 ( .A(n11700), .B(n11701), .Z(n11699) );
  XOR U11602 ( .A(n11698), .B(n11702), .Z(n11700) );
  XNOR U11603 ( .A(n11659), .B(n11666), .Z(n11680) );
  NOR U11604 ( .A(n11623), .B(n11703), .Z(n11666) );
  XOR U11605 ( .A(n11671), .B(n11670), .Z(n11659) );
  XNOR U11606 ( .A(n11704), .B(n11667), .Z(n11670) );
  XOR U11607 ( .A(n11705), .B(n11706), .Z(n11667) );
  AND U11608 ( .A(n11707), .B(n11708), .Z(n11706) );
  XOR U11609 ( .A(n11705), .B(n11709), .Z(n11707) );
  XNOR U11610 ( .A(n11710), .B(n11711), .Z(n11704) );
  NOR U11611 ( .A(n11712), .B(n11713), .Z(n11711) );
  XNOR U11612 ( .A(n11710), .B(n11714), .Z(n11712) );
  XOR U11613 ( .A(n11715), .B(n11716), .Z(n11671) );
  NOR U11614 ( .A(n11717), .B(n11718), .Z(n11716) );
  XNOR U11615 ( .A(n11715), .B(n11719), .Z(n11717) );
  XNOR U11616 ( .A(n11608), .B(n11676), .Z(n11678) );
  XOR U11617 ( .A(n11720), .B(n11721), .Z(n11608) );
  AND U11618 ( .A(n199), .B(n11722), .Z(n11721) );
  XOR U11619 ( .A(n11723), .B(n11720), .Z(n11722) );
  AND U11620 ( .A(n11620), .B(n11623), .Z(n11676) );
  XOR U11621 ( .A(n11724), .B(n11703), .Z(n11623) );
  XNOR U11622 ( .A(p_input[2048]), .B(p_input[768]), .Z(n11703) );
  XOR U11623 ( .A(n11691), .B(n11690), .Z(n11724) );
  XNOR U11624 ( .A(n11725), .B(n11697), .Z(n11690) );
  XNOR U11625 ( .A(n11686), .B(n11685), .Z(n11697) );
  XOR U11626 ( .A(n11726), .B(n11682), .Z(n11685) );
  XNOR U11627 ( .A(n6439), .B(p_input[778]), .Z(n11682) );
  XNOR U11628 ( .A(p_input[2059]), .B(p_input[779]), .Z(n11726) );
  XOR U11629 ( .A(p_input[2060]), .B(p_input[780]), .Z(n11686) );
  XNOR U11630 ( .A(n11696), .B(n11687), .Z(n11725) );
  XNOR U11631 ( .A(n6553), .B(p_input[769]), .Z(n11687) );
  XOR U11632 ( .A(n11727), .B(n11702), .Z(n11696) );
  XNOR U11633 ( .A(p_input[2063]), .B(p_input[783]), .Z(n11702) );
  XOR U11634 ( .A(n11693), .B(n11701), .Z(n11727) );
  XOR U11635 ( .A(n11728), .B(n11698), .Z(n11701) );
  XOR U11636 ( .A(p_input[2061]), .B(p_input[781]), .Z(n11698) );
  XNOR U11637 ( .A(p_input[2062]), .B(p_input[782]), .Z(n11728) );
  XNOR U11638 ( .A(n6325), .B(p_input[777]), .Z(n11693) );
  XNOR U11639 ( .A(n11709), .B(n11708), .Z(n11691) );
  XNOR U11640 ( .A(n11729), .B(n11714), .Z(n11708) );
  XOR U11641 ( .A(p_input[2056]), .B(p_input[776]), .Z(n11714) );
  XOR U11642 ( .A(n11705), .B(n11713), .Z(n11729) );
  XOR U11643 ( .A(n11730), .B(n11710), .Z(n11713) );
  XOR U11644 ( .A(p_input[2054]), .B(p_input[774]), .Z(n11710) );
  XNOR U11645 ( .A(p_input[2055]), .B(p_input[775]), .Z(n11730) );
  XNOR U11646 ( .A(n6328), .B(p_input[770]), .Z(n11705) );
  XNOR U11647 ( .A(n11719), .B(n11718), .Z(n11709) );
  XOR U11648 ( .A(n11731), .B(n11715), .Z(n11718) );
  XOR U11649 ( .A(p_input[2051]), .B(p_input[771]), .Z(n11715) );
  XNOR U11650 ( .A(p_input[2052]), .B(p_input[772]), .Z(n11731) );
  XOR U11651 ( .A(p_input[2053]), .B(p_input[773]), .Z(n11719) );
  XOR U11652 ( .A(n11732), .B(n11733), .Z(n11620) );
  AND U11653 ( .A(n199), .B(n11734), .Z(n11733) );
  XNOR U11654 ( .A(n11735), .B(n11732), .Z(n11734) );
  XNOR U11655 ( .A(n11736), .B(n11737), .Z(n199) );
  AND U11656 ( .A(n11738), .B(n11739), .Z(n11737) );
  XOR U11657 ( .A(n11633), .B(n11736), .Z(n11739) );
  AND U11658 ( .A(n11740), .B(n11741), .Z(n11633) );
  XNOR U11659 ( .A(n11630), .B(n11736), .Z(n11738) );
  XOR U11660 ( .A(n11742), .B(n11743), .Z(n11630) );
  AND U11661 ( .A(n203), .B(n11744), .Z(n11743) );
  XOR U11662 ( .A(n11745), .B(n11742), .Z(n11744) );
  XOR U11663 ( .A(n11746), .B(n11747), .Z(n11736) );
  AND U11664 ( .A(n11748), .B(n11749), .Z(n11747) );
  XNOR U11665 ( .A(n11746), .B(n11740), .Z(n11749) );
  IV U11666 ( .A(n11648), .Z(n11740) );
  XOR U11667 ( .A(n11750), .B(n11751), .Z(n11648) );
  XOR U11668 ( .A(n11752), .B(n11741), .Z(n11751) );
  AND U11669 ( .A(n11675), .B(n11753), .Z(n11741) );
  AND U11670 ( .A(n11754), .B(n11755), .Z(n11752) );
  XOR U11671 ( .A(n11756), .B(n11750), .Z(n11754) );
  XNOR U11672 ( .A(n11645), .B(n11746), .Z(n11748) );
  XOR U11673 ( .A(n11757), .B(n11758), .Z(n11645) );
  AND U11674 ( .A(n203), .B(n11759), .Z(n11758) );
  XOR U11675 ( .A(n11760), .B(n11757), .Z(n11759) );
  XOR U11676 ( .A(n11761), .B(n11762), .Z(n11746) );
  AND U11677 ( .A(n11763), .B(n11764), .Z(n11762) );
  XNOR U11678 ( .A(n11761), .B(n11675), .Z(n11764) );
  XOR U11679 ( .A(n11765), .B(n11755), .Z(n11675) );
  XNOR U11680 ( .A(n11766), .B(n11750), .Z(n11755) );
  XOR U11681 ( .A(n11767), .B(n11768), .Z(n11750) );
  AND U11682 ( .A(n11769), .B(n11770), .Z(n11768) );
  XOR U11683 ( .A(n11771), .B(n11767), .Z(n11769) );
  XNOR U11684 ( .A(n11772), .B(n11773), .Z(n11766) );
  AND U11685 ( .A(n11774), .B(n11775), .Z(n11773) );
  XOR U11686 ( .A(n11772), .B(n11776), .Z(n11774) );
  XNOR U11687 ( .A(n11756), .B(n11753), .Z(n11765) );
  AND U11688 ( .A(n11777), .B(n11778), .Z(n11753) );
  XOR U11689 ( .A(n11779), .B(n11780), .Z(n11756) );
  AND U11690 ( .A(n11781), .B(n11782), .Z(n11780) );
  XOR U11691 ( .A(n11779), .B(n11783), .Z(n11781) );
  XNOR U11692 ( .A(n11672), .B(n11761), .Z(n11763) );
  XOR U11693 ( .A(n11784), .B(n11785), .Z(n11672) );
  AND U11694 ( .A(n203), .B(n11786), .Z(n11785) );
  XNOR U11695 ( .A(n11787), .B(n11784), .Z(n11786) );
  XOR U11696 ( .A(n11788), .B(n11789), .Z(n11761) );
  AND U11697 ( .A(n11790), .B(n11791), .Z(n11789) );
  XNOR U11698 ( .A(n11788), .B(n11777), .Z(n11791) );
  IV U11699 ( .A(n11723), .Z(n11777) );
  XNOR U11700 ( .A(n11792), .B(n11770), .Z(n11723) );
  XNOR U11701 ( .A(n11793), .B(n11776), .Z(n11770) );
  XOR U11702 ( .A(n11794), .B(n11795), .Z(n11776) );
  NOR U11703 ( .A(n11796), .B(n11797), .Z(n11795) );
  XNOR U11704 ( .A(n11794), .B(n11798), .Z(n11796) );
  XNOR U11705 ( .A(n11775), .B(n11767), .Z(n11793) );
  XOR U11706 ( .A(n11799), .B(n11800), .Z(n11767) );
  AND U11707 ( .A(n11801), .B(n11802), .Z(n11800) );
  XNOR U11708 ( .A(n11799), .B(n11803), .Z(n11801) );
  XNOR U11709 ( .A(n11804), .B(n11772), .Z(n11775) );
  XOR U11710 ( .A(n11805), .B(n11806), .Z(n11772) );
  AND U11711 ( .A(n11807), .B(n11808), .Z(n11806) );
  XOR U11712 ( .A(n11805), .B(n11809), .Z(n11807) );
  XNOR U11713 ( .A(n11810), .B(n11811), .Z(n11804) );
  NOR U11714 ( .A(n11812), .B(n11813), .Z(n11811) );
  XOR U11715 ( .A(n11810), .B(n11814), .Z(n11812) );
  XNOR U11716 ( .A(n11771), .B(n11778), .Z(n11792) );
  NOR U11717 ( .A(n11735), .B(n11815), .Z(n11778) );
  XOR U11718 ( .A(n11783), .B(n11782), .Z(n11771) );
  XNOR U11719 ( .A(n11816), .B(n11779), .Z(n11782) );
  XOR U11720 ( .A(n11817), .B(n11818), .Z(n11779) );
  AND U11721 ( .A(n11819), .B(n11820), .Z(n11818) );
  XOR U11722 ( .A(n11817), .B(n11821), .Z(n11819) );
  XNOR U11723 ( .A(n11822), .B(n11823), .Z(n11816) );
  NOR U11724 ( .A(n11824), .B(n11825), .Z(n11823) );
  XNOR U11725 ( .A(n11822), .B(n11826), .Z(n11824) );
  XOR U11726 ( .A(n11827), .B(n11828), .Z(n11783) );
  NOR U11727 ( .A(n11829), .B(n11830), .Z(n11828) );
  XNOR U11728 ( .A(n11827), .B(n11831), .Z(n11829) );
  XNOR U11729 ( .A(n11720), .B(n11788), .Z(n11790) );
  XOR U11730 ( .A(n11832), .B(n11833), .Z(n11720) );
  AND U11731 ( .A(n203), .B(n11834), .Z(n11833) );
  XOR U11732 ( .A(n11835), .B(n11832), .Z(n11834) );
  AND U11733 ( .A(n11732), .B(n11735), .Z(n11788) );
  XOR U11734 ( .A(n11836), .B(n11815), .Z(n11735) );
  XNOR U11735 ( .A(p_input[2048]), .B(p_input[784]), .Z(n11815) );
  XOR U11736 ( .A(n11803), .B(n11802), .Z(n11836) );
  XNOR U11737 ( .A(n11837), .B(n11809), .Z(n11802) );
  XNOR U11738 ( .A(n11798), .B(n11797), .Z(n11809) );
  XOR U11739 ( .A(n11838), .B(n11794), .Z(n11797) );
  XNOR U11740 ( .A(n6439), .B(p_input[794]), .Z(n11794) );
  XNOR U11741 ( .A(p_input[2059]), .B(p_input[795]), .Z(n11838) );
  XOR U11742 ( .A(p_input[2060]), .B(p_input[796]), .Z(n11798) );
  XNOR U11743 ( .A(n11808), .B(n11799), .Z(n11837) );
  XNOR U11744 ( .A(n6553), .B(p_input[785]), .Z(n11799) );
  XOR U11745 ( .A(n11839), .B(n11814), .Z(n11808) );
  XNOR U11746 ( .A(p_input[2063]), .B(p_input[799]), .Z(n11814) );
  XOR U11747 ( .A(n11805), .B(n11813), .Z(n11839) );
  XOR U11748 ( .A(n11840), .B(n11810), .Z(n11813) );
  XOR U11749 ( .A(p_input[2061]), .B(p_input[797]), .Z(n11810) );
  XNOR U11750 ( .A(p_input[2062]), .B(p_input[798]), .Z(n11840) );
  XNOR U11751 ( .A(n6325), .B(p_input[793]), .Z(n11805) );
  XNOR U11752 ( .A(n11821), .B(n11820), .Z(n11803) );
  XNOR U11753 ( .A(n11841), .B(n11826), .Z(n11820) );
  XOR U11754 ( .A(p_input[2056]), .B(p_input[792]), .Z(n11826) );
  XOR U11755 ( .A(n11817), .B(n11825), .Z(n11841) );
  XOR U11756 ( .A(n11842), .B(n11822), .Z(n11825) );
  XOR U11757 ( .A(p_input[2054]), .B(p_input[790]), .Z(n11822) );
  XNOR U11758 ( .A(p_input[2055]), .B(p_input[791]), .Z(n11842) );
  XNOR U11759 ( .A(n6328), .B(p_input[786]), .Z(n11817) );
  XNOR U11760 ( .A(n11831), .B(n11830), .Z(n11821) );
  XOR U11761 ( .A(n11843), .B(n11827), .Z(n11830) );
  XOR U11762 ( .A(p_input[2051]), .B(p_input[787]), .Z(n11827) );
  XNOR U11763 ( .A(p_input[2052]), .B(p_input[788]), .Z(n11843) );
  XOR U11764 ( .A(p_input[2053]), .B(p_input[789]), .Z(n11831) );
  XOR U11765 ( .A(n11844), .B(n11845), .Z(n11732) );
  AND U11766 ( .A(n203), .B(n11846), .Z(n11845) );
  XNOR U11767 ( .A(n11847), .B(n11844), .Z(n11846) );
  XNOR U11768 ( .A(n11848), .B(n11849), .Z(n203) );
  AND U11769 ( .A(n11850), .B(n11851), .Z(n11849) );
  XOR U11770 ( .A(n11745), .B(n11848), .Z(n11851) );
  AND U11771 ( .A(n11852), .B(n11853), .Z(n11745) );
  XNOR U11772 ( .A(n11742), .B(n11848), .Z(n11850) );
  XOR U11773 ( .A(n11854), .B(n11855), .Z(n11742) );
  AND U11774 ( .A(n207), .B(n11856), .Z(n11855) );
  XOR U11775 ( .A(n11857), .B(n11854), .Z(n11856) );
  XOR U11776 ( .A(n11858), .B(n11859), .Z(n11848) );
  AND U11777 ( .A(n11860), .B(n11861), .Z(n11859) );
  XNOR U11778 ( .A(n11858), .B(n11852), .Z(n11861) );
  IV U11779 ( .A(n11760), .Z(n11852) );
  XOR U11780 ( .A(n11862), .B(n11863), .Z(n11760) );
  XOR U11781 ( .A(n11864), .B(n11853), .Z(n11863) );
  AND U11782 ( .A(n11787), .B(n11865), .Z(n11853) );
  AND U11783 ( .A(n11866), .B(n11867), .Z(n11864) );
  XOR U11784 ( .A(n11868), .B(n11862), .Z(n11866) );
  XNOR U11785 ( .A(n11757), .B(n11858), .Z(n11860) );
  XOR U11786 ( .A(n11869), .B(n11870), .Z(n11757) );
  AND U11787 ( .A(n207), .B(n11871), .Z(n11870) );
  XOR U11788 ( .A(n11872), .B(n11869), .Z(n11871) );
  XOR U11789 ( .A(n11873), .B(n11874), .Z(n11858) );
  AND U11790 ( .A(n11875), .B(n11876), .Z(n11874) );
  XNOR U11791 ( .A(n11873), .B(n11787), .Z(n11876) );
  XOR U11792 ( .A(n11877), .B(n11867), .Z(n11787) );
  XNOR U11793 ( .A(n11878), .B(n11862), .Z(n11867) );
  XOR U11794 ( .A(n11879), .B(n11880), .Z(n11862) );
  AND U11795 ( .A(n11881), .B(n11882), .Z(n11880) );
  XOR U11796 ( .A(n11883), .B(n11879), .Z(n11881) );
  XNOR U11797 ( .A(n11884), .B(n11885), .Z(n11878) );
  AND U11798 ( .A(n11886), .B(n11887), .Z(n11885) );
  XOR U11799 ( .A(n11884), .B(n11888), .Z(n11886) );
  XNOR U11800 ( .A(n11868), .B(n11865), .Z(n11877) );
  AND U11801 ( .A(n11889), .B(n11890), .Z(n11865) );
  XOR U11802 ( .A(n11891), .B(n11892), .Z(n11868) );
  AND U11803 ( .A(n11893), .B(n11894), .Z(n11892) );
  XOR U11804 ( .A(n11891), .B(n11895), .Z(n11893) );
  XNOR U11805 ( .A(n11784), .B(n11873), .Z(n11875) );
  XOR U11806 ( .A(n11896), .B(n11897), .Z(n11784) );
  AND U11807 ( .A(n207), .B(n11898), .Z(n11897) );
  XNOR U11808 ( .A(n11899), .B(n11896), .Z(n11898) );
  XOR U11809 ( .A(n11900), .B(n11901), .Z(n11873) );
  AND U11810 ( .A(n11902), .B(n11903), .Z(n11901) );
  XNOR U11811 ( .A(n11900), .B(n11889), .Z(n11903) );
  IV U11812 ( .A(n11835), .Z(n11889) );
  XNOR U11813 ( .A(n11904), .B(n11882), .Z(n11835) );
  XNOR U11814 ( .A(n11905), .B(n11888), .Z(n11882) );
  XOR U11815 ( .A(n11906), .B(n11907), .Z(n11888) );
  NOR U11816 ( .A(n11908), .B(n11909), .Z(n11907) );
  XNOR U11817 ( .A(n11906), .B(n11910), .Z(n11908) );
  XNOR U11818 ( .A(n11887), .B(n11879), .Z(n11905) );
  XOR U11819 ( .A(n11911), .B(n11912), .Z(n11879) );
  AND U11820 ( .A(n11913), .B(n11914), .Z(n11912) );
  XNOR U11821 ( .A(n11911), .B(n11915), .Z(n11913) );
  XNOR U11822 ( .A(n11916), .B(n11884), .Z(n11887) );
  XOR U11823 ( .A(n11917), .B(n11918), .Z(n11884) );
  AND U11824 ( .A(n11919), .B(n11920), .Z(n11918) );
  XOR U11825 ( .A(n11917), .B(n11921), .Z(n11919) );
  XNOR U11826 ( .A(n11922), .B(n11923), .Z(n11916) );
  NOR U11827 ( .A(n11924), .B(n11925), .Z(n11923) );
  XOR U11828 ( .A(n11922), .B(n11926), .Z(n11924) );
  XNOR U11829 ( .A(n11883), .B(n11890), .Z(n11904) );
  NOR U11830 ( .A(n11847), .B(n11927), .Z(n11890) );
  XOR U11831 ( .A(n11895), .B(n11894), .Z(n11883) );
  XNOR U11832 ( .A(n11928), .B(n11891), .Z(n11894) );
  XOR U11833 ( .A(n11929), .B(n11930), .Z(n11891) );
  AND U11834 ( .A(n11931), .B(n11932), .Z(n11930) );
  XOR U11835 ( .A(n11929), .B(n11933), .Z(n11931) );
  XNOR U11836 ( .A(n11934), .B(n11935), .Z(n11928) );
  NOR U11837 ( .A(n11936), .B(n11937), .Z(n11935) );
  XNOR U11838 ( .A(n11934), .B(n11938), .Z(n11936) );
  XOR U11839 ( .A(n11939), .B(n11940), .Z(n11895) );
  NOR U11840 ( .A(n11941), .B(n11942), .Z(n11940) );
  XNOR U11841 ( .A(n11939), .B(n11943), .Z(n11941) );
  XNOR U11842 ( .A(n11832), .B(n11900), .Z(n11902) );
  XOR U11843 ( .A(n11944), .B(n11945), .Z(n11832) );
  AND U11844 ( .A(n207), .B(n11946), .Z(n11945) );
  XOR U11845 ( .A(n11947), .B(n11944), .Z(n11946) );
  AND U11846 ( .A(n11844), .B(n11847), .Z(n11900) );
  XOR U11847 ( .A(n11948), .B(n11927), .Z(n11847) );
  XNOR U11848 ( .A(p_input[2048]), .B(p_input[800]), .Z(n11927) );
  XOR U11849 ( .A(n11915), .B(n11914), .Z(n11948) );
  XNOR U11850 ( .A(n11949), .B(n11921), .Z(n11914) );
  XNOR U11851 ( .A(n11910), .B(n11909), .Z(n11921) );
  XOR U11852 ( .A(n11950), .B(n11906), .Z(n11909) );
  XNOR U11853 ( .A(n6439), .B(p_input[810]), .Z(n11906) );
  XNOR U11854 ( .A(p_input[2059]), .B(p_input[811]), .Z(n11950) );
  XOR U11855 ( .A(p_input[2060]), .B(p_input[812]), .Z(n11910) );
  XNOR U11856 ( .A(n11920), .B(n11911), .Z(n11949) );
  XNOR U11857 ( .A(n6553), .B(p_input[801]), .Z(n11911) );
  XOR U11858 ( .A(n11951), .B(n11926), .Z(n11920) );
  XNOR U11859 ( .A(p_input[2063]), .B(p_input[815]), .Z(n11926) );
  XOR U11860 ( .A(n11917), .B(n11925), .Z(n11951) );
  XOR U11861 ( .A(n11952), .B(n11922), .Z(n11925) );
  XOR U11862 ( .A(p_input[2061]), .B(p_input[813]), .Z(n11922) );
  XNOR U11863 ( .A(p_input[2062]), .B(p_input[814]), .Z(n11952) );
  XNOR U11864 ( .A(n6325), .B(p_input[809]), .Z(n11917) );
  XNOR U11865 ( .A(n11933), .B(n11932), .Z(n11915) );
  XNOR U11866 ( .A(n11953), .B(n11938), .Z(n11932) );
  XOR U11867 ( .A(p_input[2056]), .B(p_input[808]), .Z(n11938) );
  XOR U11868 ( .A(n11929), .B(n11937), .Z(n11953) );
  XOR U11869 ( .A(n11954), .B(n11934), .Z(n11937) );
  XOR U11870 ( .A(p_input[2054]), .B(p_input[806]), .Z(n11934) );
  XNOR U11871 ( .A(p_input[2055]), .B(p_input[807]), .Z(n11954) );
  XNOR U11872 ( .A(n6328), .B(p_input[802]), .Z(n11929) );
  XNOR U11873 ( .A(n11943), .B(n11942), .Z(n11933) );
  XOR U11874 ( .A(n11955), .B(n11939), .Z(n11942) );
  XOR U11875 ( .A(p_input[2051]), .B(p_input[803]), .Z(n11939) );
  XNOR U11876 ( .A(p_input[2052]), .B(p_input[804]), .Z(n11955) );
  XOR U11877 ( .A(p_input[2053]), .B(p_input[805]), .Z(n11943) );
  XOR U11878 ( .A(n11956), .B(n11957), .Z(n11844) );
  AND U11879 ( .A(n207), .B(n11958), .Z(n11957) );
  XNOR U11880 ( .A(n11959), .B(n11956), .Z(n11958) );
  XNOR U11881 ( .A(n11960), .B(n11961), .Z(n207) );
  AND U11882 ( .A(n11962), .B(n11963), .Z(n11961) );
  XOR U11883 ( .A(n11857), .B(n11960), .Z(n11963) );
  AND U11884 ( .A(n11964), .B(n11965), .Z(n11857) );
  XNOR U11885 ( .A(n11854), .B(n11960), .Z(n11962) );
  XOR U11886 ( .A(n11966), .B(n11967), .Z(n11854) );
  AND U11887 ( .A(n211), .B(n11968), .Z(n11967) );
  XOR U11888 ( .A(n11969), .B(n11966), .Z(n11968) );
  XOR U11889 ( .A(n11970), .B(n11971), .Z(n11960) );
  AND U11890 ( .A(n11972), .B(n11973), .Z(n11971) );
  XNOR U11891 ( .A(n11970), .B(n11964), .Z(n11973) );
  IV U11892 ( .A(n11872), .Z(n11964) );
  XOR U11893 ( .A(n11974), .B(n11975), .Z(n11872) );
  XOR U11894 ( .A(n11976), .B(n11965), .Z(n11975) );
  AND U11895 ( .A(n11899), .B(n11977), .Z(n11965) );
  AND U11896 ( .A(n11978), .B(n11979), .Z(n11976) );
  XOR U11897 ( .A(n11980), .B(n11974), .Z(n11978) );
  XNOR U11898 ( .A(n11869), .B(n11970), .Z(n11972) );
  XOR U11899 ( .A(n11981), .B(n11982), .Z(n11869) );
  AND U11900 ( .A(n211), .B(n11983), .Z(n11982) );
  XOR U11901 ( .A(n11984), .B(n11981), .Z(n11983) );
  XOR U11902 ( .A(n11985), .B(n11986), .Z(n11970) );
  AND U11903 ( .A(n11987), .B(n11988), .Z(n11986) );
  XNOR U11904 ( .A(n11985), .B(n11899), .Z(n11988) );
  XOR U11905 ( .A(n11989), .B(n11979), .Z(n11899) );
  XNOR U11906 ( .A(n11990), .B(n11974), .Z(n11979) );
  XOR U11907 ( .A(n11991), .B(n11992), .Z(n11974) );
  AND U11908 ( .A(n11993), .B(n11994), .Z(n11992) );
  XOR U11909 ( .A(n11995), .B(n11991), .Z(n11993) );
  XNOR U11910 ( .A(n11996), .B(n11997), .Z(n11990) );
  AND U11911 ( .A(n11998), .B(n11999), .Z(n11997) );
  XOR U11912 ( .A(n11996), .B(n12000), .Z(n11998) );
  XNOR U11913 ( .A(n11980), .B(n11977), .Z(n11989) );
  AND U11914 ( .A(n12001), .B(n12002), .Z(n11977) );
  XOR U11915 ( .A(n12003), .B(n12004), .Z(n11980) );
  AND U11916 ( .A(n12005), .B(n12006), .Z(n12004) );
  XOR U11917 ( .A(n12003), .B(n12007), .Z(n12005) );
  XNOR U11918 ( .A(n11896), .B(n11985), .Z(n11987) );
  XOR U11919 ( .A(n12008), .B(n12009), .Z(n11896) );
  AND U11920 ( .A(n211), .B(n12010), .Z(n12009) );
  XNOR U11921 ( .A(n12011), .B(n12008), .Z(n12010) );
  XOR U11922 ( .A(n12012), .B(n12013), .Z(n11985) );
  AND U11923 ( .A(n12014), .B(n12015), .Z(n12013) );
  XNOR U11924 ( .A(n12012), .B(n12001), .Z(n12015) );
  IV U11925 ( .A(n11947), .Z(n12001) );
  XNOR U11926 ( .A(n12016), .B(n11994), .Z(n11947) );
  XNOR U11927 ( .A(n12017), .B(n12000), .Z(n11994) );
  XOR U11928 ( .A(n12018), .B(n12019), .Z(n12000) );
  NOR U11929 ( .A(n12020), .B(n12021), .Z(n12019) );
  XNOR U11930 ( .A(n12018), .B(n12022), .Z(n12020) );
  XNOR U11931 ( .A(n11999), .B(n11991), .Z(n12017) );
  XOR U11932 ( .A(n12023), .B(n12024), .Z(n11991) );
  AND U11933 ( .A(n12025), .B(n12026), .Z(n12024) );
  XNOR U11934 ( .A(n12023), .B(n12027), .Z(n12025) );
  XNOR U11935 ( .A(n12028), .B(n11996), .Z(n11999) );
  XOR U11936 ( .A(n12029), .B(n12030), .Z(n11996) );
  AND U11937 ( .A(n12031), .B(n12032), .Z(n12030) );
  XOR U11938 ( .A(n12029), .B(n12033), .Z(n12031) );
  XNOR U11939 ( .A(n12034), .B(n12035), .Z(n12028) );
  NOR U11940 ( .A(n12036), .B(n12037), .Z(n12035) );
  XOR U11941 ( .A(n12034), .B(n12038), .Z(n12036) );
  XNOR U11942 ( .A(n11995), .B(n12002), .Z(n12016) );
  NOR U11943 ( .A(n11959), .B(n12039), .Z(n12002) );
  XOR U11944 ( .A(n12007), .B(n12006), .Z(n11995) );
  XNOR U11945 ( .A(n12040), .B(n12003), .Z(n12006) );
  XOR U11946 ( .A(n12041), .B(n12042), .Z(n12003) );
  AND U11947 ( .A(n12043), .B(n12044), .Z(n12042) );
  XOR U11948 ( .A(n12041), .B(n12045), .Z(n12043) );
  XNOR U11949 ( .A(n12046), .B(n12047), .Z(n12040) );
  NOR U11950 ( .A(n12048), .B(n12049), .Z(n12047) );
  XNOR U11951 ( .A(n12046), .B(n12050), .Z(n12048) );
  XOR U11952 ( .A(n12051), .B(n12052), .Z(n12007) );
  NOR U11953 ( .A(n12053), .B(n12054), .Z(n12052) );
  XNOR U11954 ( .A(n12051), .B(n12055), .Z(n12053) );
  XNOR U11955 ( .A(n11944), .B(n12012), .Z(n12014) );
  XOR U11956 ( .A(n12056), .B(n12057), .Z(n11944) );
  AND U11957 ( .A(n211), .B(n12058), .Z(n12057) );
  XOR U11958 ( .A(n12059), .B(n12056), .Z(n12058) );
  AND U11959 ( .A(n11956), .B(n11959), .Z(n12012) );
  XOR U11960 ( .A(n12060), .B(n12039), .Z(n11959) );
  XNOR U11961 ( .A(p_input[2048]), .B(p_input[816]), .Z(n12039) );
  XOR U11962 ( .A(n12027), .B(n12026), .Z(n12060) );
  XNOR U11963 ( .A(n12061), .B(n12033), .Z(n12026) );
  XNOR U11964 ( .A(n12022), .B(n12021), .Z(n12033) );
  XOR U11965 ( .A(n12062), .B(n12018), .Z(n12021) );
  XNOR U11966 ( .A(n6439), .B(p_input[826]), .Z(n12018) );
  XNOR U11967 ( .A(p_input[2059]), .B(p_input[827]), .Z(n12062) );
  XOR U11968 ( .A(p_input[2060]), .B(p_input[828]), .Z(n12022) );
  XNOR U11969 ( .A(n12032), .B(n12023), .Z(n12061) );
  XNOR U11970 ( .A(n6553), .B(p_input[817]), .Z(n12023) );
  XOR U11971 ( .A(n12063), .B(n12038), .Z(n12032) );
  XNOR U11972 ( .A(p_input[2063]), .B(p_input[831]), .Z(n12038) );
  XOR U11973 ( .A(n12029), .B(n12037), .Z(n12063) );
  XOR U11974 ( .A(n12064), .B(n12034), .Z(n12037) );
  XOR U11975 ( .A(p_input[2061]), .B(p_input[829]), .Z(n12034) );
  XNOR U11976 ( .A(p_input[2062]), .B(p_input[830]), .Z(n12064) );
  XNOR U11977 ( .A(n6325), .B(p_input[825]), .Z(n12029) );
  XNOR U11978 ( .A(n12045), .B(n12044), .Z(n12027) );
  XNOR U11979 ( .A(n12065), .B(n12050), .Z(n12044) );
  XOR U11980 ( .A(p_input[2056]), .B(p_input[824]), .Z(n12050) );
  XOR U11981 ( .A(n12041), .B(n12049), .Z(n12065) );
  XOR U11982 ( .A(n12066), .B(n12046), .Z(n12049) );
  XOR U11983 ( .A(p_input[2054]), .B(p_input[822]), .Z(n12046) );
  XNOR U11984 ( .A(p_input[2055]), .B(p_input[823]), .Z(n12066) );
  XNOR U11985 ( .A(n6328), .B(p_input[818]), .Z(n12041) );
  XNOR U11986 ( .A(n12055), .B(n12054), .Z(n12045) );
  XOR U11987 ( .A(n12067), .B(n12051), .Z(n12054) );
  XOR U11988 ( .A(p_input[2051]), .B(p_input[819]), .Z(n12051) );
  XNOR U11989 ( .A(p_input[2052]), .B(p_input[820]), .Z(n12067) );
  XOR U11990 ( .A(p_input[2053]), .B(p_input[821]), .Z(n12055) );
  XOR U11991 ( .A(n12068), .B(n12069), .Z(n11956) );
  AND U11992 ( .A(n211), .B(n12070), .Z(n12069) );
  XNOR U11993 ( .A(n12071), .B(n12068), .Z(n12070) );
  XNOR U11994 ( .A(n12072), .B(n12073), .Z(n211) );
  AND U11995 ( .A(n12074), .B(n12075), .Z(n12073) );
  XOR U11996 ( .A(n11969), .B(n12072), .Z(n12075) );
  AND U11997 ( .A(n12076), .B(n12077), .Z(n11969) );
  XNOR U11998 ( .A(n11966), .B(n12072), .Z(n12074) );
  XOR U11999 ( .A(n12078), .B(n12079), .Z(n11966) );
  AND U12000 ( .A(n215), .B(n12080), .Z(n12079) );
  XOR U12001 ( .A(n12081), .B(n12078), .Z(n12080) );
  XOR U12002 ( .A(n12082), .B(n12083), .Z(n12072) );
  AND U12003 ( .A(n12084), .B(n12085), .Z(n12083) );
  XNOR U12004 ( .A(n12082), .B(n12076), .Z(n12085) );
  IV U12005 ( .A(n11984), .Z(n12076) );
  XOR U12006 ( .A(n12086), .B(n12087), .Z(n11984) );
  XOR U12007 ( .A(n12088), .B(n12077), .Z(n12087) );
  AND U12008 ( .A(n12011), .B(n12089), .Z(n12077) );
  AND U12009 ( .A(n12090), .B(n12091), .Z(n12088) );
  XOR U12010 ( .A(n12092), .B(n12086), .Z(n12090) );
  XNOR U12011 ( .A(n11981), .B(n12082), .Z(n12084) );
  XOR U12012 ( .A(n12093), .B(n12094), .Z(n11981) );
  AND U12013 ( .A(n215), .B(n12095), .Z(n12094) );
  XOR U12014 ( .A(n12096), .B(n12093), .Z(n12095) );
  XOR U12015 ( .A(n12097), .B(n12098), .Z(n12082) );
  AND U12016 ( .A(n12099), .B(n12100), .Z(n12098) );
  XNOR U12017 ( .A(n12097), .B(n12011), .Z(n12100) );
  XOR U12018 ( .A(n12101), .B(n12091), .Z(n12011) );
  XNOR U12019 ( .A(n12102), .B(n12086), .Z(n12091) );
  XOR U12020 ( .A(n12103), .B(n12104), .Z(n12086) );
  AND U12021 ( .A(n12105), .B(n12106), .Z(n12104) );
  XOR U12022 ( .A(n12107), .B(n12103), .Z(n12105) );
  XNOR U12023 ( .A(n12108), .B(n12109), .Z(n12102) );
  AND U12024 ( .A(n12110), .B(n12111), .Z(n12109) );
  XOR U12025 ( .A(n12108), .B(n12112), .Z(n12110) );
  XNOR U12026 ( .A(n12092), .B(n12089), .Z(n12101) );
  AND U12027 ( .A(n12113), .B(n12114), .Z(n12089) );
  XOR U12028 ( .A(n12115), .B(n12116), .Z(n12092) );
  AND U12029 ( .A(n12117), .B(n12118), .Z(n12116) );
  XOR U12030 ( .A(n12115), .B(n12119), .Z(n12117) );
  XNOR U12031 ( .A(n12008), .B(n12097), .Z(n12099) );
  XOR U12032 ( .A(n12120), .B(n12121), .Z(n12008) );
  AND U12033 ( .A(n215), .B(n12122), .Z(n12121) );
  XNOR U12034 ( .A(n12123), .B(n12120), .Z(n12122) );
  XOR U12035 ( .A(n12124), .B(n12125), .Z(n12097) );
  AND U12036 ( .A(n12126), .B(n12127), .Z(n12125) );
  XNOR U12037 ( .A(n12124), .B(n12113), .Z(n12127) );
  IV U12038 ( .A(n12059), .Z(n12113) );
  XNOR U12039 ( .A(n12128), .B(n12106), .Z(n12059) );
  XNOR U12040 ( .A(n12129), .B(n12112), .Z(n12106) );
  XOR U12041 ( .A(n12130), .B(n12131), .Z(n12112) );
  NOR U12042 ( .A(n12132), .B(n12133), .Z(n12131) );
  XNOR U12043 ( .A(n12130), .B(n12134), .Z(n12132) );
  XNOR U12044 ( .A(n12111), .B(n12103), .Z(n12129) );
  XOR U12045 ( .A(n12135), .B(n12136), .Z(n12103) );
  AND U12046 ( .A(n12137), .B(n12138), .Z(n12136) );
  XNOR U12047 ( .A(n12135), .B(n12139), .Z(n12137) );
  XNOR U12048 ( .A(n12140), .B(n12108), .Z(n12111) );
  XOR U12049 ( .A(n12141), .B(n12142), .Z(n12108) );
  AND U12050 ( .A(n12143), .B(n12144), .Z(n12142) );
  XOR U12051 ( .A(n12141), .B(n12145), .Z(n12143) );
  XNOR U12052 ( .A(n12146), .B(n12147), .Z(n12140) );
  NOR U12053 ( .A(n12148), .B(n12149), .Z(n12147) );
  XOR U12054 ( .A(n12146), .B(n12150), .Z(n12148) );
  XNOR U12055 ( .A(n12107), .B(n12114), .Z(n12128) );
  NOR U12056 ( .A(n12071), .B(n12151), .Z(n12114) );
  XOR U12057 ( .A(n12119), .B(n12118), .Z(n12107) );
  XNOR U12058 ( .A(n12152), .B(n12115), .Z(n12118) );
  XOR U12059 ( .A(n12153), .B(n12154), .Z(n12115) );
  AND U12060 ( .A(n12155), .B(n12156), .Z(n12154) );
  XOR U12061 ( .A(n12153), .B(n12157), .Z(n12155) );
  XNOR U12062 ( .A(n12158), .B(n12159), .Z(n12152) );
  NOR U12063 ( .A(n12160), .B(n12161), .Z(n12159) );
  XNOR U12064 ( .A(n12158), .B(n12162), .Z(n12160) );
  XOR U12065 ( .A(n12163), .B(n12164), .Z(n12119) );
  NOR U12066 ( .A(n12165), .B(n12166), .Z(n12164) );
  XNOR U12067 ( .A(n12163), .B(n12167), .Z(n12165) );
  XNOR U12068 ( .A(n12056), .B(n12124), .Z(n12126) );
  XOR U12069 ( .A(n12168), .B(n12169), .Z(n12056) );
  AND U12070 ( .A(n215), .B(n12170), .Z(n12169) );
  XOR U12071 ( .A(n12171), .B(n12168), .Z(n12170) );
  AND U12072 ( .A(n12068), .B(n12071), .Z(n12124) );
  XOR U12073 ( .A(n12172), .B(n12151), .Z(n12071) );
  XNOR U12074 ( .A(p_input[2048]), .B(p_input[832]), .Z(n12151) );
  XOR U12075 ( .A(n12139), .B(n12138), .Z(n12172) );
  XNOR U12076 ( .A(n12173), .B(n12145), .Z(n12138) );
  XNOR U12077 ( .A(n12134), .B(n12133), .Z(n12145) );
  XOR U12078 ( .A(n12174), .B(n12130), .Z(n12133) );
  XNOR U12079 ( .A(n6439), .B(p_input[842]), .Z(n12130) );
  XNOR U12080 ( .A(p_input[2059]), .B(p_input[843]), .Z(n12174) );
  XOR U12081 ( .A(p_input[2060]), .B(p_input[844]), .Z(n12134) );
  XNOR U12082 ( .A(n12144), .B(n12135), .Z(n12173) );
  XNOR U12083 ( .A(n6553), .B(p_input[833]), .Z(n12135) );
  XOR U12084 ( .A(n12175), .B(n12150), .Z(n12144) );
  XNOR U12085 ( .A(p_input[2063]), .B(p_input[847]), .Z(n12150) );
  XOR U12086 ( .A(n12141), .B(n12149), .Z(n12175) );
  XOR U12087 ( .A(n12176), .B(n12146), .Z(n12149) );
  XOR U12088 ( .A(p_input[2061]), .B(p_input[845]), .Z(n12146) );
  XNOR U12089 ( .A(p_input[2062]), .B(p_input[846]), .Z(n12176) );
  XNOR U12090 ( .A(n6325), .B(p_input[841]), .Z(n12141) );
  XNOR U12091 ( .A(n12157), .B(n12156), .Z(n12139) );
  XNOR U12092 ( .A(n12177), .B(n12162), .Z(n12156) );
  XOR U12093 ( .A(p_input[2056]), .B(p_input[840]), .Z(n12162) );
  XOR U12094 ( .A(n12153), .B(n12161), .Z(n12177) );
  XOR U12095 ( .A(n12178), .B(n12158), .Z(n12161) );
  XOR U12096 ( .A(p_input[2054]), .B(p_input[838]), .Z(n12158) );
  XNOR U12097 ( .A(p_input[2055]), .B(p_input[839]), .Z(n12178) );
  XNOR U12098 ( .A(n6328), .B(p_input[834]), .Z(n12153) );
  XNOR U12099 ( .A(n12167), .B(n12166), .Z(n12157) );
  XOR U12100 ( .A(n12179), .B(n12163), .Z(n12166) );
  XOR U12101 ( .A(p_input[2051]), .B(p_input[835]), .Z(n12163) );
  XNOR U12102 ( .A(p_input[2052]), .B(p_input[836]), .Z(n12179) );
  XOR U12103 ( .A(p_input[2053]), .B(p_input[837]), .Z(n12167) );
  XOR U12104 ( .A(n12180), .B(n12181), .Z(n12068) );
  AND U12105 ( .A(n215), .B(n12182), .Z(n12181) );
  XNOR U12106 ( .A(n12183), .B(n12180), .Z(n12182) );
  XNOR U12107 ( .A(n12184), .B(n12185), .Z(n215) );
  AND U12108 ( .A(n12186), .B(n12187), .Z(n12185) );
  XOR U12109 ( .A(n12081), .B(n12184), .Z(n12187) );
  AND U12110 ( .A(n12188), .B(n12189), .Z(n12081) );
  XNOR U12111 ( .A(n12078), .B(n12184), .Z(n12186) );
  XOR U12112 ( .A(n12190), .B(n12191), .Z(n12078) );
  AND U12113 ( .A(n219), .B(n12192), .Z(n12191) );
  XOR U12114 ( .A(n12193), .B(n12190), .Z(n12192) );
  XOR U12115 ( .A(n12194), .B(n12195), .Z(n12184) );
  AND U12116 ( .A(n12196), .B(n12197), .Z(n12195) );
  XNOR U12117 ( .A(n12194), .B(n12188), .Z(n12197) );
  IV U12118 ( .A(n12096), .Z(n12188) );
  XOR U12119 ( .A(n12198), .B(n12199), .Z(n12096) );
  XOR U12120 ( .A(n12200), .B(n12189), .Z(n12199) );
  AND U12121 ( .A(n12123), .B(n12201), .Z(n12189) );
  AND U12122 ( .A(n12202), .B(n12203), .Z(n12200) );
  XOR U12123 ( .A(n12204), .B(n12198), .Z(n12202) );
  XNOR U12124 ( .A(n12093), .B(n12194), .Z(n12196) );
  XOR U12125 ( .A(n12205), .B(n12206), .Z(n12093) );
  AND U12126 ( .A(n219), .B(n12207), .Z(n12206) );
  XOR U12127 ( .A(n12208), .B(n12205), .Z(n12207) );
  XOR U12128 ( .A(n12209), .B(n12210), .Z(n12194) );
  AND U12129 ( .A(n12211), .B(n12212), .Z(n12210) );
  XNOR U12130 ( .A(n12209), .B(n12123), .Z(n12212) );
  XOR U12131 ( .A(n12213), .B(n12203), .Z(n12123) );
  XNOR U12132 ( .A(n12214), .B(n12198), .Z(n12203) );
  XOR U12133 ( .A(n12215), .B(n12216), .Z(n12198) );
  AND U12134 ( .A(n12217), .B(n12218), .Z(n12216) );
  XOR U12135 ( .A(n12219), .B(n12215), .Z(n12217) );
  XNOR U12136 ( .A(n12220), .B(n12221), .Z(n12214) );
  AND U12137 ( .A(n12222), .B(n12223), .Z(n12221) );
  XOR U12138 ( .A(n12220), .B(n12224), .Z(n12222) );
  XNOR U12139 ( .A(n12204), .B(n12201), .Z(n12213) );
  AND U12140 ( .A(n12225), .B(n12226), .Z(n12201) );
  XOR U12141 ( .A(n12227), .B(n12228), .Z(n12204) );
  AND U12142 ( .A(n12229), .B(n12230), .Z(n12228) );
  XOR U12143 ( .A(n12227), .B(n12231), .Z(n12229) );
  XNOR U12144 ( .A(n12120), .B(n12209), .Z(n12211) );
  XOR U12145 ( .A(n12232), .B(n12233), .Z(n12120) );
  AND U12146 ( .A(n219), .B(n12234), .Z(n12233) );
  XNOR U12147 ( .A(n12235), .B(n12232), .Z(n12234) );
  XOR U12148 ( .A(n12236), .B(n12237), .Z(n12209) );
  AND U12149 ( .A(n12238), .B(n12239), .Z(n12237) );
  XNOR U12150 ( .A(n12236), .B(n12225), .Z(n12239) );
  IV U12151 ( .A(n12171), .Z(n12225) );
  XNOR U12152 ( .A(n12240), .B(n12218), .Z(n12171) );
  XNOR U12153 ( .A(n12241), .B(n12224), .Z(n12218) );
  XOR U12154 ( .A(n12242), .B(n12243), .Z(n12224) );
  NOR U12155 ( .A(n12244), .B(n12245), .Z(n12243) );
  XNOR U12156 ( .A(n12242), .B(n12246), .Z(n12244) );
  XNOR U12157 ( .A(n12223), .B(n12215), .Z(n12241) );
  XOR U12158 ( .A(n12247), .B(n12248), .Z(n12215) );
  AND U12159 ( .A(n12249), .B(n12250), .Z(n12248) );
  XNOR U12160 ( .A(n12247), .B(n12251), .Z(n12249) );
  XNOR U12161 ( .A(n12252), .B(n12220), .Z(n12223) );
  XOR U12162 ( .A(n12253), .B(n12254), .Z(n12220) );
  AND U12163 ( .A(n12255), .B(n12256), .Z(n12254) );
  XOR U12164 ( .A(n12253), .B(n12257), .Z(n12255) );
  XNOR U12165 ( .A(n12258), .B(n12259), .Z(n12252) );
  NOR U12166 ( .A(n12260), .B(n12261), .Z(n12259) );
  XOR U12167 ( .A(n12258), .B(n12262), .Z(n12260) );
  XNOR U12168 ( .A(n12219), .B(n12226), .Z(n12240) );
  NOR U12169 ( .A(n12183), .B(n12263), .Z(n12226) );
  XOR U12170 ( .A(n12231), .B(n12230), .Z(n12219) );
  XNOR U12171 ( .A(n12264), .B(n12227), .Z(n12230) );
  XOR U12172 ( .A(n12265), .B(n12266), .Z(n12227) );
  AND U12173 ( .A(n12267), .B(n12268), .Z(n12266) );
  XOR U12174 ( .A(n12265), .B(n12269), .Z(n12267) );
  XNOR U12175 ( .A(n12270), .B(n12271), .Z(n12264) );
  NOR U12176 ( .A(n12272), .B(n12273), .Z(n12271) );
  XNOR U12177 ( .A(n12270), .B(n12274), .Z(n12272) );
  XOR U12178 ( .A(n12275), .B(n12276), .Z(n12231) );
  NOR U12179 ( .A(n12277), .B(n12278), .Z(n12276) );
  XNOR U12180 ( .A(n12275), .B(n12279), .Z(n12277) );
  XNOR U12181 ( .A(n12168), .B(n12236), .Z(n12238) );
  XOR U12182 ( .A(n12280), .B(n12281), .Z(n12168) );
  AND U12183 ( .A(n219), .B(n12282), .Z(n12281) );
  XOR U12184 ( .A(n12283), .B(n12280), .Z(n12282) );
  AND U12185 ( .A(n12180), .B(n12183), .Z(n12236) );
  XOR U12186 ( .A(n12284), .B(n12263), .Z(n12183) );
  XNOR U12187 ( .A(p_input[2048]), .B(p_input[848]), .Z(n12263) );
  XOR U12188 ( .A(n12251), .B(n12250), .Z(n12284) );
  XNOR U12189 ( .A(n12285), .B(n12257), .Z(n12250) );
  XNOR U12190 ( .A(n12246), .B(n12245), .Z(n12257) );
  XOR U12191 ( .A(n12286), .B(n12242), .Z(n12245) );
  XNOR U12192 ( .A(n6439), .B(p_input[858]), .Z(n12242) );
  XNOR U12193 ( .A(p_input[2059]), .B(p_input[859]), .Z(n12286) );
  XOR U12194 ( .A(p_input[2060]), .B(p_input[860]), .Z(n12246) );
  XNOR U12195 ( .A(n12256), .B(n12247), .Z(n12285) );
  XNOR U12196 ( .A(n6553), .B(p_input[849]), .Z(n12247) );
  XOR U12197 ( .A(n12287), .B(n12262), .Z(n12256) );
  XNOR U12198 ( .A(p_input[2063]), .B(p_input[863]), .Z(n12262) );
  XOR U12199 ( .A(n12253), .B(n12261), .Z(n12287) );
  XOR U12200 ( .A(n12288), .B(n12258), .Z(n12261) );
  XOR U12201 ( .A(p_input[2061]), .B(p_input[861]), .Z(n12258) );
  XNOR U12202 ( .A(p_input[2062]), .B(p_input[862]), .Z(n12288) );
  XNOR U12203 ( .A(n6325), .B(p_input[857]), .Z(n12253) );
  XNOR U12204 ( .A(n12269), .B(n12268), .Z(n12251) );
  XNOR U12205 ( .A(n12289), .B(n12274), .Z(n12268) );
  XOR U12206 ( .A(p_input[2056]), .B(p_input[856]), .Z(n12274) );
  XOR U12207 ( .A(n12265), .B(n12273), .Z(n12289) );
  XOR U12208 ( .A(n12290), .B(n12270), .Z(n12273) );
  XOR U12209 ( .A(p_input[2054]), .B(p_input[854]), .Z(n12270) );
  XNOR U12210 ( .A(p_input[2055]), .B(p_input[855]), .Z(n12290) );
  XNOR U12211 ( .A(n6328), .B(p_input[850]), .Z(n12265) );
  XNOR U12212 ( .A(n12279), .B(n12278), .Z(n12269) );
  XOR U12213 ( .A(n12291), .B(n12275), .Z(n12278) );
  XOR U12214 ( .A(p_input[2051]), .B(p_input[851]), .Z(n12275) );
  XNOR U12215 ( .A(p_input[2052]), .B(p_input[852]), .Z(n12291) );
  XOR U12216 ( .A(p_input[2053]), .B(p_input[853]), .Z(n12279) );
  XOR U12217 ( .A(n12292), .B(n12293), .Z(n12180) );
  AND U12218 ( .A(n219), .B(n12294), .Z(n12293) );
  XNOR U12219 ( .A(n12295), .B(n12292), .Z(n12294) );
  XNOR U12220 ( .A(n12296), .B(n12297), .Z(n219) );
  AND U12221 ( .A(n12298), .B(n12299), .Z(n12297) );
  XOR U12222 ( .A(n12193), .B(n12296), .Z(n12299) );
  AND U12223 ( .A(n12300), .B(n12301), .Z(n12193) );
  XNOR U12224 ( .A(n12190), .B(n12296), .Z(n12298) );
  XOR U12225 ( .A(n12302), .B(n12303), .Z(n12190) );
  AND U12226 ( .A(n223), .B(n12304), .Z(n12303) );
  XOR U12227 ( .A(n12305), .B(n12302), .Z(n12304) );
  XOR U12228 ( .A(n12306), .B(n12307), .Z(n12296) );
  AND U12229 ( .A(n12308), .B(n12309), .Z(n12307) );
  XNOR U12230 ( .A(n12306), .B(n12300), .Z(n12309) );
  IV U12231 ( .A(n12208), .Z(n12300) );
  XOR U12232 ( .A(n12310), .B(n12311), .Z(n12208) );
  XOR U12233 ( .A(n12312), .B(n12301), .Z(n12311) );
  AND U12234 ( .A(n12235), .B(n12313), .Z(n12301) );
  AND U12235 ( .A(n12314), .B(n12315), .Z(n12312) );
  XOR U12236 ( .A(n12316), .B(n12310), .Z(n12314) );
  XNOR U12237 ( .A(n12205), .B(n12306), .Z(n12308) );
  XOR U12238 ( .A(n12317), .B(n12318), .Z(n12205) );
  AND U12239 ( .A(n223), .B(n12319), .Z(n12318) );
  XOR U12240 ( .A(n12320), .B(n12317), .Z(n12319) );
  XOR U12241 ( .A(n12321), .B(n12322), .Z(n12306) );
  AND U12242 ( .A(n12323), .B(n12324), .Z(n12322) );
  XNOR U12243 ( .A(n12321), .B(n12235), .Z(n12324) );
  XOR U12244 ( .A(n12325), .B(n12315), .Z(n12235) );
  XNOR U12245 ( .A(n12326), .B(n12310), .Z(n12315) );
  XOR U12246 ( .A(n12327), .B(n12328), .Z(n12310) );
  AND U12247 ( .A(n12329), .B(n12330), .Z(n12328) );
  XOR U12248 ( .A(n12331), .B(n12327), .Z(n12329) );
  XNOR U12249 ( .A(n12332), .B(n12333), .Z(n12326) );
  AND U12250 ( .A(n12334), .B(n12335), .Z(n12333) );
  XOR U12251 ( .A(n12332), .B(n12336), .Z(n12334) );
  XNOR U12252 ( .A(n12316), .B(n12313), .Z(n12325) );
  AND U12253 ( .A(n12337), .B(n12338), .Z(n12313) );
  XOR U12254 ( .A(n12339), .B(n12340), .Z(n12316) );
  AND U12255 ( .A(n12341), .B(n12342), .Z(n12340) );
  XOR U12256 ( .A(n12339), .B(n12343), .Z(n12341) );
  XNOR U12257 ( .A(n12232), .B(n12321), .Z(n12323) );
  XOR U12258 ( .A(n12344), .B(n12345), .Z(n12232) );
  AND U12259 ( .A(n223), .B(n12346), .Z(n12345) );
  XNOR U12260 ( .A(n12347), .B(n12344), .Z(n12346) );
  XOR U12261 ( .A(n12348), .B(n12349), .Z(n12321) );
  AND U12262 ( .A(n12350), .B(n12351), .Z(n12349) );
  XNOR U12263 ( .A(n12348), .B(n12337), .Z(n12351) );
  IV U12264 ( .A(n12283), .Z(n12337) );
  XNOR U12265 ( .A(n12352), .B(n12330), .Z(n12283) );
  XNOR U12266 ( .A(n12353), .B(n12336), .Z(n12330) );
  XOR U12267 ( .A(n12354), .B(n12355), .Z(n12336) );
  NOR U12268 ( .A(n12356), .B(n12357), .Z(n12355) );
  XNOR U12269 ( .A(n12354), .B(n12358), .Z(n12356) );
  XNOR U12270 ( .A(n12335), .B(n12327), .Z(n12353) );
  XOR U12271 ( .A(n12359), .B(n12360), .Z(n12327) );
  AND U12272 ( .A(n12361), .B(n12362), .Z(n12360) );
  XNOR U12273 ( .A(n12359), .B(n12363), .Z(n12361) );
  XNOR U12274 ( .A(n12364), .B(n12332), .Z(n12335) );
  XOR U12275 ( .A(n12365), .B(n12366), .Z(n12332) );
  AND U12276 ( .A(n12367), .B(n12368), .Z(n12366) );
  XOR U12277 ( .A(n12365), .B(n12369), .Z(n12367) );
  XNOR U12278 ( .A(n12370), .B(n12371), .Z(n12364) );
  NOR U12279 ( .A(n12372), .B(n12373), .Z(n12371) );
  XOR U12280 ( .A(n12370), .B(n12374), .Z(n12372) );
  XNOR U12281 ( .A(n12331), .B(n12338), .Z(n12352) );
  NOR U12282 ( .A(n12295), .B(n12375), .Z(n12338) );
  XOR U12283 ( .A(n12343), .B(n12342), .Z(n12331) );
  XNOR U12284 ( .A(n12376), .B(n12339), .Z(n12342) );
  XOR U12285 ( .A(n12377), .B(n12378), .Z(n12339) );
  AND U12286 ( .A(n12379), .B(n12380), .Z(n12378) );
  XOR U12287 ( .A(n12377), .B(n12381), .Z(n12379) );
  XNOR U12288 ( .A(n12382), .B(n12383), .Z(n12376) );
  NOR U12289 ( .A(n12384), .B(n12385), .Z(n12383) );
  XNOR U12290 ( .A(n12382), .B(n12386), .Z(n12384) );
  XOR U12291 ( .A(n12387), .B(n12388), .Z(n12343) );
  NOR U12292 ( .A(n12389), .B(n12390), .Z(n12388) );
  XNOR U12293 ( .A(n12387), .B(n12391), .Z(n12389) );
  XNOR U12294 ( .A(n12280), .B(n12348), .Z(n12350) );
  XOR U12295 ( .A(n12392), .B(n12393), .Z(n12280) );
  AND U12296 ( .A(n223), .B(n12394), .Z(n12393) );
  XOR U12297 ( .A(n12395), .B(n12392), .Z(n12394) );
  AND U12298 ( .A(n12292), .B(n12295), .Z(n12348) );
  XOR U12299 ( .A(n12396), .B(n12375), .Z(n12295) );
  XNOR U12300 ( .A(p_input[2048]), .B(p_input[864]), .Z(n12375) );
  XOR U12301 ( .A(n12363), .B(n12362), .Z(n12396) );
  XNOR U12302 ( .A(n12397), .B(n12369), .Z(n12362) );
  XNOR U12303 ( .A(n12358), .B(n12357), .Z(n12369) );
  XOR U12304 ( .A(n12398), .B(n12354), .Z(n12357) );
  XNOR U12305 ( .A(n6439), .B(p_input[874]), .Z(n12354) );
  XNOR U12306 ( .A(p_input[2059]), .B(p_input[875]), .Z(n12398) );
  XOR U12307 ( .A(p_input[2060]), .B(p_input[876]), .Z(n12358) );
  XNOR U12308 ( .A(n12368), .B(n12359), .Z(n12397) );
  XNOR U12309 ( .A(n6553), .B(p_input[865]), .Z(n12359) );
  XOR U12310 ( .A(n12399), .B(n12374), .Z(n12368) );
  XNOR U12311 ( .A(p_input[2063]), .B(p_input[879]), .Z(n12374) );
  XOR U12312 ( .A(n12365), .B(n12373), .Z(n12399) );
  XOR U12313 ( .A(n12400), .B(n12370), .Z(n12373) );
  XOR U12314 ( .A(p_input[2061]), .B(p_input[877]), .Z(n12370) );
  XNOR U12315 ( .A(p_input[2062]), .B(p_input[878]), .Z(n12400) );
  XNOR U12316 ( .A(n6325), .B(p_input[873]), .Z(n12365) );
  XNOR U12317 ( .A(n12381), .B(n12380), .Z(n12363) );
  XNOR U12318 ( .A(n12401), .B(n12386), .Z(n12380) );
  XOR U12319 ( .A(p_input[2056]), .B(p_input[872]), .Z(n12386) );
  XOR U12320 ( .A(n12377), .B(n12385), .Z(n12401) );
  XOR U12321 ( .A(n12402), .B(n12382), .Z(n12385) );
  XOR U12322 ( .A(p_input[2054]), .B(p_input[870]), .Z(n12382) );
  XNOR U12323 ( .A(p_input[2055]), .B(p_input[871]), .Z(n12402) );
  XNOR U12324 ( .A(n6328), .B(p_input[866]), .Z(n12377) );
  XNOR U12325 ( .A(n12391), .B(n12390), .Z(n12381) );
  XOR U12326 ( .A(n12403), .B(n12387), .Z(n12390) );
  XOR U12327 ( .A(p_input[2051]), .B(p_input[867]), .Z(n12387) );
  XNOR U12328 ( .A(p_input[2052]), .B(p_input[868]), .Z(n12403) );
  XOR U12329 ( .A(p_input[2053]), .B(p_input[869]), .Z(n12391) );
  XOR U12330 ( .A(n12404), .B(n12405), .Z(n12292) );
  AND U12331 ( .A(n223), .B(n12406), .Z(n12405) );
  XNOR U12332 ( .A(n12407), .B(n12404), .Z(n12406) );
  XNOR U12333 ( .A(n12408), .B(n12409), .Z(n223) );
  AND U12334 ( .A(n12410), .B(n12411), .Z(n12409) );
  XOR U12335 ( .A(n12305), .B(n12408), .Z(n12411) );
  AND U12336 ( .A(n12412), .B(n12413), .Z(n12305) );
  XNOR U12337 ( .A(n12302), .B(n12408), .Z(n12410) );
  XOR U12338 ( .A(n12414), .B(n12415), .Z(n12302) );
  AND U12339 ( .A(n227), .B(n12416), .Z(n12415) );
  XOR U12340 ( .A(n12417), .B(n12414), .Z(n12416) );
  XOR U12341 ( .A(n12418), .B(n12419), .Z(n12408) );
  AND U12342 ( .A(n12420), .B(n12421), .Z(n12419) );
  XNOR U12343 ( .A(n12418), .B(n12412), .Z(n12421) );
  IV U12344 ( .A(n12320), .Z(n12412) );
  XOR U12345 ( .A(n12422), .B(n12423), .Z(n12320) );
  XOR U12346 ( .A(n12424), .B(n12413), .Z(n12423) );
  AND U12347 ( .A(n12347), .B(n12425), .Z(n12413) );
  AND U12348 ( .A(n12426), .B(n12427), .Z(n12424) );
  XOR U12349 ( .A(n12428), .B(n12422), .Z(n12426) );
  XNOR U12350 ( .A(n12317), .B(n12418), .Z(n12420) );
  XOR U12351 ( .A(n12429), .B(n12430), .Z(n12317) );
  AND U12352 ( .A(n227), .B(n12431), .Z(n12430) );
  XOR U12353 ( .A(n12432), .B(n12429), .Z(n12431) );
  XOR U12354 ( .A(n12433), .B(n12434), .Z(n12418) );
  AND U12355 ( .A(n12435), .B(n12436), .Z(n12434) );
  XNOR U12356 ( .A(n12433), .B(n12347), .Z(n12436) );
  XOR U12357 ( .A(n12437), .B(n12427), .Z(n12347) );
  XNOR U12358 ( .A(n12438), .B(n12422), .Z(n12427) );
  XOR U12359 ( .A(n12439), .B(n12440), .Z(n12422) );
  AND U12360 ( .A(n12441), .B(n12442), .Z(n12440) );
  XOR U12361 ( .A(n12443), .B(n12439), .Z(n12441) );
  XNOR U12362 ( .A(n12444), .B(n12445), .Z(n12438) );
  AND U12363 ( .A(n12446), .B(n12447), .Z(n12445) );
  XOR U12364 ( .A(n12444), .B(n12448), .Z(n12446) );
  XNOR U12365 ( .A(n12428), .B(n12425), .Z(n12437) );
  AND U12366 ( .A(n12449), .B(n12450), .Z(n12425) );
  XOR U12367 ( .A(n12451), .B(n12452), .Z(n12428) );
  AND U12368 ( .A(n12453), .B(n12454), .Z(n12452) );
  XOR U12369 ( .A(n12451), .B(n12455), .Z(n12453) );
  XNOR U12370 ( .A(n12344), .B(n12433), .Z(n12435) );
  XOR U12371 ( .A(n12456), .B(n12457), .Z(n12344) );
  AND U12372 ( .A(n227), .B(n12458), .Z(n12457) );
  XNOR U12373 ( .A(n12459), .B(n12456), .Z(n12458) );
  XOR U12374 ( .A(n12460), .B(n12461), .Z(n12433) );
  AND U12375 ( .A(n12462), .B(n12463), .Z(n12461) );
  XNOR U12376 ( .A(n12460), .B(n12449), .Z(n12463) );
  IV U12377 ( .A(n12395), .Z(n12449) );
  XNOR U12378 ( .A(n12464), .B(n12442), .Z(n12395) );
  XNOR U12379 ( .A(n12465), .B(n12448), .Z(n12442) );
  XOR U12380 ( .A(n12466), .B(n12467), .Z(n12448) );
  NOR U12381 ( .A(n12468), .B(n12469), .Z(n12467) );
  XNOR U12382 ( .A(n12466), .B(n12470), .Z(n12468) );
  XNOR U12383 ( .A(n12447), .B(n12439), .Z(n12465) );
  XOR U12384 ( .A(n12471), .B(n12472), .Z(n12439) );
  AND U12385 ( .A(n12473), .B(n12474), .Z(n12472) );
  XNOR U12386 ( .A(n12471), .B(n12475), .Z(n12473) );
  XNOR U12387 ( .A(n12476), .B(n12444), .Z(n12447) );
  XOR U12388 ( .A(n12477), .B(n12478), .Z(n12444) );
  AND U12389 ( .A(n12479), .B(n12480), .Z(n12478) );
  XOR U12390 ( .A(n12477), .B(n12481), .Z(n12479) );
  XNOR U12391 ( .A(n12482), .B(n12483), .Z(n12476) );
  NOR U12392 ( .A(n12484), .B(n12485), .Z(n12483) );
  XOR U12393 ( .A(n12482), .B(n12486), .Z(n12484) );
  XNOR U12394 ( .A(n12443), .B(n12450), .Z(n12464) );
  NOR U12395 ( .A(n12407), .B(n12487), .Z(n12450) );
  XOR U12396 ( .A(n12455), .B(n12454), .Z(n12443) );
  XNOR U12397 ( .A(n12488), .B(n12451), .Z(n12454) );
  XOR U12398 ( .A(n12489), .B(n12490), .Z(n12451) );
  AND U12399 ( .A(n12491), .B(n12492), .Z(n12490) );
  XOR U12400 ( .A(n12489), .B(n12493), .Z(n12491) );
  XNOR U12401 ( .A(n12494), .B(n12495), .Z(n12488) );
  NOR U12402 ( .A(n12496), .B(n12497), .Z(n12495) );
  XNOR U12403 ( .A(n12494), .B(n12498), .Z(n12496) );
  XOR U12404 ( .A(n12499), .B(n12500), .Z(n12455) );
  NOR U12405 ( .A(n12501), .B(n12502), .Z(n12500) );
  XNOR U12406 ( .A(n12499), .B(n12503), .Z(n12501) );
  XNOR U12407 ( .A(n12392), .B(n12460), .Z(n12462) );
  XOR U12408 ( .A(n12504), .B(n12505), .Z(n12392) );
  AND U12409 ( .A(n227), .B(n12506), .Z(n12505) );
  XOR U12410 ( .A(n12507), .B(n12504), .Z(n12506) );
  AND U12411 ( .A(n12404), .B(n12407), .Z(n12460) );
  XOR U12412 ( .A(n12508), .B(n12487), .Z(n12407) );
  XNOR U12413 ( .A(p_input[2048]), .B(p_input[880]), .Z(n12487) );
  XOR U12414 ( .A(n12475), .B(n12474), .Z(n12508) );
  XNOR U12415 ( .A(n12509), .B(n12481), .Z(n12474) );
  XNOR U12416 ( .A(n12470), .B(n12469), .Z(n12481) );
  XOR U12417 ( .A(n12510), .B(n12466), .Z(n12469) );
  XNOR U12418 ( .A(n6439), .B(p_input[890]), .Z(n12466) );
  XNOR U12419 ( .A(p_input[2059]), .B(p_input[891]), .Z(n12510) );
  XOR U12420 ( .A(p_input[2060]), .B(p_input[892]), .Z(n12470) );
  XNOR U12421 ( .A(n12480), .B(n12471), .Z(n12509) );
  XNOR U12422 ( .A(n6553), .B(p_input[881]), .Z(n12471) );
  XOR U12423 ( .A(n12511), .B(n12486), .Z(n12480) );
  XNOR U12424 ( .A(p_input[2063]), .B(p_input[895]), .Z(n12486) );
  XOR U12425 ( .A(n12477), .B(n12485), .Z(n12511) );
  XOR U12426 ( .A(n12512), .B(n12482), .Z(n12485) );
  XOR U12427 ( .A(p_input[2061]), .B(p_input[893]), .Z(n12482) );
  XNOR U12428 ( .A(p_input[2062]), .B(p_input[894]), .Z(n12512) );
  XNOR U12429 ( .A(n6325), .B(p_input[889]), .Z(n12477) );
  XNOR U12430 ( .A(n12493), .B(n12492), .Z(n12475) );
  XNOR U12431 ( .A(n12513), .B(n12498), .Z(n12492) );
  XOR U12432 ( .A(p_input[2056]), .B(p_input[888]), .Z(n12498) );
  XOR U12433 ( .A(n12489), .B(n12497), .Z(n12513) );
  XOR U12434 ( .A(n12514), .B(n12494), .Z(n12497) );
  XOR U12435 ( .A(p_input[2054]), .B(p_input[886]), .Z(n12494) );
  XNOR U12436 ( .A(p_input[2055]), .B(p_input[887]), .Z(n12514) );
  XNOR U12437 ( .A(n6328), .B(p_input[882]), .Z(n12489) );
  XNOR U12438 ( .A(n12503), .B(n12502), .Z(n12493) );
  XOR U12439 ( .A(n12515), .B(n12499), .Z(n12502) );
  XOR U12440 ( .A(p_input[2051]), .B(p_input[883]), .Z(n12499) );
  XNOR U12441 ( .A(p_input[2052]), .B(p_input[884]), .Z(n12515) );
  XOR U12442 ( .A(p_input[2053]), .B(p_input[885]), .Z(n12503) );
  XOR U12443 ( .A(n12516), .B(n12517), .Z(n12404) );
  AND U12444 ( .A(n227), .B(n12518), .Z(n12517) );
  XNOR U12445 ( .A(n12519), .B(n12516), .Z(n12518) );
  XNOR U12446 ( .A(n12520), .B(n12521), .Z(n227) );
  AND U12447 ( .A(n12522), .B(n12523), .Z(n12521) );
  XOR U12448 ( .A(n12417), .B(n12520), .Z(n12523) );
  AND U12449 ( .A(n12524), .B(n12525), .Z(n12417) );
  XNOR U12450 ( .A(n12414), .B(n12520), .Z(n12522) );
  XOR U12451 ( .A(n12526), .B(n12527), .Z(n12414) );
  AND U12452 ( .A(n231), .B(n12528), .Z(n12527) );
  XOR U12453 ( .A(n12529), .B(n12526), .Z(n12528) );
  XOR U12454 ( .A(n12530), .B(n12531), .Z(n12520) );
  AND U12455 ( .A(n12532), .B(n12533), .Z(n12531) );
  XNOR U12456 ( .A(n12530), .B(n12524), .Z(n12533) );
  IV U12457 ( .A(n12432), .Z(n12524) );
  XOR U12458 ( .A(n12534), .B(n12535), .Z(n12432) );
  XOR U12459 ( .A(n12536), .B(n12525), .Z(n12535) );
  AND U12460 ( .A(n12459), .B(n12537), .Z(n12525) );
  AND U12461 ( .A(n12538), .B(n12539), .Z(n12536) );
  XOR U12462 ( .A(n12540), .B(n12534), .Z(n12538) );
  XNOR U12463 ( .A(n12429), .B(n12530), .Z(n12532) );
  XOR U12464 ( .A(n12541), .B(n12542), .Z(n12429) );
  AND U12465 ( .A(n231), .B(n12543), .Z(n12542) );
  XOR U12466 ( .A(n12544), .B(n12541), .Z(n12543) );
  XOR U12467 ( .A(n12545), .B(n12546), .Z(n12530) );
  AND U12468 ( .A(n12547), .B(n12548), .Z(n12546) );
  XNOR U12469 ( .A(n12545), .B(n12459), .Z(n12548) );
  XOR U12470 ( .A(n12549), .B(n12539), .Z(n12459) );
  XNOR U12471 ( .A(n12550), .B(n12534), .Z(n12539) );
  XOR U12472 ( .A(n12551), .B(n12552), .Z(n12534) );
  AND U12473 ( .A(n12553), .B(n12554), .Z(n12552) );
  XOR U12474 ( .A(n12555), .B(n12551), .Z(n12553) );
  XNOR U12475 ( .A(n12556), .B(n12557), .Z(n12550) );
  AND U12476 ( .A(n12558), .B(n12559), .Z(n12557) );
  XOR U12477 ( .A(n12556), .B(n12560), .Z(n12558) );
  XNOR U12478 ( .A(n12540), .B(n12537), .Z(n12549) );
  AND U12479 ( .A(n12561), .B(n12562), .Z(n12537) );
  XOR U12480 ( .A(n12563), .B(n12564), .Z(n12540) );
  AND U12481 ( .A(n12565), .B(n12566), .Z(n12564) );
  XOR U12482 ( .A(n12563), .B(n12567), .Z(n12565) );
  XNOR U12483 ( .A(n12456), .B(n12545), .Z(n12547) );
  XOR U12484 ( .A(n12568), .B(n12569), .Z(n12456) );
  AND U12485 ( .A(n231), .B(n12570), .Z(n12569) );
  XNOR U12486 ( .A(n12571), .B(n12568), .Z(n12570) );
  XOR U12487 ( .A(n12572), .B(n12573), .Z(n12545) );
  AND U12488 ( .A(n12574), .B(n12575), .Z(n12573) );
  XNOR U12489 ( .A(n12572), .B(n12561), .Z(n12575) );
  IV U12490 ( .A(n12507), .Z(n12561) );
  XNOR U12491 ( .A(n12576), .B(n12554), .Z(n12507) );
  XNOR U12492 ( .A(n12577), .B(n12560), .Z(n12554) );
  XOR U12493 ( .A(n12578), .B(n12579), .Z(n12560) );
  NOR U12494 ( .A(n12580), .B(n12581), .Z(n12579) );
  XNOR U12495 ( .A(n12578), .B(n12582), .Z(n12580) );
  XNOR U12496 ( .A(n12559), .B(n12551), .Z(n12577) );
  XOR U12497 ( .A(n12583), .B(n12584), .Z(n12551) );
  AND U12498 ( .A(n12585), .B(n12586), .Z(n12584) );
  XNOR U12499 ( .A(n12583), .B(n12587), .Z(n12585) );
  XNOR U12500 ( .A(n12588), .B(n12556), .Z(n12559) );
  XOR U12501 ( .A(n12589), .B(n12590), .Z(n12556) );
  AND U12502 ( .A(n12591), .B(n12592), .Z(n12590) );
  XOR U12503 ( .A(n12589), .B(n12593), .Z(n12591) );
  XNOR U12504 ( .A(n12594), .B(n12595), .Z(n12588) );
  NOR U12505 ( .A(n12596), .B(n12597), .Z(n12595) );
  XOR U12506 ( .A(n12594), .B(n12598), .Z(n12596) );
  XNOR U12507 ( .A(n12555), .B(n12562), .Z(n12576) );
  NOR U12508 ( .A(n12519), .B(n12599), .Z(n12562) );
  XOR U12509 ( .A(n12567), .B(n12566), .Z(n12555) );
  XNOR U12510 ( .A(n12600), .B(n12563), .Z(n12566) );
  XOR U12511 ( .A(n12601), .B(n12602), .Z(n12563) );
  AND U12512 ( .A(n12603), .B(n12604), .Z(n12602) );
  XOR U12513 ( .A(n12601), .B(n12605), .Z(n12603) );
  XNOR U12514 ( .A(n12606), .B(n12607), .Z(n12600) );
  NOR U12515 ( .A(n12608), .B(n12609), .Z(n12607) );
  XNOR U12516 ( .A(n12606), .B(n12610), .Z(n12608) );
  XOR U12517 ( .A(n12611), .B(n12612), .Z(n12567) );
  NOR U12518 ( .A(n12613), .B(n12614), .Z(n12612) );
  XNOR U12519 ( .A(n12611), .B(n12615), .Z(n12613) );
  XNOR U12520 ( .A(n12504), .B(n12572), .Z(n12574) );
  XOR U12521 ( .A(n12616), .B(n12617), .Z(n12504) );
  AND U12522 ( .A(n231), .B(n12618), .Z(n12617) );
  XOR U12523 ( .A(n12619), .B(n12616), .Z(n12618) );
  AND U12524 ( .A(n12516), .B(n12519), .Z(n12572) );
  XOR U12525 ( .A(n12620), .B(n12599), .Z(n12519) );
  XNOR U12526 ( .A(p_input[2048]), .B(p_input[896]), .Z(n12599) );
  XOR U12527 ( .A(n12587), .B(n12586), .Z(n12620) );
  XNOR U12528 ( .A(n12621), .B(n12593), .Z(n12586) );
  XNOR U12529 ( .A(n12582), .B(n12581), .Z(n12593) );
  XOR U12530 ( .A(n12622), .B(n12578), .Z(n12581) );
  XNOR U12531 ( .A(n6439), .B(p_input[906]), .Z(n12578) );
  XNOR U12532 ( .A(p_input[2059]), .B(p_input[907]), .Z(n12622) );
  XOR U12533 ( .A(p_input[2060]), .B(p_input[908]), .Z(n12582) );
  XNOR U12534 ( .A(n12592), .B(n12583), .Z(n12621) );
  XNOR U12535 ( .A(n6553), .B(p_input[897]), .Z(n12583) );
  XOR U12536 ( .A(n12623), .B(n12598), .Z(n12592) );
  XNOR U12537 ( .A(p_input[2063]), .B(p_input[911]), .Z(n12598) );
  XOR U12538 ( .A(n12589), .B(n12597), .Z(n12623) );
  XOR U12539 ( .A(n12624), .B(n12594), .Z(n12597) );
  XOR U12540 ( .A(p_input[2061]), .B(p_input[909]), .Z(n12594) );
  XNOR U12541 ( .A(p_input[2062]), .B(p_input[910]), .Z(n12624) );
  XNOR U12542 ( .A(n6325), .B(p_input[905]), .Z(n12589) );
  XNOR U12543 ( .A(n12605), .B(n12604), .Z(n12587) );
  XNOR U12544 ( .A(n12625), .B(n12610), .Z(n12604) );
  XOR U12545 ( .A(p_input[2056]), .B(p_input[904]), .Z(n12610) );
  XOR U12546 ( .A(n12601), .B(n12609), .Z(n12625) );
  XOR U12547 ( .A(n12626), .B(n12606), .Z(n12609) );
  XOR U12548 ( .A(p_input[2054]), .B(p_input[902]), .Z(n12606) );
  XNOR U12549 ( .A(p_input[2055]), .B(p_input[903]), .Z(n12626) );
  XNOR U12550 ( .A(n6328), .B(p_input[898]), .Z(n12601) );
  XNOR U12551 ( .A(n12615), .B(n12614), .Z(n12605) );
  XOR U12552 ( .A(n12627), .B(n12611), .Z(n12614) );
  XOR U12553 ( .A(p_input[2051]), .B(p_input[899]), .Z(n12611) );
  XNOR U12554 ( .A(p_input[2052]), .B(p_input[900]), .Z(n12627) );
  XOR U12555 ( .A(p_input[2053]), .B(p_input[901]), .Z(n12615) );
  XOR U12556 ( .A(n12628), .B(n12629), .Z(n12516) );
  AND U12557 ( .A(n231), .B(n12630), .Z(n12629) );
  XNOR U12558 ( .A(n12631), .B(n12628), .Z(n12630) );
  XNOR U12559 ( .A(n12632), .B(n12633), .Z(n231) );
  AND U12560 ( .A(n12634), .B(n12635), .Z(n12633) );
  XOR U12561 ( .A(n12529), .B(n12632), .Z(n12635) );
  AND U12562 ( .A(n12636), .B(n12637), .Z(n12529) );
  XNOR U12563 ( .A(n12526), .B(n12632), .Z(n12634) );
  XOR U12564 ( .A(n12638), .B(n12639), .Z(n12526) );
  AND U12565 ( .A(n235), .B(n12640), .Z(n12639) );
  XOR U12566 ( .A(n12641), .B(n12638), .Z(n12640) );
  XOR U12567 ( .A(n12642), .B(n12643), .Z(n12632) );
  AND U12568 ( .A(n12644), .B(n12645), .Z(n12643) );
  XNOR U12569 ( .A(n12642), .B(n12636), .Z(n12645) );
  IV U12570 ( .A(n12544), .Z(n12636) );
  XOR U12571 ( .A(n12646), .B(n12647), .Z(n12544) );
  XOR U12572 ( .A(n12648), .B(n12637), .Z(n12647) );
  AND U12573 ( .A(n12571), .B(n12649), .Z(n12637) );
  AND U12574 ( .A(n12650), .B(n12651), .Z(n12648) );
  XOR U12575 ( .A(n12652), .B(n12646), .Z(n12650) );
  XNOR U12576 ( .A(n12541), .B(n12642), .Z(n12644) );
  XOR U12577 ( .A(n12653), .B(n12654), .Z(n12541) );
  AND U12578 ( .A(n235), .B(n12655), .Z(n12654) );
  XOR U12579 ( .A(n12656), .B(n12653), .Z(n12655) );
  XOR U12580 ( .A(n12657), .B(n12658), .Z(n12642) );
  AND U12581 ( .A(n12659), .B(n12660), .Z(n12658) );
  XNOR U12582 ( .A(n12657), .B(n12571), .Z(n12660) );
  XOR U12583 ( .A(n12661), .B(n12651), .Z(n12571) );
  XNOR U12584 ( .A(n12662), .B(n12646), .Z(n12651) );
  XOR U12585 ( .A(n12663), .B(n12664), .Z(n12646) );
  AND U12586 ( .A(n12665), .B(n12666), .Z(n12664) );
  XOR U12587 ( .A(n12667), .B(n12663), .Z(n12665) );
  XNOR U12588 ( .A(n12668), .B(n12669), .Z(n12662) );
  AND U12589 ( .A(n12670), .B(n12671), .Z(n12669) );
  XOR U12590 ( .A(n12668), .B(n12672), .Z(n12670) );
  XNOR U12591 ( .A(n12652), .B(n12649), .Z(n12661) );
  AND U12592 ( .A(n12673), .B(n12674), .Z(n12649) );
  XOR U12593 ( .A(n12675), .B(n12676), .Z(n12652) );
  AND U12594 ( .A(n12677), .B(n12678), .Z(n12676) );
  XOR U12595 ( .A(n12675), .B(n12679), .Z(n12677) );
  XNOR U12596 ( .A(n12568), .B(n12657), .Z(n12659) );
  XOR U12597 ( .A(n12680), .B(n12681), .Z(n12568) );
  AND U12598 ( .A(n235), .B(n12682), .Z(n12681) );
  XNOR U12599 ( .A(n12683), .B(n12680), .Z(n12682) );
  XOR U12600 ( .A(n12684), .B(n12685), .Z(n12657) );
  AND U12601 ( .A(n12686), .B(n12687), .Z(n12685) );
  XNOR U12602 ( .A(n12684), .B(n12673), .Z(n12687) );
  IV U12603 ( .A(n12619), .Z(n12673) );
  XNOR U12604 ( .A(n12688), .B(n12666), .Z(n12619) );
  XNOR U12605 ( .A(n12689), .B(n12672), .Z(n12666) );
  XOR U12606 ( .A(n12690), .B(n12691), .Z(n12672) );
  NOR U12607 ( .A(n12692), .B(n12693), .Z(n12691) );
  XNOR U12608 ( .A(n12690), .B(n12694), .Z(n12692) );
  XNOR U12609 ( .A(n12671), .B(n12663), .Z(n12689) );
  XOR U12610 ( .A(n12695), .B(n12696), .Z(n12663) );
  AND U12611 ( .A(n12697), .B(n12698), .Z(n12696) );
  XNOR U12612 ( .A(n12695), .B(n12699), .Z(n12697) );
  XNOR U12613 ( .A(n12700), .B(n12668), .Z(n12671) );
  XOR U12614 ( .A(n12701), .B(n12702), .Z(n12668) );
  AND U12615 ( .A(n12703), .B(n12704), .Z(n12702) );
  XOR U12616 ( .A(n12701), .B(n12705), .Z(n12703) );
  XNOR U12617 ( .A(n12706), .B(n12707), .Z(n12700) );
  NOR U12618 ( .A(n12708), .B(n12709), .Z(n12707) );
  XOR U12619 ( .A(n12706), .B(n12710), .Z(n12708) );
  XNOR U12620 ( .A(n12667), .B(n12674), .Z(n12688) );
  NOR U12621 ( .A(n12631), .B(n12711), .Z(n12674) );
  XOR U12622 ( .A(n12679), .B(n12678), .Z(n12667) );
  XNOR U12623 ( .A(n12712), .B(n12675), .Z(n12678) );
  XOR U12624 ( .A(n12713), .B(n12714), .Z(n12675) );
  AND U12625 ( .A(n12715), .B(n12716), .Z(n12714) );
  XOR U12626 ( .A(n12713), .B(n12717), .Z(n12715) );
  XNOR U12627 ( .A(n12718), .B(n12719), .Z(n12712) );
  NOR U12628 ( .A(n12720), .B(n12721), .Z(n12719) );
  XNOR U12629 ( .A(n12718), .B(n12722), .Z(n12720) );
  XOR U12630 ( .A(n12723), .B(n12724), .Z(n12679) );
  NOR U12631 ( .A(n12725), .B(n12726), .Z(n12724) );
  XNOR U12632 ( .A(n12723), .B(n12727), .Z(n12725) );
  XNOR U12633 ( .A(n12616), .B(n12684), .Z(n12686) );
  XOR U12634 ( .A(n12728), .B(n12729), .Z(n12616) );
  AND U12635 ( .A(n235), .B(n12730), .Z(n12729) );
  XOR U12636 ( .A(n12731), .B(n12728), .Z(n12730) );
  AND U12637 ( .A(n12628), .B(n12631), .Z(n12684) );
  XOR U12638 ( .A(n12732), .B(n12711), .Z(n12631) );
  XNOR U12639 ( .A(p_input[2048]), .B(p_input[912]), .Z(n12711) );
  XOR U12640 ( .A(n12699), .B(n12698), .Z(n12732) );
  XNOR U12641 ( .A(n12733), .B(n12705), .Z(n12698) );
  XNOR U12642 ( .A(n12694), .B(n12693), .Z(n12705) );
  XOR U12643 ( .A(n12734), .B(n12690), .Z(n12693) );
  XNOR U12644 ( .A(n6439), .B(p_input[922]), .Z(n12690) );
  XNOR U12645 ( .A(p_input[2059]), .B(p_input[923]), .Z(n12734) );
  XOR U12646 ( .A(p_input[2060]), .B(p_input[924]), .Z(n12694) );
  XNOR U12647 ( .A(n12704), .B(n12695), .Z(n12733) );
  XNOR U12648 ( .A(n6553), .B(p_input[913]), .Z(n12695) );
  XOR U12649 ( .A(n12735), .B(n12710), .Z(n12704) );
  XNOR U12650 ( .A(p_input[2063]), .B(p_input[927]), .Z(n12710) );
  XOR U12651 ( .A(n12701), .B(n12709), .Z(n12735) );
  XOR U12652 ( .A(n12736), .B(n12706), .Z(n12709) );
  XOR U12653 ( .A(p_input[2061]), .B(p_input[925]), .Z(n12706) );
  XNOR U12654 ( .A(p_input[2062]), .B(p_input[926]), .Z(n12736) );
  XNOR U12655 ( .A(n6325), .B(p_input[921]), .Z(n12701) );
  XNOR U12656 ( .A(n12717), .B(n12716), .Z(n12699) );
  XNOR U12657 ( .A(n12737), .B(n12722), .Z(n12716) );
  XOR U12658 ( .A(p_input[2056]), .B(p_input[920]), .Z(n12722) );
  XOR U12659 ( .A(n12713), .B(n12721), .Z(n12737) );
  XOR U12660 ( .A(n12738), .B(n12718), .Z(n12721) );
  XOR U12661 ( .A(p_input[2054]), .B(p_input[918]), .Z(n12718) );
  XNOR U12662 ( .A(p_input[2055]), .B(p_input[919]), .Z(n12738) );
  XNOR U12663 ( .A(n6328), .B(p_input[914]), .Z(n12713) );
  XNOR U12664 ( .A(n12727), .B(n12726), .Z(n12717) );
  XOR U12665 ( .A(n12739), .B(n12723), .Z(n12726) );
  XOR U12666 ( .A(p_input[2051]), .B(p_input[915]), .Z(n12723) );
  XNOR U12667 ( .A(p_input[2052]), .B(p_input[916]), .Z(n12739) );
  XOR U12668 ( .A(p_input[2053]), .B(p_input[917]), .Z(n12727) );
  XOR U12669 ( .A(n12740), .B(n12741), .Z(n12628) );
  AND U12670 ( .A(n235), .B(n12742), .Z(n12741) );
  XNOR U12671 ( .A(n12743), .B(n12740), .Z(n12742) );
  XNOR U12672 ( .A(n12744), .B(n12745), .Z(n235) );
  AND U12673 ( .A(n12746), .B(n12747), .Z(n12745) );
  XOR U12674 ( .A(n12641), .B(n12744), .Z(n12747) );
  AND U12675 ( .A(n12748), .B(n12749), .Z(n12641) );
  XNOR U12676 ( .A(n12638), .B(n12744), .Z(n12746) );
  XOR U12677 ( .A(n12750), .B(n12751), .Z(n12638) );
  AND U12678 ( .A(n239), .B(n12752), .Z(n12751) );
  XOR U12679 ( .A(n12753), .B(n12750), .Z(n12752) );
  XOR U12680 ( .A(n12754), .B(n12755), .Z(n12744) );
  AND U12681 ( .A(n12756), .B(n12757), .Z(n12755) );
  XNOR U12682 ( .A(n12754), .B(n12748), .Z(n12757) );
  IV U12683 ( .A(n12656), .Z(n12748) );
  XOR U12684 ( .A(n12758), .B(n12759), .Z(n12656) );
  XOR U12685 ( .A(n12760), .B(n12749), .Z(n12759) );
  AND U12686 ( .A(n12683), .B(n12761), .Z(n12749) );
  AND U12687 ( .A(n12762), .B(n12763), .Z(n12760) );
  XOR U12688 ( .A(n12764), .B(n12758), .Z(n12762) );
  XNOR U12689 ( .A(n12653), .B(n12754), .Z(n12756) );
  XOR U12690 ( .A(n12765), .B(n12766), .Z(n12653) );
  AND U12691 ( .A(n239), .B(n12767), .Z(n12766) );
  XOR U12692 ( .A(n12768), .B(n12765), .Z(n12767) );
  XOR U12693 ( .A(n12769), .B(n12770), .Z(n12754) );
  AND U12694 ( .A(n12771), .B(n12772), .Z(n12770) );
  XNOR U12695 ( .A(n12769), .B(n12683), .Z(n12772) );
  XOR U12696 ( .A(n12773), .B(n12763), .Z(n12683) );
  XNOR U12697 ( .A(n12774), .B(n12758), .Z(n12763) );
  XOR U12698 ( .A(n12775), .B(n12776), .Z(n12758) );
  AND U12699 ( .A(n12777), .B(n12778), .Z(n12776) );
  XOR U12700 ( .A(n12779), .B(n12775), .Z(n12777) );
  XNOR U12701 ( .A(n12780), .B(n12781), .Z(n12774) );
  AND U12702 ( .A(n12782), .B(n12783), .Z(n12781) );
  XOR U12703 ( .A(n12780), .B(n12784), .Z(n12782) );
  XNOR U12704 ( .A(n12764), .B(n12761), .Z(n12773) );
  AND U12705 ( .A(n12785), .B(n12786), .Z(n12761) );
  XOR U12706 ( .A(n12787), .B(n12788), .Z(n12764) );
  AND U12707 ( .A(n12789), .B(n12790), .Z(n12788) );
  XOR U12708 ( .A(n12787), .B(n12791), .Z(n12789) );
  XNOR U12709 ( .A(n12680), .B(n12769), .Z(n12771) );
  XOR U12710 ( .A(n12792), .B(n12793), .Z(n12680) );
  AND U12711 ( .A(n239), .B(n12794), .Z(n12793) );
  XNOR U12712 ( .A(n12795), .B(n12792), .Z(n12794) );
  XOR U12713 ( .A(n12796), .B(n12797), .Z(n12769) );
  AND U12714 ( .A(n12798), .B(n12799), .Z(n12797) );
  XNOR U12715 ( .A(n12796), .B(n12785), .Z(n12799) );
  IV U12716 ( .A(n12731), .Z(n12785) );
  XNOR U12717 ( .A(n12800), .B(n12778), .Z(n12731) );
  XNOR U12718 ( .A(n12801), .B(n12784), .Z(n12778) );
  XOR U12719 ( .A(n12802), .B(n12803), .Z(n12784) );
  NOR U12720 ( .A(n12804), .B(n12805), .Z(n12803) );
  XNOR U12721 ( .A(n12802), .B(n12806), .Z(n12804) );
  XNOR U12722 ( .A(n12783), .B(n12775), .Z(n12801) );
  XOR U12723 ( .A(n12807), .B(n12808), .Z(n12775) );
  AND U12724 ( .A(n12809), .B(n12810), .Z(n12808) );
  XNOR U12725 ( .A(n12807), .B(n12811), .Z(n12809) );
  XNOR U12726 ( .A(n12812), .B(n12780), .Z(n12783) );
  XOR U12727 ( .A(n12813), .B(n12814), .Z(n12780) );
  AND U12728 ( .A(n12815), .B(n12816), .Z(n12814) );
  XOR U12729 ( .A(n12813), .B(n12817), .Z(n12815) );
  XNOR U12730 ( .A(n12818), .B(n12819), .Z(n12812) );
  NOR U12731 ( .A(n12820), .B(n12821), .Z(n12819) );
  XOR U12732 ( .A(n12818), .B(n12822), .Z(n12820) );
  XNOR U12733 ( .A(n12779), .B(n12786), .Z(n12800) );
  NOR U12734 ( .A(n12743), .B(n12823), .Z(n12786) );
  XOR U12735 ( .A(n12791), .B(n12790), .Z(n12779) );
  XNOR U12736 ( .A(n12824), .B(n12787), .Z(n12790) );
  XOR U12737 ( .A(n12825), .B(n12826), .Z(n12787) );
  AND U12738 ( .A(n12827), .B(n12828), .Z(n12826) );
  XOR U12739 ( .A(n12825), .B(n12829), .Z(n12827) );
  XNOR U12740 ( .A(n12830), .B(n12831), .Z(n12824) );
  NOR U12741 ( .A(n12832), .B(n12833), .Z(n12831) );
  XNOR U12742 ( .A(n12830), .B(n12834), .Z(n12832) );
  XOR U12743 ( .A(n12835), .B(n12836), .Z(n12791) );
  NOR U12744 ( .A(n12837), .B(n12838), .Z(n12836) );
  XNOR U12745 ( .A(n12835), .B(n12839), .Z(n12837) );
  XNOR U12746 ( .A(n12728), .B(n12796), .Z(n12798) );
  XOR U12747 ( .A(n12840), .B(n12841), .Z(n12728) );
  AND U12748 ( .A(n239), .B(n12842), .Z(n12841) );
  XOR U12749 ( .A(n12843), .B(n12840), .Z(n12842) );
  AND U12750 ( .A(n12740), .B(n12743), .Z(n12796) );
  XOR U12751 ( .A(n12844), .B(n12823), .Z(n12743) );
  XNOR U12752 ( .A(p_input[2048]), .B(p_input[928]), .Z(n12823) );
  XOR U12753 ( .A(n12811), .B(n12810), .Z(n12844) );
  XNOR U12754 ( .A(n12845), .B(n12817), .Z(n12810) );
  XNOR U12755 ( .A(n12806), .B(n12805), .Z(n12817) );
  XOR U12756 ( .A(n12846), .B(n12802), .Z(n12805) );
  XNOR U12757 ( .A(n6439), .B(p_input[938]), .Z(n12802) );
  XNOR U12758 ( .A(p_input[2059]), .B(p_input[939]), .Z(n12846) );
  XOR U12759 ( .A(p_input[2060]), .B(p_input[940]), .Z(n12806) );
  XNOR U12760 ( .A(n12816), .B(n12807), .Z(n12845) );
  XNOR U12761 ( .A(n6553), .B(p_input[929]), .Z(n12807) );
  XOR U12762 ( .A(n12847), .B(n12822), .Z(n12816) );
  XNOR U12763 ( .A(p_input[2063]), .B(p_input[943]), .Z(n12822) );
  XOR U12764 ( .A(n12813), .B(n12821), .Z(n12847) );
  XOR U12765 ( .A(n12848), .B(n12818), .Z(n12821) );
  XOR U12766 ( .A(p_input[2061]), .B(p_input[941]), .Z(n12818) );
  XNOR U12767 ( .A(p_input[2062]), .B(p_input[942]), .Z(n12848) );
  XNOR U12768 ( .A(n6325), .B(p_input[937]), .Z(n12813) );
  XNOR U12769 ( .A(n12829), .B(n12828), .Z(n12811) );
  XNOR U12770 ( .A(n12849), .B(n12834), .Z(n12828) );
  XOR U12771 ( .A(p_input[2056]), .B(p_input[936]), .Z(n12834) );
  XOR U12772 ( .A(n12825), .B(n12833), .Z(n12849) );
  XOR U12773 ( .A(n12850), .B(n12830), .Z(n12833) );
  XOR U12774 ( .A(p_input[2054]), .B(p_input[934]), .Z(n12830) );
  XNOR U12775 ( .A(p_input[2055]), .B(p_input[935]), .Z(n12850) );
  XNOR U12776 ( .A(n6328), .B(p_input[930]), .Z(n12825) );
  XNOR U12777 ( .A(n12839), .B(n12838), .Z(n12829) );
  XOR U12778 ( .A(n12851), .B(n12835), .Z(n12838) );
  XOR U12779 ( .A(p_input[2051]), .B(p_input[931]), .Z(n12835) );
  XNOR U12780 ( .A(p_input[2052]), .B(p_input[932]), .Z(n12851) );
  XOR U12781 ( .A(p_input[2053]), .B(p_input[933]), .Z(n12839) );
  XOR U12782 ( .A(n12852), .B(n12853), .Z(n12740) );
  AND U12783 ( .A(n239), .B(n12854), .Z(n12853) );
  XNOR U12784 ( .A(n12855), .B(n12852), .Z(n12854) );
  XNOR U12785 ( .A(n12856), .B(n12857), .Z(n239) );
  AND U12786 ( .A(n12858), .B(n12859), .Z(n12857) );
  XOR U12787 ( .A(n12753), .B(n12856), .Z(n12859) );
  AND U12788 ( .A(n12860), .B(n12861), .Z(n12753) );
  XNOR U12789 ( .A(n12750), .B(n12856), .Z(n12858) );
  XOR U12790 ( .A(n12862), .B(n12863), .Z(n12750) );
  AND U12791 ( .A(n243), .B(n12864), .Z(n12863) );
  XOR U12792 ( .A(n12865), .B(n12862), .Z(n12864) );
  XOR U12793 ( .A(n12866), .B(n12867), .Z(n12856) );
  AND U12794 ( .A(n12868), .B(n12869), .Z(n12867) );
  XNOR U12795 ( .A(n12866), .B(n12860), .Z(n12869) );
  IV U12796 ( .A(n12768), .Z(n12860) );
  XOR U12797 ( .A(n12870), .B(n12871), .Z(n12768) );
  XOR U12798 ( .A(n12872), .B(n12861), .Z(n12871) );
  AND U12799 ( .A(n12795), .B(n12873), .Z(n12861) );
  AND U12800 ( .A(n12874), .B(n12875), .Z(n12872) );
  XOR U12801 ( .A(n12876), .B(n12870), .Z(n12874) );
  XNOR U12802 ( .A(n12765), .B(n12866), .Z(n12868) );
  XOR U12803 ( .A(n12877), .B(n12878), .Z(n12765) );
  AND U12804 ( .A(n243), .B(n12879), .Z(n12878) );
  XOR U12805 ( .A(n12880), .B(n12877), .Z(n12879) );
  XOR U12806 ( .A(n12881), .B(n12882), .Z(n12866) );
  AND U12807 ( .A(n12883), .B(n12884), .Z(n12882) );
  XNOR U12808 ( .A(n12881), .B(n12795), .Z(n12884) );
  XOR U12809 ( .A(n12885), .B(n12875), .Z(n12795) );
  XNOR U12810 ( .A(n12886), .B(n12870), .Z(n12875) );
  XOR U12811 ( .A(n12887), .B(n12888), .Z(n12870) );
  AND U12812 ( .A(n12889), .B(n12890), .Z(n12888) );
  XOR U12813 ( .A(n12891), .B(n12887), .Z(n12889) );
  XNOR U12814 ( .A(n12892), .B(n12893), .Z(n12886) );
  AND U12815 ( .A(n12894), .B(n12895), .Z(n12893) );
  XOR U12816 ( .A(n12892), .B(n12896), .Z(n12894) );
  XNOR U12817 ( .A(n12876), .B(n12873), .Z(n12885) );
  AND U12818 ( .A(n12897), .B(n12898), .Z(n12873) );
  XOR U12819 ( .A(n12899), .B(n12900), .Z(n12876) );
  AND U12820 ( .A(n12901), .B(n12902), .Z(n12900) );
  XOR U12821 ( .A(n12899), .B(n12903), .Z(n12901) );
  XNOR U12822 ( .A(n12792), .B(n12881), .Z(n12883) );
  XOR U12823 ( .A(n12904), .B(n12905), .Z(n12792) );
  AND U12824 ( .A(n243), .B(n12906), .Z(n12905) );
  XNOR U12825 ( .A(n12907), .B(n12904), .Z(n12906) );
  XOR U12826 ( .A(n12908), .B(n12909), .Z(n12881) );
  AND U12827 ( .A(n12910), .B(n12911), .Z(n12909) );
  XNOR U12828 ( .A(n12908), .B(n12897), .Z(n12911) );
  IV U12829 ( .A(n12843), .Z(n12897) );
  XNOR U12830 ( .A(n12912), .B(n12890), .Z(n12843) );
  XNOR U12831 ( .A(n12913), .B(n12896), .Z(n12890) );
  XOR U12832 ( .A(n12914), .B(n12915), .Z(n12896) );
  NOR U12833 ( .A(n12916), .B(n12917), .Z(n12915) );
  XNOR U12834 ( .A(n12914), .B(n12918), .Z(n12916) );
  XNOR U12835 ( .A(n12895), .B(n12887), .Z(n12913) );
  XOR U12836 ( .A(n12919), .B(n12920), .Z(n12887) );
  AND U12837 ( .A(n12921), .B(n12922), .Z(n12920) );
  XNOR U12838 ( .A(n12919), .B(n12923), .Z(n12921) );
  XNOR U12839 ( .A(n12924), .B(n12892), .Z(n12895) );
  XOR U12840 ( .A(n12925), .B(n12926), .Z(n12892) );
  AND U12841 ( .A(n12927), .B(n12928), .Z(n12926) );
  XOR U12842 ( .A(n12925), .B(n12929), .Z(n12927) );
  XNOR U12843 ( .A(n12930), .B(n12931), .Z(n12924) );
  NOR U12844 ( .A(n12932), .B(n12933), .Z(n12931) );
  XOR U12845 ( .A(n12930), .B(n12934), .Z(n12932) );
  XNOR U12846 ( .A(n12891), .B(n12898), .Z(n12912) );
  NOR U12847 ( .A(n12855), .B(n12935), .Z(n12898) );
  XOR U12848 ( .A(n12903), .B(n12902), .Z(n12891) );
  XNOR U12849 ( .A(n12936), .B(n12899), .Z(n12902) );
  XOR U12850 ( .A(n12937), .B(n12938), .Z(n12899) );
  AND U12851 ( .A(n12939), .B(n12940), .Z(n12938) );
  XOR U12852 ( .A(n12937), .B(n12941), .Z(n12939) );
  XNOR U12853 ( .A(n12942), .B(n12943), .Z(n12936) );
  NOR U12854 ( .A(n12944), .B(n12945), .Z(n12943) );
  XNOR U12855 ( .A(n12942), .B(n12946), .Z(n12944) );
  XOR U12856 ( .A(n12947), .B(n12948), .Z(n12903) );
  NOR U12857 ( .A(n12949), .B(n12950), .Z(n12948) );
  XNOR U12858 ( .A(n12947), .B(n12951), .Z(n12949) );
  XNOR U12859 ( .A(n12840), .B(n12908), .Z(n12910) );
  XOR U12860 ( .A(n12952), .B(n12953), .Z(n12840) );
  AND U12861 ( .A(n243), .B(n12954), .Z(n12953) );
  XOR U12862 ( .A(n12955), .B(n12952), .Z(n12954) );
  AND U12863 ( .A(n12852), .B(n12855), .Z(n12908) );
  XOR U12864 ( .A(n12956), .B(n12935), .Z(n12855) );
  XNOR U12865 ( .A(p_input[2048]), .B(p_input[944]), .Z(n12935) );
  XOR U12866 ( .A(n12923), .B(n12922), .Z(n12956) );
  XNOR U12867 ( .A(n12957), .B(n12929), .Z(n12922) );
  XNOR U12868 ( .A(n12918), .B(n12917), .Z(n12929) );
  XOR U12869 ( .A(n12958), .B(n12914), .Z(n12917) );
  XNOR U12870 ( .A(n6439), .B(p_input[954]), .Z(n12914) );
  XNOR U12871 ( .A(p_input[2059]), .B(p_input[955]), .Z(n12958) );
  XOR U12872 ( .A(p_input[2060]), .B(p_input[956]), .Z(n12918) );
  XNOR U12873 ( .A(n12928), .B(n12919), .Z(n12957) );
  XNOR U12874 ( .A(n6553), .B(p_input[945]), .Z(n12919) );
  XOR U12875 ( .A(n12959), .B(n12934), .Z(n12928) );
  XNOR U12876 ( .A(p_input[2063]), .B(p_input[959]), .Z(n12934) );
  XOR U12877 ( .A(n12925), .B(n12933), .Z(n12959) );
  XOR U12878 ( .A(n12960), .B(n12930), .Z(n12933) );
  XOR U12879 ( .A(p_input[2061]), .B(p_input[957]), .Z(n12930) );
  XNOR U12880 ( .A(p_input[2062]), .B(p_input[958]), .Z(n12960) );
  XNOR U12881 ( .A(n6325), .B(p_input[953]), .Z(n12925) );
  XNOR U12882 ( .A(n12941), .B(n12940), .Z(n12923) );
  XNOR U12883 ( .A(n12961), .B(n12946), .Z(n12940) );
  XOR U12884 ( .A(p_input[2056]), .B(p_input[952]), .Z(n12946) );
  XOR U12885 ( .A(n12937), .B(n12945), .Z(n12961) );
  XOR U12886 ( .A(n12962), .B(n12942), .Z(n12945) );
  XOR U12887 ( .A(p_input[2054]), .B(p_input[950]), .Z(n12942) );
  XNOR U12888 ( .A(p_input[2055]), .B(p_input[951]), .Z(n12962) );
  XNOR U12889 ( .A(n6328), .B(p_input[946]), .Z(n12937) );
  XNOR U12890 ( .A(n12951), .B(n12950), .Z(n12941) );
  XOR U12891 ( .A(n12963), .B(n12947), .Z(n12950) );
  XOR U12892 ( .A(p_input[2051]), .B(p_input[947]), .Z(n12947) );
  XNOR U12893 ( .A(p_input[2052]), .B(p_input[948]), .Z(n12963) );
  XOR U12894 ( .A(p_input[2053]), .B(p_input[949]), .Z(n12951) );
  XOR U12895 ( .A(n12964), .B(n12965), .Z(n12852) );
  AND U12896 ( .A(n243), .B(n12966), .Z(n12965) );
  XNOR U12897 ( .A(n12967), .B(n12964), .Z(n12966) );
  XNOR U12898 ( .A(n12968), .B(n12969), .Z(n243) );
  AND U12899 ( .A(n12970), .B(n12971), .Z(n12969) );
  XOR U12900 ( .A(n12865), .B(n12968), .Z(n12971) );
  AND U12901 ( .A(n12972), .B(n12973), .Z(n12865) );
  XNOR U12902 ( .A(n12862), .B(n12968), .Z(n12970) );
  XOR U12903 ( .A(n12974), .B(n12975), .Z(n12862) );
  AND U12904 ( .A(n247), .B(n12976), .Z(n12975) );
  XOR U12905 ( .A(n12977), .B(n12974), .Z(n12976) );
  XOR U12906 ( .A(n12978), .B(n12979), .Z(n12968) );
  AND U12907 ( .A(n12980), .B(n12981), .Z(n12979) );
  XNOR U12908 ( .A(n12978), .B(n12972), .Z(n12981) );
  IV U12909 ( .A(n12880), .Z(n12972) );
  XOR U12910 ( .A(n12982), .B(n12983), .Z(n12880) );
  XOR U12911 ( .A(n12984), .B(n12973), .Z(n12983) );
  AND U12912 ( .A(n12907), .B(n12985), .Z(n12973) );
  AND U12913 ( .A(n12986), .B(n12987), .Z(n12984) );
  XOR U12914 ( .A(n12988), .B(n12982), .Z(n12986) );
  XNOR U12915 ( .A(n12877), .B(n12978), .Z(n12980) );
  XOR U12916 ( .A(n12989), .B(n12990), .Z(n12877) );
  AND U12917 ( .A(n247), .B(n12991), .Z(n12990) );
  XOR U12918 ( .A(n12992), .B(n12989), .Z(n12991) );
  XOR U12919 ( .A(n12993), .B(n12994), .Z(n12978) );
  AND U12920 ( .A(n12995), .B(n12996), .Z(n12994) );
  XNOR U12921 ( .A(n12993), .B(n12907), .Z(n12996) );
  XOR U12922 ( .A(n12997), .B(n12987), .Z(n12907) );
  XNOR U12923 ( .A(n12998), .B(n12982), .Z(n12987) );
  XOR U12924 ( .A(n12999), .B(n13000), .Z(n12982) );
  AND U12925 ( .A(n13001), .B(n13002), .Z(n13000) );
  XOR U12926 ( .A(n13003), .B(n12999), .Z(n13001) );
  XNOR U12927 ( .A(n13004), .B(n13005), .Z(n12998) );
  AND U12928 ( .A(n13006), .B(n13007), .Z(n13005) );
  XOR U12929 ( .A(n13004), .B(n13008), .Z(n13006) );
  XNOR U12930 ( .A(n12988), .B(n12985), .Z(n12997) );
  AND U12931 ( .A(n13009), .B(n13010), .Z(n12985) );
  XOR U12932 ( .A(n13011), .B(n13012), .Z(n12988) );
  AND U12933 ( .A(n13013), .B(n13014), .Z(n13012) );
  XOR U12934 ( .A(n13011), .B(n13015), .Z(n13013) );
  XNOR U12935 ( .A(n12904), .B(n12993), .Z(n12995) );
  XOR U12936 ( .A(n13016), .B(n13017), .Z(n12904) );
  AND U12937 ( .A(n247), .B(n13018), .Z(n13017) );
  XNOR U12938 ( .A(n13019), .B(n13016), .Z(n13018) );
  XOR U12939 ( .A(n13020), .B(n13021), .Z(n12993) );
  AND U12940 ( .A(n13022), .B(n13023), .Z(n13021) );
  XNOR U12941 ( .A(n13020), .B(n13009), .Z(n13023) );
  IV U12942 ( .A(n12955), .Z(n13009) );
  XNOR U12943 ( .A(n13024), .B(n13002), .Z(n12955) );
  XNOR U12944 ( .A(n13025), .B(n13008), .Z(n13002) );
  XOR U12945 ( .A(n13026), .B(n13027), .Z(n13008) );
  NOR U12946 ( .A(n13028), .B(n13029), .Z(n13027) );
  XNOR U12947 ( .A(n13026), .B(n13030), .Z(n13028) );
  XNOR U12948 ( .A(n13007), .B(n12999), .Z(n13025) );
  XOR U12949 ( .A(n13031), .B(n13032), .Z(n12999) );
  AND U12950 ( .A(n13033), .B(n13034), .Z(n13032) );
  XNOR U12951 ( .A(n13031), .B(n13035), .Z(n13033) );
  XNOR U12952 ( .A(n13036), .B(n13004), .Z(n13007) );
  XOR U12953 ( .A(n13037), .B(n13038), .Z(n13004) );
  AND U12954 ( .A(n13039), .B(n13040), .Z(n13038) );
  XOR U12955 ( .A(n13037), .B(n13041), .Z(n13039) );
  XNOR U12956 ( .A(n13042), .B(n13043), .Z(n13036) );
  NOR U12957 ( .A(n13044), .B(n13045), .Z(n13043) );
  XOR U12958 ( .A(n13042), .B(n13046), .Z(n13044) );
  XNOR U12959 ( .A(n13003), .B(n13010), .Z(n13024) );
  NOR U12960 ( .A(n12967), .B(n13047), .Z(n13010) );
  XOR U12961 ( .A(n13015), .B(n13014), .Z(n13003) );
  XNOR U12962 ( .A(n13048), .B(n13011), .Z(n13014) );
  XOR U12963 ( .A(n13049), .B(n13050), .Z(n13011) );
  AND U12964 ( .A(n13051), .B(n13052), .Z(n13050) );
  XOR U12965 ( .A(n13049), .B(n13053), .Z(n13051) );
  XNOR U12966 ( .A(n13054), .B(n13055), .Z(n13048) );
  NOR U12967 ( .A(n13056), .B(n13057), .Z(n13055) );
  XNOR U12968 ( .A(n13054), .B(n13058), .Z(n13056) );
  XOR U12969 ( .A(n13059), .B(n13060), .Z(n13015) );
  NOR U12970 ( .A(n13061), .B(n13062), .Z(n13060) );
  XNOR U12971 ( .A(n13059), .B(n13063), .Z(n13061) );
  XNOR U12972 ( .A(n12952), .B(n13020), .Z(n13022) );
  XOR U12973 ( .A(n13064), .B(n13065), .Z(n12952) );
  AND U12974 ( .A(n247), .B(n13066), .Z(n13065) );
  XOR U12975 ( .A(n13067), .B(n13064), .Z(n13066) );
  AND U12976 ( .A(n12964), .B(n12967), .Z(n13020) );
  XOR U12977 ( .A(n13068), .B(n13047), .Z(n12967) );
  XNOR U12978 ( .A(p_input[2048]), .B(p_input[960]), .Z(n13047) );
  XOR U12979 ( .A(n13035), .B(n13034), .Z(n13068) );
  XNOR U12980 ( .A(n13069), .B(n13041), .Z(n13034) );
  XNOR U12981 ( .A(n13030), .B(n13029), .Z(n13041) );
  XOR U12982 ( .A(n13070), .B(n13026), .Z(n13029) );
  XNOR U12983 ( .A(n6439), .B(p_input[970]), .Z(n13026) );
  XNOR U12984 ( .A(p_input[2059]), .B(p_input[971]), .Z(n13070) );
  XOR U12985 ( .A(p_input[2060]), .B(p_input[972]), .Z(n13030) );
  XNOR U12986 ( .A(n13040), .B(n13031), .Z(n13069) );
  XNOR U12987 ( .A(n6553), .B(p_input[961]), .Z(n13031) );
  XOR U12988 ( .A(n13071), .B(n13046), .Z(n13040) );
  XNOR U12989 ( .A(p_input[2063]), .B(p_input[975]), .Z(n13046) );
  XOR U12990 ( .A(n13037), .B(n13045), .Z(n13071) );
  XOR U12991 ( .A(n13072), .B(n13042), .Z(n13045) );
  XOR U12992 ( .A(p_input[2061]), .B(p_input[973]), .Z(n13042) );
  XNOR U12993 ( .A(p_input[2062]), .B(p_input[974]), .Z(n13072) );
  XNOR U12994 ( .A(n6325), .B(p_input[969]), .Z(n13037) );
  XNOR U12995 ( .A(n13053), .B(n13052), .Z(n13035) );
  XNOR U12996 ( .A(n13073), .B(n13058), .Z(n13052) );
  XOR U12997 ( .A(p_input[2056]), .B(p_input[968]), .Z(n13058) );
  XOR U12998 ( .A(n13049), .B(n13057), .Z(n13073) );
  XOR U12999 ( .A(n13074), .B(n13054), .Z(n13057) );
  XOR U13000 ( .A(p_input[2054]), .B(p_input[966]), .Z(n13054) );
  XNOR U13001 ( .A(p_input[2055]), .B(p_input[967]), .Z(n13074) );
  XNOR U13002 ( .A(n6328), .B(p_input[962]), .Z(n13049) );
  XNOR U13003 ( .A(n13063), .B(n13062), .Z(n13053) );
  XOR U13004 ( .A(n13075), .B(n13059), .Z(n13062) );
  XOR U13005 ( .A(p_input[2051]), .B(p_input[963]), .Z(n13059) );
  XNOR U13006 ( .A(p_input[2052]), .B(p_input[964]), .Z(n13075) );
  XOR U13007 ( .A(p_input[2053]), .B(p_input[965]), .Z(n13063) );
  XOR U13008 ( .A(n13076), .B(n13077), .Z(n12964) );
  AND U13009 ( .A(n247), .B(n13078), .Z(n13077) );
  XNOR U13010 ( .A(n13079), .B(n13076), .Z(n13078) );
  XNOR U13011 ( .A(n13080), .B(n13081), .Z(n247) );
  AND U13012 ( .A(n13082), .B(n13083), .Z(n13081) );
  XOR U13013 ( .A(n12977), .B(n13080), .Z(n13083) );
  AND U13014 ( .A(n13084), .B(n13085), .Z(n12977) );
  XNOR U13015 ( .A(n12974), .B(n13080), .Z(n13082) );
  XOR U13016 ( .A(n13086), .B(n13087), .Z(n12974) );
  AND U13017 ( .A(n251), .B(n13088), .Z(n13087) );
  XOR U13018 ( .A(n13089), .B(n13086), .Z(n13088) );
  XOR U13019 ( .A(n13090), .B(n13091), .Z(n13080) );
  AND U13020 ( .A(n13092), .B(n13093), .Z(n13091) );
  XNOR U13021 ( .A(n13090), .B(n13084), .Z(n13093) );
  IV U13022 ( .A(n12992), .Z(n13084) );
  XOR U13023 ( .A(n13094), .B(n13095), .Z(n12992) );
  XOR U13024 ( .A(n13096), .B(n13085), .Z(n13095) );
  AND U13025 ( .A(n13019), .B(n13097), .Z(n13085) );
  AND U13026 ( .A(n13098), .B(n13099), .Z(n13096) );
  XOR U13027 ( .A(n13100), .B(n13094), .Z(n13098) );
  XNOR U13028 ( .A(n12989), .B(n13090), .Z(n13092) );
  XOR U13029 ( .A(n13101), .B(n13102), .Z(n12989) );
  AND U13030 ( .A(n251), .B(n13103), .Z(n13102) );
  XOR U13031 ( .A(n13104), .B(n13101), .Z(n13103) );
  XOR U13032 ( .A(n13105), .B(n13106), .Z(n13090) );
  AND U13033 ( .A(n13107), .B(n13108), .Z(n13106) );
  XNOR U13034 ( .A(n13105), .B(n13019), .Z(n13108) );
  XOR U13035 ( .A(n13109), .B(n13099), .Z(n13019) );
  XNOR U13036 ( .A(n13110), .B(n13094), .Z(n13099) );
  XOR U13037 ( .A(n13111), .B(n13112), .Z(n13094) );
  AND U13038 ( .A(n13113), .B(n13114), .Z(n13112) );
  XOR U13039 ( .A(n13115), .B(n13111), .Z(n13113) );
  XNOR U13040 ( .A(n13116), .B(n13117), .Z(n13110) );
  AND U13041 ( .A(n13118), .B(n13119), .Z(n13117) );
  XOR U13042 ( .A(n13116), .B(n13120), .Z(n13118) );
  XNOR U13043 ( .A(n13100), .B(n13097), .Z(n13109) );
  AND U13044 ( .A(n13121), .B(n13122), .Z(n13097) );
  XOR U13045 ( .A(n13123), .B(n13124), .Z(n13100) );
  AND U13046 ( .A(n13125), .B(n13126), .Z(n13124) );
  XOR U13047 ( .A(n13123), .B(n13127), .Z(n13125) );
  XNOR U13048 ( .A(n13016), .B(n13105), .Z(n13107) );
  XOR U13049 ( .A(n13128), .B(n13129), .Z(n13016) );
  AND U13050 ( .A(n251), .B(n13130), .Z(n13129) );
  XNOR U13051 ( .A(n13131), .B(n13128), .Z(n13130) );
  XOR U13052 ( .A(n13132), .B(n13133), .Z(n13105) );
  AND U13053 ( .A(n13134), .B(n13135), .Z(n13133) );
  XNOR U13054 ( .A(n13132), .B(n13121), .Z(n13135) );
  IV U13055 ( .A(n13067), .Z(n13121) );
  XNOR U13056 ( .A(n13136), .B(n13114), .Z(n13067) );
  XNOR U13057 ( .A(n13137), .B(n13120), .Z(n13114) );
  XOR U13058 ( .A(n13138), .B(n13139), .Z(n13120) );
  NOR U13059 ( .A(n13140), .B(n13141), .Z(n13139) );
  XNOR U13060 ( .A(n13138), .B(n13142), .Z(n13140) );
  XNOR U13061 ( .A(n13119), .B(n13111), .Z(n13137) );
  XOR U13062 ( .A(n13143), .B(n13144), .Z(n13111) );
  AND U13063 ( .A(n13145), .B(n13146), .Z(n13144) );
  XNOR U13064 ( .A(n13143), .B(n13147), .Z(n13145) );
  XNOR U13065 ( .A(n13148), .B(n13116), .Z(n13119) );
  XOR U13066 ( .A(n13149), .B(n13150), .Z(n13116) );
  AND U13067 ( .A(n13151), .B(n13152), .Z(n13150) );
  XOR U13068 ( .A(n13149), .B(n13153), .Z(n13151) );
  XNOR U13069 ( .A(n13154), .B(n13155), .Z(n13148) );
  NOR U13070 ( .A(n13156), .B(n13157), .Z(n13155) );
  XOR U13071 ( .A(n13154), .B(n13158), .Z(n13156) );
  XNOR U13072 ( .A(n13115), .B(n13122), .Z(n13136) );
  NOR U13073 ( .A(n13079), .B(n13159), .Z(n13122) );
  XOR U13074 ( .A(n13127), .B(n13126), .Z(n13115) );
  XNOR U13075 ( .A(n13160), .B(n13123), .Z(n13126) );
  XOR U13076 ( .A(n13161), .B(n13162), .Z(n13123) );
  AND U13077 ( .A(n13163), .B(n13164), .Z(n13162) );
  XOR U13078 ( .A(n13161), .B(n13165), .Z(n13163) );
  XNOR U13079 ( .A(n13166), .B(n13167), .Z(n13160) );
  NOR U13080 ( .A(n13168), .B(n13169), .Z(n13167) );
  XNOR U13081 ( .A(n13166), .B(n13170), .Z(n13168) );
  XOR U13082 ( .A(n13171), .B(n13172), .Z(n13127) );
  NOR U13083 ( .A(n13173), .B(n13174), .Z(n13172) );
  XNOR U13084 ( .A(n13171), .B(n13175), .Z(n13173) );
  XNOR U13085 ( .A(n13064), .B(n13132), .Z(n13134) );
  XOR U13086 ( .A(n13176), .B(n13177), .Z(n13064) );
  AND U13087 ( .A(n251), .B(n13178), .Z(n13177) );
  XOR U13088 ( .A(n13179), .B(n13176), .Z(n13178) );
  AND U13089 ( .A(n13076), .B(n13079), .Z(n13132) );
  XOR U13090 ( .A(n13180), .B(n13159), .Z(n13079) );
  XNOR U13091 ( .A(p_input[2048]), .B(p_input[976]), .Z(n13159) );
  XOR U13092 ( .A(n13147), .B(n13146), .Z(n13180) );
  XNOR U13093 ( .A(n13181), .B(n13153), .Z(n13146) );
  XNOR U13094 ( .A(n13142), .B(n13141), .Z(n13153) );
  XOR U13095 ( .A(n13182), .B(n13138), .Z(n13141) );
  XNOR U13096 ( .A(n6439), .B(p_input[986]), .Z(n13138) );
  XNOR U13097 ( .A(p_input[2059]), .B(p_input[987]), .Z(n13182) );
  XOR U13098 ( .A(p_input[2060]), .B(p_input[988]), .Z(n13142) );
  XNOR U13099 ( .A(n13152), .B(n13143), .Z(n13181) );
  XNOR U13100 ( .A(n6553), .B(p_input[977]), .Z(n13143) );
  XOR U13101 ( .A(n13183), .B(n13158), .Z(n13152) );
  XNOR U13102 ( .A(p_input[2063]), .B(p_input[991]), .Z(n13158) );
  XOR U13103 ( .A(n13149), .B(n13157), .Z(n13183) );
  XOR U13104 ( .A(n13184), .B(n13154), .Z(n13157) );
  XOR U13105 ( .A(p_input[2061]), .B(p_input[989]), .Z(n13154) );
  XNOR U13106 ( .A(p_input[2062]), .B(p_input[990]), .Z(n13184) );
  XNOR U13107 ( .A(n6325), .B(p_input[985]), .Z(n13149) );
  XNOR U13108 ( .A(n13165), .B(n13164), .Z(n13147) );
  XNOR U13109 ( .A(n13185), .B(n13170), .Z(n13164) );
  XOR U13110 ( .A(p_input[2056]), .B(p_input[984]), .Z(n13170) );
  XOR U13111 ( .A(n13161), .B(n13169), .Z(n13185) );
  XOR U13112 ( .A(n13186), .B(n13166), .Z(n13169) );
  XOR U13113 ( .A(p_input[2054]), .B(p_input[982]), .Z(n13166) );
  XNOR U13114 ( .A(p_input[2055]), .B(p_input[983]), .Z(n13186) );
  XNOR U13115 ( .A(n6328), .B(p_input[978]), .Z(n13161) );
  XNOR U13116 ( .A(n13175), .B(n13174), .Z(n13165) );
  XOR U13117 ( .A(n13187), .B(n13171), .Z(n13174) );
  XOR U13118 ( .A(p_input[2051]), .B(p_input[979]), .Z(n13171) );
  XNOR U13119 ( .A(p_input[2052]), .B(p_input[980]), .Z(n13187) );
  XOR U13120 ( .A(p_input[2053]), .B(p_input[981]), .Z(n13175) );
  XOR U13121 ( .A(n13188), .B(n13189), .Z(n13076) );
  AND U13122 ( .A(n251), .B(n13190), .Z(n13189) );
  XNOR U13123 ( .A(n13191), .B(n13188), .Z(n13190) );
  XNOR U13124 ( .A(n13192), .B(n13193), .Z(n251) );
  AND U13125 ( .A(n13194), .B(n13195), .Z(n13193) );
  XOR U13126 ( .A(n13089), .B(n13192), .Z(n13195) );
  AND U13127 ( .A(n13196), .B(n13197), .Z(n13089) );
  XNOR U13128 ( .A(n13086), .B(n13192), .Z(n13194) );
  XOR U13129 ( .A(n13198), .B(n13199), .Z(n13086) );
  AND U13130 ( .A(n255), .B(n13200), .Z(n13199) );
  XOR U13131 ( .A(n13201), .B(n13198), .Z(n13200) );
  XOR U13132 ( .A(n13202), .B(n13203), .Z(n13192) );
  AND U13133 ( .A(n13204), .B(n13205), .Z(n13203) );
  XNOR U13134 ( .A(n13202), .B(n13196), .Z(n13205) );
  IV U13135 ( .A(n13104), .Z(n13196) );
  XOR U13136 ( .A(n13206), .B(n13207), .Z(n13104) );
  XOR U13137 ( .A(n13208), .B(n13197), .Z(n13207) );
  AND U13138 ( .A(n13131), .B(n13209), .Z(n13197) );
  AND U13139 ( .A(n13210), .B(n13211), .Z(n13208) );
  XOR U13140 ( .A(n13212), .B(n13206), .Z(n13210) );
  XNOR U13141 ( .A(n13101), .B(n13202), .Z(n13204) );
  XOR U13142 ( .A(n13213), .B(n13214), .Z(n13101) );
  AND U13143 ( .A(n255), .B(n13215), .Z(n13214) );
  XOR U13144 ( .A(n13216), .B(n13213), .Z(n13215) );
  XOR U13145 ( .A(n13217), .B(n13218), .Z(n13202) );
  AND U13146 ( .A(n13219), .B(n13220), .Z(n13218) );
  XNOR U13147 ( .A(n13217), .B(n13131), .Z(n13220) );
  XOR U13148 ( .A(n13221), .B(n13211), .Z(n13131) );
  XNOR U13149 ( .A(n13222), .B(n13206), .Z(n13211) );
  XOR U13150 ( .A(n13223), .B(n13224), .Z(n13206) );
  AND U13151 ( .A(n13225), .B(n13226), .Z(n13224) );
  XOR U13152 ( .A(n13227), .B(n13223), .Z(n13225) );
  XNOR U13153 ( .A(n13228), .B(n13229), .Z(n13222) );
  AND U13154 ( .A(n13230), .B(n13231), .Z(n13229) );
  XOR U13155 ( .A(n13228), .B(n13232), .Z(n13230) );
  XNOR U13156 ( .A(n13212), .B(n13209), .Z(n13221) );
  AND U13157 ( .A(n13233), .B(n13234), .Z(n13209) );
  XOR U13158 ( .A(n13235), .B(n13236), .Z(n13212) );
  AND U13159 ( .A(n13237), .B(n13238), .Z(n13236) );
  XOR U13160 ( .A(n13235), .B(n13239), .Z(n13237) );
  XNOR U13161 ( .A(n13128), .B(n13217), .Z(n13219) );
  XOR U13162 ( .A(n13240), .B(n13241), .Z(n13128) );
  AND U13163 ( .A(n255), .B(n13242), .Z(n13241) );
  XNOR U13164 ( .A(n13243), .B(n13240), .Z(n13242) );
  XOR U13165 ( .A(n13244), .B(n13245), .Z(n13217) );
  AND U13166 ( .A(n13246), .B(n13247), .Z(n13245) );
  XNOR U13167 ( .A(n13244), .B(n13233), .Z(n13247) );
  IV U13168 ( .A(n13179), .Z(n13233) );
  XNOR U13169 ( .A(n13248), .B(n13226), .Z(n13179) );
  XNOR U13170 ( .A(n13249), .B(n13232), .Z(n13226) );
  XNOR U13171 ( .A(n13250), .B(n13251), .Z(n13232) );
  NOR U13172 ( .A(n13252), .B(n13253), .Z(n13251) );
  XOR U13173 ( .A(n13250), .B(n13254), .Z(n13252) );
  XNOR U13174 ( .A(n13231), .B(n13223), .Z(n13249) );
  XOR U13175 ( .A(n13255), .B(n13256), .Z(n13223) );
  AND U13176 ( .A(n13257), .B(n13258), .Z(n13256) );
  XOR U13177 ( .A(n13255), .B(n13259), .Z(n13257) );
  XNOR U13178 ( .A(n13260), .B(n13228), .Z(n13231) );
  XOR U13179 ( .A(n13261), .B(n13262), .Z(n13228) );
  AND U13180 ( .A(n13263), .B(n13264), .Z(n13262) );
  XNOR U13181 ( .A(n13265), .B(n13266), .Z(n13263) );
  IV U13182 ( .A(n13261), .Z(n13265) );
  XNOR U13183 ( .A(n13267), .B(n13268), .Z(n13260) );
  NOR U13184 ( .A(n13269), .B(n13270), .Z(n13268) );
  XNOR U13185 ( .A(n13267), .B(n13271), .Z(n13269) );
  XNOR U13186 ( .A(n13227), .B(n13234), .Z(n13248) );
  NOR U13187 ( .A(n13191), .B(n13272), .Z(n13234) );
  XOR U13188 ( .A(n13239), .B(n13238), .Z(n13227) );
  XNOR U13189 ( .A(n13273), .B(n13235), .Z(n13238) );
  XOR U13190 ( .A(n13274), .B(n13275), .Z(n13235) );
  AND U13191 ( .A(n13276), .B(n13277), .Z(n13275) );
  XOR U13192 ( .A(n13274), .B(n13278), .Z(n13276) );
  XNOR U13193 ( .A(n13279), .B(n13280), .Z(n13273) );
  NOR U13194 ( .A(n13281), .B(n13282), .Z(n13280) );
  XNOR U13195 ( .A(n13279), .B(n13283), .Z(n13281) );
  XOR U13196 ( .A(n13284), .B(n13285), .Z(n13239) );
  NOR U13197 ( .A(n13286), .B(n13287), .Z(n13285) );
  XNOR U13198 ( .A(n13284), .B(n13288), .Z(n13286) );
  XNOR U13199 ( .A(n13176), .B(n13244), .Z(n13246) );
  XOR U13200 ( .A(n13289), .B(n13290), .Z(n13176) );
  AND U13201 ( .A(n255), .B(n13291), .Z(n13290) );
  XOR U13202 ( .A(n13292), .B(n13289), .Z(n13291) );
  AND U13203 ( .A(n13188), .B(n13191), .Z(n13244) );
  XOR U13204 ( .A(n13293), .B(n13272), .Z(n13191) );
  XNOR U13205 ( .A(p_input[2048]), .B(p_input[992]), .Z(n13272) );
  XNOR U13206 ( .A(n13259), .B(n13258), .Z(n13293) );
  XNOR U13207 ( .A(n13294), .B(n13266), .Z(n13258) );
  XNOR U13208 ( .A(n13254), .B(n13253), .Z(n13266) );
  XNOR U13209 ( .A(n13295), .B(n13250), .Z(n13253) );
  XNOR U13210 ( .A(p_input[1002]), .B(p_input[2058]), .Z(n13250) );
  XOR U13211 ( .A(p_input[1003]), .B(n6319), .Z(n13295) );
  XOR U13212 ( .A(p_input[1004]), .B(p_input[2060]), .Z(n13254) );
  XNOR U13213 ( .A(n13264), .B(n13255), .Z(n13294) );
  XNOR U13214 ( .A(n6553), .B(p_input[993]), .Z(n13255) );
  XNOR U13215 ( .A(n13296), .B(n13271), .Z(n13264) );
  XNOR U13216 ( .A(p_input[1007]), .B(n6322), .Z(n13271) );
  XOR U13217 ( .A(n13261), .B(n13270), .Z(n13296) );
  XOR U13218 ( .A(n13297), .B(n13267), .Z(n13270) );
  XOR U13219 ( .A(p_input[1005]), .B(p_input[2061]), .Z(n13267) );
  XOR U13220 ( .A(p_input[1006]), .B(n6324), .Z(n13297) );
  XOR U13221 ( .A(p_input[1001]), .B(p_input[2057]), .Z(n13261) );
  XOR U13222 ( .A(n13278), .B(n13277), .Z(n13259) );
  XNOR U13223 ( .A(n13298), .B(n13283), .Z(n13277) );
  XOR U13224 ( .A(p_input[1000]), .B(p_input[2056]), .Z(n13283) );
  XOR U13225 ( .A(n13274), .B(n13282), .Z(n13298) );
  XOR U13226 ( .A(n13299), .B(n13279), .Z(n13282) );
  XOR U13227 ( .A(p_input[2054]), .B(p_input[998]), .Z(n13279) );
  XNOR U13228 ( .A(p_input[2055]), .B(p_input[999]), .Z(n13299) );
  XNOR U13229 ( .A(n6328), .B(p_input[994]), .Z(n13274) );
  XNOR U13230 ( .A(n13288), .B(n13287), .Z(n13278) );
  XOR U13231 ( .A(n13300), .B(n13284), .Z(n13287) );
  XOR U13232 ( .A(p_input[2051]), .B(p_input[995]), .Z(n13284) );
  XNOR U13233 ( .A(p_input[2052]), .B(p_input[996]), .Z(n13300) );
  XOR U13234 ( .A(p_input[2053]), .B(p_input[997]), .Z(n13288) );
  XOR U13235 ( .A(n13301), .B(n13302), .Z(n13188) );
  AND U13236 ( .A(n255), .B(n13303), .Z(n13302) );
  XNOR U13237 ( .A(n13304), .B(n13301), .Z(n13303) );
  XNOR U13238 ( .A(n13305), .B(n13306), .Z(n255) );
  AND U13239 ( .A(n13307), .B(n13308), .Z(n13306) );
  XOR U13240 ( .A(n13201), .B(n13305), .Z(n13308) );
  AND U13241 ( .A(n13309), .B(n13310), .Z(n13201) );
  XNOR U13242 ( .A(n13198), .B(n13305), .Z(n13307) );
  XOR U13243 ( .A(n13311), .B(n13312), .Z(n13198) );
  AND U13244 ( .A(n259), .B(n13313), .Z(n13312) );
  XOR U13245 ( .A(n13314), .B(n13311), .Z(n13313) );
  XOR U13246 ( .A(n13315), .B(n13316), .Z(n13305) );
  AND U13247 ( .A(n13317), .B(n13318), .Z(n13316) );
  XNOR U13248 ( .A(n13315), .B(n13309), .Z(n13318) );
  IV U13249 ( .A(n13216), .Z(n13309) );
  XOR U13250 ( .A(n13319), .B(n13320), .Z(n13216) );
  XOR U13251 ( .A(n13321), .B(n13310), .Z(n13320) );
  AND U13252 ( .A(n13243), .B(n13322), .Z(n13310) );
  AND U13253 ( .A(n13323), .B(n13324), .Z(n13321) );
  XOR U13254 ( .A(n13325), .B(n13319), .Z(n13323) );
  XNOR U13255 ( .A(n13213), .B(n13315), .Z(n13317) );
  XOR U13256 ( .A(n13326), .B(n13327), .Z(n13213) );
  AND U13257 ( .A(n259), .B(n13328), .Z(n13327) );
  XOR U13258 ( .A(n13329), .B(n13326), .Z(n13328) );
  XOR U13259 ( .A(n13330), .B(n13331), .Z(n13315) );
  AND U13260 ( .A(n13332), .B(n13333), .Z(n13331) );
  XNOR U13261 ( .A(n13330), .B(n13243), .Z(n13333) );
  XOR U13262 ( .A(n13334), .B(n13324), .Z(n13243) );
  XNOR U13263 ( .A(n13335), .B(n13319), .Z(n13324) );
  XOR U13264 ( .A(n13336), .B(n13337), .Z(n13319) );
  AND U13265 ( .A(n13338), .B(n13339), .Z(n13337) );
  XOR U13266 ( .A(n13340), .B(n13336), .Z(n13338) );
  XNOR U13267 ( .A(n13341), .B(n13342), .Z(n13335) );
  AND U13268 ( .A(n13343), .B(n13344), .Z(n13342) );
  XOR U13269 ( .A(n13341), .B(n13345), .Z(n13343) );
  XNOR U13270 ( .A(n13325), .B(n13322), .Z(n13334) );
  AND U13271 ( .A(n13346), .B(n13347), .Z(n13322) );
  XOR U13272 ( .A(n13348), .B(n13349), .Z(n13325) );
  AND U13273 ( .A(n13350), .B(n13351), .Z(n13349) );
  XOR U13274 ( .A(n13348), .B(n13352), .Z(n13350) );
  XNOR U13275 ( .A(n13240), .B(n13330), .Z(n13332) );
  XOR U13276 ( .A(n13353), .B(n13354), .Z(n13240) );
  AND U13277 ( .A(n259), .B(n13355), .Z(n13354) );
  XNOR U13278 ( .A(n13356), .B(n13353), .Z(n13355) );
  XOR U13279 ( .A(n13357), .B(n13358), .Z(n13330) );
  AND U13280 ( .A(n13359), .B(n13360), .Z(n13358) );
  XNOR U13281 ( .A(n13357), .B(n13346), .Z(n13360) );
  IV U13282 ( .A(n13292), .Z(n13346) );
  XNOR U13283 ( .A(n13361), .B(n13339), .Z(n13292) );
  XNOR U13284 ( .A(n13362), .B(n13345), .Z(n13339) );
  XNOR U13285 ( .A(n13363), .B(n13364), .Z(n13345) );
  NOR U13286 ( .A(n13365), .B(n13366), .Z(n13364) );
  XOR U13287 ( .A(n13363), .B(n13367), .Z(n13365) );
  XNOR U13288 ( .A(n13344), .B(n13336), .Z(n13362) );
  XOR U13289 ( .A(n13368), .B(n13369), .Z(n13336) );
  AND U13290 ( .A(n13370), .B(n13371), .Z(n13369) );
  XOR U13291 ( .A(n13368), .B(n13372), .Z(n13370) );
  XNOR U13292 ( .A(n13373), .B(n13341), .Z(n13344) );
  XOR U13293 ( .A(n13374), .B(n13375), .Z(n13341) );
  AND U13294 ( .A(n13376), .B(n13377), .Z(n13375) );
  XNOR U13295 ( .A(n13378), .B(n13379), .Z(n13376) );
  IV U13296 ( .A(n13374), .Z(n13378) );
  XNOR U13297 ( .A(n13380), .B(n13381), .Z(n13373) );
  NOR U13298 ( .A(n13382), .B(n13383), .Z(n13381) );
  XNOR U13299 ( .A(n13380), .B(n13384), .Z(n13382) );
  XNOR U13300 ( .A(n13340), .B(n13347), .Z(n13361) );
  NOR U13301 ( .A(n13304), .B(n13385), .Z(n13347) );
  XOR U13302 ( .A(n13352), .B(n13351), .Z(n13340) );
  XNOR U13303 ( .A(n13386), .B(n13348), .Z(n13351) );
  XOR U13304 ( .A(n13387), .B(n13388), .Z(n13348) );
  AND U13305 ( .A(n13389), .B(n13390), .Z(n13388) );
  XNOR U13306 ( .A(n13391), .B(n13392), .Z(n13389) );
  IV U13307 ( .A(n13387), .Z(n13391) );
  XNOR U13308 ( .A(n13393), .B(n13394), .Z(n13386) );
  NOR U13309 ( .A(n13395), .B(n13396), .Z(n13394) );
  XNOR U13310 ( .A(n13393), .B(n13397), .Z(n13395) );
  XOR U13311 ( .A(n13398), .B(n13399), .Z(n13352) );
  NOR U13312 ( .A(n13400), .B(n13401), .Z(n13399) );
  XNOR U13313 ( .A(n13398), .B(n13402), .Z(n13400) );
  XNOR U13314 ( .A(n13289), .B(n13357), .Z(n13359) );
  XOR U13315 ( .A(n13403), .B(n13404), .Z(n13289) );
  AND U13316 ( .A(n259), .B(n13405), .Z(n13404) );
  XOR U13317 ( .A(n13406), .B(n13403), .Z(n13405) );
  AND U13318 ( .A(n13301), .B(n13304), .Z(n13357) );
  XOR U13319 ( .A(n13407), .B(n13385), .Z(n13304) );
  XNOR U13320 ( .A(p_input[1008]), .B(p_input[2048]), .Z(n13385) );
  XNOR U13321 ( .A(n13372), .B(n13371), .Z(n13407) );
  XNOR U13322 ( .A(n13408), .B(n13379), .Z(n13371) );
  XNOR U13323 ( .A(n13367), .B(n13366), .Z(n13379) );
  XNOR U13324 ( .A(n13409), .B(n13363), .Z(n13366) );
  XNOR U13325 ( .A(p_input[1018]), .B(p_input[2058]), .Z(n13363) );
  XOR U13326 ( .A(p_input[1019]), .B(n6319), .Z(n13409) );
  XOR U13327 ( .A(p_input[1020]), .B(p_input[2060]), .Z(n13367) );
  XOR U13328 ( .A(n13377), .B(n13410), .Z(n13408) );
  IV U13329 ( .A(n13368), .Z(n13410) );
  XOR U13330 ( .A(p_input[1009]), .B(p_input[2049]), .Z(n13368) );
  XNOR U13331 ( .A(n13411), .B(n13384), .Z(n13377) );
  XNOR U13332 ( .A(p_input[1023]), .B(n6322), .Z(n13384) );
  XOR U13333 ( .A(n13374), .B(n13383), .Z(n13411) );
  XOR U13334 ( .A(n13412), .B(n13380), .Z(n13383) );
  XOR U13335 ( .A(p_input[1021]), .B(p_input[2061]), .Z(n13380) );
  XOR U13336 ( .A(p_input[1022]), .B(n6324), .Z(n13412) );
  XOR U13337 ( .A(p_input[1017]), .B(p_input[2057]), .Z(n13374) );
  XOR U13338 ( .A(n13392), .B(n13390), .Z(n13372) );
  XNOR U13339 ( .A(n13413), .B(n13397), .Z(n13390) );
  XOR U13340 ( .A(p_input[1016]), .B(p_input[2056]), .Z(n13397) );
  XOR U13341 ( .A(n13387), .B(n13396), .Z(n13413) );
  XOR U13342 ( .A(n13414), .B(n13393), .Z(n13396) );
  XOR U13343 ( .A(p_input[1014]), .B(p_input[2054]), .Z(n13393) );
  XOR U13344 ( .A(p_input[1015]), .B(n7007), .Z(n13414) );
  XOR U13345 ( .A(p_input[1010]), .B(p_input[2050]), .Z(n13387) );
  XNOR U13346 ( .A(n13402), .B(n13401), .Z(n13392) );
  XOR U13347 ( .A(n13415), .B(n13398), .Z(n13401) );
  XOR U13348 ( .A(p_input[1011]), .B(p_input[2051]), .Z(n13398) );
  XOR U13349 ( .A(p_input[1012]), .B(n7009), .Z(n13415) );
  XOR U13350 ( .A(p_input[1013]), .B(p_input[2053]), .Z(n13402) );
  XOR U13351 ( .A(n13416), .B(n13417), .Z(n13301) );
  AND U13352 ( .A(n259), .B(n13418), .Z(n13417) );
  XNOR U13353 ( .A(n13419), .B(n13416), .Z(n13418) );
  XNOR U13354 ( .A(n13420), .B(n13421), .Z(n259) );
  AND U13355 ( .A(n13422), .B(n13423), .Z(n13421) );
  XOR U13356 ( .A(n13314), .B(n13420), .Z(n13423) );
  AND U13357 ( .A(n13424), .B(n13425), .Z(n13314) );
  XNOR U13358 ( .A(n13311), .B(n13420), .Z(n13422) );
  XOR U13359 ( .A(n13426), .B(n13427), .Z(n13311) );
  AND U13360 ( .A(n263), .B(n13428), .Z(n13427) );
  XOR U13361 ( .A(n13429), .B(n13426), .Z(n13428) );
  XOR U13362 ( .A(n13430), .B(n13431), .Z(n13420) );
  AND U13363 ( .A(n13432), .B(n13433), .Z(n13431) );
  XNOR U13364 ( .A(n13430), .B(n13424), .Z(n13433) );
  IV U13365 ( .A(n13329), .Z(n13424) );
  XOR U13366 ( .A(n13434), .B(n13435), .Z(n13329) );
  XOR U13367 ( .A(n13436), .B(n13425), .Z(n13435) );
  AND U13368 ( .A(n13356), .B(n13437), .Z(n13425) );
  AND U13369 ( .A(n13438), .B(n13439), .Z(n13436) );
  XOR U13370 ( .A(n13440), .B(n13434), .Z(n13438) );
  XNOR U13371 ( .A(n13326), .B(n13430), .Z(n13432) );
  XOR U13372 ( .A(n13441), .B(n13442), .Z(n13326) );
  AND U13373 ( .A(n263), .B(n13443), .Z(n13442) );
  XOR U13374 ( .A(n13444), .B(n13441), .Z(n13443) );
  XOR U13375 ( .A(n13445), .B(n13446), .Z(n13430) );
  AND U13376 ( .A(n13447), .B(n13448), .Z(n13446) );
  XNOR U13377 ( .A(n13445), .B(n13356), .Z(n13448) );
  XOR U13378 ( .A(n13449), .B(n13439), .Z(n13356) );
  XNOR U13379 ( .A(n13450), .B(n13434), .Z(n13439) );
  XOR U13380 ( .A(n13451), .B(n13452), .Z(n13434) );
  AND U13381 ( .A(n13453), .B(n13454), .Z(n13452) );
  XOR U13382 ( .A(n13455), .B(n13451), .Z(n13453) );
  XNOR U13383 ( .A(n13456), .B(n13457), .Z(n13450) );
  AND U13384 ( .A(n13458), .B(n13459), .Z(n13457) );
  XOR U13385 ( .A(n13456), .B(n13460), .Z(n13458) );
  XNOR U13386 ( .A(n13440), .B(n13437), .Z(n13449) );
  AND U13387 ( .A(n13461), .B(n13462), .Z(n13437) );
  XOR U13388 ( .A(n13463), .B(n13464), .Z(n13440) );
  AND U13389 ( .A(n13465), .B(n13466), .Z(n13464) );
  XOR U13390 ( .A(n13463), .B(n13467), .Z(n13465) );
  XNOR U13391 ( .A(n13353), .B(n13445), .Z(n13447) );
  XOR U13392 ( .A(n13468), .B(n13469), .Z(n13353) );
  AND U13393 ( .A(n263), .B(n13470), .Z(n13469) );
  XNOR U13394 ( .A(n13471), .B(n13468), .Z(n13470) );
  XOR U13395 ( .A(n13472), .B(n13473), .Z(n13445) );
  AND U13396 ( .A(n13474), .B(n13475), .Z(n13473) );
  XNOR U13397 ( .A(n13472), .B(n13461), .Z(n13475) );
  IV U13398 ( .A(n13406), .Z(n13461) );
  XNOR U13399 ( .A(n13476), .B(n13454), .Z(n13406) );
  XNOR U13400 ( .A(n13477), .B(n13460), .Z(n13454) );
  XNOR U13401 ( .A(n13478), .B(n13479), .Z(n13460) );
  NOR U13402 ( .A(n13480), .B(n13481), .Z(n13479) );
  XOR U13403 ( .A(n13478), .B(n13482), .Z(n13480) );
  XNOR U13404 ( .A(n13459), .B(n13451), .Z(n13477) );
  XOR U13405 ( .A(n13483), .B(n13484), .Z(n13451) );
  AND U13406 ( .A(n13485), .B(n13486), .Z(n13484) );
  XOR U13407 ( .A(n13483), .B(n13487), .Z(n13485) );
  XNOR U13408 ( .A(n13488), .B(n13456), .Z(n13459) );
  XOR U13409 ( .A(n13489), .B(n13490), .Z(n13456) );
  AND U13410 ( .A(n13491), .B(n13492), .Z(n13490) );
  XNOR U13411 ( .A(n13493), .B(n13494), .Z(n13491) );
  IV U13412 ( .A(n13489), .Z(n13493) );
  XNOR U13413 ( .A(n13495), .B(n13496), .Z(n13488) );
  NOR U13414 ( .A(n13497), .B(n13498), .Z(n13496) );
  XNOR U13415 ( .A(n13495), .B(n13499), .Z(n13497) );
  XNOR U13416 ( .A(n13455), .B(n13462), .Z(n13476) );
  NOR U13417 ( .A(n13419), .B(n13500), .Z(n13462) );
  XOR U13418 ( .A(n13467), .B(n13466), .Z(n13455) );
  XNOR U13419 ( .A(n13501), .B(n13463), .Z(n13466) );
  XOR U13420 ( .A(n13502), .B(n13503), .Z(n13463) );
  AND U13421 ( .A(n13504), .B(n13505), .Z(n13503) );
  XNOR U13422 ( .A(n13506), .B(n13507), .Z(n13504) );
  IV U13423 ( .A(n13502), .Z(n13506) );
  XNOR U13424 ( .A(n13508), .B(n13509), .Z(n13501) );
  NOR U13425 ( .A(n13510), .B(n13511), .Z(n13509) );
  XNOR U13426 ( .A(n13508), .B(n13512), .Z(n13510) );
  XOR U13427 ( .A(n13513), .B(n13514), .Z(n13467) );
  NOR U13428 ( .A(n13515), .B(n13516), .Z(n13514) );
  XNOR U13429 ( .A(n13513), .B(n13517), .Z(n13515) );
  XNOR U13430 ( .A(n13403), .B(n13472), .Z(n13474) );
  XOR U13431 ( .A(n13518), .B(n13519), .Z(n13403) );
  AND U13432 ( .A(n263), .B(n13520), .Z(n13519) );
  XOR U13433 ( .A(n13521), .B(n13518), .Z(n13520) );
  AND U13434 ( .A(n13416), .B(n13419), .Z(n13472) );
  XOR U13435 ( .A(n13522), .B(n13500), .Z(n13419) );
  XNOR U13436 ( .A(p_input[1024]), .B(p_input[2048]), .Z(n13500) );
  XNOR U13437 ( .A(n13487), .B(n13486), .Z(n13522) );
  XNOR U13438 ( .A(n13523), .B(n13494), .Z(n13486) );
  XNOR U13439 ( .A(n13482), .B(n13481), .Z(n13494) );
  XNOR U13440 ( .A(n13524), .B(n13478), .Z(n13481) );
  XNOR U13441 ( .A(p_input[1034]), .B(p_input[2058]), .Z(n13478) );
  XOR U13442 ( .A(p_input[1035]), .B(n6319), .Z(n13524) );
  XOR U13443 ( .A(p_input[1036]), .B(p_input[2060]), .Z(n13482) );
  XOR U13444 ( .A(n13492), .B(n13525), .Z(n13523) );
  IV U13445 ( .A(n13483), .Z(n13525) );
  XOR U13446 ( .A(p_input[1025]), .B(p_input[2049]), .Z(n13483) );
  XNOR U13447 ( .A(n13526), .B(n13499), .Z(n13492) );
  XNOR U13448 ( .A(p_input[1039]), .B(n6322), .Z(n13499) );
  XOR U13449 ( .A(n13489), .B(n13498), .Z(n13526) );
  XOR U13450 ( .A(n13527), .B(n13495), .Z(n13498) );
  XOR U13451 ( .A(p_input[1037]), .B(p_input[2061]), .Z(n13495) );
  XOR U13452 ( .A(p_input[1038]), .B(n6324), .Z(n13527) );
  XOR U13453 ( .A(p_input[1033]), .B(p_input[2057]), .Z(n13489) );
  XOR U13454 ( .A(n13507), .B(n13505), .Z(n13487) );
  XNOR U13455 ( .A(n13528), .B(n13512), .Z(n13505) );
  XOR U13456 ( .A(p_input[1032]), .B(p_input[2056]), .Z(n13512) );
  XOR U13457 ( .A(n13502), .B(n13511), .Z(n13528) );
  XOR U13458 ( .A(n13529), .B(n13508), .Z(n13511) );
  XOR U13459 ( .A(p_input[1030]), .B(p_input[2054]), .Z(n13508) );
  XOR U13460 ( .A(p_input[1031]), .B(n7007), .Z(n13529) );
  XOR U13461 ( .A(p_input[1026]), .B(p_input[2050]), .Z(n13502) );
  XNOR U13462 ( .A(n13517), .B(n13516), .Z(n13507) );
  XOR U13463 ( .A(n13530), .B(n13513), .Z(n13516) );
  XOR U13464 ( .A(p_input[1027]), .B(p_input[2051]), .Z(n13513) );
  XOR U13465 ( .A(p_input[1028]), .B(n7009), .Z(n13530) );
  XOR U13466 ( .A(p_input[1029]), .B(p_input[2053]), .Z(n13517) );
  XOR U13467 ( .A(n13531), .B(n13532), .Z(n13416) );
  AND U13468 ( .A(n263), .B(n13533), .Z(n13532) );
  XNOR U13469 ( .A(n13534), .B(n13531), .Z(n13533) );
  XNOR U13470 ( .A(n13535), .B(n13536), .Z(n263) );
  AND U13471 ( .A(n13537), .B(n13538), .Z(n13536) );
  XOR U13472 ( .A(n13429), .B(n13535), .Z(n13538) );
  AND U13473 ( .A(n13539), .B(n13540), .Z(n13429) );
  XNOR U13474 ( .A(n13426), .B(n13535), .Z(n13537) );
  XOR U13475 ( .A(n13541), .B(n13542), .Z(n13426) );
  AND U13476 ( .A(n267), .B(n13543), .Z(n13542) );
  XOR U13477 ( .A(n13544), .B(n13541), .Z(n13543) );
  XOR U13478 ( .A(n13545), .B(n13546), .Z(n13535) );
  AND U13479 ( .A(n13547), .B(n13548), .Z(n13546) );
  XNOR U13480 ( .A(n13545), .B(n13539), .Z(n13548) );
  IV U13481 ( .A(n13444), .Z(n13539) );
  XOR U13482 ( .A(n13549), .B(n13550), .Z(n13444) );
  XOR U13483 ( .A(n13551), .B(n13540), .Z(n13550) );
  AND U13484 ( .A(n13471), .B(n13552), .Z(n13540) );
  AND U13485 ( .A(n13553), .B(n13554), .Z(n13551) );
  XOR U13486 ( .A(n13555), .B(n13549), .Z(n13553) );
  XNOR U13487 ( .A(n13441), .B(n13545), .Z(n13547) );
  XOR U13488 ( .A(n13556), .B(n13557), .Z(n13441) );
  AND U13489 ( .A(n267), .B(n13558), .Z(n13557) );
  XOR U13490 ( .A(n13559), .B(n13556), .Z(n13558) );
  XOR U13491 ( .A(n13560), .B(n13561), .Z(n13545) );
  AND U13492 ( .A(n13562), .B(n13563), .Z(n13561) );
  XNOR U13493 ( .A(n13560), .B(n13471), .Z(n13563) );
  XOR U13494 ( .A(n13564), .B(n13554), .Z(n13471) );
  XNOR U13495 ( .A(n13565), .B(n13549), .Z(n13554) );
  XOR U13496 ( .A(n13566), .B(n13567), .Z(n13549) );
  AND U13497 ( .A(n13568), .B(n13569), .Z(n13567) );
  XOR U13498 ( .A(n13570), .B(n13566), .Z(n13568) );
  XNOR U13499 ( .A(n13571), .B(n13572), .Z(n13565) );
  AND U13500 ( .A(n13573), .B(n13574), .Z(n13572) );
  XOR U13501 ( .A(n13571), .B(n13575), .Z(n13573) );
  XNOR U13502 ( .A(n13555), .B(n13552), .Z(n13564) );
  AND U13503 ( .A(n13576), .B(n13577), .Z(n13552) );
  XOR U13504 ( .A(n13578), .B(n13579), .Z(n13555) );
  AND U13505 ( .A(n13580), .B(n13581), .Z(n13579) );
  XOR U13506 ( .A(n13578), .B(n13582), .Z(n13580) );
  XNOR U13507 ( .A(n13468), .B(n13560), .Z(n13562) );
  XOR U13508 ( .A(n13583), .B(n13584), .Z(n13468) );
  AND U13509 ( .A(n267), .B(n13585), .Z(n13584) );
  XNOR U13510 ( .A(n13586), .B(n13583), .Z(n13585) );
  XOR U13511 ( .A(n13587), .B(n13588), .Z(n13560) );
  AND U13512 ( .A(n13589), .B(n13590), .Z(n13588) );
  XNOR U13513 ( .A(n13587), .B(n13576), .Z(n13590) );
  IV U13514 ( .A(n13521), .Z(n13576) );
  XNOR U13515 ( .A(n13591), .B(n13569), .Z(n13521) );
  XNOR U13516 ( .A(n13592), .B(n13575), .Z(n13569) );
  XNOR U13517 ( .A(n13593), .B(n13594), .Z(n13575) );
  NOR U13518 ( .A(n13595), .B(n13596), .Z(n13594) );
  XOR U13519 ( .A(n13593), .B(n13597), .Z(n13595) );
  XNOR U13520 ( .A(n13574), .B(n13566), .Z(n13592) );
  XOR U13521 ( .A(n13598), .B(n13599), .Z(n13566) );
  AND U13522 ( .A(n13600), .B(n13601), .Z(n13599) );
  XOR U13523 ( .A(n13598), .B(n13602), .Z(n13600) );
  XNOR U13524 ( .A(n13603), .B(n13571), .Z(n13574) );
  XOR U13525 ( .A(n13604), .B(n13605), .Z(n13571) );
  AND U13526 ( .A(n13606), .B(n13607), .Z(n13605) );
  XNOR U13527 ( .A(n13608), .B(n13609), .Z(n13606) );
  IV U13528 ( .A(n13604), .Z(n13608) );
  XNOR U13529 ( .A(n13610), .B(n13611), .Z(n13603) );
  NOR U13530 ( .A(n13612), .B(n13613), .Z(n13611) );
  XNOR U13531 ( .A(n13610), .B(n13614), .Z(n13612) );
  XNOR U13532 ( .A(n13570), .B(n13577), .Z(n13591) );
  NOR U13533 ( .A(n13534), .B(n13615), .Z(n13577) );
  XOR U13534 ( .A(n13582), .B(n13581), .Z(n13570) );
  XNOR U13535 ( .A(n13616), .B(n13578), .Z(n13581) );
  XOR U13536 ( .A(n13617), .B(n13618), .Z(n13578) );
  AND U13537 ( .A(n13619), .B(n13620), .Z(n13618) );
  XNOR U13538 ( .A(n13621), .B(n13622), .Z(n13619) );
  IV U13539 ( .A(n13617), .Z(n13621) );
  XNOR U13540 ( .A(n13623), .B(n13624), .Z(n13616) );
  NOR U13541 ( .A(n13625), .B(n13626), .Z(n13624) );
  XNOR U13542 ( .A(n13623), .B(n13627), .Z(n13625) );
  XOR U13543 ( .A(n13628), .B(n13629), .Z(n13582) );
  NOR U13544 ( .A(n13630), .B(n13631), .Z(n13629) );
  XNOR U13545 ( .A(n13628), .B(n13632), .Z(n13630) );
  XNOR U13546 ( .A(n13518), .B(n13587), .Z(n13589) );
  XOR U13547 ( .A(n13633), .B(n13634), .Z(n13518) );
  AND U13548 ( .A(n267), .B(n13635), .Z(n13634) );
  XOR U13549 ( .A(n13636), .B(n13633), .Z(n13635) );
  AND U13550 ( .A(n13531), .B(n13534), .Z(n13587) );
  XOR U13551 ( .A(n13637), .B(n13615), .Z(n13534) );
  XNOR U13552 ( .A(p_input[1040]), .B(p_input[2048]), .Z(n13615) );
  XNOR U13553 ( .A(n13602), .B(n13601), .Z(n13637) );
  XNOR U13554 ( .A(n13638), .B(n13609), .Z(n13601) );
  XNOR U13555 ( .A(n13597), .B(n13596), .Z(n13609) );
  XNOR U13556 ( .A(n13639), .B(n13593), .Z(n13596) );
  XNOR U13557 ( .A(p_input[1050]), .B(p_input[2058]), .Z(n13593) );
  XOR U13558 ( .A(p_input[1051]), .B(n6319), .Z(n13639) );
  XOR U13559 ( .A(p_input[1052]), .B(p_input[2060]), .Z(n13597) );
  XOR U13560 ( .A(n13607), .B(n13640), .Z(n13638) );
  IV U13561 ( .A(n13598), .Z(n13640) );
  XOR U13562 ( .A(p_input[1041]), .B(p_input[2049]), .Z(n13598) );
  XNOR U13563 ( .A(n13641), .B(n13614), .Z(n13607) );
  XNOR U13564 ( .A(p_input[1055]), .B(n6322), .Z(n13614) );
  XOR U13565 ( .A(n13604), .B(n13613), .Z(n13641) );
  XOR U13566 ( .A(n13642), .B(n13610), .Z(n13613) );
  XOR U13567 ( .A(p_input[1053]), .B(p_input[2061]), .Z(n13610) );
  XOR U13568 ( .A(p_input[1054]), .B(n6324), .Z(n13642) );
  XOR U13569 ( .A(p_input[1049]), .B(p_input[2057]), .Z(n13604) );
  XOR U13570 ( .A(n13622), .B(n13620), .Z(n13602) );
  XNOR U13571 ( .A(n13643), .B(n13627), .Z(n13620) );
  XOR U13572 ( .A(p_input[1048]), .B(p_input[2056]), .Z(n13627) );
  XOR U13573 ( .A(n13617), .B(n13626), .Z(n13643) );
  XOR U13574 ( .A(n13644), .B(n13623), .Z(n13626) );
  XOR U13575 ( .A(p_input[1046]), .B(p_input[2054]), .Z(n13623) );
  XOR U13576 ( .A(p_input[1047]), .B(n7007), .Z(n13644) );
  XOR U13577 ( .A(p_input[1042]), .B(p_input[2050]), .Z(n13617) );
  XNOR U13578 ( .A(n13632), .B(n13631), .Z(n13622) );
  XOR U13579 ( .A(n13645), .B(n13628), .Z(n13631) );
  XOR U13580 ( .A(p_input[1043]), .B(p_input[2051]), .Z(n13628) );
  XOR U13581 ( .A(p_input[1044]), .B(n7009), .Z(n13645) );
  XOR U13582 ( .A(p_input[1045]), .B(p_input[2053]), .Z(n13632) );
  XOR U13583 ( .A(n13646), .B(n13647), .Z(n13531) );
  AND U13584 ( .A(n267), .B(n13648), .Z(n13647) );
  XNOR U13585 ( .A(n13649), .B(n13646), .Z(n13648) );
  XNOR U13586 ( .A(n13650), .B(n13651), .Z(n267) );
  AND U13587 ( .A(n13652), .B(n13653), .Z(n13651) );
  XOR U13588 ( .A(n13544), .B(n13650), .Z(n13653) );
  AND U13589 ( .A(n13654), .B(n13655), .Z(n13544) );
  XNOR U13590 ( .A(n13541), .B(n13650), .Z(n13652) );
  XOR U13591 ( .A(n13656), .B(n13657), .Z(n13541) );
  AND U13592 ( .A(n271), .B(n13658), .Z(n13657) );
  XOR U13593 ( .A(n13659), .B(n13656), .Z(n13658) );
  XOR U13594 ( .A(n13660), .B(n13661), .Z(n13650) );
  AND U13595 ( .A(n13662), .B(n13663), .Z(n13661) );
  XNOR U13596 ( .A(n13660), .B(n13654), .Z(n13663) );
  IV U13597 ( .A(n13559), .Z(n13654) );
  XOR U13598 ( .A(n13664), .B(n13665), .Z(n13559) );
  XOR U13599 ( .A(n13666), .B(n13655), .Z(n13665) );
  AND U13600 ( .A(n13586), .B(n13667), .Z(n13655) );
  AND U13601 ( .A(n13668), .B(n13669), .Z(n13666) );
  XOR U13602 ( .A(n13670), .B(n13664), .Z(n13668) );
  XNOR U13603 ( .A(n13556), .B(n13660), .Z(n13662) );
  XOR U13604 ( .A(n13671), .B(n13672), .Z(n13556) );
  AND U13605 ( .A(n271), .B(n13673), .Z(n13672) );
  XOR U13606 ( .A(n13674), .B(n13671), .Z(n13673) );
  XOR U13607 ( .A(n13675), .B(n13676), .Z(n13660) );
  AND U13608 ( .A(n13677), .B(n13678), .Z(n13676) );
  XNOR U13609 ( .A(n13675), .B(n13586), .Z(n13678) );
  XOR U13610 ( .A(n13679), .B(n13669), .Z(n13586) );
  XNOR U13611 ( .A(n13680), .B(n13664), .Z(n13669) );
  XOR U13612 ( .A(n13681), .B(n13682), .Z(n13664) );
  AND U13613 ( .A(n13683), .B(n13684), .Z(n13682) );
  XOR U13614 ( .A(n13685), .B(n13681), .Z(n13683) );
  XNOR U13615 ( .A(n13686), .B(n13687), .Z(n13680) );
  AND U13616 ( .A(n13688), .B(n13689), .Z(n13687) );
  XOR U13617 ( .A(n13686), .B(n13690), .Z(n13688) );
  XNOR U13618 ( .A(n13670), .B(n13667), .Z(n13679) );
  AND U13619 ( .A(n13691), .B(n13692), .Z(n13667) );
  XOR U13620 ( .A(n13693), .B(n13694), .Z(n13670) );
  AND U13621 ( .A(n13695), .B(n13696), .Z(n13694) );
  XOR U13622 ( .A(n13693), .B(n13697), .Z(n13695) );
  XNOR U13623 ( .A(n13583), .B(n13675), .Z(n13677) );
  XOR U13624 ( .A(n13698), .B(n13699), .Z(n13583) );
  AND U13625 ( .A(n271), .B(n13700), .Z(n13699) );
  XNOR U13626 ( .A(n13701), .B(n13698), .Z(n13700) );
  XOR U13627 ( .A(n13702), .B(n13703), .Z(n13675) );
  AND U13628 ( .A(n13704), .B(n13705), .Z(n13703) );
  XNOR U13629 ( .A(n13702), .B(n13691), .Z(n13705) );
  IV U13630 ( .A(n13636), .Z(n13691) );
  XNOR U13631 ( .A(n13706), .B(n13684), .Z(n13636) );
  XNOR U13632 ( .A(n13707), .B(n13690), .Z(n13684) );
  XNOR U13633 ( .A(n13708), .B(n13709), .Z(n13690) );
  NOR U13634 ( .A(n13710), .B(n13711), .Z(n13709) );
  XOR U13635 ( .A(n13708), .B(n13712), .Z(n13710) );
  XNOR U13636 ( .A(n13689), .B(n13681), .Z(n13707) );
  XOR U13637 ( .A(n13713), .B(n13714), .Z(n13681) );
  AND U13638 ( .A(n13715), .B(n13716), .Z(n13714) );
  XOR U13639 ( .A(n13713), .B(n13717), .Z(n13715) );
  XNOR U13640 ( .A(n13718), .B(n13686), .Z(n13689) );
  XOR U13641 ( .A(n13719), .B(n13720), .Z(n13686) );
  AND U13642 ( .A(n13721), .B(n13722), .Z(n13720) );
  XNOR U13643 ( .A(n13723), .B(n13724), .Z(n13721) );
  IV U13644 ( .A(n13719), .Z(n13723) );
  XNOR U13645 ( .A(n13725), .B(n13726), .Z(n13718) );
  NOR U13646 ( .A(n13727), .B(n13728), .Z(n13726) );
  XNOR U13647 ( .A(n13725), .B(n13729), .Z(n13727) );
  XNOR U13648 ( .A(n13685), .B(n13692), .Z(n13706) );
  NOR U13649 ( .A(n13649), .B(n13730), .Z(n13692) );
  XOR U13650 ( .A(n13697), .B(n13696), .Z(n13685) );
  XNOR U13651 ( .A(n13731), .B(n13693), .Z(n13696) );
  XOR U13652 ( .A(n13732), .B(n13733), .Z(n13693) );
  AND U13653 ( .A(n13734), .B(n13735), .Z(n13733) );
  XNOR U13654 ( .A(n13736), .B(n13737), .Z(n13734) );
  IV U13655 ( .A(n13732), .Z(n13736) );
  XNOR U13656 ( .A(n13738), .B(n13739), .Z(n13731) );
  NOR U13657 ( .A(n13740), .B(n13741), .Z(n13739) );
  XNOR U13658 ( .A(n13738), .B(n13742), .Z(n13740) );
  XOR U13659 ( .A(n13743), .B(n13744), .Z(n13697) );
  NOR U13660 ( .A(n13745), .B(n13746), .Z(n13744) );
  XNOR U13661 ( .A(n13743), .B(n13747), .Z(n13745) );
  XNOR U13662 ( .A(n13633), .B(n13702), .Z(n13704) );
  XOR U13663 ( .A(n13748), .B(n13749), .Z(n13633) );
  AND U13664 ( .A(n271), .B(n13750), .Z(n13749) );
  XOR U13665 ( .A(n13751), .B(n13748), .Z(n13750) );
  AND U13666 ( .A(n13646), .B(n13649), .Z(n13702) );
  XOR U13667 ( .A(n13752), .B(n13730), .Z(n13649) );
  XNOR U13668 ( .A(p_input[1056]), .B(p_input[2048]), .Z(n13730) );
  XNOR U13669 ( .A(n13717), .B(n13716), .Z(n13752) );
  XNOR U13670 ( .A(n13753), .B(n13724), .Z(n13716) );
  XNOR U13671 ( .A(n13712), .B(n13711), .Z(n13724) );
  XNOR U13672 ( .A(n13754), .B(n13708), .Z(n13711) );
  XNOR U13673 ( .A(p_input[1066]), .B(p_input[2058]), .Z(n13708) );
  XOR U13674 ( .A(p_input[1067]), .B(n6319), .Z(n13754) );
  XOR U13675 ( .A(p_input[1068]), .B(p_input[2060]), .Z(n13712) );
  XOR U13676 ( .A(n13722), .B(n13755), .Z(n13753) );
  IV U13677 ( .A(n13713), .Z(n13755) );
  XOR U13678 ( .A(p_input[1057]), .B(p_input[2049]), .Z(n13713) );
  XNOR U13679 ( .A(n13756), .B(n13729), .Z(n13722) );
  XNOR U13680 ( .A(p_input[1071]), .B(n6322), .Z(n13729) );
  XOR U13681 ( .A(n13719), .B(n13728), .Z(n13756) );
  XOR U13682 ( .A(n13757), .B(n13725), .Z(n13728) );
  XOR U13683 ( .A(p_input[1069]), .B(p_input[2061]), .Z(n13725) );
  XOR U13684 ( .A(p_input[1070]), .B(n6324), .Z(n13757) );
  XOR U13685 ( .A(p_input[1065]), .B(p_input[2057]), .Z(n13719) );
  XOR U13686 ( .A(n13737), .B(n13735), .Z(n13717) );
  XNOR U13687 ( .A(n13758), .B(n13742), .Z(n13735) );
  XOR U13688 ( .A(p_input[1064]), .B(p_input[2056]), .Z(n13742) );
  XOR U13689 ( .A(n13732), .B(n13741), .Z(n13758) );
  XOR U13690 ( .A(n13759), .B(n13738), .Z(n13741) );
  XOR U13691 ( .A(p_input[1062]), .B(p_input[2054]), .Z(n13738) );
  XOR U13692 ( .A(p_input[1063]), .B(n7007), .Z(n13759) );
  XOR U13693 ( .A(p_input[1058]), .B(p_input[2050]), .Z(n13732) );
  XNOR U13694 ( .A(n13747), .B(n13746), .Z(n13737) );
  XOR U13695 ( .A(n13760), .B(n13743), .Z(n13746) );
  XOR U13696 ( .A(p_input[1059]), .B(p_input[2051]), .Z(n13743) );
  XOR U13697 ( .A(p_input[1060]), .B(n7009), .Z(n13760) );
  XOR U13698 ( .A(p_input[1061]), .B(p_input[2053]), .Z(n13747) );
  XOR U13699 ( .A(n13761), .B(n13762), .Z(n13646) );
  AND U13700 ( .A(n271), .B(n13763), .Z(n13762) );
  XNOR U13701 ( .A(n13764), .B(n13761), .Z(n13763) );
  XNOR U13702 ( .A(n13765), .B(n13766), .Z(n271) );
  AND U13703 ( .A(n13767), .B(n13768), .Z(n13766) );
  XOR U13704 ( .A(n13659), .B(n13765), .Z(n13768) );
  AND U13705 ( .A(n13769), .B(n13770), .Z(n13659) );
  XNOR U13706 ( .A(n13656), .B(n13765), .Z(n13767) );
  XOR U13707 ( .A(n13771), .B(n13772), .Z(n13656) );
  AND U13708 ( .A(n275), .B(n13773), .Z(n13772) );
  XOR U13709 ( .A(n13774), .B(n13771), .Z(n13773) );
  XOR U13710 ( .A(n13775), .B(n13776), .Z(n13765) );
  AND U13711 ( .A(n13777), .B(n13778), .Z(n13776) );
  XNOR U13712 ( .A(n13775), .B(n13769), .Z(n13778) );
  IV U13713 ( .A(n13674), .Z(n13769) );
  XOR U13714 ( .A(n13779), .B(n13780), .Z(n13674) );
  XOR U13715 ( .A(n13781), .B(n13770), .Z(n13780) );
  AND U13716 ( .A(n13701), .B(n13782), .Z(n13770) );
  AND U13717 ( .A(n13783), .B(n13784), .Z(n13781) );
  XOR U13718 ( .A(n13785), .B(n13779), .Z(n13783) );
  XNOR U13719 ( .A(n13671), .B(n13775), .Z(n13777) );
  XOR U13720 ( .A(n13786), .B(n13787), .Z(n13671) );
  AND U13721 ( .A(n275), .B(n13788), .Z(n13787) );
  XOR U13722 ( .A(n13789), .B(n13786), .Z(n13788) );
  XOR U13723 ( .A(n13790), .B(n13791), .Z(n13775) );
  AND U13724 ( .A(n13792), .B(n13793), .Z(n13791) );
  XNOR U13725 ( .A(n13790), .B(n13701), .Z(n13793) );
  XOR U13726 ( .A(n13794), .B(n13784), .Z(n13701) );
  XNOR U13727 ( .A(n13795), .B(n13779), .Z(n13784) );
  XOR U13728 ( .A(n13796), .B(n13797), .Z(n13779) );
  AND U13729 ( .A(n13798), .B(n13799), .Z(n13797) );
  XOR U13730 ( .A(n13800), .B(n13796), .Z(n13798) );
  XNOR U13731 ( .A(n13801), .B(n13802), .Z(n13795) );
  AND U13732 ( .A(n13803), .B(n13804), .Z(n13802) );
  XOR U13733 ( .A(n13801), .B(n13805), .Z(n13803) );
  XNOR U13734 ( .A(n13785), .B(n13782), .Z(n13794) );
  AND U13735 ( .A(n13806), .B(n13807), .Z(n13782) );
  XOR U13736 ( .A(n13808), .B(n13809), .Z(n13785) );
  AND U13737 ( .A(n13810), .B(n13811), .Z(n13809) );
  XOR U13738 ( .A(n13808), .B(n13812), .Z(n13810) );
  XNOR U13739 ( .A(n13698), .B(n13790), .Z(n13792) );
  XOR U13740 ( .A(n13813), .B(n13814), .Z(n13698) );
  AND U13741 ( .A(n275), .B(n13815), .Z(n13814) );
  XNOR U13742 ( .A(n13816), .B(n13813), .Z(n13815) );
  XOR U13743 ( .A(n13817), .B(n13818), .Z(n13790) );
  AND U13744 ( .A(n13819), .B(n13820), .Z(n13818) );
  XNOR U13745 ( .A(n13817), .B(n13806), .Z(n13820) );
  IV U13746 ( .A(n13751), .Z(n13806) );
  XNOR U13747 ( .A(n13821), .B(n13799), .Z(n13751) );
  XNOR U13748 ( .A(n13822), .B(n13805), .Z(n13799) );
  XNOR U13749 ( .A(n13823), .B(n13824), .Z(n13805) );
  NOR U13750 ( .A(n13825), .B(n13826), .Z(n13824) );
  XOR U13751 ( .A(n13823), .B(n13827), .Z(n13825) );
  XNOR U13752 ( .A(n13804), .B(n13796), .Z(n13822) );
  XOR U13753 ( .A(n13828), .B(n13829), .Z(n13796) );
  AND U13754 ( .A(n13830), .B(n13831), .Z(n13829) );
  XOR U13755 ( .A(n13828), .B(n13832), .Z(n13830) );
  XNOR U13756 ( .A(n13833), .B(n13801), .Z(n13804) );
  XOR U13757 ( .A(n13834), .B(n13835), .Z(n13801) );
  AND U13758 ( .A(n13836), .B(n13837), .Z(n13835) );
  XNOR U13759 ( .A(n13838), .B(n13839), .Z(n13836) );
  IV U13760 ( .A(n13834), .Z(n13838) );
  XNOR U13761 ( .A(n13840), .B(n13841), .Z(n13833) );
  NOR U13762 ( .A(n13842), .B(n13843), .Z(n13841) );
  XNOR U13763 ( .A(n13840), .B(n13844), .Z(n13842) );
  XNOR U13764 ( .A(n13800), .B(n13807), .Z(n13821) );
  NOR U13765 ( .A(n13764), .B(n13845), .Z(n13807) );
  XOR U13766 ( .A(n13812), .B(n13811), .Z(n13800) );
  XNOR U13767 ( .A(n13846), .B(n13808), .Z(n13811) );
  XOR U13768 ( .A(n13847), .B(n13848), .Z(n13808) );
  AND U13769 ( .A(n13849), .B(n13850), .Z(n13848) );
  XNOR U13770 ( .A(n13851), .B(n13852), .Z(n13849) );
  IV U13771 ( .A(n13847), .Z(n13851) );
  XNOR U13772 ( .A(n13853), .B(n13854), .Z(n13846) );
  NOR U13773 ( .A(n13855), .B(n13856), .Z(n13854) );
  XNOR U13774 ( .A(n13853), .B(n13857), .Z(n13855) );
  XOR U13775 ( .A(n13858), .B(n13859), .Z(n13812) );
  NOR U13776 ( .A(n13860), .B(n13861), .Z(n13859) );
  XNOR U13777 ( .A(n13858), .B(n13862), .Z(n13860) );
  XNOR U13778 ( .A(n13748), .B(n13817), .Z(n13819) );
  XOR U13779 ( .A(n13863), .B(n13864), .Z(n13748) );
  AND U13780 ( .A(n275), .B(n13865), .Z(n13864) );
  XOR U13781 ( .A(n13866), .B(n13863), .Z(n13865) );
  AND U13782 ( .A(n13761), .B(n13764), .Z(n13817) );
  XOR U13783 ( .A(n13867), .B(n13845), .Z(n13764) );
  XNOR U13784 ( .A(p_input[1072]), .B(p_input[2048]), .Z(n13845) );
  XNOR U13785 ( .A(n13832), .B(n13831), .Z(n13867) );
  XNOR U13786 ( .A(n13868), .B(n13839), .Z(n13831) );
  XNOR U13787 ( .A(n13827), .B(n13826), .Z(n13839) );
  XNOR U13788 ( .A(n13869), .B(n13823), .Z(n13826) );
  XNOR U13789 ( .A(p_input[1082]), .B(p_input[2058]), .Z(n13823) );
  XOR U13790 ( .A(p_input[1083]), .B(n6319), .Z(n13869) );
  XOR U13791 ( .A(p_input[1084]), .B(p_input[2060]), .Z(n13827) );
  XOR U13792 ( .A(n13837), .B(n13870), .Z(n13868) );
  IV U13793 ( .A(n13828), .Z(n13870) );
  XOR U13794 ( .A(p_input[1073]), .B(p_input[2049]), .Z(n13828) );
  XNOR U13795 ( .A(n13871), .B(n13844), .Z(n13837) );
  XNOR U13796 ( .A(p_input[1087]), .B(n6322), .Z(n13844) );
  XOR U13797 ( .A(n13834), .B(n13843), .Z(n13871) );
  XOR U13798 ( .A(n13872), .B(n13840), .Z(n13843) );
  XOR U13799 ( .A(p_input[1085]), .B(p_input[2061]), .Z(n13840) );
  XOR U13800 ( .A(p_input[1086]), .B(n6324), .Z(n13872) );
  XOR U13801 ( .A(p_input[1081]), .B(p_input[2057]), .Z(n13834) );
  XOR U13802 ( .A(n13852), .B(n13850), .Z(n13832) );
  XNOR U13803 ( .A(n13873), .B(n13857), .Z(n13850) );
  XOR U13804 ( .A(p_input[1080]), .B(p_input[2056]), .Z(n13857) );
  XOR U13805 ( .A(n13847), .B(n13856), .Z(n13873) );
  XOR U13806 ( .A(n13874), .B(n13853), .Z(n13856) );
  XOR U13807 ( .A(p_input[1078]), .B(p_input[2054]), .Z(n13853) );
  XOR U13808 ( .A(p_input[1079]), .B(n7007), .Z(n13874) );
  XOR U13809 ( .A(p_input[1074]), .B(p_input[2050]), .Z(n13847) );
  XNOR U13810 ( .A(n13862), .B(n13861), .Z(n13852) );
  XOR U13811 ( .A(n13875), .B(n13858), .Z(n13861) );
  XOR U13812 ( .A(p_input[1075]), .B(p_input[2051]), .Z(n13858) );
  XOR U13813 ( .A(p_input[1076]), .B(n7009), .Z(n13875) );
  XOR U13814 ( .A(p_input[1077]), .B(p_input[2053]), .Z(n13862) );
  XOR U13815 ( .A(n13876), .B(n13877), .Z(n13761) );
  AND U13816 ( .A(n275), .B(n13878), .Z(n13877) );
  XNOR U13817 ( .A(n13879), .B(n13876), .Z(n13878) );
  XNOR U13818 ( .A(n13880), .B(n13881), .Z(n275) );
  AND U13819 ( .A(n13882), .B(n13883), .Z(n13881) );
  XOR U13820 ( .A(n13774), .B(n13880), .Z(n13883) );
  AND U13821 ( .A(n13884), .B(n13885), .Z(n13774) );
  XNOR U13822 ( .A(n13771), .B(n13880), .Z(n13882) );
  XOR U13823 ( .A(n13886), .B(n13887), .Z(n13771) );
  AND U13824 ( .A(n279), .B(n13888), .Z(n13887) );
  XOR U13825 ( .A(n13889), .B(n13886), .Z(n13888) );
  XOR U13826 ( .A(n13890), .B(n13891), .Z(n13880) );
  AND U13827 ( .A(n13892), .B(n13893), .Z(n13891) );
  XNOR U13828 ( .A(n13890), .B(n13884), .Z(n13893) );
  IV U13829 ( .A(n13789), .Z(n13884) );
  XOR U13830 ( .A(n13894), .B(n13895), .Z(n13789) );
  XOR U13831 ( .A(n13896), .B(n13885), .Z(n13895) );
  AND U13832 ( .A(n13816), .B(n13897), .Z(n13885) );
  AND U13833 ( .A(n13898), .B(n13899), .Z(n13896) );
  XOR U13834 ( .A(n13900), .B(n13894), .Z(n13898) );
  XNOR U13835 ( .A(n13786), .B(n13890), .Z(n13892) );
  XOR U13836 ( .A(n13901), .B(n13902), .Z(n13786) );
  AND U13837 ( .A(n279), .B(n13903), .Z(n13902) );
  XOR U13838 ( .A(n13904), .B(n13901), .Z(n13903) );
  XOR U13839 ( .A(n13905), .B(n13906), .Z(n13890) );
  AND U13840 ( .A(n13907), .B(n13908), .Z(n13906) );
  XNOR U13841 ( .A(n13905), .B(n13816), .Z(n13908) );
  XOR U13842 ( .A(n13909), .B(n13899), .Z(n13816) );
  XNOR U13843 ( .A(n13910), .B(n13894), .Z(n13899) );
  XOR U13844 ( .A(n13911), .B(n13912), .Z(n13894) );
  AND U13845 ( .A(n13913), .B(n13914), .Z(n13912) );
  XOR U13846 ( .A(n13915), .B(n13911), .Z(n13913) );
  XNOR U13847 ( .A(n13916), .B(n13917), .Z(n13910) );
  AND U13848 ( .A(n13918), .B(n13919), .Z(n13917) );
  XOR U13849 ( .A(n13916), .B(n13920), .Z(n13918) );
  XNOR U13850 ( .A(n13900), .B(n13897), .Z(n13909) );
  AND U13851 ( .A(n13921), .B(n13922), .Z(n13897) );
  XOR U13852 ( .A(n13923), .B(n13924), .Z(n13900) );
  AND U13853 ( .A(n13925), .B(n13926), .Z(n13924) );
  XOR U13854 ( .A(n13923), .B(n13927), .Z(n13925) );
  XNOR U13855 ( .A(n13813), .B(n13905), .Z(n13907) );
  XOR U13856 ( .A(n13928), .B(n13929), .Z(n13813) );
  AND U13857 ( .A(n279), .B(n13930), .Z(n13929) );
  XNOR U13858 ( .A(n13931), .B(n13928), .Z(n13930) );
  XOR U13859 ( .A(n13932), .B(n13933), .Z(n13905) );
  AND U13860 ( .A(n13934), .B(n13935), .Z(n13933) );
  XNOR U13861 ( .A(n13932), .B(n13921), .Z(n13935) );
  IV U13862 ( .A(n13866), .Z(n13921) );
  XNOR U13863 ( .A(n13936), .B(n13914), .Z(n13866) );
  XNOR U13864 ( .A(n13937), .B(n13920), .Z(n13914) );
  XNOR U13865 ( .A(n13938), .B(n13939), .Z(n13920) );
  NOR U13866 ( .A(n13940), .B(n13941), .Z(n13939) );
  XOR U13867 ( .A(n13938), .B(n13942), .Z(n13940) );
  XNOR U13868 ( .A(n13919), .B(n13911), .Z(n13937) );
  XOR U13869 ( .A(n13943), .B(n13944), .Z(n13911) );
  AND U13870 ( .A(n13945), .B(n13946), .Z(n13944) );
  XOR U13871 ( .A(n13943), .B(n13947), .Z(n13945) );
  XNOR U13872 ( .A(n13948), .B(n13916), .Z(n13919) );
  XOR U13873 ( .A(n13949), .B(n13950), .Z(n13916) );
  AND U13874 ( .A(n13951), .B(n13952), .Z(n13950) );
  XNOR U13875 ( .A(n13953), .B(n13954), .Z(n13951) );
  IV U13876 ( .A(n13949), .Z(n13953) );
  XNOR U13877 ( .A(n13955), .B(n13956), .Z(n13948) );
  NOR U13878 ( .A(n13957), .B(n13958), .Z(n13956) );
  XNOR U13879 ( .A(n13955), .B(n13959), .Z(n13957) );
  XNOR U13880 ( .A(n13915), .B(n13922), .Z(n13936) );
  NOR U13881 ( .A(n13879), .B(n13960), .Z(n13922) );
  XOR U13882 ( .A(n13927), .B(n13926), .Z(n13915) );
  XNOR U13883 ( .A(n13961), .B(n13923), .Z(n13926) );
  XOR U13884 ( .A(n13962), .B(n13963), .Z(n13923) );
  AND U13885 ( .A(n13964), .B(n13965), .Z(n13963) );
  XNOR U13886 ( .A(n13966), .B(n13967), .Z(n13964) );
  IV U13887 ( .A(n13962), .Z(n13966) );
  XNOR U13888 ( .A(n13968), .B(n13969), .Z(n13961) );
  NOR U13889 ( .A(n13970), .B(n13971), .Z(n13969) );
  XNOR U13890 ( .A(n13968), .B(n13972), .Z(n13970) );
  XOR U13891 ( .A(n13973), .B(n13974), .Z(n13927) );
  NOR U13892 ( .A(n13975), .B(n13976), .Z(n13974) );
  XNOR U13893 ( .A(n13973), .B(n13977), .Z(n13975) );
  XNOR U13894 ( .A(n13863), .B(n13932), .Z(n13934) );
  XOR U13895 ( .A(n13978), .B(n13979), .Z(n13863) );
  AND U13896 ( .A(n279), .B(n13980), .Z(n13979) );
  XOR U13897 ( .A(n13981), .B(n13978), .Z(n13980) );
  AND U13898 ( .A(n13876), .B(n13879), .Z(n13932) );
  XOR U13899 ( .A(n13982), .B(n13960), .Z(n13879) );
  XNOR U13900 ( .A(p_input[1088]), .B(p_input[2048]), .Z(n13960) );
  XNOR U13901 ( .A(n13947), .B(n13946), .Z(n13982) );
  XNOR U13902 ( .A(n13983), .B(n13954), .Z(n13946) );
  XNOR U13903 ( .A(n13942), .B(n13941), .Z(n13954) );
  XNOR U13904 ( .A(n13984), .B(n13938), .Z(n13941) );
  XNOR U13905 ( .A(p_input[1098]), .B(p_input[2058]), .Z(n13938) );
  XOR U13906 ( .A(p_input[1099]), .B(n6319), .Z(n13984) );
  XOR U13907 ( .A(p_input[1100]), .B(p_input[2060]), .Z(n13942) );
  XOR U13908 ( .A(n13952), .B(n13985), .Z(n13983) );
  IV U13909 ( .A(n13943), .Z(n13985) );
  XOR U13910 ( .A(p_input[1089]), .B(p_input[2049]), .Z(n13943) );
  XNOR U13911 ( .A(n13986), .B(n13959), .Z(n13952) );
  XNOR U13912 ( .A(p_input[1103]), .B(n6322), .Z(n13959) );
  XOR U13913 ( .A(n13949), .B(n13958), .Z(n13986) );
  XOR U13914 ( .A(n13987), .B(n13955), .Z(n13958) );
  XOR U13915 ( .A(p_input[1101]), .B(p_input[2061]), .Z(n13955) );
  XOR U13916 ( .A(p_input[1102]), .B(n6324), .Z(n13987) );
  XOR U13917 ( .A(p_input[1097]), .B(p_input[2057]), .Z(n13949) );
  XOR U13918 ( .A(n13967), .B(n13965), .Z(n13947) );
  XNOR U13919 ( .A(n13988), .B(n13972), .Z(n13965) );
  XOR U13920 ( .A(p_input[1096]), .B(p_input[2056]), .Z(n13972) );
  XOR U13921 ( .A(n13962), .B(n13971), .Z(n13988) );
  XOR U13922 ( .A(n13989), .B(n13968), .Z(n13971) );
  XOR U13923 ( .A(p_input[1094]), .B(p_input[2054]), .Z(n13968) );
  XOR U13924 ( .A(p_input[1095]), .B(n7007), .Z(n13989) );
  XOR U13925 ( .A(p_input[1090]), .B(p_input[2050]), .Z(n13962) );
  XNOR U13926 ( .A(n13977), .B(n13976), .Z(n13967) );
  XOR U13927 ( .A(n13990), .B(n13973), .Z(n13976) );
  XOR U13928 ( .A(p_input[1091]), .B(p_input[2051]), .Z(n13973) );
  XOR U13929 ( .A(p_input[1092]), .B(n7009), .Z(n13990) );
  XOR U13930 ( .A(p_input[1093]), .B(p_input[2053]), .Z(n13977) );
  XOR U13931 ( .A(n13991), .B(n13992), .Z(n13876) );
  AND U13932 ( .A(n279), .B(n13993), .Z(n13992) );
  XNOR U13933 ( .A(n13994), .B(n13991), .Z(n13993) );
  XNOR U13934 ( .A(n13995), .B(n13996), .Z(n279) );
  AND U13935 ( .A(n13997), .B(n13998), .Z(n13996) );
  XOR U13936 ( .A(n13889), .B(n13995), .Z(n13998) );
  AND U13937 ( .A(n13999), .B(n14000), .Z(n13889) );
  XNOR U13938 ( .A(n13886), .B(n13995), .Z(n13997) );
  XOR U13939 ( .A(n14001), .B(n14002), .Z(n13886) );
  AND U13940 ( .A(n283), .B(n14003), .Z(n14002) );
  XOR U13941 ( .A(n14004), .B(n14001), .Z(n14003) );
  XOR U13942 ( .A(n14005), .B(n14006), .Z(n13995) );
  AND U13943 ( .A(n14007), .B(n14008), .Z(n14006) );
  XNOR U13944 ( .A(n14005), .B(n13999), .Z(n14008) );
  IV U13945 ( .A(n13904), .Z(n13999) );
  XOR U13946 ( .A(n14009), .B(n14010), .Z(n13904) );
  XOR U13947 ( .A(n14011), .B(n14000), .Z(n14010) );
  AND U13948 ( .A(n13931), .B(n14012), .Z(n14000) );
  AND U13949 ( .A(n14013), .B(n14014), .Z(n14011) );
  XOR U13950 ( .A(n14015), .B(n14009), .Z(n14013) );
  XNOR U13951 ( .A(n13901), .B(n14005), .Z(n14007) );
  XOR U13952 ( .A(n14016), .B(n14017), .Z(n13901) );
  AND U13953 ( .A(n283), .B(n14018), .Z(n14017) );
  XOR U13954 ( .A(n14019), .B(n14016), .Z(n14018) );
  XOR U13955 ( .A(n14020), .B(n14021), .Z(n14005) );
  AND U13956 ( .A(n14022), .B(n14023), .Z(n14021) );
  XNOR U13957 ( .A(n14020), .B(n13931), .Z(n14023) );
  XOR U13958 ( .A(n14024), .B(n14014), .Z(n13931) );
  XNOR U13959 ( .A(n14025), .B(n14009), .Z(n14014) );
  XOR U13960 ( .A(n14026), .B(n14027), .Z(n14009) );
  AND U13961 ( .A(n14028), .B(n14029), .Z(n14027) );
  XOR U13962 ( .A(n14030), .B(n14026), .Z(n14028) );
  XNOR U13963 ( .A(n14031), .B(n14032), .Z(n14025) );
  AND U13964 ( .A(n14033), .B(n14034), .Z(n14032) );
  XOR U13965 ( .A(n14031), .B(n14035), .Z(n14033) );
  XNOR U13966 ( .A(n14015), .B(n14012), .Z(n14024) );
  AND U13967 ( .A(n14036), .B(n14037), .Z(n14012) );
  XOR U13968 ( .A(n14038), .B(n14039), .Z(n14015) );
  AND U13969 ( .A(n14040), .B(n14041), .Z(n14039) );
  XOR U13970 ( .A(n14038), .B(n14042), .Z(n14040) );
  XNOR U13971 ( .A(n13928), .B(n14020), .Z(n14022) );
  XOR U13972 ( .A(n14043), .B(n14044), .Z(n13928) );
  AND U13973 ( .A(n283), .B(n14045), .Z(n14044) );
  XNOR U13974 ( .A(n14046), .B(n14043), .Z(n14045) );
  XOR U13975 ( .A(n14047), .B(n14048), .Z(n14020) );
  AND U13976 ( .A(n14049), .B(n14050), .Z(n14048) );
  XNOR U13977 ( .A(n14047), .B(n14036), .Z(n14050) );
  IV U13978 ( .A(n13981), .Z(n14036) );
  XNOR U13979 ( .A(n14051), .B(n14029), .Z(n13981) );
  XNOR U13980 ( .A(n14052), .B(n14035), .Z(n14029) );
  XNOR U13981 ( .A(n14053), .B(n14054), .Z(n14035) );
  NOR U13982 ( .A(n14055), .B(n14056), .Z(n14054) );
  XOR U13983 ( .A(n14053), .B(n14057), .Z(n14055) );
  XNOR U13984 ( .A(n14034), .B(n14026), .Z(n14052) );
  XOR U13985 ( .A(n14058), .B(n14059), .Z(n14026) );
  AND U13986 ( .A(n14060), .B(n14061), .Z(n14059) );
  XOR U13987 ( .A(n14058), .B(n14062), .Z(n14060) );
  XNOR U13988 ( .A(n14063), .B(n14031), .Z(n14034) );
  XOR U13989 ( .A(n14064), .B(n14065), .Z(n14031) );
  AND U13990 ( .A(n14066), .B(n14067), .Z(n14065) );
  XNOR U13991 ( .A(n14068), .B(n14069), .Z(n14066) );
  IV U13992 ( .A(n14064), .Z(n14068) );
  XNOR U13993 ( .A(n14070), .B(n14071), .Z(n14063) );
  NOR U13994 ( .A(n14072), .B(n14073), .Z(n14071) );
  XNOR U13995 ( .A(n14070), .B(n14074), .Z(n14072) );
  XNOR U13996 ( .A(n14030), .B(n14037), .Z(n14051) );
  NOR U13997 ( .A(n13994), .B(n14075), .Z(n14037) );
  XOR U13998 ( .A(n14042), .B(n14041), .Z(n14030) );
  XNOR U13999 ( .A(n14076), .B(n14038), .Z(n14041) );
  XOR U14000 ( .A(n14077), .B(n14078), .Z(n14038) );
  AND U14001 ( .A(n14079), .B(n14080), .Z(n14078) );
  XNOR U14002 ( .A(n14081), .B(n14082), .Z(n14079) );
  IV U14003 ( .A(n14077), .Z(n14081) );
  XNOR U14004 ( .A(n14083), .B(n14084), .Z(n14076) );
  NOR U14005 ( .A(n14085), .B(n14086), .Z(n14084) );
  XNOR U14006 ( .A(n14083), .B(n14087), .Z(n14085) );
  XOR U14007 ( .A(n14088), .B(n14089), .Z(n14042) );
  NOR U14008 ( .A(n14090), .B(n14091), .Z(n14089) );
  XNOR U14009 ( .A(n14088), .B(n14092), .Z(n14090) );
  XNOR U14010 ( .A(n13978), .B(n14047), .Z(n14049) );
  XOR U14011 ( .A(n14093), .B(n14094), .Z(n13978) );
  AND U14012 ( .A(n283), .B(n14095), .Z(n14094) );
  XOR U14013 ( .A(n14096), .B(n14093), .Z(n14095) );
  AND U14014 ( .A(n13991), .B(n13994), .Z(n14047) );
  XOR U14015 ( .A(n14097), .B(n14075), .Z(n13994) );
  XNOR U14016 ( .A(p_input[1104]), .B(p_input[2048]), .Z(n14075) );
  XNOR U14017 ( .A(n14062), .B(n14061), .Z(n14097) );
  XNOR U14018 ( .A(n14098), .B(n14069), .Z(n14061) );
  XNOR U14019 ( .A(n14057), .B(n14056), .Z(n14069) );
  XNOR U14020 ( .A(n14099), .B(n14053), .Z(n14056) );
  XNOR U14021 ( .A(p_input[1114]), .B(p_input[2058]), .Z(n14053) );
  XOR U14022 ( .A(p_input[1115]), .B(n6319), .Z(n14099) );
  XOR U14023 ( .A(p_input[1116]), .B(p_input[2060]), .Z(n14057) );
  XOR U14024 ( .A(n14067), .B(n14100), .Z(n14098) );
  IV U14025 ( .A(n14058), .Z(n14100) );
  XOR U14026 ( .A(p_input[1105]), .B(p_input[2049]), .Z(n14058) );
  XNOR U14027 ( .A(n14101), .B(n14074), .Z(n14067) );
  XNOR U14028 ( .A(p_input[1119]), .B(n6322), .Z(n14074) );
  XOR U14029 ( .A(n14064), .B(n14073), .Z(n14101) );
  XOR U14030 ( .A(n14102), .B(n14070), .Z(n14073) );
  XOR U14031 ( .A(p_input[1117]), .B(p_input[2061]), .Z(n14070) );
  XOR U14032 ( .A(p_input[1118]), .B(n6324), .Z(n14102) );
  XOR U14033 ( .A(p_input[1113]), .B(p_input[2057]), .Z(n14064) );
  XOR U14034 ( .A(n14082), .B(n14080), .Z(n14062) );
  XNOR U14035 ( .A(n14103), .B(n14087), .Z(n14080) );
  XOR U14036 ( .A(p_input[1112]), .B(p_input[2056]), .Z(n14087) );
  XOR U14037 ( .A(n14077), .B(n14086), .Z(n14103) );
  XOR U14038 ( .A(n14104), .B(n14083), .Z(n14086) );
  XOR U14039 ( .A(p_input[1110]), .B(p_input[2054]), .Z(n14083) );
  XOR U14040 ( .A(p_input[1111]), .B(n7007), .Z(n14104) );
  XOR U14041 ( .A(p_input[1106]), .B(p_input[2050]), .Z(n14077) );
  XNOR U14042 ( .A(n14092), .B(n14091), .Z(n14082) );
  XOR U14043 ( .A(n14105), .B(n14088), .Z(n14091) );
  XOR U14044 ( .A(p_input[1107]), .B(p_input[2051]), .Z(n14088) );
  XOR U14045 ( .A(p_input[1108]), .B(n7009), .Z(n14105) );
  XOR U14046 ( .A(p_input[1109]), .B(p_input[2053]), .Z(n14092) );
  XOR U14047 ( .A(n14106), .B(n14107), .Z(n13991) );
  AND U14048 ( .A(n283), .B(n14108), .Z(n14107) );
  XNOR U14049 ( .A(n14109), .B(n14106), .Z(n14108) );
  XNOR U14050 ( .A(n14110), .B(n14111), .Z(n283) );
  AND U14051 ( .A(n14112), .B(n14113), .Z(n14111) );
  XOR U14052 ( .A(n14004), .B(n14110), .Z(n14113) );
  AND U14053 ( .A(n14114), .B(n14115), .Z(n14004) );
  XNOR U14054 ( .A(n14001), .B(n14110), .Z(n14112) );
  XOR U14055 ( .A(n14116), .B(n14117), .Z(n14001) );
  AND U14056 ( .A(n287), .B(n14118), .Z(n14117) );
  XOR U14057 ( .A(n14119), .B(n14116), .Z(n14118) );
  XOR U14058 ( .A(n14120), .B(n14121), .Z(n14110) );
  AND U14059 ( .A(n14122), .B(n14123), .Z(n14121) );
  XNOR U14060 ( .A(n14120), .B(n14114), .Z(n14123) );
  IV U14061 ( .A(n14019), .Z(n14114) );
  XOR U14062 ( .A(n14124), .B(n14125), .Z(n14019) );
  XOR U14063 ( .A(n14126), .B(n14115), .Z(n14125) );
  AND U14064 ( .A(n14046), .B(n14127), .Z(n14115) );
  AND U14065 ( .A(n14128), .B(n14129), .Z(n14126) );
  XOR U14066 ( .A(n14130), .B(n14124), .Z(n14128) );
  XNOR U14067 ( .A(n14016), .B(n14120), .Z(n14122) );
  XOR U14068 ( .A(n14131), .B(n14132), .Z(n14016) );
  AND U14069 ( .A(n287), .B(n14133), .Z(n14132) );
  XOR U14070 ( .A(n14134), .B(n14131), .Z(n14133) );
  XOR U14071 ( .A(n14135), .B(n14136), .Z(n14120) );
  AND U14072 ( .A(n14137), .B(n14138), .Z(n14136) );
  XNOR U14073 ( .A(n14135), .B(n14046), .Z(n14138) );
  XOR U14074 ( .A(n14139), .B(n14129), .Z(n14046) );
  XNOR U14075 ( .A(n14140), .B(n14124), .Z(n14129) );
  XOR U14076 ( .A(n14141), .B(n14142), .Z(n14124) );
  AND U14077 ( .A(n14143), .B(n14144), .Z(n14142) );
  XOR U14078 ( .A(n14145), .B(n14141), .Z(n14143) );
  XNOR U14079 ( .A(n14146), .B(n14147), .Z(n14140) );
  AND U14080 ( .A(n14148), .B(n14149), .Z(n14147) );
  XOR U14081 ( .A(n14146), .B(n14150), .Z(n14148) );
  XNOR U14082 ( .A(n14130), .B(n14127), .Z(n14139) );
  AND U14083 ( .A(n14151), .B(n14152), .Z(n14127) );
  XOR U14084 ( .A(n14153), .B(n14154), .Z(n14130) );
  AND U14085 ( .A(n14155), .B(n14156), .Z(n14154) );
  XOR U14086 ( .A(n14153), .B(n14157), .Z(n14155) );
  XNOR U14087 ( .A(n14043), .B(n14135), .Z(n14137) );
  XOR U14088 ( .A(n14158), .B(n14159), .Z(n14043) );
  AND U14089 ( .A(n287), .B(n14160), .Z(n14159) );
  XNOR U14090 ( .A(n14161), .B(n14158), .Z(n14160) );
  XOR U14091 ( .A(n14162), .B(n14163), .Z(n14135) );
  AND U14092 ( .A(n14164), .B(n14165), .Z(n14163) );
  XNOR U14093 ( .A(n14162), .B(n14151), .Z(n14165) );
  IV U14094 ( .A(n14096), .Z(n14151) );
  XNOR U14095 ( .A(n14166), .B(n14144), .Z(n14096) );
  XNOR U14096 ( .A(n14167), .B(n14150), .Z(n14144) );
  XNOR U14097 ( .A(n14168), .B(n14169), .Z(n14150) );
  NOR U14098 ( .A(n14170), .B(n14171), .Z(n14169) );
  XOR U14099 ( .A(n14168), .B(n14172), .Z(n14170) );
  XNOR U14100 ( .A(n14149), .B(n14141), .Z(n14167) );
  XOR U14101 ( .A(n14173), .B(n14174), .Z(n14141) );
  AND U14102 ( .A(n14175), .B(n14176), .Z(n14174) );
  XOR U14103 ( .A(n14173), .B(n14177), .Z(n14175) );
  XNOR U14104 ( .A(n14178), .B(n14146), .Z(n14149) );
  XOR U14105 ( .A(n14179), .B(n14180), .Z(n14146) );
  AND U14106 ( .A(n14181), .B(n14182), .Z(n14180) );
  XNOR U14107 ( .A(n14183), .B(n14184), .Z(n14181) );
  IV U14108 ( .A(n14179), .Z(n14183) );
  XNOR U14109 ( .A(n14185), .B(n14186), .Z(n14178) );
  NOR U14110 ( .A(n14187), .B(n14188), .Z(n14186) );
  XNOR U14111 ( .A(n14185), .B(n14189), .Z(n14187) );
  XNOR U14112 ( .A(n14145), .B(n14152), .Z(n14166) );
  NOR U14113 ( .A(n14109), .B(n14190), .Z(n14152) );
  XOR U14114 ( .A(n14157), .B(n14156), .Z(n14145) );
  XNOR U14115 ( .A(n14191), .B(n14153), .Z(n14156) );
  XOR U14116 ( .A(n14192), .B(n14193), .Z(n14153) );
  AND U14117 ( .A(n14194), .B(n14195), .Z(n14193) );
  XNOR U14118 ( .A(n14196), .B(n14197), .Z(n14194) );
  IV U14119 ( .A(n14192), .Z(n14196) );
  XNOR U14120 ( .A(n14198), .B(n14199), .Z(n14191) );
  NOR U14121 ( .A(n14200), .B(n14201), .Z(n14199) );
  XNOR U14122 ( .A(n14198), .B(n14202), .Z(n14200) );
  XOR U14123 ( .A(n14203), .B(n14204), .Z(n14157) );
  NOR U14124 ( .A(n14205), .B(n14206), .Z(n14204) );
  XNOR U14125 ( .A(n14203), .B(n14207), .Z(n14205) );
  XNOR U14126 ( .A(n14093), .B(n14162), .Z(n14164) );
  XOR U14127 ( .A(n14208), .B(n14209), .Z(n14093) );
  AND U14128 ( .A(n287), .B(n14210), .Z(n14209) );
  XOR U14129 ( .A(n14211), .B(n14208), .Z(n14210) );
  AND U14130 ( .A(n14106), .B(n14109), .Z(n14162) );
  XOR U14131 ( .A(n14212), .B(n14190), .Z(n14109) );
  XNOR U14132 ( .A(p_input[1120]), .B(p_input[2048]), .Z(n14190) );
  XNOR U14133 ( .A(n14177), .B(n14176), .Z(n14212) );
  XNOR U14134 ( .A(n14213), .B(n14184), .Z(n14176) );
  XNOR U14135 ( .A(n14172), .B(n14171), .Z(n14184) );
  XNOR U14136 ( .A(n14214), .B(n14168), .Z(n14171) );
  XNOR U14137 ( .A(p_input[1130]), .B(p_input[2058]), .Z(n14168) );
  XOR U14138 ( .A(p_input[1131]), .B(n6319), .Z(n14214) );
  XOR U14139 ( .A(p_input[1132]), .B(p_input[2060]), .Z(n14172) );
  XOR U14140 ( .A(n14182), .B(n14215), .Z(n14213) );
  IV U14141 ( .A(n14173), .Z(n14215) );
  XOR U14142 ( .A(p_input[1121]), .B(p_input[2049]), .Z(n14173) );
  XNOR U14143 ( .A(n14216), .B(n14189), .Z(n14182) );
  XNOR U14144 ( .A(p_input[1135]), .B(n6322), .Z(n14189) );
  XOR U14145 ( .A(n14179), .B(n14188), .Z(n14216) );
  XOR U14146 ( .A(n14217), .B(n14185), .Z(n14188) );
  XOR U14147 ( .A(p_input[1133]), .B(p_input[2061]), .Z(n14185) );
  XOR U14148 ( .A(p_input[1134]), .B(n6324), .Z(n14217) );
  XOR U14149 ( .A(p_input[1129]), .B(p_input[2057]), .Z(n14179) );
  XOR U14150 ( .A(n14197), .B(n14195), .Z(n14177) );
  XNOR U14151 ( .A(n14218), .B(n14202), .Z(n14195) );
  XOR U14152 ( .A(p_input[1128]), .B(p_input[2056]), .Z(n14202) );
  XOR U14153 ( .A(n14192), .B(n14201), .Z(n14218) );
  XOR U14154 ( .A(n14219), .B(n14198), .Z(n14201) );
  XOR U14155 ( .A(p_input[1126]), .B(p_input[2054]), .Z(n14198) );
  XOR U14156 ( .A(p_input[1127]), .B(n7007), .Z(n14219) );
  XOR U14157 ( .A(p_input[1122]), .B(p_input[2050]), .Z(n14192) );
  XNOR U14158 ( .A(n14207), .B(n14206), .Z(n14197) );
  XOR U14159 ( .A(n14220), .B(n14203), .Z(n14206) );
  XOR U14160 ( .A(p_input[1123]), .B(p_input[2051]), .Z(n14203) );
  XOR U14161 ( .A(p_input[1124]), .B(n7009), .Z(n14220) );
  XOR U14162 ( .A(p_input[1125]), .B(p_input[2053]), .Z(n14207) );
  XOR U14163 ( .A(n14221), .B(n14222), .Z(n14106) );
  AND U14164 ( .A(n287), .B(n14223), .Z(n14222) );
  XNOR U14165 ( .A(n14224), .B(n14221), .Z(n14223) );
  XNOR U14166 ( .A(n14225), .B(n14226), .Z(n287) );
  AND U14167 ( .A(n14227), .B(n14228), .Z(n14226) );
  XOR U14168 ( .A(n14119), .B(n14225), .Z(n14228) );
  AND U14169 ( .A(n14229), .B(n14230), .Z(n14119) );
  XNOR U14170 ( .A(n14116), .B(n14225), .Z(n14227) );
  XOR U14171 ( .A(n14231), .B(n14232), .Z(n14116) );
  AND U14172 ( .A(n291), .B(n14233), .Z(n14232) );
  XOR U14173 ( .A(n14234), .B(n14231), .Z(n14233) );
  XOR U14174 ( .A(n14235), .B(n14236), .Z(n14225) );
  AND U14175 ( .A(n14237), .B(n14238), .Z(n14236) );
  XNOR U14176 ( .A(n14235), .B(n14229), .Z(n14238) );
  IV U14177 ( .A(n14134), .Z(n14229) );
  XOR U14178 ( .A(n14239), .B(n14240), .Z(n14134) );
  XOR U14179 ( .A(n14241), .B(n14230), .Z(n14240) );
  AND U14180 ( .A(n14161), .B(n14242), .Z(n14230) );
  AND U14181 ( .A(n14243), .B(n14244), .Z(n14241) );
  XOR U14182 ( .A(n14245), .B(n14239), .Z(n14243) );
  XNOR U14183 ( .A(n14131), .B(n14235), .Z(n14237) );
  XOR U14184 ( .A(n14246), .B(n14247), .Z(n14131) );
  AND U14185 ( .A(n291), .B(n14248), .Z(n14247) );
  XOR U14186 ( .A(n14249), .B(n14246), .Z(n14248) );
  XOR U14187 ( .A(n14250), .B(n14251), .Z(n14235) );
  AND U14188 ( .A(n14252), .B(n14253), .Z(n14251) );
  XNOR U14189 ( .A(n14250), .B(n14161), .Z(n14253) );
  XOR U14190 ( .A(n14254), .B(n14244), .Z(n14161) );
  XNOR U14191 ( .A(n14255), .B(n14239), .Z(n14244) );
  XOR U14192 ( .A(n14256), .B(n14257), .Z(n14239) );
  AND U14193 ( .A(n14258), .B(n14259), .Z(n14257) );
  XOR U14194 ( .A(n14260), .B(n14256), .Z(n14258) );
  XNOR U14195 ( .A(n14261), .B(n14262), .Z(n14255) );
  AND U14196 ( .A(n14263), .B(n14264), .Z(n14262) );
  XOR U14197 ( .A(n14261), .B(n14265), .Z(n14263) );
  XNOR U14198 ( .A(n14245), .B(n14242), .Z(n14254) );
  AND U14199 ( .A(n14266), .B(n14267), .Z(n14242) );
  XOR U14200 ( .A(n14268), .B(n14269), .Z(n14245) );
  AND U14201 ( .A(n14270), .B(n14271), .Z(n14269) );
  XOR U14202 ( .A(n14268), .B(n14272), .Z(n14270) );
  XNOR U14203 ( .A(n14158), .B(n14250), .Z(n14252) );
  XOR U14204 ( .A(n14273), .B(n14274), .Z(n14158) );
  AND U14205 ( .A(n291), .B(n14275), .Z(n14274) );
  XNOR U14206 ( .A(n14276), .B(n14273), .Z(n14275) );
  XOR U14207 ( .A(n14277), .B(n14278), .Z(n14250) );
  AND U14208 ( .A(n14279), .B(n14280), .Z(n14278) );
  XNOR U14209 ( .A(n14277), .B(n14266), .Z(n14280) );
  IV U14210 ( .A(n14211), .Z(n14266) );
  XNOR U14211 ( .A(n14281), .B(n14259), .Z(n14211) );
  XNOR U14212 ( .A(n14282), .B(n14265), .Z(n14259) );
  XNOR U14213 ( .A(n14283), .B(n14284), .Z(n14265) );
  NOR U14214 ( .A(n14285), .B(n14286), .Z(n14284) );
  XOR U14215 ( .A(n14283), .B(n14287), .Z(n14285) );
  XNOR U14216 ( .A(n14264), .B(n14256), .Z(n14282) );
  XOR U14217 ( .A(n14288), .B(n14289), .Z(n14256) );
  AND U14218 ( .A(n14290), .B(n14291), .Z(n14289) );
  XOR U14219 ( .A(n14288), .B(n14292), .Z(n14290) );
  XNOR U14220 ( .A(n14293), .B(n14261), .Z(n14264) );
  XOR U14221 ( .A(n14294), .B(n14295), .Z(n14261) );
  AND U14222 ( .A(n14296), .B(n14297), .Z(n14295) );
  XNOR U14223 ( .A(n14298), .B(n14299), .Z(n14296) );
  IV U14224 ( .A(n14294), .Z(n14298) );
  XNOR U14225 ( .A(n14300), .B(n14301), .Z(n14293) );
  NOR U14226 ( .A(n14302), .B(n14303), .Z(n14301) );
  XNOR U14227 ( .A(n14300), .B(n14304), .Z(n14302) );
  XNOR U14228 ( .A(n14260), .B(n14267), .Z(n14281) );
  NOR U14229 ( .A(n14224), .B(n14305), .Z(n14267) );
  XOR U14230 ( .A(n14272), .B(n14271), .Z(n14260) );
  XNOR U14231 ( .A(n14306), .B(n14268), .Z(n14271) );
  XOR U14232 ( .A(n14307), .B(n14308), .Z(n14268) );
  AND U14233 ( .A(n14309), .B(n14310), .Z(n14308) );
  XNOR U14234 ( .A(n14311), .B(n14312), .Z(n14309) );
  IV U14235 ( .A(n14307), .Z(n14311) );
  XNOR U14236 ( .A(n14313), .B(n14314), .Z(n14306) );
  NOR U14237 ( .A(n14315), .B(n14316), .Z(n14314) );
  XNOR U14238 ( .A(n14313), .B(n14317), .Z(n14315) );
  XOR U14239 ( .A(n14318), .B(n14319), .Z(n14272) );
  NOR U14240 ( .A(n14320), .B(n14321), .Z(n14319) );
  XNOR U14241 ( .A(n14318), .B(n14322), .Z(n14320) );
  XNOR U14242 ( .A(n14208), .B(n14277), .Z(n14279) );
  XOR U14243 ( .A(n14323), .B(n14324), .Z(n14208) );
  AND U14244 ( .A(n291), .B(n14325), .Z(n14324) );
  XOR U14245 ( .A(n14326), .B(n14323), .Z(n14325) );
  AND U14246 ( .A(n14221), .B(n14224), .Z(n14277) );
  XOR U14247 ( .A(n14327), .B(n14305), .Z(n14224) );
  XNOR U14248 ( .A(p_input[1136]), .B(p_input[2048]), .Z(n14305) );
  XNOR U14249 ( .A(n14292), .B(n14291), .Z(n14327) );
  XNOR U14250 ( .A(n14328), .B(n14299), .Z(n14291) );
  XNOR U14251 ( .A(n14287), .B(n14286), .Z(n14299) );
  XNOR U14252 ( .A(n14329), .B(n14283), .Z(n14286) );
  XNOR U14253 ( .A(p_input[1146]), .B(p_input[2058]), .Z(n14283) );
  XOR U14254 ( .A(p_input[1147]), .B(n6319), .Z(n14329) );
  XOR U14255 ( .A(p_input[1148]), .B(p_input[2060]), .Z(n14287) );
  XOR U14256 ( .A(n14297), .B(n14330), .Z(n14328) );
  IV U14257 ( .A(n14288), .Z(n14330) );
  XOR U14258 ( .A(p_input[1137]), .B(p_input[2049]), .Z(n14288) );
  XNOR U14259 ( .A(n14331), .B(n14304), .Z(n14297) );
  XNOR U14260 ( .A(p_input[1151]), .B(n6322), .Z(n14304) );
  XOR U14261 ( .A(n14294), .B(n14303), .Z(n14331) );
  XOR U14262 ( .A(n14332), .B(n14300), .Z(n14303) );
  XOR U14263 ( .A(p_input[1149]), .B(p_input[2061]), .Z(n14300) );
  XOR U14264 ( .A(p_input[1150]), .B(n6324), .Z(n14332) );
  XOR U14265 ( .A(p_input[1145]), .B(p_input[2057]), .Z(n14294) );
  XOR U14266 ( .A(n14312), .B(n14310), .Z(n14292) );
  XNOR U14267 ( .A(n14333), .B(n14317), .Z(n14310) );
  XOR U14268 ( .A(p_input[1144]), .B(p_input[2056]), .Z(n14317) );
  XOR U14269 ( .A(n14307), .B(n14316), .Z(n14333) );
  XOR U14270 ( .A(n14334), .B(n14313), .Z(n14316) );
  XOR U14271 ( .A(p_input[1142]), .B(p_input[2054]), .Z(n14313) );
  XOR U14272 ( .A(p_input[1143]), .B(n7007), .Z(n14334) );
  XOR U14273 ( .A(p_input[1138]), .B(p_input[2050]), .Z(n14307) );
  XNOR U14274 ( .A(n14322), .B(n14321), .Z(n14312) );
  XOR U14275 ( .A(n14335), .B(n14318), .Z(n14321) );
  XOR U14276 ( .A(p_input[1139]), .B(p_input[2051]), .Z(n14318) );
  XOR U14277 ( .A(p_input[1140]), .B(n7009), .Z(n14335) );
  XOR U14278 ( .A(p_input[1141]), .B(p_input[2053]), .Z(n14322) );
  XOR U14279 ( .A(n14336), .B(n14337), .Z(n14221) );
  AND U14280 ( .A(n291), .B(n14338), .Z(n14337) );
  XNOR U14281 ( .A(n14339), .B(n14336), .Z(n14338) );
  XNOR U14282 ( .A(n14340), .B(n14341), .Z(n291) );
  AND U14283 ( .A(n14342), .B(n14343), .Z(n14341) );
  XOR U14284 ( .A(n14234), .B(n14340), .Z(n14343) );
  AND U14285 ( .A(n14344), .B(n14345), .Z(n14234) );
  XNOR U14286 ( .A(n14231), .B(n14340), .Z(n14342) );
  XOR U14287 ( .A(n14346), .B(n14347), .Z(n14231) );
  AND U14288 ( .A(n295), .B(n14348), .Z(n14347) );
  XOR U14289 ( .A(n14349), .B(n14346), .Z(n14348) );
  XOR U14290 ( .A(n14350), .B(n14351), .Z(n14340) );
  AND U14291 ( .A(n14352), .B(n14353), .Z(n14351) );
  XNOR U14292 ( .A(n14350), .B(n14344), .Z(n14353) );
  IV U14293 ( .A(n14249), .Z(n14344) );
  XOR U14294 ( .A(n14354), .B(n14355), .Z(n14249) );
  XOR U14295 ( .A(n14356), .B(n14345), .Z(n14355) );
  AND U14296 ( .A(n14276), .B(n14357), .Z(n14345) );
  AND U14297 ( .A(n14358), .B(n14359), .Z(n14356) );
  XOR U14298 ( .A(n14360), .B(n14354), .Z(n14358) );
  XNOR U14299 ( .A(n14246), .B(n14350), .Z(n14352) );
  XOR U14300 ( .A(n14361), .B(n14362), .Z(n14246) );
  AND U14301 ( .A(n295), .B(n14363), .Z(n14362) );
  XOR U14302 ( .A(n14364), .B(n14361), .Z(n14363) );
  XOR U14303 ( .A(n14365), .B(n14366), .Z(n14350) );
  AND U14304 ( .A(n14367), .B(n14368), .Z(n14366) );
  XNOR U14305 ( .A(n14365), .B(n14276), .Z(n14368) );
  XOR U14306 ( .A(n14369), .B(n14359), .Z(n14276) );
  XNOR U14307 ( .A(n14370), .B(n14354), .Z(n14359) );
  XOR U14308 ( .A(n14371), .B(n14372), .Z(n14354) );
  AND U14309 ( .A(n14373), .B(n14374), .Z(n14372) );
  XOR U14310 ( .A(n14375), .B(n14371), .Z(n14373) );
  XNOR U14311 ( .A(n14376), .B(n14377), .Z(n14370) );
  AND U14312 ( .A(n14378), .B(n14379), .Z(n14377) );
  XOR U14313 ( .A(n14376), .B(n14380), .Z(n14378) );
  XNOR U14314 ( .A(n14360), .B(n14357), .Z(n14369) );
  AND U14315 ( .A(n14381), .B(n14382), .Z(n14357) );
  XOR U14316 ( .A(n14383), .B(n14384), .Z(n14360) );
  AND U14317 ( .A(n14385), .B(n14386), .Z(n14384) );
  XOR U14318 ( .A(n14383), .B(n14387), .Z(n14385) );
  XNOR U14319 ( .A(n14273), .B(n14365), .Z(n14367) );
  XOR U14320 ( .A(n14388), .B(n14389), .Z(n14273) );
  AND U14321 ( .A(n295), .B(n14390), .Z(n14389) );
  XNOR U14322 ( .A(n14391), .B(n14388), .Z(n14390) );
  XOR U14323 ( .A(n14392), .B(n14393), .Z(n14365) );
  AND U14324 ( .A(n14394), .B(n14395), .Z(n14393) );
  XNOR U14325 ( .A(n14392), .B(n14381), .Z(n14395) );
  IV U14326 ( .A(n14326), .Z(n14381) );
  XNOR U14327 ( .A(n14396), .B(n14374), .Z(n14326) );
  XNOR U14328 ( .A(n14397), .B(n14380), .Z(n14374) );
  XNOR U14329 ( .A(n14398), .B(n14399), .Z(n14380) );
  NOR U14330 ( .A(n14400), .B(n14401), .Z(n14399) );
  XOR U14331 ( .A(n14398), .B(n14402), .Z(n14400) );
  XNOR U14332 ( .A(n14379), .B(n14371), .Z(n14397) );
  XOR U14333 ( .A(n14403), .B(n14404), .Z(n14371) );
  AND U14334 ( .A(n14405), .B(n14406), .Z(n14404) );
  XOR U14335 ( .A(n14403), .B(n14407), .Z(n14405) );
  XNOR U14336 ( .A(n14408), .B(n14376), .Z(n14379) );
  XOR U14337 ( .A(n14409), .B(n14410), .Z(n14376) );
  AND U14338 ( .A(n14411), .B(n14412), .Z(n14410) );
  XNOR U14339 ( .A(n14413), .B(n14414), .Z(n14411) );
  IV U14340 ( .A(n14409), .Z(n14413) );
  XNOR U14341 ( .A(n14415), .B(n14416), .Z(n14408) );
  NOR U14342 ( .A(n14417), .B(n14418), .Z(n14416) );
  XNOR U14343 ( .A(n14415), .B(n14419), .Z(n14417) );
  XNOR U14344 ( .A(n14375), .B(n14382), .Z(n14396) );
  NOR U14345 ( .A(n14339), .B(n14420), .Z(n14382) );
  XOR U14346 ( .A(n14387), .B(n14386), .Z(n14375) );
  XNOR U14347 ( .A(n14421), .B(n14383), .Z(n14386) );
  XOR U14348 ( .A(n14422), .B(n14423), .Z(n14383) );
  AND U14349 ( .A(n14424), .B(n14425), .Z(n14423) );
  XNOR U14350 ( .A(n14426), .B(n14427), .Z(n14424) );
  IV U14351 ( .A(n14422), .Z(n14426) );
  XNOR U14352 ( .A(n14428), .B(n14429), .Z(n14421) );
  NOR U14353 ( .A(n14430), .B(n14431), .Z(n14429) );
  XNOR U14354 ( .A(n14428), .B(n14432), .Z(n14430) );
  XOR U14355 ( .A(n14433), .B(n14434), .Z(n14387) );
  NOR U14356 ( .A(n14435), .B(n14436), .Z(n14434) );
  XNOR U14357 ( .A(n14433), .B(n14437), .Z(n14435) );
  XNOR U14358 ( .A(n14323), .B(n14392), .Z(n14394) );
  XOR U14359 ( .A(n14438), .B(n14439), .Z(n14323) );
  AND U14360 ( .A(n295), .B(n14440), .Z(n14439) );
  XOR U14361 ( .A(n14441), .B(n14438), .Z(n14440) );
  AND U14362 ( .A(n14336), .B(n14339), .Z(n14392) );
  XOR U14363 ( .A(n14442), .B(n14420), .Z(n14339) );
  XNOR U14364 ( .A(p_input[1152]), .B(p_input[2048]), .Z(n14420) );
  XNOR U14365 ( .A(n14407), .B(n14406), .Z(n14442) );
  XNOR U14366 ( .A(n14443), .B(n14414), .Z(n14406) );
  XNOR U14367 ( .A(n14402), .B(n14401), .Z(n14414) );
  XNOR U14368 ( .A(n14444), .B(n14398), .Z(n14401) );
  XNOR U14369 ( .A(p_input[1162]), .B(p_input[2058]), .Z(n14398) );
  XOR U14370 ( .A(p_input[1163]), .B(n6319), .Z(n14444) );
  XOR U14371 ( .A(p_input[1164]), .B(p_input[2060]), .Z(n14402) );
  XOR U14372 ( .A(n14412), .B(n14445), .Z(n14443) );
  IV U14373 ( .A(n14403), .Z(n14445) );
  XOR U14374 ( .A(p_input[1153]), .B(p_input[2049]), .Z(n14403) );
  XNOR U14375 ( .A(n14446), .B(n14419), .Z(n14412) );
  XNOR U14376 ( .A(p_input[1167]), .B(n6322), .Z(n14419) );
  XOR U14377 ( .A(n14409), .B(n14418), .Z(n14446) );
  XOR U14378 ( .A(n14447), .B(n14415), .Z(n14418) );
  XOR U14379 ( .A(p_input[1165]), .B(p_input[2061]), .Z(n14415) );
  XOR U14380 ( .A(p_input[1166]), .B(n6324), .Z(n14447) );
  XOR U14381 ( .A(p_input[1161]), .B(p_input[2057]), .Z(n14409) );
  XOR U14382 ( .A(n14427), .B(n14425), .Z(n14407) );
  XNOR U14383 ( .A(n14448), .B(n14432), .Z(n14425) );
  XOR U14384 ( .A(p_input[1160]), .B(p_input[2056]), .Z(n14432) );
  XOR U14385 ( .A(n14422), .B(n14431), .Z(n14448) );
  XOR U14386 ( .A(n14449), .B(n14428), .Z(n14431) );
  XOR U14387 ( .A(p_input[1158]), .B(p_input[2054]), .Z(n14428) );
  XOR U14388 ( .A(p_input[1159]), .B(n7007), .Z(n14449) );
  XOR U14389 ( .A(p_input[1154]), .B(p_input[2050]), .Z(n14422) );
  XNOR U14390 ( .A(n14437), .B(n14436), .Z(n14427) );
  XOR U14391 ( .A(n14450), .B(n14433), .Z(n14436) );
  XOR U14392 ( .A(p_input[1155]), .B(p_input[2051]), .Z(n14433) );
  XOR U14393 ( .A(p_input[1156]), .B(n7009), .Z(n14450) );
  XOR U14394 ( .A(p_input[1157]), .B(p_input[2053]), .Z(n14437) );
  XOR U14395 ( .A(n14451), .B(n14452), .Z(n14336) );
  AND U14396 ( .A(n295), .B(n14453), .Z(n14452) );
  XNOR U14397 ( .A(n14454), .B(n14451), .Z(n14453) );
  XNOR U14398 ( .A(n14455), .B(n14456), .Z(n295) );
  AND U14399 ( .A(n14457), .B(n14458), .Z(n14456) );
  XOR U14400 ( .A(n14349), .B(n14455), .Z(n14458) );
  AND U14401 ( .A(n14459), .B(n14460), .Z(n14349) );
  XNOR U14402 ( .A(n14346), .B(n14455), .Z(n14457) );
  XOR U14403 ( .A(n14461), .B(n14462), .Z(n14346) );
  AND U14404 ( .A(n299), .B(n14463), .Z(n14462) );
  XOR U14405 ( .A(n14464), .B(n14461), .Z(n14463) );
  XOR U14406 ( .A(n14465), .B(n14466), .Z(n14455) );
  AND U14407 ( .A(n14467), .B(n14468), .Z(n14466) );
  XNOR U14408 ( .A(n14465), .B(n14459), .Z(n14468) );
  IV U14409 ( .A(n14364), .Z(n14459) );
  XOR U14410 ( .A(n14469), .B(n14470), .Z(n14364) );
  XOR U14411 ( .A(n14471), .B(n14460), .Z(n14470) );
  AND U14412 ( .A(n14391), .B(n14472), .Z(n14460) );
  AND U14413 ( .A(n14473), .B(n14474), .Z(n14471) );
  XOR U14414 ( .A(n14475), .B(n14469), .Z(n14473) );
  XNOR U14415 ( .A(n14361), .B(n14465), .Z(n14467) );
  XOR U14416 ( .A(n14476), .B(n14477), .Z(n14361) );
  AND U14417 ( .A(n299), .B(n14478), .Z(n14477) );
  XOR U14418 ( .A(n14479), .B(n14476), .Z(n14478) );
  XOR U14419 ( .A(n14480), .B(n14481), .Z(n14465) );
  AND U14420 ( .A(n14482), .B(n14483), .Z(n14481) );
  XNOR U14421 ( .A(n14480), .B(n14391), .Z(n14483) );
  XOR U14422 ( .A(n14484), .B(n14474), .Z(n14391) );
  XNOR U14423 ( .A(n14485), .B(n14469), .Z(n14474) );
  XOR U14424 ( .A(n14486), .B(n14487), .Z(n14469) );
  AND U14425 ( .A(n14488), .B(n14489), .Z(n14487) );
  XOR U14426 ( .A(n14490), .B(n14486), .Z(n14488) );
  XNOR U14427 ( .A(n14491), .B(n14492), .Z(n14485) );
  AND U14428 ( .A(n14493), .B(n14494), .Z(n14492) );
  XOR U14429 ( .A(n14491), .B(n14495), .Z(n14493) );
  XNOR U14430 ( .A(n14475), .B(n14472), .Z(n14484) );
  AND U14431 ( .A(n14496), .B(n14497), .Z(n14472) );
  XOR U14432 ( .A(n14498), .B(n14499), .Z(n14475) );
  AND U14433 ( .A(n14500), .B(n14501), .Z(n14499) );
  XOR U14434 ( .A(n14498), .B(n14502), .Z(n14500) );
  XNOR U14435 ( .A(n14388), .B(n14480), .Z(n14482) );
  XOR U14436 ( .A(n14503), .B(n14504), .Z(n14388) );
  AND U14437 ( .A(n299), .B(n14505), .Z(n14504) );
  XNOR U14438 ( .A(n14506), .B(n14503), .Z(n14505) );
  XOR U14439 ( .A(n14507), .B(n14508), .Z(n14480) );
  AND U14440 ( .A(n14509), .B(n14510), .Z(n14508) );
  XNOR U14441 ( .A(n14507), .B(n14496), .Z(n14510) );
  IV U14442 ( .A(n14441), .Z(n14496) );
  XNOR U14443 ( .A(n14511), .B(n14489), .Z(n14441) );
  XNOR U14444 ( .A(n14512), .B(n14495), .Z(n14489) );
  XNOR U14445 ( .A(n14513), .B(n14514), .Z(n14495) );
  NOR U14446 ( .A(n14515), .B(n14516), .Z(n14514) );
  XOR U14447 ( .A(n14513), .B(n14517), .Z(n14515) );
  XNOR U14448 ( .A(n14494), .B(n14486), .Z(n14512) );
  XOR U14449 ( .A(n14518), .B(n14519), .Z(n14486) );
  AND U14450 ( .A(n14520), .B(n14521), .Z(n14519) );
  XOR U14451 ( .A(n14518), .B(n14522), .Z(n14520) );
  XNOR U14452 ( .A(n14523), .B(n14491), .Z(n14494) );
  XOR U14453 ( .A(n14524), .B(n14525), .Z(n14491) );
  AND U14454 ( .A(n14526), .B(n14527), .Z(n14525) );
  XNOR U14455 ( .A(n14528), .B(n14529), .Z(n14526) );
  IV U14456 ( .A(n14524), .Z(n14528) );
  XNOR U14457 ( .A(n14530), .B(n14531), .Z(n14523) );
  NOR U14458 ( .A(n14532), .B(n14533), .Z(n14531) );
  XNOR U14459 ( .A(n14530), .B(n14534), .Z(n14532) );
  XNOR U14460 ( .A(n14490), .B(n14497), .Z(n14511) );
  NOR U14461 ( .A(n14454), .B(n14535), .Z(n14497) );
  XOR U14462 ( .A(n14502), .B(n14501), .Z(n14490) );
  XNOR U14463 ( .A(n14536), .B(n14498), .Z(n14501) );
  XOR U14464 ( .A(n14537), .B(n14538), .Z(n14498) );
  AND U14465 ( .A(n14539), .B(n14540), .Z(n14538) );
  XNOR U14466 ( .A(n14541), .B(n14542), .Z(n14539) );
  IV U14467 ( .A(n14537), .Z(n14541) );
  XNOR U14468 ( .A(n14543), .B(n14544), .Z(n14536) );
  NOR U14469 ( .A(n14545), .B(n14546), .Z(n14544) );
  XNOR U14470 ( .A(n14543), .B(n14547), .Z(n14545) );
  XOR U14471 ( .A(n14548), .B(n14549), .Z(n14502) );
  NOR U14472 ( .A(n14550), .B(n14551), .Z(n14549) );
  XNOR U14473 ( .A(n14548), .B(n14552), .Z(n14550) );
  XNOR U14474 ( .A(n14438), .B(n14507), .Z(n14509) );
  XOR U14475 ( .A(n14553), .B(n14554), .Z(n14438) );
  AND U14476 ( .A(n299), .B(n14555), .Z(n14554) );
  XOR U14477 ( .A(n14556), .B(n14553), .Z(n14555) );
  AND U14478 ( .A(n14451), .B(n14454), .Z(n14507) );
  XOR U14479 ( .A(n14557), .B(n14535), .Z(n14454) );
  XNOR U14480 ( .A(p_input[1168]), .B(p_input[2048]), .Z(n14535) );
  XNOR U14481 ( .A(n14522), .B(n14521), .Z(n14557) );
  XNOR U14482 ( .A(n14558), .B(n14529), .Z(n14521) );
  XNOR U14483 ( .A(n14517), .B(n14516), .Z(n14529) );
  XNOR U14484 ( .A(n14559), .B(n14513), .Z(n14516) );
  XNOR U14485 ( .A(p_input[1178]), .B(p_input[2058]), .Z(n14513) );
  XOR U14486 ( .A(p_input[1179]), .B(n6319), .Z(n14559) );
  XOR U14487 ( .A(p_input[1180]), .B(p_input[2060]), .Z(n14517) );
  XOR U14488 ( .A(n14527), .B(n14560), .Z(n14558) );
  IV U14489 ( .A(n14518), .Z(n14560) );
  XOR U14490 ( .A(p_input[1169]), .B(p_input[2049]), .Z(n14518) );
  XNOR U14491 ( .A(n14561), .B(n14534), .Z(n14527) );
  XNOR U14492 ( .A(p_input[1183]), .B(n6322), .Z(n14534) );
  XOR U14493 ( .A(n14524), .B(n14533), .Z(n14561) );
  XOR U14494 ( .A(n14562), .B(n14530), .Z(n14533) );
  XOR U14495 ( .A(p_input[1181]), .B(p_input[2061]), .Z(n14530) );
  XOR U14496 ( .A(p_input[1182]), .B(n6324), .Z(n14562) );
  XOR U14497 ( .A(p_input[1177]), .B(p_input[2057]), .Z(n14524) );
  XOR U14498 ( .A(n14542), .B(n14540), .Z(n14522) );
  XNOR U14499 ( .A(n14563), .B(n14547), .Z(n14540) );
  XOR U14500 ( .A(p_input[1176]), .B(p_input[2056]), .Z(n14547) );
  XOR U14501 ( .A(n14537), .B(n14546), .Z(n14563) );
  XOR U14502 ( .A(n14564), .B(n14543), .Z(n14546) );
  XOR U14503 ( .A(p_input[1174]), .B(p_input[2054]), .Z(n14543) );
  XOR U14504 ( .A(p_input[1175]), .B(n7007), .Z(n14564) );
  XOR U14505 ( .A(p_input[1170]), .B(p_input[2050]), .Z(n14537) );
  XNOR U14506 ( .A(n14552), .B(n14551), .Z(n14542) );
  XOR U14507 ( .A(n14565), .B(n14548), .Z(n14551) );
  XOR U14508 ( .A(p_input[1171]), .B(p_input[2051]), .Z(n14548) );
  XOR U14509 ( .A(p_input[1172]), .B(n7009), .Z(n14565) );
  XOR U14510 ( .A(p_input[1173]), .B(p_input[2053]), .Z(n14552) );
  XOR U14511 ( .A(n14566), .B(n14567), .Z(n14451) );
  AND U14512 ( .A(n299), .B(n14568), .Z(n14567) );
  XNOR U14513 ( .A(n14569), .B(n14566), .Z(n14568) );
  XNOR U14514 ( .A(n14570), .B(n14571), .Z(n299) );
  AND U14515 ( .A(n14572), .B(n14573), .Z(n14571) );
  XOR U14516 ( .A(n14464), .B(n14570), .Z(n14573) );
  AND U14517 ( .A(n14574), .B(n14575), .Z(n14464) );
  XNOR U14518 ( .A(n14461), .B(n14570), .Z(n14572) );
  XOR U14519 ( .A(n14576), .B(n14577), .Z(n14461) );
  AND U14520 ( .A(n303), .B(n14578), .Z(n14577) );
  XOR U14521 ( .A(n14579), .B(n14576), .Z(n14578) );
  XOR U14522 ( .A(n14580), .B(n14581), .Z(n14570) );
  AND U14523 ( .A(n14582), .B(n14583), .Z(n14581) );
  XNOR U14524 ( .A(n14580), .B(n14574), .Z(n14583) );
  IV U14525 ( .A(n14479), .Z(n14574) );
  XOR U14526 ( .A(n14584), .B(n14585), .Z(n14479) );
  XOR U14527 ( .A(n14586), .B(n14575), .Z(n14585) );
  AND U14528 ( .A(n14506), .B(n14587), .Z(n14575) );
  AND U14529 ( .A(n14588), .B(n14589), .Z(n14586) );
  XOR U14530 ( .A(n14590), .B(n14584), .Z(n14588) );
  XNOR U14531 ( .A(n14476), .B(n14580), .Z(n14582) );
  XOR U14532 ( .A(n14591), .B(n14592), .Z(n14476) );
  AND U14533 ( .A(n303), .B(n14593), .Z(n14592) );
  XOR U14534 ( .A(n14594), .B(n14591), .Z(n14593) );
  XOR U14535 ( .A(n14595), .B(n14596), .Z(n14580) );
  AND U14536 ( .A(n14597), .B(n14598), .Z(n14596) );
  XNOR U14537 ( .A(n14595), .B(n14506), .Z(n14598) );
  XOR U14538 ( .A(n14599), .B(n14589), .Z(n14506) );
  XNOR U14539 ( .A(n14600), .B(n14584), .Z(n14589) );
  XOR U14540 ( .A(n14601), .B(n14602), .Z(n14584) );
  AND U14541 ( .A(n14603), .B(n14604), .Z(n14602) );
  XOR U14542 ( .A(n14605), .B(n14601), .Z(n14603) );
  XNOR U14543 ( .A(n14606), .B(n14607), .Z(n14600) );
  AND U14544 ( .A(n14608), .B(n14609), .Z(n14607) );
  XOR U14545 ( .A(n14606), .B(n14610), .Z(n14608) );
  XNOR U14546 ( .A(n14590), .B(n14587), .Z(n14599) );
  AND U14547 ( .A(n14611), .B(n14612), .Z(n14587) );
  XOR U14548 ( .A(n14613), .B(n14614), .Z(n14590) );
  AND U14549 ( .A(n14615), .B(n14616), .Z(n14614) );
  XOR U14550 ( .A(n14613), .B(n14617), .Z(n14615) );
  XNOR U14551 ( .A(n14503), .B(n14595), .Z(n14597) );
  XOR U14552 ( .A(n14618), .B(n14619), .Z(n14503) );
  AND U14553 ( .A(n303), .B(n14620), .Z(n14619) );
  XNOR U14554 ( .A(n14621), .B(n14618), .Z(n14620) );
  XOR U14555 ( .A(n14622), .B(n14623), .Z(n14595) );
  AND U14556 ( .A(n14624), .B(n14625), .Z(n14623) );
  XNOR U14557 ( .A(n14622), .B(n14611), .Z(n14625) );
  IV U14558 ( .A(n14556), .Z(n14611) );
  XNOR U14559 ( .A(n14626), .B(n14604), .Z(n14556) );
  XNOR U14560 ( .A(n14627), .B(n14610), .Z(n14604) );
  XNOR U14561 ( .A(n14628), .B(n14629), .Z(n14610) );
  NOR U14562 ( .A(n14630), .B(n14631), .Z(n14629) );
  XOR U14563 ( .A(n14628), .B(n14632), .Z(n14630) );
  XNOR U14564 ( .A(n14609), .B(n14601), .Z(n14627) );
  XOR U14565 ( .A(n14633), .B(n14634), .Z(n14601) );
  AND U14566 ( .A(n14635), .B(n14636), .Z(n14634) );
  XOR U14567 ( .A(n14633), .B(n14637), .Z(n14635) );
  XNOR U14568 ( .A(n14638), .B(n14606), .Z(n14609) );
  XOR U14569 ( .A(n14639), .B(n14640), .Z(n14606) );
  AND U14570 ( .A(n14641), .B(n14642), .Z(n14640) );
  XNOR U14571 ( .A(n14643), .B(n14644), .Z(n14641) );
  IV U14572 ( .A(n14639), .Z(n14643) );
  XNOR U14573 ( .A(n14645), .B(n14646), .Z(n14638) );
  NOR U14574 ( .A(n14647), .B(n14648), .Z(n14646) );
  XNOR U14575 ( .A(n14645), .B(n14649), .Z(n14647) );
  XNOR U14576 ( .A(n14605), .B(n14612), .Z(n14626) );
  NOR U14577 ( .A(n14569), .B(n14650), .Z(n14612) );
  XOR U14578 ( .A(n14617), .B(n14616), .Z(n14605) );
  XNOR U14579 ( .A(n14651), .B(n14613), .Z(n14616) );
  XOR U14580 ( .A(n14652), .B(n14653), .Z(n14613) );
  AND U14581 ( .A(n14654), .B(n14655), .Z(n14653) );
  XNOR U14582 ( .A(n14656), .B(n14657), .Z(n14654) );
  IV U14583 ( .A(n14652), .Z(n14656) );
  XNOR U14584 ( .A(n14658), .B(n14659), .Z(n14651) );
  NOR U14585 ( .A(n14660), .B(n14661), .Z(n14659) );
  XNOR U14586 ( .A(n14658), .B(n14662), .Z(n14660) );
  XOR U14587 ( .A(n14663), .B(n14664), .Z(n14617) );
  NOR U14588 ( .A(n14665), .B(n14666), .Z(n14664) );
  XNOR U14589 ( .A(n14663), .B(n14667), .Z(n14665) );
  XNOR U14590 ( .A(n14553), .B(n14622), .Z(n14624) );
  XOR U14591 ( .A(n14668), .B(n14669), .Z(n14553) );
  AND U14592 ( .A(n303), .B(n14670), .Z(n14669) );
  XOR U14593 ( .A(n14671), .B(n14668), .Z(n14670) );
  AND U14594 ( .A(n14566), .B(n14569), .Z(n14622) );
  XOR U14595 ( .A(n14672), .B(n14650), .Z(n14569) );
  XNOR U14596 ( .A(p_input[1184]), .B(p_input[2048]), .Z(n14650) );
  XNOR U14597 ( .A(n14637), .B(n14636), .Z(n14672) );
  XNOR U14598 ( .A(n14673), .B(n14644), .Z(n14636) );
  XNOR U14599 ( .A(n14632), .B(n14631), .Z(n14644) );
  XNOR U14600 ( .A(n14674), .B(n14628), .Z(n14631) );
  XNOR U14601 ( .A(p_input[1194]), .B(p_input[2058]), .Z(n14628) );
  XOR U14602 ( .A(p_input[1195]), .B(n6319), .Z(n14674) );
  XOR U14603 ( .A(p_input[1196]), .B(p_input[2060]), .Z(n14632) );
  XOR U14604 ( .A(n14642), .B(n14675), .Z(n14673) );
  IV U14605 ( .A(n14633), .Z(n14675) );
  XOR U14606 ( .A(p_input[1185]), .B(p_input[2049]), .Z(n14633) );
  XNOR U14607 ( .A(n14676), .B(n14649), .Z(n14642) );
  XNOR U14608 ( .A(p_input[1199]), .B(n6322), .Z(n14649) );
  XOR U14609 ( .A(n14639), .B(n14648), .Z(n14676) );
  XOR U14610 ( .A(n14677), .B(n14645), .Z(n14648) );
  XOR U14611 ( .A(p_input[1197]), .B(p_input[2061]), .Z(n14645) );
  XOR U14612 ( .A(p_input[1198]), .B(n6324), .Z(n14677) );
  XOR U14613 ( .A(p_input[1193]), .B(p_input[2057]), .Z(n14639) );
  XOR U14614 ( .A(n14657), .B(n14655), .Z(n14637) );
  XNOR U14615 ( .A(n14678), .B(n14662), .Z(n14655) );
  XOR U14616 ( .A(p_input[1192]), .B(p_input[2056]), .Z(n14662) );
  XOR U14617 ( .A(n14652), .B(n14661), .Z(n14678) );
  XOR U14618 ( .A(n14679), .B(n14658), .Z(n14661) );
  XOR U14619 ( .A(p_input[1190]), .B(p_input[2054]), .Z(n14658) );
  XOR U14620 ( .A(p_input[1191]), .B(n7007), .Z(n14679) );
  XOR U14621 ( .A(p_input[1186]), .B(p_input[2050]), .Z(n14652) );
  XNOR U14622 ( .A(n14667), .B(n14666), .Z(n14657) );
  XOR U14623 ( .A(n14680), .B(n14663), .Z(n14666) );
  XOR U14624 ( .A(p_input[1187]), .B(p_input[2051]), .Z(n14663) );
  XOR U14625 ( .A(p_input[1188]), .B(n7009), .Z(n14680) );
  XOR U14626 ( .A(p_input[1189]), .B(p_input[2053]), .Z(n14667) );
  XOR U14627 ( .A(n14681), .B(n14682), .Z(n14566) );
  AND U14628 ( .A(n303), .B(n14683), .Z(n14682) );
  XNOR U14629 ( .A(n14684), .B(n14681), .Z(n14683) );
  XNOR U14630 ( .A(n14685), .B(n14686), .Z(n303) );
  AND U14631 ( .A(n14687), .B(n14688), .Z(n14686) );
  XOR U14632 ( .A(n14579), .B(n14685), .Z(n14688) );
  AND U14633 ( .A(n14689), .B(n14690), .Z(n14579) );
  XNOR U14634 ( .A(n14576), .B(n14685), .Z(n14687) );
  XOR U14635 ( .A(n14691), .B(n14692), .Z(n14576) );
  AND U14636 ( .A(n307), .B(n14693), .Z(n14692) );
  XOR U14637 ( .A(n14694), .B(n14691), .Z(n14693) );
  XOR U14638 ( .A(n14695), .B(n14696), .Z(n14685) );
  AND U14639 ( .A(n14697), .B(n14698), .Z(n14696) );
  XNOR U14640 ( .A(n14695), .B(n14689), .Z(n14698) );
  IV U14641 ( .A(n14594), .Z(n14689) );
  XOR U14642 ( .A(n14699), .B(n14700), .Z(n14594) );
  XOR U14643 ( .A(n14701), .B(n14690), .Z(n14700) );
  AND U14644 ( .A(n14621), .B(n14702), .Z(n14690) );
  AND U14645 ( .A(n14703), .B(n14704), .Z(n14701) );
  XOR U14646 ( .A(n14705), .B(n14699), .Z(n14703) );
  XNOR U14647 ( .A(n14591), .B(n14695), .Z(n14697) );
  XOR U14648 ( .A(n14706), .B(n14707), .Z(n14591) );
  AND U14649 ( .A(n307), .B(n14708), .Z(n14707) );
  XOR U14650 ( .A(n14709), .B(n14706), .Z(n14708) );
  XOR U14651 ( .A(n14710), .B(n14711), .Z(n14695) );
  AND U14652 ( .A(n14712), .B(n14713), .Z(n14711) );
  XNOR U14653 ( .A(n14710), .B(n14621), .Z(n14713) );
  XOR U14654 ( .A(n14714), .B(n14704), .Z(n14621) );
  XNOR U14655 ( .A(n14715), .B(n14699), .Z(n14704) );
  XOR U14656 ( .A(n14716), .B(n14717), .Z(n14699) );
  AND U14657 ( .A(n14718), .B(n14719), .Z(n14717) );
  XOR U14658 ( .A(n14720), .B(n14716), .Z(n14718) );
  XNOR U14659 ( .A(n14721), .B(n14722), .Z(n14715) );
  AND U14660 ( .A(n14723), .B(n14724), .Z(n14722) );
  XOR U14661 ( .A(n14721), .B(n14725), .Z(n14723) );
  XNOR U14662 ( .A(n14705), .B(n14702), .Z(n14714) );
  AND U14663 ( .A(n14726), .B(n14727), .Z(n14702) );
  XOR U14664 ( .A(n14728), .B(n14729), .Z(n14705) );
  AND U14665 ( .A(n14730), .B(n14731), .Z(n14729) );
  XOR U14666 ( .A(n14728), .B(n14732), .Z(n14730) );
  XNOR U14667 ( .A(n14618), .B(n14710), .Z(n14712) );
  XOR U14668 ( .A(n14733), .B(n14734), .Z(n14618) );
  AND U14669 ( .A(n307), .B(n14735), .Z(n14734) );
  XNOR U14670 ( .A(n14736), .B(n14733), .Z(n14735) );
  XOR U14671 ( .A(n14737), .B(n14738), .Z(n14710) );
  AND U14672 ( .A(n14739), .B(n14740), .Z(n14738) );
  XNOR U14673 ( .A(n14737), .B(n14726), .Z(n14740) );
  IV U14674 ( .A(n14671), .Z(n14726) );
  XNOR U14675 ( .A(n14741), .B(n14719), .Z(n14671) );
  XNOR U14676 ( .A(n14742), .B(n14725), .Z(n14719) );
  XNOR U14677 ( .A(n14743), .B(n14744), .Z(n14725) );
  NOR U14678 ( .A(n14745), .B(n14746), .Z(n14744) );
  XOR U14679 ( .A(n14743), .B(n14747), .Z(n14745) );
  XNOR U14680 ( .A(n14724), .B(n14716), .Z(n14742) );
  XOR U14681 ( .A(n14748), .B(n14749), .Z(n14716) );
  AND U14682 ( .A(n14750), .B(n14751), .Z(n14749) );
  XOR U14683 ( .A(n14748), .B(n14752), .Z(n14750) );
  XNOR U14684 ( .A(n14753), .B(n14721), .Z(n14724) );
  XOR U14685 ( .A(n14754), .B(n14755), .Z(n14721) );
  AND U14686 ( .A(n14756), .B(n14757), .Z(n14755) );
  XNOR U14687 ( .A(n14758), .B(n14759), .Z(n14756) );
  IV U14688 ( .A(n14754), .Z(n14758) );
  XNOR U14689 ( .A(n14760), .B(n14761), .Z(n14753) );
  NOR U14690 ( .A(n14762), .B(n14763), .Z(n14761) );
  XNOR U14691 ( .A(n14760), .B(n14764), .Z(n14762) );
  XNOR U14692 ( .A(n14720), .B(n14727), .Z(n14741) );
  NOR U14693 ( .A(n14684), .B(n14765), .Z(n14727) );
  XOR U14694 ( .A(n14732), .B(n14731), .Z(n14720) );
  XNOR U14695 ( .A(n14766), .B(n14728), .Z(n14731) );
  XOR U14696 ( .A(n14767), .B(n14768), .Z(n14728) );
  AND U14697 ( .A(n14769), .B(n14770), .Z(n14768) );
  XNOR U14698 ( .A(n14771), .B(n14772), .Z(n14769) );
  IV U14699 ( .A(n14767), .Z(n14771) );
  XNOR U14700 ( .A(n14773), .B(n14774), .Z(n14766) );
  NOR U14701 ( .A(n14775), .B(n14776), .Z(n14774) );
  XNOR U14702 ( .A(n14773), .B(n14777), .Z(n14775) );
  XOR U14703 ( .A(n14778), .B(n14779), .Z(n14732) );
  NOR U14704 ( .A(n14780), .B(n14781), .Z(n14779) );
  XNOR U14705 ( .A(n14778), .B(n14782), .Z(n14780) );
  XNOR U14706 ( .A(n14668), .B(n14737), .Z(n14739) );
  XOR U14707 ( .A(n14783), .B(n14784), .Z(n14668) );
  AND U14708 ( .A(n307), .B(n14785), .Z(n14784) );
  XOR U14709 ( .A(n14786), .B(n14783), .Z(n14785) );
  AND U14710 ( .A(n14681), .B(n14684), .Z(n14737) );
  XOR U14711 ( .A(n14787), .B(n14765), .Z(n14684) );
  XNOR U14712 ( .A(p_input[1200]), .B(p_input[2048]), .Z(n14765) );
  XNOR U14713 ( .A(n14752), .B(n14751), .Z(n14787) );
  XNOR U14714 ( .A(n14788), .B(n14759), .Z(n14751) );
  XNOR U14715 ( .A(n14747), .B(n14746), .Z(n14759) );
  XNOR U14716 ( .A(n14789), .B(n14743), .Z(n14746) );
  XNOR U14717 ( .A(p_input[1210]), .B(p_input[2058]), .Z(n14743) );
  XOR U14718 ( .A(p_input[1211]), .B(n6319), .Z(n14789) );
  XOR U14719 ( .A(p_input[1212]), .B(p_input[2060]), .Z(n14747) );
  XOR U14720 ( .A(n14757), .B(n14790), .Z(n14788) );
  IV U14721 ( .A(n14748), .Z(n14790) );
  XOR U14722 ( .A(p_input[1201]), .B(p_input[2049]), .Z(n14748) );
  XNOR U14723 ( .A(n14791), .B(n14764), .Z(n14757) );
  XNOR U14724 ( .A(p_input[1215]), .B(n6322), .Z(n14764) );
  XOR U14725 ( .A(n14754), .B(n14763), .Z(n14791) );
  XOR U14726 ( .A(n14792), .B(n14760), .Z(n14763) );
  XOR U14727 ( .A(p_input[1213]), .B(p_input[2061]), .Z(n14760) );
  XOR U14728 ( .A(p_input[1214]), .B(n6324), .Z(n14792) );
  XOR U14729 ( .A(p_input[1209]), .B(p_input[2057]), .Z(n14754) );
  XOR U14730 ( .A(n14772), .B(n14770), .Z(n14752) );
  XNOR U14731 ( .A(n14793), .B(n14777), .Z(n14770) );
  XOR U14732 ( .A(p_input[1208]), .B(p_input[2056]), .Z(n14777) );
  XOR U14733 ( .A(n14767), .B(n14776), .Z(n14793) );
  XOR U14734 ( .A(n14794), .B(n14773), .Z(n14776) );
  XOR U14735 ( .A(p_input[1206]), .B(p_input[2054]), .Z(n14773) );
  XOR U14736 ( .A(p_input[1207]), .B(n7007), .Z(n14794) );
  XOR U14737 ( .A(p_input[1202]), .B(p_input[2050]), .Z(n14767) );
  XNOR U14738 ( .A(n14782), .B(n14781), .Z(n14772) );
  XOR U14739 ( .A(n14795), .B(n14778), .Z(n14781) );
  XOR U14740 ( .A(p_input[1203]), .B(p_input[2051]), .Z(n14778) );
  XOR U14741 ( .A(p_input[1204]), .B(n7009), .Z(n14795) );
  XOR U14742 ( .A(p_input[1205]), .B(p_input[2053]), .Z(n14782) );
  XOR U14743 ( .A(n14796), .B(n14797), .Z(n14681) );
  AND U14744 ( .A(n307), .B(n14798), .Z(n14797) );
  XNOR U14745 ( .A(n14799), .B(n14796), .Z(n14798) );
  XNOR U14746 ( .A(n14800), .B(n14801), .Z(n307) );
  AND U14747 ( .A(n14802), .B(n14803), .Z(n14801) );
  XOR U14748 ( .A(n14694), .B(n14800), .Z(n14803) );
  AND U14749 ( .A(n14804), .B(n14805), .Z(n14694) );
  XNOR U14750 ( .A(n14691), .B(n14800), .Z(n14802) );
  XOR U14751 ( .A(n14806), .B(n14807), .Z(n14691) );
  AND U14752 ( .A(n311), .B(n14808), .Z(n14807) );
  XOR U14753 ( .A(n14809), .B(n14806), .Z(n14808) );
  XOR U14754 ( .A(n14810), .B(n14811), .Z(n14800) );
  AND U14755 ( .A(n14812), .B(n14813), .Z(n14811) );
  XNOR U14756 ( .A(n14810), .B(n14804), .Z(n14813) );
  IV U14757 ( .A(n14709), .Z(n14804) );
  XOR U14758 ( .A(n14814), .B(n14815), .Z(n14709) );
  XOR U14759 ( .A(n14816), .B(n14805), .Z(n14815) );
  AND U14760 ( .A(n14736), .B(n14817), .Z(n14805) );
  AND U14761 ( .A(n14818), .B(n14819), .Z(n14816) );
  XOR U14762 ( .A(n14820), .B(n14814), .Z(n14818) );
  XNOR U14763 ( .A(n14706), .B(n14810), .Z(n14812) );
  XOR U14764 ( .A(n14821), .B(n14822), .Z(n14706) );
  AND U14765 ( .A(n311), .B(n14823), .Z(n14822) );
  XOR U14766 ( .A(n14824), .B(n14821), .Z(n14823) );
  XOR U14767 ( .A(n14825), .B(n14826), .Z(n14810) );
  AND U14768 ( .A(n14827), .B(n14828), .Z(n14826) );
  XNOR U14769 ( .A(n14825), .B(n14736), .Z(n14828) );
  XOR U14770 ( .A(n14829), .B(n14819), .Z(n14736) );
  XNOR U14771 ( .A(n14830), .B(n14814), .Z(n14819) );
  XOR U14772 ( .A(n14831), .B(n14832), .Z(n14814) );
  AND U14773 ( .A(n14833), .B(n14834), .Z(n14832) );
  XOR U14774 ( .A(n14835), .B(n14831), .Z(n14833) );
  XNOR U14775 ( .A(n14836), .B(n14837), .Z(n14830) );
  AND U14776 ( .A(n14838), .B(n14839), .Z(n14837) );
  XOR U14777 ( .A(n14836), .B(n14840), .Z(n14838) );
  XNOR U14778 ( .A(n14820), .B(n14817), .Z(n14829) );
  AND U14779 ( .A(n14841), .B(n14842), .Z(n14817) );
  XOR U14780 ( .A(n14843), .B(n14844), .Z(n14820) );
  AND U14781 ( .A(n14845), .B(n14846), .Z(n14844) );
  XOR U14782 ( .A(n14843), .B(n14847), .Z(n14845) );
  XNOR U14783 ( .A(n14733), .B(n14825), .Z(n14827) );
  XOR U14784 ( .A(n14848), .B(n14849), .Z(n14733) );
  AND U14785 ( .A(n311), .B(n14850), .Z(n14849) );
  XNOR U14786 ( .A(n14851), .B(n14848), .Z(n14850) );
  XOR U14787 ( .A(n14852), .B(n14853), .Z(n14825) );
  AND U14788 ( .A(n14854), .B(n14855), .Z(n14853) );
  XNOR U14789 ( .A(n14852), .B(n14841), .Z(n14855) );
  IV U14790 ( .A(n14786), .Z(n14841) );
  XNOR U14791 ( .A(n14856), .B(n14834), .Z(n14786) );
  XNOR U14792 ( .A(n14857), .B(n14840), .Z(n14834) );
  XNOR U14793 ( .A(n14858), .B(n14859), .Z(n14840) );
  NOR U14794 ( .A(n14860), .B(n14861), .Z(n14859) );
  XOR U14795 ( .A(n14858), .B(n14862), .Z(n14860) );
  XNOR U14796 ( .A(n14839), .B(n14831), .Z(n14857) );
  XOR U14797 ( .A(n14863), .B(n14864), .Z(n14831) );
  AND U14798 ( .A(n14865), .B(n14866), .Z(n14864) );
  XOR U14799 ( .A(n14863), .B(n14867), .Z(n14865) );
  XNOR U14800 ( .A(n14868), .B(n14836), .Z(n14839) );
  XOR U14801 ( .A(n14869), .B(n14870), .Z(n14836) );
  AND U14802 ( .A(n14871), .B(n14872), .Z(n14870) );
  XNOR U14803 ( .A(n14873), .B(n14874), .Z(n14871) );
  IV U14804 ( .A(n14869), .Z(n14873) );
  XNOR U14805 ( .A(n14875), .B(n14876), .Z(n14868) );
  NOR U14806 ( .A(n14877), .B(n14878), .Z(n14876) );
  XNOR U14807 ( .A(n14875), .B(n14879), .Z(n14877) );
  XNOR U14808 ( .A(n14835), .B(n14842), .Z(n14856) );
  NOR U14809 ( .A(n14799), .B(n14880), .Z(n14842) );
  XOR U14810 ( .A(n14847), .B(n14846), .Z(n14835) );
  XNOR U14811 ( .A(n14881), .B(n14843), .Z(n14846) );
  XOR U14812 ( .A(n14882), .B(n14883), .Z(n14843) );
  AND U14813 ( .A(n14884), .B(n14885), .Z(n14883) );
  XNOR U14814 ( .A(n14886), .B(n14887), .Z(n14884) );
  IV U14815 ( .A(n14882), .Z(n14886) );
  XNOR U14816 ( .A(n14888), .B(n14889), .Z(n14881) );
  NOR U14817 ( .A(n14890), .B(n14891), .Z(n14889) );
  XNOR U14818 ( .A(n14888), .B(n14892), .Z(n14890) );
  XOR U14819 ( .A(n14893), .B(n14894), .Z(n14847) );
  NOR U14820 ( .A(n14895), .B(n14896), .Z(n14894) );
  XNOR U14821 ( .A(n14893), .B(n14897), .Z(n14895) );
  XNOR U14822 ( .A(n14783), .B(n14852), .Z(n14854) );
  XOR U14823 ( .A(n14898), .B(n14899), .Z(n14783) );
  AND U14824 ( .A(n311), .B(n14900), .Z(n14899) );
  XOR U14825 ( .A(n14901), .B(n14898), .Z(n14900) );
  AND U14826 ( .A(n14796), .B(n14799), .Z(n14852) );
  XOR U14827 ( .A(n14902), .B(n14880), .Z(n14799) );
  XNOR U14828 ( .A(p_input[1216]), .B(p_input[2048]), .Z(n14880) );
  XNOR U14829 ( .A(n14867), .B(n14866), .Z(n14902) );
  XNOR U14830 ( .A(n14903), .B(n14874), .Z(n14866) );
  XNOR U14831 ( .A(n14862), .B(n14861), .Z(n14874) );
  XNOR U14832 ( .A(n14904), .B(n14858), .Z(n14861) );
  XNOR U14833 ( .A(p_input[1226]), .B(p_input[2058]), .Z(n14858) );
  XOR U14834 ( .A(p_input[1227]), .B(n6319), .Z(n14904) );
  XOR U14835 ( .A(p_input[1228]), .B(p_input[2060]), .Z(n14862) );
  XOR U14836 ( .A(n14872), .B(n14905), .Z(n14903) );
  IV U14837 ( .A(n14863), .Z(n14905) );
  XOR U14838 ( .A(p_input[1217]), .B(p_input[2049]), .Z(n14863) );
  XNOR U14839 ( .A(n14906), .B(n14879), .Z(n14872) );
  XNOR U14840 ( .A(p_input[1231]), .B(n6322), .Z(n14879) );
  XOR U14841 ( .A(n14869), .B(n14878), .Z(n14906) );
  XOR U14842 ( .A(n14907), .B(n14875), .Z(n14878) );
  XOR U14843 ( .A(p_input[1229]), .B(p_input[2061]), .Z(n14875) );
  XOR U14844 ( .A(p_input[1230]), .B(n6324), .Z(n14907) );
  XOR U14845 ( .A(p_input[1225]), .B(p_input[2057]), .Z(n14869) );
  XOR U14846 ( .A(n14887), .B(n14885), .Z(n14867) );
  XNOR U14847 ( .A(n14908), .B(n14892), .Z(n14885) );
  XOR U14848 ( .A(p_input[1224]), .B(p_input[2056]), .Z(n14892) );
  XOR U14849 ( .A(n14882), .B(n14891), .Z(n14908) );
  XOR U14850 ( .A(n14909), .B(n14888), .Z(n14891) );
  XOR U14851 ( .A(p_input[1222]), .B(p_input[2054]), .Z(n14888) );
  XOR U14852 ( .A(p_input[1223]), .B(n7007), .Z(n14909) );
  XOR U14853 ( .A(p_input[1218]), .B(p_input[2050]), .Z(n14882) );
  XNOR U14854 ( .A(n14897), .B(n14896), .Z(n14887) );
  XOR U14855 ( .A(n14910), .B(n14893), .Z(n14896) );
  XOR U14856 ( .A(p_input[1219]), .B(p_input[2051]), .Z(n14893) );
  XOR U14857 ( .A(p_input[1220]), .B(n7009), .Z(n14910) );
  XOR U14858 ( .A(p_input[1221]), .B(p_input[2053]), .Z(n14897) );
  XOR U14859 ( .A(n14911), .B(n14912), .Z(n14796) );
  AND U14860 ( .A(n311), .B(n14913), .Z(n14912) );
  XNOR U14861 ( .A(n14914), .B(n14911), .Z(n14913) );
  XNOR U14862 ( .A(n14915), .B(n14916), .Z(n311) );
  AND U14863 ( .A(n14917), .B(n14918), .Z(n14916) );
  XOR U14864 ( .A(n14809), .B(n14915), .Z(n14918) );
  AND U14865 ( .A(n14919), .B(n14920), .Z(n14809) );
  XNOR U14866 ( .A(n14806), .B(n14915), .Z(n14917) );
  XOR U14867 ( .A(n14921), .B(n14922), .Z(n14806) );
  AND U14868 ( .A(n315), .B(n14923), .Z(n14922) );
  XOR U14869 ( .A(n14924), .B(n14921), .Z(n14923) );
  XOR U14870 ( .A(n14925), .B(n14926), .Z(n14915) );
  AND U14871 ( .A(n14927), .B(n14928), .Z(n14926) );
  XNOR U14872 ( .A(n14925), .B(n14919), .Z(n14928) );
  IV U14873 ( .A(n14824), .Z(n14919) );
  XOR U14874 ( .A(n14929), .B(n14930), .Z(n14824) );
  XOR U14875 ( .A(n14931), .B(n14920), .Z(n14930) );
  AND U14876 ( .A(n14851), .B(n14932), .Z(n14920) );
  AND U14877 ( .A(n14933), .B(n14934), .Z(n14931) );
  XOR U14878 ( .A(n14935), .B(n14929), .Z(n14933) );
  XNOR U14879 ( .A(n14821), .B(n14925), .Z(n14927) );
  XOR U14880 ( .A(n14936), .B(n14937), .Z(n14821) );
  AND U14881 ( .A(n315), .B(n14938), .Z(n14937) );
  XOR U14882 ( .A(n14939), .B(n14936), .Z(n14938) );
  XOR U14883 ( .A(n14940), .B(n14941), .Z(n14925) );
  AND U14884 ( .A(n14942), .B(n14943), .Z(n14941) );
  XNOR U14885 ( .A(n14940), .B(n14851), .Z(n14943) );
  XOR U14886 ( .A(n14944), .B(n14934), .Z(n14851) );
  XNOR U14887 ( .A(n14945), .B(n14929), .Z(n14934) );
  XOR U14888 ( .A(n14946), .B(n14947), .Z(n14929) );
  AND U14889 ( .A(n14948), .B(n14949), .Z(n14947) );
  XOR U14890 ( .A(n14950), .B(n14946), .Z(n14948) );
  XNOR U14891 ( .A(n14951), .B(n14952), .Z(n14945) );
  AND U14892 ( .A(n14953), .B(n14954), .Z(n14952) );
  XOR U14893 ( .A(n14951), .B(n14955), .Z(n14953) );
  XNOR U14894 ( .A(n14935), .B(n14932), .Z(n14944) );
  AND U14895 ( .A(n14956), .B(n14957), .Z(n14932) );
  XOR U14896 ( .A(n14958), .B(n14959), .Z(n14935) );
  AND U14897 ( .A(n14960), .B(n14961), .Z(n14959) );
  XOR U14898 ( .A(n14958), .B(n14962), .Z(n14960) );
  XNOR U14899 ( .A(n14848), .B(n14940), .Z(n14942) );
  XOR U14900 ( .A(n14963), .B(n14964), .Z(n14848) );
  AND U14901 ( .A(n315), .B(n14965), .Z(n14964) );
  XNOR U14902 ( .A(n14966), .B(n14963), .Z(n14965) );
  XOR U14903 ( .A(n14967), .B(n14968), .Z(n14940) );
  AND U14904 ( .A(n14969), .B(n14970), .Z(n14968) );
  XNOR U14905 ( .A(n14967), .B(n14956), .Z(n14970) );
  IV U14906 ( .A(n14901), .Z(n14956) );
  XNOR U14907 ( .A(n14971), .B(n14949), .Z(n14901) );
  XNOR U14908 ( .A(n14972), .B(n14955), .Z(n14949) );
  XNOR U14909 ( .A(n14973), .B(n14974), .Z(n14955) );
  NOR U14910 ( .A(n14975), .B(n14976), .Z(n14974) );
  XOR U14911 ( .A(n14973), .B(n14977), .Z(n14975) );
  XNOR U14912 ( .A(n14954), .B(n14946), .Z(n14972) );
  XOR U14913 ( .A(n14978), .B(n14979), .Z(n14946) );
  AND U14914 ( .A(n14980), .B(n14981), .Z(n14979) );
  XOR U14915 ( .A(n14978), .B(n14982), .Z(n14980) );
  XNOR U14916 ( .A(n14983), .B(n14951), .Z(n14954) );
  XOR U14917 ( .A(n14984), .B(n14985), .Z(n14951) );
  AND U14918 ( .A(n14986), .B(n14987), .Z(n14985) );
  XNOR U14919 ( .A(n14988), .B(n14989), .Z(n14986) );
  IV U14920 ( .A(n14984), .Z(n14988) );
  XNOR U14921 ( .A(n14990), .B(n14991), .Z(n14983) );
  NOR U14922 ( .A(n14992), .B(n14993), .Z(n14991) );
  XNOR U14923 ( .A(n14990), .B(n14994), .Z(n14992) );
  XNOR U14924 ( .A(n14950), .B(n14957), .Z(n14971) );
  NOR U14925 ( .A(n14914), .B(n14995), .Z(n14957) );
  XOR U14926 ( .A(n14962), .B(n14961), .Z(n14950) );
  XNOR U14927 ( .A(n14996), .B(n14958), .Z(n14961) );
  XOR U14928 ( .A(n14997), .B(n14998), .Z(n14958) );
  AND U14929 ( .A(n14999), .B(n15000), .Z(n14998) );
  XNOR U14930 ( .A(n15001), .B(n15002), .Z(n14999) );
  IV U14931 ( .A(n14997), .Z(n15001) );
  XNOR U14932 ( .A(n15003), .B(n15004), .Z(n14996) );
  NOR U14933 ( .A(n15005), .B(n15006), .Z(n15004) );
  XNOR U14934 ( .A(n15003), .B(n15007), .Z(n15005) );
  XOR U14935 ( .A(n15008), .B(n15009), .Z(n14962) );
  NOR U14936 ( .A(n15010), .B(n15011), .Z(n15009) );
  XNOR U14937 ( .A(n15008), .B(n15012), .Z(n15010) );
  XNOR U14938 ( .A(n14898), .B(n14967), .Z(n14969) );
  XOR U14939 ( .A(n15013), .B(n15014), .Z(n14898) );
  AND U14940 ( .A(n315), .B(n15015), .Z(n15014) );
  XOR U14941 ( .A(n15016), .B(n15013), .Z(n15015) );
  AND U14942 ( .A(n14911), .B(n14914), .Z(n14967) );
  XOR U14943 ( .A(n15017), .B(n14995), .Z(n14914) );
  XNOR U14944 ( .A(p_input[1232]), .B(p_input[2048]), .Z(n14995) );
  XNOR U14945 ( .A(n14982), .B(n14981), .Z(n15017) );
  XNOR U14946 ( .A(n15018), .B(n14989), .Z(n14981) );
  XNOR U14947 ( .A(n14977), .B(n14976), .Z(n14989) );
  XNOR U14948 ( .A(n15019), .B(n14973), .Z(n14976) );
  XNOR U14949 ( .A(p_input[1242]), .B(p_input[2058]), .Z(n14973) );
  XOR U14950 ( .A(p_input[1243]), .B(n6319), .Z(n15019) );
  XOR U14951 ( .A(p_input[1244]), .B(p_input[2060]), .Z(n14977) );
  XOR U14952 ( .A(n14987), .B(n15020), .Z(n15018) );
  IV U14953 ( .A(n14978), .Z(n15020) );
  XOR U14954 ( .A(p_input[1233]), .B(p_input[2049]), .Z(n14978) );
  XNOR U14955 ( .A(n15021), .B(n14994), .Z(n14987) );
  XNOR U14956 ( .A(p_input[1247]), .B(n6322), .Z(n14994) );
  XOR U14957 ( .A(n14984), .B(n14993), .Z(n15021) );
  XOR U14958 ( .A(n15022), .B(n14990), .Z(n14993) );
  XOR U14959 ( .A(p_input[1245]), .B(p_input[2061]), .Z(n14990) );
  XOR U14960 ( .A(p_input[1246]), .B(n6324), .Z(n15022) );
  XOR U14961 ( .A(p_input[1241]), .B(p_input[2057]), .Z(n14984) );
  XOR U14962 ( .A(n15002), .B(n15000), .Z(n14982) );
  XNOR U14963 ( .A(n15023), .B(n15007), .Z(n15000) );
  XOR U14964 ( .A(p_input[1240]), .B(p_input[2056]), .Z(n15007) );
  XOR U14965 ( .A(n14997), .B(n15006), .Z(n15023) );
  XOR U14966 ( .A(n15024), .B(n15003), .Z(n15006) );
  XOR U14967 ( .A(p_input[1238]), .B(p_input[2054]), .Z(n15003) );
  XOR U14968 ( .A(p_input[1239]), .B(n7007), .Z(n15024) );
  XOR U14969 ( .A(p_input[1234]), .B(p_input[2050]), .Z(n14997) );
  XNOR U14970 ( .A(n15012), .B(n15011), .Z(n15002) );
  XOR U14971 ( .A(n15025), .B(n15008), .Z(n15011) );
  XOR U14972 ( .A(p_input[1235]), .B(p_input[2051]), .Z(n15008) );
  XOR U14973 ( .A(p_input[1236]), .B(n7009), .Z(n15025) );
  XOR U14974 ( .A(p_input[1237]), .B(p_input[2053]), .Z(n15012) );
  XOR U14975 ( .A(n15026), .B(n15027), .Z(n14911) );
  AND U14976 ( .A(n315), .B(n15028), .Z(n15027) );
  XNOR U14977 ( .A(n15029), .B(n15026), .Z(n15028) );
  XNOR U14978 ( .A(n15030), .B(n15031), .Z(n315) );
  AND U14979 ( .A(n15032), .B(n15033), .Z(n15031) );
  XOR U14980 ( .A(n14924), .B(n15030), .Z(n15033) );
  AND U14981 ( .A(n15034), .B(n15035), .Z(n14924) );
  XNOR U14982 ( .A(n14921), .B(n15030), .Z(n15032) );
  XOR U14983 ( .A(n15036), .B(n15037), .Z(n14921) );
  AND U14984 ( .A(n319), .B(n15038), .Z(n15037) );
  XOR U14985 ( .A(n15039), .B(n15036), .Z(n15038) );
  XOR U14986 ( .A(n15040), .B(n15041), .Z(n15030) );
  AND U14987 ( .A(n15042), .B(n15043), .Z(n15041) );
  XNOR U14988 ( .A(n15040), .B(n15034), .Z(n15043) );
  IV U14989 ( .A(n14939), .Z(n15034) );
  XOR U14990 ( .A(n15044), .B(n15045), .Z(n14939) );
  XOR U14991 ( .A(n15046), .B(n15035), .Z(n15045) );
  AND U14992 ( .A(n14966), .B(n15047), .Z(n15035) );
  AND U14993 ( .A(n15048), .B(n15049), .Z(n15046) );
  XOR U14994 ( .A(n15050), .B(n15044), .Z(n15048) );
  XNOR U14995 ( .A(n14936), .B(n15040), .Z(n15042) );
  XOR U14996 ( .A(n15051), .B(n15052), .Z(n14936) );
  AND U14997 ( .A(n319), .B(n15053), .Z(n15052) );
  XOR U14998 ( .A(n15054), .B(n15051), .Z(n15053) );
  XOR U14999 ( .A(n15055), .B(n15056), .Z(n15040) );
  AND U15000 ( .A(n15057), .B(n15058), .Z(n15056) );
  XNOR U15001 ( .A(n15055), .B(n14966), .Z(n15058) );
  XOR U15002 ( .A(n15059), .B(n15049), .Z(n14966) );
  XNOR U15003 ( .A(n15060), .B(n15044), .Z(n15049) );
  XOR U15004 ( .A(n15061), .B(n15062), .Z(n15044) );
  AND U15005 ( .A(n15063), .B(n15064), .Z(n15062) );
  XOR U15006 ( .A(n15065), .B(n15061), .Z(n15063) );
  XNOR U15007 ( .A(n15066), .B(n15067), .Z(n15060) );
  AND U15008 ( .A(n15068), .B(n15069), .Z(n15067) );
  XOR U15009 ( .A(n15066), .B(n15070), .Z(n15068) );
  XNOR U15010 ( .A(n15050), .B(n15047), .Z(n15059) );
  AND U15011 ( .A(n15071), .B(n15072), .Z(n15047) );
  XOR U15012 ( .A(n15073), .B(n15074), .Z(n15050) );
  AND U15013 ( .A(n15075), .B(n15076), .Z(n15074) );
  XOR U15014 ( .A(n15073), .B(n15077), .Z(n15075) );
  XNOR U15015 ( .A(n14963), .B(n15055), .Z(n15057) );
  XOR U15016 ( .A(n15078), .B(n15079), .Z(n14963) );
  AND U15017 ( .A(n319), .B(n15080), .Z(n15079) );
  XNOR U15018 ( .A(n15081), .B(n15078), .Z(n15080) );
  XOR U15019 ( .A(n15082), .B(n15083), .Z(n15055) );
  AND U15020 ( .A(n15084), .B(n15085), .Z(n15083) );
  XNOR U15021 ( .A(n15082), .B(n15071), .Z(n15085) );
  IV U15022 ( .A(n15016), .Z(n15071) );
  XNOR U15023 ( .A(n15086), .B(n15064), .Z(n15016) );
  XNOR U15024 ( .A(n15087), .B(n15070), .Z(n15064) );
  XNOR U15025 ( .A(n15088), .B(n15089), .Z(n15070) );
  NOR U15026 ( .A(n15090), .B(n15091), .Z(n15089) );
  XOR U15027 ( .A(n15088), .B(n15092), .Z(n15090) );
  XNOR U15028 ( .A(n15069), .B(n15061), .Z(n15087) );
  XOR U15029 ( .A(n15093), .B(n15094), .Z(n15061) );
  AND U15030 ( .A(n15095), .B(n15096), .Z(n15094) );
  XOR U15031 ( .A(n15093), .B(n15097), .Z(n15095) );
  XNOR U15032 ( .A(n15098), .B(n15066), .Z(n15069) );
  XOR U15033 ( .A(n15099), .B(n15100), .Z(n15066) );
  AND U15034 ( .A(n15101), .B(n15102), .Z(n15100) );
  XNOR U15035 ( .A(n15103), .B(n15104), .Z(n15101) );
  IV U15036 ( .A(n15099), .Z(n15103) );
  XNOR U15037 ( .A(n15105), .B(n15106), .Z(n15098) );
  NOR U15038 ( .A(n15107), .B(n15108), .Z(n15106) );
  XNOR U15039 ( .A(n15105), .B(n15109), .Z(n15107) );
  XNOR U15040 ( .A(n15065), .B(n15072), .Z(n15086) );
  NOR U15041 ( .A(n15029), .B(n15110), .Z(n15072) );
  XOR U15042 ( .A(n15077), .B(n15076), .Z(n15065) );
  XNOR U15043 ( .A(n15111), .B(n15073), .Z(n15076) );
  XOR U15044 ( .A(n15112), .B(n15113), .Z(n15073) );
  AND U15045 ( .A(n15114), .B(n15115), .Z(n15113) );
  XNOR U15046 ( .A(n15116), .B(n15117), .Z(n15114) );
  IV U15047 ( .A(n15112), .Z(n15116) );
  XNOR U15048 ( .A(n15118), .B(n15119), .Z(n15111) );
  NOR U15049 ( .A(n15120), .B(n15121), .Z(n15119) );
  XNOR U15050 ( .A(n15118), .B(n15122), .Z(n15120) );
  XOR U15051 ( .A(n15123), .B(n15124), .Z(n15077) );
  NOR U15052 ( .A(n15125), .B(n15126), .Z(n15124) );
  XNOR U15053 ( .A(n15123), .B(n15127), .Z(n15125) );
  XNOR U15054 ( .A(n15013), .B(n15082), .Z(n15084) );
  XOR U15055 ( .A(n15128), .B(n15129), .Z(n15013) );
  AND U15056 ( .A(n319), .B(n15130), .Z(n15129) );
  XOR U15057 ( .A(n15131), .B(n15128), .Z(n15130) );
  AND U15058 ( .A(n15026), .B(n15029), .Z(n15082) );
  XOR U15059 ( .A(n15132), .B(n15110), .Z(n15029) );
  XNOR U15060 ( .A(p_input[1248]), .B(p_input[2048]), .Z(n15110) );
  XNOR U15061 ( .A(n15097), .B(n15096), .Z(n15132) );
  XNOR U15062 ( .A(n15133), .B(n15104), .Z(n15096) );
  XNOR U15063 ( .A(n15092), .B(n15091), .Z(n15104) );
  XNOR U15064 ( .A(n15134), .B(n15088), .Z(n15091) );
  XNOR U15065 ( .A(p_input[1258]), .B(p_input[2058]), .Z(n15088) );
  XOR U15066 ( .A(p_input[1259]), .B(n6319), .Z(n15134) );
  XOR U15067 ( .A(p_input[1260]), .B(p_input[2060]), .Z(n15092) );
  XOR U15068 ( .A(n15102), .B(n15135), .Z(n15133) );
  IV U15069 ( .A(n15093), .Z(n15135) );
  XOR U15070 ( .A(p_input[1249]), .B(p_input[2049]), .Z(n15093) );
  XNOR U15071 ( .A(n15136), .B(n15109), .Z(n15102) );
  XNOR U15072 ( .A(p_input[1263]), .B(n6322), .Z(n15109) );
  XOR U15073 ( .A(n15099), .B(n15108), .Z(n15136) );
  XOR U15074 ( .A(n15137), .B(n15105), .Z(n15108) );
  XOR U15075 ( .A(p_input[1261]), .B(p_input[2061]), .Z(n15105) );
  XOR U15076 ( .A(p_input[1262]), .B(n6324), .Z(n15137) );
  XOR U15077 ( .A(p_input[1257]), .B(p_input[2057]), .Z(n15099) );
  XOR U15078 ( .A(n15117), .B(n15115), .Z(n15097) );
  XNOR U15079 ( .A(n15138), .B(n15122), .Z(n15115) );
  XOR U15080 ( .A(p_input[1256]), .B(p_input[2056]), .Z(n15122) );
  XOR U15081 ( .A(n15112), .B(n15121), .Z(n15138) );
  XOR U15082 ( .A(n15139), .B(n15118), .Z(n15121) );
  XOR U15083 ( .A(p_input[1254]), .B(p_input[2054]), .Z(n15118) );
  XOR U15084 ( .A(p_input[1255]), .B(n7007), .Z(n15139) );
  XOR U15085 ( .A(p_input[1250]), .B(p_input[2050]), .Z(n15112) );
  XNOR U15086 ( .A(n15127), .B(n15126), .Z(n15117) );
  XOR U15087 ( .A(n15140), .B(n15123), .Z(n15126) );
  XOR U15088 ( .A(p_input[1251]), .B(p_input[2051]), .Z(n15123) );
  XOR U15089 ( .A(p_input[1252]), .B(n7009), .Z(n15140) );
  XOR U15090 ( .A(p_input[1253]), .B(p_input[2053]), .Z(n15127) );
  XOR U15091 ( .A(n15141), .B(n15142), .Z(n15026) );
  AND U15092 ( .A(n319), .B(n15143), .Z(n15142) );
  XNOR U15093 ( .A(n15144), .B(n15141), .Z(n15143) );
  XNOR U15094 ( .A(n15145), .B(n15146), .Z(n319) );
  AND U15095 ( .A(n15147), .B(n15148), .Z(n15146) );
  XOR U15096 ( .A(n15039), .B(n15145), .Z(n15148) );
  AND U15097 ( .A(n15149), .B(n15150), .Z(n15039) );
  XNOR U15098 ( .A(n15036), .B(n15145), .Z(n15147) );
  XOR U15099 ( .A(n15151), .B(n15152), .Z(n15036) );
  AND U15100 ( .A(n323), .B(n15153), .Z(n15152) );
  XOR U15101 ( .A(n15154), .B(n15151), .Z(n15153) );
  XOR U15102 ( .A(n15155), .B(n15156), .Z(n15145) );
  AND U15103 ( .A(n15157), .B(n15158), .Z(n15156) );
  XNOR U15104 ( .A(n15155), .B(n15149), .Z(n15158) );
  IV U15105 ( .A(n15054), .Z(n15149) );
  XOR U15106 ( .A(n15159), .B(n15160), .Z(n15054) );
  XOR U15107 ( .A(n15161), .B(n15150), .Z(n15160) );
  AND U15108 ( .A(n15081), .B(n15162), .Z(n15150) );
  AND U15109 ( .A(n15163), .B(n15164), .Z(n15161) );
  XOR U15110 ( .A(n15165), .B(n15159), .Z(n15163) );
  XNOR U15111 ( .A(n15051), .B(n15155), .Z(n15157) );
  XOR U15112 ( .A(n15166), .B(n15167), .Z(n15051) );
  AND U15113 ( .A(n323), .B(n15168), .Z(n15167) );
  XOR U15114 ( .A(n15169), .B(n15166), .Z(n15168) );
  XOR U15115 ( .A(n15170), .B(n15171), .Z(n15155) );
  AND U15116 ( .A(n15172), .B(n15173), .Z(n15171) );
  XNOR U15117 ( .A(n15170), .B(n15081), .Z(n15173) );
  XOR U15118 ( .A(n15174), .B(n15164), .Z(n15081) );
  XNOR U15119 ( .A(n15175), .B(n15159), .Z(n15164) );
  XOR U15120 ( .A(n15176), .B(n15177), .Z(n15159) );
  AND U15121 ( .A(n15178), .B(n15179), .Z(n15177) );
  XOR U15122 ( .A(n15180), .B(n15176), .Z(n15178) );
  XNOR U15123 ( .A(n15181), .B(n15182), .Z(n15175) );
  AND U15124 ( .A(n15183), .B(n15184), .Z(n15182) );
  XOR U15125 ( .A(n15181), .B(n15185), .Z(n15183) );
  XNOR U15126 ( .A(n15165), .B(n15162), .Z(n15174) );
  AND U15127 ( .A(n15186), .B(n15187), .Z(n15162) );
  XOR U15128 ( .A(n15188), .B(n15189), .Z(n15165) );
  AND U15129 ( .A(n15190), .B(n15191), .Z(n15189) );
  XOR U15130 ( .A(n15188), .B(n15192), .Z(n15190) );
  XNOR U15131 ( .A(n15078), .B(n15170), .Z(n15172) );
  XOR U15132 ( .A(n15193), .B(n15194), .Z(n15078) );
  AND U15133 ( .A(n323), .B(n15195), .Z(n15194) );
  XNOR U15134 ( .A(n15196), .B(n15193), .Z(n15195) );
  XOR U15135 ( .A(n15197), .B(n15198), .Z(n15170) );
  AND U15136 ( .A(n15199), .B(n15200), .Z(n15198) );
  XNOR U15137 ( .A(n15197), .B(n15186), .Z(n15200) );
  IV U15138 ( .A(n15131), .Z(n15186) );
  XNOR U15139 ( .A(n15201), .B(n15179), .Z(n15131) );
  XNOR U15140 ( .A(n15202), .B(n15185), .Z(n15179) );
  XNOR U15141 ( .A(n15203), .B(n15204), .Z(n15185) );
  NOR U15142 ( .A(n15205), .B(n15206), .Z(n15204) );
  XOR U15143 ( .A(n15203), .B(n15207), .Z(n15205) );
  XNOR U15144 ( .A(n15184), .B(n15176), .Z(n15202) );
  XOR U15145 ( .A(n15208), .B(n15209), .Z(n15176) );
  AND U15146 ( .A(n15210), .B(n15211), .Z(n15209) );
  XOR U15147 ( .A(n15208), .B(n15212), .Z(n15210) );
  XNOR U15148 ( .A(n15213), .B(n15181), .Z(n15184) );
  XOR U15149 ( .A(n15214), .B(n15215), .Z(n15181) );
  AND U15150 ( .A(n15216), .B(n15217), .Z(n15215) );
  XNOR U15151 ( .A(n15218), .B(n15219), .Z(n15216) );
  IV U15152 ( .A(n15214), .Z(n15218) );
  XNOR U15153 ( .A(n15220), .B(n15221), .Z(n15213) );
  NOR U15154 ( .A(n15222), .B(n15223), .Z(n15221) );
  XNOR U15155 ( .A(n15220), .B(n15224), .Z(n15222) );
  XNOR U15156 ( .A(n15180), .B(n15187), .Z(n15201) );
  NOR U15157 ( .A(n15144), .B(n15225), .Z(n15187) );
  XOR U15158 ( .A(n15192), .B(n15191), .Z(n15180) );
  XNOR U15159 ( .A(n15226), .B(n15188), .Z(n15191) );
  XOR U15160 ( .A(n15227), .B(n15228), .Z(n15188) );
  AND U15161 ( .A(n15229), .B(n15230), .Z(n15228) );
  XNOR U15162 ( .A(n15231), .B(n15232), .Z(n15229) );
  IV U15163 ( .A(n15227), .Z(n15231) );
  XNOR U15164 ( .A(n15233), .B(n15234), .Z(n15226) );
  NOR U15165 ( .A(n15235), .B(n15236), .Z(n15234) );
  XNOR U15166 ( .A(n15233), .B(n15237), .Z(n15235) );
  XOR U15167 ( .A(n15238), .B(n15239), .Z(n15192) );
  NOR U15168 ( .A(n15240), .B(n15241), .Z(n15239) );
  XNOR U15169 ( .A(n15238), .B(n15242), .Z(n15240) );
  XNOR U15170 ( .A(n15128), .B(n15197), .Z(n15199) );
  XOR U15171 ( .A(n15243), .B(n15244), .Z(n15128) );
  AND U15172 ( .A(n323), .B(n15245), .Z(n15244) );
  XOR U15173 ( .A(n15246), .B(n15243), .Z(n15245) );
  AND U15174 ( .A(n15141), .B(n15144), .Z(n15197) );
  XOR U15175 ( .A(n15247), .B(n15225), .Z(n15144) );
  XNOR U15176 ( .A(p_input[1264]), .B(p_input[2048]), .Z(n15225) );
  XNOR U15177 ( .A(n15212), .B(n15211), .Z(n15247) );
  XNOR U15178 ( .A(n15248), .B(n15219), .Z(n15211) );
  XNOR U15179 ( .A(n15207), .B(n15206), .Z(n15219) );
  XNOR U15180 ( .A(n15249), .B(n15203), .Z(n15206) );
  XNOR U15181 ( .A(p_input[1274]), .B(p_input[2058]), .Z(n15203) );
  XOR U15182 ( .A(p_input[1275]), .B(n6319), .Z(n15249) );
  XOR U15183 ( .A(p_input[1276]), .B(p_input[2060]), .Z(n15207) );
  XOR U15184 ( .A(n15217), .B(n15250), .Z(n15248) );
  IV U15185 ( .A(n15208), .Z(n15250) );
  XOR U15186 ( .A(p_input[1265]), .B(p_input[2049]), .Z(n15208) );
  XNOR U15187 ( .A(n15251), .B(n15224), .Z(n15217) );
  XNOR U15188 ( .A(p_input[1279]), .B(n6322), .Z(n15224) );
  XOR U15189 ( .A(n15214), .B(n15223), .Z(n15251) );
  XOR U15190 ( .A(n15252), .B(n15220), .Z(n15223) );
  XOR U15191 ( .A(p_input[1277]), .B(p_input[2061]), .Z(n15220) );
  XOR U15192 ( .A(p_input[1278]), .B(n6324), .Z(n15252) );
  XOR U15193 ( .A(p_input[1273]), .B(p_input[2057]), .Z(n15214) );
  XOR U15194 ( .A(n15232), .B(n15230), .Z(n15212) );
  XNOR U15195 ( .A(n15253), .B(n15237), .Z(n15230) );
  XOR U15196 ( .A(p_input[1272]), .B(p_input[2056]), .Z(n15237) );
  XOR U15197 ( .A(n15227), .B(n15236), .Z(n15253) );
  XOR U15198 ( .A(n15254), .B(n15233), .Z(n15236) );
  XOR U15199 ( .A(p_input[1270]), .B(p_input[2054]), .Z(n15233) );
  XOR U15200 ( .A(p_input[1271]), .B(n7007), .Z(n15254) );
  XOR U15201 ( .A(p_input[1266]), .B(p_input[2050]), .Z(n15227) );
  XNOR U15202 ( .A(n15242), .B(n15241), .Z(n15232) );
  XOR U15203 ( .A(n15255), .B(n15238), .Z(n15241) );
  XOR U15204 ( .A(p_input[1267]), .B(p_input[2051]), .Z(n15238) );
  XOR U15205 ( .A(p_input[1268]), .B(n7009), .Z(n15255) );
  XOR U15206 ( .A(p_input[1269]), .B(p_input[2053]), .Z(n15242) );
  XOR U15207 ( .A(n15256), .B(n15257), .Z(n15141) );
  AND U15208 ( .A(n323), .B(n15258), .Z(n15257) );
  XNOR U15209 ( .A(n15259), .B(n15256), .Z(n15258) );
  XNOR U15210 ( .A(n15260), .B(n15261), .Z(n323) );
  AND U15211 ( .A(n15262), .B(n15263), .Z(n15261) );
  XOR U15212 ( .A(n15154), .B(n15260), .Z(n15263) );
  AND U15213 ( .A(n15264), .B(n15265), .Z(n15154) );
  XNOR U15214 ( .A(n15151), .B(n15260), .Z(n15262) );
  XOR U15215 ( .A(n15266), .B(n15267), .Z(n15151) );
  AND U15216 ( .A(n327), .B(n15268), .Z(n15267) );
  XOR U15217 ( .A(n15269), .B(n15266), .Z(n15268) );
  XOR U15218 ( .A(n15270), .B(n15271), .Z(n15260) );
  AND U15219 ( .A(n15272), .B(n15273), .Z(n15271) );
  XNOR U15220 ( .A(n15270), .B(n15264), .Z(n15273) );
  IV U15221 ( .A(n15169), .Z(n15264) );
  XOR U15222 ( .A(n15274), .B(n15275), .Z(n15169) );
  XOR U15223 ( .A(n15276), .B(n15265), .Z(n15275) );
  AND U15224 ( .A(n15196), .B(n15277), .Z(n15265) );
  AND U15225 ( .A(n15278), .B(n15279), .Z(n15276) );
  XOR U15226 ( .A(n15280), .B(n15274), .Z(n15278) );
  XNOR U15227 ( .A(n15166), .B(n15270), .Z(n15272) );
  XOR U15228 ( .A(n15281), .B(n15282), .Z(n15166) );
  AND U15229 ( .A(n327), .B(n15283), .Z(n15282) );
  XOR U15230 ( .A(n15284), .B(n15281), .Z(n15283) );
  XOR U15231 ( .A(n15285), .B(n15286), .Z(n15270) );
  AND U15232 ( .A(n15287), .B(n15288), .Z(n15286) );
  XNOR U15233 ( .A(n15285), .B(n15196), .Z(n15288) );
  XOR U15234 ( .A(n15289), .B(n15279), .Z(n15196) );
  XNOR U15235 ( .A(n15290), .B(n15274), .Z(n15279) );
  XOR U15236 ( .A(n15291), .B(n15292), .Z(n15274) );
  AND U15237 ( .A(n15293), .B(n15294), .Z(n15292) );
  XOR U15238 ( .A(n15295), .B(n15291), .Z(n15293) );
  XNOR U15239 ( .A(n15296), .B(n15297), .Z(n15290) );
  AND U15240 ( .A(n15298), .B(n15299), .Z(n15297) );
  XOR U15241 ( .A(n15296), .B(n15300), .Z(n15298) );
  XNOR U15242 ( .A(n15280), .B(n15277), .Z(n15289) );
  AND U15243 ( .A(n15301), .B(n15302), .Z(n15277) );
  XOR U15244 ( .A(n15303), .B(n15304), .Z(n15280) );
  AND U15245 ( .A(n15305), .B(n15306), .Z(n15304) );
  XOR U15246 ( .A(n15303), .B(n15307), .Z(n15305) );
  XNOR U15247 ( .A(n15193), .B(n15285), .Z(n15287) );
  XOR U15248 ( .A(n15308), .B(n15309), .Z(n15193) );
  AND U15249 ( .A(n327), .B(n15310), .Z(n15309) );
  XNOR U15250 ( .A(n15311), .B(n15308), .Z(n15310) );
  XOR U15251 ( .A(n15312), .B(n15313), .Z(n15285) );
  AND U15252 ( .A(n15314), .B(n15315), .Z(n15313) );
  XNOR U15253 ( .A(n15312), .B(n15301), .Z(n15315) );
  IV U15254 ( .A(n15246), .Z(n15301) );
  XNOR U15255 ( .A(n15316), .B(n15294), .Z(n15246) );
  XNOR U15256 ( .A(n15317), .B(n15300), .Z(n15294) );
  XNOR U15257 ( .A(n15318), .B(n15319), .Z(n15300) );
  NOR U15258 ( .A(n15320), .B(n15321), .Z(n15319) );
  XOR U15259 ( .A(n15318), .B(n15322), .Z(n15320) );
  XNOR U15260 ( .A(n15299), .B(n15291), .Z(n15317) );
  XOR U15261 ( .A(n15323), .B(n15324), .Z(n15291) );
  AND U15262 ( .A(n15325), .B(n15326), .Z(n15324) );
  XOR U15263 ( .A(n15323), .B(n15327), .Z(n15325) );
  XNOR U15264 ( .A(n15328), .B(n15296), .Z(n15299) );
  XOR U15265 ( .A(n15329), .B(n15330), .Z(n15296) );
  AND U15266 ( .A(n15331), .B(n15332), .Z(n15330) );
  XNOR U15267 ( .A(n15333), .B(n15334), .Z(n15331) );
  IV U15268 ( .A(n15329), .Z(n15333) );
  XNOR U15269 ( .A(n15335), .B(n15336), .Z(n15328) );
  NOR U15270 ( .A(n15337), .B(n15338), .Z(n15336) );
  XNOR U15271 ( .A(n15335), .B(n15339), .Z(n15337) );
  XNOR U15272 ( .A(n15295), .B(n15302), .Z(n15316) );
  NOR U15273 ( .A(n15259), .B(n15340), .Z(n15302) );
  XOR U15274 ( .A(n15307), .B(n15306), .Z(n15295) );
  XNOR U15275 ( .A(n15341), .B(n15303), .Z(n15306) );
  XOR U15276 ( .A(n15342), .B(n15343), .Z(n15303) );
  AND U15277 ( .A(n15344), .B(n15345), .Z(n15343) );
  XNOR U15278 ( .A(n15346), .B(n15347), .Z(n15344) );
  IV U15279 ( .A(n15342), .Z(n15346) );
  XNOR U15280 ( .A(n15348), .B(n15349), .Z(n15341) );
  NOR U15281 ( .A(n15350), .B(n15351), .Z(n15349) );
  XNOR U15282 ( .A(n15348), .B(n15352), .Z(n15350) );
  XOR U15283 ( .A(n15353), .B(n15354), .Z(n15307) );
  NOR U15284 ( .A(n15355), .B(n15356), .Z(n15354) );
  XNOR U15285 ( .A(n15353), .B(n15357), .Z(n15355) );
  XNOR U15286 ( .A(n15243), .B(n15312), .Z(n15314) );
  XOR U15287 ( .A(n15358), .B(n15359), .Z(n15243) );
  AND U15288 ( .A(n327), .B(n15360), .Z(n15359) );
  XOR U15289 ( .A(n15361), .B(n15358), .Z(n15360) );
  AND U15290 ( .A(n15256), .B(n15259), .Z(n15312) );
  XOR U15291 ( .A(n15362), .B(n15340), .Z(n15259) );
  XNOR U15292 ( .A(p_input[1280]), .B(p_input[2048]), .Z(n15340) );
  XNOR U15293 ( .A(n15327), .B(n15326), .Z(n15362) );
  XNOR U15294 ( .A(n15363), .B(n15334), .Z(n15326) );
  XNOR U15295 ( .A(n15322), .B(n15321), .Z(n15334) );
  XNOR U15296 ( .A(n15364), .B(n15318), .Z(n15321) );
  XNOR U15297 ( .A(p_input[1290]), .B(p_input[2058]), .Z(n15318) );
  XOR U15298 ( .A(p_input[1291]), .B(n6319), .Z(n15364) );
  XOR U15299 ( .A(p_input[1292]), .B(p_input[2060]), .Z(n15322) );
  XOR U15300 ( .A(n15332), .B(n15365), .Z(n15363) );
  IV U15301 ( .A(n15323), .Z(n15365) );
  XOR U15302 ( .A(p_input[1281]), .B(p_input[2049]), .Z(n15323) );
  XNOR U15303 ( .A(n15366), .B(n15339), .Z(n15332) );
  XNOR U15304 ( .A(p_input[1295]), .B(n6322), .Z(n15339) );
  XOR U15305 ( .A(n15329), .B(n15338), .Z(n15366) );
  XOR U15306 ( .A(n15367), .B(n15335), .Z(n15338) );
  XOR U15307 ( .A(p_input[1293]), .B(p_input[2061]), .Z(n15335) );
  XOR U15308 ( .A(p_input[1294]), .B(n6324), .Z(n15367) );
  XOR U15309 ( .A(p_input[1289]), .B(p_input[2057]), .Z(n15329) );
  XOR U15310 ( .A(n15347), .B(n15345), .Z(n15327) );
  XNOR U15311 ( .A(n15368), .B(n15352), .Z(n15345) );
  XOR U15312 ( .A(p_input[1288]), .B(p_input[2056]), .Z(n15352) );
  XOR U15313 ( .A(n15342), .B(n15351), .Z(n15368) );
  XOR U15314 ( .A(n15369), .B(n15348), .Z(n15351) );
  XOR U15315 ( .A(p_input[1286]), .B(p_input[2054]), .Z(n15348) );
  XOR U15316 ( .A(p_input[1287]), .B(n7007), .Z(n15369) );
  XOR U15317 ( .A(p_input[1282]), .B(p_input[2050]), .Z(n15342) );
  XNOR U15318 ( .A(n15357), .B(n15356), .Z(n15347) );
  XOR U15319 ( .A(n15370), .B(n15353), .Z(n15356) );
  XOR U15320 ( .A(p_input[1283]), .B(p_input[2051]), .Z(n15353) );
  XOR U15321 ( .A(p_input[1284]), .B(n7009), .Z(n15370) );
  XOR U15322 ( .A(p_input[1285]), .B(p_input[2053]), .Z(n15357) );
  XOR U15323 ( .A(n15371), .B(n15372), .Z(n15256) );
  AND U15324 ( .A(n327), .B(n15373), .Z(n15372) );
  XNOR U15325 ( .A(n15374), .B(n15371), .Z(n15373) );
  XNOR U15326 ( .A(n15375), .B(n15376), .Z(n327) );
  AND U15327 ( .A(n15377), .B(n15378), .Z(n15376) );
  XOR U15328 ( .A(n15269), .B(n15375), .Z(n15378) );
  AND U15329 ( .A(n15379), .B(n15380), .Z(n15269) );
  XNOR U15330 ( .A(n15266), .B(n15375), .Z(n15377) );
  XOR U15331 ( .A(n15381), .B(n15382), .Z(n15266) );
  AND U15332 ( .A(n331), .B(n15383), .Z(n15382) );
  XOR U15333 ( .A(n15384), .B(n15381), .Z(n15383) );
  XOR U15334 ( .A(n15385), .B(n15386), .Z(n15375) );
  AND U15335 ( .A(n15387), .B(n15388), .Z(n15386) );
  XNOR U15336 ( .A(n15385), .B(n15379), .Z(n15388) );
  IV U15337 ( .A(n15284), .Z(n15379) );
  XOR U15338 ( .A(n15389), .B(n15390), .Z(n15284) );
  XOR U15339 ( .A(n15391), .B(n15380), .Z(n15390) );
  AND U15340 ( .A(n15311), .B(n15392), .Z(n15380) );
  AND U15341 ( .A(n15393), .B(n15394), .Z(n15391) );
  XOR U15342 ( .A(n15395), .B(n15389), .Z(n15393) );
  XNOR U15343 ( .A(n15281), .B(n15385), .Z(n15387) );
  XOR U15344 ( .A(n15396), .B(n15397), .Z(n15281) );
  AND U15345 ( .A(n331), .B(n15398), .Z(n15397) );
  XOR U15346 ( .A(n15399), .B(n15396), .Z(n15398) );
  XOR U15347 ( .A(n15400), .B(n15401), .Z(n15385) );
  AND U15348 ( .A(n15402), .B(n15403), .Z(n15401) );
  XNOR U15349 ( .A(n15400), .B(n15311), .Z(n15403) );
  XOR U15350 ( .A(n15404), .B(n15394), .Z(n15311) );
  XNOR U15351 ( .A(n15405), .B(n15389), .Z(n15394) );
  XOR U15352 ( .A(n15406), .B(n15407), .Z(n15389) );
  AND U15353 ( .A(n15408), .B(n15409), .Z(n15407) );
  XOR U15354 ( .A(n15410), .B(n15406), .Z(n15408) );
  XNOR U15355 ( .A(n15411), .B(n15412), .Z(n15405) );
  AND U15356 ( .A(n15413), .B(n15414), .Z(n15412) );
  XOR U15357 ( .A(n15411), .B(n15415), .Z(n15413) );
  XNOR U15358 ( .A(n15395), .B(n15392), .Z(n15404) );
  AND U15359 ( .A(n15416), .B(n15417), .Z(n15392) );
  XOR U15360 ( .A(n15418), .B(n15419), .Z(n15395) );
  AND U15361 ( .A(n15420), .B(n15421), .Z(n15419) );
  XOR U15362 ( .A(n15418), .B(n15422), .Z(n15420) );
  XNOR U15363 ( .A(n15308), .B(n15400), .Z(n15402) );
  XOR U15364 ( .A(n15423), .B(n15424), .Z(n15308) );
  AND U15365 ( .A(n331), .B(n15425), .Z(n15424) );
  XNOR U15366 ( .A(n15426), .B(n15423), .Z(n15425) );
  XOR U15367 ( .A(n15427), .B(n15428), .Z(n15400) );
  AND U15368 ( .A(n15429), .B(n15430), .Z(n15428) );
  XNOR U15369 ( .A(n15427), .B(n15416), .Z(n15430) );
  IV U15370 ( .A(n15361), .Z(n15416) );
  XNOR U15371 ( .A(n15431), .B(n15409), .Z(n15361) );
  XNOR U15372 ( .A(n15432), .B(n15415), .Z(n15409) );
  XNOR U15373 ( .A(n15433), .B(n15434), .Z(n15415) );
  NOR U15374 ( .A(n15435), .B(n15436), .Z(n15434) );
  XOR U15375 ( .A(n15433), .B(n15437), .Z(n15435) );
  XNOR U15376 ( .A(n15414), .B(n15406), .Z(n15432) );
  XOR U15377 ( .A(n15438), .B(n15439), .Z(n15406) );
  AND U15378 ( .A(n15440), .B(n15441), .Z(n15439) );
  XOR U15379 ( .A(n15438), .B(n15442), .Z(n15440) );
  XNOR U15380 ( .A(n15443), .B(n15411), .Z(n15414) );
  XOR U15381 ( .A(n15444), .B(n15445), .Z(n15411) );
  AND U15382 ( .A(n15446), .B(n15447), .Z(n15445) );
  XNOR U15383 ( .A(n15448), .B(n15449), .Z(n15446) );
  IV U15384 ( .A(n15444), .Z(n15448) );
  XNOR U15385 ( .A(n15450), .B(n15451), .Z(n15443) );
  NOR U15386 ( .A(n15452), .B(n15453), .Z(n15451) );
  XNOR U15387 ( .A(n15450), .B(n15454), .Z(n15452) );
  XNOR U15388 ( .A(n15410), .B(n15417), .Z(n15431) );
  NOR U15389 ( .A(n15374), .B(n15455), .Z(n15417) );
  XOR U15390 ( .A(n15422), .B(n15421), .Z(n15410) );
  XNOR U15391 ( .A(n15456), .B(n15418), .Z(n15421) );
  XOR U15392 ( .A(n15457), .B(n15458), .Z(n15418) );
  AND U15393 ( .A(n15459), .B(n15460), .Z(n15458) );
  XNOR U15394 ( .A(n15461), .B(n15462), .Z(n15459) );
  IV U15395 ( .A(n15457), .Z(n15461) );
  XNOR U15396 ( .A(n15463), .B(n15464), .Z(n15456) );
  NOR U15397 ( .A(n15465), .B(n15466), .Z(n15464) );
  XNOR U15398 ( .A(n15463), .B(n15467), .Z(n15465) );
  XOR U15399 ( .A(n15468), .B(n15469), .Z(n15422) );
  NOR U15400 ( .A(n15470), .B(n15471), .Z(n15469) );
  XNOR U15401 ( .A(n15468), .B(n15472), .Z(n15470) );
  XNOR U15402 ( .A(n15358), .B(n15427), .Z(n15429) );
  XOR U15403 ( .A(n15473), .B(n15474), .Z(n15358) );
  AND U15404 ( .A(n331), .B(n15475), .Z(n15474) );
  XOR U15405 ( .A(n15476), .B(n15473), .Z(n15475) );
  AND U15406 ( .A(n15371), .B(n15374), .Z(n15427) );
  XOR U15407 ( .A(n15477), .B(n15455), .Z(n15374) );
  XNOR U15408 ( .A(p_input[1296]), .B(p_input[2048]), .Z(n15455) );
  XNOR U15409 ( .A(n15442), .B(n15441), .Z(n15477) );
  XNOR U15410 ( .A(n15478), .B(n15449), .Z(n15441) );
  XNOR U15411 ( .A(n15437), .B(n15436), .Z(n15449) );
  XNOR U15412 ( .A(n15479), .B(n15433), .Z(n15436) );
  XNOR U15413 ( .A(p_input[1306]), .B(p_input[2058]), .Z(n15433) );
  XOR U15414 ( .A(p_input[1307]), .B(n6319), .Z(n15479) );
  XOR U15415 ( .A(p_input[1308]), .B(p_input[2060]), .Z(n15437) );
  XOR U15416 ( .A(n15447), .B(n15480), .Z(n15478) );
  IV U15417 ( .A(n15438), .Z(n15480) );
  XOR U15418 ( .A(p_input[1297]), .B(p_input[2049]), .Z(n15438) );
  XNOR U15419 ( .A(n15481), .B(n15454), .Z(n15447) );
  XNOR U15420 ( .A(p_input[1311]), .B(n6322), .Z(n15454) );
  XOR U15421 ( .A(n15444), .B(n15453), .Z(n15481) );
  XOR U15422 ( .A(n15482), .B(n15450), .Z(n15453) );
  XOR U15423 ( .A(p_input[1309]), .B(p_input[2061]), .Z(n15450) );
  XOR U15424 ( .A(p_input[1310]), .B(n6324), .Z(n15482) );
  XOR U15425 ( .A(p_input[1305]), .B(p_input[2057]), .Z(n15444) );
  XOR U15426 ( .A(n15462), .B(n15460), .Z(n15442) );
  XNOR U15427 ( .A(n15483), .B(n15467), .Z(n15460) );
  XOR U15428 ( .A(p_input[1304]), .B(p_input[2056]), .Z(n15467) );
  XOR U15429 ( .A(n15457), .B(n15466), .Z(n15483) );
  XOR U15430 ( .A(n15484), .B(n15463), .Z(n15466) );
  XOR U15431 ( .A(p_input[1302]), .B(p_input[2054]), .Z(n15463) );
  XOR U15432 ( .A(p_input[1303]), .B(n7007), .Z(n15484) );
  XOR U15433 ( .A(p_input[1298]), .B(p_input[2050]), .Z(n15457) );
  XNOR U15434 ( .A(n15472), .B(n15471), .Z(n15462) );
  XOR U15435 ( .A(n15485), .B(n15468), .Z(n15471) );
  XOR U15436 ( .A(p_input[1299]), .B(p_input[2051]), .Z(n15468) );
  XOR U15437 ( .A(p_input[1300]), .B(n7009), .Z(n15485) );
  XOR U15438 ( .A(p_input[1301]), .B(p_input[2053]), .Z(n15472) );
  XOR U15439 ( .A(n15486), .B(n15487), .Z(n15371) );
  AND U15440 ( .A(n331), .B(n15488), .Z(n15487) );
  XNOR U15441 ( .A(n15489), .B(n15486), .Z(n15488) );
  XNOR U15442 ( .A(n15490), .B(n15491), .Z(n331) );
  AND U15443 ( .A(n15492), .B(n15493), .Z(n15491) );
  XOR U15444 ( .A(n15384), .B(n15490), .Z(n15493) );
  AND U15445 ( .A(n15494), .B(n15495), .Z(n15384) );
  XNOR U15446 ( .A(n15381), .B(n15490), .Z(n15492) );
  XOR U15447 ( .A(n15496), .B(n15497), .Z(n15381) );
  AND U15448 ( .A(n335), .B(n15498), .Z(n15497) );
  XOR U15449 ( .A(n15499), .B(n15496), .Z(n15498) );
  XOR U15450 ( .A(n15500), .B(n15501), .Z(n15490) );
  AND U15451 ( .A(n15502), .B(n15503), .Z(n15501) );
  XNOR U15452 ( .A(n15500), .B(n15494), .Z(n15503) );
  IV U15453 ( .A(n15399), .Z(n15494) );
  XOR U15454 ( .A(n15504), .B(n15505), .Z(n15399) );
  XOR U15455 ( .A(n15506), .B(n15495), .Z(n15505) );
  AND U15456 ( .A(n15426), .B(n15507), .Z(n15495) );
  AND U15457 ( .A(n15508), .B(n15509), .Z(n15506) );
  XOR U15458 ( .A(n15510), .B(n15504), .Z(n15508) );
  XNOR U15459 ( .A(n15396), .B(n15500), .Z(n15502) );
  XOR U15460 ( .A(n15511), .B(n15512), .Z(n15396) );
  AND U15461 ( .A(n335), .B(n15513), .Z(n15512) );
  XOR U15462 ( .A(n15514), .B(n15511), .Z(n15513) );
  XOR U15463 ( .A(n15515), .B(n15516), .Z(n15500) );
  AND U15464 ( .A(n15517), .B(n15518), .Z(n15516) );
  XNOR U15465 ( .A(n15515), .B(n15426), .Z(n15518) );
  XOR U15466 ( .A(n15519), .B(n15509), .Z(n15426) );
  XNOR U15467 ( .A(n15520), .B(n15504), .Z(n15509) );
  XOR U15468 ( .A(n15521), .B(n15522), .Z(n15504) );
  AND U15469 ( .A(n15523), .B(n15524), .Z(n15522) );
  XOR U15470 ( .A(n15525), .B(n15521), .Z(n15523) );
  XNOR U15471 ( .A(n15526), .B(n15527), .Z(n15520) );
  AND U15472 ( .A(n15528), .B(n15529), .Z(n15527) );
  XOR U15473 ( .A(n15526), .B(n15530), .Z(n15528) );
  XNOR U15474 ( .A(n15510), .B(n15507), .Z(n15519) );
  AND U15475 ( .A(n15531), .B(n15532), .Z(n15507) );
  XOR U15476 ( .A(n15533), .B(n15534), .Z(n15510) );
  AND U15477 ( .A(n15535), .B(n15536), .Z(n15534) );
  XOR U15478 ( .A(n15533), .B(n15537), .Z(n15535) );
  XNOR U15479 ( .A(n15423), .B(n15515), .Z(n15517) );
  XOR U15480 ( .A(n15538), .B(n15539), .Z(n15423) );
  AND U15481 ( .A(n335), .B(n15540), .Z(n15539) );
  XNOR U15482 ( .A(n15541), .B(n15538), .Z(n15540) );
  XOR U15483 ( .A(n15542), .B(n15543), .Z(n15515) );
  AND U15484 ( .A(n15544), .B(n15545), .Z(n15543) );
  XNOR U15485 ( .A(n15542), .B(n15531), .Z(n15545) );
  IV U15486 ( .A(n15476), .Z(n15531) );
  XNOR U15487 ( .A(n15546), .B(n15524), .Z(n15476) );
  XNOR U15488 ( .A(n15547), .B(n15530), .Z(n15524) );
  XNOR U15489 ( .A(n15548), .B(n15549), .Z(n15530) );
  NOR U15490 ( .A(n15550), .B(n15551), .Z(n15549) );
  XOR U15491 ( .A(n15548), .B(n15552), .Z(n15550) );
  XNOR U15492 ( .A(n15529), .B(n15521), .Z(n15547) );
  XOR U15493 ( .A(n15553), .B(n15554), .Z(n15521) );
  AND U15494 ( .A(n15555), .B(n15556), .Z(n15554) );
  XOR U15495 ( .A(n15553), .B(n15557), .Z(n15555) );
  XNOR U15496 ( .A(n15558), .B(n15526), .Z(n15529) );
  XOR U15497 ( .A(n15559), .B(n15560), .Z(n15526) );
  AND U15498 ( .A(n15561), .B(n15562), .Z(n15560) );
  XNOR U15499 ( .A(n15563), .B(n15564), .Z(n15561) );
  IV U15500 ( .A(n15559), .Z(n15563) );
  XNOR U15501 ( .A(n15565), .B(n15566), .Z(n15558) );
  NOR U15502 ( .A(n15567), .B(n15568), .Z(n15566) );
  XNOR U15503 ( .A(n15565), .B(n15569), .Z(n15567) );
  XNOR U15504 ( .A(n15525), .B(n15532), .Z(n15546) );
  NOR U15505 ( .A(n15489), .B(n15570), .Z(n15532) );
  XOR U15506 ( .A(n15537), .B(n15536), .Z(n15525) );
  XNOR U15507 ( .A(n15571), .B(n15533), .Z(n15536) );
  XOR U15508 ( .A(n15572), .B(n15573), .Z(n15533) );
  AND U15509 ( .A(n15574), .B(n15575), .Z(n15573) );
  XNOR U15510 ( .A(n15576), .B(n15577), .Z(n15574) );
  IV U15511 ( .A(n15572), .Z(n15576) );
  XNOR U15512 ( .A(n15578), .B(n15579), .Z(n15571) );
  NOR U15513 ( .A(n15580), .B(n15581), .Z(n15579) );
  XNOR U15514 ( .A(n15578), .B(n15582), .Z(n15580) );
  XOR U15515 ( .A(n15583), .B(n15584), .Z(n15537) );
  NOR U15516 ( .A(n15585), .B(n15586), .Z(n15584) );
  XNOR U15517 ( .A(n15583), .B(n15587), .Z(n15585) );
  XNOR U15518 ( .A(n15473), .B(n15542), .Z(n15544) );
  XOR U15519 ( .A(n15588), .B(n15589), .Z(n15473) );
  AND U15520 ( .A(n335), .B(n15590), .Z(n15589) );
  XOR U15521 ( .A(n15591), .B(n15588), .Z(n15590) );
  AND U15522 ( .A(n15486), .B(n15489), .Z(n15542) );
  XOR U15523 ( .A(n15592), .B(n15570), .Z(n15489) );
  XNOR U15524 ( .A(p_input[1312]), .B(p_input[2048]), .Z(n15570) );
  XNOR U15525 ( .A(n15557), .B(n15556), .Z(n15592) );
  XNOR U15526 ( .A(n15593), .B(n15564), .Z(n15556) );
  XNOR U15527 ( .A(n15552), .B(n15551), .Z(n15564) );
  XNOR U15528 ( .A(n15594), .B(n15548), .Z(n15551) );
  XNOR U15529 ( .A(p_input[1322]), .B(p_input[2058]), .Z(n15548) );
  XOR U15530 ( .A(p_input[1323]), .B(n6319), .Z(n15594) );
  XOR U15531 ( .A(p_input[1324]), .B(p_input[2060]), .Z(n15552) );
  XOR U15532 ( .A(n15562), .B(n15595), .Z(n15593) );
  IV U15533 ( .A(n15553), .Z(n15595) );
  XOR U15534 ( .A(p_input[1313]), .B(p_input[2049]), .Z(n15553) );
  XNOR U15535 ( .A(n15596), .B(n15569), .Z(n15562) );
  XNOR U15536 ( .A(p_input[1327]), .B(n6322), .Z(n15569) );
  XOR U15537 ( .A(n15559), .B(n15568), .Z(n15596) );
  XOR U15538 ( .A(n15597), .B(n15565), .Z(n15568) );
  XOR U15539 ( .A(p_input[1325]), .B(p_input[2061]), .Z(n15565) );
  XOR U15540 ( .A(p_input[1326]), .B(n6324), .Z(n15597) );
  XOR U15541 ( .A(p_input[1321]), .B(p_input[2057]), .Z(n15559) );
  XOR U15542 ( .A(n15577), .B(n15575), .Z(n15557) );
  XNOR U15543 ( .A(n15598), .B(n15582), .Z(n15575) );
  XOR U15544 ( .A(p_input[1320]), .B(p_input[2056]), .Z(n15582) );
  XOR U15545 ( .A(n15572), .B(n15581), .Z(n15598) );
  XOR U15546 ( .A(n15599), .B(n15578), .Z(n15581) );
  XOR U15547 ( .A(p_input[1318]), .B(p_input[2054]), .Z(n15578) );
  XOR U15548 ( .A(p_input[1319]), .B(n7007), .Z(n15599) );
  XOR U15549 ( .A(p_input[1314]), .B(p_input[2050]), .Z(n15572) );
  XNOR U15550 ( .A(n15587), .B(n15586), .Z(n15577) );
  XOR U15551 ( .A(n15600), .B(n15583), .Z(n15586) );
  XOR U15552 ( .A(p_input[1315]), .B(p_input[2051]), .Z(n15583) );
  XOR U15553 ( .A(p_input[1316]), .B(n7009), .Z(n15600) );
  XOR U15554 ( .A(p_input[1317]), .B(p_input[2053]), .Z(n15587) );
  XOR U15555 ( .A(n15601), .B(n15602), .Z(n15486) );
  AND U15556 ( .A(n335), .B(n15603), .Z(n15602) );
  XNOR U15557 ( .A(n15604), .B(n15601), .Z(n15603) );
  XNOR U15558 ( .A(n15605), .B(n15606), .Z(n335) );
  AND U15559 ( .A(n15607), .B(n15608), .Z(n15606) );
  XOR U15560 ( .A(n15499), .B(n15605), .Z(n15608) );
  AND U15561 ( .A(n15609), .B(n15610), .Z(n15499) );
  XNOR U15562 ( .A(n15496), .B(n15605), .Z(n15607) );
  XOR U15563 ( .A(n15611), .B(n15612), .Z(n15496) );
  AND U15564 ( .A(n339), .B(n15613), .Z(n15612) );
  XOR U15565 ( .A(n15614), .B(n15611), .Z(n15613) );
  XOR U15566 ( .A(n15615), .B(n15616), .Z(n15605) );
  AND U15567 ( .A(n15617), .B(n15618), .Z(n15616) );
  XNOR U15568 ( .A(n15615), .B(n15609), .Z(n15618) );
  IV U15569 ( .A(n15514), .Z(n15609) );
  XOR U15570 ( .A(n15619), .B(n15620), .Z(n15514) );
  XOR U15571 ( .A(n15621), .B(n15610), .Z(n15620) );
  AND U15572 ( .A(n15541), .B(n15622), .Z(n15610) );
  AND U15573 ( .A(n15623), .B(n15624), .Z(n15621) );
  XOR U15574 ( .A(n15625), .B(n15619), .Z(n15623) );
  XNOR U15575 ( .A(n15511), .B(n15615), .Z(n15617) );
  XOR U15576 ( .A(n15626), .B(n15627), .Z(n15511) );
  AND U15577 ( .A(n339), .B(n15628), .Z(n15627) );
  XOR U15578 ( .A(n15629), .B(n15626), .Z(n15628) );
  XOR U15579 ( .A(n15630), .B(n15631), .Z(n15615) );
  AND U15580 ( .A(n15632), .B(n15633), .Z(n15631) );
  XNOR U15581 ( .A(n15630), .B(n15541), .Z(n15633) );
  XOR U15582 ( .A(n15634), .B(n15624), .Z(n15541) );
  XNOR U15583 ( .A(n15635), .B(n15619), .Z(n15624) );
  XOR U15584 ( .A(n15636), .B(n15637), .Z(n15619) );
  AND U15585 ( .A(n15638), .B(n15639), .Z(n15637) );
  XOR U15586 ( .A(n15640), .B(n15636), .Z(n15638) );
  XNOR U15587 ( .A(n15641), .B(n15642), .Z(n15635) );
  AND U15588 ( .A(n15643), .B(n15644), .Z(n15642) );
  XOR U15589 ( .A(n15641), .B(n15645), .Z(n15643) );
  XNOR U15590 ( .A(n15625), .B(n15622), .Z(n15634) );
  AND U15591 ( .A(n15646), .B(n15647), .Z(n15622) );
  XOR U15592 ( .A(n15648), .B(n15649), .Z(n15625) );
  AND U15593 ( .A(n15650), .B(n15651), .Z(n15649) );
  XOR U15594 ( .A(n15648), .B(n15652), .Z(n15650) );
  XNOR U15595 ( .A(n15538), .B(n15630), .Z(n15632) );
  XOR U15596 ( .A(n15653), .B(n15654), .Z(n15538) );
  AND U15597 ( .A(n339), .B(n15655), .Z(n15654) );
  XNOR U15598 ( .A(n15656), .B(n15653), .Z(n15655) );
  XOR U15599 ( .A(n15657), .B(n15658), .Z(n15630) );
  AND U15600 ( .A(n15659), .B(n15660), .Z(n15658) );
  XNOR U15601 ( .A(n15657), .B(n15646), .Z(n15660) );
  IV U15602 ( .A(n15591), .Z(n15646) );
  XNOR U15603 ( .A(n15661), .B(n15639), .Z(n15591) );
  XNOR U15604 ( .A(n15662), .B(n15645), .Z(n15639) );
  XNOR U15605 ( .A(n15663), .B(n15664), .Z(n15645) );
  NOR U15606 ( .A(n15665), .B(n15666), .Z(n15664) );
  XOR U15607 ( .A(n15663), .B(n15667), .Z(n15665) );
  XNOR U15608 ( .A(n15644), .B(n15636), .Z(n15662) );
  XOR U15609 ( .A(n15668), .B(n15669), .Z(n15636) );
  AND U15610 ( .A(n15670), .B(n15671), .Z(n15669) );
  XOR U15611 ( .A(n15668), .B(n15672), .Z(n15670) );
  XNOR U15612 ( .A(n15673), .B(n15641), .Z(n15644) );
  XOR U15613 ( .A(n15674), .B(n15675), .Z(n15641) );
  AND U15614 ( .A(n15676), .B(n15677), .Z(n15675) );
  XNOR U15615 ( .A(n15678), .B(n15679), .Z(n15676) );
  IV U15616 ( .A(n15674), .Z(n15678) );
  XNOR U15617 ( .A(n15680), .B(n15681), .Z(n15673) );
  NOR U15618 ( .A(n15682), .B(n15683), .Z(n15681) );
  XNOR U15619 ( .A(n15680), .B(n15684), .Z(n15682) );
  XNOR U15620 ( .A(n15640), .B(n15647), .Z(n15661) );
  NOR U15621 ( .A(n15604), .B(n15685), .Z(n15647) );
  XOR U15622 ( .A(n15652), .B(n15651), .Z(n15640) );
  XNOR U15623 ( .A(n15686), .B(n15648), .Z(n15651) );
  XOR U15624 ( .A(n15687), .B(n15688), .Z(n15648) );
  AND U15625 ( .A(n15689), .B(n15690), .Z(n15688) );
  XNOR U15626 ( .A(n15691), .B(n15692), .Z(n15689) );
  IV U15627 ( .A(n15687), .Z(n15691) );
  XNOR U15628 ( .A(n15693), .B(n15694), .Z(n15686) );
  NOR U15629 ( .A(n15695), .B(n15696), .Z(n15694) );
  XNOR U15630 ( .A(n15693), .B(n15697), .Z(n15695) );
  XOR U15631 ( .A(n15698), .B(n15699), .Z(n15652) );
  NOR U15632 ( .A(n15700), .B(n15701), .Z(n15699) );
  XNOR U15633 ( .A(n15698), .B(n15702), .Z(n15700) );
  XNOR U15634 ( .A(n15588), .B(n15657), .Z(n15659) );
  XOR U15635 ( .A(n15703), .B(n15704), .Z(n15588) );
  AND U15636 ( .A(n339), .B(n15705), .Z(n15704) );
  XOR U15637 ( .A(n15706), .B(n15703), .Z(n15705) );
  AND U15638 ( .A(n15601), .B(n15604), .Z(n15657) );
  XOR U15639 ( .A(n15707), .B(n15685), .Z(n15604) );
  XNOR U15640 ( .A(p_input[1328]), .B(p_input[2048]), .Z(n15685) );
  XNOR U15641 ( .A(n15672), .B(n15671), .Z(n15707) );
  XNOR U15642 ( .A(n15708), .B(n15679), .Z(n15671) );
  XNOR U15643 ( .A(n15667), .B(n15666), .Z(n15679) );
  XNOR U15644 ( .A(n15709), .B(n15663), .Z(n15666) );
  XNOR U15645 ( .A(p_input[1338]), .B(p_input[2058]), .Z(n15663) );
  XOR U15646 ( .A(p_input[1339]), .B(n6319), .Z(n15709) );
  XOR U15647 ( .A(p_input[1340]), .B(p_input[2060]), .Z(n15667) );
  XOR U15648 ( .A(n15677), .B(n15710), .Z(n15708) );
  IV U15649 ( .A(n15668), .Z(n15710) );
  XOR U15650 ( .A(p_input[1329]), .B(p_input[2049]), .Z(n15668) );
  XNOR U15651 ( .A(n15711), .B(n15684), .Z(n15677) );
  XNOR U15652 ( .A(p_input[1343]), .B(n6322), .Z(n15684) );
  XOR U15653 ( .A(n15674), .B(n15683), .Z(n15711) );
  XOR U15654 ( .A(n15712), .B(n15680), .Z(n15683) );
  XOR U15655 ( .A(p_input[1341]), .B(p_input[2061]), .Z(n15680) );
  XOR U15656 ( .A(p_input[1342]), .B(n6324), .Z(n15712) );
  XOR U15657 ( .A(p_input[1337]), .B(p_input[2057]), .Z(n15674) );
  XOR U15658 ( .A(n15692), .B(n15690), .Z(n15672) );
  XNOR U15659 ( .A(n15713), .B(n15697), .Z(n15690) );
  XOR U15660 ( .A(p_input[1336]), .B(p_input[2056]), .Z(n15697) );
  XOR U15661 ( .A(n15687), .B(n15696), .Z(n15713) );
  XOR U15662 ( .A(n15714), .B(n15693), .Z(n15696) );
  XOR U15663 ( .A(p_input[1334]), .B(p_input[2054]), .Z(n15693) );
  XOR U15664 ( .A(p_input[1335]), .B(n7007), .Z(n15714) );
  XOR U15665 ( .A(p_input[1330]), .B(p_input[2050]), .Z(n15687) );
  XNOR U15666 ( .A(n15702), .B(n15701), .Z(n15692) );
  XOR U15667 ( .A(n15715), .B(n15698), .Z(n15701) );
  XOR U15668 ( .A(p_input[1331]), .B(p_input[2051]), .Z(n15698) );
  XOR U15669 ( .A(p_input[1332]), .B(n7009), .Z(n15715) );
  XOR U15670 ( .A(p_input[1333]), .B(p_input[2053]), .Z(n15702) );
  XOR U15671 ( .A(n15716), .B(n15717), .Z(n15601) );
  AND U15672 ( .A(n339), .B(n15718), .Z(n15717) );
  XNOR U15673 ( .A(n15719), .B(n15716), .Z(n15718) );
  XNOR U15674 ( .A(n15720), .B(n15721), .Z(n339) );
  AND U15675 ( .A(n15722), .B(n15723), .Z(n15721) );
  XOR U15676 ( .A(n15614), .B(n15720), .Z(n15723) );
  AND U15677 ( .A(n15724), .B(n15725), .Z(n15614) );
  XNOR U15678 ( .A(n15611), .B(n15720), .Z(n15722) );
  XOR U15679 ( .A(n15726), .B(n15727), .Z(n15611) );
  AND U15680 ( .A(n343), .B(n15728), .Z(n15727) );
  XOR U15681 ( .A(n15729), .B(n15726), .Z(n15728) );
  XOR U15682 ( .A(n15730), .B(n15731), .Z(n15720) );
  AND U15683 ( .A(n15732), .B(n15733), .Z(n15731) );
  XNOR U15684 ( .A(n15730), .B(n15724), .Z(n15733) );
  IV U15685 ( .A(n15629), .Z(n15724) );
  XOR U15686 ( .A(n15734), .B(n15735), .Z(n15629) );
  XOR U15687 ( .A(n15736), .B(n15725), .Z(n15735) );
  AND U15688 ( .A(n15656), .B(n15737), .Z(n15725) );
  AND U15689 ( .A(n15738), .B(n15739), .Z(n15736) );
  XOR U15690 ( .A(n15740), .B(n15734), .Z(n15738) );
  XNOR U15691 ( .A(n15626), .B(n15730), .Z(n15732) );
  XOR U15692 ( .A(n15741), .B(n15742), .Z(n15626) );
  AND U15693 ( .A(n343), .B(n15743), .Z(n15742) );
  XOR U15694 ( .A(n15744), .B(n15741), .Z(n15743) );
  XOR U15695 ( .A(n15745), .B(n15746), .Z(n15730) );
  AND U15696 ( .A(n15747), .B(n15748), .Z(n15746) );
  XNOR U15697 ( .A(n15745), .B(n15656), .Z(n15748) );
  XOR U15698 ( .A(n15749), .B(n15739), .Z(n15656) );
  XNOR U15699 ( .A(n15750), .B(n15734), .Z(n15739) );
  XOR U15700 ( .A(n15751), .B(n15752), .Z(n15734) );
  AND U15701 ( .A(n15753), .B(n15754), .Z(n15752) );
  XOR U15702 ( .A(n15755), .B(n15751), .Z(n15753) );
  XNOR U15703 ( .A(n15756), .B(n15757), .Z(n15750) );
  AND U15704 ( .A(n15758), .B(n15759), .Z(n15757) );
  XOR U15705 ( .A(n15756), .B(n15760), .Z(n15758) );
  XNOR U15706 ( .A(n15740), .B(n15737), .Z(n15749) );
  AND U15707 ( .A(n15761), .B(n15762), .Z(n15737) );
  XOR U15708 ( .A(n15763), .B(n15764), .Z(n15740) );
  AND U15709 ( .A(n15765), .B(n15766), .Z(n15764) );
  XOR U15710 ( .A(n15763), .B(n15767), .Z(n15765) );
  XNOR U15711 ( .A(n15653), .B(n15745), .Z(n15747) );
  XOR U15712 ( .A(n15768), .B(n15769), .Z(n15653) );
  AND U15713 ( .A(n343), .B(n15770), .Z(n15769) );
  XNOR U15714 ( .A(n15771), .B(n15768), .Z(n15770) );
  XOR U15715 ( .A(n15772), .B(n15773), .Z(n15745) );
  AND U15716 ( .A(n15774), .B(n15775), .Z(n15773) );
  XNOR U15717 ( .A(n15772), .B(n15761), .Z(n15775) );
  IV U15718 ( .A(n15706), .Z(n15761) );
  XNOR U15719 ( .A(n15776), .B(n15754), .Z(n15706) );
  XNOR U15720 ( .A(n15777), .B(n15760), .Z(n15754) );
  XNOR U15721 ( .A(n15778), .B(n15779), .Z(n15760) );
  NOR U15722 ( .A(n15780), .B(n15781), .Z(n15779) );
  XOR U15723 ( .A(n15778), .B(n15782), .Z(n15780) );
  XNOR U15724 ( .A(n15759), .B(n15751), .Z(n15777) );
  XOR U15725 ( .A(n15783), .B(n15784), .Z(n15751) );
  AND U15726 ( .A(n15785), .B(n15786), .Z(n15784) );
  XOR U15727 ( .A(n15783), .B(n15787), .Z(n15785) );
  XNOR U15728 ( .A(n15788), .B(n15756), .Z(n15759) );
  XOR U15729 ( .A(n15789), .B(n15790), .Z(n15756) );
  AND U15730 ( .A(n15791), .B(n15792), .Z(n15790) );
  XNOR U15731 ( .A(n15793), .B(n15794), .Z(n15791) );
  IV U15732 ( .A(n15789), .Z(n15793) );
  XNOR U15733 ( .A(n15795), .B(n15796), .Z(n15788) );
  NOR U15734 ( .A(n15797), .B(n15798), .Z(n15796) );
  XNOR U15735 ( .A(n15795), .B(n15799), .Z(n15797) );
  XNOR U15736 ( .A(n15755), .B(n15762), .Z(n15776) );
  NOR U15737 ( .A(n15719), .B(n15800), .Z(n15762) );
  XOR U15738 ( .A(n15767), .B(n15766), .Z(n15755) );
  XNOR U15739 ( .A(n15801), .B(n15763), .Z(n15766) );
  XOR U15740 ( .A(n15802), .B(n15803), .Z(n15763) );
  AND U15741 ( .A(n15804), .B(n15805), .Z(n15803) );
  XNOR U15742 ( .A(n15806), .B(n15807), .Z(n15804) );
  IV U15743 ( .A(n15802), .Z(n15806) );
  XNOR U15744 ( .A(n15808), .B(n15809), .Z(n15801) );
  NOR U15745 ( .A(n15810), .B(n15811), .Z(n15809) );
  XNOR U15746 ( .A(n15808), .B(n15812), .Z(n15810) );
  XOR U15747 ( .A(n15813), .B(n15814), .Z(n15767) );
  NOR U15748 ( .A(n15815), .B(n15816), .Z(n15814) );
  XNOR U15749 ( .A(n15813), .B(n15817), .Z(n15815) );
  XNOR U15750 ( .A(n15703), .B(n15772), .Z(n15774) );
  XOR U15751 ( .A(n15818), .B(n15819), .Z(n15703) );
  AND U15752 ( .A(n343), .B(n15820), .Z(n15819) );
  XOR U15753 ( .A(n15821), .B(n15818), .Z(n15820) );
  AND U15754 ( .A(n15716), .B(n15719), .Z(n15772) );
  XOR U15755 ( .A(n15822), .B(n15800), .Z(n15719) );
  XNOR U15756 ( .A(p_input[1344]), .B(p_input[2048]), .Z(n15800) );
  XNOR U15757 ( .A(n15787), .B(n15786), .Z(n15822) );
  XNOR U15758 ( .A(n15823), .B(n15794), .Z(n15786) );
  XNOR U15759 ( .A(n15782), .B(n15781), .Z(n15794) );
  XNOR U15760 ( .A(n15824), .B(n15778), .Z(n15781) );
  XNOR U15761 ( .A(p_input[1354]), .B(p_input[2058]), .Z(n15778) );
  XOR U15762 ( .A(p_input[1355]), .B(n6319), .Z(n15824) );
  XOR U15763 ( .A(p_input[1356]), .B(p_input[2060]), .Z(n15782) );
  XOR U15764 ( .A(n15792), .B(n15825), .Z(n15823) );
  IV U15765 ( .A(n15783), .Z(n15825) );
  XOR U15766 ( .A(p_input[1345]), .B(p_input[2049]), .Z(n15783) );
  XNOR U15767 ( .A(n15826), .B(n15799), .Z(n15792) );
  XNOR U15768 ( .A(p_input[1359]), .B(n6322), .Z(n15799) );
  XOR U15769 ( .A(n15789), .B(n15798), .Z(n15826) );
  XOR U15770 ( .A(n15827), .B(n15795), .Z(n15798) );
  XOR U15771 ( .A(p_input[1357]), .B(p_input[2061]), .Z(n15795) );
  XOR U15772 ( .A(p_input[1358]), .B(n6324), .Z(n15827) );
  XOR U15773 ( .A(p_input[1353]), .B(p_input[2057]), .Z(n15789) );
  XOR U15774 ( .A(n15807), .B(n15805), .Z(n15787) );
  XNOR U15775 ( .A(n15828), .B(n15812), .Z(n15805) );
  XOR U15776 ( .A(p_input[1352]), .B(p_input[2056]), .Z(n15812) );
  XOR U15777 ( .A(n15802), .B(n15811), .Z(n15828) );
  XOR U15778 ( .A(n15829), .B(n15808), .Z(n15811) );
  XOR U15779 ( .A(p_input[1350]), .B(p_input[2054]), .Z(n15808) );
  XOR U15780 ( .A(p_input[1351]), .B(n7007), .Z(n15829) );
  XOR U15781 ( .A(p_input[1346]), .B(p_input[2050]), .Z(n15802) );
  XNOR U15782 ( .A(n15817), .B(n15816), .Z(n15807) );
  XOR U15783 ( .A(n15830), .B(n15813), .Z(n15816) );
  XOR U15784 ( .A(p_input[1347]), .B(p_input[2051]), .Z(n15813) );
  XOR U15785 ( .A(p_input[1348]), .B(n7009), .Z(n15830) );
  XOR U15786 ( .A(p_input[1349]), .B(p_input[2053]), .Z(n15817) );
  XOR U15787 ( .A(n15831), .B(n15832), .Z(n15716) );
  AND U15788 ( .A(n343), .B(n15833), .Z(n15832) );
  XNOR U15789 ( .A(n15834), .B(n15831), .Z(n15833) );
  XNOR U15790 ( .A(n15835), .B(n15836), .Z(n343) );
  AND U15791 ( .A(n15837), .B(n15838), .Z(n15836) );
  XOR U15792 ( .A(n15729), .B(n15835), .Z(n15838) );
  AND U15793 ( .A(n15839), .B(n15840), .Z(n15729) );
  XNOR U15794 ( .A(n15726), .B(n15835), .Z(n15837) );
  XOR U15795 ( .A(n15841), .B(n15842), .Z(n15726) );
  AND U15796 ( .A(n347), .B(n15843), .Z(n15842) );
  XOR U15797 ( .A(n15844), .B(n15841), .Z(n15843) );
  XOR U15798 ( .A(n15845), .B(n15846), .Z(n15835) );
  AND U15799 ( .A(n15847), .B(n15848), .Z(n15846) );
  XNOR U15800 ( .A(n15845), .B(n15839), .Z(n15848) );
  IV U15801 ( .A(n15744), .Z(n15839) );
  XOR U15802 ( .A(n15849), .B(n15850), .Z(n15744) );
  XOR U15803 ( .A(n15851), .B(n15840), .Z(n15850) );
  AND U15804 ( .A(n15771), .B(n15852), .Z(n15840) );
  AND U15805 ( .A(n15853), .B(n15854), .Z(n15851) );
  XOR U15806 ( .A(n15855), .B(n15849), .Z(n15853) );
  XNOR U15807 ( .A(n15741), .B(n15845), .Z(n15847) );
  XOR U15808 ( .A(n15856), .B(n15857), .Z(n15741) );
  AND U15809 ( .A(n347), .B(n15858), .Z(n15857) );
  XOR U15810 ( .A(n15859), .B(n15856), .Z(n15858) );
  XOR U15811 ( .A(n15860), .B(n15861), .Z(n15845) );
  AND U15812 ( .A(n15862), .B(n15863), .Z(n15861) );
  XNOR U15813 ( .A(n15860), .B(n15771), .Z(n15863) );
  XOR U15814 ( .A(n15864), .B(n15854), .Z(n15771) );
  XNOR U15815 ( .A(n15865), .B(n15849), .Z(n15854) );
  XOR U15816 ( .A(n15866), .B(n15867), .Z(n15849) );
  AND U15817 ( .A(n15868), .B(n15869), .Z(n15867) );
  XOR U15818 ( .A(n15870), .B(n15866), .Z(n15868) );
  XNOR U15819 ( .A(n15871), .B(n15872), .Z(n15865) );
  AND U15820 ( .A(n15873), .B(n15874), .Z(n15872) );
  XOR U15821 ( .A(n15871), .B(n15875), .Z(n15873) );
  XNOR U15822 ( .A(n15855), .B(n15852), .Z(n15864) );
  AND U15823 ( .A(n15876), .B(n15877), .Z(n15852) );
  XOR U15824 ( .A(n15878), .B(n15879), .Z(n15855) );
  AND U15825 ( .A(n15880), .B(n15881), .Z(n15879) );
  XOR U15826 ( .A(n15878), .B(n15882), .Z(n15880) );
  XNOR U15827 ( .A(n15768), .B(n15860), .Z(n15862) );
  XOR U15828 ( .A(n15883), .B(n15884), .Z(n15768) );
  AND U15829 ( .A(n347), .B(n15885), .Z(n15884) );
  XNOR U15830 ( .A(n15886), .B(n15883), .Z(n15885) );
  XOR U15831 ( .A(n15887), .B(n15888), .Z(n15860) );
  AND U15832 ( .A(n15889), .B(n15890), .Z(n15888) );
  XNOR U15833 ( .A(n15887), .B(n15876), .Z(n15890) );
  IV U15834 ( .A(n15821), .Z(n15876) );
  XNOR U15835 ( .A(n15891), .B(n15869), .Z(n15821) );
  XNOR U15836 ( .A(n15892), .B(n15875), .Z(n15869) );
  XNOR U15837 ( .A(n15893), .B(n15894), .Z(n15875) );
  NOR U15838 ( .A(n15895), .B(n15896), .Z(n15894) );
  XOR U15839 ( .A(n15893), .B(n15897), .Z(n15895) );
  XNOR U15840 ( .A(n15874), .B(n15866), .Z(n15892) );
  XOR U15841 ( .A(n15898), .B(n15899), .Z(n15866) );
  AND U15842 ( .A(n15900), .B(n15901), .Z(n15899) );
  XOR U15843 ( .A(n15898), .B(n15902), .Z(n15900) );
  XNOR U15844 ( .A(n15903), .B(n15871), .Z(n15874) );
  XOR U15845 ( .A(n15904), .B(n15905), .Z(n15871) );
  AND U15846 ( .A(n15906), .B(n15907), .Z(n15905) );
  XNOR U15847 ( .A(n15908), .B(n15909), .Z(n15906) );
  IV U15848 ( .A(n15904), .Z(n15908) );
  XNOR U15849 ( .A(n15910), .B(n15911), .Z(n15903) );
  NOR U15850 ( .A(n15912), .B(n15913), .Z(n15911) );
  XNOR U15851 ( .A(n15910), .B(n15914), .Z(n15912) );
  XNOR U15852 ( .A(n15870), .B(n15877), .Z(n15891) );
  NOR U15853 ( .A(n15834), .B(n15915), .Z(n15877) );
  XOR U15854 ( .A(n15882), .B(n15881), .Z(n15870) );
  XNOR U15855 ( .A(n15916), .B(n15878), .Z(n15881) );
  XOR U15856 ( .A(n15917), .B(n15918), .Z(n15878) );
  AND U15857 ( .A(n15919), .B(n15920), .Z(n15918) );
  XNOR U15858 ( .A(n15921), .B(n15922), .Z(n15919) );
  IV U15859 ( .A(n15917), .Z(n15921) );
  XNOR U15860 ( .A(n15923), .B(n15924), .Z(n15916) );
  NOR U15861 ( .A(n15925), .B(n15926), .Z(n15924) );
  XNOR U15862 ( .A(n15923), .B(n15927), .Z(n15925) );
  XOR U15863 ( .A(n15928), .B(n15929), .Z(n15882) );
  NOR U15864 ( .A(n15930), .B(n15931), .Z(n15929) );
  XNOR U15865 ( .A(n15928), .B(n15932), .Z(n15930) );
  XNOR U15866 ( .A(n15818), .B(n15887), .Z(n15889) );
  XOR U15867 ( .A(n15933), .B(n15934), .Z(n15818) );
  AND U15868 ( .A(n347), .B(n15935), .Z(n15934) );
  XOR U15869 ( .A(n15936), .B(n15933), .Z(n15935) );
  AND U15870 ( .A(n15831), .B(n15834), .Z(n15887) );
  XOR U15871 ( .A(n15937), .B(n15915), .Z(n15834) );
  XNOR U15872 ( .A(p_input[1360]), .B(p_input[2048]), .Z(n15915) );
  XNOR U15873 ( .A(n15902), .B(n15901), .Z(n15937) );
  XNOR U15874 ( .A(n15938), .B(n15909), .Z(n15901) );
  XNOR U15875 ( .A(n15897), .B(n15896), .Z(n15909) );
  XNOR U15876 ( .A(n15939), .B(n15893), .Z(n15896) );
  XNOR U15877 ( .A(p_input[1370]), .B(p_input[2058]), .Z(n15893) );
  XOR U15878 ( .A(p_input[1371]), .B(n6319), .Z(n15939) );
  XOR U15879 ( .A(p_input[1372]), .B(p_input[2060]), .Z(n15897) );
  XOR U15880 ( .A(n15907), .B(n15940), .Z(n15938) );
  IV U15881 ( .A(n15898), .Z(n15940) );
  XOR U15882 ( .A(p_input[1361]), .B(p_input[2049]), .Z(n15898) );
  XNOR U15883 ( .A(n15941), .B(n15914), .Z(n15907) );
  XNOR U15884 ( .A(p_input[1375]), .B(n6322), .Z(n15914) );
  XOR U15885 ( .A(n15904), .B(n15913), .Z(n15941) );
  XOR U15886 ( .A(n15942), .B(n15910), .Z(n15913) );
  XOR U15887 ( .A(p_input[1373]), .B(p_input[2061]), .Z(n15910) );
  XOR U15888 ( .A(p_input[1374]), .B(n6324), .Z(n15942) );
  XOR U15889 ( .A(p_input[1369]), .B(p_input[2057]), .Z(n15904) );
  XOR U15890 ( .A(n15922), .B(n15920), .Z(n15902) );
  XNOR U15891 ( .A(n15943), .B(n15927), .Z(n15920) );
  XOR U15892 ( .A(p_input[1368]), .B(p_input[2056]), .Z(n15927) );
  XOR U15893 ( .A(n15917), .B(n15926), .Z(n15943) );
  XOR U15894 ( .A(n15944), .B(n15923), .Z(n15926) );
  XOR U15895 ( .A(p_input[1366]), .B(p_input[2054]), .Z(n15923) );
  XOR U15896 ( .A(p_input[1367]), .B(n7007), .Z(n15944) );
  XOR U15897 ( .A(p_input[1362]), .B(p_input[2050]), .Z(n15917) );
  XNOR U15898 ( .A(n15932), .B(n15931), .Z(n15922) );
  XOR U15899 ( .A(n15945), .B(n15928), .Z(n15931) );
  XOR U15900 ( .A(p_input[1363]), .B(p_input[2051]), .Z(n15928) );
  XOR U15901 ( .A(p_input[1364]), .B(n7009), .Z(n15945) );
  XOR U15902 ( .A(p_input[1365]), .B(p_input[2053]), .Z(n15932) );
  XOR U15903 ( .A(n15946), .B(n15947), .Z(n15831) );
  AND U15904 ( .A(n347), .B(n15948), .Z(n15947) );
  XNOR U15905 ( .A(n15949), .B(n15946), .Z(n15948) );
  XNOR U15906 ( .A(n15950), .B(n15951), .Z(n347) );
  AND U15907 ( .A(n15952), .B(n15953), .Z(n15951) );
  XOR U15908 ( .A(n15844), .B(n15950), .Z(n15953) );
  AND U15909 ( .A(n15954), .B(n15955), .Z(n15844) );
  XNOR U15910 ( .A(n15841), .B(n15950), .Z(n15952) );
  XOR U15911 ( .A(n15956), .B(n15957), .Z(n15841) );
  AND U15912 ( .A(n351), .B(n15958), .Z(n15957) );
  XOR U15913 ( .A(n15959), .B(n15956), .Z(n15958) );
  XOR U15914 ( .A(n15960), .B(n15961), .Z(n15950) );
  AND U15915 ( .A(n15962), .B(n15963), .Z(n15961) );
  XNOR U15916 ( .A(n15960), .B(n15954), .Z(n15963) );
  IV U15917 ( .A(n15859), .Z(n15954) );
  XOR U15918 ( .A(n15964), .B(n15965), .Z(n15859) );
  XOR U15919 ( .A(n15966), .B(n15955), .Z(n15965) );
  AND U15920 ( .A(n15886), .B(n15967), .Z(n15955) );
  AND U15921 ( .A(n15968), .B(n15969), .Z(n15966) );
  XOR U15922 ( .A(n15970), .B(n15964), .Z(n15968) );
  XNOR U15923 ( .A(n15856), .B(n15960), .Z(n15962) );
  XOR U15924 ( .A(n15971), .B(n15972), .Z(n15856) );
  AND U15925 ( .A(n351), .B(n15973), .Z(n15972) );
  XOR U15926 ( .A(n15974), .B(n15971), .Z(n15973) );
  XOR U15927 ( .A(n15975), .B(n15976), .Z(n15960) );
  AND U15928 ( .A(n15977), .B(n15978), .Z(n15976) );
  XNOR U15929 ( .A(n15975), .B(n15886), .Z(n15978) );
  XOR U15930 ( .A(n15979), .B(n15969), .Z(n15886) );
  XNOR U15931 ( .A(n15980), .B(n15964), .Z(n15969) );
  XOR U15932 ( .A(n15981), .B(n15982), .Z(n15964) );
  AND U15933 ( .A(n15983), .B(n15984), .Z(n15982) );
  XOR U15934 ( .A(n15985), .B(n15981), .Z(n15983) );
  XNOR U15935 ( .A(n15986), .B(n15987), .Z(n15980) );
  AND U15936 ( .A(n15988), .B(n15989), .Z(n15987) );
  XOR U15937 ( .A(n15986), .B(n15990), .Z(n15988) );
  XNOR U15938 ( .A(n15970), .B(n15967), .Z(n15979) );
  AND U15939 ( .A(n15991), .B(n15992), .Z(n15967) );
  XOR U15940 ( .A(n15993), .B(n15994), .Z(n15970) );
  AND U15941 ( .A(n15995), .B(n15996), .Z(n15994) );
  XOR U15942 ( .A(n15993), .B(n15997), .Z(n15995) );
  XNOR U15943 ( .A(n15883), .B(n15975), .Z(n15977) );
  XOR U15944 ( .A(n15998), .B(n15999), .Z(n15883) );
  AND U15945 ( .A(n351), .B(n16000), .Z(n15999) );
  XNOR U15946 ( .A(n16001), .B(n15998), .Z(n16000) );
  XOR U15947 ( .A(n16002), .B(n16003), .Z(n15975) );
  AND U15948 ( .A(n16004), .B(n16005), .Z(n16003) );
  XNOR U15949 ( .A(n16002), .B(n15991), .Z(n16005) );
  IV U15950 ( .A(n15936), .Z(n15991) );
  XNOR U15951 ( .A(n16006), .B(n15984), .Z(n15936) );
  XNOR U15952 ( .A(n16007), .B(n15990), .Z(n15984) );
  XNOR U15953 ( .A(n16008), .B(n16009), .Z(n15990) );
  NOR U15954 ( .A(n16010), .B(n16011), .Z(n16009) );
  XOR U15955 ( .A(n16008), .B(n16012), .Z(n16010) );
  XNOR U15956 ( .A(n15989), .B(n15981), .Z(n16007) );
  XOR U15957 ( .A(n16013), .B(n16014), .Z(n15981) );
  AND U15958 ( .A(n16015), .B(n16016), .Z(n16014) );
  XOR U15959 ( .A(n16013), .B(n16017), .Z(n16015) );
  XNOR U15960 ( .A(n16018), .B(n15986), .Z(n15989) );
  XOR U15961 ( .A(n16019), .B(n16020), .Z(n15986) );
  AND U15962 ( .A(n16021), .B(n16022), .Z(n16020) );
  XNOR U15963 ( .A(n16023), .B(n16024), .Z(n16021) );
  IV U15964 ( .A(n16019), .Z(n16023) );
  XNOR U15965 ( .A(n16025), .B(n16026), .Z(n16018) );
  NOR U15966 ( .A(n16027), .B(n16028), .Z(n16026) );
  XNOR U15967 ( .A(n16025), .B(n16029), .Z(n16027) );
  XNOR U15968 ( .A(n15985), .B(n15992), .Z(n16006) );
  NOR U15969 ( .A(n15949), .B(n16030), .Z(n15992) );
  XOR U15970 ( .A(n15997), .B(n15996), .Z(n15985) );
  XNOR U15971 ( .A(n16031), .B(n15993), .Z(n15996) );
  XOR U15972 ( .A(n16032), .B(n16033), .Z(n15993) );
  AND U15973 ( .A(n16034), .B(n16035), .Z(n16033) );
  XNOR U15974 ( .A(n16036), .B(n16037), .Z(n16034) );
  IV U15975 ( .A(n16032), .Z(n16036) );
  XNOR U15976 ( .A(n16038), .B(n16039), .Z(n16031) );
  NOR U15977 ( .A(n16040), .B(n16041), .Z(n16039) );
  XNOR U15978 ( .A(n16038), .B(n16042), .Z(n16040) );
  XOR U15979 ( .A(n16043), .B(n16044), .Z(n15997) );
  NOR U15980 ( .A(n16045), .B(n16046), .Z(n16044) );
  XNOR U15981 ( .A(n16043), .B(n16047), .Z(n16045) );
  XNOR U15982 ( .A(n15933), .B(n16002), .Z(n16004) );
  XOR U15983 ( .A(n16048), .B(n16049), .Z(n15933) );
  AND U15984 ( .A(n351), .B(n16050), .Z(n16049) );
  XOR U15985 ( .A(n16051), .B(n16048), .Z(n16050) );
  AND U15986 ( .A(n15946), .B(n15949), .Z(n16002) );
  XOR U15987 ( .A(n16052), .B(n16030), .Z(n15949) );
  XNOR U15988 ( .A(p_input[1376]), .B(p_input[2048]), .Z(n16030) );
  XNOR U15989 ( .A(n16017), .B(n16016), .Z(n16052) );
  XNOR U15990 ( .A(n16053), .B(n16024), .Z(n16016) );
  XNOR U15991 ( .A(n16012), .B(n16011), .Z(n16024) );
  XNOR U15992 ( .A(n16054), .B(n16008), .Z(n16011) );
  XNOR U15993 ( .A(p_input[1386]), .B(p_input[2058]), .Z(n16008) );
  XOR U15994 ( .A(p_input[1387]), .B(n6319), .Z(n16054) );
  XOR U15995 ( .A(p_input[1388]), .B(p_input[2060]), .Z(n16012) );
  XOR U15996 ( .A(n16022), .B(n16055), .Z(n16053) );
  IV U15997 ( .A(n16013), .Z(n16055) );
  XOR U15998 ( .A(p_input[1377]), .B(p_input[2049]), .Z(n16013) );
  XNOR U15999 ( .A(n16056), .B(n16029), .Z(n16022) );
  XNOR U16000 ( .A(p_input[1391]), .B(n6322), .Z(n16029) );
  XOR U16001 ( .A(n16019), .B(n16028), .Z(n16056) );
  XOR U16002 ( .A(n16057), .B(n16025), .Z(n16028) );
  XOR U16003 ( .A(p_input[1389]), .B(p_input[2061]), .Z(n16025) );
  XOR U16004 ( .A(p_input[1390]), .B(n6324), .Z(n16057) );
  XOR U16005 ( .A(p_input[1385]), .B(p_input[2057]), .Z(n16019) );
  XOR U16006 ( .A(n16037), .B(n16035), .Z(n16017) );
  XNOR U16007 ( .A(n16058), .B(n16042), .Z(n16035) );
  XOR U16008 ( .A(p_input[1384]), .B(p_input[2056]), .Z(n16042) );
  XOR U16009 ( .A(n16032), .B(n16041), .Z(n16058) );
  XOR U16010 ( .A(n16059), .B(n16038), .Z(n16041) );
  XOR U16011 ( .A(p_input[1382]), .B(p_input[2054]), .Z(n16038) );
  XOR U16012 ( .A(p_input[1383]), .B(n7007), .Z(n16059) );
  XOR U16013 ( .A(p_input[1378]), .B(p_input[2050]), .Z(n16032) );
  XNOR U16014 ( .A(n16047), .B(n16046), .Z(n16037) );
  XOR U16015 ( .A(n16060), .B(n16043), .Z(n16046) );
  XOR U16016 ( .A(p_input[1379]), .B(p_input[2051]), .Z(n16043) );
  XOR U16017 ( .A(p_input[1380]), .B(n7009), .Z(n16060) );
  XOR U16018 ( .A(p_input[1381]), .B(p_input[2053]), .Z(n16047) );
  XOR U16019 ( .A(n16061), .B(n16062), .Z(n15946) );
  AND U16020 ( .A(n351), .B(n16063), .Z(n16062) );
  XNOR U16021 ( .A(n16064), .B(n16061), .Z(n16063) );
  XNOR U16022 ( .A(n16065), .B(n16066), .Z(n351) );
  AND U16023 ( .A(n16067), .B(n16068), .Z(n16066) );
  XOR U16024 ( .A(n15959), .B(n16065), .Z(n16068) );
  AND U16025 ( .A(n16069), .B(n16070), .Z(n15959) );
  XNOR U16026 ( .A(n15956), .B(n16065), .Z(n16067) );
  XOR U16027 ( .A(n16071), .B(n16072), .Z(n15956) );
  AND U16028 ( .A(n355), .B(n16073), .Z(n16072) );
  XOR U16029 ( .A(n16074), .B(n16071), .Z(n16073) );
  XOR U16030 ( .A(n16075), .B(n16076), .Z(n16065) );
  AND U16031 ( .A(n16077), .B(n16078), .Z(n16076) );
  XNOR U16032 ( .A(n16075), .B(n16069), .Z(n16078) );
  IV U16033 ( .A(n15974), .Z(n16069) );
  XOR U16034 ( .A(n16079), .B(n16080), .Z(n15974) );
  XOR U16035 ( .A(n16081), .B(n16070), .Z(n16080) );
  AND U16036 ( .A(n16001), .B(n16082), .Z(n16070) );
  AND U16037 ( .A(n16083), .B(n16084), .Z(n16081) );
  XOR U16038 ( .A(n16085), .B(n16079), .Z(n16083) );
  XNOR U16039 ( .A(n15971), .B(n16075), .Z(n16077) );
  XOR U16040 ( .A(n16086), .B(n16087), .Z(n15971) );
  AND U16041 ( .A(n355), .B(n16088), .Z(n16087) );
  XOR U16042 ( .A(n16089), .B(n16086), .Z(n16088) );
  XOR U16043 ( .A(n16090), .B(n16091), .Z(n16075) );
  AND U16044 ( .A(n16092), .B(n16093), .Z(n16091) );
  XNOR U16045 ( .A(n16090), .B(n16001), .Z(n16093) );
  XOR U16046 ( .A(n16094), .B(n16084), .Z(n16001) );
  XNOR U16047 ( .A(n16095), .B(n16079), .Z(n16084) );
  XOR U16048 ( .A(n16096), .B(n16097), .Z(n16079) );
  AND U16049 ( .A(n16098), .B(n16099), .Z(n16097) );
  XOR U16050 ( .A(n16100), .B(n16096), .Z(n16098) );
  XNOR U16051 ( .A(n16101), .B(n16102), .Z(n16095) );
  AND U16052 ( .A(n16103), .B(n16104), .Z(n16102) );
  XOR U16053 ( .A(n16101), .B(n16105), .Z(n16103) );
  XNOR U16054 ( .A(n16085), .B(n16082), .Z(n16094) );
  AND U16055 ( .A(n16106), .B(n16107), .Z(n16082) );
  XOR U16056 ( .A(n16108), .B(n16109), .Z(n16085) );
  AND U16057 ( .A(n16110), .B(n16111), .Z(n16109) );
  XOR U16058 ( .A(n16108), .B(n16112), .Z(n16110) );
  XNOR U16059 ( .A(n15998), .B(n16090), .Z(n16092) );
  XOR U16060 ( .A(n16113), .B(n16114), .Z(n15998) );
  AND U16061 ( .A(n355), .B(n16115), .Z(n16114) );
  XNOR U16062 ( .A(n16116), .B(n16113), .Z(n16115) );
  XOR U16063 ( .A(n16117), .B(n16118), .Z(n16090) );
  AND U16064 ( .A(n16119), .B(n16120), .Z(n16118) );
  XNOR U16065 ( .A(n16117), .B(n16106), .Z(n16120) );
  IV U16066 ( .A(n16051), .Z(n16106) );
  XNOR U16067 ( .A(n16121), .B(n16099), .Z(n16051) );
  XNOR U16068 ( .A(n16122), .B(n16105), .Z(n16099) );
  XNOR U16069 ( .A(n16123), .B(n16124), .Z(n16105) );
  NOR U16070 ( .A(n16125), .B(n16126), .Z(n16124) );
  XOR U16071 ( .A(n16123), .B(n16127), .Z(n16125) );
  XNOR U16072 ( .A(n16104), .B(n16096), .Z(n16122) );
  XOR U16073 ( .A(n16128), .B(n16129), .Z(n16096) );
  AND U16074 ( .A(n16130), .B(n16131), .Z(n16129) );
  XOR U16075 ( .A(n16128), .B(n16132), .Z(n16130) );
  XNOR U16076 ( .A(n16133), .B(n16101), .Z(n16104) );
  XOR U16077 ( .A(n16134), .B(n16135), .Z(n16101) );
  AND U16078 ( .A(n16136), .B(n16137), .Z(n16135) );
  XNOR U16079 ( .A(n16138), .B(n16139), .Z(n16136) );
  IV U16080 ( .A(n16134), .Z(n16138) );
  XNOR U16081 ( .A(n16140), .B(n16141), .Z(n16133) );
  NOR U16082 ( .A(n16142), .B(n16143), .Z(n16141) );
  XNOR U16083 ( .A(n16140), .B(n16144), .Z(n16142) );
  XNOR U16084 ( .A(n16100), .B(n16107), .Z(n16121) );
  NOR U16085 ( .A(n16064), .B(n16145), .Z(n16107) );
  XOR U16086 ( .A(n16112), .B(n16111), .Z(n16100) );
  XNOR U16087 ( .A(n16146), .B(n16108), .Z(n16111) );
  XOR U16088 ( .A(n16147), .B(n16148), .Z(n16108) );
  AND U16089 ( .A(n16149), .B(n16150), .Z(n16148) );
  XNOR U16090 ( .A(n16151), .B(n16152), .Z(n16149) );
  IV U16091 ( .A(n16147), .Z(n16151) );
  XNOR U16092 ( .A(n16153), .B(n16154), .Z(n16146) );
  NOR U16093 ( .A(n16155), .B(n16156), .Z(n16154) );
  XNOR U16094 ( .A(n16153), .B(n16157), .Z(n16155) );
  XOR U16095 ( .A(n16158), .B(n16159), .Z(n16112) );
  NOR U16096 ( .A(n16160), .B(n16161), .Z(n16159) );
  XNOR U16097 ( .A(n16158), .B(n16162), .Z(n16160) );
  XNOR U16098 ( .A(n16048), .B(n16117), .Z(n16119) );
  XOR U16099 ( .A(n16163), .B(n16164), .Z(n16048) );
  AND U16100 ( .A(n355), .B(n16165), .Z(n16164) );
  XOR U16101 ( .A(n16166), .B(n16163), .Z(n16165) );
  AND U16102 ( .A(n16061), .B(n16064), .Z(n16117) );
  XOR U16103 ( .A(n16167), .B(n16145), .Z(n16064) );
  XNOR U16104 ( .A(p_input[1392]), .B(p_input[2048]), .Z(n16145) );
  XNOR U16105 ( .A(n16132), .B(n16131), .Z(n16167) );
  XNOR U16106 ( .A(n16168), .B(n16139), .Z(n16131) );
  XNOR U16107 ( .A(n16127), .B(n16126), .Z(n16139) );
  XNOR U16108 ( .A(n16169), .B(n16123), .Z(n16126) );
  XNOR U16109 ( .A(p_input[1402]), .B(p_input[2058]), .Z(n16123) );
  XOR U16110 ( .A(p_input[1403]), .B(n6319), .Z(n16169) );
  XOR U16111 ( .A(p_input[1404]), .B(p_input[2060]), .Z(n16127) );
  XOR U16112 ( .A(n16137), .B(n16170), .Z(n16168) );
  IV U16113 ( .A(n16128), .Z(n16170) );
  XOR U16114 ( .A(p_input[1393]), .B(p_input[2049]), .Z(n16128) );
  XNOR U16115 ( .A(n16171), .B(n16144), .Z(n16137) );
  XNOR U16116 ( .A(p_input[1407]), .B(n6322), .Z(n16144) );
  XOR U16117 ( .A(n16134), .B(n16143), .Z(n16171) );
  XOR U16118 ( .A(n16172), .B(n16140), .Z(n16143) );
  XOR U16119 ( .A(p_input[1405]), .B(p_input[2061]), .Z(n16140) );
  XOR U16120 ( .A(p_input[1406]), .B(n6324), .Z(n16172) );
  XOR U16121 ( .A(p_input[1401]), .B(p_input[2057]), .Z(n16134) );
  XOR U16122 ( .A(n16152), .B(n16150), .Z(n16132) );
  XNOR U16123 ( .A(n16173), .B(n16157), .Z(n16150) );
  XOR U16124 ( .A(p_input[1400]), .B(p_input[2056]), .Z(n16157) );
  XOR U16125 ( .A(n16147), .B(n16156), .Z(n16173) );
  XOR U16126 ( .A(n16174), .B(n16153), .Z(n16156) );
  XOR U16127 ( .A(p_input[1398]), .B(p_input[2054]), .Z(n16153) );
  XOR U16128 ( .A(p_input[1399]), .B(n7007), .Z(n16174) );
  XOR U16129 ( .A(p_input[1394]), .B(p_input[2050]), .Z(n16147) );
  XNOR U16130 ( .A(n16162), .B(n16161), .Z(n16152) );
  XOR U16131 ( .A(n16175), .B(n16158), .Z(n16161) );
  XOR U16132 ( .A(p_input[1395]), .B(p_input[2051]), .Z(n16158) );
  XOR U16133 ( .A(p_input[1396]), .B(n7009), .Z(n16175) );
  XOR U16134 ( .A(p_input[1397]), .B(p_input[2053]), .Z(n16162) );
  XOR U16135 ( .A(n16176), .B(n16177), .Z(n16061) );
  AND U16136 ( .A(n355), .B(n16178), .Z(n16177) );
  XNOR U16137 ( .A(n16179), .B(n16176), .Z(n16178) );
  XNOR U16138 ( .A(n16180), .B(n16181), .Z(n355) );
  AND U16139 ( .A(n16182), .B(n16183), .Z(n16181) );
  XOR U16140 ( .A(n16074), .B(n16180), .Z(n16183) );
  AND U16141 ( .A(n16184), .B(n16185), .Z(n16074) );
  XNOR U16142 ( .A(n16071), .B(n16180), .Z(n16182) );
  XOR U16143 ( .A(n16186), .B(n16187), .Z(n16071) );
  AND U16144 ( .A(n359), .B(n16188), .Z(n16187) );
  XOR U16145 ( .A(n16189), .B(n16186), .Z(n16188) );
  XOR U16146 ( .A(n16190), .B(n16191), .Z(n16180) );
  AND U16147 ( .A(n16192), .B(n16193), .Z(n16191) );
  XNOR U16148 ( .A(n16190), .B(n16184), .Z(n16193) );
  IV U16149 ( .A(n16089), .Z(n16184) );
  XOR U16150 ( .A(n16194), .B(n16195), .Z(n16089) );
  XOR U16151 ( .A(n16196), .B(n16185), .Z(n16195) );
  AND U16152 ( .A(n16116), .B(n16197), .Z(n16185) );
  AND U16153 ( .A(n16198), .B(n16199), .Z(n16196) );
  XOR U16154 ( .A(n16200), .B(n16194), .Z(n16198) );
  XNOR U16155 ( .A(n16086), .B(n16190), .Z(n16192) );
  XOR U16156 ( .A(n16201), .B(n16202), .Z(n16086) );
  AND U16157 ( .A(n359), .B(n16203), .Z(n16202) );
  XOR U16158 ( .A(n16204), .B(n16201), .Z(n16203) );
  XOR U16159 ( .A(n16205), .B(n16206), .Z(n16190) );
  AND U16160 ( .A(n16207), .B(n16208), .Z(n16206) );
  XNOR U16161 ( .A(n16205), .B(n16116), .Z(n16208) );
  XOR U16162 ( .A(n16209), .B(n16199), .Z(n16116) );
  XNOR U16163 ( .A(n16210), .B(n16194), .Z(n16199) );
  XOR U16164 ( .A(n16211), .B(n16212), .Z(n16194) );
  AND U16165 ( .A(n16213), .B(n16214), .Z(n16212) );
  XOR U16166 ( .A(n16215), .B(n16211), .Z(n16213) );
  XNOR U16167 ( .A(n16216), .B(n16217), .Z(n16210) );
  AND U16168 ( .A(n16218), .B(n16219), .Z(n16217) );
  XOR U16169 ( .A(n16216), .B(n16220), .Z(n16218) );
  XNOR U16170 ( .A(n16200), .B(n16197), .Z(n16209) );
  AND U16171 ( .A(n16221), .B(n16222), .Z(n16197) );
  XOR U16172 ( .A(n16223), .B(n16224), .Z(n16200) );
  AND U16173 ( .A(n16225), .B(n16226), .Z(n16224) );
  XOR U16174 ( .A(n16223), .B(n16227), .Z(n16225) );
  XNOR U16175 ( .A(n16113), .B(n16205), .Z(n16207) );
  XOR U16176 ( .A(n16228), .B(n16229), .Z(n16113) );
  AND U16177 ( .A(n359), .B(n16230), .Z(n16229) );
  XNOR U16178 ( .A(n16231), .B(n16228), .Z(n16230) );
  XOR U16179 ( .A(n16232), .B(n16233), .Z(n16205) );
  AND U16180 ( .A(n16234), .B(n16235), .Z(n16233) );
  XNOR U16181 ( .A(n16232), .B(n16221), .Z(n16235) );
  IV U16182 ( .A(n16166), .Z(n16221) );
  XNOR U16183 ( .A(n16236), .B(n16214), .Z(n16166) );
  XNOR U16184 ( .A(n16237), .B(n16220), .Z(n16214) );
  XNOR U16185 ( .A(n16238), .B(n16239), .Z(n16220) );
  NOR U16186 ( .A(n16240), .B(n16241), .Z(n16239) );
  XOR U16187 ( .A(n16238), .B(n16242), .Z(n16240) );
  XNOR U16188 ( .A(n16219), .B(n16211), .Z(n16237) );
  XOR U16189 ( .A(n16243), .B(n16244), .Z(n16211) );
  AND U16190 ( .A(n16245), .B(n16246), .Z(n16244) );
  XOR U16191 ( .A(n16243), .B(n16247), .Z(n16245) );
  XNOR U16192 ( .A(n16248), .B(n16216), .Z(n16219) );
  XOR U16193 ( .A(n16249), .B(n16250), .Z(n16216) );
  AND U16194 ( .A(n16251), .B(n16252), .Z(n16250) );
  XNOR U16195 ( .A(n16253), .B(n16254), .Z(n16251) );
  IV U16196 ( .A(n16249), .Z(n16253) );
  XNOR U16197 ( .A(n16255), .B(n16256), .Z(n16248) );
  NOR U16198 ( .A(n16257), .B(n16258), .Z(n16256) );
  XNOR U16199 ( .A(n16255), .B(n16259), .Z(n16257) );
  XNOR U16200 ( .A(n16215), .B(n16222), .Z(n16236) );
  NOR U16201 ( .A(n16179), .B(n16260), .Z(n16222) );
  XOR U16202 ( .A(n16227), .B(n16226), .Z(n16215) );
  XNOR U16203 ( .A(n16261), .B(n16223), .Z(n16226) );
  XOR U16204 ( .A(n16262), .B(n16263), .Z(n16223) );
  AND U16205 ( .A(n16264), .B(n16265), .Z(n16263) );
  XNOR U16206 ( .A(n16266), .B(n16267), .Z(n16264) );
  IV U16207 ( .A(n16262), .Z(n16266) );
  XNOR U16208 ( .A(n16268), .B(n16269), .Z(n16261) );
  NOR U16209 ( .A(n16270), .B(n16271), .Z(n16269) );
  XNOR U16210 ( .A(n16268), .B(n16272), .Z(n16270) );
  XOR U16211 ( .A(n16273), .B(n16274), .Z(n16227) );
  NOR U16212 ( .A(n16275), .B(n16276), .Z(n16274) );
  XNOR U16213 ( .A(n16273), .B(n16277), .Z(n16275) );
  XNOR U16214 ( .A(n16163), .B(n16232), .Z(n16234) );
  XOR U16215 ( .A(n16278), .B(n16279), .Z(n16163) );
  AND U16216 ( .A(n359), .B(n16280), .Z(n16279) );
  XOR U16217 ( .A(n16281), .B(n16278), .Z(n16280) );
  AND U16218 ( .A(n16176), .B(n16179), .Z(n16232) );
  XOR U16219 ( .A(n16282), .B(n16260), .Z(n16179) );
  XNOR U16220 ( .A(p_input[1408]), .B(p_input[2048]), .Z(n16260) );
  XNOR U16221 ( .A(n16247), .B(n16246), .Z(n16282) );
  XNOR U16222 ( .A(n16283), .B(n16254), .Z(n16246) );
  XNOR U16223 ( .A(n16242), .B(n16241), .Z(n16254) );
  XNOR U16224 ( .A(n16284), .B(n16238), .Z(n16241) );
  XNOR U16225 ( .A(p_input[1418]), .B(p_input[2058]), .Z(n16238) );
  XOR U16226 ( .A(p_input[1419]), .B(n6319), .Z(n16284) );
  XOR U16227 ( .A(p_input[1420]), .B(p_input[2060]), .Z(n16242) );
  XOR U16228 ( .A(n16252), .B(n16285), .Z(n16283) );
  IV U16229 ( .A(n16243), .Z(n16285) );
  XOR U16230 ( .A(p_input[1409]), .B(p_input[2049]), .Z(n16243) );
  XNOR U16231 ( .A(n16286), .B(n16259), .Z(n16252) );
  XNOR U16232 ( .A(p_input[1423]), .B(n6322), .Z(n16259) );
  XOR U16233 ( .A(n16249), .B(n16258), .Z(n16286) );
  XOR U16234 ( .A(n16287), .B(n16255), .Z(n16258) );
  XOR U16235 ( .A(p_input[1421]), .B(p_input[2061]), .Z(n16255) );
  XOR U16236 ( .A(p_input[1422]), .B(n6324), .Z(n16287) );
  XOR U16237 ( .A(p_input[1417]), .B(p_input[2057]), .Z(n16249) );
  XOR U16238 ( .A(n16267), .B(n16265), .Z(n16247) );
  XNOR U16239 ( .A(n16288), .B(n16272), .Z(n16265) );
  XOR U16240 ( .A(p_input[1416]), .B(p_input[2056]), .Z(n16272) );
  XOR U16241 ( .A(n16262), .B(n16271), .Z(n16288) );
  XOR U16242 ( .A(n16289), .B(n16268), .Z(n16271) );
  XOR U16243 ( .A(p_input[1414]), .B(p_input[2054]), .Z(n16268) );
  XOR U16244 ( .A(p_input[1415]), .B(n7007), .Z(n16289) );
  XOR U16245 ( .A(p_input[1410]), .B(p_input[2050]), .Z(n16262) );
  XNOR U16246 ( .A(n16277), .B(n16276), .Z(n16267) );
  XOR U16247 ( .A(n16290), .B(n16273), .Z(n16276) );
  XOR U16248 ( .A(p_input[1411]), .B(p_input[2051]), .Z(n16273) );
  XOR U16249 ( .A(p_input[1412]), .B(n7009), .Z(n16290) );
  XOR U16250 ( .A(p_input[1413]), .B(p_input[2053]), .Z(n16277) );
  XOR U16251 ( .A(n16291), .B(n16292), .Z(n16176) );
  AND U16252 ( .A(n359), .B(n16293), .Z(n16292) );
  XNOR U16253 ( .A(n16294), .B(n16291), .Z(n16293) );
  XNOR U16254 ( .A(n16295), .B(n16296), .Z(n359) );
  AND U16255 ( .A(n16297), .B(n16298), .Z(n16296) );
  XOR U16256 ( .A(n16189), .B(n16295), .Z(n16298) );
  AND U16257 ( .A(n16299), .B(n16300), .Z(n16189) );
  XNOR U16258 ( .A(n16186), .B(n16295), .Z(n16297) );
  XOR U16259 ( .A(n16301), .B(n16302), .Z(n16186) );
  AND U16260 ( .A(n363), .B(n16303), .Z(n16302) );
  XOR U16261 ( .A(n16304), .B(n16301), .Z(n16303) );
  XOR U16262 ( .A(n16305), .B(n16306), .Z(n16295) );
  AND U16263 ( .A(n16307), .B(n16308), .Z(n16306) );
  XNOR U16264 ( .A(n16305), .B(n16299), .Z(n16308) );
  IV U16265 ( .A(n16204), .Z(n16299) );
  XOR U16266 ( .A(n16309), .B(n16310), .Z(n16204) );
  XOR U16267 ( .A(n16311), .B(n16300), .Z(n16310) );
  AND U16268 ( .A(n16231), .B(n16312), .Z(n16300) );
  AND U16269 ( .A(n16313), .B(n16314), .Z(n16311) );
  XOR U16270 ( .A(n16315), .B(n16309), .Z(n16313) );
  XNOR U16271 ( .A(n16201), .B(n16305), .Z(n16307) );
  XOR U16272 ( .A(n16316), .B(n16317), .Z(n16201) );
  AND U16273 ( .A(n363), .B(n16318), .Z(n16317) );
  XOR U16274 ( .A(n16319), .B(n16316), .Z(n16318) );
  XOR U16275 ( .A(n16320), .B(n16321), .Z(n16305) );
  AND U16276 ( .A(n16322), .B(n16323), .Z(n16321) );
  XNOR U16277 ( .A(n16320), .B(n16231), .Z(n16323) );
  XOR U16278 ( .A(n16324), .B(n16314), .Z(n16231) );
  XNOR U16279 ( .A(n16325), .B(n16309), .Z(n16314) );
  XOR U16280 ( .A(n16326), .B(n16327), .Z(n16309) );
  AND U16281 ( .A(n16328), .B(n16329), .Z(n16327) );
  XOR U16282 ( .A(n16330), .B(n16326), .Z(n16328) );
  XNOR U16283 ( .A(n16331), .B(n16332), .Z(n16325) );
  AND U16284 ( .A(n16333), .B(n16334), .Z(n16332) );
  XOR U16285 ( .A(n16331), .B(n16335), .Z(n16333) );
  XNOR U16286 ( .A(n16315), .B(n16312), .Z(n16324) );
  AND U16287 ( .A(n16336), .B(n16337), .Z(n16312) );
  XOR U16288 ( .A(n16338), .B(n16339), .Z(n16315) );
  AND U16289 ( .A(n16340), .B(n16341), .Z(n16339) );
  XOR U16290 ( .A(n16338), .B(n16342), .Z(n16340) );
  XNOR U16291 ( .A(n16228), .B(n16320), .Z(n16322) );
  XOR U16292 ( .A(n16343), .B(n16344), .Z(n16228) );
  AND U16293 ( .A(n363), .B(n16345), .Z(n16344) );
  XNOR U16294 ( .A(n16346), .B(n16343), .Z(n16345) );
  XOR U16295 ( .A(n16347), .B(n16348), .Z(n16320) );
  AND U16296 ( .A(n16349), .B(n16350), .Z(n16348) );
  XNOR U16297 ( .A(n16347), .B(n16336), .Z(n16350) );
  IV U16298 ( .A(n16281), .Z(n16336) );
  XNOR U16299 ( .A(n16351), .B(n16329), .Z(n16281) );
  XNOR U16300 ( .A(n16352), .B(n16335), .Z(n16329) );
  XNOR U16301 ( .A(n16353), .B(n16354), .Z(n16335) );
  NOR U16302 ( .A(n16355), .B(n16356), .Z(n16354) );
  XOR U16303 ( .A(n16353), .B(n16357), .Z(n16355) );
  XNOR U16304 ( .A(n16334), .B(n16326), .Z(n16352) );
  XOR U16305 ( .A(n16358), .B(n16359), .Z(n16326) );
  AND U16306 ( .A(n16360), .B(n16361), .Z(n16359) );
  XOR U16307 ( .A(n16358), .B(n16362), .Z(n16360) );
  XNOR U16308 ( .A(n16363), .B(n16331), .Z(n16334) );
  XOR U16309 ( .A(n16364), .B(n16365), .Z(n16331) );
  AND U16310 ( .A(n16366), .B(n16367), .Z(n16365) );
  XNOR U16311 ( .A(n16368), .B(n16369), .Z(n16366) );
  IV U16312 ( .A(n16364), .Z(n16368) );
  XNOR U16313 ( .A(n16370), .B(n16371), .Z(n16363) );
  NOR U16314 ( .A(n16372), .B(n16373), .Z(n16371) );
  XNOR U16315 ( .A(n16370), .B(n16374), .Z(n16372) );
  XNOR U16316 ( .A(n16330), .B(n16337), .Z(n16351) );
  NOR U16317 ( .A(n16294), .B(n16375), .Z(n16337) );
  XOR U16318 ( .A(n16342), .B(n16341), .Z(n16330) );
  XNOR U16319 ( .A(n16376), .B(n16338), .Z(n16341) );
  XOR U16320 ( .A(n16377), .B(n16378), .Z(n16338) );
  AND U16321 ( .A(n16379), .B(n16380), .Z(n16378) );
  XNOR U16322 ( .A(n16381), .B(n16382), .Z(n16379) );
  IV U16323 ( .A(n16377), .Z(n16381) );
  XNOR U16324 ( .A(n16383), .B(n16384), .Z(n16376) );
  NOR U16325 ( .A(n16385), .B(n16386), .Z(n16384) );
  XNOR U16326 ( .A(n16383), .B(n16387), .Z(n16385) );
  XOR U16327 ( .A(n16388), .B(n16389), .Z(n16342) );
  NOR U16328 ( .A(n16390), .B(n16391), .Z(n16389) );
  XNOR U16329 ( .A(n16388), .B(n16392), .Z(n16390) );
  XNOR U16330 ( .A(n16278), .B(n16347), .Z(n16349) );
  XOR U16331 ( .A(n16393), .B(n16394), .Z(n16278) );
  AND U16332 ( .A(n363), .B(n16395), .Z(n16394) );
  XOR U16333 ( .A(n16396), .B(n16393), .Z(n16395) );
  AND U16334 ( .A(n16291), .B(n16294), .Z(n16347) );
  XOR U16335 ( .A(n16397), .B(n16375), .Z(n16294) );
  XNOR U16336 ( .A(p_input[1424]), .B(p_input[2048]), .Z(n16375) );
  XNOR U16337 ( .A(n16362), .B(n16361), .Z(n16397) );
  XNOR U16338 ( .A(n16398), .B(n16369), .Z(n16361) );
  XNOR U16339 ( .A(n16357), .B(n16356), .Z(n16369) );
  XNOR U16340 ( .A(n16399), .B(n16353), .Z(n16356) );
  XNOR U16341 ( .A(p_input[1434]), .B(p_input[2058]), .Z(n16353) );
  XOR U16342 ( .A(p_input[1435]), .B(n6319), .Z(n16399) );
  XOR U16343 ( .A(p_input[1436]), .B(p_input[2060]), .Z(n16357) );
  XOR U16344 ( .A(n16367), .B(n16400), .Z(n16398) );
  IV U16345 ( .A(n16358), .Z(n16400) );
  XOR U16346 ( .A(p_input[1425]), .B(p_input[2049]), .Z(n16358) );
  XNOR U16347 ( .A(n16401), .B(n16374), .Z(n16367) );
  XNOR U16348 ( .A(p_input[1439]), .B(n6322), .Z(n16374) );
  XOR U16349 ( .A(n16364), .B(n16373), .Z(n16401) );
  XOR U16350 ( .A(n16402), .B(n16370), .Z(n16373) );
  XOR U16351 ( .A(p_input[1437]), .B(p_input[2061]), .Z(n16370) );
  XOR U16352 ( .A(p_input[1438]), .B(n6324), .Z(n16402) );
  XOR U16353 ( .A(p_input[1433]), .B(p_input[2057]), .Z(n16364) );
  XOR U16354 ( .A(n16382), .B(n16380), .Z(n16362) );
  XNOR U16355 ( .A(n16403), .B(n16387), .Z(n16380) );
  XOR U16356 ( .A(p_input[1432]), .B(p_input[2056]), .Z(n16387) );
  XOR U16357 ( .A(n16377), .B(n16386), .Z(n16403) );
  XOR U16358 ( .A(n16404), .B(n16383), .Z(n16386) );
  XOR U16359 ( .A(p_input[1430]), .B(p_input[2054]), .Z(n16383) );
  XOR U16360 ( .A(p_input[1431]), .B(n7007), .Z(n16404) );
  XOR U16361 ( .A(p_input[1426]), .B(p_input[2050]), .Z(n16377) );
  XNOR U16362 ( .A(n16392), .B(n16391), .Z(n16382) );
  XOR U16363 ( .A(n16405), .B(n16388), .Z(n16391) );
  XOR U16364 ( .A(p_input[1427]), .B(p_input[2051]), .Z(n16388) );
  XOR U16365 ( .A(p_input[1428]), .B(n7009), .Z(n16405) );
  XOR U16366 ( .A(p_input[1429]), .B(p_input[2053]), .Z(n16392) );
  XOR U16367 ( .A(n16406), .B(n16407), .Z(n16291) );
  AND U16368 ( .A(n363), .B(n16408), .Z(n16407) );
  XNOR U16369 ( .A(n16409), .B(n16406), .Z(n16408) );
  XNOR U16370 ( .A(n16410), .B(n16411), .Z(n363) );
  AND U16371 ( .A(n16412), .B(n16413), .Z(n16411) );
  XOR U16372 ( .A(n16304), .B(n16410), .Z(n16413) );
  AND U16373 ( .A(n16414), .B(n16415), .Z(n16304) );
  XNOR U16374 ( .A(n16301), .B(n16410), .Z(n16412) );
  XOR U16375 ( .A(n16416), .B(n16417), .Z(n16301) );
  AND U16376 ( .A(n367), .B(n16418), .Z(n16417) );
  XOR U16377 ( .A(n16419), .B(n16416), .Z(n16418) );
  XOR U16378 ( .A(n16420), .B(n16421), .Z(n16410) );
  AND U16379 ( .A(n16422), .B(n16423), .Z(n16421) );
  XNOR U16380 ( .A(n16420), .B(n16414), .Z(n16423) );
  IV U16381 ( .A(n16319), .Z(n16414) );
  XOR U16382 ( .A(n16424), .B(n16425), .Z(n16319) );
  XOR U16383 ( .A(n16426), .B(n16415), .Z(n16425) );
  AND U16384 ( .A(n16346), .B(n16427), .Z(n16415) );
  AND U16385 ( .A(n16428), .B(n16429), .Z(n16426) );
  XOR U16386 ( .A(n16430), .B(n16424), .Z(n16428) );
  XNOR U16387 ( .A(n16316), .B(n16420), .Z(n16422) );
  XOR U16388 ( .A(n16431), .B(n16432), .Z(n16316) );
  AND U16389 ( .A(n367), .B(n16433), .Z(n16432) );
  XOR U16390 ( .A(n16434), .B(n16431), .Z(n16433) );
  XOR U16391 ( .A(n16435), .B(n16436), .Z(n16420) );
  AND U16392 ( .A(n16437), .B(n16438), .Z(n16436) );
  XNOR U16393 ( .A(n16435), .B(n16346), .Z(n16438) );
  XOR U16394 ( .A(n16439), .B(n16429), .Z(n16346) );
  XNOR U16395 ( .A(n16440), .B(n16424), .Z(n16429) );
  XOR U16396 ( .A(n16441), .B(n16442), .Z(n16424) );
  AND U16397 ( .A(n16443), .B(n16444), .Z(n16442) );
  XOR U16398 ( .A(n16445), .B(n16441), .Z(n16443) );
  XNOR U16399 ( .A(n16446), .B(n16447), .Z(n16440) );
  AND U16400 ( .A(n16448), .B(n16449), .Z(n16447) );
  XOR U16401 ( .A(n16446), .B(n16450), .Z(n16448) );
  XNOR U16402 ( .A(n16430), .B(n16427), .Z(n16439) );
  AND U16403 ( .A(n16451), .B(n16452), .Z(n16427) );
  XOR U16404 ( .A(n16453), .B(n16454), .Z(n16430) );
  AND U16405 ( .A(n16455), .B(n16456), .Z(n16454) );
  XOR U16406 ( .A(n16453), .B(n16457), .Z(n16455) );
  XNOR U16407 ( .A(n16343), .B(n16435), .Z(n16437) );
  XOR U16408 ( .A(n16458), .B(n16459), .Z(n16343) );
  AND U16409 ( .A(n367), .B(n16460), .Z(n16459) );
  XNOR U16410 ( .A(n16461), .B(n16458), .Z(n16460) );
  XOR U16411 ( .A(n16462), .B(n16463), .Z(n16435) );
  AND U16412 ( .A(n16464), .B(n16465), .Z(n16463) );
  XNOR U16413 ( .A(n16462), .B(n16451), .Z(n16465) );
  IV U16414 ( .A(n16396), .Z(n16451) );
  XNOR U16415 ( .A(n16466), .B(n16444), .Z(n16396) );
  XNOR U16416 ( .A(n16467), .B(n16450), .Z(n16444) );
  XNOR U16417 ( .A(n16468), .B(n16469), .Z(n16450) );
  NOR U16418 ( .A(n16470), .B(n16471), .Z(n16469) );
  XOR U16419 ( .A(n16468), .B(n16472), .Z(n16470) );
  XNOR U16420 ( .A(n16449), .B(n16441), .Z(n16467) );
  XOR U16421 ( .A(n16473), .B(n16474), .Z(n16441) );
  AND U16422 ( .A(n16475), .B(n16476), .Z(n16474) );
  XOR U16423 ( .A(n16473), .B(n16477), .Z(n16475) );
  XNOR U16424 ( .A(n16478), .B(n16446), .Z(n16449) );
  XOR U16425 ( .A(n16479), .B(n16480), .Z(n16446) );
  AND U16426 ( .A(n16481), .B(n16482), .Z(n16480) );
  XNOR U16427 ( .A(n16483), .B(n16484), .Z(n16481) );
  IV U16428 ( .A(n16479), .Z(n16483) );
  XNOR U16429 ( .A(n16485), .B(n16486), .Z(n16478) );
  NOR U16430 ( .A(n16487), .B(n16488), .Z(n16486) );
  XNOR U16431 ( .A(n16485), .B(n16489), .Z(n16487) );
  XNOR U16432 ( .A(n16445), .B(n16452), .Z(n16466) );
  NOR U16433 ( .A(n16409), .B(n16490), .Z(n16452) );
  XOR U16434 ( .A(n16457), .B(n16456), .Z(n16445) );
  XNOR U16435 ( .A(n16491), .B(n16453), .Z(n16456) );
  XOR U16436 ( .A(n16492), .B(n16493), .Z(n16453) );
  AND U16437 ( .A(n16494), .B(n16495), .Z(n16493) );
  XNOR U16438 ( .A(n16496), .B(n16497), .Z(n16494) );
  IV U16439 ( .A(n16492), .Z(n16496) );
  XNOR U16440 ( .A(n16498), .B(n16499), .Z(n16491) );
  NOR U16441 ( .A(n16500), .B(n16501), .Z(n16499) );
  XNOR U16442 ( .A(n16498), .B(n16502), .Z(n16500) );
  XOR U16443 ( .A(n16503), .B(n16504), .Z(n16457) );
  NOR U16444 ( .A(n16505), .B(n16506), .Z(n16504) );
  XNOR U16445 ( .A(n16503), .B(n16507), .Z(n16505) );
  XNOR U16446 ( .A(n16393), .B(n16462), .Z(n16464) );
  XOR U16447 ( .A(n16508), .B(n16509), .Z(n16393) );
  AND U16448 ( .A(n367), .B(n16510), .Z(n16509) );
  XOR U16449 ( .A(n16511), .B(n16508), .Z(n16510) );
  AND U16450 ( .A(n16406), .B(n16409), .Z(n16462) );
  XOR U16451 ( .A(n16512), .B(n16490), .Z(n16409) );
  XNOR U16452 ( .A(p_input[1440]), .B(p_input[2048]), .Z(n16490) );
  XNOR U16453 ( .A(n16477), .B(n16476), .Z(n16512) );
  XNOR U16454 ( .A(n16513), .B(n16484), .Z(n16476) );
  XNOR U16455 ( .A(n16472), .B(n16471), .Z(n16484) );
  XNOR U16456 ( .A(n16514), .B(n16468), .Z(n16471) );
  XNOR U16457 ( .A(p_input[1450]), .B(p_input[2058]), .Z(n16468) );
  XOR U16458 ( .A(p_input[1451]), .B(n6319), .Z(n16514) );
  XOR U16459 ( .A(p_input[1452]), .B(p_input[2060]), .Z(n16472) );
  XOR U16460 ( .A(n16482), .B(n16515), .Z(n16513) );
  IV U16461 ( .A(n16473), .Z(n16515) );
  XOR U16462 ( .A(p_input[1441]), .B(p_input[2049]), .Z(n16473) );
  XNOR U16463 ( .A(n16516), .B(n16489), .Z(n16482) );
  XNOR U16464 ( .A(p_input[1455]), .B(n6322), .Z(n16489) );
  XOR U16465 ( .A(n16479), .B(n16488), .Z(n16516) );
  XOR U16466 ( .A(n16517), .B(n16485), .Z(n16488) );
  XOR U16467 ( .A(p_input[1453]), .B(p_input[2061]), .Z(n16485) );
  XOR U16468 ( .A(p_input[1454]), .B(n6324), .Z(n16517) );
  XOR U16469 ( .A(p_input[1449]), .B(p_input[2057]), .Z(n16479) );
  XOR U16470 ( .A(n16497), .B(n16495), .Z(n16477) );
  XNOR U16471 ( .A(n16518), .B(n16502), .Z(n16495) );
  XOR U16472 ( .A(p_input[1448]), .B(p_input[2056]), .Z(n16502) );
  XOR U16473 ( .A(n16492), .B(n16501), .Z(n16518) );
  XOR U16474 ( .A(n16519), .B(n16498), .Z(n16501) );
  XOR U16475 ( .A(p_input[1446]), .B(p_input[2054]), .Z(n16498) );
  XOR U16476 ( .A(p_input[1447]), .B(n7007), .Z(n16519) );
  XOR U16477 ( .A(p_input[1442]), .B(p_input[2050]), .Z(n16492) );
  XNOR U16478 ( .A(n16507), .B(n16506), .Z(n16497) );
  XOR U16479 ( .A(n16520), .B(n16503), .Z(n16506) );
  XOR U16480 ( .A(p_input[1443]), .B(p_input[2051]), .Z(n16503) );
  XOR U16481 ( .A(p_input[1444]), .B(n7009), .Z(n16520) );
  XOR U16482 ( .A(p_input[1445]), .B(p_input[2053]), .Z(n16507) );
  XOR U16483 ( .A(n16521), .B(n16522), .Z(n16406) );
  AND U16484 ( .A(n367), .B(n16523), .Z(n16522) );
  XNOR U16485 ( .A(n16524), .B(n16521), .Z(n16523) );
  XNOR U16486 ( .A(n16525), .B(n16526), .Z(n367) );
  AND U16487 ( .A(n16527), .B(n16528), .Z(n16526) );
  XOR U16488 ( .A(n16419), .B(n16525), .Z(n16528) );
  AND U16489 ( .A(n16529), .B(n16530), .Z(n16419) );
  XNOR U16490 ( .A(n16416), .B(n16525), .Z(n16527) );
  XOR U16491 ( .A(n16531), .B(n16532), .Z(n16416) );
  AND U16492 ( .A(n371), .B(n16533), .Z(n16532) );
  XOR U16493 ( .A(n16534), .B(n16531), .Z(n16533) );
  XOR U16494 ( .A(n16535), .B(n16536), .Z(n16525) );
  AND U16495 ( .A(n16537), .B(n16538), .Z(n16536) );
  XNOR U16496 ( .A(n16535), .B(n16529), .Z(n16538) );
  IV U16497 ( .A(n16434), .Z(n16529) );
  XOR U16498 ( .A(n16539), .B(n16540), .Z(n16434) );
  XOR U16499 ( .A(n16541), .B(n16530), .Z(n16540) );
  AND U16500 ( .A(n16461), .B(n16542), .Z(n16530) );
  AND U16501 ( .A(n16543), .B(n16544), .Z(n16541) );
  XOR U16502 ( .A(n16545), .B(n16539), .Z(n16543) );
  XNOR U16503 ( .A(n16431), .B(n16535), .Z(n16537) );
  XOR U16504 ( .A(n16546), .B(n16547), .Z(n16431) );
  AND U16505 ( .A(n371), .B(n16548), .Z(n16547) );
  XOR U16506 ( .A(n16549), .B(n16546), .Z(n16548) );
  XOR U16507 ( .A(n16550), .B(n16551), .Z(n16535) );
  AND U16508 ( .A(n16552), .B(n16553), .Z(n16551) );
  XNOR U16509 ( .A(n16550), .B(n16461), .Z(n16553) );
  XOR U16510 ( .A(n16554), .B(n16544), .Z(n16461) );
  XNOR U16511 ( .A(n16555), .B(n16539), .Z(n16544) );
  XOR U16512 ( .A(n16556), .B(n16557), .Z(n16539) );
  AND U16513 ( .A(n16558), .B(n16559), .Z(n16557) );
  XOR U16514 ( .A(n16560), .B(n16556), .Z(n16558) );
  XNOR U16515 ( .A(n16561), .B(n16562), .Z(n16555) );
  AND U16516 ( .A(n16563), .B(n16564), .Z(n16562) );
  XOR U16517 ( .A(n16561), .B(n16565), .Z(n16563) );
  XNOR U16518 ( .A(n16545), .B(n16542), .Z(n16554) );
  AND U16519 ( .A(n16566), .B(n16567), .Z(n16542) );
  XOR U16520 ( .A(n16568), .B(n16569), .Z(n16545) );
  AND U16521 ( .A(n16570), .B(n16571), .Z(n16569) );
  XOR U16522 ( .A(n16568), .B(n16572), .Z(n16570) );
  XNOR U16523 ( .A(n16458), .B(n16550), .Z(n16552) );
  XOR U16524 ( .A(n16573), .B(n16574), .Z(n16458) );
  AND U16525 ( .A(n371), .B(n16575), .Z(n16574) );
  XNOR U16526 ( .A(n16576), .B(n16573), .Z(n16575) );
  XOR U16527 ( .A(n16577), .B(n16578), .Z(n16550) );
  AND U16528 ( .A(n16579), .B(n16580), .Z(n16578) );
  XNOR U16529 ( .A(n16577), .B(n16566), .Z(n16580) );
  IV U16530 ( .A(n16511), .Z(n16566) );
  XNOR U16531 ( .A(n16581), .B(n16559), .Z(n16511) );
  XNOR U16532 ( .A(n16582), .B(n16565), .Z(n16559) );
  XNOR U16533 ( .A(n16583), .B(n16584), .Z(n16565) );
  NOR U16534 ( .A(n16585), .B(n16586), .Z(n16584) );
  XOR U16535 ( .A(n16583), .B(n16587), .Z(n16585) );
  XNOR U16536 ( .A(n16564), .B(n16556), .Z(n16582) );
  XOR U16537 ( .A(n16588), .B(n16589), .Z(n16556) );
  AND U16538 ( .A(n16590), .B(n16591), .Z(n16589) );
  XOR U16539 ( .A(n16588), .B(n16592), .Z(n16590) );
  XNOR U16540 ( .A(n16593), .B(n16561), .Z(n16564) );
  XOR U16541 ( .A(n16594), .B(n16595), .Z(n16561) );
  AND U16542 ( .A(n16596), .B(n16597), .Z(n16595) );
  XNOR U16543 ( .A(n16598), .B(n16599), .Z(n16596) );
  IV U16544 ( .A(n16594), .Z(n16598) );
  XNOR U16545 ( .A(n16600), .B(n16601), .Z(n16593) );
  NOR U16546 ( .A(n16602), .B(n16603), .Z(n16601) );
  XNOR U16547 ( .A(n16600), .B(n16604), .Z(n16602) );
  XNOR U16548 ( .A(n16560), .B(n16567), .Z(n16581) );
  NOR U16549 ( .A(n16524), .B(n16605), .Z(n16567) );
  XOR U16550 ( .A(n16572), .B(n16571), .Z(n16560) );
  XNOR U16551 ( .A(n16606), .B(n16568), .Z(n16571) );
  XOR U16552 ( .A(n16607), .B(n16608), .Z(n16568) );
  AND U16553 ( .A(n16609), .B(n16610), .Z(n16608) );
  XNOR U16554 ( .A(n16611), .B(n16612), .Z(n16609) );
  IV U16555 ( .A(n16607), .Z(n16611) );
  XNOR U16556 ( .A(n16613), .B(n16614), .Z(n16606) );
  NOR U16557 ( .A(n16615), .B(n16616), .Z(n16614) );
  XNOR U16558 ( .A(n16613), .B(n16617), .Z(n16615) );
  XOR U16559 ( .A(n16618), .B(n16619), .Z(n16572) );
  NOR U16560 ( .A(n16620), .B(n16621), .Z(n16619) );
  XNOR U16561 ( .A(n16618), .B(n16622), .Z(n16620) );
  XNOR U16562 ( .A(n16508), .B(n16577), .Z(n16579) );
  XOR U16563 ( .A(n16623), .B(n16624), .Z(n16508) );
  AND U16564 ( .A(n371), .B(n16625), .Z(n16624) );
  XOR U16565 ( .A(n16626), .B(n16623), .Z(n16625) );
  AND U16566 ( .A(n16521), .B(n16524), .Z(n16577) );
  XOR U16567 ( .A(n16627), .B(n16605), .Z(n16524) );
  XNOR U16568 ( .A(p_input[1456]), .B(p_input[2048]), .Z(n16605) );
  XNOR U16569 ( .A(n16592), .B(n16591), .Z(n16627) );
  XNOR U16570 ( .A(n16628), .B(n16599), .Z(n16591) );
  XNOR U16571 ( .A(n16587), .B(n16586), .Z(n16599) );
  XNOR U16572 ( .A(n16629), .B(n16583), .Z(n16586) );
  XNOR U16573 ( .A(p_input[1466]), .B(p_input[2058]), .Z(n16583) );
  XOR U16574 ( .A(p_input[1467]), .B(n6319), .Z(n16629) );
  XOR U16575 ( .A(p_input[1468]), .B(p_input[2060]), .Z(n16587) );
  XOR U16576 ( .A(n16597), .B(n16630), .Z(n16628) );
  IV U16577 ( .A(n16588), .Z(n16630) );
  XOR U16578 ( .A(p_input[1457]), .B(p_input[2049]), .Z(n16588) );
  XNOR U16579 ( .A(n16631), .B(n16604), .Z(n16597) );
  XNOR U16580 ( .A(p_input[1471]), .B(n6322), .Z(n16604) );
  XOR U16581 ( .A(n16594), .B(n16603), .Z(n16631) );
  XOR U16582 ( .A(n16632), .B(n16600), .Z(n16603) );
  XOR U16583 ( .A(p_input[1469]), .B(p_input[2061]), .Z(n16600) );
  XOR U16584 ( .A(p_input[1470]), .B(n6324), .Z(n16632) );
  XOR U16585 ( .A(p_input[1465]), .B(p_input[2057]), .Z(n16594) );
  XOR U16586 ( .A(n16612), .B(n16610), .Z(n16592) );
  XNOR U16587 ( .A(n16633), .B(n16617), .Z(n16610) );
  XOR U16588 ( .A(p_input[1464]), .B(p_input[2056]), .Z(n16617) );
  XOR U16589 ( .A(n16607), .B(n16616), .Z(n16633) );
  XOR U16590 ( .A(n16634), .B(n16613), .Z(n16616) );
  XOR U16591 ( .A(p_input[1462]), .B(p_input[2054]), .Z(n16613) );
  XOR U16592 ( .A(p_input[1463]), .B(n7007), .Z(n16634) );
  XOR U16593 ( .A(p_input[1458]), .B(p_input[2050]), .Z(n16607) );
  XNOR U16594 ( .A(n16622), .B(n16621), .Z(n16612) );
  XOR U16595 ( .A(n16635), .B(n16618), .Z(n16621) );
  XOR U16596 ( .A(p_input[1459]), .B(p_input[2051]), .Z(n16618) );
  XOR U16597 ( .A(p_input[1460]), .B(n7009), .Z(n16635) );
  XOR U16598 ( .A(p_input[1461]), .B(p_input[2053]), .Z(n16622) );
  XOR U16599 ( .A(n16636), .B(n16637), .Z(n16521) );
  AND U16600 ( .A(n371), .B(n16638), .Z(n16637) );
  XNOR U16601 ( .A(n16639), .B(n16636), .Z(n16638) );
  XNOR U16602 ( .A(n16640), .B(n16641), .Z(n371) );
  AND U16603 ( .A(n16642), .B(n16643), .Z(n16641) );
  XOR U16604 ( .A(n16534), .B(n16640), .Z(n16643) );
  AND U16605 ( .A(n16644), .B(n16645), .Z(n16534) );
  XNOR U16606 ( .A(n16531), .B(n16640), .Z(n16642) );
  XOR U16607 ( .A(n16646), .B(n16647), .Z(n16531) );
  AND U16608 ( .A(n375), .B(n16648), .Z(n16647) );
  XOR U16609 ( .A(n16649), .B(n16646), .Z(n16648) );
  XOR U16610 ( .A(n16650), .B(n16651), .Z(n16640) );
  AND U16611 ( .A(n16652), .B(n16653), .Z(n16651) );
  XNOR U16612 ( .A(n16650), .B(n16644), .Z(n16653) );
  IV U16613 ( .A(n16549), .Z(n16644) );
  XOR U16614 ( .A(n16654), .B(n16655), .Z(n16549) );
  XOR U16615 ( .A(n16656), .B(n16645), .Z(n16655) );
  AND U16616 ( .A(n16576), .B(n16657), .Z(n16645) );
  AND U16617 ( .A(n16658), .B(n16659), .Z(n16656) );
  XOR U16618 ( .A(n16660), .B(n16654), .Z(n16658) );
  XNOR U16619 ( .A(n16546), .B(n16650), .Z(n16652) );
  XOR U16620 ( .A(n16661), .B(n16662), .Z(n16546) );
  AND U16621 ( .A(n375), .B(n16663), .Z(n16662) );
  XOR U16622 ( .A(n16664), .B(n16661), .Z(n16663) );
  XOR U16623 ( .A(n16665), .B(n16666), .Z(n16650) );
  AND U16624 ( .A(n16667), .B(n16668), .Z(n16666) );
  XNOR U16625 ( .A(n16665), .B(n16576), .Z(n16668) );
  XOR U16626 ( .A(n16669), .B(n16659), .Z(n16576) );
  XNOR U16627 ( .A(n16670), .B(n16654), .Z(n16659) );
  XOR U16628 ( .A(n16671), .B(n16672), .Z(n16654) );
  AND U16629 ( .A(n16673), .B(n16674), .Z(n16672) );
  XOR U16630 ( .A(n16675), .B(n16671), .Z(n16673) );
  XNOR U16631 ( .A(n16676), .B(n16677), .Z(n16670) );
  AND U16632 ( .A(n16678), .B(n16679), .Z(n16677) );
  XOR U16633 ( .A(n16676), .B(n16680), .Z(n16678) );
  XNOR U16634 ( .A(n16660), .B(n16657), .Z(n16669) );
  AND U16635 ( .A(n16681), .B(n16682), .Z(n16657) );
  XOR U16636 ( .A(n16683), .B(n16684), .Z(n16660) );
  AND U16637 ( .A(n16685), .B(n16686), .Z(n16684) );
  XOR U16638 ( .A(n16683), .B(n16687), .Z(n16685) );
  XNOR U16639 ( .A(n16573), .B(n16665), .Z(n16667) );
  XOR U16640 ( .A(n16688), .B(n16689), .Z(n16573) );
  AND U16641 ( .A(n375), .B(n16690), .Z(n16689) );
  XNOR U16642 ( .A(n16691), .B(n16688), .Z(n16690) );
  XOR U16643 ( .A(n16692), .B(n16693), .Z(n16665) );
  AND U16644 ( .A(n16694), .B(n16695), .Z(n16693) );
  XNOR U16645 ( .A(n16692), .B(n16681), .Z(n16695) );
  IV U16646 ( .A(n16626), .Z(n16681) );
  XNOR U16647 ( .A(n16696), .B(n16674), .Z(n16626) );
  XNOR U16648 ( .A(n16697), .B(n16680), .Z(n16674) );
  XNOR U16649 ( .A(n16698), .B(n16699), .Z(n16680) );
  NOR U16650 ( .A(n16700), .B(n16701), .Z(n16699) );
  XOR U16651 ( .A(n16698), .B(n16702), .Z(n16700) );
  XNOR U16652 ( .A(n16679), .B(n16671), .Z(n16697) );
  XOR U16653 ( .A(n16703), .B(n16704), .Z(n16671) );
  AND U16654 ( .A(n16705), .B(n16706), .Z(n16704) );
  XOR U16655 ( .A(n16703), .B(n16707), .Z(n16705) );
  XNOR U16656 ( .A(n16708), .B(n16676), .Z(n16679) );
  XOR U16657 ( .A(n16709), .B(n16710), .Z(n16676) );
  AND U16658 ( .A(n16711), .B(n16712), .Z(n16710) );
  XNOR U16659 ( .A(n16713), .B(n16714), .Z(n16711) );
  IV U16660 ( .A(n16709), .Z(n16713) );
  XNOR U16661 ( .A(n16715), .B(n16716), .Z(n16708) );
  NOR U16662 ( .A(n16717), .B(n16718), .Z(n16716) );
  XNOR U16663 ( .A(n16715), .B(n16719), .Z(n16717) );
  XNOR U16664 ( .A(n16675), .B(n16682), .Z(n16696) );
  NOR U16665 ( .A(n16639), .B(n16720), .Z(n16682) );
  XOR U16666 ( .A(n16687), .B(n16686), .Z(n16675) );
  XNOR U16667 ( .A(n16721), .B(n16683), .Z(n16686) );
  XOR U16668 ( .A(n16722), .B(n16723), .Z(n16683) );
  AND U16669 ( .A(n16724), .B(n16725), .Z(n16723) );
  XNOR U16670 ( .A(n16726), .B(n16727), .Z(n16724) );
  IV U16671 ( .A(n16722), .Z(n16726) );
  XNOR U16672 ( .A(n16728), .B(n16729), .Z(n16721) );
  NOR U16673 ( .A(n16730), .B(n16731), .Z(n16729) );
  XNOR U16674 ( .A(n16728), .B(n16732), .Z(n16730) );
  XOR U16675 ( .A(n16733), .B(n16734), .Z(n16687) );
  NOR U16676 ( .A(n16735), .B(n16736), .Z(n16734) );
  XNOR U16677 ( .A(n16733), .B(n16737), .Z(n16735) );
  XNOR U16678 ( .A(n16623), .B(n16692), .Z(n16694) );
  XOR U16679 ( .A(n16738), .B(n16739), .Z(n16623) );
  AND U16680 ( .A(n375), .B(n16740), .Z(n16739) );
  XOR U16681 ( .A(n16741), .B(n16738), .Z(n16740) );
  AND U16682 ( .A(n16636), .B(n16639), .Z(n16692) );
  XOR U16683 ( .A(n16742), .B(n16720), .Z(n16639) );
  XNOR U16684 ( .A(p_input[1472]), .B(p_input[2048]), .Z(n16720) );
  XNOR U16685 ( .A(n16707), .B(n16706), .Z(n16742) );
  XNOR U16686 ( .A(n16743), .B(n16714), .Z(n16706) );
  XNOR U16687 ( .A(n16702), .B(n16701), .Z(n16714) );
  XNOR U16688 ( .A(n16744), .B(n16698), .Z(n16701) );
  XNOR U16689 ( .A(p_input[1482]), .B(p_input[2058]), .Z(n16698) );
  XOR U16690 ( .A(p_input[1483]), .B(n6319), .Z(n16744) );
  XOR U16691 ( .A(p_input[1484]), .B(p_input[2060]), .Z(n16702) );
  XOR U16692 ( .A(n16712), .B(n16745), .Z(n16743) );
  IV U16693 ( .A(n16703), .Z(n16745) );
  XOR U16694 ( .A(p_input[1473]), .B(p_input[2049]), .Z(n16703) );
  XNOR U16695 ( .A(n16746), .B(n16719), .Z(n16712) );
  XNOR U16696 ( .A(p_input[1487]), .B(n6322), .Z(n16719) );
  XOR U16697 ( .A(n16709), .B(n16718), .Z(n16746) );
  XOR U16698 ( .A(n16747), .B(n16715), .Z(n16718) );
  XOR U16699 ( .A(p_input[1485]), .B(p_input[2061]), .Z(n16715) );
  XOR U16700 ( .A(p_input[1486]), .B(n6324), .Z(n16747) );
  XOR U16701 ( .A(p_input[1481]), .B(p_input[2057]), .Z(n16709) );
  XOR U16702 ( .A(n16727), .B(n16725), .Z(n16707) );
  XNOR U16703 ( .A(n16748), .B(n16732), .Z(n16725) );
  XOR U16704 ( .A(p_input[1480]), .B(p_input[2056]), .Z(n16732) );
  XOR U16705 ( .A(n16722), .B(n16731), .Z(n16748) );
  XOR U16706 ( .A(n16749), .B(n16728), .Z(n16731) );
  XOR U16707 ( .A(p_input[1478]), .B(p_input[2054]), .Z(n16728) );
  XOR U16708 ( .A(p_input[1479]), .B(n7007), .Z(n16749) );
  XOR U16709 ( .A(p_input[1474]), .B(p_input[2050]), .Z(n16722) );
  XNOR U16710 ( .A(n16737), .B(n16736), .Z(n16727) );
  XOR U16711 ( .A(n16750), .B(n16733), .Z(n16736) );
  XOR U16712 ( .A(p_input[1475]), .B(p_input[2051]), .Z(n16733) );
  XOR U16713 ( .A(p_input[1476]), .B(n7009), .Z(n16750) );
  XOR U16714 ( .A(p_input[1477]), .B(p_input[2053]), .Z(n16737) );
  XOR U16715 ( .A(n16751), .B(n16752), .Z(n16636) );
  AND U16716 ( .A(n375), .B(n16753), .Z(n16752) );
  XNOR U16717 ( .A(n16754), .B(n16751), .Z(n16753) );
  XNOR U16718 ( .A(n16755), .B(n16756), .Z(n375) );
  AND U16719 ( .A(n16757), .B(n16758), .Z(n16756) );
  XOR U16720 ( .A(n16649), .B(n16755), .Z(n16758) );
  AND U16721 ( .A(n16759), .B(n16760), .Z(n16649) );
  XNOR U16722 ( .A(n16646), .B(n16755), .Z(n16757) );
  XOR U16723 ( .A(n16761), .B(n16762), .Z(n16646) );
  AND U16724 ( .A(n379), .B(n16763), .Z(n16762) );
  XOR U16725 ( .A(n16764), .B(n16761), .Z(n16763) );
  XOR U16726 ( .A(n16765), .B(n16766), .Z(n16755) );
  AND U16727 ( .A(n16767), .B(n16768), .Z(n16766) );
  XNOR U16728 ( .A(n16765), .B(n16759), .Z(n16768) );
  IV U16729 ( .A(n16664), .Z(n16759) );
  XOR U16730 ( .A(n16769), .B(n16770), .Z(n16664) );
  XOR U16731 ( .A(n16771), .B(n16760), .Z(n16770) );
  AND U16732 ( .A(n16691), .B(n16772), .Z(n16760) );
  AND U16733 ( .A(n16773), .B(n16774), .Z(n16771) );
  XOR U16734 ( .A(n16775), .B(n16769), .Z(n16773) );
  XNOR U16735 ( .A(n16661), .B(n16765), .Z(n16767) );
  XOR U16736 ( .A(n16776), .B(n16777), .Z(n16661) );
  AND U16737 ( .A(n379), .B(n16778), .Z(n16777) );
  XOR U16738 ( .A(n16779), .B(n16776), .Z(n16778) );
  XOR U16739 ( .A(n16780), .B(n16781), .Z(n16765) );
  AND U16740 ( .A(n16782), .B(n16783), .Z(n16781) );
  XNOR U16741 ( .A(n16780), .B(n16691), .Z(n16783) );
  XOR U16742 ( .A(n16784), .B(n16774), .Z(n16691) );
  XNOR U16743 ( .A(n16785), .B(n16769), .Z(n16774) );
  XOR U16744 ( .A(n16786), .B(n16787), .Z(n16769) );
  AND U16745 ( .A(n16788), .B(n16789), .Z(n16787) );
  XOR U16746 ( .A(n16790), .B(n16786), .Z(n16788) );
  XNOR U16747 ( .A(n16791), .B(n16792), .Z(n16785) );
  AND U16748 ( .A(n16793), .B(n16794), .Z(n16792) );
  XOR U16749 ( .A(n16791), .B(n16795), .Z(n16793) );
  XNOR U16750 ( .A(n16775), .B(n16772), .Z(n16784) );
  AND U16751 ( .A(n16796), .B(n16797), .Z(n16772) );
  XOR U16752 ( .A(n16798), .B(n16799), .Z(n16775) );
  AND U16753 ( .A(n16800), .B(n16801), .Z(n16799) );
  XOR U16754 ( .A(n16798), .B(n16802), .Z(n16800) );
  XNOR U16755 ( .A(n16688), .B(n16780), .Z(n16782) );
  XOR U16756 ( .A(n16803), .B(n16804), .Z(n16688) );
  AND U16757 ( .A(n379), .B(n16805), .Z(n16804) );
  XNOR U16758 ( .A(n16806), .B(n16803), .Z(n16805) );
  XOR U16759 ( .A(n16807), .B(n16808), .Z(n16780) );
  AND U16760 ( .A(n16809), .B(n16810), .Z(n16808) );
  XNOR U16761 ( .A(n16807), .B(n16796), .Z(n16810) );
  IV U16762 ( .A(n16741), .Z(n16796) );
  XNOR U16763 ( .A(n16811), .B(n16789), .Z(n16741) );
  XNOR U16764 ( .A(n16812), .B(n16795), .Z(n16789) );
  XNOR U16765 ( .A(n16813), .B(n16814), .Z(n16795) );
  NOR U16766 ( .A(n16815), .B(n16816), .Z(n16814) );
  XOR U16767 ( .A(n16813), .B(n16817), .Z(n16815) );
  XNOR U16768 ( .A(n16794), .B(n16786), .Z(n16812) );
  XOR U16769 ( .A(n16818), .B(n16819), .Z(n16786) );
  AND U16770 ( .A(n16820), .B(n16821), .Z(n16819) );
  XOR U16771 ( .A(n16818), .B(n16822), .Z(n16820) );
  XNOR U16772 ( .A(n16823), .B(n16791), .Z(n16794) );
  XOR U16773 ( .A(n16824), .B(n16825), .Z(n16791) );
  AND U16774 ( .A(n16826), .B(n16827), .Z(n16825) );
  XNOR U16775 ( .A(n16828), .B(n16829), .Z(n16826) );
  IV U16776 ( .A(n16824), .Z(n16828) );
  XNOR U16777 ( .A(n16830), .B(n16831), .Z(n16823) );
  NOR U16778 ( .A(n16832), .B(n16833), .Z(n16831) );
  XNOR U16779 ( .A(n16830), .B(n16834), .Z(n16832) );
  XNOR U16780 ( .A(n16790), .B(n16797), .Z(n16811) );
  NOR U16781 ( .A(n16754), .B(n16835), .Z(n16797) );
  XOR U16782 ( .A(n16802), .B(n16801), .Z(n16790) );
  XNOR U16783 ( .A(n16836), .B(n16798), .Z(n16801) );
  XOR U16784 ( .A(n16837), .B(n16838), .Z(n16798) );
  AND U16785 ( .A(n16839), .B(n16840), .Z(n16838) );
  XNOR U16786 ( .A(n16841), .B(n16842), .Z(n16839) );
  IV U16787 ( .A(n16837), .Z(n16841) );
  XNOR U16788 ( .A(n16843), .B(n16844), .Z(n16836) );
  NOR U16789 ( .A(n16845), .B(n16846), .Z(n16844) );
  XNOR U16790 ( .A(n16843), .B(n16847), .Z(n16845) );
  XOR U16791 ( .A(n16848), .B(n16849), .Z(n16802) );
  NOR U16792 ( .A(n16850), .B(n16851), .Z(n16849) );
  XNOR U16793 ( .A(n16848), .B(n16852), .Z(n16850) );
  XNOR U16794 ( .A(n16738), .B(n16807), .Z(n16809) );
  XOR U16795 ( .A(n16853), .B(n16854), .Z(n16738) );
  AND U16796 ( .A(n379), .B(n16855), .Z(n16854) );
  XOR U16797 ( .A(n16856), .B(n16853), .Z(n16855) );
  AND U16798 ( .A(n16751), .B(n16754), .Z(n16807) );
  XOR U16799 ( .A(n16857), .B(n16835), .Z(n16754) );
  XNOR U16800 ( .A(p_input[1488]), .B(p_input[2048]), .Z(n16835) );
  XNOR U16801 ( .A(n16822), .B(n16821), .Z(n16857) );
  XNOR U16802 ( .A(n16858), .B(n16829), .Z(n16821) );
  XNOR U16803 ( .A(n16817), .B(n16816), .Z(n16829) );
  XNOR U16804 ( .A(n16859), .B(n16813), .Z(n16816) );
  XNOR U16805 ( .A(p_input[1498]), .B(p_input[2058]), .Z(n16813) );
  XOR U16806 ( .A(p_input[1499]), .B(n6319), .Z(n16859) );
  XOR U16807 ( .A(p_input[1500]), .B(p_input[2060]), .Z(n16817) );
  XOR U16808 ( .A(n16827), .B(n16860), .Z(n16858) );
  IV U16809 ( .A(n16818), .Z(n16860) );
  XOR U16810 ( .A(p_input[1489]), .B(p_input[2049]), .Z(n16818) );
  XNOR U16811 ( .A(n16861), .B(n16834), .Z(n16827) );
  XNOR U16812 ( .A(p_input[1503]), .B(n6322), .Z(n16834) );
  XOR U16813 ( .A(n16824), .B(n16833), .Z(n16861) );
  XOR U16814 ( .A(n16862), .B(n16830), .Z(n16833) );
  XOR U16815 ( .A(p_input[1501]), .B(p_input[2061]), .Z(n16830) );
  XOR U16816 ( .A(p_input[1502]), .B(n6324), .Z(n16862) );
  XOR U16817 ( .A(p_input[1497]), .B(p_input[2057]), .Z(n16824) );
  XOR U16818 ( .A(n16842), .B(n16840), .Z(n16822) );
  XNOR U16819 ( .A(n16863), .B(n16847), .Z(n16840) );
  XOR U16820 ( .A(p_input[1496]), .B(p_input[2056]), .Z(n16847) );
  XOR U16821 ( .A(n16837), .B(n16846), .Z(n16863) );
  XOR U16822 ( .A(n16864), .B(n16843), .Z(n16846) );
  XOR U16823 ( .A(p_input[1494]), .B(p_input[2054]), .Z(n16843) );
  XOR U16824 ( .A(p_input[1495]), .B(n7007), .Z(n16864) );
  XOR U16825 ( .A(p_input[1490]), .B(p_input[2050]), .Z(n16837) );
  XNOR U16826 ( .A(n16852), .B(n16851), .Z(n16842) );
  XOR U16827 ( .A(n16865), .B(n16848), .Z(n16851) );
  XOR U16828 ( .A(p_input[1491]), .B(p_input[2051]), .Z(n16848) );
  XOR U16829 ( .A(p_input[1492]), .B(n7009), .Z(n16865) );
  XOR U16830 ( .A(p_input[1493]), .B(p_input[2053]), .Z(n16852) );
  XOR U16831 ( .A(n16866), .B(n16867), .Z(n16751) );
  AND U16832 ( .A(n379), .B(n16868), .Z(n16867) );
  XNOR U16833 ( .A(n16869), .B(n16866), .Z(n16868) );
  XNOR U16834 ( .A(n16870), .B(n16871), .Z(n379) );
  AND U16835 ( .A(n16872), .B(n16873), .Z(n16871) );
  XOR U16836 ( .A(n16764), .B(n16870), .Z(n16873) );
  AND U16837 ( .A(n16874), .B(n16875), .Z(n16764) );
  XNOR U16838 ( .A(n16761), .B(n16870), .Z(n16872) );
  XOR U16839 ( .A(n16876), .B(n16877), .Z(n16761) );
  AND U16840 ( .A(n383), .B(n16878), .Z(n16877) );
  XOR U16841 ( .A(n16879), .B(n16876), .Z(n16878) );
  XOR U16842 ( .A(n16880), .B(n16881), .Z(n16870) );
  AND U16843 ( .A(n16882), .B(n16883), .Z(n16881) );
  XNOR U16844 ( .A(n16880), .B(n16874), .Z(n16883) );
  IV U16845 ( .A(n16779), .Z(n16874) );
  XOR U16846 ( .A(n16884), .B(n16885), .Z(n16779) );
  XOR U16847 ( .A(n16886), .B(n16875), .Z(n16885) );
  AND U16848 ( .A(n16806), .B(n16887), .Z(n16875) );
  AND U16849 ( .A(n16888), .B(n16889), .Z(n16886) );
  XOR U16850 ( .A(n16890), .B(n16884), .Z(n16888) );
  XNOR U16851 ( .A(n16776), .B(n16880), .Z(n16882) );
  XOR U16852 ( .A(n16891), .B(n16892), .Z(n16776) );
  AND U16853 ( .A(n383), .B(n16893), .Z(n16892) );
  XOR U16854 ( .A(n16894), .B(n16891), .Z(n16893) );
  XOR U16855 ( .A(n16895), .B(n16896), .Z(n16880) );
  AND U16856 ( .A(n16897), .B(n16898), .Z(n16896) );
  XNOR U16857 ( .A(n16895), .B(n16806), .Z(n16898) );
  XOR U16858 ( .A(n16899), .B(n16889), .Z(n16806) );
  XNOR U16859 ( .A(n16900), .B(n16884), .Z(n16889) );
  XOR U16860 ( .A(n16901), .B(n16902), .Z(n16884) );
  AND U16861 ( .A(n16903), .B(n16904), .Z(n16902) );
  XOR U16862 ( .A(n16905), .B(n16901), .Z(n16903) );
  XNOR U16863 ( .A(n16906), .B(n16907), .Z(n16900) );
  AND U16864 ( .A(n16908), .B(n16909), .Z(n16907) );
  XOR U16865 ( .A(n16906), .B(n16910), .Z(n16908) );
  XNOR U16866 ( .A(n16890), .B(n16887), .Z(n16899) );
  AND U16867 ( .A(n16911), .B(n16912), .Z(n16887) );
  XOR U16868 ( .A(n16913), .B(n16914), .Z(n16890) );
  AND U16869 ( .A(n16915), .B(n16916), .Z(n16914) );
  XOR U16870 ( .A(n16913), .B(n16917), .Z(n16915) );
  XNOR U16871 ( .A(n16803), .B(n16895), .Z(n16897) );
  XOR U16872 ( .A(n16918), .B(n16919), .Z(n16803) );
  AND U16873 ( .A(n383), .B(n16920), .Z(n16919) );
  XNOR U16874 ( .A(n16921), .B(n16918), .Z(n16920) );
  XOR U16875 ( .A(n16922), .B(n16923), .Z(n16895) );
  AND U16876 ( .A(n16924), .B(n16925), .Z(n16923) );
  XNOR U16877 ( .A(n16922), .B(n16911), .Z(n16925) );
  IV U16878 ( .A(n16856), .Z(n16911) );
  XNOR U16879 ( .A(n16926), .B(n16904), .Z(n16856) );
  XNOR U16880 ( .A(n16927), .B(n16910), .Z(n16904) );
  XNOR U16881 ( .A(n16928), .B(n16929), .Z(n16910) );
  NOR U16882 ( .A(n16930), .B(n16931), .Z(n16929) );
  XOR U16883 ( .A(n16928), .B(n16932), .Z(n16930) );
  XNOR U16884 ( .A(n16909), .B(n16901), .Z(n16927) );
  XOR U16885 ( .A(n16933), .B(n16934), .Z(n16901) );
  AND U16886 ( .A(n16935), .B(n16936), .Z(n16934) );
  XOR U16887 ( .A(n16933), .B(n16937), .Z(n16935) );
  XNOR U16888 ( .A(n16938), .B(n16906), .Z(n16909) );
  XOR U16889 ( .A(n16939), .B(n16940), .Z(n16906) );
  AND U16890 ( .A(n16941), .B(n16942), .Z(n16940) );
  XNOR U16891 ( .A(n16943), .B(n16944), .Z(n16941) );
  IV U16892 ( .A(n16939), .Z(n16943) );
  XNOR U16893 ( .A(n16945), .B(n16946), .Z(n16938) );
  NOR U16894 ( .A(n16947), .B(n16948), .Z(n16946) );
  XNOR U16895 ( .A(n16945), .B(n16949), .Z(n16947) );
  XNOR U16896 ( .A(n16905), .B(n16912), .Z(n16926) );
  NOR U16897 ( .A(n16869), .B(n16950), .Z(n16912) );
  XOR U16898 ( .A(n16917), .B(n16916), .Z(n16905) );
  XNOR U16899 ( .A(n16951), .B(n16913), .Z(n16916) );
  XOR U16900 ( .A(n16952), .B(n16953), .Z(n16913) );
  AND U16901 ( .A(n16954), .B(n16955), .Z(n16953) );
  XNOR U16902 ( .A(n16956), .B(n16957), .Z(n16954) );
  IV U16903 ( .A(n16952), .Z(n16956) );
  XNOR U16904 ( .A(n16958), .B(n16959), .Z(n16951) );
  NOR U16905 ( .A(n16960), .B(n16961), .Z(n16959) );
  XNOR U16906 ( .A(n16958), .B(n16962), .Z(n16960) );
  XOR U16907 ( .A(n16963), .B(n16964), .Z(n16917) );
  NOR U16908 ( .A(n16965), .B(n16966), .Z(n16964) );
  XNOR U16909 ( .A(n16963), .B(n16967), .Z(n16965) );
  XNOR U16910 ( .A(n16853), .B(n16922), .Z(n16924) );
  XOR U16911 ( .A(n16968), .B(n16969), .Z(n16853) );
  AND U16912 ( .A(n383), .B(n16970), .Z(n16969) );
  XOR U16913 ( .A(n16971), .B(n16968), .Z(n16970) );
  AND U16914 ( .A(n16866), .B(n16869), .Z(n16922) );
  XOR U16915 ( .A(n16972), .B(n16950), .Z(n16869) );
  XNOR U16916 ( .A(p_input[1504]), .B(p_input[2048]), .Z(n16950) );
  XNOR U16917 ( .A(n16937), .B(n16936), .Z(n16972) );
  XNOR U16918 ( .A(n16973), .B(n16944), .Z(n16936) );
  XNOR U16919 ( .A(n16932), .B(n16931), .Z(n16944) );
  XNOR U16920 ( .A(n16974), .B(n16928), .Z(n16931) );
  XNOR U16921 ( .A(p_input[1514]), .B(p_input[2058]), .Z(n16928) );
  XOR U16922 ( .A(p_input[1515]), .B(n6319), .Z(n16974) );
  XOR U16923 ( .A(p_input[1516]), .B(p_input[2060]), .Z(n16932) );
  XOR U16924 ( .A(n16942), .B(n16975), .Z(n16973) );
  IV U16925 ( .A(n16933), .Z(n16975) );
  XOR U16926 ( .A(p_input[1505]), .B(p_input[2049]), .Z(n16933) );
  XNOR U16927 ( .A(n16976), .B(n16949), .Z(n16942) );
  XNOR U16928 ( .A(p_input[1519]), .B(n6322), .Z(n16949) );
  XOR U16929 ( .A(n16939), .B(n16948), .Z(n16976) );
  XOR U16930 ( .A(n16977), .B(n16945), .Z(n16948) );
  XOR U16931 ( .A(p_input[1517]), .B(p_input[2061]), .Z(n16945) );
  XOR U16932 ( .A(p_input[1518]), .B(n6324), .Z(n16977) );
  XOR U16933 ( .A(p_input[1513]), .B(p_input[2057]), .Z(n16939) );
  XOR U16934 ( .A(n16957), .B(n16955), .Z(n16937) );
  XNOR U16935 ( .A(n16978), .B(n16962), .Z(n16955) );
  XOR U16936 ( .A(p_input[1512]), .B(p_input[2056]), .Z(n16962) );
  XOR U16937 ( .A(n16952), .B(n16961), .Z(n16978) );
  XOR U16938 ( .A(n16979), .B(n16958), .Z(n16961) );
  XOR U16939 ( .A(p_input[1510]), .B(p_input[2054]), .Z(n16958) );
  XOR U16940 ( .A(p_input[1511]), .B(n7007), .Z(n16979) );
  XOR U16941 ( .A(p_input[1506]), .B(p_input[2050]), .Z(n16952) );
  XNOR U16942 ( .A(n16967), .B(n16966), .Z(n16957) );
  XOR U16943 ( .A(n16980), .B(n16963), .Z(n16966) );
  XOR U16944 ( .A(p_input[1507]), .B(p_input[2051]), .Z(n16963) );
  XOR U16945 ( .A(p_input[1508]), .B(n7009), .Z(n16980) );
  XOR U16946 ( .A(p_input[1509]), .B(p_input[2053]), .Z(n16967) );
  XOR U16947 ( .A(n16981), .B(n16982), .Z(n16866) );
  AND U16948 ( .A(n383), .B(n16983), .Z(n16982) );
  XNOR U16949 ( .A(n16984), .B(n16981), .Z(n16983) );
  XNOR U16950 ( .A(n16985), .B(n16986), .Z(n383) );
  AND U16951 ( .A(n16987), .B(n16988), .Z(n16986) );
  XOR U16952 ( .A(n16879), .B(n16985), .Z(n16988) );
  AND U16953 ( .A(n16989), .B(n16990), .Z(n16879) );
  XNOR U16954 ( .A(n16876), .B(n16985), .Z(n16987) );
  XOR U16955 ( .A(n16991), .B(n16992), .Z(n16876) );
  AND U16956 ( .A(n387), .B(n16993), .Z(n16992) );
  XOR U16957 ( .A(n16994), .B(n16991), .Z(n16993) );
  XOR U16958 ( .A(n16995), .B(n16996), .Z(n16985) );
  AND U16959 ( .A(n16997), .B(n16998), .Z(n16996) );
  XNOR U16960 ( .A(n16995), .B(n16989), .Z(n16998) );
  IV U16961 ( .A(n16894), .Z(n16989) );
  XOR U16962 ( .A(n16999), .B(n17000), .Z(n16894) );
  XOR U16963 ( .A(n17001), .B(n16990), .Z(n17000) );
  AND U16964 ( .A(n16921), .B(n17002), .Z(n16990) );
  AND U16965 ( .A(n17003), .B(n17004), .Z(n17001) );
  XOR U16966 ( .A(n17005), .B(n16999), .Z(n17003) );
  XNOR U16967 ( .A(n16891), .B(n16995), .Z(n16997) );
  XOR U16968 ( .A(n17006), .B(n17007), .Z(n16891) );
  AND U16969 ( .A(n387), .B(n17008), .Z(n17007) );
  XOR U16970 ( .A(n17009), .B(n17006), .Z(n17008) );
  XOR U16971 ( .A(n17010), .B(n17011), .Z(n16995) );
  AND U16972 ( .A(n17012), .B(n17013), .Z(n17011) );
  XNOR U16973 ( .A(n17010), .B(n16921), .Z(n17013) );
  XOR U16974 ( .A(n17014), .B(n17004), .Z(n16921) );
  XNOR U16975 ( .A(n17015), .B(n16999), .Z(n17004) );
  XOR U16976 ( .A(n17016), .B(n17017), .Z(n16999) );
  AND U16977 ( .A(n17018), .B(n17019), .Z(n17017) );
  XOR U16978 ( .A(n17020), .B(n17016), .Z(n17018) );
  XNOR U16979 ( .A(n17021), .B(n17022), .Z(n17015) );
  AND U16980 ( .A(n17023), .B(n17024), .Z(n17022) );
  XOR U16981 ( .A(n17021), .B(n17025), .Z(n17023) );
  XNOR U16982 ( .A(n17005), .B(n17002), .Z(n17014) );
  AND U16983 ( .A(n17026), .B(n17027), .Z(n17002) );
  XOR U16984 ( .A(n17028), .B(n17029), .Z(n17005) );
  AND U16985 ( .A(n17030), .B(n17031), .Z(n17029) );
  XOR U16986 ( .A(n17028), .B(n17032), .Z(n17030) );
  XNOR U16987 ( .A(n16918), .B(n17010), .Z(n17012) );
  XOR U16988 ( .A(n17033), .B(n17034), .Z(n16918) );
  AND U16989 ( .A(n387), .B(n17035), .Z(n17034) );
  XNOR U16990 ( .A(n17036), .B(n17033), .Z(n17035) );
  XOR U16991 ( .A(n17037), .B(n17038), .Z(n17010) );
  AND U16992 ( .A(n17039), .B(n17040), .Z(n17038) );
  XNOR U16993 ( .A(n17037), .B(n17026), .Z(n17040) );
  IV U16994 ( .A(n16971), .Z(n17026) );
  XNOR U16995 ( .A(n17041), .B(n17019), .Z(n16971) );
  XNOR U16996 ( .A(n17042), .B(n17025), .Z(n17019) );
  XNOR U16997 ( .A(n17043), .B(n17044), .Z(n17025) );
  NOR U16998 ( .A(n17045), .B(n17046), .Z(n17044) );
  XOR U16999 ( .A(n17043), .B(n17047), .Z(n17045) );
  XNOR U17000 ( .A(n17024), .B(n17016), .Z(n17042) );
  XOR U17001 ( .A(n17048), .B(n17049), .Z(n17016) );
  AND U17002 ( .A(n17050), .B(n17051), .Z(n17049) );
  XOR U17003 ( .A(n17048), .B(n17052), .Z(n17050) );
  XNOR U17004 ( .A(n17053), .B(n17021), .Z(n17024) );
  XOR U17005 ( .A(n17054), .B(n17055), .Z(n17021) );
  AND U17006 ( .A(n17056), .B(n17057), .Z(n17055) );
  XNOR U17007 ( .A(n17058), .B(n17059), .Z(n17056) );
  IV U17008 ( .A(n17054), .Z(n17058) );
  XNOR U17009 ( .A(n17060), .B(n17061), .Z(n17053) );
  NOR U17010 ( .A(n17062), .B(n17063), .Z(n17061) );
  XNOR U17011 ( .A(n17060), .B(n17064), .Z(n17062) );
  XNOR U17012 ( .A(n17020), .B(n17027), .Z(n17041) );
  NOR U17013 ( .A(n16984), .B(n17065), .Z(n17027) );
  XOR U17014 ( .A(n17032), .B(n17031), .Z(n17020) );
  XNOR U17015 ( .A(n17066), .B(n17028), .Z(n17031) );
  XOR U17016 ( .A(n17067), .B(n17068), .Z(n17028) );
  AND U17017 ( .A(n17069), .B(n17070), .Z(n17068) );
  XNOR U17018 ( .A(n17071), .B(n17072), .Z(n17069) );
  IV U17019 ( .A(n17067), .Z(n17071) );
  XNOR U17020 ( .A(n17073), .B(n17074), .Z(n17066) );
  NOR U17021 ( .A(n17075), .B(n17076), .Z(n17074) );
  XNOR U17022 ( .A(n17073), .B(n17077), .Z(n17075) );
  XOR U17023 ( .A(n17078), .B(n17079), .Z(n17032) );
  NOR U17024 ( .A(n17080), .B(n17081), .Z(n17079) );
  XNOR U17025 ( .A(n17078), .B(n17082), .Z(n17080) );
  XNOR U17026 ( .A(n16968), .B(n17037), .Z(n17039) );
  XOR U17027 ( .A(n17083), .B(n17084), .Z(n16968) );
  AND U17028 ( .A(n387), .B(n17085), .Z(n17084) );
  XOR U17029 ( .A(n17086), .B(n17083), .Z(n17085) );
  AND U17030 ( .A(n16981), .B(n16984), .Z(n17037) );
  XOR U17031 ( .A(n17087), .B(n17065), .Z(n16984) );
  XNOR U17032 ( .A(p_input[1520]), .B(p_input[2048]), .Z(n17065) );
  XNOR U17033 ( .A(n17052), .B(n17051), .Z(n17087) );
  XNOR U17034 ( .A(n17088), .B(n17059), .Z(n17051) );
  XNOR U17035 ( .A(n17047), .B(n17046), .Z(n17059) );
  XNOR U17036 ( .A(n17089), .B(n17043), .Z(n17046) );
  XNOR U17037 ( .A(p_input[1530]), .B(p_input[2058]), .Z(n17043) );
  XOR U17038 ( .A(p_input[1531]), .B(n6319), .Z(n17089) );
  XOR U17039 ( .A(p_input[1532]), .B(p_input[2060]), .Z(n17047) );
  XOR U17040 ( .A(n17057), .B(n17090), .Z(n17088) );
  IV U17041 ( .A(n17048), .Z(n17090) );
  XOR U17042 ( .A(p_input[1521]), .B(p_input[2049]), .Z(n17048) );
  XNOR U17043 ( .A(n17091), .B(n17064), .Z(n17057) );
  XNOR U17044 ( .A(p_input[1535]), .B(n6322), .Z(n17064) );
  XOR U17045 ( .A(n17054), .B(n17063), .Z(n17091) );
  XOR U17046 ( .A(n17092), .B(n17060), .Z(n17063) );
  XOR U17047 ( .A(p_input[1533]), .B(p_input[2061]), .Z(n17060) );
  XOR U17048 ( .A(p_input[1534]), .B(n6324), .Z(n17092) );
  XOR U17049 ( .A(p_input[1529]), .B(p_input[2057]), .Z(n17054) );
  XOR U17050 ( .A(n17072), .B(n17070), .Z(n17052) );
  XNOR U17051 ( .A(n17093), .B(n17077), .Z(n17070) );
  XOR U17052 ( .A(p_input[1528]), .B(p_input[2056]), .Z(n17077) );
  XOR U17053 ( .A(n17067), .B(n17076), .Z(n17093) );
  XOR U17054 ( .A(n17094), .B(n17073), .Z(n17076) );
  XOR U17055 ( .A(p_input[1526]), .B(p_input[2054]), .Z(n17073) );
  XOR U17056 ( .A(p_input[1527]), .B(n7007), .Z(n17094) );
  XOR U17057 ( .A(p_input[1522]), .B(p_input[2050]), .Z(n17067) );
  XNOR U17058 ( .A(n17082), .B(n17081), .Z(n17072) );
  XOR U17059 ( .A(n17095), .B(n17078), .Z(n17081) );
  XOR U17060 ( .A(p_input[1523]), .B(p_input[2051]), .Z(n17078) );
  XOR U17061 ( .A(p_input[1524]), .B(n7009), .Z(n17095) );
  XOR U17062 ( .A(p_input[1525]), .B(p_input[2053]), .Z(n17082) );
  XOR U17063 ( .A(n17096), .B(n17097), .Z(n16981) );
  AND U17064 ( .A(n387), .B(n17098), .Z(n17097) );
  XNOR U17065 ( .A(n17099), .B(n17096), .Z(n17098) );
  XNOR U17066 ( .A(n17100), .B(n17101), .Z(n387) );
  AND U17067 ( .A(n17102), .B(n17103), .Z(n17101) );
  XOR U17068 ( .A(n16994), .B(n17100), .Z(n17103) );
  AND U17069 ( .A(n17104), .B(n17105), .Z(n16994) );
  XNOR U17070 ( .A(n16991), .B(n17100), .Z(n17102) );
  XOR U17071 ( .A(n17106), .B(n17107), .Z(n16991) );
  AND U17072 ( .A(n391), .B(n17108), .Z(n17107) );
  XOR U17073 ( .A(n17109), .B(n17106), .Z(n17108) );
  XOR U17074 ( .A(n17110), .B(n17111), .Z(n17100) );
  AND U17075 ( .A(n17112), .B(n17113), .Z(n17111) );
  XNOR U17076 ( .A(n17110), .B(n17104), .Z(n17113) );
  IV U17077 ( .A(n17009), .Z(n17104) );
  XOR U17078 ( .A(n17114), .B(n17115), .Z(n17009) );
  XOR U17079 ( .A(n17116), .B(n17105), .Z(n17115) );
  AND U17080 ( .A(n17036), .B(n17117), .Z(n17105) );
  AND U17081 ( .A(n17118), .B(n17119), .Z(n17116) );
  XOR U17082 ( .A(n17120), .B(n17114), .Z(n17118) );
  XNOR U17083 ( .A(n17006), .B(n17110), .Z(n17112) );
  XOR U17084 ( .A(n17121), .B(n17122), .Z(n17006) );
  AND U17085 ( .A(n391), .B(n17123), .Z(n17122) );
  XOR U17086 ( .A(n17124), .B(n17121), .Z(n17123) );
  XOR U17087 ( .A(n17125), .B(n17126), .Z(n17110) );
  AND U17088 ( .A(n17127), .B(n17128), .Z(n17126) );
  XNOR U17089 ( .A(n17125), .B(n17036), .Z(n17128) );
  XOR U17090 ( .A(n17129), .B(n17119), .Z(n17036) );
  XNOR U17091 ( .A(n17130), .B(n17114), .Z(n17119) );
  XOR U17092 ( .A(n17131), .B(n17132), .Z(n17114) );
  AND U17093 ( .A(n17133), .B(n17134), .Z(n17132) );
  XOR U17094 ( .A(n17135), .B(n17131), .Z(n17133) );
  XNOR U17095 ( .A(n17136), .B(n17137), .Z(n17130) );
  AND U17096 ( .A(n17138), .B(n17139), .Z(n17137) );
  XOR U17097 ( .A(n17136), .B(n17140), .Z(n17138) );
  XNOR U17098 ( .A(n17120), .B(n17117), .Z(n17129) );
  AND U17099 ( .A(n17141), .B(n17142), .Z(n17117) );
  XOR U17100 ( .A(n17143), .B(n17144), .Z(n17120) );
  AND U17101 ( .A(n17145), .B(n17146), .Z(n17144) );
  XOR U17102 ( .A(n17143), .B(n17147), .Z(n17145) );
  XNOR U17103 ( .A(n17033), .B(n17125), .Z(n17127) );
  XOR U17104 ( .A(n17148), .B(n17149), .Z(n17033) );
  AND U17105 ( .A(n391), .B(n17150), .Z(n17149) );
  XNOR U17106 ( .A(n17151), .B(n17148), .Z(n17150) );
  XOR U17107 ( .A(n17152), .B(n17153), .Z(n17125) );
  AND U17108 ( .A(n17154), .B(n17155), .Z(n17153) );
  XNOR U17109 ( .A(n17152), .B(n17141), .Z(n17155) );
  IV U17110 ( .A(n17086), .Z(n17141) );
  XNOR U17111 ( .A(n17156), .B(n17134), .Z(n17086) );
  XNOR U17112 ( .A(n17157), .B(n17140), .Z(n17134) );
  XNOR U17113 ( .A(n17158), .B(n17159), .Z(n17140) );
  NOR U17114 ( .A(n17160), .B(n17161), .Z(n17159) );
  XOR U17115 ( .A(n17158), .B(n17162), .Z(n17160) );
  XNOR U17116 ( .A(n17139), .B(n17131), .Z(n17157) );
  XOR U17117 ( .A(n17163), .B(n17164), .Z(n17131) );
  AND U17118 ( .A(n17165), .B(n17166), .Z(n17164) );
  XOR U17119 ( .A(n17163), .B(n17167), .Z(n17165) );
  XNOR U17120 ( .A(n17168), .B(n17136), .Z(n17139) );
  XOR U17121 ( .A(n17169), .B(n17170), .Z(n17136) );
  AND U17122 ( .A(n17171), .B(n17172), .Z(n17170) );
  XNOR U17123 ( .A(n17173), .B(n17174), .Z(n17171) );
  IV U17124 ( .A(n17169), .Z(n17173) );
  XNOR U17125 ( .A(n17175), .B(n17176), .Z(n17168) );
  NOR U17126 ( .A(n17177), .B(n17178), .Z(n17176) );
  XNOR U17127 ( .A(n17175), .B(n17179), .Z(n17177) );
  XNOR U17128 ( .A(n17135), .B(n17142), .Z(n17156) );
  NOR U17129 ( .A(n17099), .B(n17180), .Z(n17142) );
  XOR U17130 ( .A(n17147), .B(n17146), .Z(n17135) );
  XNOR U17131 ( .A(n17181), .B(n17143), .Z(n17146) );
  XOR U17132 ( .A(n17182), .B(n17183), .Z(n17143) );
  AND U17133 ( .A(n17184), .B(n17185), .Z(n17183) );
  XNOR U17134 ( .A(n17186), .B(n17187), .Z(n17184) );
  IV U17135 ( .A(n17182), .Z(n17186) );
  XNOR U17136 ( .A(n17188), .B(n17189), .Z(n17181) );
  NOR U17137 ( .A(n17190), .B(n17191), .Z(n17189) );
  XNOR U17138 ( .A(n17188), .B(n17192), .Z(n17190) );
  XOR U17139 ( .A(n17193), .B(n17194), .Z(n17147) );
  NOR U17140 ( .A(n17195), .B(n17196), .Z(n17194) );
  XNOR U17141 ( .A(n17193), .B(n17197), .Z(n17195) );
  XNOR U17142 ( .A(n17083), .B(n17152), .Z(n17154) );
  XOR U17143 ( .A(n17198), .B(n17199), .Z(n17083) );
  AND U17144 ( .A(n391), .B(n17200), .Z(n17199) );
  XOR U17145 ( .A(n17201), .B(n17198), .Z(n17200) );
  AND U17146 ( .A(n17096), .B(n17099), .Z(n17152) );
  XOR U17147 ( .A(n17202), .B(n17180), .Z(n17099) );
  XNOR U17148 ( .A(p_input[1536]), .B(p_input[2048]), .Z(n17180) );
  XNOR U17149 ( .A(n17167), .B(n17166), .Z(n17202) );
  XNOR U17150 ( .A(n17203), .B(n17174), .Z(n17166) );
  XNOR U17151 ( .A(n17162), .B(n17161), .Z(n17174) );
  XNOR U17152 ( .A(n17204), .B(n17158), .Z(n17161) );
  XNOR U17153 ( .A(p_input[1546]), .B(p_input[2058]), .Z(n17158) );
  XOR U17154 ( .A(p_input[1547]), .B(n6319), .Z(n17204) );
  XOR U17155 ( .A(p_input[1548]), .B(p_input[2060]), .Z(n17162) );
  XOR U17156 ( .A(n17172), .B(n17205), .Z(n17203) );
  IV U17157 ( .A(n17163), .Z(n17205) );
  XOR U17158 ( .A(p_input[1537]), .B(p_input[2049]), .Z(n17163) );
  XNOR U17159 ( .A(n17206), .B(n17179), .Z(n17172) );
  XNOR U17160 ( .A(p_input[1551]), .B(n6322), .Z(n17179) );
  XOR U17161 ( .A(n17169), .B(n17178), .Z(n17206) );
  XOR U17162 ( .A(n17207), .B(n17175), .Z(n17178) );
  XOR U17163 ( .A(p_input[1549]), .B(p_input[2061]), .Z(n17175) );
  XOR U17164 ( .A(p_input[1550]), .B(n6324), .Z(n17207) );
  XOR U17165 ( .A(p_input[1545]), .B(p_input[2057]), .Z(n17169) );
  XOR U17166 ( .A(n17187), .B(n17185), .Z(n17167) );
  XNOR U17167 ( .A(n17208), .B(n17192), .Z(n17185) );
  XOR U17168 ( .A(p_input[1544]), .B(p_input[2056]), .Z(n17192) );
  XOR U17169 ( .A(n17182), .B(n17191), .Z(n17208) );
  XOR U17170 ( .A(n17209), .B(n17188), .Z(n17191) );
  XOR U17171 ( .A(p_input[1542]), .B(p_input[2054]), .Z(n17188) );
  XOR U17172 ( .A(p_input[1543]), .B(n7007), .Z(n17209) );
  XOR U17173 ( .A(p_input[1538]), .B(p_input[2050]), .Z(n17182) );
  XNOR U17174 ( .A(n17197), .B(n17196), .Z(n17187) );
  XOR U17175 ( .A(n17210), .B(n17193), .Z(n17196) );
  XOR U17176 ( .A(p_input[1539]), .B(p_input[2051]), .Z(n17193) );
  XOR U17177 ( .A(p_input[1540]), .B(n7009), .Z(n17210) );
  XOR U17178 ( .A(p_input[1541]), .B(p_input[2053]), .Z(n17197) );
  XOR U17179 ( .A(n17211), .B(n17212), .Z(n17096) );
  AND U17180 ( .A(n391), .B(n17213), .Z(n17212) );
  XNOR U17181 ( .A(n17214), .B(n17211), .Z(n17213) );
  XNOR U17182 ( .A(n17215), .B(n17216), .Z(n391) );
  AND U17183 ( .A(n17217), .B(n17218), .Z(n17216) );
  XOR U17184 ( .A(n17109), .B(n17215), .Z(n17218) );
  AND U17185 ( .A(n17219), .B(n17220), .Z(n17109) );
  XNOR U17186 ( .A(n17106), .B(n17215), .Z(n17217) );
  XOR U17187 ( .A(n17221), .B(n17222), .Z(n17106) );
  AND U17188 ( .A(n395), .B(n17223), .Z(n17222) );
  XOR U17189 ( .A(n17224), .B(n17221), .Z(n17223) );
  XOR U17190 ( .A(n17225), .B(n17226), .Z(n17215) );
  AND U17191 ( .A(n17227), .B(n17228), .Z(n17226) );
  XNOR U17192 ( .A(n17225), .B(n17219), .Z(n17228) );
  IV U17193 ( .A(n17124), .Z(n17219) );
  XOR U17194 ( .A(n17229), .B(n17230), .Z(n17124) );
  XOR U17195 ( .A(n17231), .B(n17220), .Z(n17230) );
  AND U17196 ( .A(n17151), .B(n17232), .Z(n17220) );
  AND U17197 ( .A(n17233), .B(n17234), .Z(n17231) );
  XOR U17198 ( .A(n17235), .B(n17229), .Z(n17233) );
  XNOR U17199 ( .A(n17121), .B(n17225), .Z(n17227) );
  XOR U17200 ( .A(n17236), .B(n17237), .Z(n17121) );
  AND U17201 ( .A(n395), .B(n17238), .Z(n17237) );
  XOR U17202 ( .A(n17239), .B(n17236), .Z(n17238) );
  XOR U17203 ( .A(n17240), .B(n17241), .Z(n17225) );
  AND U17204 ( .A(n17242), .B(n17243), .Z(n17241) );
  XNOR U17205 ( .A(n17240), .B(n17151), .Z(n17243) );
  XOR U17206 ( .A(n17244), .B(n17234), .Z(n17151) );
  XNOR U17207 ( .A(n17245), .B(n17229), .Z(n17234) );
  XOR U17208 ( .A(n17246), .B(n17247), .Z(n17229) );
  AND U17209 ( .A(n17248), .B(n17249), .Z(n17247) );
  XOR U17210 ( .A(n17250), .B(n17246), .Z(n17248) );
  XNOR U17211 ( .A(n17251), .B(n17252), .Z(n17245) );
  AND U17212 ( .A(n17253), .B(n17254), .Z(n17252) );
  XOR U17213 ( .A(n17251), .B(n17255), .Z(n17253) );
  XNOR U17214 ( .A(n17235), .B(n17232), .Z(n17244) );
  AND U17215 ( .A(n17256), .B(n17257), .Z(n17232) );
  XOR U17216 ( .A(n17258), .B(n17259), .Z(n17235) );
  AND U17217 ( .A(n17260), .B(n17261), .Z(n17259) );
  XOR U17218 ( .A(n17258), .B(n17262), .Z(n17260) );
  XNOR U17219 ( .A(n17148), .B(n17240), .Z(n17242) );
  XOR U17220 ( .A(n17263), .B(n17264), .Z(n17148) );
  AND U17221 ( .A(n395), .B(n17265), .Z(n17264) );
  XNOR U17222 ( .A(n17266), .B(n17263), .Z(n17265) );
  XOR U17223 ( .A(n17267), .B(n17268), .Z(n17240) );
  AND U17224 ( .A(n17269), .B(n17270), .Z(n17268) );
  XNOR U17225 ( .A(n17267), .B(n17256), .Z(n17270) );
  IV U17226 ( .A(n17201), .Z(n17256) );
  XNOR U17227 ( .A(n17271), .B(n17249), .Z(n17201) );
  XNOR U17228 ( .A(n17272), .B(n17255), .Z(n17249) );
  XNOR U17229 ( .A(n17273), .B(n17274), .Z(n17255) );
  NOR U17230 ( .A(n17275), .B(n17276), .Z(n17274) );
  XOR U17231 ( .A(n17273), .B(n17277), .Z(n17275) );
  XNOR U17232 ( .A(n17254), .B(n17246), .Z(n17272) );
  XOR U17233 ( .A(n17278), .B(n17279), .Z(n17246) );
  AND U17234 ( .A(n17280), .B(n17281), .Z(n17279) );
  XOR U17235 ( .A(n17278), .B(n17282), .Z(n17280) );
  XNOR U17236 ( .A(n17283), .B(n17251), .Z(n17254) );
  XOR U17237 ( .A(n17284), .B(n17285), .Z(n17251) );
  AND U17238 ( .A(n17286), .B(n17287), .Z(n17285) );
  XNOR U17239 ( .A(n17288), .B(n17289), .Z(n17286) );
  IV U17240 ( .A(n17284), .Z(n17288) );
  XNOR U17241 ( .A(n17290), .B(n17291), .Z(n17283) );
  NOR U17242 ( .A(n17292), .B(n17293), .Z(n17291) );
  XNOR U17243 ( .A(n17290), .B(n17294), .Z(n17292) );
  XNOR U17244 ( .A(n17250), .B(n17257), .Z(n17271) );
  NOR U17245 ( .A(n17214), .B(n17295), .Z(n17257) );
  XOR U17246 ( .A(n17262), .B(n17261), .Z(n17250) );
  XNOR U17247 ( .A(n17296), .B(n17258), .Z(n17261) );
  XOR U17248 ( .A(n17297), .B(n17298), .Z(n17258) );
  AND U17249 ( .A(n17299), .B(n17300), .Z(n17298) );
  XNOR U17250 ( .A(n17301), .B(n17302), .Z(n17299) );
  IV U17251 ( .A(n17297), .Z(n17301) );
  XNOR U17252 ( .A(n17303), .B(n17304), .Z(n17296) );
  NOR U17253 ( .A(n17305), .B(n17306), .Z(n17304) );
  XNOR U17254 ( .A(n17303), .B(n17307), .Z(n17305) );
  XOR U17255 ( .A(n17308), .B(n17309), .Z(n17262) );
  NOR U17256 ( .A(n17310), .B(n17311), .Z(n17309) );
  XNOR U17257 ( .A(n17308), .B(n17312), .Z(n17310) );
  XNOR U17258 ( .A(n17198), .B(n17267), .Z(n17269) );
  XOR U17259 ( .A(n17313), .B(n17314), .Z(n17198) );
  AND U17260 ( .A(n395), .B(n17315), .Z(n17314) );
  XOR U17261 ( .A(n17316), .B(n17313), .Z(n17315) );
  AND U17262 ( .A(n17211), .B(n17214), .Z(n17267) );
  XOR U17263 ( .A(n17317), .B(n17295), .Z(n17214) );
  XNOR U17264 ( .A(p_input[1552]), .B(p_input[2048]), .Z(n17295) );
  XNOR U17265 ( .A(n17282), .B(n17281), .Z(n17317) );
  XNOR U17266 ( .A(n17318), .B(n17289), .Z(n17281) );
  XNOR U17267 ( .A(n17277), .B(n17276), .Z(n17289) );
  XNOR U17268 ( .A(n17319), .B(n17273), .Z(n17276) );
  XNOR U17269 ( .A(p_input[1562]), .B(p_input[2058]), .Z(n17273) );
  XOR U17270 ( .A(p_input[1563]), .B(n6319), .Z(n17319) );
  XOR U17271 ( .A(p_input[1564]), .B(p_input[2060]), .Z(n17277) );
  XOR U17272 ( .A(n17287), .B(n17320), .Z(n17318) );
  IV U17273 ( .A(n17278), .Z(n17320) );
  XOR U17274 ( .A(p_input[1553]), .B(p_input[2049]), .Z(n17278) );
  XNOR U17275 ( .A(n17321), .B(n17294), .Z(n17287) );
  XNOR U17276 ( .A(p_input[1567]), .B(n6322), .Z(n17294) );
  XOR U17277 ( .A(n17284), .B(n17293), .Z(n17321) );
  XOR U17278 ( .A(n17322), .B(n17290), .Z(n17293) );
  XOR U17279 ( .A(p_input[1565]), .B(p_input[2061]), .Z(n17290) );
  XOR U17280 ( .A(p_input[1566]), .B(n6324), .Z(n17322) );
  XOR U17281 ( .A(p_input[1561]), .B(p_input[2057]), .Z(n17284) );
  XOR U17282 ( .A(n17302), .B(n17300), .Z(n17282) );
  XNOR U17283 ( .A(n17323), .B(n17307), .Z(n17300) );
  XOR U17284 ( .A(p_input[1560]), .B(p_input[2056]), .Z(n17307) );
  XOR U17285 ( .A(n17297), .B(n17306), .Z(n17323) );
  XOR U17286 ( .A(n17324), .B(n17303), .Z(n17306) );
  XOR U17287 ( .A(p_input[1558]), .B(p_input[2054]), .Z(n17303) );
  XOR U17288 ( .A(p_input[1559]), .B(n7007), .Z(n17324) );
  XOR U17289 ( .A(p_input[1554]), .B(p_input[2050]), .Z(n17297) );
  XNOR U17290 ( .A(n17312), .B(n17311), .Z(n17302) );
  XOR U17291 ( .A(n17325), .B(n17308), .Z(n17311) );
  XOR U17292 ( .A(p_input[1555]), .B(p_input[2051]), .Z(n17308) );
  XOR U17293 ( .A(p_input[1556]), .B(n7009), .Z(n17325) );
  XOR U17294 ( .A(p_input[1557]), .B(p_input[2053]), .Z(n17312) );
  XOR U17295 ( .A(n17326), .B(n17327), .Z(n17211) );
  AND U17296 ( .A(n395), .B(n17328), .Z(n17327) );
  XNOR U17297 ( .A(n17329), .B(n17326), .Z(n17328) );
  XNOR U17298 ( .A(n17330), .B(n17331), .Z(n395) );
  AND U17299 ( .A(n17332), .B(n17333), .Z(n17331) );
  XOR U17300 ( .A(n17224), .B(n17330), .Z(n17333) );
  AND U17301 ( .A(n17334), .B(n17335), .Z(n17224) );
  XNOR U17302 ( .A(n17221), .B(n17330), .Z(n17332) );
  XOR U17303 ( .A(n17336), .B(n17337), .Z(n17221) );
  AND U17304 ( .A(n399), .B(n17338), .Z(n17337) );
  XOR U17305 ( .A(n17339), .B(n17336), .Z(n17338) );
  XOR U17306 ( .A(n17340), .B(n17341), .Z(n17330) );
  AND U17307 ( .A(n17342), .B(n17343), .Z(n17341) );
  XNOR U17308 ( .A(n17340), .B(n17334), .Z(n17343) );
  IV U17309 ( .A(n17239), .Z(n17334) );
  XOR U17310 ( .A(n17344), .B(n17345), .Z(n17239) );
  XOR U17311 ( .A(n17346), .B(n17335), .Z(n17345) );
  AND U17312 ( .A(n17266), .B(n17347), .Z(n17335) );
  AND U17313 ( .A(n17348), .B(n17349), .Z(n17346) );
  XOR U17314 ( .A(n17350), .B(n17344), .Z(n17348) );
  XNOR U17315 ( .A(n17236), .B(n17340), .Z(n17342) );
  XOR U17316 ( .A(n17351), .B(n17352), .Z(n17236) );
  AND U17317 ( .A(n399), .B(n17353), .Z(n17352) );
  XOR U17318 ( .A(n17354), .B(n17351), .Z(n17353) );
  XOR U17319 ( .A(n17355), .B(n17356), .Z(n17340) );
  AND U17320 ( .A(n17357), .B(n17358), .Z(n17356) );
  XNOR U17321 ( .A(n17355), .B(n17266), .Z(n17358) );
  XOR U17322 ( .A(n17359), .B(n17349), .Z(n17266) );
  XNOR U17323 ( .A(n17360), .B(n17344), .Z(n17349) );
  XOR U17324 ( .A(n17361), .B(n17362), .Z(n17344) );
  AND U17325 ( .A(n17363), .B(n17364), .Z(n17362) );
  XOR U17326 ( .A(n17365), .B(n17361), .Z(n17363) );
  XNOR U17327 ( .A(n17366), .B(n17367), .Z(n17360) );
  AND U17328 ( .A(n17368), .B(n17369), .Z(n17367) );
  XOR U17329 ( .A(n17366), .B(n17370), .Z(n17368) );
  XNOR U17330 ( .A(n17350), .B(n17347), .Z(n17359) );
  AND U17331 ( .A(n17371), .B(n17372), .Z(n17347) );
  XOR U17332 ( .A(n17373), .B(n17374), .Z(n17350) );
  AND U17333 ( .A(n17375), .B(n17376), .Z(n17374) );
  XOR U17334 ( .A(n17373), .B(n17377), .Z(n17375) );
  XNOR U17335 ( .A(n17263), .B(n17355), .Z(n17357) );
  XOR U17336 ( .A(n17378), .B(n17379), .Z(n17263) );
  AND U17337 ( .A(n399), .B(n17380), .Z(n17379) );
  XNOR U17338 ( .A(n17381), .B(n17378), .Z(n17380) );
  XOR U17339 ( .A(n17382), .B(n17383), .Z(n17355) );
  AND U17340 ( .A(n17384), .B(n17385), .Z(n17383) );
  XNOR U17341 ( .A(n17382), .B(n17371), .Z(n17385) );
  IV U17342 ( .A(n17316), .Z(n17371) );
  XNOR U17343 ( .A(n17386), .B(n17364), .Z(n17316) );
  XNOR U17344 ( .A(n17387), .B(n17370), .Z(n17364) );
  XNOR U17345 ( .A(n17388), .B(n17389), .Z(n17370) );
  NOR U17346 ( .A(n17390), .B(n17391), .Z(n17389) );
  XOR U17347 ( .A(n17388), .B(n17392), .Z(n17390) );
  XNOR U17348 ( .A(n17369), .B(n17361), .Z(n17387) );
  XOR U17349 ( .A(n17393), .B(n17394), .Z(n17361) );
  AND U17350 ( .A(n17395), .B(n17396), .Z(n17394) );
  XOR U17351 ( .A(n17393), .B(n17397), .Z(n17395) );
  XNOR U17352 ( .A(n17398), .B(n17366), .Z(n17369) );
  XOR U17353 ( .A(n17399), .B(n17400), .Z(n17366) );
  AND U17354 ( .A(n17401), .B(n17402), .Z(n17400) );
  XNOR U17355 ( .A(n17403), .B(n17404), .Z(n17401) );
  IV U17356 ( .A(n17399), .Z(n17403) );
  XNOR U17357 ( .A(n17405), .B(n17406), .Z(n17398) );
  NOR U17358 ( .A(n17407), .B(n17408), .Z(n17406) );
  XNOR U17359 ( .A(n17405), .B(n17409), .Z(n17407) );
  XNOR U17360 ( .A(n17365), .B(n17372), .Z(n17386) );
  NOR U17361 ( .A(n17329), .B(n17410), .Z(n17372) );
  XOR U17362 ( .A(n17377), .B(n17376), .Z(n17365) );
  XNOR U17363 ( .A(n17411), .B(n17373), .Z(n17376) );
  XOR U17364 ( .A(n17412), .B(n17413), .Z(n17373) );
  AND U17365 ( .A(n17414), .B(n17415), .Z(n17413) );
  XNOR U17366 ( .A(n17416), .B(n17417), .Z(n17414) );
  IV U17367 ( .A(n17412), .Z(n17416) );
  XNOR U17368 ( .A(n17418), .B(n17419), .Z(n17411) );
  NOR U17369 ( .A(n17420), .B(n17421), .Z(n17419) );
  XNOR U17370 ( .A(n17418), .B(n17422), .Z(n17420) );
  XOR U17371 ( .A(n17423), .B(n17424), .Z(n17377) );
  NOR U17372 ( .A(n17425), .B(n17426), .Z(n17424) );
  XNOR U17373 ( .A(n17423), .B(n17427), .Z(n17425) );
  XNOR U17374 ( .A(n17313), .B(n17382), .Z(n17384) );
  XOR U17375 ( .A(n17428), .B(n17429), .Z(n17313) );
  AND U17376 ( .A(n399), .B(n17430), .Z(n17429) );
  XOR U17377 ( .A(n17431), .B(n17428), .Z(n17430) );
  AND U17378 ( .A(n17326), .B(n17329), .Z(n17382) );
  XOR U17379 ( .A(n17432), .B(n17410), .Z(n17329) );
  XNOR U17380 ( .A(p_input[1568]), .B(p_input[2048]), .Z(n17410) );
  XNOR U17381 ( .A(n17397), .B(n17396), .Z(n17432) );
  XNOR U17382 ( .A(n17433), .B(n17404), .Z(n17396) );
  XNOR U17383 ( .A(n17392), .B(n17391), .Z(n17404) );
  XNOR U17384 ( .A(n17434), .B(n17388), .Z(n17391) );
  XNOR U17385 ( .A(p_input[1578]), .B(p_input[2058]), .Z(n17388) );
  XOR U17386 ( .A(p_input[1579]), .B(n6319), .Z(n17434) );
  XOR U17387 ( .A(p_input[1580]), .B(p_input[2060]), .Z(n17392) );
  XOR U17388 ( .A(n17402), .B(n17435), .Z(n17433) );
  IV U17389 ( .A(n17393), .Z(n17435) );
  XOR U17390 ( .A(p_input[1569]), .B(p_input[2049]), .Z(n17393) );
  XNOR U17391 ( .A(n17436), .B(n17409), .Z(n17402) );
  XNOR U17392 ( .A(p_input[1583]), .B(n6322), .Z(n17409) );
  XOR U17393 ( .A(n17399), .B(n17408), .Z(n17436) );
  XOR U17394 ( .A(n17437), .B(n17405), .Z(n17408) );
  XOR U17395 ( .A(p_input[1581]), .B(p_input[2061]), .Z(n17405) );
  XOR U17396 ( .A(p_input[1582]), .B(n6324), .Z(n17437) );
  XOR U17397 ( .A(p_input[1577]), .B(p_input[2057]), .Z(n17399) );
  XOR U17398 ( .A(n17417), .B(n17415), .Z(n17397) );
  XNOR U17399 ( .A(n17438), .B(n17422), .Z(n17415) );
  XOR U17400 ( .A(p_input[1576]), .B(p_input[2056]), .Z(n17422) );
  XOR U17401 ( .A(n17412), .B(n17421), .Z(n17438) );
  XOR U17402 ( .A(n17439), .B(n17418), .Z(n17421) );
  XOR U17403 ( .A(p_input[1574]), .B(p_input[2054]), .Z(n17418) );
  XOR U17404 ( .A(p_input[1575]), .B(n7007), .Z(n17439) );
  XOR U17405 ( .A(p_input[1570]), .B(p_input[2050]), .Z(n17412) );
  XNOR U17406 ( .A(n17427), .B(n17426), .Z(n17417) );
  XOR U17407 ( .A(n17440), .B(n17423), .Z(n17426) );
  XOR U17408 ( .A(p_input[1571]), .B(p_input[2051]), .Z(n17423) );
  XOR U17409 ( .A(p_input[1572]), .B(n7009), .Z(n17440) );
  XOR U17410 ( .A(p_input[1573]), .B(p_input[2053]), .Z(n17427) );
  XOR U17411 ( .A(n17441), .B(n17442), .Z(n17326) );
  AND U17412 ( .A(n399), .B(n17443), .Z(n17442) );
  XNOR U17413 ( .A(n17444), .B(n17441), .Z(n17443) );
  XNOR U17414 ( .A(n17445), .B(n17446), .Z(n399) );
  AND U17415 ( .A(n17447), .B(n17448), .Z(n17446) );
  XOR U17416 ( .A(n17339), .B(n17445), .Z(n17448) );
  AND U17417 ( .A(n17449), .B(n17450), .Z(n17339) );
  XNOR U17418 ( .A(n17336), .B(n17445), .Z(n17447) );
  XOR U17419 ( .A(n17451), .B(n17452), .Z(n17336) );
  AND U17420 ( .A(n403), .B(n17453), .Z(n17452) );
  XOR U17421 ( .A(n17454), .B(n17451), .Z(n17453) );
  XOR U17422 ( .A(n17455), .B(n17456), .Z(n17445) );
  AND U17423 ( .A(n17457), .B(n17458), .Z(n17456) );
  XNOR U17424 ( .A(n17455), .B(n17449), .Z(n17458) );
  IV U17425 ( .A(n17354), .Z(n17449) );
  XOR U17426 ( .A(n17459), .B(n17460), .Z(n17354) );
  XOR U17427 ( .A(n17461), .B(n17450), .Z(n17460) );
  AND U17428 ( .A(n17381), .B(n17462), .Z(n17450) );
  AND U17429 ( .A(n17463), .B(n17464), .Z(n17461) );
  XOR U17430 ( .A(n17465), .B(n17459), .Z(n17463) );
  XNOR U17431 ( .A(n17351), .B(n17455), .Z(n17457) );
  XOR U17432 ( .A(n17466), .B(n17467), .Z(n17351) );
  AND U17433 ( .A(n403), .B(n17468), .Z(n17467) );
  XOR U17434 ( .A(n17469), .B(n17466), .Z(n17468) );
  XOR U17435 ( .A(n17470), .B(n17471), .Z(n17455) );
  AND U17436 ( .A(n17472), .B(n17473), .Z(n17471) );
  XNOR U17437 ( .A(n17470), .B(n17381), .Z(n17473) );
  XOR U17438 ( .A(n17474), .B(n17464), .Z(n17381) );
  XNOR U17439 ( .A(n17475), .B(n17459), .Z(n17464) );
  XOR U17440 ( .A(n17476), .B(n17477), .Z(n17459) );
  AND U17441 ( .A(n17478), .B(n17479), .Z(n17477) );
  XOR U17442 ( .A(n17480), .B(n17476), .Z(n17478) );
  XNOR U17443 ( .A(n17481), .B(n17482), .Z(n17475) );
  AND U17444 ( .A(n17483), .B(n17484), .Z(n17482) );
  XOR U17445 ( .A(n17481), .B(n17485), .Z(n17483) );
  XNOR U17446 ( .A(n17465), .B(n17462), .Z(n17474) );
  AND U17447 ( .A(n17486), .B(n17487), .Z(n17462) );
  XOR U17448 ( .A(n17488), .B(n17489), .Z(n17465) );
  AND U17449 ( .A(n17490), .B(n17491), .Z(n17489) );
  XOR U17450 ( .A(n17488), .B(n17492), .Z(n17490) );
  XNOR U17451 ( .A(n17378), .B(n17470), .Z(n17472) );
  XOR U17452 ( .A(n17493), .B(n17494), .Z(n17378) );
  AND U17453 ( .A(n403), .B(n17495), .Z(n17494) );
  XNOR U17454 ( .A(n17496), .B(n17493), .Z(n17495) );
  XOR U17455 ( .A(n17497), .B(n17498), .Z(n17470) );
  AND U17456 ( .A(n17499), .B(n17500), .Z(n17498) );
  XNOR U17457 ( .A(n17497), .B(n17486), .Z(n17500) );
  IV U17458 ( .A(n17431), .Z(n17486) );
  XNOR U17459 ( .A(n17501), .B(n17479), .Z(n17431) );
  XNOR U17460 ( .A(n17502), .B(n17485), .Z(n17479) );
  XNOR U17461 ( .A(n17503), .B(n17504), .Z(n17485) );
  NOR U17462 ( .A(n17505), .B(n17506), .Z(n17504) );
  XOR U17463 ( .A(n17503), .B(n17507), .Z(n17505) );
  XNOR U17464 ( .A(n17484), .B(n17476), .Z(n17502) );
  XOR U17465 ( .A(n17508), .B(n17509), .Z(n17476) );
  AND U17466 ( .A(n17510), .B(n17511), .Z(n17509) );
  XOR U17467 ( .A(n17508), .B(n17512), .Z(n17510) );
  XNOR U17468 ( .A(n17513), .B(n17481), .Z(n17484) );
  XOR U17469 ( .A(n17514), .B(n17515), .Z(n17481) );
  AND U17470 ( .A(n17516), .B(n17517), .Z(n17515) );
  XNOR U17471 ( .A(n17518), .B(n17519), .Z(n17516) );
  IV U17472 ( .A(n17514), .Z(n17518) );
  XNOR U17473 ( .A(n17520), .B(n17521), .Z(n17513) );
  NOR U17474 ( .A(n17522), .B(n17523), .Z(n17521) );
  XNOR U17475 ( .A(n17520), .B(n17524), .Z(n17522) );
  XNOR U17476 ( .A(n17480), .B(n17487), .Z(n17501) );
  NOR U17477 ( .A(n17444), .B(n17525), .Z(n17487) );
  XOR U17478 ( .A(n17492), .B(n17491), .Z(n17480) );
  XNOR U17479 ( .A(n17526), .B(n17488), .Z(n17491) );
  XOR U17480 ( .A(n17527), .B(n17528), .Z(n17488) );
  AND U17481 ( .A(n17529), .B(n17530), .Z(n17528) );
  XNOR U17482 ( .A(n17531), .B(n17532), .Z(n17529) );
  IV U17483 ( .A(n17527), .Z(n17531) );
  XNOR U17484 ( .A(n17533), .B(n17534), .Z(n17526) );
  NOR U17485 ( .A(n17535), .B(n17536), .Z(n17534) );
  XNOR U17486 ( .A(n17533), .B(n17537), .Z(n17535) );
  XOR U17487 ( .A(n17538), .B(n17539), .Z(n17492) );
  NOR U17488 ( .A(n17540), .B(n17541), .Z(n17539) );
  XNOR U17489 ( .A(n17538), .B(n17542), .Z(n17540) );
  XNOR U17490 ( .A(n17428), .B(n17497), .Z(n17499) );
  XOR U17491 ( .A(n17543), .B(n17544), .Z(n17428) );
  AND U17492 ( .A(n403), .B(n17545), .Z(n17544) );
  XOR U17493 ( .A(n17546), .B(n17543), .Z(n17545) );
  AND U17494 ( .A(n17441), .B(n17444), .Z(n17497) );
  XOR U17495 ( .A(n17547), .B(n17525), .Z(n17444) );
  XNOR U17496 ( .A(p_input[1584]), .B(p_input[2048]), .Z(n17525) );
  XNOR U17497 ( .A(n17512), .B(n17511), .Z(n17547) );
  XNOR U17498 ( .A(n17548), .B(n17519), .Z(n17511) );
  XNOR U17499 ( .A(n17507), .B(n17506), .Z(n17519) );
  XNOR U17500 ( .A(n17549), .B(n17503), .Z(n17506) );
  XNOR U17501 ( .A(p_input[1594]), .B(p_input[2058]), .Z(n17503) );
  XOR U17502 ( .A(p_input[1595]), .B(n6319), .Z(n17549) );
  XOR U17503 ( .A(p_input[1596]), .B(p_input[2060]), .Z(n17507) );
  XOR U17504 ( .A(n17517), .B(n17550), .Z(n17548) );
  IV U17505 ( .A(n17508), .Z(n17550) );
  XOR U17506 ( .A(p_input[1585]), .B(p_input[2049]), .Z(n17508) );
  XNOR U17507 ( .A(n17551), .B(n17524), .Z(n17517) );
  XNOR U17508 ( .A(p_input[1599]), .B(n6322), .Z(n17524) );
  XOR U17509 ( .A(n17514), .B(n17523), .Z(n17551) );
  XOR U17510 ( .A(n17552), .B(n17520), .Z(n17523) );
  XOR U17511 ( .A(p_input[1597]), .B(p_input[2061]), .Z(n17520) );
  XOR U17512 ( .A(p_input[1598]), .B(n6324), .Z(n17552) );
  XOR U17513 ( .A(p_input[1593]), .B(p_input[2057]), .Z(n17514) );
  XOR U17514 ( .A(n17532), .B(n17530), .Z(n17512) );
  XNOR U17515 ( .A(n17553), .B(n17537), .Z(n17530) );
  XOR U17516 ( .A(p_input[1592]), .B(p_input[2056]), .Z(n17537) );
  XOR U17517 ( .A(n17527), .B(n17536), .Z(n17553) );
  XOR U17518 ( .A(n17554), .B(n17533), .Z(n17536) );
  XOR U17519 ( .A(p_input[1590]), .B(p_input[2054]), .Z(n17533) );
  XOR U17520 ( .A(p_input[1591]), .B(n7007), .Z(n17554) );
  XOR U17521 ( .A(p_input[1586]), .B(p_input[2050]), .Z(n17527) );
  XNOR U17522 ( .A(n17542), .B(n17541), .Z(n17532) );
  XOR U17523 ( .A(n17555), .B(n17538), .Z(n17541) );
  XOR U17524 ( .A(p_input[1587]), .B(p_input[2051]), .Z(n17538) );
  XOR U17525 ( .A(p_input[1588]), .B(n7009), .Z(n17555) );
  XOR U17526 ( .A(p_input[1589]), .B(p_input[2053]), .Z(n17542) );
  XOR U17527 ( .A(n17556), .B(n17557), .Z(n17441) );
  AND U17528 ( .A(n403), .B(n17558), .Z(n17557) );
  XNOR U17529 ( .A(n17559), .B(n17556), .Z(n17558) );
  XNOR U17530 ( .A(n17560), .B(n17561), .Z(n403) );
  AND U17531 ( .A(n17562), .B(n17563), .Z(n17561) );
  XOR U17532 ( .A(n17454), .B(n17560), .Z(n17563) );
  AND U17533 ( .A(n17564), .B(n17565), .Z(n17454) );
  XNOR U17534 ( .A(n17451), .B(n17560), .Z(n17562) );
  XOR U17535 ( .A(n17566), .B(n17567), .Z(n17451) );
  AND U17536 ( .A(n407), .B(n17568), .Z(n17567) );
  XOR U17537 ( .A(n17569), .B(n17566), .Z(n17568) );
  XOR U17538 ( .A(n17570), .B(n17571), .Z(n17560) );
  AND U17539 ( .A(n17572), .B(n17573), .Z(n17571) );
  XNOR U17540 ( .A(n17570), .B(n17564), .Z(n17573) );
  IV U17541 ( .A(n17469), .Z(n17564) );
  XOR U17542 ( .A(n17574), .B(n17575), .Z(n17469) );
  XOR U17543 ( .A(n17576), .B(n17565), .Z(n17575) );
  AND U17544 ( .A(n17496), .B(n17577), .Z(n17565) );
  AND U17545 ( .A(n17578), .B(n17579), .Z(n17576) );
  XOR U17546 ( .A(n17580), .B(n17574), .Z(n17578) );
  XNOR U17547 ( .A(n17466), .B(n17570), .Z(n17572) );
  XOR U17548 ( .A(n17581), .B(n17582), .Z(n17466) );
  AND U17549 ( .A(n407), .B(n17583), .Z(n17582) );
  XOR U17550 ( .A(n17584), .B(n17581), .Z(n17583) );
  XOR U17551 ( .A(n17585), .B(n17586), .Z(n17570) );
  AND U17552 ( .A(n17587), .B(n17588), .Z(n17586) );
  XNOR U17553 ( .A(n17585), .B(n17496), .Z(n17588) );
  XOR U17554 ( .A(n17589), .B(n17579), .Z(n17496) );
  XNOR U17555 ( .A(n17590), .B(n17574), .Z(n17579) );
  XOR U17556 ( .A(n17591), .B(n17592), .Z(n17574) );
  AND U17557 ( .A(n17593), .B(n17594), .Z(n17592) );
  XOR U17558 ( .A(n17595), .B(n17591), .Z(n17593) );
  XNOR U17559 ( .A(n17596), .B(n17597), .Z(n17590) );
  AND U17560 ( .A(n17598), .B(n17599), .Z(n17597) );
  XOR U17561 ( .A(n17596), .B(n17600), .Z(n17598) );
  XNOR U17562 ( .A(n17580), .B(n17577), .Z(n17589) );
  AND U17563 ( .A(n17601), .B(n17602), .Z(n17577) );
  XOR U17564 ( .A(n17603), .B(n17604), .Z(n17580) );
  AND U17565 ( .A(n17605), .B(n17606), .Z(n17604) );
  XOR U17566 ( .A(n17603), .B(n17607), .Z(n17605) );
  XNOR U17567 ( .A(n17493), .B(n17585), .Z(n17587) );
  XOR U17568 ( .A(n17608), .B(n17609), .Z(n17493) );
  AND U17569 ( .A(n407), .B(n17610), .Z(n17609) );
  XNOR U17570 ( .A(n17611), .B(n17608), .Z(n17610) );
  XOR U17571 ( .A(n17612), .B(n17613), .Z(n17585) );
  AND U17572 ( .A(n17614), .B(n17615), .Z(n17613) );
  XNOR U17573 ( .A(n17612), .B(n17601), .Z(n17615) );
  IV U17574 ( .A(n17546), .Z(n17601) );
  XNOR U17575 ( .A(n17616), .B(n17594), .Z(n17546) );
  XNOR U17576 ( .A(n17617), .B(n17600), .Z(n17594) );
  XNOR U17577 ( .A(n17618), .B(n17619), .Z(n17600) );
  NOR U17578 ( .A(n17620), .B(n17621), .Z(n17619) );
  XOR U17579 ( .A(n17618), .B(n17622), .Z(n17620) );
  XNOR U17580 ( .A(n17599), .B(n17591), .Z(n17617) );
  XOR U17581 ( .A(n17623), .B(n17624), .Z(n17591) );
  AND U17582 ( .A(n17625), .B(n17626), .Z(n17624) );
  XOR U17583 ( .A(n17623), .B(n17627), .Z(n17625) );
  XNOR U17584 ( .A(n17628), .B(n17596), .Z(n17599) );
  XOR U17585 ( .A(n17629), .B(n17630), .Z(n17596) );
  AND U17586 ( .A(n17631), .B(n17632), .Z(n17630) );
  XNOR U17587 ( .A(n17633), .B(n17634), .Z(n17631) );
  IV U17588 ( .A(n17629), .Z(n17633) );
  XNOR U17589 ( .A(n17635), .B(n17636), .Z(n17628) );
  NOR U17590 ( .A(n17637), .B(n17638), .Z(n17636) );
  XNOR U17591 ( .A(n17635), .B(n17639), .Z(n17637) );
  XNOR U17592 ( .A(n17595), .B(n17602), .Z(n17616) );
  NOR U17593 ( .A(n17559), .B(n17640), .Z(n17602) );
  XOR U17594 ( .A(n17607), .B(n17606), .Z(n17595) );
  XNOR U17595 ( .A(n17641), .B(n17603), .Z(n17606) );
  XOR U17596 ( .A(n17642), .B(n17643), .Z(n17603) );
  AND U17597 ( .A(n17644), .B(n17645), .Z(n17643) );
  XNOR U17598 ( .A(n17646), .B(n17647), .Z(n17644) );
  IV U17599 ( .A(n17642), .Z(n17646) );
  XNOR U17600 ( .A(n17648), .B(n17649), .Z(n17641) );
  NOR U17601 ( .A(n17650), .B(n17651), .Z(n17649) );
  XNOR U17602 ( .A(n17648), .B(n17652), .Z(n17650) );
  XOR U17603 ( .A(n17653), .B(n17654), .Z(n17607) );
  NOR U17604 ( .A(n17655), .B(n17656), .Z(n17654) );
  XNOR U17605 ( .A(n17653), .B(n17657), .Z(n17655) );
  XNOR U17606 ( .A(n17543), .B(n17612), .Z(n17614) );
  XOR U17607 ( .A(n17658), .B(n17659), .Z(n17543) );
  AND U17608 ( .A(n407), .B(n17660), .Z(n17659) );
  XOR U17609 ( .A(n17661), .B(n17658), .Z(n17660) );
  AND U17610 ( .A(n17556), .B(n17559), .Z(n17612) );
  XOR U17611 ( .A(n17662), .B(n17640), .Z(n17559) );
  XNOR U17612 ( .A(p_input[1600]), .B(p_input[2048]), .Z(n17640) );
  XNOR U17613 ( .A(n17627), .B(n17626), .Z(n17662) );
  XNOR U17614 ( .A(n17663), .B(n17634), .Z(n17626) );
  XNOR U17615 ( .A(n17622), .B(n17621), .Z(n17634) );
  XNOR U17616 ( .A(n17664), .B(n17618), .Z(n17621) );
  XNOR U17617 ( .A(p_input[1610]), .B(p_input[2058]), .Z(n17618) );
  XOR U17618 ( .A(p_input[1611]), .B(n6319), .Z(n17664) );
  XOR U17619 ( .A(p_input[1612]), .B(p_input[2060]), .Z(n17622) );
  XOR U17620 ( .A(n17632), .B(n17665), .Z(n17663) );
  IV U17621 ( .A(n17623), .Z(n17665) );
  XOR U17622 ( .A(p_input[1601]), .B(p_input[2049]), .Z(n17623) );
  XNOR U17623 ( .A(n17666), .B(n17639), .Z(n17632) );
  XNOR U17624 ( .A(p_input[1615]), .B(n6322), .Z(n17639) );
  XOR U17625 ( .A(n17629), .B(n17638), .Z(n17666) );
  XOR U17626 ( .A(n17667), .B(n17635), .Z(n17638) );
  XOR U17627 ( .A(p_input[1613]), .B(p_input[2061]), .Z(n17635) );
  XOR U17628 ( .A(p_input[1614]), .B(n6324), .Z(n17667) );
  XOR U17629 ( .A(p_input[1609]), .B(p_input[2057]), .Z(n17629) );
  XOR U17630 ( .A(n17647), .B(n17645), .Z(n17627) );
  XNOR U17631 ( .A(n17668), .B(n17652), .Z(n17645) );
  XOR U17632 ( .A(p_input[1608]), .B(p_input[2056]), .Z(n17652) );
  XOR U17633 ( .A(n17642), .B(n17651), .Z(n17668) );
  XOR U17634 ( .A(n17669), .B(n17648), .Z(n17651) );
  XOR U17635 ( .A(p_input[1606]), .B(p_input[2054]), .Z(n17648) );
  XOR U17636 ( .A(p_input[1607]), .B(n7007), .Z(n17669) );
  XOR U17637 ( .A(p_input[1602]), .B(p_input[2050]), .Z(n17642) );
  XNOR U17638 ( .A(n17657), .B(n17656), .Z(n17647) );
  XOR U17639 ( .A(n17670), .B(n17653), .Z(n17656) );
  XOR U17640 ( .A(p_input[1603]), .B(p_input[2051]), .Z(n17653) );
  XOR U17641 ( .A(p_input[1604]), .B(n7009), .Z(n17670) );
  XOR U17642 ( .A(p_input[1605]), .B(p_input[2053]), .Z(n17657) );
  XOR U17643 ( .A(n17671), .B(n17672), .Z(n17556) );
  AND U17644 ( .A(n407), .B(n17673), .Z(n17672) );
  XNOR U17645 ( .A(n17674), .B(n17671), .Z(n17673) );
  XNOR U17646 ( .A(n17675), .B(n17676), .Z(n407) );
  AND U17647 ( .A(n17677), .B(n17678), .Z(n17676) );
  XOR U17648 ( .A(n17569), .B(n17675), .Z(n17678) );
  AND U17649 ( .A(n17679), .B(n17680), .Z(n17569) );
  XNOR U17650 ( .A(n17566), .B(n17675), .Z(n17677) );
  XOR U17651 ( .A(n17681), .B(n17682), .Z(n17566) );
  AND U17652 ( .A(n411), .B(n17683), .Z(n17682) );
  XOR U17653 ( .A(n17684), .B(n17681), .Z(n17683) );
  XOR U17654 ( .A(n17685), .B(n17686), .Z(n17675) );
  AND U17655 ( .A(n17687), .B(n17688), .Z(n17686) );
  XNOR U17656 ( .A(n17685), .B(n17679), .Z(n17688) );
  IV U17657 ( .A(n17584), .Z(n17679) );
  XOR U17658 ( .A(n17689), .B(n17690), .Z(n17584) );
  XOR U17659 ( .A(n17691), .B(n17680), .Z(n17690) );
  AND U17660 ( .A(n17611), .B(n17692), .Z(n17680) );
  AND U17661 ( .A(n17693), .B(n17694), .Z(n17691) );
  XOR U17662 ( .A(n17695), .B(n17689), .Z(n17693) );
  XNOR U17663 ( .A(n17581), .B(n17685), .Z(n17687) );
  XOR U17664 ( .A(n17696), .B(n17697), .Z(n17581) );
  AND U17665 ( .A(n411), .B(n17698), .Z(n17697) );
  XOR U17666 ( .A(n17699), .B(n17696), .Z(n17698) );
  XOR U17667 ( .A(n17700), .B(n17701), .Z(n17685) );
  AND U17668 ( .A(n17702), .B(n17703), .Z(n17701) );
  XNOR U17669 ( .A(n17700), .B(n17611), .Z(n17703) );
  XOR U17670 ( .A(n17704), .B(n17694), .Z(n17611) );
  XNOR U17671 ( .A(n17705), .B(n17689), .Z(n17694) );
  XOR U17672 ( .A(n17706), .B(n17707), .Z(n17689) );
  AND U17673 ( .A(n17708), .B(n17709), .Z(n17707) );
  XOR U17674 ( .A(n17710), .B(n17706), .Z(n17708) );
  XNOR U17675 ( .A(n17711), .B(n17712), .Z(n17705) );
  AND U17676 ( .A(n17713), .B(n17714), .Z(n17712) );
  XOR U17677 ( .A(n17711), .B(n17715), .Z(n17713) );
  XNOR U17678 ( .A(n17695), .B(n17692), .Z(n17704) );
  AND U17679 ( .A(n17716), .B(n17717), .Z(n17692) );
  XOR U17680 ( .A(n17718), .B(n17719), .Z(n17695) );
  AND U17681 ( .A(n17720), .B(n17721), .Z(n17719) );
  XOR U17682 ( .A(n17718), .B(n17722), .Z(n17720) );
  XNOR U17683 ( .A(n17608), .B(n17700), .Z(n17702) );
  XOR U17684 ( .A(n17723), .B(n17724), .Z(n17608) );
  AND U17685 ( .A(n411), .B(n17725), .Z(n17724) );
  XNOR U17686 ( .A(n17726), .B(n17723), .Z(n17725) );
  XOR U17687 ( .A(n17727), .B(n17728), .Z(n17700) );
  AND U17688 ( .A(n17729), .B(n17730), .Z(n17728) );
  XNOR U17689 ( .A(n17727), .B(n17716), .Z(n17730) );
  IV U17690 ( .A(n17661), .Z(n17716) );
  XNOR U17691 ( .A(n17731), .B(n17709), .Z(n17661) );
  XNOR U17692 ( .A(n17732), .B(n17715), .Z(n17709) );
  XNOR U17693 ( .A(n17733), .B(n17734), .Z(n17715) );
  NOR U17694 ( .A(n17735), .B(n17736), .Z(n17734) );
  XOR U17695 ( .A(n17733), .B(n17737), .Z(n17735) );
  XNOR U17696 ( .A(n17714), .B(n17706), .Z(n17732) );
  XOR U17697 ( .A(n17738), .B(n17739), .Z(n17706) );
  AND U17698 ( .A(n17740), .B(n17741), .Z(n17739) );
  XOR U17699 ( .A(n17738), .B(n17742), .Z(n17740) );
  XNOR U17700 ( .A(n17743), .B(n17711), .Z(n17714) );
  XOR U17701 ( .A(n17744), .B(n17745), .Z(n17711) );
  AND U17702 ( .A(n17746), .B(n17747), .Z(n17745) );
  XNOR U17703 ( .A(n17748), .B(n17749), .Z(n17746) );
  IV U17704 ( .A(n17744), .Z(n17748) );
  XNOR U17705 ( .A(n17750), .B(n17751), .Z(n17743) );
  NOR U17706 ( .A(n17752), .B(n17753), .Z(n17751) );
  XNOR U17707 ( .A(n17750), .B(n17754), .Z(n17752) );
  XNOR U17708 ( .A(n17710), .B(n17717), .Z(n17731) );
  NOR U17709 ( .A(n17674), .B(n17755), .Z(n17717) );
  XOR U17710 ( .A(n17722), .B(n17721), .Z(n17710) );
  XNOR U17711 ( .A(n17756), .B(n17718), .Z(n17721) );
  XOR U17712 ( .A(n17757), .B(n17758), .Z(n17718) );
  AND U17713 ( .A(n17759), .B(n17760), .Z(n17758) );
  XNOR U17714 ( .A(n17761), .B(n17762), .Z(n17759) );
  IV U17715 ( .A(n17757), .Z(n17761) );
  XNOR U17716 ( .A(n17763), .B(n17764), .Z(n17756) );
  NOR U17717 ( .A(n17765), .B(n17766), .Z(n17764) );
  XNOR U17718 ( .A(n17763), .B(n17767), .Z(n17765) );
  XOR U17719 ( .A(n17768), .B(n17769), .Z(n17722) );
  NOR U17720 ( .A(n17770), .B(n17771), .Z(n17769) );
  XNOR U17721 ( .A(n17768), .B(n17772), .Z(n17770) );
  XNOR U17722 ( .A(n17658), .B(n17727), .Z(n17729) );
  XOR U17723 ( .A(n17773), .B(n17774), .Z(n17658) );
  AND U17724 ( .A(n411), .B(n17775), .Z(n17774) );
  XOR U17725 ( .A(n17776), .B(n17773), .Z(n17775) );
  AND U17726 ( .A(n17671), .B(n17674), .Z(n17727) );
  XOR U17727 ( .A(n17777), .B(n17755), .Z(n17674) );
  XNOR U17728 ( .A(p_input[1616]), .B(p_input[2048]), .Z(n17755) );
  XNOR U17729 ( .A(n17742), .B(n17741), .Z(n17777) );
  XNOR U17730 ( .A(n17778), .B(n17749), .Z(n17741) );
  XNOR U17731 ( .A(n17737), .B(n17736), .Z(n17749) );
  XNOR U17732 ( .A(n17779), .B(n17733), .Z(n17736) );
  XNOR U17733 ( .A(p_input[1626]), .B(p_input[2058]), .Z(n17733) );
  XOR U17734 ( .A(p_input[1627]), .B(n6319), .Z(n17779) );
  XOR U17735 ( .A(p_input[1628]), .B(p_input[2060]), .Z(n17737) );
  XOR U17736 ( .A(n17747), .B(n17780), .Z(n17778) );
  IV U17737 ( .A(n17738), .Z(n17780) );
  XOR U17738 ( .A(p_input[1617]), .B(p_input[2049]), .Z(n17738) );
  XNOR U17739 ( .A(n17781), .B(n17754), .Z(n17747) );
  XNOR U17740 ( .A(p_input[1631]), .B(n6322), .Z(n17754) );
  XOR U17741 ( .A(n17744), .B(n17753), .Z(n17781) );
  XOR U17742 ( .A(n17782), .B(n17750), .Z(n17753) );
  XOR U17743 ( .A(p_input[1629]), .B(p_input[2061]), .Z(n17750) );
  XOR U17744 ( .A(p_input[1630]), .B(n6324), .Z(n17782) );
  XOR U17745 ( .A(p_input[1625]), .B(p_input[2057]), .Z(n17744) );
  XOR U17746 ( .A(n17762), .B(n17760), .Z(n17742) );
  XNOR U17747 ( .A(n17783), .B(n17767), .Z(n17760) );
  XOR U17748 ( .A(p_input[1624]), .B(p_input[2056]), .Z(n17767) );
  XOR U17749 ( .A(n17757), .B(n17766), .Z(n17783) );
  XOR U17750 ( .A(n17784), .B(n17763), .Z(n17766) );
  XOR U17751 ( .A(p_input[1622]), .B(p_input[2054]), .Z(n17763) );
  XOR U17752 ( .A(p_input[1623]), .B(n7007), .Z(n17784) );
  XOR U17753 ( .A(p_input[1618]), .B(p_input[2050]), .Z(n17757) );
  XNOR U17754 ( .A(n17772), .B(n17771), .Z(n17762) );
  XOR U17755 ( .A(n17785), .B(n17768), .Z(n17771) );
  XOR U17756 ( .A(p_input[1619]), .B(p_input[2051]), .Z(n17768) );
  XOR U17757 ( .A(p_input[1620]), .B(n7009), .Z(n17785) );
  XOR U17758 ( .A(p_input[1621]), .B(p_input[2053]), .Z(n17772) );
  XOR U17759 ( .A(n17786), .B(n17787), .Z(n17671) );
  AND U17760 ( .A(n411), .B(n17788), .Z(n17787) );
  XNOR U17761 ( .A(n17789), .B(n17786), .Z(n17788) );
  XNOR U17762 ( .A(n17790), .B(n17791), .Z(n411) );
  AND U17763 ( .A(n17792), .B(n17793), .Z(n17791) );
  XOR U17764 ( .A(n17684), .B(n17790), .Z(n17793) );
  AND U17765 ( .A(n17794), .B(n17795), .Z(n17684) );
  XNOR U17766 ( .A(n17681), .B(n17790), .Z(n17792) );
  XOR U17767 ( .A(n17796), .B(n17797), .Z(n17681) );
  AND U17768 ( .A(n415), .B(n17798), .Z(n17797) );
  XOR U17769 ( .A(n17799), .B(n17796), .Z(n17798) );
  XOR U17770 ( .A(n17800), .B(n17801), .Z(n17790) );
  AND U17771 ( .A(n17802), .B(n17803), .Z(n17801) );
  XNOR U17772 ( .A(n17800), .B(n17794), .Z(n17803) );
  IV U17773 ( .A(n17699), .Z(n17794) );
  XOR U17774 ( .A(n17804), .B(n17805), .Z(n17699) );
  XOR U17775 ( .A(n17806), .B(n17795), .Z(n17805) );
  AND U17776 ( .A(n17726), .B(n17807), .Z(n17795) );
  AND U17777 ( .A(n17808), .B(n17809), .Z(n17806) );
  XOR U17778 ( .A(n17810), .B(n17804), .Z(n17808) );
  XNOR U17779 ( .A(n17696), .B(n17800), .Z(n17802) );
  XOR U17780 ( .A(n17811), .B(n17812), .Z(n17696) );
  AND U17781 ( .A(n415), .B(n17813), .Z(n17812) );
  XOR U17782 ( .A(n17814), .B(n17811), .Z(n17813) );
  XOR U17783 ( .A(n17815), .B(n17816), .Z(n17800) );
  AND U17784 ( .A(n17817), .B(n17818), .Z(n17816) );
  XNOR U17785 ( .A(n17815), .B(n17726), .Z(n17818) );
  XOR U17786 ( .A(n17819), .B(n17809), .Z(n17726) );
  XNOR U17787 ( .A(n17820), .B(n17804), .Z(n17809) );
  XOR U17788 ( .A(n17821), .B(n17822), .Z(n17804) );
  AND U17789 ( .A(n17823), .B(n17824), .Z(n17822) );
  XOR U17790 ( .A(n17825), .B(n17821), .Z(n17823) );
  XNOR U17791 ( .A(n17826), .B(n17827), .Z(n17820) );
  AND U17792 ( .A(n17828), .B(n17829), .Z(n17827) );
  XOR U17793 ( .A(n17826), .B(n17830), .Z(n17828) );
  XNOR U17794 ( .A(n17810), .B(n17807), .Z(n17819) );
  AND U17795 ( .A(n17831), .B(n17832), .Z(n17807) );
  XOR U17796 ( .A(n17833), .B(n17834), .Z(n17810) );
  AND U17797 ( .A(n17835), .B(n17836), .Z(n17834) );
  XOR U17798 ( .A(n17833), .B(n17837), .Z(n17835) );
  XNOR U17799 ( .A(n17723), .B(n17815), .Z(n17817) );
  XOR U17800 ( .A(n17838), .B(n17839), .Z(n17723) );
  AND U17801 ( .A(n415), .B(n17840), .Z(n17839) );
  XNOR U17802 ( .A(n17841), .B(n17838), .Z(n17840) );
  XOR U17803 ( .A(n17842), .B(n17843), .Z(n17815) );
  AND U17804 ( .A(n17844), .B(n17845), .Z(n17843) );
  XNOR U17805 ( .A(n17842), .B(n17831), .Z(n17845) );
  IV U17806 ( .A(n17776), .Z(n17831) );
  XNOR U17807 ( .A(n17846), .B(n17824), .Z(n17776) );
  XNOR U17808 ( .A(n17847), .B(n17830), .Z(n17824) );
  XNOR U17809 ( .A(n17848), .B(n17849), .Z(n17830) );
  NOR U17810 ( .A(n17850), .B(n17851), .Z(n17849) );
  XOR U17811 ( .A(n17848), .B(n17852), .Z(n17850) );
  XNOR U17812 ( .A(n17829), .B(n17821), .Z(n17847) );
  XOR U17813 ( .A(n17853), .B(n17854), .Z(n17821) );
  AND U17814 ( .A(n17855), .B(n17856), .Z(n17854) );
  XOR U17815 ( .A(n17853), .B(n17857), .Z(n17855) );
  XNOR U17816 ( .A(n17858), .B(n17826), .Z(n17829) );
  XOR U17817 ( .A(n17859), .B(n17860), .Z(n17826) );
  AND U17818 ( .A(n17861), .B(n17862), .Z(n17860) );
  XNOR U17819 ( .A(n17863), .B(n17864), .Z(n17861) );
  IV U17820 ( .A(n17859), .Z(n17863) );
  XNOR U17821 ( .A(n17865), .B(n17866), .Z(n17858) );
  NOR U17822 ( .A(n17867), .B(n17868), .Z(n17866) );
  XNOR U17823 ( .A(n17865), .B(n17869), .Z(n17867) );
  XNOR U17824 ( .A(n17825), .B(n17832), .Z(n17846) );
  NOR U17825 ( .A(n17789), .B(n17870), .Z(n17832) );
  XOR U17826 ( .A(n17837), .B(n17836), .Z(n17825) );
  XNOR U17827 ( .A(n17871), .B(n17833), .Z(n17836) );
  XOR U17828 ( .A(n17872), .B(n17873), .Z(n17833) );
  AND U17829 ( .A(n17874), .B(n17875), .Z(n17873) );
  XNOR U17830 ( .A(n17876), .B(n17877), .Z(n17874) );
  IV U17831 ( .A(n17872), .Z(n17876) );
  XNOR U17832 ( .A(n17878), .B(n17879), .Z(n17871) );
  NOR U17833 ( .A(n17880), .B(n17881), .Z(n17879) );
  XNOR U17834 ( .A(n17878), .B(n17882), .Z(n17880) );
  XOR U17835 ( .A(n17883), .B(n17884), .Z(n17837) );
  NOR U17836 ( .A(n17885), .B(n17886), .Z(n17884) );
  XNOR U17837 ( .A(n17883), .B(n17887), .Z(n17885) );
  XNOR U17838 ( .A(n17773), .B(n17842), .Z(n17844) );
  XOR U17839 ( .A(n17888), .B(n17889), .Z(n17773) );
  AND U17840 ( .A(n415), .B(n17890), .Z(n17889) );
  XOR U17841 ( .A(n17891), .B(n17888), .Z(n17890) );
  AND U17842 ( .A(n17786), .B(n17789), .Z(n17842) );
  XOR U17843 ( .A(n17892), .B(n17870), .Z(n17789) );
  XNOR U17844 ( .A(p_input[1632]), .B(p_input[2048]), .Z(n17870) );
  XNOR U17845 ( .A(n17857), .B(n17856), .Z(n17892) );
  XNOR U17846 ( .A(n17893), .B(n17864), .Z(n17856) );
  XNOR U17847 ( .A(n17852), .B(n17851), .Z(n17864) );
  XNOR U17848 ( .A(n17894), .B(n17848), .Z(n17851) );
  XNOR U17849 ( .A(p_input[1642]), .B(p_input[2058]), .Z(n17848) );
  XOR U17850 ( .A(p_input[1643]), .B(n6319), .Z(n17894) );
  XOR U17851 ( .A(p_input[1644]), .B(p_input[2060]), .Z(n17852) );
  XOR U17852 ( .A(n17862), .B(n17895), .Z(n17893) );
  IV U17853 ( .A(n17853), .Z(n17895) );
  XOR U17854 ( .A(p_input[1633]), .B(p_input[2049]), .Z(n17853) );
  XNOR U17855 ( .A(n17896), .B(n17869), .Z(n17862) );
  XNOR U17856 ( .A(p_input[1647]), .B(n6322), .Z(n17869) );
  XOR U17857 ( .A(n17859), .B(n17868), .Z(n17896) );
  XOR U17858 ( .A(n17897), .B(n17865), .Z(n17868) );
  XOR U17859 ( .A(p_input[1645]), .B(p_input[2061]), .Z(n17865) );
  XOR U17860 ( .A(p_input[1646]), .B(n6324), .Z(n17897) );
  XOR U17861 ( .A(p_input[1641]), .B(p_input[2057]), .Z(n17859) );
  XOR U17862 ( .A(n17877), .B(n17875), .Z(n17857) );
  XNOR U17863 ( .A(n17898), .B(n17882), .Z(n17875) );
  XOR U17864 ( .A(p_input[1640]), .B(p_input[2056]), .Z(n17882) );
  XOR U17865 ( .A(n17872), .B(n17881), .Z(n17898) );
  XOR U17866 ( .A(n17899), .B(n17878), .Z(n17881) );
  XOR U17867 ( .A(p_input[1638]), .B(p_input[2054]), .Z(n17878) );
  XOR U17868 ( .A(p_input[1639]), .B(n7007), .Z(n17899) );
  XOR U17869 ( .A(p_input[1634]), .B(p_input[2050]), .Z(n17872) );
  XNOR U17870 ( .A(n17887), .B(n17886), .Z(n17877) );
  XOR U17871 ( .A(n17900), .B(n17883), .Z(n17886) );
  XOR U17872 ( .A(p_input[1635]), .B(p_input[2051]), .Z(n17883) );
  XOR U17873 ( .A(p_input[1636]), .B(n7009), .Z(n17900) );
  XOR U17874 ( .A(p_input[1637]), .B(p_input[2053]), .Z(n17887) );
  XOR U17875 ( .A(n17901), .B(n17902), .Z(n17786) );
  AND U17876 ( .A(n415), .B(n17903), .Z(n17902) );
  XNOR U17877 ( .A(n17904), .B(n17901), .Z(n17903) );
  XNOR U17878 ( .A(n17905), .B(n17906), .Z(n415) );
  AND U17879 ( .A(n17907), .B(n17908), .Z(n17906) );
  XOR U17880 ( .A(n17799), .B(n17905), .Z(n17908) );
  AND U17881 ( .A(n17909), .B(n17910), .Z(n17799) );
  XNOR U17882 ( .A(n17796), .B(n17905), .Z(n17907) );
  XOR U17883 ( .A(n17911), .B(n17912), .Z(n17796) );
  AND U17884 ( .A(n419), .B(n17913), .Z(n17912) );
  XOR U17885 ( .A(n17914), .B(n17911), .Z(n17913) );
  XOR U17886 ( .A(n17915), .B(n17916), .Z(n17905) );
  AND U17887 ( .A(n17917), .B(n17918), .Z(n17916) );
  XNOR U17888 ( .A(n17915), .B(n17909), .Z(n17918) );
  IV U17889 ( .A(n17814), .Z(n17909) );
  XOR U17890 ( .A(n17919), .B(n17920), .Z(n17814) );
  XOR U17891 ( .A(n17921), .B(n17910), .Z(n17920) );
  AND U17892 ( .A(n17841), .B(n17922), .Z(n17910) );
  AND U17893 ( .A(n17923), .B(n17924), .Z(n17921) );
  XOR U17894 ( .A(n17925), .B(n17919), .Z(n17923) );
  XNOR U17895 ( .A(n17811), .B(n17915), .Z(n17917) );
  XOR U17896 ( .A(n17926), .B(n17927), .Z(n17811) );
  AND U17897 ( .A(n419), .B(n17928), .Z(n17927) );
  XOR U17898 ( .A(n17929), .B(n17926), .Z(n17928) );
  XOR U17899 ( .A(n17930), .B(n17931), .Z(n17915) );
  AND U17900 ( .A(n17932), .B(n17933), .Z(n17931) );
  XNOR U17901 ( .A(n17930), .B(n17841), .Z(n17933) );
  XOR U17902 ( .A(n17934), .B(n17924), .Z(n17841) );
  XNOR U17903 ( .A(n17935), .B(n17919), .Z(n17924) );
  XOR U17904 ( .A(n17936), .B(n17937), .Z(n17919) );
  AND U17905 ( .A(n17938), .B(n17939), .Z(n17937) );
  XOR U17906 ( .A(n17940), .B(n17936), .Z(n17938) );
  XNOR U17907 ( .A(n17941), .B(n17942), .Z(n17935) );
  AND U17908 ( .A(n17943), .B(n17944), .Z(n17942) );
  XOR U17909 ( .A(n17941), .B(n17945), .Z(n17943) );
  XNOR U17910 ( .A(n17925), .B(n17922), .Z(n17934) );
  AND U17911 ( .A(n17946), .B(n17947), .Z(n17922) );
  XOR U17912 ( .A(n17948), .B(n17949), .Z(n17925) );
  AND U17913 ( .A(n17950), .B(n17951), .Z(n17949) );
  XOR U17914 ( .A(n17948), .B(n17952), .Z(n17950) );
  XNOR U17915 ( .A(n17838), .B(n17930), .Z(n17932) );
  XOR U17916 ( .A(n17953), .B(n17954), .Z(n17838) );
  AND U17917 ( .A(n419), .B(n17955), .Z(n17954) );
  XNOR U17918 ( .A(n17956), .B(n17953), .Z(n17955) );
  XOR U17919 ( .A(n17957), .B(n17958), .Z(n17930) );
  AND U17920 ( .A(n17959), .B(n17960), .Z(n17958) );
  XNOR U17921 ( .A(n17957), .B(n17946), .Z(n17960) );
  IV U17922 ( .A(n17891), .Z(n17946) );
  XNOR U17923 ( .A(n17961), .B(n17939), .Z(n17891) );
  XNOR U17924 ( .A(n17962), .B(n17945), .Z(n17939) );
  XNOR U17925 ( .A(n17963), .B(n17964), .Z(n17945) );
  NOR U17926 ( .A(n17965), .B(n17966), .Z(n17964) );
  XOR U17927 ( .A(n17963), .B(n17967), .Z(n17965) );
  XNOR U17928 ( .A(n17944), .B(n17936), .Z(n17962) );
  XOR U17929 ( .A(n17968), .B(n17969), .Z(n17936) );
  AND U17930 ( .A(n17970), .B(n17971), .Z(n17969) );
  XOR U17931 ( .A(n17968), .B(n17972), .Z(n17970) );
  XNOR U17932 ( .A(n17973), .B(n17941), .Z(n17944) );
  XOR U17933 ( .A(n17974), .B(n17975), .Z(n17941) );
  AND U17934 ( .A(n17976), .B(n17977), .Z(n17975) );
  XNOR U17935 ( .A(n17978), .B(n17979), .Z(n17976) );
  IV U17936 ( .A(n17974), .Z(n17978) );
  XNOR U17937 ( .A(n17980), .B(n17981), .Z(n17973) );
  NOR U17938 ( .A(n17982), .B(n17983), .Z(n17981) );
  XNOR U17939 ( .A(n17980), .B(n17984), .Z(n17982) );
  XNOR U17940 ( .A(n17940), .B(n17947), .Z(n17961) );
  NOR U17941 ( .A(n17904), .B(n17985), .Z(n17947) );
  XOR U17942 ( .A(n17952), .B(n17951), .Z(n17940) );
  XNOR U17943 ( .A(n17986), .B(n17948), .Z(n17951) );
  XOR U17944 ( .A(n17987), .B(n17988), .Z(n17948) );
  AND U17945 ( .A(n17989), .B(n17990), .Z(n17988) );
  XNOR U17946 ( .A(n17991), .B(n17992), .Z(n17989) );
  IV U17947 ( .A(n17987), .Z(n17991) );
  XNOR U17948 ( .A(n17993), .B(n17994), .Z(n17986) );
  NOR U17949 ( .A(n17995), .B(n17996), .Z(n17994) );
  XNOR U17950 ( .A(n17993), .B(n17997), .Z(n17995) );
  XOR U17951 ( .A(n17998), .B(n17999), .Z(n17952) );
  NOR U17952 ( .A(n18000), .B(n18001), .Z(n17999) );
  XNOR U17953 ( .A(n17998), .B(n18002), .Z(n18000) );
  XNOR U17954 ( .A(n17888), .B(n17957), .Z(n17959) );
  XOR U17955 ( .A(n18003), .B(n18004), .Z(n17888) );
  AND U17956 ( .A(n419), .B(n18005), .Z(n18004) );
  XOR U17957 ( .A(n18006), .B(n18003), .Z(n18005) );
  AND U17958 ( .A(n17901), .B(n17904), .Z(n17957) );
  XOR U17959 ( .A(n18007), .B(n17985), .Z(n17904) );
  XNOR U17960 ( .A(p_input[1648]), .B(p_input[2048]), .Z(n17985) );
  XNOR U17961 ( .A(n17972), .B(n17971), .Z(n18007) );
  XNOR U17962 ( .A(n18008), .B(n17979), .Z(n17971) );
  XNOR U17963 ( .A(n17967), .B(n17966), .Z(n17979) );
  XNOR U17964 ( .A(n18009), .B(n17963), .Z(n17966) );
  XNOR U17965 ( .A(p_input[1658]), .B(p_input[2058]), .Z(n17963) );
  XOR U17966 ( .A(p_input[1659]), .B(n6319), .Z(n18009) );
  XOR U17967 ( .A(p_input[1660]), .B(p_input[2060]), .Z(n17967) );
  XOR U17968 ( .A(n17977), .B(n18010), .Z(n18008) );
  IV U17969 ( .A(n17968), .Z(n18010) );
  XOR U17970 ( .A(p_input[1649]), .B(p_input[2049]), .Z(n17968) );
  XNOR U17971 ( .A(n18011), .B(n17984), .Z(n17977) );
  XNOR U17972 ( .A(p_input[1663]), .B(n6322), .Z(n17984) );
  XOR U17973 ( .A(n17974), .B(n17983), .Z(n18011) );
  XOR U17974 ( .A(n18012), .B(n17980), .Z(n17983) );
  XOR U17975 ( .A(p_input[1661]), .B(p_input[2061]), .Z(n17980) );
  XOR U17976 ( .A(p_input[1662]), .B(n6324), .Z(n18012) );
  XOR U17977 ( .A(p_input[1657]), .B(p_input[2057]), .Z(n17974) );
  XOR U17978 ( .A(n17992), .B(n17990), .Z(n17972) );
  XNOR U17979 ( .A(n18013), .B(n17997), .Z(n17990) );
  XOR U17980 ( .A(p_input[1656]), .B(p_input[2056]), .Z(n17997) );
  XOR U17981 ( .A(n17987), .B(n17996), .Z(n18013) );
  XOR U17982 ( .A(n18014), .B(n17993), .Z(n17996) );
  XOR U17983 ( .A(p_input[1654]), .B(p_input[2054]), .Z(n17993) );
  XOR U17984 ( .A(p_input[1655]), .B(n7007), .Z(n18014) );
  XOR U17985 ( .A(p_input[1650]), .B(p_input[2050]), .Z(n17987) );
  XNOR U17986 ( .A(n18002), .B(n18001), .Z(n17992) );
  XOR U17987 ( .A(n18015), .B(n17998), .Z(n18001) );
  XOR U17988 ( .A(p_input[1651]), .B(p_input[2051]), .Z(n17998) );
  XOR U17989 ( .A(p_input[1652]), .B(n7009), .Z(n18015) );
  XOR U17990 ( .A(p_input[1653]), .B(p_input[2053]), .Z(n18002) );
  XOR U17991 ( .A(n18016), .B(n18017), .Z(n17901) );
  AND U17992 ( .A(n419), .B(n18018), .Z(n18017) );
  XNOR U17993 ( .A(n18019), .B(n18016), .Z(n18018) );
  XNOR U17994 ( .A(n18020), .B(n18021), .Z(n419) );
  AND U17995 ( .A(n18022), .B(n18023), .Z(n18021) );
  XOR U17996 ( .A(n17914), .B(n18020), .Z(n18023) );
  AND U17997 ( .A(n18024), .B(n18025), .Z(n17914) );
  XNOR U17998 ( .A(n17911), .B(n18020), .Z(n18022) );
  XOR U17999 ( .A(n18026), .B(n18027), .Z(n17911) );
  AND U18000 ( .A(n423), .B(n18028), .Z(n18027) );
  XOR U18001 ( .A(n18029), .B(n18026), .Z(n18028) );
  XOR U18002 ( .A(n18030), .B(n18031), .Z(n18020) );
  AND U18003 ( .A(n18032), .B(n18033), .Z(n18031) );
  XNOR U18004 ( .A(n18030), .B(n18024), .Z(n18033) );
  IV U18005 ( .A(n17929), .Z(n18024) );
  XOR U18006 ( .A(n18034), .B(n18035), .Z(n17929) );
  XOR U18007 ( .A(n18036), .B(n18025), .Z(n18035) );
  AND U18008 ( .A(n17956), .B(n18037), .Z(n18025) );
  AND U18009 ( .A(n18038), .B(n18039), .Z(n18036) );
  XOR U18010 ( .A(n18040), .B(n18034), .Z(n18038) );
  XNOR U18011 ( .A(n17926), .B(n18030), .Z(n18032) );
  XOR U18012 ( .A(n18041), .B(n18042), .Z(n17926) );
  AND U18013 ( .A(n423), .B(n18043), .Z(n18042) );
  XOR U18014 ( .A(n18044), .B(n18041), .Z(n18043) );
  XOR U18015 ( .A(n18045), .B(n18046), .Z(n18030) );
  AND U18016 ( .A(n18047), .B(n18048), .Z(n18046) );
  XNOR U18017 ( .A(n18045), .B(n17956), .Z(n18048) );
  XOR U18018 ( .A(n18049), .B(n18039), .Z(n17956) );
  XNOR U18019 ( .A(n18050), .B(n18034), .Z(n18039) );
  XOR U18020 ( .A(n18051), .B(n18052), .Z(n18034) );
  AND U18021 ( .A(n18053), .B(n18054), .Z(n18052) );
  XOR U18022 ( .A(n18055), .B(n18051), .Z(n18053) );
  XNOR U18023 ( .A(n18056), .B(n18057), .Z(n18050) );
  AND U18024 ( .A(n18058), .B(n18059), .Z(n18057) );
  XOR U18025 ( .A(n18056), .B(n18060), .Z(n18058) );
  XNOR U18026 ( .A(n18040), .B(n18037), .Z(n18049) );
  AND U18027 ( .A(n18061), .B(n18062), .Z(n18037) );
  XOR U18028 ( .A(n18063), .B(n18064), .Z(n18040) );
  AND U18029 ( .A(n18065), .B(n18066), .Z(n18064) );
  XOR U18030 ( .A(n18063), .B(n18067), .Z(n18065) );
  XNOR U18031 ( .A(n17953), .B(n18045), .Z(n18047) );
  XOR U18032 ( .A(n18068), .B(n18069), .Z(n17953) );
  AND U18033 ( .A(n423), .B(n18070), .Z(n18069) );
  XNOR U18034 ( .A(n18071), .B(n18068), .Z(n18070) );
  XOR U18035 ( .A(n18072), .B(n18073), .Z(n18045) );
  AND U18036 ( .A(n18074), .B(n18075), .Z(n18073) );
  XNOR U18037 ( .A(n18072), .B(n18061), .Z(n18075) );
  IV U18038 ( .A(n18006), .Z(n18061) );
  XNOR U18039 ( .A(n18076), .B(n18054), .Z(n18006) );
  XNOR U18040 ( .A(n18077), .B(n18060), .Z(n18054) );
  XNOR U18041 ( .A(n18078), .B(n18079), .Z(n18060) );
  NOR U18042 ( .A(n18080), .B(n18081), .Z(n18079) );
  XOR U18043 ( .A(n18078), .B(n18082), .Z(n18080) );
  XNOR U18044 ( .A(n18059), .B(n18051), .Z(n18077) );
  XOR U18045 ( .A(n18083), .B(n18084), .Z(n18051) );
  AND U18046 ( .A(n18085), .B(n18086), .Z(n18084) );
  XOR U18047 ( .A(n18083), .B(n18087), .Z(n18085) );
  XNOR U18048 ( .A(n18088), .B(n18056), .Z(n18059) );
  XOR U18049 ( .A(n18089), .B(n18090), .Z(n18056) );
  AND U18050 ( .A(n18091), .B(n18092), .Z(n18090) );
  XNOR U18051 ( .A(n18093), .B(n18094), .Z(n18091) );
  IV U18052 ( .A(n18089), .Z(n18093) );
  XNOR U18053 ( .A(n18095), .B(n18096), .Z(n18088) );
  NOR U18054 ( .A(n18097), .B(n18098), .Z(n18096) );
  XNOR U18055 ( .A(n18095), .B(n18099), .Z(n18097) );
  XNOR U18056 ( .A(n18055), .B(n18062), .Z(n18076) );
  NOR U18057 ( .A(n18019), .B(n18100), .Z(n18062) );
  XOR U18058 ( .A(n18067), .B(n18066), .Z(n18055) );
  XNOR U18059 ( .A(n18101), .B(n18063), .Z(n18066) );
  XOR U18060 ( .A(n18102), .B(n18103), .Z(n18063) );
  AND U18061 ( .A(n18104), .B(n18105), .Z(n18103) );
  XNOR U18062 ( .A(n18106), .B(n18107), .Z(n18104) );
  IV U18063 ( .A(n18102), .Z(n18106) );
  XNOR U18064 ( .A(n18108), .B(n18109), .Z(n18101) );
  NOR U18065 ( .A(n18110), .B(n18111), .Z(n18109) );
  XNOR U18066 ( .A(n18108), .B(n18112), .Z(n18110) );
  XOR U18067 ( .A(n18113), .B(n18114), .Z(n18067) );
  NOR U18068 ( .A(n18115), .B(n18116), .Z(n18114) );
  XNOR U18069 ( .A(n18113), .B(n18117), .Z(n18115) );
  XNOR U18070 ( .A(n18003), .B(n18072), .Z(n18074) );
  XOR U18071 ( .A(n18118), .B(n18119), .Z(n18003) );
  AND U18072 ( .A(n423), .B(n18120), .Z(n18119) );
  XOR U18073 ( .A(n18121), .B(n18118), .Z(n18120) );
  AND U18074 ( .A(n18016), .B(n18019), .Z(n18072) );
  XOR U18075 ( .A(n18122), .B(n18100), .Z(n18019) );
  XNOR U18076 ( .A(p_input[1664]), .B(p_input[2048]), .Z(n18100) );
  XNOR U18077 ( .A(n18087), .B(n18086), .Z(n18122) );
  XNOR U18078 ( .A(n18123), .B(n18094), .Z(n18086) );
  XNOR U18079 ( .A(n18082), .B(n18081), .Z(n18094) );
  XNOR U18080 ( .A(n18124), .B(n18078), .Z(n18081) );
  XNOR U18081 ( .A(p_input[1674]), .B(p_input[2058]), .Z(n18078) );
  XOR U18082 ( .A(p_input[1675]), .B(n6319), .Z(n18124) );
  XOR U18083 ( .A(p_input[1676]), .B(p_input[2060]), .Z(n18082) );
  XOR U18084 ( .A(n18092), .B(n18125), .Z(n18123) );
  IV U18085 ( .A(n18083), .Z(n18125) );
  XOR U18086 ( .A(p_input[1665]), .B(p_input[2049]), .Z(n18083) );
  XNOR U18087 ( .A(n18126), .B(n18099), .Z(n18092) );
  XNOR U18088 ( .A(p_input[1679]), .B(n6322), .Z(n18099) );
  XOR U18089 ( .A(n18089), .B(n18098), .Z(n18126) );
  XOR U18090 ( .A(n18127), .B(n18095), .Z(n18098) );
  XOR U18091 ( .A(p_input[1677]), .B(p_input[2061]), .Z(n18095) );
  XOR U18092 ( .A(p_input[1678]), .B(n6324), .Z(n18127) );
  XOR U18093 ( .A(p_input[1673]), .B(p_input[2057]), .Z(n18089) );
  XOR U18094 ( .A(n18107), .B(n18105), .Z(n18087) );
  XNOR U18095 ( .A(n18128), .B(n18112), .Z(n18105) );
  XOR U18096 ( .A(p_input[1672]), .B(p_input[2056]), .Z(n18112) );
  XOR U18097 ( .A(n18102), .B(n18111), .Z(n18128) );
  XOR U18098 ( .A(n18129), .B(n18108), .Z(n18111) );
  XOR U18099 ( .A(p_input[1670]), .B(p_input[2054]), .Z(n18108) );
  XOR U18100 ( .A(p_input[1671]), .B(n7007), .Z(n18129) );
  XOR U18101 ( .A(p_input[1666]), .B(p_input[2050]), .Z(n18102) );
  XNOR U18102 ( .A(n18117), .B(n18116), .Z(n18107) );
  XOR U18103 ( .A(n18130), .B(n18113), .Z(n18116) );
  XOR U18104 ( .A(p_input[1667]), .B(p_input[2051]), .Z(n18113) );
  XOR U18105 ( .A(p_input[1668]), .B(n7009), .Z(n18130) );
  XOR U18106 ( .A(p_input[1669]), .B(p_input[2053]), .Z(n18117) );
  XOR U18107 ( .A(n18131), .B(n18132), .Z(n18016) );
  AND U18108 ( .A(n423), .B(n18133), .Z(n18132) );
  XNOR U18109 ( .A(n18134), .B(n18131), .Z(n18133) );
  XNOR U18110 ( .A(n18135), .B(n18136), .Z(n423) );
  AND U18111 ( .A(n18137), .B(n18138), .Z(n18136) );
  XOR U18112 ( .A(n18029), .B(n18135), .Z(n18138) );
  AND U18113 ( .A(n18139), .B(n18140), .Z(n18029) );
  XNOR U18114 ( .A(n18026), .B(n18135), .Z(n18137) );
  XOR U18115 ( .A(n18141), .B(n18142), .Z(n18026) );
  AND U18116 ( .A(n427), .B(n18143), .Z(n18142) );
  XOR U18117 ( .A(n18144), .B(n18141), .Z(n18143) );
  XOR U18118 ( .A(n18145), .B(n18146), .Z(n18135) );
  AND U18119 ( .A(n18147), .B(n18148), .Z(n18146) );
  XNOR U18120 ( .A(n18145), .B(n18139), .Z(n18148) );
  IV U18121 ( .A(n18044), .Z(n18139) );
  XOR U18122 ( .A(n18149), .B(n18150), .Z(n18044) );
  XOR U18123 ( .A(n18151), .B(n18140), .Z(n18150) );
  AND U18124 ( .A(n18071), .B(n18152), .Z(n18140) );
  AND U18125 ( .A(n18153), .B(n18154), .Z(n18151) );
  XOR U18126 ( .A(n18155), .B(n18149), .Z(n18153) );
  XNOR U18127 ( .A(n18041), .B(n18145), .Z(n18147) );
  XOR U18128 ( .A(n18156), .B(n18157), .Z(n18041) );
  AND U18129 ( .A(n427), .B(n18158), .Z(n18157) );
  XOR U18130 ( .A(n18159), .B(n18156), .Z(n18158) );
  XOR U18131 ( .A(n18160), .B(n18161), .Z(n18145) );
  AND U18132 ( .A(n18162), .B(n18163), .Z(n18161) );
  XNOR U18133 ( .A(n18160), .B(n18071), .Z(n18163) );
  XOR U18134 ( .A(n18164), .B(n18154), .Z(n18071) );
  XNOR U18135 ( .A(n18165), .B(n18149), .Z(n18154) );
  XOR U18136 ( .A(n18166), .B(n18167), .Z(n18149) );
  AND U18137 ( .A(n18168), .B(n18169), .Z(n18167) );
  XOR U18138 ( .A(n18170), .B(n18166), .Z(n18168) );
  XNOR U18139 ( .A(n18171), .B(n18172), .Z(n18165) );
  AND U18140 ( .A(n18173), .B(n18174), .Z(n18172) );
  XOR U18141 ( .A(n18171), .B(n18175), .Z(n18173) );
  XNOR U18142 ( .A(n18155), .B(n18152), .Z(n18164) );
  AND U18143 ( .A(n18176), .B(n18177), .Z(n18152) );
  XOR U18144 ( .A(n18178), .B(n18179), .Z(n18155) );
  AND U18145 ( .A(n18180), .B(n18181), .Z(n18179) );
  XOR U18146 ( .A(n18178), .B(n18182), .Z(n18180) );
  XNOR U18147 ( .A(n18068), .B(n18160), .Z(n18162) );
  XOR U18148 ( .A(n18183), .B(n18184), .Z(n18068) );
  AND U18149 ( .A(n427), .B(n18185), .Z(n18184) );
  XNOR U18150 ( .A(n18186), .B(n18183), .Z(n18185) );
  XOR U18151 ( .A(n18187), .B(n18188), .Z(n18160) );
  AND U18152 ( .A(n18189), .B(n18190), .Z(n18188) );
  XNOR U18153 ( .A(n18187), .B(n18176), .Z(n18190) );
  IV U18154 ( .A(n18121), .Z(n18176) );
  XNOR U18155 ( .A(n18191), .B(n18169), .Z(n18121) );
  XNOR U18156 ( .A(n18192), .B(n18175), .Z(n18169) );
  XNOR U18157 ( .A(n18193), .B(n18194), .Z(n18175) );
  NOR U18158 ( .A(n18195), .B(n18196), .Z(n18194) );
  XOR U18159 ( .A(n18193), .B(n18197), .Z(n18195) );
  XNOR U18160 ( .A(n18174), .B(n18166), .Z(n18192) );
  XOR U18161 ( .A(n18198), .B(n18199), .Z(n18166) );
  AND U18162 ( .A(n18200), .B(n18201), .Z(n18199) );
  XOR U18163 ( .A(n18198), .B(n18202), .Z(n18200) );
  XNOR U18164 ( .A(n18203), .B(n18171), .Z(n18174) );
  XOR U18165 ( .A(n18204), .B(n18205), .Z(n18171) );
  AND U18166 ( .A(n18206), .B(n18207), .Z(n18205) );
  XNOR U18167 ( .A(n18208), .B(n18209), .Z(n18206) );
  IV U18168 ( .A(n18204), .Z(n18208) );
  XNOR U18169 ( .A(n18210), .B(n18211), .Z(n18203) );
  NOR U18170 ( .A(n18212), .B(n18213), .Z(n18211) );
  XNOR U18171 ( .A(n18210), .B(n18214), .Z(n18212) );
  XNOR U18172 ( .A(n18170), .B(n18177), .Z(n18191) );
  NOR U18173 ( .A(n18134), .B(n18215), .Z(n18177) );
  XOR U18174 ( .A(n18182), .B(n18181), .Z(n18170) );
  XNOR U18175 ( .A(n18216), .B(n18178), .Z(n18181) );
  XOR U18176 ( .A(n18217), .B(n18218), .Z(n18178) );
  AND U18177 ( .A(n18219), .B(n18220), .Z(n18218) );
  XNOR U18178 ( .A(n18221), .B(n18222), .Z(n18219) );
  IV U18179 ( .A(n18217), .Z(n18221) );
  XNOR U18180 ( .A(n18223), .B(n18224), .Z(n18216) );
  NOR U18181 ( .A(n18225), .B(n18226), .Z(n18224) );
  XNOR U18182 ( .A(n18223), .B(n18227), .Z(n18225) );
  XOR U18183 ( .A(n18228), .B(n18229), .Z(n18182) );
  NOR U18184 ( .A(n18230), .B(n18231), .Z(n18229) );
  XNOR U18185 ( .A(n18228), .B(n18232), .Z(n18230) );
  XNOR U18186 ( .A(n18118), .B(n18187), .Z(n18189) );
  XOR U18187 ( .A(n18233), .B(n18234), .Z(n18118) );
  AND U18188 ( .A(n427), .B(n18235), .Z(n18234) );
  XOR U18189 ( .A(n18236), .B(n18233), .Z(n18235) );
  AND U18190 ( .A(n18131), .B(n18134), .Z(n18187) );
  XOR U18191 ( .A(n18237), .B(n18215), .Z(n18134) );
  XNOR U18192 ( .A(p_input[1680]), .B(p_input[2048]), .Z(n18215) );
  XNOR U18193 ( .A(n18202), .B(n18201), .Z(n18237) );
  XNOR U18194 ( .A(n18238), .B(n18209), .Z(n18201) );
  XNOR U18195 ( .A(n18197), .B(n18196), .Z(n18209) );
  XNOR U18196 ( .A(n18239), .B(n18193), .Z(n18196) );
  XNOR U18197 ( .A(p_input[1690]), .B(p_input[2058]), .Z(n18193) );
  XOR U18198 ( .A(p_input[1691]), .B(n6319), .Z(n18239) );
  XOR U18199 ( .A(p_input[1692]), .B(p_input[2060]), .Z(n18197) );
  XOR U18200 ( .A(n18207), .B(n18240), .Z(n18238) );
  IV U18201 ( .A(n18198), .Z(n18240) );
  XOR U18202 ( .A(p_input[1681]), .B(p_input[2049]), .Z(n18198) );
  XNOR U18203 ( .A(n18241), .B(n18214), .Z(n18207) );
  XNOR U18204 ( .A(p_input[1695]), .B(n6322), .Z(n18214) );
  XOR U18205 ( .A(n18204), .B(n18213), .Z(n18241) );
  XOR U18206 ( .A(n18242), .B(n18210), .Z(n18213) );
  XOR U18207 ( .A(p_input[1693]), .B(p_input[2061]), .Z(n18210) );
  XOR U18208 ( .A(p_input[1694]), .B(n6324), .Z(n18242) );
  XOR U18209 ( .A(p_input[1689]), .B(p_input[2057]), .Z(n18204) );
  XOR U18210 ( .A(n18222), .B(n18220), .Z(n18202) );
  XNOR U18211 ( .A(n18243), .B(n18227), .Z(n18220) );
  XOR U18212 ( .A(p_input[1688]), .B(p_input[2056]), .Z(n18227) );
  XOR U18213 ( .A(n18217), .B(n18226), .Z(n18243) );
  XOR U18214 ( .A(n18244), .B(n18223), .Z(n18226) );
  XOR U18215 ( .A(p_input[1686]), .B(p_input[2054]), .Z(n18223) );
  XOR U18216 ( .A(p_input[1687]), .B(n7007), .Z(n18244) );
  XOR U18217 ( .A(p_input[1682]), .B(p_input[2050]), .Z(n18217) );
  XNOR U18218 ( .A(n18232), .B(n18231), .Z(n18222) );
  XOR U18219 ( .A(n18245), .B(n18228), .Z(n18231) );
  XOR U18220 ( .A(p_input[1683]), .B(p_input[2051]), .Z(n18228) );
  XOR U18221 ( .A(p_input[1684]), .B(n7009), .Z(n18245) );
  XOR U18222 ( .A(p_input[1685]), .B(p_input[2053]), .Z(n18232) );
  XOR U18223 ( .A(n18246), .B(n18247), .Z(n18131) );
  AND U18224 ( .A(n427), .B(n18248), .Z(n18247) );
  XNOR U18225 ( .A(n18249), .B(n18246), .Z(n18248) );
  XNOR U18226 ( .A(n18250), .B(n18251), .Z(n427) );
  AND U18227 ( .A(n18252), .B(n18253), .Z(n18251) );
  XOR U18228 ( .A(n18144), .B(n18250), .Z(n18253) );
  AND U18229 ( .A(n18254), .B(n18255), .Z(n18144) );
  XNOR U18230 ( .A(n18141), .B(n18250), .Z(n18252) );
  XOR U18231 ( .A(n18256), .B(n18257), .Z(n18141) );
  AND U18232 ( .A(n431), .B(n18258), .Z(n18257) );
  XOR U18233 ( .A(n18259), .B(n18256), .Z(n18258) );
  XOR U18234 ( .A(n18260), .B(n18261), .Z(n18250) );
  AND U18235 ( .A(n18262), .B(n18263), .Z(n18261) );
  XNOR U18236 ( .A(n18260), .B(n18254), .Z(n18263) );
  IV U18237 ( .A(n18159), .Z(n18254) );
  XOR U18238 ( .A(n18264), .B(n18265), .Z(n18159) );
  XOR U18239 ( .A(n18266), .B(n18255), .Z(n18265) );
  AND U18240 ( .A(n18186), .B(n18267), .Z(n18255) );
  AND U18241 ( .A(n18268), .B(n18269), .Z(n18266) );
  XOR U18242 ( .A(n18270), .B(n18264), .Z(n18268) );
  XNOR U18243 ( .A(n18156), .B(n18260), .Z(n18262) );
  XOR U18244 ( .A(n18271), .B(n18272), .Z(n18156) );
  AND U18245 ( .A(n431), .B(n18273), .Z(n18272) );
  XOR U18246 ( .A(n18274), .B(n18271), .Z(n18273) );
  XOR U18247 ( .A(n18275), .B(n18276), .Z(n18260) );
  AND U18248 ( .A(n18277), .B(n18278), .Z(n18276) );
  XNOR U18249 ( .A(n18275), .B(n18186), .Z(n18278) );
  XOR U18250 ( .A(n18279), .B(n18269), .Z(n18186) );
  XNOR U18251 ( .A(n18280), .B(n18264), .Z(n18269) );
  XOR U18252 ( .A(n18281), .B(n18282), .Z(n18264) );
  AND U18253 ( .A(n18283), .B(n18284), .Z(n18282) );
  XOR U18254 ( .A(n18285), .B(n18281), .Z(n18283) );
  XNOR U18255 ( .A(n18286), .B(n18287), .Z(n18280) );
  AND U18256 ( .A(n18288), .B(n18289), .Z(n18287) );
  XOR U18257 ( .A(n18286), .B(n18290), .Z(n18288) );
  XNOR U18258 ( .A(n18270), .B(n18267), .Z(n18279) );
  AND U18259 ( .A(n18291), .B(n18292), .Z(n18267) );
  XOR U18260 ( .A(n18293), .B(n18294), .Z(n18270) );
  AND U18261 ( .A(n18295), .B(n18296), .Z(n18294) );
  XOR U18262 ( .A(n18293), .B(n18297), .Z(n18295) );
  XNOR U18263 ( .A(n18183), .B(n18275), .Z(n18277) );
  XOR U18264 ( .A(n18298), .B(n18299), .Z(n18183) );
  AND U18265 ( .A(n431), .B(n18300), .Z(n18299) );
  XNOR U18266 ( .A(n18301), .B(n18298), .Z(n18300) );
  XOR U18267 ( .A(n18302), .B(n18303), .Z(n18275) );
  AND U18268 ( .A(n18304), .B(n18305), .Z(n18303) );
  XNOR U18269 ( .A(n18302), .B(n18291), .Z(n18305) );
  IV U18270 ( .A(n18236), .Z(n18291) );
  XNOR U18271 ( .A(n18306), .B(n18284), .Z(n18236) );
  XNOR U18272 ( .A(n18307), .B(n18290), .Z(n18284) );
  XNOR U18273 ( .A(n18308), .B(n18309), .Z(n18290) );
  NOR U18274 ( .A(n18310), .B(n18311), .Z(n18309) );
  XOR U18275 ( .A(n18308), .B(n18312), .Z(n18310) );
  XNOR U18276 ( .A(n18289), .B(n18281), .Z(n18307) );
  XOR U18277 ( .A(n18313), .B(n18314), .Z(n18281) );
  AND U18278 ( .A(n18315), .B(n18316), .Z(n18314) );
  XOR U18279 ( .A(n18313), .B(n18317), .Z(n18315) );
  XNOR U18280 ( .A(n18318), .B(n18286), .Z(n18289) );
  XOR U18281 ( .A(n18319), .B(n18320), .Z(n18286) );
  AND U18282 ( .A(n18321), .B(n18322), .Z(n18320) );
  XNOR U18283 ( .A(n18323), .B(n18324), .Z(n18321) );
  IV U18284 ( .A(n18319), .Z(n18323) );
  XNOR U18285 ( .A(n18325), .B(n18326), .Z(n18318) );
  NOR U18286 ( .A(n18327), .B(n18328), .Z(n18326) );
  XNOR U18287 ( .A(n18325), .B(n18329), .Z(n18327) );
  XNOR U18288 ( .A(n18285), .B(n18292), .Z(n18306) );
  NOR U18289 ( .A(n18249), .B(n18330), .Z(n18292) );
  XOR U18290 ( .A(n18297), .B(n18296), .Z(n18285) );
  XNOR U18291 ( .A(n18331), .B(n18293), .Z(n18296) );
  XOR U18292 ( .A(n18332), .B(n18333), .Z(n18293) );
  AND U18293 ( .A(n18334), .B(n18335), .Z(n18333) );
  XNOR U18294 ( .A(n18336), .B(n18337), .Z(n18334) );
  IV U18295 ( .A(n18332), .Z(n18336) );
  XNOR U18296 ( .A(n18338), .B(n18339), .Z(n18331) );
  NOR U18297 ( .A(n18340), .B(n18341), .Z(n18339) );
  XNOR U18298 ( .A(n18338), .B(n18342), .Z(n18340) );
  XOR U18299 ( .A(n18343), .B(n18344), .Z(n18297) );
  NOR U18300 ( .A(n18345), .B(n18346), .Z(n18344) );
  XNOR U18301 ( .A(n18343), .B(n18347), .Z(n18345) );
  XNOR U18302 ( .A(n18233), .B(n18302), .Z(n18304) );
  XOR U18303 ( .A(n18348), .B(n18349), .Z(n18233) );
  AND U18304 ( .A(n431), .B(n18350), .Z(n18349) );
  XOR U18305 ( .A(n18351), .B(n18348), .Z(n18350) );
  AND U18306 ( .A(n18246), .B(n18249), .Z(n18302) );
  XOR U18307 ( .A(n18352), .B(n18330), .Z(n18249) );
  XNOR U18308 ( .A(p_input[1696]), .B(p_input[2048]), .Z(n18330) );
  XNOR U18309 ( .A(n18317), .B(n18316), .Z(n18352) );
  XNOR U18310 ( .A(n18353), .B(n18324), .Z(n18316) );
  XNOR U18311 ( .A(n18312), .B(n18311), .Z(n18324) );
  XNOR U18312 ( .A(n18354), .B(n18308), .Z(n18311) );
  XNOR U18313 ( .A(p_input[1706]), .B(p_input[2058]), .Z(n18308) );
  XOR U18314 ( .A(p_input[1707]), .B(n6319), .Z(n18354) );
  XOR U18315 ( .A(p_input[1708]), .B(p_input[2060]), .Z(n18312) );
  XOR U18316 ( .A(n18322), .B(n18355), .Z(n18353) );
  IV U18317 ( .A(n18313), .Z(n18355) );
  XOR U18318 ( .A(p_input[1697]), .B(p_input[2049]), .Z(n18313) );
  XNOR U18319 ( .A(n18356), .B(n18329), .Z(n18322) );
  XNOR U18320 ( .A(p_input[1711]), .B(n6322), .Z(n18329) );
  XOR U18321 ( .A(n18319), .B(n18328), .Z(n18356) );
  XOR U18322 ( .A(n18357), .B(n18325), .Z(n18328) );
  XOR U18323 ( .A(p_input[1709]), .B(p_input[2061]), .Z(n18325) );
  XOR U18324 ( .A(p_input[1710]), .B(n6324), .Z(n18357) );
  XOR U18325 ( .A(p_input[1705]), .B(p_input[2057]), .Z(n18319) );
  XOR U18326 ( .A(n18337), .B(n18335), .Z(n18317) );
  XNOR U18327 ( .A(n18358), .B(n18342), .Z(n18335) );
  XOR U18328 ( .A(p_input[1704]), .B(p_input[2056]), .Z(n18342) );
  XOR U18329 ( .A(n18332), .B(n18341), .Z(n18358) );
  XOR U18330 ( .A(n18359), .B(n18338), .Z(n18341) );
  XOR U18331 ( .A(p_input[1702]), .B(p_input[2054]), .Z(n18338) );
  XOR U18332 ( .A(p_input[1703]), .B(n7007), .Z(n18359) );
  XOR U18333 ( .A(p_input[1698]), .B(p_input[2050]), .Z(n18332) );
  XNOR U18334 ( .A(n18347), .B(n18346), .Z(n18337) );
  XOR U18335 ( .A(n18360), .B(n18343), .Z(n18346) );
  XOR U18336 ( .A(p_input[1699]), .B(p_input[2051]), .Z(n18343) );
  XOR U18337 ( .A(p_input[1700]), .B(n7009), .Z(n18360) );
  XOR U18338 ( .A(p_input[1701]), .B(p_input[2053]), .Z(n18347) );
  XOR U18339 ( .A(n18361), .B(n18362), .Z(n18246) );
  AND U18340 ( .A(n431), .B(n18363), .Z(n18362) );
  XNOR U18341 ( .A(n18364), .B(n18361), .Z(n18363) );
  XNOR U18342 ( .A(n18365), .B(n18366), .Z(n431) );
  AND U18343 ( .A(n18367), .B(n18368), .Z(n18366) );
  XOR U18344 ( .A(n18259), .B(n18365), .Z(n18368) );
  AND U18345 ( .A(n18369), .B(n18370), .Z(n18259) );
  XNOR U18346 ( .A(n18256), .B(n18365), .Z(n18367) );
  XOR U18347 ( .A(n18371), .B(n18372), .Z(n18256) );
  AND U18348 ( .A(n435), .B(n18373), .Z(n18372) );
  XOR U18349 ( .A(n18374), .B(n18371), .Z(n18373) );
  XOR U18350 ( .A(n18375), .B(n18376), .Z(n18365) );
  AND U18351 ( .A(n18377), .B(n18378), .Z(n18376) );
  XNOR U18352 ( .A(n18375), .B(n18369), .Z(n18378) );
  IV U18353 ( .A(n18274), .Z(n18369) );
  XOR U18354 ( .A(n18379), .B(n18380), .Z(n18274) );
  XOR U18355 ( .A(n18381), .B(n18370), .Z(n18380) );
  AND U18356 ( .A(n18301), .B(n18382), .Z(n18370) );
  AND U18357 ( .A(n18383), .B(n18384), .Z(n18381) );
  XOR U18358 ( .A(n18385), .B(n18379), .Z(n18383) );
  XNOR U18359 ( .A(n18271), .B(n18375), .Z(n18377) );
  XOR U18360 ( .A(n18386), .B(n18387), .Z(n18271) );
  AND U18361 ( .A(n435), .B(n18388), .Z(n18387) );
  XOR U18362 ( .A(n18389), .B(n18386), .Z(n18388) );
  XOR U18363 ( .A(n18390), .B(n18391), .Z(n18375) );
  AND U18364 ( .A(n18392), .B(n18393), .Z(n18391) );
  XNOR U18365 ( .A(n18390), .B(n18301), .Z(n18393) );
  XOR U18366 ( .A(n18394), .B(n18384), .Z(n18301) );
  XNOR U18367 ( .A(n18395), .B(n18379), .Z(n18384) );
  XOR U18368 ( .A(n18396), .B(n18397), .Z(n18379) );
  AND U18369 ( .A(n18398), .B(n18399), .Z(n18397) );
  XOR U18370 ( .A(n18400), .B(n18396), .Z(n18398) );
  XNOR U18371 ( .A(n18401), .B(n18402), .Z(n18395) );
  AND U18372 ( .A(n18403), .B(n18404), .Z(n18402) );
  XOR U18373 ( .A(n18401), .B(n18405), .Z(n18403) );
  XNOR U18374 ( .A(n18385), .B(n18382), .Z(n18394) );
  AND U18375 ( .A(n18406), .B(n18407), .Z(n18382) );
  XOR U18376 ( .A(n18408), .B(n18409), .Z(n18385) );
  AND U18377 ( .A(n18410), .B(n18411), .Z(n18409) );
  XOR U18378 ( .A(n18408), .B(n18412), .Z(n18410) );
  XNOR U18379 ( .A(n18298), .B(n18390), .Z(n18392) );
  XOR U18380 ( .A(n18413), .B(n18414), .Z(n18298) );
  AND U18381 ( .A(n435), .B(n18415), .Z(n18414) );
  XNOR U18382 ( .A(n18416), .B(n18413), .Z(n18415) );
  XOR U18383 ( .A(n18417), .B(n18418), .Z(n18390) );
  AND U18384 ( .A(n18419), .B(n18420), .Z(n18418) );
  XNOR U18385 ( .A(n18417), .B(n18406), .Z(n18420) );
  IV U18386 ( .A(n18351), .Z(n18406) );
  XNOR U18387 ( .A(n18421), .B(n18399), .Z(n18351) );
  XNOR U18388 ( .A(n18422), .B(n18405), .Z(n18399) );
  XNOR U18389 ( .A(n18423), .B(n18424), .Z(n18405) );
  NOR U18390 ( .A(n18425), .B(n18426), .Z(n18424) );
  XOR U18391 ( .A(n18423), .B(n18427), .Z(n18425) );
  XNOR U18392 ( .A(n18404), .B(n18396), .Z(n18422) );
  XOR U18393 ( .A(n18428), .B(n18429), .Z(n18396) );
  AND U18394 ( .A(n18430), .B(n18431), .Z(n18429) );
  XOR U18395 ( .A(n18428), .B(n18432), .Z(n18430) );
  XNOR U18396 ( .A(n18433), .B(n18401), .Z(n18404) );
  XOR U18397 ( .A(n18434), .B(n18435), .Z(n18401) );
  AND U18398 ( .A(n18436), .B(n18437), .Z(n18435) );
  XNOR U18399 ( .A(n18438), .B(n18439), .Z(n18436) );
  IV U18400 ( .A(n18434), .Z(n18438) );
  XNOR U18401 ( .A(n18440), .B(n18441), .Z(n18433) );
  NOR U18402 ( .A(n18442), .B(n18443), .Z(n18441) );
  XNOR U18403 ( .A(n18440), .B(n18444), .Z(n18442) );
  XNOR U18404 ( .A(n18400), .B(n18407), .Z(n18421) );
  NOR U18405 ( .A(n18364), .B(n18445), .Z(n18407) );
  XOR U18406 ( .A(n18412), .B(n18411), .Z(n18400) );
  XNOR U18407 ( .A(n18446), .B(n18408), .Z(n18411) );
  XOR U18408 ( .A(n18447), .B(n18448), .Z(n18408) );
  AND U18409 ( .A(n18449), .B(n18450), .Z(n18448) );
  XNOR U18410 ( .A(n18451), .B(n18452), .Z(n18449) );
  IV U18411 ( .A(n18447), .Z(n18451) );
  XNOR U18412 ( .A(n18453), .B(n18454), .Z(n18446) );
  NOR U18413 ( .A(n18455), .B(n18456), .Z(n18454) );
  XNOR U18414 ( .A(n18453), .B(n18457), .Z(n18455) );
  XOR U18415 ( .A(n18458), .B(n18459), .Z(n18412) );
  NOR U18416 ( .A(n18460), .B(n18461), .Z(n18459) );
  XNOR U18417 ( .A(n18458), .B(n18462), .Z(n18460) );
  XNOR U18418 ( .A(n18348), .B(n18417), .Z(n18419) );
  XOR U18419 ( .A(n18463), .B(n18464), .Z(n18348) );
  AND U18420 ( .A(n435), .B(n18465), .Z(n18464) );
  XOR U18421 ( .A(n18466), .B(n18463), .Z(n18465) );
  AND U18422 ( .A(n18361), .B(n18364), .Z(n18417) );
  XOR U18423 ( .A(n18467), .B(n18445), .Z(n18364) );
  XNOR U18424 ( .A(p_input[1712]), .B(p_input[2048]), .Z(n18445) );
  XNOR U18425 ( .A(n18432), .B(n18431), .Z(n18467) );
  XNOR U18426 ( .A(n18468), .B(n18439), .Z(n18431) );
  XNOR U18427 ( .A(n18427), .B(n18426), .Z(n18439) );
  XNOR U18428 ( .A(n18469), .B(n18423), .Z(n18426) );
  XNOR U18429 ( .A(p_input[1722]), .B(p_input[2058]), .Z(n18423) );
  XOR U18430 ( .A(p_input[1723]), .B(n6319), .Z(n18469) );
  XOR U18431 ( .A(p_input[1724]), .B(p_input[2060]), .Z(n18427) );
  XOR U18432 ( .A(n18437), .B(n18470), .Z(n18468) );
  IV U18433 ( .A(n18428), .Z(n18470) );
  XOR U18434 ( .A(p_input[1713]), .B(p_input[2049]), .Z(n18428) );
  XNOR U18435 ( .A(n18471), .B(n18444), .Z(n18437) );
  XNOR U18436 ( .A(p_input[1727]), .B(n6322), .Z(n18444) );
  XOR U18437 ( .A(n18434), .B(n18443), .Z(n18471) );
  XOR U18438 ( .A(n18472), .B(n18440), .Z(n18443) );
  XOR U18439 ( .A(p_input[1725]), .B(p_input[2061]), .Z(n18440) );
  XOR U18440 ( .A(p_input[1726]), .B(n6324), .Z(n18472) );
  XOR U18441 ( .A(p_input[1721]), .B(p_input[2057]), .Z(n18434) );
  XOR U18442 ( .A(n18452), .B(n18450), .Z(n18432) );
  XNOR U18443 ( .A(n18473), .B(n18457), .Z(n18450) );
  XOR U18444 ( .A(p_input[1720]), .B(p_input[2056]), .Z(n18457) );
  XOR U18445 ( .A(n18447), .B(n18456), .Z(n18473) );
  XOR U18446 ( .A(n18474), .B(n18453), .Z(n18456) );
  XOR U18447 ( .A(p_input[1718]), .B(p_input[2054]), .Z(n18453) );
  XOR U18448 ( .A(p_input[1719]), .B(n7007), .Z(n18474) );
  XOR U18449 ( .A(p_input[1714]), .B(p_input[2050]), .Z(n18447) );
  XNOR U18450 ( .A(n18462), .B(n18461), .Z(n18452) );
  XOR U18451 ( .A(n18475), .B(n18458), .Z(n18461) );
  XOR U18452 ( .A(p_input[1715]), .B(p_input[2051]), .Z(n18458) );
  XOR U18453 ( .A(p_input[1716]), .B(n7009), .Z(n18475) );
  XOR U18454 ( .A(p_input[1717]), .B(p_input[2053]), .Z(n18462) );
  XOR U18455 ( .A(n18476), .B(n18477), .Z(n18361) );
  AND U18456 ( .A(n435), .B(n18478), .Z(n18477) );
  XNOR U18457 ( .A(n18479), .B(n18476), .Z(n18478) );
  XNOR U18458 ( .A(n18480), .B(n18481), .Z(n435) );
  AND U18459 ( .A(n18482), .B(n18483), .Z(n18481) );
  XOR U18460 ( .A(n18374), .B(n18480), .Z(n18483) );
  AND U18461 ( .A(n18484), .B(n18485), .Z(n18374) );
  XNOR U18462 ( .A(n18371), .B(n18480), .Z(n18482) );
  XOR U18463 ( .A(n18486), .B(n18487), .Z(n18371) );
  AND U18464 ( .A(n439), .B(n18488), .Z(n18487) );
  XOR U18465 ( .A(n18489), .B(n18486), .Z(n18488) );
  XOR U18466 ( .A(n18490), .B(n18491), .Z(n18480) );
  AND U18467 ( .A(n18492), .B(n18493), .Z(n18491) );
  XNOR U18468 ( .A(n18490), .B(n18484), .Z(n18493) );
  IV U18469 ( .A(n18389), .Z(n18484) );
  XOR U18470 ( .A(n18494), .B(n18495), .Z(n18389) );
  XOR U18471 ( .A(n18496), .B(n18485), .Z(n18495) );
  AND U18472 ( .A(n18416), .B(n18497), .Z(n18485) );
  AND U18473 ( .A(n18498), .B(n18499), .Z(n18496) );
  XOR U18474 ( .A(n18500), .B(n18494), .Z(n18498) );
  XNOR U18475 ( .A(n18386), .B(n18490), .Z(n18492) );
  XOR U18476 ( .A(n18501), .B(n18502), .Z(n18386) );
  AND U18477 ( .A(n439), .B(n18503), .Z(n18502) );
  XOR U18478 ( .A(n18504), .B(n18501), .Z(n18503) );
  XOR U18479 ( .A(n18505), .B(n18506), .Z(n18490) );
  AND U18480 ( .A(n18507), .B(n18508), .Z(n18506) );
  XNOR U18481 ( .A(n18505), .B(n18416), .Z(n18508) );
  XOR U18482 ( .A(n18509), .B(n18499), .Z(n18416) );
  XNOR U18483 ( .A(n18510), .B(n18494), .Z(n18499) );
  XOR U18484 ( .A(n18511), .B(n18512), .Z(n18494) );
  AND U18485 ( .A(n18513), .B(n18514), .Z(n18512) );
  XOR U18486 ( .A(n18515), .B(n18511), .Z(n18513) );
  XNOR U18487 ( .A(n18516), .B(n18517), .Z(n18510) );
  AND U18488 ( .A(n18518), .B(n18519), .Z(n18517) );
  XOR U18489 ( .A(n18516), .B(n18520), .Z(n18518) );
  XNOR U18490 ( .A(n18500), .B(n18497), .Z(n18509) );
  AND U18491 ( .A(n18521), .B(n18522), .Z(n18497) );
  XOR U18492 ( .A(n18523), .B(n18524), .Z(n18500) );
  AND U18493 ( .A(n18525), .B(n18526), .Z(n18524) );
  XOR U18494 ( .A(n18523), .B(n18527), .Z(n18525) );
  XNOR U18495 ( .A(n18413), .B(n18505), .Z(n18507) );
  XOR U18496 ( .A(n18528), .B(n18529), .Z(n18413) );
  AND U18497 ( .A(n439), .B(n18530), .Z(n18529) );
  XNOR U18498 ( .A(n18531), .B(n18528), .Z(n18530) );
  XOR U18499 ( .A(n18532), .B(n18533), .Z(n18505) );
  AND U18500 ( .A(n18534), .B(n18535), .Z(n18533) );
  XNOR U18501 ( .A(n18532), .B(n18521), .Z(n18535) );
  IV U18502 ( .A(n18466), .Z(n18521) );
  XNOR U18503 ( .A(n18536), .B(n18514), .Z(n18466) );
  XNOR U18504 ( .A(n18537), .B(n18520), .Z(n18514) );
  XNOR U18505 ( .A(n18538), .B(n18539), .Z(n18520) );
  NOR U18506 ( .A(n18540), .B(n18541), .Z(n18539) );
  XOR U18507 ( .A(n18538), .B(n18542), .Z(n18540) );
  XNOR U18508 ( .A(n18519), .B(n18511), .Z(n18537) );
  XOR U18509 ( .A(n18543), .B(n18544), .Z(n18511) );
  AND U18510 ( .A(n18545), .B(n18546), .Z(n18544) );
  XOR U18511 ( .A(n18543), .B(n18547), .Z(n18545) );
  XNOR U18512 ( .A(n18548), .B(n18516), .Z(n18519) );
  XOR U18513 ( .A(n18549), .B(n18550), .Z(n18516) );
  AND U18514 ( .A(n18551), .B(n18552), .Z(n18550) );
  XNOR U18515 ( .A(n18553), .B(n18554), .Z(n18551) );
  IV U18516 ( .A(n18549), .Z(n18553) );
  XNOR U18517 ( .A(n18555), .B(n18556), .Z(n18548) );
  NOR U18518 ( .A(n18557), .B(n18558), .Z(n18556) );
  XNOR U18519 ( .A(n18555), .B(n18559), .Z(n18557) );
  XNOR U18520 ( .A(n18515), .B(n18522), .Z(n18536) );
  NOR U18521 ( .A(n18479), .B(n18560), .Z(n18522) );
  XOR U18522 ( .A(n18527), .B(n18526), .Z(n18515) );
  XNOR U18523 ( .A(n18561), .B(n18523), .Z(n18526) );
  XOR U18524 ( .A(n18562), .B(n18563), .Z(n18523) );
  AND U18525 ( .A(n18564), .B(n18565), .Z(n18563) );
  XNOR U18526 ( .A(n18566), .B(n18567), .Z(n18564) );
  IV U18527 ( .A(n18562), .Z(n18566) );
  XNOR U18528 ( .A(n18568), .B(n18569), .Z(n18561) );
  NOR U18529 ( .A(n18570), .B(n18571), .Z(n18569) );
  XNOR U18530 ( .A(n18568), .B(n18572), .Z(n18570) );
  XOR U18531 ( .A(n18573), .B(n18574), .Z(n18527) );
  NOR U18532 ( .A(n18575), .B(n18576), .Z(n18574) );
  XNOR U18533 ( .A(n18573), .B(n18577), .Z(n18575) );
  XNOR U18534 ( .A(n18463), .B(n18532), .Z(n18534) );
  XOR U18535 ( .A(n18578), .B(n18579), .Z(n18463) );
  AND U18536 ( .A(n439), .B(n18580), .Z(n18579) );
  XOR U18537 ( .A(n18581), .B(n18578), .Z(n18580) );
  AND U18538 ( .A(n18476), .B(n18479), .Z(n18532) );
  XOR U18539 ( .A(n18582), .B(n18560), .Z(n18479) );
  XNOR U18540 ( .A(p_input[1728]), .B(p_input[2048]), .Z(n18560) );
  XNOR U18541 ( .A(n18547), .B(n18546), .Z(n18582) );
  XNOR U18542 ( .A(n18583), .B(n18554), .Z(n18546) );
  XNOR U18543 ( .A(n18542), .B(n18541), .Z(n18554) );
  XNOR U18544 ( .A(n18584), .B(n18538), .Z(n18541) );
  XNOR U18545 ( .A(p_input[1738]), .B(p_input[2058]), .Z(n18538) );
  XOR U18546 ( .A(p_input[1739]), .B(n6319), .Z(n18584) );
  XOR U18547 ( .A(p_input[1740]), .B(p_input[2060]), .Z(n18542) );
  XOR U18548 ( .A(n18552), .B(n18585), .Z(n18583) );
  IV U18549 ( .A(n18543), .Z(n18585) );
  XOR U18550 ( .A(p_input[1729]), .B(p_input[2049]), .Z(n18543) );
  XNOR U18551 ( .A(n18586), .B(n18559), .Z(n18552) );
  XNOR U18552 ( .A(p_input[1743]), .B(n6322), .Z(n18559) );
  XOR U18553 ( .A(n18549), .B(n18558), .Z(n18586) );
  XOR U18554 ( .A(n18587), .B(n18555), .Z(n18558) );
  XOR U18555 ( .A(p_input[1741]), .B(p_input[2061]), .Z(n18555) );
  XOR U18556 ( .A(p_input[1742]), .B(n6324), .Z(n18587) );
  XOR U18557 ( .A(p_input[1737]), .B(p_input[2057]), .Z(n18549) );
  XOR U18558 ( .A(n18567), .B(n18565), .Z(n18547) );
  XNOR U18559 ( .A(n18588), .B(n18572), .Z(n18565) );
  XOR U18560 ( .A(p_input[1736]), .B(p_input[2056]), .Z(n18572) );
  XOR U18561 ( .A(n18562), .B(n18571), .Z(n18588) );
  XOR U18562 ( .A(n18589), .B(n18568), .Z(n18571) );
  XOR U18563 ( .A(p_input[1734]), .B(p_input[2054]), .Z(n18568) );
  XOR U18564 ( .A(p_input[1735]), .B(n7007), .Z(n18589) );
  XOR U18565 ( .A(p_input[1730]), .B(p_input[2050]), .Z(n18562) );
  XNOR U18566 ( .A(n18577), .B(n18576), .Z(n18567) );
  XOR U18567 ( .A(n18590), .B(n18573), .Z(n18576) );
  XOR U18568 ( .A(p_input[1731]), .B(p_input[2051]), .Z(n18573) );
  XOR U18569 ( .A(p_input[1732]), .B(n7009), .Z(n18590) );
  XOR U18570 ( .A(p_input[1733]), .B(p_input[2053]), .Z(n18577) );
  XOR U18571 ( .A(n18591), .B(n18592), .Z(n18476) );
  AND U18572 ( .A(n439), .B(n18593), .Z(n18592) );
  XNOR U18573 ( .A(n18594), .B(n18591), .Z(n18593) );
  XNOR U18574 ( .A(n18595), .B(n18596), .Z(n439) );
  AND U18575 ( .A(n18597), .B(n18598), .Z(n18596) );
  XOR U18576 ( .A(n18489), .B(n18595), .Z(n18598) );
  AND U18577 ( .A(n18599), .B(n18600), .Z(n18489) );
  XNOR U18578 ( .A(n18486), .B(n18595), .Z(n18597) );
  XOR U18579 ( .A(n18601), .B(n18602), .Z(n18486) );
  AND U18580 ( .A(n443), .B(n18603), .Z(n18602) );
  XOR U18581 ( .A(n18604), .B(n18601), .Z(n18603) );
  XOR U18582 ( .A(n18605), .B(n18606), .Z(n18595) );
  AND U18583 ( .A(n18607), .B(n18608), .Z(n18606) );
  XNOR U18584 ( .A(n18605), .B(n18599), .Z(n18608) );
  IV U18585 ( .A(n18504), .Z(n18599) );
  XOR U18586 ( .A(n18609), .B(n18610), .Z(n18504) );
  XOR U18587 ( .A(n18611), .B(n18600), .Z(n18610) );
  AND U18588 ( .A(n18531), .B(n18612), .Z(n18600) );
  AND U18589 ( .A(n18613), .B(n18614), .Z(n18611) );
  XOR U18590 ( .A(n18615), .B(n18609), .Z(n18613) );
  XNOR U18591 ( .A(n18501), .B(n18605), .Z(n18607) );
  XOR U18592 ( .A(n18616), .B(n18617), .Z(n18501) );
  AND U18593 ( .A(n443), .B(n18618), .Z(n18617) );
  XOR U18594 ( .A(n18619), .B(n18616), .Z(n18618) );
  XOR U18595 ( .A(n18620), .B(n18621), .Z(n18605) );
  AND U18596 ( .A(n18622), .B(n18623), .Z(n18621) );
  XNOR U18597 ( .A(n18620), .B(n18531), .Z(n18623) );
  XOR U18598 ( .A(n18624), .B(n18614), .Z(n18531) );
  XNOR U18599 ( .A(n18625), .B(n18609), .Z(n18614) );
  XOR U18600 ( .A(n18626), .B(n18627), .Z(n18609) );
  AND U18601 ( .A(n18628), .B(n18629), .Z(n18627) );
  XOR U18602 ( .A(n18630), .B(n18626), .Z(n18628) );
  XNOR U18603 ( .A(n18631), .B(n18632), .Z(n18625) );
  AND U18604 ( .A(n18633), .B(n18634), .Z(n18632) );
  XOR U18605 ( .A(n18631), .B(n18635), .Z(n18633) );
  XNOR U18606 ( .A(n18615), .B(n18612), .Z(n18624) );
  AND U18607 ( .A(n18636), .B(n18637), .Z(n18612) );
  XOR U18608 ( .A(n18638), .B(n18639), .Z(n18615) );
  AND U18609 ( .A(n18640), .B(n18641), .Z(n18639) );
  XOR U18610 ( .A(n18638), .B(n18642), .Z(n18640) );
  XNOR U18611 ( .A(n18528), .B(n18620), .Z(n18622) );
  XOR U18612 ( .A(n18643), .B(n18644), .Z(n18528) );
  AND U18613 ( .A(n443), .B(n18645), .Z(n18644) );
  XNOR U18614 ( .A(n18646), .B(n18643), .Z(n18645) );
  XOR U18615 ( .A(n18647), .B(n18648), .Z(n18620) );
  AND U18616 ( .A(n18649), .B(n18650), .Z(n18648) );
  XNOR U18617 ( .A(n18647), .B(n18636), .Z(n18650) );
  IV U18618 ( .A(n18581), .Z(n18636) );
  XNOR U18619 ( .A(n18651), .B(n18629), .Z(n18581) );
  XNOR U18620 ( .A(n18652), .B(n18635), .Z(n18629) );
  XNOR U18621 ( .A(n18653), .B(n18654), .Z(n18635) );
  NOR U18622 ( .A(n18655), .B(n18656), .Z(n18654) );
  XOR U18623 ( .A(n18653), .B(n18657), .Z(n18655) );
  XNOR U18624 ( .A(n18634), .B(n18626), .Z(n18652) );
  XOR U18625 ( .A(n18658), .B(n18659), .Z(n18626) );
  AND U18626 ( .A(n18660), .B(n18661), .Z(n18659) );
  XOR U18627 ( .A(n18658), .B(n18662), .Z(n18660) );
  XNOR U18628 ( .A(n18663), .B(n18631), .Z(n18634) );
  XOR U18629 ( .A(n18664), .B(n18665), .Z(n18631) );
  AND U18630 ( .A(n18666), .B(n18667), .Z(n18665) );
  XNOR U18631 ( .A(n18668), .B(n18669), .Z(n18666) );
  IV U18632 ( .A(n18664), .Z(n18668) );
  XNOR U18633 ( .A(n18670), .B(n18671), .Z(n18663) );
  NOR U18634 ( .A(n18672), .B(n18673), .Z(n18671) );
  XNOR U18635 ( .A(n18670), .B(n18674), .Z(n18672) );
  XNOR U18636 ( .A(n18630), .B(n18637), .Z(n18651) );
  NOR U18637 ( .A(n18594), .B(n18675), .Z(n18637) );
  XOR U18638 ( .A(n18642), .B(n18641), .Z(n18630) );
  XNOR U18639 ( .A(n18676), .B(n18638), .Z(n18641) );
  XOR U18640 ( .A(n18677), .B(n18678), .Z(n18638) );
  AND U18641 ( .A(n18679), .B(n18680), .Z(n18678) );
  XNOR U18642 ( .A(n18681), .B(n18682), .Z(n18679) );
  IV U18643 ( .A(n18677), .Z(n18681) );
  XNOR U18644 ( .A(n18683), .B(n18684), .Z(n18676) );
  NOR U18645 ( .A(n18685), .B(n18686), .Z(n18684) );
  XNOR U18646 ( .A(n18683), .B(n18687), .Z(n18685) );
  XOR U18647 ( .A(n18688), .B(n18689), .Z(n18642) );
  NOR U18648 ( .A(n18690), .B(n18691), .Z(n18689) );
  XNOR U18649 ( .A(n18688), .B(n18692), .Z(n18690) );
  XNOR U18650 ( .A(n18578), .B(n18647), .Z(n18649) );
  XOR U18651 ( .A(n18693), .B(n18694), .Z(n18578) );
  AND U18652 ( .A(n443), .B(n18695), .Z(n18694) );
  XOR U18653 ( .A(n18696), .B(n18693), .Z(n18695) );
  AND U18654 ( .A(n18591), .B(n18594), .Z(n18647) );
  XOR U18655 ( .A(n18697), .B(n18675), .Z(n18594) );
  XNOR U18656 ( .A(p_input[1744]), .B(p_input[2048]), .Z(n18675) );
  XNOR U18657 ( .A(n18662), .B(n18661), .Z(n18697) );
  XNOR U18658 ( .A(n18698), .B(n18669), .Z(n18661) );
  XNOR U18659 ( .A(n18657), .B(n18656), .Z(n18669) );
  XNOR U18660 ( .A(n18699), .B(n18653), .Z(n18656) );
  XNOR U18661 ( .A(p_input[1754]), .B(p_input[2058]), .Z(n18653) );
  XOR U18662 ( .A(p_input[1755]), .B(n6319), .Z(n18699) );
  XOR U18663 ( .A(p_input[1756]), .B(p_input[2060]), .Z(n18657) );
  XOR U18664 ( .A(n18667), .B(n18700), .Z(n18698) );
  IV U18665 ( .A(n18658), .Z(n18700) );
  XOR U18666 ( .A(p_input[1745]), .B(p_input[2049]), .Z(n18658) );
  XNOR U18667 ( .A(n18701), .B(n18674), .Z(n18667) );
  XNOR U18668 ( .A(p_input[1759]), .B(n6322), .Z(n18674) );
  XOR U18669 ( .A(n18664), .B(n18673), .Z(n18701) );
  XOR U18670 ( .A(n18702), .B(n18670), .Z(n18673) );
  XOR U18671 ( .A(p_input[1757]), .B(p_input[2061]), .Z(n18670) );
  XOR U18672 ( .A(p_input[1758]), .B(n6324), .Z(n18702) );
  XOR U18673 ( .A(p_input[1753]), .B(p_input[2057]), .Z(n18664) );
  XOR U18674 ( .A(n18682), .B(n18680), .Z(n18662) );
  XNOR U18675 ( .A(n18703), .B(n18687), .Z(n18680) );
  XOR U18676 ( .A(p_input[1752]), .B(p_input[2056]), .Z(n18687) );
  XOR U18677 ( .A(n18677), .B(n18686), .Z(n18703) );
  XOR U18678 ( .A(n18704), .B(n18683), .Z(n18686) );
  XOR U18679 ( .A(p_input[1750]), .B(p_input[2054]), .Z(n18683) );
  XOR U18680 ( .A(p_input[1751]), .B(n7007), .Z(n18704) );
  XOR U18681 ( .A(p_input[1746]), .B(p_input[2050]), .Z(n18677) );
  XNOR U18682 ( .A(n18692), .B(n18691), .Z(n18682) );
  XOR U18683 ( .A(n18705), .B(n18688), .Z(n18691) );
  XOR U18684 ( .A(p_input[1747]), .B(p_input[2051]), .Z(n18688) );
  XOR U18685 ( .A(p_input[1748]), .B(n7009), .Z(n18705) );
  XOR U18686 ( .A(p_input[1749]), .B(p_input[2053]), .Z(n18692) );
  XOR U18687 ( .A(n18706), .B(n18707), .Z(n18591) );
  AND U18688 ( .A(n443), .B(n18708), .Z(n18707) );
  XNOR U18689 ( .A(n18709), .B(n18706), .Z(n18708) );
  XNOR U18690 ( .A(n18710), .B(n18711), .Z(n443) );
  AND U18691 ( .A(n18712), .B(n18713), .Z(n18711) );
  XOR U18692 ( .A(n18604), .B(n18710), .Z(n18713) );
  AND U18693 ( .A(n18714), .B(n18715), .Z(n18604) );
  XNOR U18694 ( .A(n18601), .B(n18710), .Z(n18712) );
  XOR U18695 ( .A(n18716), .B(n18717), .Z(n18601) );
  AND U18696 ( .A(n447), .B(n18718), .Z(n18717) );
  XOR U18697 ( .A(n18719), .B(n18716), .Z(n18718) );
  XOR U18698 ( .A(n18720), .B(n18721), .Z(n18710) );
  AND U18699 ( .A(n18722), .B(n18723), .Z(n18721) );
  XNOR U18700 ( .A(n18720), .B(n18714), .Z(n18723) );
  IV U18701 ( .A(n18619), .Z(n18714) );
  XOR U18702 ( .A(n18724), .B(n18725), .Z(n18619) );
  XOR U18703 ( .A(n18726), .B(n18715), .Z(n18725) );
  AND U18704 ( .A(n18646), .B(n18727), .Z(n18715) );
  AND U18705 ( .A(n18728), .B(n18729), .Z(n18726) );
  XOR U18706 ( .A(n18730), .B(n18724), .Z(n18728) );
  XNOR U18707 ( .A(n18616), .B(n18720), .Z(n18722) );
  XOR U18708 ( .A(n18731), .B(n18732), .Z(n18616) );
  AND U18709 ( .A(n447), .B(n18733), .Z(n18732) );
  XOR U18710 ( .A(n18734), .B(n18731), .Z(n18733) );
  XOR U18711 ( .A(n18735), .B(n18736), .Z(n18720) );
  AND U18712 ( .A(n18737), .B(n18738), .Z(n18736) );
  XNOR U18713 ( .A(n18735), .B(n18646), .Z(n18738) );
  XOR U18714 ( .A(n18739), .B(n18729), .Z(n18646) );
  XNOR U18715 ( .A(n18740), .B(n18724), .Z(n18729) );
  XOR U18716 ( .A(n18741), .B(n18742), .Z(n18724) );
  AND U18717 ( .A(n18743), .B(n18744), .Z(n18742) );
  XOR U18718 ( .A(n18745), .B(n18741), .Z(n18743) );
  XNOR U18719 ( .A(n18746), .B(n18747), .Z(n18740) );
  AND U18720 ( .A(n18748), .B(n18749), .Z(n18747) );
  XOR U18721 ( .A(n18746), .B(n18750), .Z(n18748) );
  XNOR U18722 ( .A(n18730), .B(n18727), .Z(n18739) );
  AND U18723 ( .A(n18751), .B(n18752), .Z(n18727) );
  XOR U18724 ( .A(n18753), .B(n18754), .Z(n18730) );
  AND U18725 ( .A(n18755), .B(n18756), .Z(n18754) );
  XOR U18726 ( .A(n18753), .B(n18757), .Z(n18755) );
  XNOR U18727 ( .A(n18643), .B(n18735), .Z(n18737) );
  XOR U18728 ( .A(n18758), .B(n18759), .Z(n18643) );
  AND U18729 ( .A(n447), .B(n18760), .Z(n18759) );
  XNOR U18730 ( .A(n18761), .B(n18758), .Z(n18760) );
  XOR U18731 ( .A(n18762), .B(n18763), .Z(n18735) );
  AND U18732 ( .A(n18764), .B(n18765), .Z(n18763) );
  XNOR U18733 ( .A(n18762), .B(n18751), .Z(n18765) );
  IV U18734 ( .A(n18696), .Z(n18751) );
  XNOR U18735 ( .A(n18766), .B(n18744), .Z(n18696) );
  XNOR U18736 ( .A(n18767), .B(n18750), .Z(n18744) );
  XNOR U18737 ( .A(n18768), .B(n18769), .Z(n18750) );
  NOR U18738 ( .A(n18770), .B(n18771), .Z(n18769) );
  XOR U18739 ( .A(n18768), .B(n18772), .Z(n18770) );
  XNOR U18740 ( .A(n18749), .B(n18741), .Z(n18767) );
  XOR U18741 ( .A(n18773), .B(n18774), .Z(n18741) );
  AND U18742 ( .A(n18775), .B(n18776), .Z(n18774) );
  XOR U18743 ( .A(n18773), .B(n18777), .Z(n18775) );
  XNOR U18744 ( .A(n18778), .B(n18746), .Z(n18749) );
  XOR U18745 ( .A(n18779), .B(n18780), .Z(n18746) );
  AND U18746 ( .A(n18781), .B(n18782), .Z(n18780) );
  XNOR U18747 ( .A(n18783), .B(n18784), .Z(n18781) );
  IV U18748 ( .A(n18779), .Z(n18783) );
  XNOR U18749 ( .A(n18785), .B(n18786), .Z(n18778) );
  NOR U18750 ( .A(n18787), .B(n18788), .Z(n18786) );
  XNOR U18751 ( .A(n18785), .B(n18789), .Z(n18787) );
  XNOR U18752 ( .A(n18745), .B(n18752), .Z(n18766) );
  NOR U18753 ( .A(n18709), .B(n18790), .Z(n18752) );
  XOR U18754 ( .A(n18757), .B(n18756), .Z(n18745) );
  XNOR U18755 ( .A(n18791), .B(n18753), .Z(n18756) );
  XOR U18756 ( .A(n18792), .B(n18793), .Z(n18753) );
  AND U18757 ( .A(n18794), .B(n18795), .Z(n18793) );
  XNOR U18758 ( .A(n18796), .B(n18797), .Z(n18794) );
  IV U18759 ( .A(n18792), .Z(n18796) );
  XNOR U18760 ( .A(n18798), .B(n18799), .Z(n18791) );
  NOR U18761 ( .A(n18800), .B(n18801), .Z(n18799) );
  XNOR U18762 ( .A(n18798), .B(n18802), .Z(n18800) );
  XOR U18763 ( .A(n18803), .B(n18804), .Z(n18757) );
  NOR U18764 ( .A(n18805), .B(n18806), .Z(n18804) );
  XNOR U18765 ( .A(n18803), .B(n18807), .Z(n18805) );
  XNOR U18766 ( .A(n18693), .B(n18762), .Z(n18764) );
  XOR U18767 ( .A(n18808), .B(n18809), .Z(n18693) );
  AND U18768 ( .A(n447), .B(n18810), .Z(n18809) );
  XOR U18769 ( .A(n18811), .B(n18808), .Z(n18810) );
  AND U18770 ( .A(n18706), .B(n18709), .Z(n18762) );
  XOR U18771 ( .A(n18812), .B(n18790), .Z(n18709) );
  XNOR U18772 ( .A(p_input[1760]), .B(p_input[2048]), .Z(n18790) );
  XNOR U18773 ( .A(n18777), .B(n18776), .Z(n18812) );
  XNOR U18774 ( .A(n18813), .B(n18784), .Z(n18776) );
  XNOR U18775 ( .A(n18772), .B(n18771), .Z(n18784) );
  XNOR U18776 ( .A(n18814), .B(n18768), .Z(n18771) );
  XNOR U18777 ( .A(p_input[1770]), .B(p_input[2058]), .Z(n18768) );
  XOR U18778 ( .A(p_input[1771]), .B(n6319), .Z(n18814) );
  XOR U18779 ( .A(p_input[1772]), .B(p_input[2060]), .Z(n18772) );
  XOR U18780 ( .A(n18782), .B(n18815), .Z(n18813) );
  IV U18781 ( .A(n18773), .Z(n18815) );
  XOR U18782 ( .A(p_input[1761]), .B(p_input[2049]), .Z(n18773) );
  XNOR U18783 ( .A(n18816), .B(n18789), .Z(n18782) );
  XNOR U18784 ( .A(p_input[1775]), .B(n6322), .Z(n18789) );
  XOR U18785 ( .A(n18779), .B(n18788), .Z(n18816) );
  XOR U18786 ( .A(n18817), .B(n18785), .Z(n18788) );
  XOR U18787 ( .A(p_input[1773]), .B(p_input[2061]), .Z(n18785) );
  XOR U18788 ( .A(p_input[1774]), .B(n6324), .Z(n18817) );
  XOR U18789 ( .A(p_input[1769]), .B(p_input[2057]), .Z(n18779) );
  XOR U18790 ( .A(n18797), .B(n18795), .Z(n18777) );
  XNOR U18791 ( .A(n18818), .B(n18802), .Z(n18795) );
  XOR U18792 ( .A(p_input[1768]), .B(p_input[2056]), .Z(n18802) );
  XOR U18793 ( .A(n18792), .B(n18801), .Z(n18818) );
  XOR U18794 ( .A(n18819), .B(n18798), .Z(n18801) );
  XOR U18795 ( .A(p_input[1766]), .B(p_input[2054]), .Z(n18798) );
  XOR U18796 ( .A(p_input[1767]), .B(n7007), .Z(n18819) );
  XOR U18797 ( .A(p_input[1762]), .B(p_input[2050]), .Z(n18792) );
  XNOR U18798 ( .A(n18807), .B(n18806), .Z(n18797) );
  XOR U18799 ( .A(n18820), .B(n18803), .Z(n18806) );
  XOR U18800 ( .A(p_input[1763]), .B(p_input[2051]), .Z(n18803) );
  XOR U18801 ( .A(p_input[1764]), .B(n7009), .Z(n18820) );
  XOR U18802 ( .A(p_input[1765]), .B(p_input[2053]), .Z(n18807) );
  XOR U18803 ( .A(n18821), .B(n18822), .Z(n18706) );
  AND U18804 ( .A(n447), .B(n18823), .Z(n18822) );
  XNOR U18805 ( .A(n18824), .B(n18821), .Z(n18823) );
  XNOR U18806 ( .A(n18825), .B(n18826), .Z(n447) );
  AND U18807 ( .A(n18827), .B(n18828), .Z(n18826) );
  XOR U18808 ( .A(n18719), .B(n18825), .Z(n18828) );
  AND U18809 ( .A(n18829), .B(n18830), .Z(n18719) );
  XNOR U18810 ( .A(n18716), .B(n18825), .Z(n18827) );
  XOR U18811 ( .A(n18831), .B(n18832), .Z(n18716) );
  AND U18812 ( .A(n451), .B(n18833), .Z(n18832) );
  XOR U18813 ( .A(n18834), .B(n18831), .Z(n18833) );
  XOR U18814 ( .A(n18835), .B(n18836), .Z(n18825) );
  AND U18815 ( .A(n18837), .B(n18838), .Z(n18836) );
  XNOR U18816 ( .A(n18835), .B(n18829), .Z(n18838) );
  IV U18817 ( .A(n18734), .Z(n18829) );
  XOR U18818 ( .A(n18839), .B(n18840), .Z(n18734) );
  XOR U18819 ( .A(n18841), .B(n18830), .Z(n18840) );
  AND U18820 ( .A(n18761), .B(n18842), .Z(n18830) );
  AND U18821 ( .A(n18843), .B(n18844), .Z(n18841) );
  XOR U18822 ( .A(n18845), .B(n18839), .Z(n18843) );
  XNOR U18823 ( .A(n18731), .B(n18835), .Z(n18837) );
  XOR U18824 ( .A(n18846), .B(n18847), .Z(n18731) );
  AND U18825 ( .A(n451), .B(n18848), .Z(n18847) );
  XOR U18826 ( .A(n18849), .B(n18846), .Z(n18848) );
  XOR U18827 ( .A(n18850), .B(n18851), .Z(n18835) );
  AND U18828 ( .A(n18852), .B(n18853), .Z(n18851) );
  XNOR U18829 ( .A(n18850), .B(n18761), .Z(n18853) );
  XOR U18830 ( .A(n18854), .B(n18844), .Z(n18761) );
  XNOR U18831 ( .A(n18855), .B(n18839), .Z(n18844) );
  XOR U18832 ( .A(n18856), .B(n18857), .Z(n18839) );
  AND U18833 ( .A(n18858), .B(n18859), .Z(n18857) );
  XOR U18834 ( .A(n18860), .B(n18856), .Z(n18858) );
  XNOR U18835 ( .A(n18861), .B(n18862), .Z(n18855) );
  AND U18836 ( .A(n18863), .B(n18864), .Z(n18862) );
  XOR U18837 ( .A(n18861), .B(n18865), .Z(n18863) );
  XNOR U18838 ( .A(n18845), .B(n18842), .Z(n18854) );
  AND U18839 ( .A(n18866), .B(n18867), .Z(n18842) );
  XOR U18840 ( .A(n18868), .B(n18869), .Z(n18845) );
  AND U18841 ( .A(n18870), .B(n18871), .Z(n18869) );
  XOR U18842 ( .A(n18868), .B(n18872), .Z(n18870) );
  XNOR U18843 ( .A(n18758), .B(n18850), .Z(n18852) );
  XOR U18844 ( .A(n18873), .B(n18874), .Z(n18758) );
  AND U18845 ( .A(n451), .B(n18875), .Z(n18874) );
  XNOR U18846 ( .A(n18876), .B(n18873), .Z(n18875) );
  XOR U18847 ( .A(n18877), .B(n18878), .Z(n18850) );
  AND U18848 ( .A(n18879), .B(n18880), .Z(n18878) );
  XNOR U18849 ( .A(n18877), .B(n18866), .Z(n18880) );
  IV U18850 ( .A(n18811), .Z(n18866) );
  XNOR U18851 ( .A(n18881), .B(n18859), .Z(n18811) );
  XNOR U18852 ( .A(n18882), .B(n18865), .Z(n18859) );
  XNOR U18853 ( .A(n18883), .B(n18884), .Z(n18865) );
  NOR U18854 ( .A(n18885), .B(n18886), .Z(n18884) );
  XOR U18855 ( .A(n18883), .B(n18887), .Z(n18885) );
  XNOR U18856 ( .A(n18864), .B(n18856), .Z(n18882) );
  XOR U18857 ( .A(n18888), .B(n18889), .Z(n18856) );
  AND U18858 ( .A(n18890), .B(n18891), .Z(n18889) );
  XOR U18859 ( .A(n18888), .B(n18892), .Z(n18890) );
  XNOR U18860 ( .A(n18893), .B(n18861), .Z(n18864) );
  XOR U18861 ( .A(n18894), .B(n18895), .Z(n18861) );
  AND U18862 ( .A(n18896), .B(n18897), .Z(n18895) );
  XNOR U18863 ( .A(n18898), .B(n18899), .Z(n18896) );
  IV U18864 ( .A(n18894), .Z(n18898) );
  XNOR U18865 ( .A(n18900), .B(n18901), .Z(n18893) );
  NOR U18866 ( .A(n18902), .B(n18903), .Z(n18901) );
  XNOR U18867 ( .A(n18900), .B(n18904), .Z(n18902) );
  XNOR U18868 ( .A(n18860), .B(n18867), .Z(n18881) );
  NOR U18869 ( .A(n18824), .B(n18905), .Z(n18867) );
  XOR U18870 ( .A(n18872), .B(n18871), .Z(n18860) );
  XNOR U18871 ( .A(n18906), .B(n18868), .Z(n18871) );
  XOR U18872 ( .A(n18907), .B(n18908), .Z(n18868) );
  AND U18873 ( .A(n18909), .B(n18910), .Z(n18908) );
  XNOR U18874 ( .A(n18911), .B(n18912), .Z(n18909) );
  IV U18875 ( .A(n18907), .Z(n18911) );
  XNOR U18876 ( .A(n18913), .B(n18914), .Z(n18906) );
  NOR U18877 ( .A(n18915), .B(n18916), .Z(n18914) );
  XNOR U18878 ( .A(n18913), .B(n18917), .Z(n18915) );
  XOR U18879 ( .A(n18918), .B(n18919), .Z(n18872) );
  NOR U18880 ( .A(n18920), .B(n18921), .Z(n18919) );
  XNOR U18881 ( .A(n18918), .B(n18922), .Z(n18920) );
  XNOR U18882 ( .A(n18808), .B(n18877), .Z(n18879) );
  XOR U18883 ( .A(n18923), .B(n18924), .Z(n18808) );
  AND U18884 ( .A(n451), .B(n18925), .Z(n18924) );
  XOR U18885 ( .A(n18926), .B(n18923), .Z(n18925) );
  AND U18886 ( .A(n18821), .B(n18824), .Z(n18877) );
  XOR U18887 ( .A(n18927), .B(n18905), .Z(n18824) );
  XNOR U18888 ( .A(p_input[1776]), .B(p_input[2048]), .Z(n18905) );
  XNOR U18889 ( .A(n18892), .B(n18891), .Z(n18927) );
  XNOR U18890 ( .A(n18928), .B(n18899), .Z(n18891) );
  XNOR U18891 ( .A(n18887), .B(n18886), .Z(n18899) );
  XNOR U18892 ( .A(n18929), .B(n18883), .Z(n18886) );
  XNOR U18893 ( .A(p_input[1786]), .B(p_input[2058]), .Z(n18883) );
  XOR U18894 ( .A(p_input[1787]), .B(n6319), .Z(n18929) );
  XOR U18895 ( .A(p_input[1788]), .B(p_input[2060]), .Z(n18887) );
  XOR U18896 ( .A(n18897), .B(n18930), .Z(n18928) );
  IV U18897 ( .A(n18888), .Z(n18930) );
  XOR U18898 ( .A(p_input[1777]), .B(p_input[2049]), .Z(n18888) );
  XNOR U18899 ( .A(n18931), .B(n18904), .Z(n18897) );
  XNOR U18900 ( .A(p_input[1791]), .B(n6322), .Z(n18904) );
  XOR U18901 ( .A(n18894), .B(n18903), .Z(n18931) );
  XOR U18902 ( .A(n18932), .B(n18900), .Z(n18903) );
  XOR U18903 ( .A(p_input[1789]), .B(p_input[2061]), .Z(n18900) );
  XOR U18904 ( .A(p_input[1790]), .B(n6324), .Z(n18932) );
  XOR U18905 ( .A(p_input[1785]), .B(p_input[2057]), .Z(n18894) );
  XOR U18906 ( .A(n18912), .B(n18910), .Z(n18892) );
  XNOR U18907 ( .A(n18933), .B(n18917), .Z(n18910) );
  XOR U18908 ( .A(p_input[1784]), .B(p_input[2056]), .Z(n18917) );
  XOR U18909 ( .A(n18907), .B(n18916), .Z(n18933) );
  XOR U18910 ( .A(n18934), .B(n18913), .Z(n18916) );
  XOR U18911 ( .A(p_input[1782]), .B(p_input[2054]), .Z(n18913) );
  XOR U18912 ( .A(p_input[1783]), .B(n7007), .Z(n18934) );
  XOR U18913 ( .A(p_input[1778]), .B(p_input[2050]), .Z(n18907) );
  XNOR U18914 ( .A(n18922), .B(n18921), .Z(n18912) );
  XOR U18915 ( .A(n18935), .B(n18918), .Z(n18921) );
  XOR U18916 ( .A(p_input[1779]), .B(p_input[2051]), .Z(n18918) );
  XOR U18917 ( .A(p_input[1780]), .B(n7009), .Z(n18935) );
  XOR U18918 ( .A(p_input[1781]), .B(p_input[2053]), .Z(n18922) );
  XOR U18919 ( .A(n18936), .B(n18937), .Z(n18821) );
  AND U18920 ( .A(n451), .B(n18938), .Z(n18937) );
  XNOR U18921 ( .A(n18939), .B(n18936), .Z(n18938) );
  XNOR U18922 ( .A(n18940), .B(n18941), .Z(n451) );
  AND U18923 ( .A(n18942), .B(n18943), .Z(n18941) );
  XOR U18924 ( .A(n18834), .B(n18940), .Z(n18943) );
  AND U18925 ( .A(n18944), .B(n18945), .Z(n18834) );
  XNOR U18926 ( .A(n18831), .B(n18940), .Z(n18942) );
  XOR U18927 ( .A(n18946), .B(n18947), .Z(n18831) );
  AND U18928 ( .A(n455), .B(n18948), .Z(n18947) );
  XOR U18929 ( .A(n18949), .B(n18946), .Z(n18948) );
  XOR U18930 ( .A(n18950), .B(n18951), .Z(n18940) );
  AND U18931 ( .A(n18952), .B(n18953), .Z(n18951) );
  XNOR U18932 ( .A(n18950), .B(n18944), .Z(n18953) );
  IV U18933 ( .A(n18849), .Z(n18944) );
  XOR U18934 ( .A(n18954), .B(n18955), .Z(n18849) );
  XOR U18935 ( .A(n18956), .B(n18945), .Z(n18955) );
  AND U18936 ( .A(n18876), .B(n18957), .Z(n18945) );
  AND U18937 ( .A(n18958), .B(n18959), .Z(n18956) );
  XOR U18938 ( .A(n18960), .B(n18954), .Z(n18958) );
  XNOR U18939 ( .A(n18846), .B(n18950), .Z(n18952) );
  XOR U18940 ( .A(n18961), .B(n18962), .Z(n18846) );
  AND U18941 ( .A(n455), .B(n18963), .Z(n18962) );
  XOR U18942 ( .A(n18964), .B(n18961), .Z(n18963) );
  XOR U18943 ( .A(n18965), .B(n18966), .Z(n18950) );
  AND U18944 ( .A(n18967), .B(n18968), .Z(n18966) );
  XNOR U18945 ( .A(n18965), .B(n18876), .Z(n18968) );
  XOR U18946 ( .A(n18969), .B(n18959), .Z(n18876) );
  XNOR U18947 ( .A(n18970), .B(n18954), .Z(n18959) );
  XOR U18948 ( .A(n18971), .B(n18972), .Z(n18954) );
  AND U18949 ( .A(n18973), .B(n18974), .Z(n18972) );
  XOR U18950 ( .A(n18975), .B(n18971), .Z(n18973) );
  XNOR U18951 ( .A(n18976), .B(n18977), .Z(n18970) );
  AND U18952 ( .A(n18978), .B(n18979), .Z(n18977) );
  XOR U18953 ( .A(n18976), .B(n18980), .Z(n18978) );
  XNOR U18954 ( .A(n18960), .B(n18957), .Z(n18969) );
  AND U18955 ( .A(n18981), .B(n18982), .Z(n18957) );
  XOR U18956 ( .A(n18983), .B(n18984), .Z(n18960) );
  AND U18957 ( .A(n18985), .B(n18986), .Z(n18984) );
  XOR U18958 ( .A(n18983), .B(n18987), .Z(n18985) );
  XNOR U18959 ( .A(n18873), .B(n18965), .Z(n18967) );
  XOR U18960 ( .A(n18988), .B(n18989), .Z(n18873) );
  AND U18961 ( .A(n455), .B(n18990), .Z(n18989) );
  XNOR U18962 ( .A(n18991), .B(n18988), .Z(n18990) );
  XOR U18963 ( .A(n18992), .B(n18993), .Z(n18965) );
  AND U18964 ( .A(n18994), .B(n18995), .Z(n18993) );
  XNOR U18965 ( .A(n18992), .B(n18981), .Z(n18995) );
  IV U18966 ( .A(n18926), .Z(n18981) );
  XNOR U18967 ( .A(n18996), .B(n18974), .Z(n18926) );
  XNOR U18968 ( .A(n18997), .B(n18980), .Z(n18974) );
  XNOR U18969 ( .A(n18998), .B(n18999), .Z(n18980) );
  NOR U18970 ( .A(n19000), .B(n19001), .Z(n18999) );
  XOR U18971 ( .A(n18998), .B(n19002), .Z(n19000) );
  XNOR U18972 ( .A(n18979), .B(n18971), .Z(n18997) );
  XOR U18973 ( .A(n19003), .B(n19004), .Z(n18971) );
  AND U18974 ( .A(n19005), .B(n19006), .Z(n19004) );
  XOR U18975 ( .A(n19003), .B(n19007), .Z(n19005) );
  XNOR U18976 ( .A(n19008), .B(n18976), .Z(n18979) );
  XOR U18977 ( .A(n19009), .B(n19010), .Z(n18976) );
  AND U18978 ( .A(n19011), .B(n19012), .Z(n19010) );
  XNOR U18979 ( .A(n19013), .B(n19014), .Z(n19011) );
  IV U18980 ( .A(n19009), .Z(n19013) );
  XNOR U18981 ( .A(n19015), .B(n19016), .Z(n19008) );
  NOR U18982 ( .A(n19017), .B(n19018), .Z(n19016) );
  XNOR U18983 ( .A(n19015), .B(n19019), .Z(n19017) );
  XNOR U18984 ( .A(n18975), .B(n18982), .Z(n18996) );
  NOR U18985 ( .A(n18939), .B(n19020), .Z(n18982) );
  XOR U18986 ( .A(n18987), .B(n18986), .Z(n18975) );
  XNOR U18987 ( .A(n19021), .B(n18983), .Z(n18986) );
  XOR U18988 ( .A(n19022), .B(n19023), .Z(n18983) );
  AND U18989 ( .A(n19024), .B(n19025), .Z(n19023) );
  XNOR U18990 ( .A(n19026), .B(n19027), .Z(n19024) );
  IV U18991 ( .A(n19022), .Z(n19026) );
  XNOR U18992 ( .A(n19028), .B(n19029), .Z(n19021) );
  NOR U18993 ( .A(n19030), .B(n19031), .Z(n19029) );
  XNOR U18994 ( .A(n19028), .B(n19032), .Z(n19030) );
  XOR U18995 ( .A(n19033), .B(n19034), .Z(n18987) );
  NOR U18996 ( .A(n19035), .B(n19036), .Z(n19034) );
  XNOR U18997 ( .A(n19033), .B(n19037), .Z(n19035) );
  XNOR U18998 ( .A(n18923), .B(n18992), .Z(n18994) );
  XOR U18999 ( .A(n19038), .B(n19039), .Z(n18923) );
  AND U19000 ( .A(n455), .B(n19040), .Z(n19039) );
  XOR U19001 ( .A(n19041), .B(n19038), .Z(n19040) );
  AND U19002 ( .A(n18936), .B(n18939), .Z(n18992) );
  XOR U19003 ( .A(n19042), .B(n19020), .Z(n18939) );
  XNOR U19004 ( .A(p_input[1792]), .B(p_input[2048]), .Z(n19020) );
  XNOR U19005 ( .A(n19007), .B(n19006), .Z(n19042) );
  XNOR U19006 ( .A(n19043), .B(n19014), .Z(n19006) );
  XNOR U19007 ( .A(n19002), .B(n19001), .Z(n19014) );
  XNOR U19008 ( .A(n19044), .B(n18998), .Z(n19001) );
  XNOR U19009 ( .A(p_input[1802]), .B(p_input[2058]), .Z(n18998) );
  XOR U19010 ( .A(p_input[1803]), .B(n6319), .Z(n19044) );
  XOR U19011 ( .A(p_input[1804]), .B(p_input[2060]), .Z(n19002) );
  XOR U19012 ( .A(n19012), .B(n19045), .Z(n19043) );
  IV U19013 ( .A(n19003), .Z(n19045) );
  XOR U19014 ( .A(p_input[1793]), .B(p_input[2049]), .Z(n19003) );
  XNOR U19015 ( .A(n19046), .B(n19019), .Z(n19012) );
  XNOR U19016 ( .A(p_input[1807]), .B(n6322), .Z(n19019) );
  XOR U19017 ( .A(n19009), .B(n19018), .Z(n19046) );
  XOR U19018 ( .A(n19047), .B(n19015), .Z(n19018) );
  XOR U19019 ( .A(p_input[1805]), .B(p_input[2061]), .Z(n19015) );
  XOR U19020 ( .A(p_input[1806]), .B(n6324), .Z(n19047) );
  XOR U19021 ( .A(p_input[1801]), .B(p_input[2057]), .Z(n19009) );
  XOR U19022 ( .A(n19027), .B(n19025), .Z(n19007) );
  XNOR U19023 ( .A(n19048), .B(n19032), .Z(n19025) );
  XOR U19024 ( .A(p_input[1800]), .B(p_input[2056]), .Z(n19032) );
  XOR U19025 ( .A(n19022), .B(n19031), .Z(n19048) );
  XOR U19026 ( .A(n19049), .B(n19028), .Z(n19031) );
  XOR U19027 ( .A(p_input[1798]), .B(p_input[2054]), .Z(n19028) );
  XOR U19028 ( .A(p_input[1799]), .B(n7007), .Z(n19049) );
  XOR U19029 ( .A(p_input[1794]), .B(p_input[2050]), .Z(n19022) );
  XNOR U19030 ( .A(n19037), .B(n19036), .Z(n19027) );
  XOR U19031 ( .A(n19050), .B(n19033), .Z(n19036) );
  XOR U19032 ( .A(p_input[1795]), .B(p_input[2051]), .Z(n19033) );
  XOR U19033 ( .A(p_input[1796]), .B(n7009), .Z(n19050) );
  XOR U19034 ( .A(p_input[1797]), .B(p_input[2053]), .Z(n19037) );
  XOR U19035 ( .A(n19051), .B(n19052), .Z(n18936) );
  AND U19036 ( .A(n455), .B(n19053), .Z(n19052) );
  XNOR U19037 ( .A(n19054), .B(n19051), .Z(n19053) );
  XNOR U19038 ( .A(n19055), .B(n19056), .Z(n455) );
  AND U19039 ( .A(n19057), .B(n19058), .Z(n19056) );
  XOR U19040 ( .A(n18949), .B(n19055), .Z(n19058) );
  AND U19041 ( .A(n19059), .B(n19060), .Z(n18949) );
  XNOR U19042 ( .A(n18946), .B(n19055), .Z(n19057) );
  XOR U19043 ( .A(n19061), .B(n19062), .Z(n18946) );
  AND U19044 ( .A(n459), .B(n19063), .Z(n19062) );
  XOR U19045 ( .A(n19064), .B(n19061), .Z(n19063) );
  XOR U19046 ( .A(n19065), .B(n19066), .Z(n19055) );
  AND U19047 ( .A(n19067), .B(n19068), .Z(n19066) );
  XNOR U19048 ( .A(n19065), .B(n19059), .Z(n19068) );
  IV U19049 ( .A(n18964), .Z(n19059) );
  XOR U19050 ( .A(n19069), .B(n19070), .Z(n18964) );
  XOR U19051 ( .A(n19071), .B(n19060), .Z(n19070) );
  AND U19052 ( .A(n18991), .B(n19072), .Z(n19060) );
  AND U19053 ( .A(n19073), .B(n19074), .Z(n19071) );
  XOR U19054 ( .A(n19075), .B(n19069), .Z(n19073) );
  XNOR U19055 ( .A(n18961), .B(n19065), .Z(n19067) );
  XOR U19056 ( .A(n19076), .B(n19077), .Z(n18961) );
  AND U19057 ( .A(n459), .B(n19078), .Z(n19077) );
  XOR U19058 ( .A(n19079), .B(n19076), .Z(n19078) );
  XOR U19059 ( .A(n19080), .B(n19081), .Z(n19065) );
  AND U19060 ( .A(n19082), .B(n19083), .Z(n19081) );
  XNOR U19061 ( .A(n19080), .B(n18991), .Z(n19083) );
  XOR U19062 ( .A(n19084), .B(n19074), .Z(n18991) );
  XNOR U19063 ( .A(n19085), .B(n19069), .Z(n19074) );
  XOR U19064 ( .A(n19086), .B(n19087), .Z(n19069) );
  AND U19065 ( .A(n19088), .B(n19089), .Z(n19087) );
  XOR U19066 ( .A(n19090), .B(n19086), .Z(n19088) );
  XNOR U19067 ( .A(n19091), .B(n19092), .Z(n19085) );
  AND U19068 ( .A(n19093), .B(n19094), .Z(n19092) );
  XOR U19069 ( .A(n19091), .B(n19095), .Z(n19093) );
  XNOR U19070 ( .A(n19075), .B(n19072), .Z(n19084) );
  AND U19071 ( .A(n19096), .B(n19097), .Z(n19072) );
  XOR U19072 ( .A(n19098), .B(n19099), .Z(n19075) );
  AND U19073 ( .A(n19100), .B(n19101), .Z(n19099) );
  XOR U19074 ( .A(n19098), .B(n19102), .Z(n19100) );
  XNOR U19075 ( .A(n18988), .B(n19080), .Z(n19082) );
  XOR U19076 ( .A(n19103), .B(n19104), .Z(n18988) );
  AND U19077 ( .A(n459), .B(n19105), .Z(n19104) );
  XNOR U19078 ( .A(n19106), .B(n19103), .Z(n19105) );
  XOR U19079 ( .A(n19107), .B(n19108), .Z(n19080) );
  AND U19080 ( .A(n19109), .B(n19110), .Z(n19108) );
  XNOR U19081 ( .A(n19107), .B(n19096), .Z(n19110) );
  IV U19082 ( .A(n19041), .Z(n19096) );
  XNOR U19083 ( .A(n19111), .B(n19089), .Z(n19041) );
  XNOR U19084 ( .A(n19112), .B(n19095), .Z(n19089) );
  XNOR U19085 ( .A(n19113), .B(n19114), .Z(n19095) );
  NOR U19086 ( .A(n19115), .B(n19116), .Z(n19114) );
  XOR U19087 ( .A(n19113), .B(n19117), .Z(n19115) );
  XNOR U19088 ( .A(n19094), .B(n19086), .Z(n19112) );
  XOR U19089 ( .A(n19118), .B(n19119), .Z(n19086) );
  AND U19090 ( .A(n19120), .B(n19121), .Z(n19119) );
  XOR U19091 ( .A(n19118), .B(n19122), .Z(n19120) );
  XNOR U19092 ( .A(n19123), .B(n19091), .Z(n19094) );
  XOR U19093 ( .A(n19124), .B(n19125), .Z(n19091) );
  AND U19094 ( .A(n19126), .B(n19127), .Z(n19125) );
  XNOR U19095 ( .A(n19128), .B(n19129), .Z(n19126) );
  IV U19096 ( .A(n19124), .Z(n19128) );
  XNOR U19097 ( .A(n19130), .B(n19131), .Z(n19123) );
  NOR U19098 ( .A(n19132), .B(n19133), .Z(n19131) );
  XNOR U19099 ( .A(n19130), .B(n19134), .Z(n19132) );
  XNOR U19100 ( .A(n19090), .B(n19097), .Z(n19111) );
  NOR U19101 ( .A(n19054), .B(n19135), .Z(n19097) );
  XOR U19102 ( .A(n19102), .B(n19101), .Z(n19090) );
  XNOR U19103 ( .A(n19136), .B(n19098), .Z(n19101) );
  XOR U19104 ( .A(n19137), .B(n19138), .Z(n19098) );
  AND U19105 ( .A(n19139), .B(n19140), .Z(n19138) );
  XNOR U19106 ( .A(n19141), .B(n19142), .Z(n19139) );
  IV U19107 ( .A(n19137), .Z(n19141) );
  XNOR U19108 ( .A(n19143), .B(n19144), .Z(n19136) );
  NOR U19109 ( .A(n19145), .B(n19146), .Z(n19144) );
  XNOR U19110 ( .A(n19143), .B(n19147), .Z(n19145) );
  XOR U19111 ( .A(n19148), .B(n19149), .Z(n19102) );
  NOR U19112 ( .A(n19150), .B(n19151), .Z(n19149) );
  XNOR U19113 ( .A(n19148), .B(n19152), .Z(n19150) );
  XNOR U19114 ( .A(n19038), .B(n19107), .Z(n19109) );
  XOR U19115 ( .A(n19153), .B(n19154), .Z(n19038) );
  AND U19116 ( .A(n459), .B(n19155), .Z(n19154) );
  XOR U19117 ( .A(n19156), .B(n19153), .Z(n19155) );
  AND U19118 ( .A(n19051), .B(n19054), .Z(n19107) );
  XOR U19119 ( .A(n19157), .B(n19135), .Z(n19054) );
  XNOR U19120 ( .A(p_input[1808]), .B(p_input[2048]), .Z(n19135) );
  XNOR U19121 ( .A(n19122), .B(n19121), .Z(n19157) );
  XNOR U19122 ( .A(n19158), .B(n19129), .Z(n19121) );
  XNOR U19123 ( .A(n19117), .B(n19116), .Z(n19129) );
  XNOR U19124 ( .A(n19159), .B(n19113), .Z(n19116) );
  XNOR U19125 ( .A(p_input[1818]), .B(p_input[2058]), .Z(n19113) );
  XOR U19126 ( .A(p_input[1819]), .B(n6319), .Z(n19159) );
  XOR U19127 ( .A(p_input[1820]), .B(p_input[2060]), .Z(n19117) );
  XOR U19128 ( .A(n19127), .B(n19160), .Z(n19158) );
  IV U19129 ( .A(n19118), .Z(n19160) );
  XOR U19130 ( .A(p_input[1809]), .B(p_input[2049]), .Z(n19118) );
  XNOR U19131 ( .A(n19161), .B(n19134), .Z(n19127) );
  XNOR U19132 ( .A(p_input[1823]), .B(n6322), .Z(n19134) );
  XOR U19133 ( .A(n19124), .B(n19133), .Z(n19161) );
  XOR U19134 ( .A(n19162), .B(n19130), .Z(n19133) );
  XOR U19135 ( .A(p_input[1821]), .B(p_input[2061]), .Z(n19130) );
  XOR U19136 ( .A(p_input[1822]), .B(n6324), .Z(n19162) );
  XOR U19137 ( .A(p_input[1817]), .B(p_input[2057]), .Z(n19124) );
  XOR U19138 ( .A(n19142), .B(n19140), .Z(n19122) );
  XNOR U19139 ( .A(n19163), .B(n19147), .Z(n19140) );
  XOR U19140 ( .A(p_input[1816]), .B(p_input[2056]), .Z(n19147) );
  XOR U19141 ( .A(n19137), .B(n19146), .Z(n19163) );
  XOR U19142 ( .A(n19164), .B(n19143), .Z(n19146) );
  XOR U19143 ( .A(p_input[1814]), .B(p_input[2054]), .Z(n19143) );
  XOR U19144 ( .A(p_input[1815]), .B(n7007), .Z(n19164) );
  XOR U19145 ( .A(p_input[1810]), .B(p_input[2050]), .Z(n19137) );
  XNOR U19146 ( .A(n19152), .B(n19151), .Z(n19142) );
  XOR U19147 ( .A(n19165), .B(n19148), .Z(n19151) );
  XOR U19148 ( .A(p_input[1811]), .B(p_input[2051]), .Z(n19148) );
  XOR U19149 ( .A(p_input[1812]), .B(n7009), .Z(n19165) );
  XOR U19150 ( .A(p_input[1813]), .B(p_input[2053]), .Z(n19152) );
  XOR U19151 ( .A(n19166), .B(n19167), .Z(n19051) );
  AND U19152 ( .A(n459), .B(n19168), .Z(n19167) );
  XNOR U19153 ( .A(n19169), .B(n19166), .Z(n19168) );
  XNOR U19154 ( .A(n19170), .B(n19171), .Z(n459) );
  AND U19155 ( .A(n19172), .B(n19173), .Z(n19171) );
  XOR U19156 ( .A(n19064), .B(n19170), .Z(n19173) );
  AND U19157 ( .A(n19174), .B(n19175), .Z(n19064) );
  XNOR U19158 ( .A(n19061), .B(n19170), .Z(n19172) );
  XOR U19159 ( .A(n19176), .B(n19177), .Z(n19061) );
  AND U19160 ( .A(n463), .B(n19178), .Z(n19177) );
  XOR U19161 ( .A(n19179), .B(n19176), .Z(n19178) );
  XOR U19162 ( .A(n19180), .B(n19181), .Z(n19170) );
  AND U19163 ( .A(n19182), .B(n19183), .Z(n19181) );
  XNOR U19164 ( .A(n19180), .B(n19174), .Z(n19183) );
  IV U19165 ( .A(n19079), .Z(n19174) );
  XOR U19166 ( .A(n19184), .B(n19185), .Z(n19079) );
  XOR U19167 ( .A(n19186), .B(n19175), .Z(n19185) );
  AND U19168 ( .A(n19106), .B(n19187), .Z(n19175) );
  AND U19169 ( .A(n19188), .B(n19189), .Z(n19186) );
  XOR U19170 ( .A(n19190), .B(n19184), .Z(n19188) );
  XNOR U19171 ( .A(n19076), .B(n19180), .Z(n19182) );
  XOR U19172 ( .A(n19191), .B(n19192), .Z(n19076) );
  AND U19173 ( .A(n463), .B(n19193), .Z(n19192) );
  XOR U19174 ( .A(n19194), .B(n19191), .Z(n19193) );
  XOR U19175 ( .A(n19195), .B(n19196), .Z(n19180) );
  AND U19176 ( .A(n19197), .B(n19198), .Z(n19196) );
  XNOR U19177 ( .A(n19195), .B(n19106), .Z(n19198) );
  XOR U19178 ( .A(n19199), .B(n19189), .Z(n19106) );
  XNOR U19179 ( .A(n19200), .B(n19184), .Z(n19189) );
  XOR U19180 ( .A(n19201), .B(n19202), .Z(n19184) );
  AND U19181 ( .A(n19203), .B(n19204), .Z(n19202) );
  XOR U19182 ( .A(n19205), .B(n19201), .Z(n19203) );
  XNOR U19183 ( .A(n19206), .B(n19207), .Z(n19200) );
  AND U19184 ( .A(n19208), .B(n19209), .Z(n19207) );
  XOR U19185 ( .A(n19206), .B(n19210), .Z(n19208) );
  XNOR U19186 ( .A(n19190), .B(n19187), .Z(n19199) );
  AND U19187 ( .A(n19211), .B(n19212), .Z(n19187) );
  XOR U19188 ( .A(n19213), .B(n19214), .Z(n19190) );
  AND U19189 ( .A(n19215), .B(n19216), .Z(n19214) );
  XOR U19190 ( .A(n19213), .B(n19217), .Z(n19215) );
  XNOR U19191 ( .A(n19103), .B(n19195), .Z(n19197) );
  XOR U19192 ( .A(n19218), .B(n19219), .Z(n19103) );
  AND U19193 ( .A(n463), .B(n19220), .Z(n19219) );
  XNOR U19194 ( .A(n19221), .B(n19218), .Z(n19220) );
  XOR U19195 ( .A(n19222), .B(n19223), .Z(n19195) );
  AND U19196 ( .A(n19224), .B(n19225), .Z(n19223) );
  XNOR U19197 ( .A(n19222), .B(n19211), .Z(n19225) );
  IV U19198 ( .A(n19156), .Z(n19211) );
  XNOR U19199 ( .A(n19226), .B(n19204), .Z(n19156) );
  XNOR U19200 ( .A(n19227), .B(n19210), .Z(n19204) );
  XNOR U19201 ( .A(n19228), .B(n19229), .Z(n19210) );
  NOR U19202 ( .A(n19230), .B(n19231), .Z(n19229) );
  XOR U19203 ( .A(n19228), .B(n19232), .Z(n19230) );
  XNOR U19204 ( .A(n19209), .B(n19201), .Z(n19227) );
  XOR U19205 ( .A(n19233), .B(n19234), .Z(n19201) );
  AND U19206 ( .A(n19235), .B(n19236), .Z(n19234) );
  XOR U19207 ( .A(n19233), .B(n19237), .Z(n19235) );
  XNOR U19208 ( .A(n19238), .B(n19206), .Z(n19209) );
  XOR U19209 ( .A(n19239), .B(n19240), .Z(n19206) );
  AND U19210 ( .A(n19241), .B(n19242), .Z(n19240) );
  XNOR U19211 ( .A(n19243), .B(n19244), .Z(n19241) );
  IV U19212 ( .A(n19239), .Z(n19243) );
  XNOR U19213 ( .A(n19245), .B(n19246), .Z(n19238) );
  NOR U19214 ( .A(n19247), .B(n19248), .Z(n19246) );
  XNOR U19215 ( .A(n19245), .B(n19249), .Z(n19247) );
  XNOR U19216 ( .A(n19205), .B(n19212), .Z(n19226) );
  NOR U19217 ( .A(n19169), .B(n19250), .Z(n19212) );
  XOR U19218 ( .A(n19217), .B(n19216), .Z(n19205) );
  XNOR U19219 ( .A(n19251), .B(n19213), .Z(n19216) );
  XOR U19220 ( .A(n19252), .B(n19253), .Z(n19213) );
  AND U19221 ( .A(n19254), .B(n19255), .Z(n19253) );
  XNOR U19222 ( .A(n19256), .B(n19257), .Z(n19254) );
  IV U19223 ( .A(n19252), .Z(n19256) );
  XNOR U19224 ( .A(n19258), .B(n19259), .Z(n19251) );
  NOR U19225 ( .A(n19260), .B(n19261), .Z(n19259) );
  XNOR U19226 ( .A(n19258), .B(n19262), .Z(n19260) );
  XOR U19227 ( .A(n19263), .B(n19264), .Z(n19217) );
  NOR U19228 ( .A(n19265), .B(n19266), .Z(n19264) );
  XNOR U19229 ( .A(n19263), .B(n19267), .Z(n19265) );
  XNOR U19230 ( .A(n19153), .B(n19222), .Z(n19224) );
  XOR U19231 ( .A(n19268), .B(n19269), .Z(n19153) );
  AND U19232 ( .A(n463), .B(n19270), .Z(n19269) );
  XOR U19233 ( .A(n19271), .B(n19268), .Z(n19270) );
  AND U19234 ( .A(n19166), .B(n19169), .Z(n19222) );
  XOR U19235 ( .A(n19272), .B(n19250), .Z(n19169) );
  XNOR U19236 ( .A(p_input[1824]), .B(p_input[2048]), .Z(n19250) );
  XNOR U19237 ( .A(n19237), .B(n19236), .Z(n19272) );
  XNOR U19238 ( .A(n19273), .B(n19244), .Z(n19236) );
  XNOR U19239 ( .A(n19232), .B(n19231), .Z(n19244) );
  XNOR U19240 ( .A(n19274), .B(n19228), .Z(n19231) );
  XNOR U19241 ( .A(p_input[1834]), .B(p_input[2058]), .Z(n19228) );
  XOR U19242 ( .A(p_input[1835]), .B(n6319), .Z(n19274) );
  XOR U19243 ( .A(p_input[1836]), .B(p_input[2060]), .Z(n19232) );
  XOR U19244 ( .A(n19242), .B(n19275), .Z(n19273) );
  IV U19245 ( .A(n19233), .Z(n19275) );
  XOR U19246 ( .A(p_input[1825]), .B(p_input[2049]), .Z(n19233) );
  XNOR U19247 ( .A(n19276), .B(n19249), .Z(n19242) );
  XNOR U19248 ( .A(p_input[1839]), .B(n6322), .Z(n19249) );
  XOR U19249 ( .A(n19239), .B(n19248), .Z(n19276) );
  XOR U19250 ( .A(n19277), .B(n19245), .Z(n19248) );
  XOR U19251 ( .A(p_input[1837]), .B(p_input[2061]), .Z(n19245) );
  XOR U19252 ( .A(p_input[1838]), .B(n6324), .Z(n19277) );
  XOR U19253 ( .A(p_input[1833]), .B(p_input[2057]), .Z(n19239) );
  XOR U19254 ( .A(n19257), .B(n19255), .Z(n19237) );
  XNOR U19255 ( .A(n19278), .B(n19262), .Z(n19255) );
  XOR U19256 ( .A(p_input[1832]), .B(p_input[2056]), .Z(n19262) );
  XOR U19257 ( .A(n19252), .B(n19261), .Z(n19278) );
  XOR U19258 ( .A(n19279), .B(n19258), .Z(n19261) );
  XOR U19259 ( .A(p_input[1830]), .B(p_input[2054]), .Z(n19258) );
  XOR U19260 ( .A(p_input[1831]), .B(n7007), .Z(n19279) );
  XOR U19261 ( .A(p_input[1826]), .B(p_input[2050]), .Z(n19252) );
  XNOR U19262 ( .A(n19267), .B(n19266), .Z(n19257) );
  XOR U19263 ( .A(n19280), .B(n19263), .Z(n19266) );
  XOR U19264 ( .A(p_input[1827]), .B(p_input[2051]), .Z(n19263) );
  XOR U19265 ( .A(p_input[1828]), .B(n7009), .Z(n19280) );
  XOR U19266 ( .A(p_input[1829]), .B(p_input[2053]), .Z(n19267) );
  XOR U19267 ( .A(n19281), .B(n19282), .Z(n19166) );
  AND U19268 ( .A(n463), .B(n19283), .Z(n19282) );
  XNOR U19269 ( .A(n19284), .B(n19281), .Z(n19283) );
  XNOR U19270 ( .A(n19285), .B(n19286), .Z(n463) );
  AND U19271 ( .A(n19287), .B(n19288), .Z(n19286) );
  XOR U19272 ( .A(n19179), .B(n19285), .Z(n19288) );
  AND U19273 ( .A(n19289), .B(n19290), .Z(n19179) );
  XNOR U19274 ( .A(n19176), .B(n19285), .Z(n19287) );
  XOR U19275 ( .A(n19291), .B(n19292), .Z(n19176) );
  AND U19276 ( .A(n467), .B(n19293), .Z(n19292) );
  XOR U19277 ( .A(n19294), .B(n19291), .Z(n19293) );
  XOR U19278 ( .A(n19295), .B(n19296), .Z(n19285) );
  AND U19279 ( .A(n19297), .B(n19298), .Z(n19296) );
  XNOR U19280 ( .A(n19295), .B(n19289), .Z(n19298) );
  IV U19281 ( .A(n19194), .Z(n19289) );
  XOR U19282 ( .A(n19299), .B(n19300), .Z(n19194) );
  XOR U19283 ( .A(n19301), .B(n19290), .Z(n19300) );
  AND U19284 ( .A(n19221), .B(n19302), .Z(n19290) );
  AND U19285 ( .A(n19303), .B(n19304), .Z(n19301) );
  XOR U19286 ( .A(n19305), .B(n19299), .Z(n19303) );
  XNOR U19287 ( .A(n19191), .B(n19295), .Z(n19297) );
  XOR U19288 ( .A(n19306), .B(n19307), .Z(n19191) );
  AND U19289 ( .A(n467), .B(n19308), .Z(n19307) );
  XOR U19290 ( .A(n19309), .B(n19306), .Z(n19308) );
  XOR U19291 ( .A(n19310), .B(n19311), .Z(n19295) );
  AND U19292 ( .A(n19312), .B(n19313), .Z(n19311) );
  XNOR U19293 ( .A(n19310), .B(n19221), .Z(n19313) );
  XOR U19294 ( .A(n19314), .B(n19304), .Z(n19221) );
  XNOR U19295 ( .A(n19315), .B(n19299), .Z(n19304) );
  XOR U19296 ( .A(n19316), .B(n19317), .Z(n19299) );
  AND U19297 ( .A(n19318), .B(n19319), .Z(n19317) );
  XOR U19298 ( .A(n19320), .B(n19316), .Z(n19318) );
  XNOR U19299 ( .A(n19321), .B(n19322), .Z(n19315) );
  AND U19300 ( .A(n19323), .B(n19324), .Z(n19322) );
  XOR U19301 ( .A(n19321), .B(n19325), .Z(n19323) );
  XNOR U19302 ( .A(n19305), .B(n19302), .Z(n19314) );
  AND U19303 ( .A(n19326), .B(n19327), .Z(n19302) );
  XOR U19304 ( .A(n19328), .B(n19329), .Z(n19305) );
  AND U19305 ( .A(n19330), .B(n19331), .Z(n19329) );
  XOR U19306 ( .A(n19328), .B(n19332), .Z(n19330) );
  XNOR U19307 ( .A(n19218), .B(n19310), .Z(n19312) );
  XOR U19308 ( .A(n19333), .B(n19334), .Z(n19218) );
  AND U19309 ( .A(n467), .B(n19335), .Z(n19334) );
  XNOR U19310 ( .A(n19336), .B(n19333), .Z(n19335) );
  XOR U19311 ( .A(n19337), .B(n19338), .Z(n19310) );
  AND U19312 ( .A(n19339), .B(n19340), .Z(n19338) );
  XNOR U19313 ( .A(n19337), .B(n19326), .Z(n19340) );
  IV U19314 ( .A(n19271), .Z(n19326) );
  XNOR U19315 ( .A(n19341), .B(n19319), .Z(n19271) );
  XNOR U19316 ( .A(n19342), .B(n19325), .Z(n19319) );
  XNOR U19317 ( .A(n19343), .B(n19344), .Z(n19325) );
  NOR U19318 ( .A(n19345), .B(n19346), .Z(n19344) );
  XOR U19319 ( .A(n19343), .B(n19347), .Z(n19345) );
  XNOR U19320 ( .A(n19324), .B(n19316), .Z(n19342) );
  XOR U19321 ( .A(n19348), .B(n19349), .Z(n19316) );
  AND U19322 ( .A(n19350), .B(n19351), .Z(n19349) );
  XOR U19323 ( .A(n19348), .B(n19352), .Z(n19350) );
  XNOR U19324 ( .A(n19353), .B(n19321), .Z(n19324) );
  XOR U19325 ( .A(n19354), .B(n19355), .Z(n19321) );
  AND U19326 ( .A(n19356), .B(n19357), .Z(n19355) );
  XNOR U19327 ( .A(n19358), .B(n19359), .Z(n19356) );
  IV U19328 ( .A(n19354), .Z(n19358) );
  XNOR U19329 ( .A(n19360), .B(n19361), .Z(n19353) );
  NOR U19330 ( .A(n19362), .B(n19363), .Z(n19361) );
  XNOR U19331 ( .A(n19360), .B(n19364), .Z(n19362) );
  XNOR U19332 ( .A(n19320), .B(n19327), .Z(n19341) );
  NOR U19333 ( .A(n19284), .B(n19365), .Z(n19327) );
  XOR U19334 ( .A(n19332), .B(n19331), .Z(n19320) );
  XNOR U19335 ( .A(n19366), .B(n19328), .Z(n19331) );
  XOR U19336 ( .A(n19367), .B(n19368), .Z(n19328) );
  AND U19337 ( .A(n19369), .B(n19370), .Z(n19368) );
  XNOR U19338 ( .A(n19371), .B(n19372), .Z(n19369) );
  IV U19339 ( .A(n19367), .Z(n19371) );
  XNOR U19340 ( .A(n19373), .B(n19374), .Z(n19366) );
  NOR U19341 ( .A(n19375), .B(n19376), .Z(n19374) );
  XNOR U19342 ( .A(n19373), .B(n19377), .Z(n19375) );
  XOR U19343 ( .A(n19378), .B(n19379), .Z(n19332) );
  NOR U19344 ( .A(n19380), .B(n19381), .Z(n19379) );
  XNOR U19345 ( .A(n19378), .B(n19382), .Z(n19380) );
  XNOR U19346 ( .A(n19268), .B(n19337), .Z(n19339) );
  XOR U19347 ( .A(n19383), .B(n19384), .Z(n19268) );
  AND U19348 ( .A(n467), .B(n19385), .Z(n19384) );
  XOR U19349 ( .A(n19386), .B(n19383), .Z(n19385) );
  AND U19350 ( .A(n19281), .B(n19284), .Z(n19337) );
  XOR U19351 ( .A(n19387), .B(n19365), .Z(n19284) );
  XNOR U19352 ( .A(p_input[1840]), .B(p_input[2048]), .Z(n19365) );
  XNOR U19353 ( .A(n19352), .B(n19351), .Z(n19387) );
  XNOR U19354 ( .A(n19388), .B(n19359), .Z(n19351) );
  XNOR U19355 ( .A(n19347), .B(n19346), .Z(n19359) );
  XNOR U19356 ( .A(n19389), .B(n19343), .Z(n19346) );
  XNOR U19357 ( .A(p_input[1850]), .B(p_input[2058]), .Z(n19343) );
  XOR U19358 ( .A(p_input[1851]), .B(n6319), .Z(n19389) );
  XOR U19359 ( .A(p_input[1852]), .B(p_input[2060]), .Z(n19347) );
  XOR U19360 ( .A(n19357), .B(n19390), .Z(n19388) );
  IV U19361 ( .A(n19348), .Z(n19390) );
  XOR U19362 ( .A(p_input[1841]), .B(p_input[2049]), .Z(n19348) );
  XNOR U19363 ( .A(n19391), .B(n19364), .Z(n19357) );
  XNOR U19364 ( .A(p_input[1855]), .B(n6322), .Z(n19364) );
  XOR U19365 ( .A(n19354), .B(n19363), .Z(n19391) );
  XOR U19366 ( .A(n19392), .B(n19360), .Z(n19363) );
  XOR U19367 ( .A(p_input[1853]), .B(p_input[2061]), .Z(n19360) );
  XOR U19368 ( .A(p_input[1854]), .B(n6324), .Z(n19392) );
  XOR U19369 ( .A(p_input[1849]), .B(p_input[2057]), .Z(n19354) );
  XOR U19370 ( .A(n19372), .B(n19370), .Z(n19352) );
  XNOR U19371 ( .A(n19393), .B(n19377), .Z(n19370) );
  XOR U19372 ( .A(p_input[1848]), .B(p_input[2056]), .Z(n19377) );
  XOR U19373 ( .A(n19367), .B(n19376), .Z(n19393) );
  XOR U19374 ( .A(n19394), .B(n19373), .Z(n19376) );
  XOR U19375 ( .A(p_input[1846]), .B(p_input[2054]), .Z(n19373) );
  XOR U19376 ( .A(p_input[1847]), .B(n7007), .Z(n19394) );
  XOR U19377 ( .A(p_input[1842]), .B(p_input[2050]), .Z(n19367) );
  XNOR U19378 ( .A(n19382), .B(n19381), .Z(n19372) );
  XOR U19379 ( .A(n19395), .B(n19378), .Z(n19381) );
  XOR U19380 ( .A(p_input[1843]), .B(p_input[2051]), .Z(n19378) );
  XOR U19381 ( .A(p_input[1844]), .B(n7009), .Z(n19395) );
  XOR U19382 ( .A(p_input[1845]), .B(p_input[2053]), .Z(n19382) );
  XOR U19383 ( .A(n19396), .B(n19397), .Z(n19281) );
  AND U19384 ( .A(n467), .B(n19398), .Z(n19397) );
  XNOR U19385 ( .A(n19399), .B(n19396), .Z(n19398) );
  XNOR U19386 ( .A(n19400), .B(n19401), .Z(n467) );
  AND U19387 ( .A(n19402), .B(n19403), .Z(n19401) );
  XOR U19388 ( .A(n19294), .B(n19400), .Z(n19403) );
  AND U19389 ( .A(n19404), .B(n19405), .Z(n19294) );
  XNOR U19390 ( .A(n19291), .B(n19400), .Z(n19402) );
  XOR U19391 ( .A(n19406), .B(n19407), .Z(n19291) );
  AND U19392 ( .A(n19408), .B(n471), .Z(n19407) );
  AND U19393 ( .A(n19406), .B(n19409), .Z(n19408) );
  XOR U19394 ( .A(n19410), .B(n19411), .Z(n19400) );
  AND U19395 ( .A(n19412), .B(n19413), .Z(n19411) );
  XNOR U19396 ( .A(n19410), .B(n19404), .Z(n19413) );
  IV U19397 ( .A(n19309), .Z(n19404) );
  XOR U19398 ( .A(n19414), .B(n19415), .Z(n19309) );
  XOR U19399 ( .A(n19416), .B(n19405), .Z(n19415) );
  AND U19400 ( .A(n19336), .B(n19417), .Z(n19405) );
  AND U19401 ( .A(n19418), .B(n19419), .Z(n19416) );
  XOR U19402 ( .A(n19420), .B(n19414), .Z(n19418) );
  XNOR U19403 ( .A(n19306), .B(n19410), .Z(n19412) );
  XOR U19404 ( .A(n19421), .B(n19422), .Z(n19306) );
  AND U19405 ( .A(n471), .B(n19423), .Z(n19422) );
  XOR U19406 ( .A(n19424), .B(n19421), .Z(n19423) );
  XOR U19407 ( .A(n19425), .B(n19426), .Z(n19410) );
  AND U19408 ( .A(n19427), .B(n19428), .Z(n19426) );
  XNOR U19409 ( .A(n19425), .B(n19336), .Z(n19428) );
  XOR U19410 ( .A(n19429), .B(n19419), .Z(n19336) );
  XNOR U19411 ( .A(n19430), .B(n19414), .Z(n19419) );
  XOR U19412 ( .A(n19431), .B(n19432), .Z(n19414) );
  AND U19413 ( .A(n19433), .B(n19434), .Z(n19432) );
  XOR U19414 ( .A(n19435), .B(n19431), .Z(n19433) );
  XNOR U19415 ( .A(n19436), .B(n19437), .Z(n19430) );
  AND U19416 ( .A(n19438), .B(n19439), .Z(n19437) );
  XOR U19417 ( .A(n19436), .B(n19440), .Z(n19438) );
  XNOR U19418 ( .A(n19420), .B(n19417), .Z(n19429) );
  AND U19419 ( .A(n19441), .B(n19442), .Z(n19417) );
  XOR U19420 ( .A(n19443), .B(n19444), .Z(n19420) );
  AND U19421 ( .A(n19445), .B(n19446), .Z(n19444) );
  XOR U19422 ( .A(n19443), .B(n19447), .Z(n19445) );
  XNOR U19423 ( .A(n19333), .B(n19425), .Z(n19427) );
  XOR U19424 ( .A(n19448), .B(n19449), .Z(n19333) );
  AND U19425 ( .A(n471), .B(n19450), .Z(n19449) );
  XNOR U19426 ( .A(n19451), .B(n19448), .Z(n19450) );
  XOR U19427 ( .A(n19452), .B(n19453), .Z(n19425) );
  AND U19428 ( .A(n19454), .B(n19455), .Z(n19453) );
  XNOR U19429 ( .A(n19452), .B(n19441), .Z(n19455) );
  IV U19430 ( .A(n19386), .Z(n19441) );
  XNOR U19431 ( .A(n19456), .B(n19434), .Z(n19386) );
  XNOR U19432 ( .A(n19457), .B(n19440), .Z(n19434) );
  XNOR U19433 ( .A(n19458), .B(n19459), .Z(n19440) );
  NOR U19434 ( .A(n19460), .B(n19461), .Z(n19459) );
  XOR U19435 ( .A(n19458), .B(n19462), .Z(n19460) );
  XNOR U19436 ( .A(n19439), .B(n19431), .Z(n19457) );
  XOR U19437 ( .A(n19463), .B(n19464), .Z(n19431) );
  AND U19438 ( .A(n19465), .B(n19466), .Z(n19464) );
  XOR U19439 ( .A(n19463), .B(n19467), .Z(n19465) );
  XNOR U19440 ( .A(n19468), .B(n19436), .Z(n19439) );
  XOR U19441 ( .A(n19469), .B(n19470), .Z(n19436) );
  AND U19442 ( .A(n19471), .B(n19472), .Z(n19470) );
  XNOR U19443 ( .A(n19473), .B(n19474), .Z(n19471) );
  IV U19444 ( .A(n19469), .Z(n19473) );
  XNOR U19445 ( .A(n19475), .B(n19476), .Z(n19468) );
  NOR U19446 ( .A(n19477), .B(n19478), .Z(n19476) );
  XNOR U19447 ( .A(n19475), .B(n19479), .Z(n19477) );
  XNOR U19448 ( .A(n19435), .B(n19442), .Z(n19456) );
  NOR U19449 ( .A(n19399), .B(n19480), .Z(n19442) );
  XOR U19450 ( .A(n19447), .B(n19446), .Z(n19435) );
  XNOR U19451 ( .A(n19481), .B(n19443), .Z(n19446) );
  XOR U19452 ( .A(n19482), .B(n19483), .Z(n19443) );
  AND U19453 ( .A(n19484), .B(n19485), .Z(n19483) );
  XNOR U19454 ( .A(n19486), .B(n19487), .Z(n19484) );
  IV U19455 ( .A(n19482), .Z(n19486) );
  XNOR U19456 ( .A(n19488), .B(n19489), .Z(n19481) );
  NOR U19457 ( .A(n19490), .B(n19491), .Z(n19489) );
  XNOR U19458 ( .A(n19488), .B(n19492), .Z(n19490) );
  XOR U19459 ( .A(n19493), .B(n19494), .Z(n19447) );
  NOR U19460 ( .A(n19495), .B(n19496), .Z(n19494) );
  XNOR U19461 ( .A(n19493), .B(n19497), .Z(n19495) );
  XNOR U19462 ( .A(n19383), .B(n19452), .Z(n19454) );
  XOR U19463 ( .A(n19498), .B(n19499), .Z(n19383) );
  AND U19464 ( .A(n471), .B(n19500), .Z(n19499) );
  XOR U19465 ( .A(n19501), .B(n19498), .Z(n19500) );
  AND U19466 ( .A(n19396), .B(n19399), .Z(n19452) );
  XOR U19467 ( .A(n19502), .B(n19480), .Z(n19399) );
  XNOR U19468 ( .A(p_input[1856]), .B(p_input[2048]), .Z(n19480) );
  XNOR U19469 ( .A(n19467), .B(n19466), .Z(n19502) );
  XNOR U19470 ( .A(n19503), .B(n19474), .Z(n19466) );
  XNOR U19471 ( .A(n19462), .B(n19461), .Z(n19474) );
  XNOR U19472 ( .A(n19504), .B(n19458), .Z(n19461) );
  XNOR U19473 ( .A(p_input[1866]), .B(p_input[2058]), .Z(n19458) );
  XOR U19474 ( .A(p_input[1867]), .B(n6319), .Z(n19504) );
  XOR U19475 ( .A(p_input[1868]), .B(p_input[2060]), .Z(n19462) );
  XOR U19476 ( .A(n19472), .B(n19505), .Z(n19503) );
  IV U19477 ( .A(n19463), .Z(n19505) );
  XOR U19478 ( .A(p_input[1857]), .B(p_input[2049]), .Z(n19463) );
  XNOR U19479 ( .A(n19506), .B(n19479), .Z(n19472) );
  XNOR U19480 ( .A(p_input[1871]), .B(n6322), .Z(n19479) );
  XOR U19481 ( .A(n19469), .B(n19478), .Z(n19506) );
  XOR U19482 ( .A(n19507), .B(n19475), .Z(n19478) );
  XOR U19483 ( .A(p_input[1869]), .B(p_input[2061]), .Z(n19475) );
  XOR U19484 ( .A(p_input[1870]), .B(n6324), .Z(n19507) );
  XOR U19485 ( .A(p_input[1865]), .B(p_input[2057]), .Z(n19469) );
  XOR U19486 ( .A(n19487), .B(n19485), .Z(n19467) );
  XNOR U19487 ( .A(n19508), .B(n19492), .Z(n19485) );
  XOR U19488 ( .A(p_input[1864]), .B(p_input[2056]), .Z(n19492) );
  XOR U19489 ( .A(n19482), .B(n19491), .Z(n19508) );
  XOR U19490 ( .A(n19509), .B(n19488), .Z(n19491) );
  XOR U19491 ( .A(p_input[1862]), .B(p_input[2054]), .Z(n19488) );
  XOR U19492 ( .A(p_input[1863]), .B(n7007), .Z(n19509) );
  XOR U19493 ( .A(p_input[1858]), .B(p_input[2050]), .Z(n19482) );
  XNOR U19494 ( .A(n19497), .B(n19496), .Z(n19487) );
  XOR U19495 ( .A(n19510), .B(n19493), .Z(n19496) );
  XOR U19496 ( .A(p_input[1859]), .B(p_input[2051]), .Z(n19493) );
  XOR U19497 ( .A(p_input[1860]), .B(n7009), .Z(n19510) );
  XOR U19498 ( .A(p_input[1861]), .B(p_input[2053]), .Z(n19497) );
  XOR U19499 ( .A(n19511), .B(n19512), .Z(n19396) );
  AND U19500 ( .A(n471), .B(n19513), .Z(n19512) );
  XNOR U19501 ( .A(n19514), .B(n19511), .Z(n19513) );
  XNOR U19502 ( .A(n19515), .B(n19516), .Z(n471) );
  AND U19503 ( .A(n19517), .B(n19518), .Z(n19516) );
  XNOR U19504 ( .A(n19409), .B(n19515), .Z(n19518) );
  IV U19505 ( .A(n19519), .Z(n19409) );
  AND U19506 ( .A(n19520), .B(n19521), .Z(n19519) );
  XNOR U19507 ( .A(n19515), .B(n19406), .Z(n19517) );
  AND U19508 ( .A(n19522), .B(n19523), .Z(n19406) );
  XOR U19509 ( .A(n19524), .B(n19525), .Z(n19515) );
  AND U19510 ( .A(n19526), .B(n19527), .Z(n19525) );
  XNOR U19511 ( .A(n19524), .B(n19520), .Z(n19527) );
  IV U19512 ( .A(n19424), .Z(n19520) );
  XOR U19513 ( .A(n19528), .B(n19529), .Z(n19424) );
  XOR U19514 ( .A(n19530), .B(n19521), .Z(n19529) );
  AND U19515 ( .A(n19451), .B(n19531), .Z(n19521) );
  AND U19516 ( .A(n19532), .B(n19533), .Z(n19530) );
  XOR U19517 ( .A(n19534), .B(n19528), .Z(n19532) );
  XNOR U19518 ( .A(n19421), .B(n19524), .Z(n19526) );
  XOR U19519 ( .A(n19535), .B(n19536), .Z(n19421) );
  AND U19520 ( .A(n475), .B(n19537), .Z(n19536) );
  XOR U19521 ( .A(n19538), .B(n19535), .Z(n19537) );
  XOR U19522 ( .A(n19539), .B(n19540), .Z(n19524) );
  AND U19523 ( .A(n19541), .B(n19542), .Z(n19540) );
  XNOR U19524 ( .A(n19539), .B(n19451), .Z(n19542) );
  XOR U19525 ( .A(n19543), .B(n19533), .Z(n19451) );
  XNOR U19526 ( .A(n19544), .B(n19528), .Z(n19533) );
  XOR U19527 ( .A(n19545), .B(n19546), .Z(n19528) );
  AND U19528 ( .A(n19547), .B(n19548), .Z(n19546) );
  XOR U19529 ( .A(n19549), .B(n19545), .Z(n19547) );
  XNOR U19530 ( .A(n19550), .B(n19551), .Z(n19544) );
  AND U19531 ( .A(n19552), .B(n19553), .Z(n19551) );
  XOR U19532 ( .A(n19550), .B(n19554), .Z(n19552) );
  XNOR U19533 ( .A(n19534), .B(n19531), .Z(n19543) );
  AND U19534 ( .A(n19555), .B(n19556), .Z(n19531) );
  XOR U19535 ( .A(n19557), .B(n19558), .Z(n19534) );
  AND U19536 ( .A(n19559), .B(n19560), .Z(n19558) );
  XOR U19537 ( .A(n19557), .B(n19561), .Z(n19559) );
  XNOR U19538 ( .A(n19448), .B(n19539), .Z(n19541) );
  XOR U19539 ( .A(n19562), .B(n19563), .Z(n19448) );
  AND U19540 ( .A(n475), .B(n19564), .Z(n19563) );
  XNOR U19541 ( .A(n19565), .B(n19562), .Z(n19564) );
  XOR U19542 ( .A(n19566), .B(n19567), .Z(n19539) );
  AND U19543 ( .A(n19568), .B(n19569), .Z(n19567) );
  XNOR U19544 ( .A(n19566), .B(n19555), .Z(n19569) );
  IV U19545 ( .A(n19501), .Z(n19555) );
  XNOR U19546 ( .A(n19570), .B(n19548), .Z(n19501) );
  XNOR U19547 ( .A(n19571), .B(n19554), .Z(n19548) );
  XNOR U19548 ( .A(n19572), .B(n19573), .Z(n19554) );
  NOR U19549 ( .A(n19574), .B(n19575), .Z(n19573) );
  XOR U19550 ( .A(n19572), .B(n19576), .Z(n19574) );
  XNOR U19551 ( .A(n19553), .B(n19545), .Z(n19571) );
  XOR U19552 ( .A(n19577), .B(n19578), .Z(n19545) );
  AND U19553 ( .A(n19579), .B(n19580), .Z(n19578) );
  XOR U19554 ( .A(n19577), .B(n19581), .Z(n19579) );
  XNOR U19555 ( .A(n19582), .B(n19550), .Z(n19553) );
  XOR U19556 ( .A(n19583), .B(n19584), .Z(n19550) );
  AND U19557 ( .A(n19585), .B(n19586), .Z(n19584) );
  XNOR U19558 ( .A(n19587), .B(n19588), .Z(n19585) );
  IV U19559 ( .A(n19583), .Z(n19587) );
  XNOR U19560 ( .A(n19589), .B(n19590), .Z(n19582) );
  NOR U19561 ( .A(n19591), .B(n19592), .Z(n19590) );
  XNOR U19562 ( .A(n19589), .B(n19593), .Z(n19591) );
  XNOR U19563 ( .A(n19549), .B(n19556), .Z(n19570) );
  NOR U19564 ( .A(n19514), .B(n19594), .Z(n19556) );
  XOR U19565 ( .A(n19561), .B(n19560), .Z(n19549) );
  XNOR U19566 ( .A(n19595), .B(n19557), .Z(n19560) );
  XOR U19567 ( .A(n19596), .B(n19597), .Z(n19557) );
  AND U19568 ( .A(n19598), .B(n19599), .Z(n19597) );
  XNOR U19569 ( .A(n19600), .B(n19601), .Z(n19598) );
  IV U19570 ( .A(n19596), .Z(n19600) );
  XNOR U19571 ( .A(n19602), .B(n19603), .Z(n19595) );
  NOR U19572 ( .A(n19604), .B(n19605), .Z(n19603) );
  XNOR U19573 ( .A(n19602), .B(n19606), .Z(n19604) );
  XOR U19574 ( .A(n19607), .B(n19608), .Z(n19561) );
  NOR U19575 ( .A(n19609), .B(n19610), .Z(n19608) );
  XNOR U19576 ( .A(n19607), .B(n19611), .Z(n19609) );
  XNOR U19577 ( .A(n19498), .B(n19566), .Z(n19568) );
  XOR U19578 ( .A(n19612), .B(n19613), .Z(n19498) );
  AND U19579 ( .A(n475), .B(n19614), .Z(n19613) );
  XOR U19580 ( .A(n19615), .B(n19612), .Z(n19614) );
  AND U19581 ( .A(n19511), .B(n19514), .Z(n19566) );
  XOR U19582 ( .A(n19616), .B(n19594), .Z(n19514) );
  XNOR U19583 ( .A(p_input[1872]), .B(p_input[2048]), .Z(n19594) );
  XNOR U19584 ( .A(n19581), .B(n19580), .Z(n19616) );
  XNOR U19585 ( .A(n19617), .B(n19588), .Z(n19580) );
  XNOR U19586 ( .A(n19576), .B(n19575), .Z(n19588) );
  XNOR U19587 ( .A(n19618), .B(n19572), .Z(n19575) );
  XNOR U19588 ( .A(p_input[1882]), .B(p_input[2058]), .Z(n19572) );
  XOR U19589 ( .A(p_input[1883]), .B(n6319), .Z(n19618) );
  XOR U19590 ( .A(p_input[1884]), .B(p_input[2060]), .Z(n19576) );
  XOR U19591 ( .A(n19586), .B(n19619), .Z(n19617) );
  IV U19592 ( .A(n19577), .Z(n19619) );
  XOR U19593 ( .A(p_input[1873]), .B(p_input[2049]), .Z(n19577) );
  XNOR U19594 ( .A(n19620), .B(n19593), .Z(n19586) );
  XNOR U19595 ( .A(p_input[1887]), .B(n6322), .Z(n19593) );
  XOR U19596 ( .A(n19583), .B(n19592), .Z(n19620) );
  XOR U19597 ( .A(n19621), .B(n19589), .Z(n19592) );
  XOR U19598 ( .A(p_input[1885]), .B(p_input[2061]), .Z(n19589) );
  XOR U19599 ( .A(p_input[1886]), .B(n6324), .Z(n19621) );
  XOR U19600 ( .A(p_input[1881]), .B(p_input[2057]), .Z(n19583) );
  XOR U19601 ( .A(n19601), .B(n19599), .Z(n19581) );
  XNOR U19602 ( .A(n19622), .B(n19606), .Z(n19599) );
  XOR U19603 ( .A(p_input[1880]), .B(p_input[2056]), .Z(n19606) );
  XOR U19604 ( .A(n19596), .B(n19605), .Z(n19622) );
  XOR U19605 ( .A(n19623), .B(n19602), .Z(n19605) );
  XOR U19606 ( .A(p_input[1878]), .B(p_input[2054]), .Z(n19602) );
  XOR U19607 ( .A(p_input[1879]), .B(n7007), .Z(n19623) );
  XOR U19608 ( .A(p_input[1874]), .B(p_input[2050]), .Z(n19596) );
  XNOR U19609 ( .A(n19611), .B(n19610), .Z(n19601) );
  XOR U19610 ( .A(n19624), .B(n19607), .Z(n19610) );
  XOR U19611 ( .A(p_input[1875]), .B(p_input[2051]), .Z(n19607) );
  XOR U19612 ( .A(p_input[1876]), .B(n7009), .Z(n19624) );
  XOR U19613 ( .A(p_input[1877]), .B(p_input[2053]), .Z(n19611) );
  XOR U19614 ( .A(n19625), .B(n19626), .Z(n19511) );
  AND U19615 ( .A(n475), .B(n19627), .Z(n19626) );
  XNOR U19616 ( .A(n19628), .B(n19625), .Z(n19627) );
  XNOR U19617 ( .A(n19629), .B(n19630), .Z(n475) );
  NOR U19618 ( .A(n19631), .B(n19632), .Z(n19630) );
  XOR U19619 ( .A(n19523), .B(n19629), .Z(n19632) );
  AND U19620 ( .A(n19633), .B(n19634), .Z(n19523) );
  NOR U19621 ( .A(n19629), .B(n19522), .Z(n19631) );
  AND U19622 ( .A(n19635), .B(n19636), .Z(n19522) );
  XOR U19623 ( .A(n19637), .B(n19638), .Z(n19629) );
  AND U19624 ( .A(n19639), .B(n19640), .Z(n19638) );
  XNOR U19625 ( .A(n19637), .B(n19635), .Z(n19640) );
  IV U19626 ( .A(n19538), .Z(n19635) );
  XOR U19627 ( .A(n19641), .B(n19642), .Z(n19538) );
  XOR U19628 ( .A(n19643), .B(n19636), .Z(n19642) );
  AND U19629 ( .A(n19565), .B(n19644), .Z(n19636) );
  AND U19630 ( .A(n19645), .B(n19646), .Z(n19643) );
  XOR U19631 ( .A(n19647), .B(n19641), .Z(n19645) );
  XNOR U19632 ( .A(n19535), .B(n19637), .Z(n19639) );
  XOR U19633 ( .A(n19648), .B(n19649), .Z(n19535) );
  AND U19634 ( .A(n479), .B(n19650), .Z(n19649) );
  XOR U19635 ( .A(n19651), .B(n19648), .Z(n19650) );
  XOR U19636 ( .A(n19652), .B(n19653), .Z(n19637) );
  AND U19637 ( .A(n19654), .B(n19655), .Z(n19653) );
  XNOR U19638 ( .A(n19652), .B(n19565), .Z(n19655) );
  XOR U19639 ( .A(n19656), .B(n19646), .Z(n19565) );
  XNOR U19640 ( .A(n19657), .B(n19641), .Z(n19646) );
  XOR U19641 ( .A(n19658), .B(n19659), .Z(n19641) );
  AND U19642 ( .A(n19660), .B(n19661), .Z(n19659) );
  XOR U19643 ( .A(n19662), .B(n19658), .Z(n19660) );
  XNOR U19644 ( .A(n19663), .B(n19664), .Z(n19657) );
  AND U19645 ( .A(n19665), .B(n19666), .Z(n19664) );
  XOR U19646 ( .A(n19663), .B(n19667), .Z(n19665) );
  XNOR U19647 ( .A(n19647), .B(n19644), .Z(n19656) );
  AND U19648 ( .A(n19668), .B(n19669), .Z(n19644) );
  XOR U19649 ( .A(n19670), .B(n19671), .Z(n19647) );
  AND U19650 ( .A(n19672), .B(n19673), .Z(n19671) );
  XOR U19651 ( .A(n19670), .B(n19674), .Z(n19672) );
  XNOR U19652 ( .A(n19562), .B(n19652), .Z(n19654) );
  XOR U19653 ( .A(n19675), .B(n19676), .Z(n19562) );
  AND U19654 ( .A(n479), .B(n19677), .Z(n19676) );
  XNOR U19655 ( .A(n19678), .B(n19675), .Z(n19677) );
  XOR U19656 ( .A(n19679), .B(n19680), .Z(n19652) );
  AND U19657 ( .A(n19681), .B(n19682), .Z(n19680) );
  XNOR U19658 ( .A(n19679), .B(n19668), .Z(n19682) );
  IV U19659 ( .A(n19615), .Z(n19668) );
  XNOR U19660 ( .A(n19683), .B(n19661), .Z(n19615) );
  XNOR U19661 ( .A(n19684), .B(n19667), .Z(n19661) );
  XNOR U19662 ( .A(n19685), .B(n19686), .Z(n19667) );
  NOR U19663 ( .A(n19687), .B(n19688), .Z(n19686) );
  XOR U19664 ( .A(n19685), .B(n19689), .Z(n19687) );
  XNOR U19665 ( .A(n19666), .B(n19658), .Z(n19684) );
  XOR U19666 ( .A(n19690), .B(n19691), .Z(n19658) );
  AND U19667 ( .A(n19692), .B(n19693), .Z(n19691) );
  XOR U19668 ( .A(n19690), .B(n19694), .Z(n19692) );
  XNOR U19669 ( .A(n19695), .B(n19663), .Z(n19666) );
  XOR U19670 ( .A(n19696), .B(n19697), .Z(n19663) );
  AND U19671 ( .A(n19698), .B(n19699), .Z(n19697) );
  XNOR U19672 ( .A(n19700), .B(n19701), .Z(n19698) );
  IV U19673 ( .A(n19696), .Z(n19700) );
  XNOR U19674 ( .A(n19702), .B(n19703), .Z(n19695) );
  NOR U19675 ( .A(n19704), .B(n19705), .Z(n19703) );
  XNOR U19676 ( .A(n19702), .B(n19706), .Z(n19704) );
  XNOR U19677 ( .A(n19662), .B(n19669), .Z(n19683) );
  NOR U19678 ( .A(n19628), .B(n19707), .Z(n19669) );
  XOR U19679 ( .A(n19674), .B(n19673), .Z(n19662) );
  XNOR U19680 ( .A(n19708), .B(n19670), .Z(n19673) );
  XOR U19681 ( .A(n19709), .B(n19710), .Z(n19670) );
  AND U19682 ( .A(n19711), .B(n19712), .Z(n19710) );
  XNOR U19683 ( .A(n19713), .B(n19714), .Z(n19711) );
  IV U19684 ( .A(n19709), .Z(n19713) );
  XNOR U19685 ( .A(n19715), .B(n19716), .Z(n19708) );
  NOR U19686 ( .A(n19717), .B(n19718), .Z(n19716) );
  XNOR U19687 ( .A(n19715), .B(n19719), .Z(n19717) );
  XOR U19688 ( .A(n19720), .B(n19721), .Z(n19674) );
  NOR U19689 ( .A(n19722), .B(n19723), .Z(n19721) );
  XNOR U19690 ( .A(n19720), .B(n19724), .Z(n19722) );
  XNOR U19691 ( .A(n19612), .B(n19679), .Z(n19681) );
  XOR U19692 ( .A(n19725), .B(n19726), .Z(n19612) );
  AND U19693 ( .A(n479), .B(n19727), .Z(n19726) );
  XOR U19694 ( .A(n19728), .B(n19725), .Z(n19727) );
  AND U19695 ( .A(n19625), .B(n19628), .Z(n19679) );
  XOR U19696 ( .A(n19729), .B(n19707), .Z(n19628) );
  XNOR U19697 ( .A(p_input[1888]), .B(p_input[2048]), .Z(n19707) );
  XNOR U19698 ( .A(n19694), .B(n19693), .Z(n19729) );
  XNOR U19699 ( .A(n19730), .B(n19701), .Z(n19693) );
  XNOR U19700 ( .A(n19689), .B(n19688), .Z(n19701) );
  XNOR U19701 ( .A(n19731), .B(n19685), .Z(n19688) );
  XNOR U19702 ( .A(p_input[1898]), .B(p_input[2058]), .Z(n19685) );
  XOR U19703 ( .A(p_input[1899]), .B(n6319), .Z(n19731) );
  XOR U19704 ( .A(p_input[1900]), .B(p_input[2060]), .Z(n19689) );
  XOR U19705 ( .A(n19699), .B(n19732), .Z(n19730) );
  IV U19706 ( .A(n19690), .Z(n19732) );
  XOR U19707 ( .A(p_input[1889]), .B(p_input[2049]), .Z(n19690) );
  XNOR U19708 ( .A(n19733), .B(n19706), .Z(n19699) );
  XNOR U19709 ( .A(p_input[1903]), .B(n6322), .Z(n19706) );
  XOR U19710 ( .A(n19696), .B(n19705), .Z(n19733) );
  XOR U19711 ( .A(n19734), .B(n19702), .Z(n19705) );
  XOR U19712 ( .A(p_input[1901]), .B(p_input[2061]), .Z(n19702) );
  XOR U19713 ( .A(p_input[1902]), .B(n6324), .Z(n19734) );
  XOR U19714 ( .A(p_input[1897]), .B(p_input[2057]), .Z(n19696) );
  XOR U19715 ( .A(n19714), .B(n19712), .Z(n19694) );
  XNOR U19716 ( .A(n19735), .B(n19719), .Z(n19712) );
  XOR U19717 ( .A(p_input[1896]), .B(p_input[2056]), .Z(n19719) );
  XOR U19718 ( .A(n19709), .B(n19718), .Z(n19735) );
  XOR U19719 ( .A(n19736), .B(n19715), .Z(n19718) );
  XOR U19720 ( .A(p_input[1894]), .B(p_input[2054]), .Z(n19715) );
  XOR U19721 ( .A(p_input[1895]), .B(n7007), .Z(n19736) );
  XOR U19722 ( .A(p_input[1890]), .B(p_input[2050]), .Z(n19709) );
  XNOR U19723 ( .A(n19724), .B(n19723), .Z(n19714) );
  XOR U19724 ( .A(n19737), .B(n19720), .Z(n19723) );
  XOR U19725 ( .A(p_input[1891]), .B(p_input[2051]), .Z(n19720) );
  XOR U19726 ( .A(p_input[1892]), .B(n7009), .Z(n19737) );
  XOR U19727 ( .A(p_input[1893]), .B(p_input[2053]), .Z(n19724) );
  XOR U19728 ( .A(n19738), .B(n19739), .Z(n19625) );
  AND U19729 ( .A(n479), .B(n19740), .Z(n19739) );
  XNOR U19730 ( .A(n19741), .B(n19738), .Z(n19740) );
  XNOR U19731 ( .A(n19742), .B(n19743), .Z(n479) );
  NOR U19732 ( .A(n19744), .B(n19745), .Z(n19743) );
  XOR U19733 ( .A(n19634), .B(n19742), .Z(n19745) );
  AND U19734 ( .A(n19746), .B(n19747), .Z(n19634) );
  NOR U19735 ( .A(n19742), .B(n19633), .Z(n19744) );
  AND U19736 ( .A(n19748), .B(n19749), .Z(n19633) );
  XOR U19737 ( .A(n19750), .B(n19751), .Z(n19742) );
  AND U19738 ( .A(n19752), .B(n19753), .Z(n19751) );
  XNOR U19739 ( .A(n19750), .B(n19748), .Z(n19753) );
  IV U19740 ( .A(n19651), .Z(n19748) );
  XOR U19741 ( .A(n19754), .B(n19755), .Z(n19651) );
  XOR U19742 ( .A(n19756), .B(n19749), .Z(n19755) );
  AND U19743 ( .A(n19678), .B(n19757), .Z(n19749) );
  AND U19744 ( .A(n19758), .B(n19759), .Z(n19756) );
  XOR U19745 ( .A(n19760), .B(n19754), .Z(n19758) );
  XNOR U19746 ( .A(n19648), .B(n19750), .Z(n19752) );
  XOR U19747 ( .A(n19761), .B(n19762), .Z(n19648) );
  AND U19748 ( .A(n483), .B(n19763), .Z(n19762) );
  XOR U19749 ( .A(n19764), .B(n19761), .Z(n19763) );
  XOR U19750 ( .A(n19765), .B(n19766), .Z(n19750) );
  AND U19751 ( .A(n19767), .B(n19768), .Z(n19766) );
  XNOR U19752 ( .A(n19765), .B(n19678), .Z(n19768) );
  XOR U19753 ( .A(n19769), .B(n19759), .Z(n19678) );
  XNOR U19754 ( .A(n19770), .B(n19754), .Z(n19759) );
  XOR U19755 ( .A(n19771), .B(n19772), .Z(n19754) );
  AND U19756 ( .A(n19773), .B(n19774), .Z(n19772) );
  XOR U19757 ( .A(n19775), .B(n19771), .Z(n19773) );
  XNOR U19758 ( .A(n19776), .B(n19777), .Z(n19770) );
  AND U19759 ( .A(n19778), .B(n19779), .Z(n19777) );
  XOR U19760 ( .A(n19776), .B(n19780), .Z(n19778) );
  XNOR U19761 ( .A(n19760), .B(n19757), .Z(n19769) );
  AND U19762 ( .A(n19781), .B(n19782), .Z(n19757) );
  XOR U19763 ( .A(n19783), .B(n19784), .Z(n19760) );
  AND U19764 ( .A(n19785), .B(n19786), .Z(n19784) );
  XOR U19765 ( .A(n19783), .B(n19787), .Z(n19785) );
  XNOR U19766 ( .A(n19675), .B(n19765), .Z(n19767) );
  XOR U19767 ( .A(n19788), .B(n19789), .Z(n19675) );
  AND U19768 ( .A(n483), .B(n19790), .Z(n19789) );
  XNOR U19769 ( .A(n19791), .B(n19788), .Z(n19790) );
  XOR U19770 ( .A(n19792), .B(n19793), .Z(n19765) );
  AND U19771 ( .A(n19794), .B(n19795), .Z(n19793) );
  XNOR U19772 ( .A(n19792), .B(n19781), .Z(n19795) );
  IV U19773 ( .A(n19728), .Z(n19781) );
  XNOR U19774 ( .A(n19796), .B(n19774), .Z(n19728) );
  XNOR U19775 ( .A(n19797), .B(n19780), .Z(n19774) );
  XNOR U19776 ( .A(n19798), .B(n19799), .Z(n19780) );
  NOR U19777 ( .A(n19800), .B(n19801), .Z(n19799) );
  XOR U19778 ( .A(n19798), .B(n19802), .Z(n19800) );
  XNOR U19779 ( .A(n19779), .B(n19771), .Z(n19797) );
  XOR U19780 ( .A(n19803), .B(n19804), .Z(n19771) );
  AND U19781 ( .A(n19805), .B(n19806), .Z(n19804) );
  XOR U19782 ( .A(n19803), .B(n19807), .Z(n19805) );
  XNOR U19783 ( .A(n19808), .B(n19776), .Z(n19779) );
  XOR U19784 ( .A(n19809), .B(n19810), .Z(n19776) );
  AND U19785 ( .A(n19811), .B(n19812), .Z(n19810) );
  XNOR U19786 ( .A(n19813), .B(n19814), .Z(n19811) );
  IV U19787 ( .A(n19809), .Z(n19813) );
  XNOR U19788 ( .A(n19815), .B(n19816), .Z(n19808) );
  NOR U19789 ( .A(n19817), .B(n19818), .Z(n19816) );
  XNOR U19790 ( .A(n19815), .B(n19819), .Z(n19817) );
  XNOR U19791 ( .A(n19775), .B(n19782), .Z(n19796) );
  NOR U19792 ( .A(n19741), .B(n19820), .Z(n19782) );
  XOR U19793 ( .A(n19787), .B(n19786), .Z(n19775) );
  XNOR U19794 ( .A(n19821), .B(n19783), .Z(n19786) );
  XOR U19795 ( .A(n19822), .B(n19823), .Z(n19783) );
  AND U19796 ( .A(n19824), .B(n19825), .Z(n19823) );
  XNOR U19797 ( .A(n19826), .B(n19827), .Z(n19824) );
  IV U19798 ( .A(n19822), .Z(n19826) );
  XNOR U19799 ( .A(n19828), .B(n19829), .Z(n19821) );
  NOR U19800 ( .A(n19830), .B(n19831), .Z(n19829) );
  XNOR U19801 ( .A(n19828), .B(n19832), .Z(n19830) );
  XOR U19802 ( .A(n19833), .B(n19834), .Z(n19787) );
  NOR U19803 ( .A(n19835), .B(n19836), .Z(n19834) );
  XNOR U19804 ( .A(n19833), .B(n19837), .Z(n19835) );
  XNOR U19805 ( .A(n19725), .B(n19792), .Z(n19794) );
  XOR U19806 ( .A(n19838), .B(n19839), .Z(n19725) );
  AND U19807 ( .A(n483), .B(n19840), .Z(n19839) );
  XOR U19808 ( .A(n19841), .B(n19838), .Z(n19840) );
  AND U19809 ( .A(n19738), .B(n19741), .Z(n19792) );
  XOR U19810 ( .A(n19842), .B(n19820), .Z(n19741) );
  XNOR U19811 ( .A(p_input[1904]), .B(p_input[2048]), .Z(n19820) );
  XNOR U19812 ( .A(n19807), .B(n19806), .Z(n19842) );
  XNOR U19813 ( .A(n19843), .B(n19814), .Z(n19806) );
  XNOR U19814 ( .A(n19802), .B(n19801), .Z(n19814) );
  XNOR U19815 ( .A(n19844), .B(n19798), .Z(n19801) );
  XNOR U19816 ( .A(p_input[1914]), .B(p_input[2058]), .Z(n19798) );
  XOR U19817 ( .A(p_input[1915]), .B(n6319), .Z(n19844) );
  XOR U19818 ( .A(p_input[1916]), .B(p_input[2060]), .Z(n19802) );
  XOR U19819 ( .A(n19812), .B(n19845), .Z(n19843) );
  IV U19820 ( .A(n19803), .Z(n19845) );
  XOR U19821 ( .A(p_input[1905]), .B(p_input[2049]), .Z(n19803) );
  XNOR U19822 ( .A(n19846), .B(n19819), .Z(n19812) );
  XNOR U19823 ( .A(p_input[1919]), .B(n6322), .Z(n19819) );
  XOR U19824 ( .A(n19809), .B(n19818), .Z(n19846) );
  XOR U19825 ( .A(n19847), .B(n19815), .Z(n19818) );
  XOR U19826 ( .A(p_input[1917]), .B(p_input[2061]), .Z(n19815) );
  XOR U19827 ( .A(p_input[1918]), .B(n6324), .Z(n19847) );
  XOR U19828 ( .A(p_input[1913]), .B(p_input[2057]), .Z(n19809) );
  XOR U19829 ( .A(n19827), .B(n19825), .Z(n19807) );
  XNOR U19830 ( .A(n19848), .B(n19832), .Z(n19825) );
  XOR U19831 ( .A(p_input[1912]), .B(p_input[2056]), .Z(n19832) );
  XOR U19832 ( .A(n19822), .B(n19831), .Z(n19848) );
  XOR U19833 ( .A(n19849), .B(n19828), .Z(n19831) );
  XOR U19834 ( .A(p_input[1910]), .B(p_input[2054]), .Z(n19828) );
  XOR U19835 ( .A(p_input[1911]), .B(n7007), .Z(n19849) );
  XOR U19836 ( .A(p_input[1906]), .B(p_input[2050]), .Z(n19822) );
  XNOR U19837 ( .A(n19837), .B(n19836), .Z(n19827) );
  XOR U19838 ( .A(n19850), .B(n19833), .Z(n19836) );
  XOR U19839 ( .A(p_input[1907]), .B(p_input[2051]), .Z(n19833) );
  XOR U19840 ( .A(p_input[1908]), .B(n7009), .Z(n19850) );
  XOR U19841 ( .A(p_input[1909]), .B(p_input[2053]), .Z(n19837) );
  XOR U19842 ( .A(n19851), .B(n19852), .Z(n19738) );
  AND U19843 ( .A(n483), .B(n19853), .Z(n19852) );
  XNOR U19844 ( .A(n19854), .B(n19851), .Z(n19853) );
  XNOR U19845 ( .A(n19855), .B(n19856), .Z(n483) );
  NOR U19846 ( .A(n19857), .B(n19858), .Z(n19856) );
  XOR U19847 ( .A(n19747), .B(n19855), .Z(n19858) );
  AND U19848 ( .A(n19859), .B(n19860), .Z(n19747) );
  NOR U19849 ( .A(n19855), .B(n19746), .Z(n19857) );
  AND U19850 ( .A(n19861), .B(n19862), .Z(n19746) );
  XOR U19851 ( .A(n19863), .B(n19864), .Z(n19855) );
  AND U19852 ( .A(n19865), .B(n19866), .Z(n19864) );
  XNOR U19853 ( .A(n19863), .B(n19861), .Z(n19866) );
  IV U19854 ( .A(n19764), .Z(n19861) );
  XOR U19855 ( .A(n19867), .B(n19868), .Z(n19764) );
  XOR U19856 ( .A(n19869), .B(n19862), .Z(n19868) );
  AND U19857 ( .A(n19791), .B(n19870), .Z(n19862) );
  AND U19858 ( .A(n19871), .B(n19872), .Z(n19869) );
  XOR U19859 ( .A(n19873), .B(n19867), .Z(n19871) );
  XNOR U19860 ( .A(n19761), .B(n19863), .Z(n19865) );
  XOR U19861 ( .A(n19874), .B(n19875), .Z(n19761) );
  AND U19862 ( .A(n487), .B(n19876), .Z(n19875) );
  XOR U19863 ( .A(n19877), .B(n19874), .Z(n19876) );
  XOR U19864 ( .A(n19878), .B(n19879), .Z(n19863) );
  AND U19865 ( .A(n19880), .B(n19881), .Z(n19879) );
  XNOR U19866 ( .A(n19878), .B(n19791), .Z(n19881) );
  XOR U19867 ( .A(n19882), .B(n19872), .Z(n19791) );
  XNOR U19868 ( .A(n19883), .B(n19867), .Z(n19872) );
  XOR U19869 ( .A(n19884), .B(n19885), .Z(n19867) );
  AND U19870 ( .A(n19886), .B(n19887), .Z(n19885) );
  XOR U19871 ( .A(n19888), .B(n19884), .Z(n19886) );
  XNOR U19872 ( .A(n19889), .B(n19890), .Z(n19883) );
  AND U19873 ( .A(n19891), .B(n19892), .Z(n19890) );
  XOR U19874 ( .A(n19889), .B(n19893), .Z(n19891) );
  XNOR U19875 ( .A(n19873), .B(n19870), .Z(n19882) );
  AND U19876 ( .A(n19894), .B(n19895), .Z(n19870) );
  XOR U19877 ( .A(n19896), .B(n19897), .Z(n19873) );
  AND U19878 ( .A(n19898), .B(n19899), .Z(n19897) );
  XOR U19879 ( .A(n19896), .B(n19900), .Z(n19898) );
  XNOR U19880 ( .A(n19788), .B(n19878), .Z(n19880) );
  XOR U19881 ( .A(n19901), .B(n19902), .Z(n19788) );
  AND U19882 ( .A(n487), .B(n19903), .Z(n19902) );
  XNOR U19883 ( .A(n19904), .B(n19901), .Z(n19903) );
  XOR U19884 ( .A(n19905), .B(n19906), .Z(n19878) );
  AND U19885 ( .A(n19907), .B(n19908), .Z(n19906) );
  XNOR U19886 ( .A(n19905), .B(n19894), .Z(n19908) );
  IV U19887 ( .A(n19841), .Z(n19894) );
  XNOR U19888 ( .A(n19909), .B(n19887), .Z(n19841) );
  XNOR U19889 ( .A(n19910), .B(n19893), .Z(n19887) );
  XNOR U19890 ( .A(n19911), .B(n19912), .Z(n19893) );
  NOR U19891 ( .A(n19913), .B(n19914), .Z(n19912) );
  XOR U19892 ( .A(n19911), .B(n19915), .Z(n19913) );
  XNOR U19893 ( .A(n19892), .B(n19884), .Z(n19910) );
  XOR U19894 ( .A(n19916), .B(n19917), .Z(n19884) );
  AND U19895 ( .A(n19918), .B(n19919), .Z(n19917) );
  XOR U19896 ( .A(n19916), .B(n19920), .Z(n19918) );
  XNOR U19897 ( .A(n19921), .B(n19889), .Z(n19892) );
  XOR U19898 ( .A(n19922), .B(n19923), .Z(n19889) );
  AND U19899 ( .A(n19924), .B(n19925), .Z(n19923) );
  XNOR U19900 ( .A(n19926), .B(n19927), .Z(n19924) );
  IV U19901 ( .A(n19922), .Z(n19926) );
  XNOR U19902 ( .A(n19928), .B(n19929), .Z(n19921) );
  NOR U19903 ( .A(n19930), .B(n19931), .Z(n19929) );
  XNOR U19904 ( .A(n19928), .B(n19932), .Z(n19930) );
  XNOR U19905 ( .A(n19888), .B(n19895), .Z(n19909) );
  NOR U19906 ( .A(n19854), .B(n19933), .Z(n19895) );
  XOR U19907 ( .A(n19900), .B(n19899), .Z(n19888) );
  XNOR U19908 ( .A(n19934), .B(n19896), .Z(n19899) );
  XOR U19909 ( .A(n19935), .B(n19936), .Z(n19896) );
  AND U19910 ( .A(n19937), .B(n19938), .Z(n19936) );
  XNOR U19911 ( .A(n19939), .B(n19940), .Z(n19937) );
  IV U19912 ( .A(n19935), .Z(n19939) );
  XNOR U19913 ( .A(n19941), .B(n19942), .Z(n19934) );
  NOR U19914 ( .A(n19943), .B(n19944), .Z(n19942) );
  XNOR U19915 ( .A(n19941), .B(n19945), .Z(n19943) );
  XOR U19916 ( .A(n19946), .B(n19947), .Z(n19900) );
  NOR U19917 ( .A(n19948), .B(n19949), .Z(n19947) );
  XNOR U19918 ( .A(n19946), .B(n19950), .Z(n19948) );
  XNOR U19919 ( .A(n19838), .B(n19905), .Z(n19907) );
  XOR U19920 ( .A(n19951), .B(n19952), .Z(n19838) );
  AND U19921 ( .A(n487), .B(n19953), .Z(n19952) );
  XOR U19922 ( .A(n19954), .B(n19951), .Z(n19953) );
  AND U19923 ( .A(n19851), .B(n19854), .Z(n19905) );
  XOR U19924 ( .A(n19955), .B(n19933), .Z(n19854) );
  XNOR U19925 ( .A(p_input[1920]), .B(p_input[2048]), .Z(n19933) );
  XNOR U19926 ( .A(n19920), .B(n19919), .Z(n19955) );
  XNOR U19927 ( .A(n19956), .B(n19927), .Z(n19919) );
  XNOR U19928 ( .A(n19915), .B(n19914), .Z(n19927) );
  XNOR U19929 ( .A(n19957), .B(n19911), .Z(n19914) );
  XNOR U19930 ( .A(p_input[1930]), .B(p_input[2058]), .Z(n19911) );
  XOR U19931 ( .A(p_input[1931]), .B(n6319), .Z(n19957) );
  XOR U19932 ( .A(p_input[1932]), .B(p_input[2060]), .Z(n19915) );
  XOR U19933 ( .A(n19925), .B(n19958), .Z(n19956) );
  IV U19934 ( .A(n19916), .Z(n19958) );
  XOR U19935 ( .A(p_input[1921]), .B(p_input[2049]), .Z(n19916) );
  XNOR U19936 ( .A(n19959), .B(n19932), .Z(n19925) );
  XNOR U19937 ( .A(p_input[1935]), .B(n6322), .Z(n19932) );
  XOR U19938 ( .A(n19922), .B(n19931), .Z(n19959) );
  XOR U19939 ( .A(n19960), .B(n19928), .Z(n19931) );
  XOR U19940 ( .A(p_input[1933]), .B(p_input[2061]), .Z(n19928) );
  XOR U19941 ( .A(p_input[1934]), .B(n6324), .Z(n19960) );
  XOR U19942 ( .A(p_input[1929]), .B(p_input[2057]), .Z(n19922) );
  XOR U19943 ( .A(n19940), .B(n19938), .Z(n19920) );
  XNOR U19944 ( .A(n19961), .B(n19945), .Z(n19938) );
  XOR U19945 ( .A(p_input[1928]), .B(p_input[2056]), .Z(n19945) );
  XOR U19946 ( .A(n19935), .B(n19944), .Z(n19961) );
  XOR U19947 ( .A(n19962), .B(n19941), .Z(n19944) );
  XOR U19948 ( .A(p_input[1926]), .B(p_input[2054]), .Z(n19941) );
  XOR U19949 ( .A(p_input[1927]), .B(n7007), .Z(n19962) );
  XOR U19950 ( .A(p_input[1922]), .B(p_input[2050]), .Z(n19935) );
  XNOR U19951 ( .A(n19950), .B(n19949), .Z(n19940) );
  XOR U19952 ( .A(n19963), .B(n19946), .Z(n19949) );
  XOR U19953 ( .A(p_input[1923]), .B(p_input[2051]), .Z(n19946) );
  XOR U19954 ( .A(p_input[1924]), .B(n7009), .Z(n19963) );
  XOR U19955 ( .A(p_input[1925]), .B(p_input[2053]), .Z(n19950) );
  XOR U19956 ( .A(n19964), .B(n19965), .Z(n19851) );
  AND U19957 ( .A(n487), .B(n19966), .Z(n19965) );
  XNOR U19958 ( .A(n19967), .B(n19964), .Z(n19966) );
  XNOR U19959 ( .A(n19968), .B(n19969), .Z(n487) );
  NOR U19960 ( .A(n19970), .B(n19971), .Z(n19969) );
  XOR U19961 ( .A(n19860), .B(n19968), .Z(n19971) );
  AND U19962 ( .A(n19972), .B(n19973), .Z(n19860) );
  NOR U19963 ( .A(n19968), .B(n19859), .Z(n19970) );
  AND U19964 ( .A(n19974), .B(n19975), .Z(n19859) );
  XOR U19965 ( .A(n19976), .B(n19977), .Z(n19968) );
  AND U19966 ( .A(n19978), .B(n19979), .Z(n19977) );
  XNOR U19967 ( .A(n19976), .B(n19974), .Z(n19979) );
  IV U19968 ( .A(n19877), .Z(n19974) );
  XOR U19969 ( .A(n19980), .B(n19981), .Z(n19877) );
  XOR U19970 ( .A(n19982), .B(n19975), .Z(n19981) );
  AND U19971 ( .A(n19904), .B(n19983), .Z(n19975) );
  AND U19972 ( .A(n19984), .B(n19985), .Z(n19982) );
  XOR U19973 ( .A(n19986), .B(n19980), .Z(n19984) );
  XNOR U19974 ( .A(n19874), .B(n19976), .Z(n19978) );
  XOR U19975 ( .A(n19987), .B(n19988), .Z(n19874) );
  AND U19976 ( .A(n491), .B(n19989), .Z(n19988) );
  XOR U19977 ( .A(n19990), .B(n19987), .Z(n19989) );
  XOR U19978 ( .A(n19991), .B(n19992), .Z(n19976) );
  AND U19979 ( .A(n19993), .B(n19994), .Z(n19992) );
  XNOR U19980 ( .A(n19991), .B(n19904), .Z(n19994) );
  XOR U19981 ( .A(n19995), .B(n19985), .Z(n19904) );
  XNOR U19982 ( .A(n19996), .B(n19980), .Z(n19985) );
  XOR U19983 ( .A(n19997), .B(n19998), .Z(n19980) );
  AND U19984 ( .A(n19999), .B(n20000), .Z(n19998) );
  XOR U19985 ( .A(n20001), .B(n19997), .Z(n19999) );
  XNOR U19986 ( .A(n20002), .B(n20003), .Z(n19996) );
  AND U19987 ( .A(n20004), .B(n20005), .Z(n20003) );
  XOR U19988 ( .A(n20002), .B(n20006), .Z(n20004) );
  XNOR U19989 ( .A(n19986), .B(n19983), .Z(n19995) );
  AND U19990 ( .A(n20007), .B(n20008), .Z(n19983) );
  XOR U19991 ( .A(n20009), .B(n20010), .Z(n19986) );
  AND U19992 ( .A(n20011), .B(n20012), .Z(n20010) );
  XOR U19993 ( .A(n20009), .B(n20013), .Z(n20011) );
  XNOR U19994 ( .A(n19901), .B(n19991), .Z(n19993) );
  XOR U19995 ( .A(n20014), .B(n20015), .Z(n19901) );
  AND U19996 ( .A(n491), .B(n20016), .Z(n20015) );
  XNOR U19997 ( .A(n20017), .B(n20014), .Z(n20016) );
  XOR U19998 ( .A(n20018), .B(n20019), .Z(n19991) );
  AND U19999 ( .A(n20020), .B(n20021), .Z(n20019) );
  XNOR U20000 ( .A(n20018), .B(n20007), .Z(n20021) );
  IV U20001 ( .A(n19954), .Z(n20007) );
  XNOR U20002 ( .A(n20022), .B(n20000), .Z(n19954) );
  XNOR U20003 ( .A(n20023), .B(n20006), .Z(n20000) );
  XNOR U20004 ( .A(n20024), .B(n20025), .Z(n20006) );
  NOR U20005 ( .A(n20026), .B(n20027), .Z(n20025) );
  XOR U20006 ( .A(n20024), .B(n20028), .Z(n20026) );
  XNOR U20007 ( .A(n20005), .B(n19997), .Z(n20023) );
  XOR U20008 ( .A(n20029), .B(n20030), .Z(n19997) );
  AND U20009 ( .A(n20031), .B(n20032), .Z(n20030) );
  XOR U20010 ( .A(n20029), .B(n20033), .Z(n20031) );
  XNOR U20011 ( .A(n20034), .B(n20002), .Z(n20005) );
  XOR U20012 ( .A(n20035), .B(n20036), .Z(n20002) );
  AND U20013 ( .A(n20037), .B(n20038), .Z(n20036) );
  XNOR U20014 ( .A(n20039), .B(n20040), .Z(n20037) );
  IV U20015 ( .A(n20035), .Z(n20039) );
  XNOR U20016 ( .A(n20041), .B(n20042), .Z(n20034) );
  NOR U20017 ( .A(n20043), .B(n20044), .Z(n20042) );
  XNOR U20018 ( .A(n20041), .B(n20045), .Z(n20043) );
  XNOR U20019 ( .A(n20001), .B(n20008), .Z(n20022) );
  NOR U20020 ( .A(n19967), .B(n20046), .Z(n20008) );
  XOR U20021 ( .A(n20013), .B(n20012), .Z(n20001) );
  XNOR U20022 ( .A(n20047), .B(n20009), .Z(n20012) );
  XOR U20023 ( .A(n20048), .B(n20049), .Z(n20009) );
  AND U20024 ( .A(n20050), .B(n20051), .Z(n20049) );
  XNOR U20025 ( .A(n20052), .B(n20053), .Z(n20050) );
  IV U20026 ( .A(n20048), .Z(n20052) );
  XNOR U20027 ( .A(n20054), .B(n20055), .Z(n20047) );
  NOR U20028 ( .A(n20056), .B(n20057), .Z(n20055) );
  XNOR U20029 ( .A(n20054), .B(n20058), .Z(n20056) );
  XOR U20030 ( .A(n20059), .B(n20060), .Z(n20013) );
  NOR U20031 ( .A(n20061), .B(n20062), .Z(n20060) );
  XNOR U20032 ( .A(n20059), .B(n20063), .Z(n20061) );
  XNOR U20033 ( .A(n19951), .B(n20018), .Z(n20020) );
  XOR U20034 ( .A(n20064), .B(n20065), .Z(n19951) );
  AND U20035 ( .A(n491), .B(n20066), .Z(n20065) );
  XOR U20036 ( .A(n20067), .B(n20064), .Z(n20066) );
  AND U20037 ( .A(n19964), .B(n19967), .Z(n20018) );
  XOR U20038 ( .A(n20068), .B(n20046), .Z(n19967) );
  XNOR U20039 ( .A(p_input[1936]), .B(p_input[2048]), .Z(n20046) );
  XNOR U20040 ( .A(n20033), .B(n20032), .Z(n20068) );
  XNOR U20041 ( .A(n20069), .B(n20040), .Z(n20032) );
  XNOR U20042 ( .A(n20028), .B(n20027), .Z(n20040) );
  XNOR U20043 ( .A(n20070), .B(n20024), .Z(n20027) );
  XNOR U20044 ( .A(p_input[1946]), .B(p_input[2058]), .Z(n20024) );
  XOR U20045 ( .A(p_input[1947]), .B(n6319), .Z(n20070) );
  XOR U20046 ( .A(p_input[1948]), .B(p_input[2060]), .Z(n20028) );
  XOR U20047 ( .A(n20038), .B(n20071), .Z(n20069) );
  IV U20048 ( .A(n20029), .Z(n20071) );
  XOR U20049 ( .A(p_input[1937]), .B(p_input[2049]), .Z(n20029) );
  XNOR U20050 ( .A(n20072), .B(n20045), .Z(n20038) );
  XNOR U20051 ( .A(p_input[1951]), .B(n6322), .Z(n20045) );
  XOR U20052 ( .A(n20035), .B(n20044), .Z(n20072) );
  XOR U20053 ( .A(n20073), .B(n20041), .Z(n20044) );
  XOR U20054 ( .A(p_input[1949]), .B(p_input[2061]), .Z(n20041) );
  XOR U20055 ( .A(p_input[1950]), .B(n6324), .Z(n20073) );
  XOR U20056 ( .A(p_input[1945]), .B(p_input[2057]), .Z(n20035) );
  XOR U20057 ( .A(n20053), .B(n20051), .Z(n20033) );
  XNOR U20058 ( .A(n20074), .B(n20058), .Z(n20051) );
  XOR U20059 ( .A(p_input[1944]), .B(p_input[2056]), .Z(n20058) );
  XOR U20060 ( .A(n20048), .B(n20057), .Z(n20074) );
  XOR U20061 ( .A(n20075), .B(n20054), .Z(n20057) );
  XOR U20062 ( .A(p_input[1942]), .B(p_input[2054]), .Z(n20054) );
  XOR U20063 ( .A(p_input[1943]), .B(n7007), .Z(n20075) );
  XOR U20064 ( .A(p_input[1938]), .B(p_input[2050]), .Z(n20048) );
  XNOR U20065 ( .A(n20063), .B(n20062), .Z(n20053) );
  XOR U20066 ( .A(n20076), .B(n20059), .Z(n20062) );
  XOR U20067 ( .A(p_input[1939]), .B(p_input[2051]), .Z(n20059) );
  XOR U20068 ( .A(p_input[1940]), .B(n7009), .Z(n20076) );
  XOR U20069 ( .A(p_input[1941]), .B(p_input[2053]), .Z(n20063) );
  XOR U20070 ( .A(n20077), .B(n20078), .Z(n19964) );
  AND U20071 ( .A(n491), .B(n20079), .Z(n20078) );
  XNOR U20072 ( .A(n20080), .B(n20077), .Z(n20079) );
  XNOR U20073 ( .A(n20081), .B(n20082), .Z(n491) );
  NOR U20074 ( .A(n20083), .B(n20084), .Z(n20082) );
  XOR U20075 ( .A(n19973), .B(n20081), .Z(n20084) );
  AND U20076 ( .A(n20085), .B(n20086), .Z(n19973) );
  NOR U20077 ( .A(n20081), .B(n19972), .Z(n20083) );
  AND U20078 ( .A(n20087), .B(n20088), .Z(n19972) );
  XOR U20079 ( .A(n20089), .B(n20090), .Z(n20081) );
  AND U20080 ( .A(n20091), .B(n20092), .Z(n20090) );
  XNOR U20081 ( .A(n20089), .B(n20087), .Z(n20092) );
  IV U20082 ( .A(n19990), .Z(n20087) );
  XOR U20083 ( .A(n20093), .B(n20094), .Z(n19990) );
  XOR U20084 ( .A(n20095), .B(n20088), .Z(n20094) );
  AND U20085 ( .A(n20017), .B(n20096), .Z(n20088) );
  AND U20086 ( .A(n20097), .B(n20098), .Z(n20095) );
  XOR U20087 ( .A(n20099), .B(n20093), .Z(n20097) );
  XNOR U20088 ( .A(n19987), .B(n20089), .Z(n20091) );
  XOR U20089 ( .A(n20100), .B(n20101), .Z(n19987) );
  AND U20090 ( .A(n495), .B(n20102), .Z(n20101) );
  XOR U20091 ( .A(n20103), .B(n20100), .Z(n20102) );
  XOR U20092 ( .A(n20104), .B(n20105), .Z(n20089) );
  AND U20093 ( .A(n20106), .B(n20107), .Z(n20105) );
  XNOR U20094 ( .A(n20104), .B(n20017), .Z(n20107) );
  XOR U20095 ( .A(n20108), .B(n20098), .Z(n20017) );
  XNOR U20096 ( .A(n20109), .B(n20093), .Z(n20098) );
  XOR U20097 ( .A(n20110), .B(n20111), .Z(n20093) );
  AND U20098 ( .A(n20112), .B(n20113), .Z(n20111) );
  XOR U20099 ( .A(n20114), .B(n20110), .Z(n20112) );
  XNOR U20100 ( .A(n20115), .B(n20116), .Z(n20109) );
  AND U20101 ( .A(n20117), .B(n20118), .Z(n20116) );
  XOR U20102 ( .A(n20115), .B(n20119), .Z(n20117) );
  XNOR U20103 ( .A(n20099), .B(n20096), .Z(n20108) );
  AND U20104 ( .A(n20120), .B(n20121), .Z(n20096) );
  XOR U20105 ( .A(n20122), .B(n20123), .Z(n20099) );
  AND U20106 ( .A(n20124), .B(n20125), .Z(n20123) );
  XOR U20107 ( .A(n20122), .B(n20126), .Z(n20124) );
  XNOR U20108 ( .A(n20014), .B(n20104), .Z(n20106) );
  XOR U20109 ( .A(n20127), .B(n20128), .Z(n20014) );
  AND U20110 ( .A(n495), .B(n20129), .Z(n20128) );
  XNOR U20111 ( .A(n20130), .B(n20127), .Z(n20129) );
  XOR U20112 ( .A(n20131), .B(n20132), .Z(n20104) );
  AND U20113 ( .A(n20133), .B(n20134), .Z(n20132) );
  XNOR U20114 ( .A(n20131), .B(n20120), .Z(n20134) );
  IV U20115 ( .A(n20067), .Z(n20120) );
  XNOR U20116 ( .A(n20135), .B(n20113), .Z(n20067) );
  XNOR U20117 ( .A(n20136), .B(n20119), .Z(n20113) );
  XNOR U20118 ( .A(n20137), .B(n20138), .Z(n20119) );
  NOR U20119 ( .A(n20139), .B(n20140), .Z(n20138) );
  XOR U20120 ( .A(n20137), .B(n20141), .Z(n20139) );
  XNOR U20121 ( .A(n20118), .B(n20110), .Z(n20136) );
  XOR U20122 ( .A(n20142), .B(n20143), .Z(n20110) );
  AND U20123 ( .A(n20144), .B(n20145), .Z(n20143) );
  XOR U20124 ( .A(n20142), .B(n20146), .Z(n20144) );
  XNOR U20125 ( .A(n20147), .B(n20115), .Z(n20118) );
  XOR U20126 ( .A(n20148), .B(n20149), .Z(n20115) );
  AND U20127 ( .A(n20150), .B(n20151), .Z(n20149) );
  XNOR U20128 ( .A(n20152), .B(n20153), .Z(n20150) );
  IV U20129 ( .A(n20148), .Z(n20152) );
  XNOR U20130 ( .A(n20154), .B(n20155), .Z(n20147) );
  NOR U20131 ( .A(n20156), .B(n20157), .Z(n20155) );
  XNOR U20132 ( .A(n20154), .B(n20158), .Z(n20156) );
  XNOR U20133 ( .A(n20114), .B(n20121), .Z(n20135) );
  NOR U20134 ( .A(n20080), .B(n20159), .Z(n20121) );
  XOR U20135 ( .A(n20126), .B(n20125), .Z(n20114) );
  XNOR U20136 ( .A(n20160), .B(n20122), .Z(n20125) );
  XOR U20137 ( .A(n20161), .B(n20162), .Z(n20122) );
  AND U20138 ( .A(n20163), .B(n20164), .Z(n20162) );
  XNOR U20139 ( .A(n20165), .B(n20166), .Z(n20163) );
  IV U20140 ( .A(n20161), .Z(n20165) );
  XNOR U20141 ( .A(n20167), .B(n20168), .Z(n20160) );
  NOR U20142 ( .A(n20169), .B(n20170), .Z(n20168) );
  XNOR U20143 ( .A(n20167), .B(n20171), .Z(n20169) );
  XOR U20144 ( .A(n20172), .B(n20173), .Z(n20126) );
  NOR U20145 ( .A(n20174), .B(n20175), .Z(n20173) );
  XNOR U20146 ( .A(n20172), .B(n20176), .Z(n20174) );
  XNOR U20147 ( .A(n20064), .B(n20131), .Z(n20133) );
  XOR U20148 ( .A(n20177), .B(n20178), .Z(n20064) );
  AND U20149 ( .A(n495), .B(n20179), .Z(n20178) );
  XOR U20150 ( .A(n20180), .B(n20177), .Z(n20179) );
  AND U20151 ( .A(n20077), .B(n20080), .Z(n20131) );
  XOR U20152 ( .A(n20181), .B(n20159), .Z(n20080) );
  XNOR U20153 ( .A(p_input[1952]), .B(p_input[2048]), .Z(n20159) );
  XNOR U20154 ( .A(n20146), .B(n20145), .Z(n20181) );
  XNOR U20155 ( .A(n20182), .B(n20153), .Z(n20145) );
  XNOR U20156 ( .A(n20141), .B(n20140), .Z(n20153) );
  XNOR U20157 ( .A(n20183), .B(n20137), .Z(n20140) );
  XNOR U20158 ( .A(p_input[1962]), .B(p_input[2058]), .Z(n20137) );
  XOR U20159 ( .A(p_input[1963]), .B(n6319), .Z(n20183) );
  XOR U20160 ( .A(p_input[1964]), .B(p_input[2060]), .Z(n20141) );
  XOR U20161 ( .A(n20151), .B(n20184), .Z(n20182) );
  IV U20162 ( .A(n20142), .Z(n20184) );
  XOR U20163 ( .A(p_input[1953]), .B(p_input[2049]), .Z(n20142) );
  XNOR U20164 ( .A(n20185), .B(n20158), .Z(n20151) );
  XNOR U20165 ( .A(p_input[1967]), .B(n6322), .Z(n20158) );
  XOR U20166 ( .A(n20148), .B(n20157), .Z(n20185) );
  XOR U20167 ( .A(n20186), .B(n20154), .Z(n20157) );
  XOR U20168 ( .A(p_input[1965]), .B(p_input[2061]), .Z(n20154) );
  XOR U20169 ( .A(p_input[1966]), .B(n6324), .Z(n20186) );
  XOR U20170 ( .A(p_input[1961]), .B(p_input[2057]), .Z(n20148) );
  XOR U20171 ( .A(n20166), .B(n20164), .Z(n20146) );
  XNOR U20172 ( .A(n20187), .B(n20171), .Z(n20164) );
  XOR U20173 ( .A(p_input[1960]), .B(p_input[2056]), .Z(n20171) );
  XOR U20174 ( .A(n20161), .B(n20170), .Z(n20187) );
  XOR U20175 ( .A(n20188), .B(n20167), .Z(n20170) );
  XOR U20176 ( .A(p_input[1958]), .B(p_input[2054]), .Z(n20167) );
  XOR U20177 ( .A(p_input[1959]), .B(n7007), .Z(n20188) );
  XOR U20178 ( .A(p_input[1954]), .B(p_input[2050]), .Z(n20161) );
  XNOR U20179 ( .A(n20176), .B(n20175), .Z(n20166) );
  XOR U20180 ( .A(n20189), .B(n20172), .Z(n20175) );
  XOR U20181 ( .A(p_input[1955]), .B(p_input[2051]), .Z(n20172) );
  XOR U20182 ( .A(p_input[1956]), .B(n7009), .Z(n20189) );
  XOR U20183 ( .A(p_input[1957]), .B(p_input[2053]), .Z(n20176) );
  XOR U20184 ( .A(n20190), .B(n20191), .Z(n20077) );
  AND U20185 ( .A(n495), .B(n20192), .Z(n20191) );
  XNOR U20186 ( .A(n20193), .B(n20190), .Z(n20192) );
  XNOR U20187 ( .A(n20194), .B(n20195), .Z(n495) );
  NOR U20188 ( .A(n20196), .B(n20197), .Z(n20195) );
  XOR U20189 ( .A(n20086), .B(n20194), .Z(n20197) );
  AND U20190 ( .A(n20198), .B(n20199), .Z(n20086) );
  NOR U20191 ( .A(n20194), .B(n20085), .Z(n20196) );
  AND U20192 ( .A(n20200), .B(n20201), .Z(n20085) );
  XOR U20193 ( .A(n20202), .B(n20203), .Z(n20194) );
  AND U20194 ( .A(n20204), .B(n20205), .Z(n20203) );
  XNOR U20195 ( .A(n20202), .B(n20200), .Z(n20205) );
  IV U20196 ( .A(n20103), .Z(n20200) );
  XOR U20197 ( .A(n20206), .B(n20207), .Z(n20103) );
  XOR U20198 ( .A(n20208), .B(n20201), .Z(n20207) );
  AND U20199 ( .A(n20130), .B(n20209), .Z(n20201) );
  AND U20200 ( .A(n20210), .B(n20211), .Z(n20208) );
  XOR U20201 ( .A(n20212), .B(n20206), .Z(n20210) );
  XNOR U20202 ( .A(n20100), .B(n20202), .Z(n20204) );
  XOR U20203 ( .A(n20213), .B(n20214), .Z(n20100) );
  AND U20204 ( .A(n499), .B(n20215), .Z(n20214) );
  XOR U20205 ( .A(n20216), .B(n20213), .Z(n20215) );
  XOR U20206 ( .A(n20217), .B(n20218), .Z(n20202) );
  AND U20207 ( .A(n20219), .B(n20220), .Z(n20218) );
  XNOR U20208 ( .A(n20217), .B(n20130), .Z(n20220) );
  XOR U20209 ( .A(n20221), .B(n20211), .Z(n20130) );
  XNOR U20210 ( .A(n20222), .B(n20206), .Z(n20211) );
  XOR U20211 ( .A(n20223), .B(n20224), .Z(n20206) );
  AND U20212 ( .A(n20225), .B(n20226), .Z(n20224) );
  XOR U20213 ( .A(n20227), .B(n20223), .Z(n20225) );
  XNOR U20214 ( .A(n20228), .B(n20229), .Z(n20222) );
  AND U20215 ( .A(n20230), .B(n20231), .Z(n20229) );
  XOR U20216 ( .A(n20228), .B(n20232), .Z(n20230) );
  XNOR U20217 ( .A(n20212), .B(n20209), .Z(n20221) );
  AND U20218 ( .A(n20233), .B(n20234), .Z(n20209) );
  XOR U20219 ( .A(n20235), .B(n20236), .Z(n20212) );
  AND U20220 ( .A(n20237), .B(n20238), .Z(n20236) );
  XOR U20221 ( .A(n20235), .B(n20239), .Z(n20237) );
  XNOR U20222 ( .A(n20127), .B(n20217), .Z(n20219) );
  XOR U20223 ( .A(n20240), .B(n20241), .Z(n20127) );
  AND U20224 ( .A(n499), .B(n20242), .Z(n20241) );
  XNOR U20225 ( .A(n20243), .B(n20240), .Z(n20242) );
  XOR U20226 ( .A(n20244), .B(n20245), .Z(n20217) );
  AND U20227 ( .A(n20246), .B(n20247), .Z(n20245) );
  XNOR U20228 ( .A(n20244), .B(n20233), .Z(n20247) );
  IV U20229 ( .A(n20180), .Z(n20233) );
  XNOR U20230 ( .A(n20248), .B(n20226), .Z(n20180) );
  XNOR U20231 ( .A(n20249), .B(n20232), .Z(n20226) );
  XNOR U20232 ( .A(n20250), .B(n20251), .Z(n20232) );
  NOR U20233 ( .A(n20252), .B(n20253), .Z(n20251) );
  XOR U20234 ( .A(n20250), .B(n20254), .Z(n20252) );
  XNOR U20235 ( .A(n20231), .B(n20223), .Z(n20249) );
  XOR U20236 ( .A(n20255), .B(n20256), .Z(n20223) );
  AND U20237 ( .A(n20257), .B(n20258), .Z(n20256) );
  XOR U20238 ( .A(n20255), .B(n20259), .Z(n20257) );
  XNOR U20239 ( .A(n20260), .B(n20228), .Z(n20231) );
  XOR U20240 ( .A(n20261), .B(n20262), .Z(n20228) );
  AND U20241 ( .A(n20263), .B(n20264), .Z(n20262) );
  XNOR U20242 ( .A(n20265), .B(n20266), .Z(n20263) );
  IV U20243 ( .A(n20261), .Z(n20265) );
  XNOR U20244 ( .A(n20267), .B(n20268), .Z(n20260) );
  NOR U20245 ( .A(n20269), .B(n20270), .Z(n20268) );
  XNOR U20246 ( .A(n20267), .B(n20271), .Z(n20269) );
  XNOR U20247 ( .A(n20227), .B(n20234), .Z(n20248) );
  NOR U20248 ( .A(n20193), .B(n20272), .Z(n20234) );
  XOR U20249 ( .A(n20239), .B(n20238), .Z(n20227) );
  XNOR U20250 ( .A(n20273), .B(n20235), .Z(n20238) );
  XOR U20251 ( .A(n20274), .B(n20275), .Z(n20235) );
  AND U20252 ( .A(n20276), .B(n20277), .Z(n20275) );
  XNOR U20253 ( .A(n20278), .B(n20279), .Z(n20276) );
  IV U20254 ( .A(n20274), .Z(n20278) );
  XNOR U20255 ( .A(n20280), .B(n20281), .Z(n20273) );
  NOR U20256 ( .A(n20282), .B(n20283), .Z(n20281) );
  XNOR U20257 ( .A(n20280), .B(n20284), .Z(n20282) );
  XOR U20258 ( .A(n20285), .B(n20286), .Z(n20239) );
  NOR U20259 ( .A(n20287), .B(n20288), .Z(n20286) );
  XNOR U20260 ( .A(n20285), .B(n20289), .Z(n20287) );
  XNOR U20261 ( .A(n20177), .B(n20244), .Z(n20246) );
  XOR U20262 ( .A(n20290), .B(n20291), .Z(n20177) );
  AND U20263 ( .A(n499), .B(n20292), .Z(n20291) );
  XOR U20264 ( .A(n20293), .B(n20290), .Z(n20292) );
  AND U20265 ( .A(n20190), .B(n20193), .Z(n20244) );
  XOR U20266 ( .A(n20294), .B(n20272), .Z(n20193) );
  XNOR U20267 ( .A(p_input[1968]), .B(p_input[2048]), .Z(n20272) );
  XNOR U20268 ( .A(n20259), .B(n20258), .Z(n20294) );
  XNOR U20269 ( .A(n20295), .B(n20266), .Z(n20258) );
  XNOR U20270 ( .A(n20254), .B(n20253), .Z(n20266) );
  XNOR U20271 ( .A(n20296), .B(n20250), .Z(n20253) );
  XNOR U20272 ( .A(p_input[1978]), .B(p_input[2058]), .Z(n20250) );
  XOR U20273 ( .A(p_input[1979]), .B(n6319), .Z(n20296) );
  XOR U20274 ( .A(p_input[1980]), .B(p_input[2060]), .Z(n20254) );
  XOR U20275 ( .A(n20264), .B(n20297), .Z(n20295) );
  IV U20276 ( .A(n20255), .Z(n20297) );
  XOR U20277 ( .A(p_input[1969]), .B(p_input[2049]), .Z(n20255) );
  XNOR U20278 ( .A(n20298), .B(n20271), .Z(n20264) );
  XNOR U20279 ( .A(p_input[1983]), .B(n6322), .Z(n20271) );
  XOR U20280 ( .A(n20261), .B(n20270), .Z(n20298) );
  XOR U20281 ( .A(n20299), .B(n20267), .Z(n20270) );
  XOR U20282 ( .A(p_input[1981]), .B(p_input[2061]), .Z(n20267) );
  XOR U20283 ( .A(p_input[1982]), .B(n6324), .Z(n20299) );
  XOR U20284 ( .A(p_input[1977]), .B(p_input[2057]), .Z(n20261) );
  XOR U20285 ( .A(n20279), .B(n20277), .Z(n20259) );
  XNOR U20286 ( .A(n20300), .B(n20284), .Z(n20277) );
  XOR U20287 ( .A(p_input[1976]), .B(p_input[2056]), .Z(n20284) );
  XOR U20288 ( .A(n20274), .B(n20283), .Z(n20300) );
  XOR U20289 ( .A(n20301), .B(n20280), .Z(n20283) );
  XOR U20290 ( .A(p_input[1974]), .B(p_input[2054]), .Z(n20280) );
  XOR U20291 ( .A(p_input[1975]), .B(n7007), .Z(n20301) );
  XOR U20292 ( .A(p_input[1970]), .B(p_input[2050]), .Z(n20274) );
  XNOR U20293 ( .A(n20289), .B(n20288), .Z(n20279) );
  XOR U20294 ( .A(n20302), .B(n20285), .Z(n20288) );
  XOR U20295 ( .A(p_input[1971]), .B(p_input[2051]), .Z(n20285) );
  XOR U20296 ( .A(p_input[1972]), .B(n7009), .Z(n20302) );
  XOR U20297 ( .A(p_input[1973]), .B(p_input[2053]), .Z(n20289) );
  XOR U20298 ( .A(n20303), .B(n20304), .Z(n20190) );
  AND U20299 ( .A(n499), .B(n20305), .Z(n20304) );
  XNOR U20300 ( .A(n20306), .B(n20303), .Z(n20305) );
  XNOR U20301 ( .A(n20307), .B(n20308), .Z(n499) );
  NOR U20302 ( .A(n20309), .B(n20310), .Z(n20308) );
  XOR U20303 ( .A(n20199), .B(n20307), .Z(n20310) );
  AND U20304 ( .A(n20311), .B(n20312), .Z(n20199) );
  NOR U20305 ( .A(n20307), .B(n20198), .Z(n20309) );
  AND U20306 ( .A(n20313), .B(n20314), .Z(n20198) );
  XOR U20307 ( .A(n20315), .B(n20316), .Z(n20307) );
  AND U20308 ( .A(n20317), .B(n20318), .Z(n20316) );
  XNOR U20309 ( .A(n20315), .B(n20313), .Z(n20318) );
  IV U20310 ( .A(n20216), .Z(n20313) );
  XOR U20311 ( .A(n20319), .B(n20320), .Z(n20216) );
  XOR U20312 ( .A(n20321), .B(n20314), .Z(n20320) );
  AND U20313 ( .A(n20243), .B(n20322), .Z(n20314) );
  AND U20314 ( .A(n20323), .B(n20324), .Z(n20321) );
  XOR U20315 ( .A(n20325), .B(n20319), .Z(n20323) );
  XNOR U20316 ( .A(n20213), .B(n20315), .Z(n20317) );
  XOR U20317 ( .A(n20326), .B(n20327), .Z(n20213) );
  AND U20318 ( .A(n503), .B(n20328), .Z(n20327) );
  XOR U20319 ( .A(n20329), .B(n20326), .Z(n20328) );
  XOR U20320 ( .A(n20330), .B(n20331), .Z(n20315) );
  AND U20321 ( .A(n20332), .B(n20333), .Z(n20331) );
  XNOR U20322 ( .A(n20330), .B(n20243), .Z(n20333) );
  XOR U20323 ( .A(n20334), .B(n20324), .Z(n20243) );
  XNOR U20324 ( .A(n20335), .B(n20319), .Z(n20324) );
  XOR U20325 ( .A(n20336), .B(n20337), .Z(n20319) );
  AND U20326 ( .A(n20338), .B(n20339), .Z(n20337) );
  XOR U20327 ( .A(n20340), .B(n20336), .Z(n20338) );
  XNOR U20328 ( .A(n20341), .B(n20342), .Z(n20335) );
  AND U20329 ( .A(n20343), .B(n20344), .Z(n20342) );
  XOR U20330 ( .A(n20341), .B(n20345), .Z(n20343) );
  XNOR U20331 ( .A(n20325), .B(n20322), .Z(n20334) );
  AND U20332 ( .A(n20346), .B(n20347), .Z(n20322) );
  XOR U20333 ( .A(n20348), .B(n20349), .Z(n20325) );
  AND U20334 ( .A(n20350), .B(n20351), .Z(n20349) );
  XOR U20335 ( .A(n20348), .B(n20352), .Z(n20350) );
  XNOR U20336 ( .A(n20240), .B(n20330), .Z(n20332) );
  XOR U20337 ( .A(n20353), .B(n20354), .Z(n20240) );
  AND U20338 ( .A(n503), .B(n20355), .Z(n20354) );
  XNOR U20339 ( .A(n20356), .B(n20353), .Z(n20355) );
  XOR U20340 ( .A(n20357), .B(n20358), .Z(n20330) );
  AND U20341 ( .A(n20359), .B(n20360), .Z(n20358) );
  XNOR U20342 ( .A(n20357), .B(n20346), .Z(n20360) );
  IV U20343 ( .A(n20293), .Z(n20346) );
  XNOR U20344 ( .A(n20361), .B(n20339), .Z(n20293) );
  XNOR U20345 ( .A(n20362), .B(n20345), .Z(n20339) );
  XNOR U20346 ( .A(n20363), .B(n20364), .Z(n20345) );
  NOR U20347 ( .A(n20365), .B(n20366), .Z(n20364) );
  XOR U20348 ( .A(n20363), .B(n20367), .Z(n20365) );
  XNOR U20349 ( .A(n20344), .B(n20336), .Z(n20362) );
  XOR U20350 ( .A(n20368), .B(n20369), .Z(n20336) );
  AND U20351 ( .A(n20370), .B(n20371), .Z(n20369) );
  XOR U20352 ( .A(n20368), .B(n20372), .Z(n20370) );
  XNOR U20353 ( .A(n20373), .B(n20341), .Z(n20344) );
  XOR U20354 ( .A(n20374), .B(n20375), .Z(n20341) );
  AND U20355 ( .A(n20376), .B(n20377), .Z(n20375) );
  XNOR U20356 ( .A(n20378), .B(n20379), .Z(n20376) );
  IV U20357 ( .A(n20374), .Z(n20378) );
  XNOR U20358 ( .A(n20380), .B(n20381), .Z(n20373) );
  NOR U20359 ( .A(n20382), .B(n20383), .Z(n20381) );
  XNOR U20360 ( .A(n20380), .B(n20384), .Z(n20382) );
  XNOR U20361 ( .A(n20340), .B(n20347), .Z(n20361) );
  NOR U20362 ( .A(n20306), .B(n20385), .Z(n20347) );
  XOR U20363 ( .A(n20352), .B(n20351), .Z(n20340) );
  XNOR U20364 ( .A(n20386), .B(n20348), .Z(n20351) );
  XOR U20365 ( .A(n20387), .B(n20388), .Z(n20348) );
  AND U20366 ( .A(n20389), .B(n20390), .Z(n20388) );
  XNOR U20367 ( .A(n20391), .B(n20392), .Z(n20389) );
  IV U20368 ( .A(n20387), .Z(n20391) );
  XNOR U20369 ( .A(n20393), .B(n20394), .Z(n20386) );
  NOR U20370 ( .A(n20395), .B(n20396), .Z(n20394) );
  XNOR U20371 ( .A(n20393), .B(n20397), .Z(n20395) );
  XOR U20372 ( .A(n20398), .B(n20399), .Z(n20352) );
  NOR U20373 ( .A(n20400), .B(n20401), .Z(n20399) );
  XNOR U20374 ( .A(n20398), .B(n20402), .Z(n20400) );
  XNOR U20375 ( .A(n20290), .B(n20357), .Z(n20359) );
  XOR U20376 ( .A(n20403), .B(n20404), .Z(n20290) );
  AND U20377 ( .A(n503), .B(n20405), .Z(n20404) );
  XOR U20378 ( .A(n20406), .B(n20403), .Z(n20405) );
  AND U20379 ( .A(n20303), .B(n20306), .Z(n20357) );
  XOR U20380 ( .A(n20407), .B(n20385), .Z(n20306) );
  XNOR U20381 ( .A(p_input[1984]), .B(p_input[2048]), .Z(n20385) );
  XNOR U20382 ( .A(n20372), .B(n20371), .Z(n20407) );
  XNOR U20383 ( .A(n20408), .B(n20379), .Z(n20371) );
  XNOR U20384 ( .A(n20367), .B(n20366), .Z(n20379) );
  XNOR U20385 ( .A(n20409), .B(n20363), .Z(n20366) );
  XNOR U20386 ( .A(p_input[1994]), .B(p_input[2058]), .Z(n20363) );
  XOR U20387 ( .A(p_input[1995]), .B(n6319), .Z(n20409) );
  XOR U20388 ( .A(p_input[1996]), .B(p_input[2060]), .Z(n20367) );
  XOR U20389 ( .A(n20377), .B(n20410), .Z(n20408) );
  IV U20390 ( .A(n20368), .Z(n20410) );
  XOR U20391 ( .A(p_input[1985]), .B(p_input[2049]), .Z(n20368) );
  XNOR U20392 ( .A(n20411), .B(n20384), .Z(n20377) );
  XNOR U20393 ( .A(p_input[1999]), .B(n6322), .Z(n20384) );
  XOR U20394 ( .A(n20374), .B(n20383), .Z(n20411) );
  XOR U20395 ( .A(n20412), .B(n20380), .Z(n20383) );
  XOR U20396 ( .A(p_input[1997]), .B(p_input[2061]), .Z(n20380) );
  XOR U20397 ( .A(p_input[1998]), .B(n6324), .Z(n20412) );
  XOR U20398 ( .A(p_input[1993]), .B(p_input[2057]), .Z(n20374) );
  XOR U20399 ( .A(n20392), .B(n20390), .Z(n20372) );
  XNOR U20400 ( .A(n20413), .B(n20397), .Z(n20390) );
  XOR U20401 ( .A(p_input[1992]), .B(p_input[2056]), .Z(n20397) );
  XOR U20402 ( .A(n20387), .B(n20396), .Z(n20413) );
  XOR U20403 ( .A(n20414), .B(n20393), .Z(n20396) );
  XOR U20404 ( .A(p_input[1990]), .B(p_input[2054]), .Z(n20393) );
  XOR U20405 ( .A(p_input[1991]), .B(n7007), .Z(n20414) );
  XOR U20406 ( .A(p_input[1986]), .B(p_input[2050]), .Z(n20387) );
  XNOR U20407 ( .A(n20402), .B(n20401), .Z(n20392) );
  XOR U20408 ( .A(n20415), .B(n20398), .Z(n20401) );
  XOR U20409 ( .A(p_input[1987]), .B(p_input[2051]), .Z(n20398) );
  XOR U20410 ( .A(p_input[1988]), .B(n7009), .Z(n20415) );
  XOR U20411 ( .A(p_input[1989]), .B(p_input[2053]), .Z(n20402) );
  XOR U20412 ( .A(n20416), .B(n20417), .Z(n20303) );
  AND U20413 ( .A(n503), .B(n20418), .Z(n20417) );
  XNOR U20414 ( .A(n20419), .B(n20416), .Z(n20418) );
  XNOR U20415 ( .A(n20420), .B(n20421), .Z(n503) );
  NOR U20416 ( .A(n20422), .B(n20423), .Z(n20421) );
  XOR U20417 ( .A(n20312), .B(n20420), .Z(n20423) );
  AND U20418 ( .A(n20424), .B(n20425), .Z(n20312) );
  NOR U20419 ( .A(n20420), .B(n20311), .Z(n20422) );
  AND U20420 ( .A(n20426), .B(n20427), .Z(n20311) );
  XOR U20421 ( .A(n20428), .B(n20429), .Z(n20420) );
  AND U20422 ( .A(n20430), .B(n20431), .Z(n20429) );
  XNOR U20423 ( .A(n20428), .B(n20426), .Z(n20431) );
  IV U20424 ( .A(n20329), .Z(n20426) );
  XOR U20425 ( .A(n20432), .B(n20433), .Z(n20329) );
  XOR U20426 ( .A(n20434), .B(n20427), .Z(n20433) );
  AND U20427 ( .A(n20356), .B(n20435), .Z(n20427) );
  AND U20428 ( .A(n20436), .B(n20437), .Z(n20434) );
  XOR U20429 ( .A(n20438), .B(n20432), .Z(n20436) );
  XNOR U20430 ( .A(n20326), .B(n20428), .Z(n20430) );
  XNOR U20431 ( .A(n20439), .B(n20440), .Z(n20326) );
  AND U20432 ( .A(n506), .B(n20441), .Z(n20440) );
  XNOR U20433 ( .A(n20442), .B(n20439), .Z(n20441) );
  XOR U20434 ( .A(n20443), .B(n20444), .Z(n20428) );
  AND U20435 ( .A(n20445), .B(n20446), .Z(n20444) );
  XNOR U20436 ( .A(n20443), .B(n20356), .Z(n20446) );
  XOR U20437 ( .A(n20447), .B(n20437), .Z(n20356) );
  XNOR U20438 ( .A(n20448), .B(n20432), .Z(n20437) );
  XOR U20439 ( .A(n20449), .B(n20450), .Z(n20432) );
  AND U20440 ( .A(n20451), .B(n20452), .Z(n20450) );
  XOR U20441 ( .A(n20453), .B(n20449), .Z(n20451) );
  XNOR U20442 ( .A(n20454), .B(n20455), .Z(n20448) );
  AND U20443 ( .A(n20456), .B(n20457), .Z(n20455) );
  XOR U20444 ( .A(n20454), .B(n20458), .Z(n20456) );
  XNOR U20445 ( .A(n20438), .B(n20435), .Z(n20447) );
  AND U20446 ( .A(n20459), .B(n20460), .Z(n20435) );
  XOR U20447 ( .A(n20461), .B(n20462), .Z(n20438) );
  AND U20448 ( .A(n20463), .B(n20464), .Z(n20462) );
  XOR U20449 ( .A(n20461), .B(n20465), .Z(n20463) );
  XNOR U20450 ( .A(n20353), .B(n20443), .Z(n20445) );
  XNOR U20451 ( .A(n20466), .B(n20467), .Z(n20353) );
  AND U20452 ( .A(n506), .B(n20468), .Z(n20467) );
  XOR U20453 ( .A(n20469), .B(n20466), .Z(n20468) );
  XOR U20454 ( .A(n20470), .B(n20471), .Z(n20443) );
  AND U20455 ( .A(n20472), .B(n20473), .Z(n20471) );
  XNOR U20456 ( .A(n20470), .B(n20459), .Z(n20473) );
  IV U20457 ( .A(n20406), .Z(n20459) );
  XNOR U20458 ( .A(n20474), .B(n20452), .Z(n20406) );
  XNOR U20459 ( .A(n20475), .B(n20458), .Z(n20452) );
  XNOR U20460 ( .A(n20476), .B(n20477), .Z(n20458) );
  NOR U20461 ( .A(n20478), .B(n20479), .Z(n20477) );
  XOR U20462 ( .A(n20476), .B(n20480), .Z(n20478) );
  XNOR U20463 ( .A(n20457), .B(n20449), .Z(n20475) );
  XOR U20464 ( .A(n20481), .B(n20482), .Z(n20449) );
  AND U20465 ( .A(n20483), .B(n20484), .Z(n20482) );
  XOR U20466 ( .A(n20481), .B(n20485), .Z(n20483) );
  XNOR U20467 ( .A(n20486), .B(n20454), .Z(n20457) );
  XOR U20468 ( .A(n20487), .B(n20488), .Z(n20454) );
  AND U20469 ( .A(n20489), .B(n20490), .Z(n20488) );
  XNOR U20470 ( .A(n20491), .B(n20492), .Z(n20489) );
  IV U20471 ( .A(n20487), .Z(n20491) );
  XNOR U20472 ( .A(n20493), .B(n20494), .Z(n20486) );
  NOR U20473 ( .A(n20495), .B(n20496), .Z(n20494) );
  XNOR U20474 ( .A(n20493), .B(n20497), .Z(n20495) );
  XNOR U20475 ( .A(n20453), .B(n20460), .Z(n20474) );
  NOR U20476 ( .A(n20419), .B(n20498), .Z(n20460) );
  XOR U20477 ( .A(n20465), .B(n20464), .Z(n20453) );
  XNOR U20478 ( .A(n20499), .B(n20461), .Z(n20464) );
  XOR U20479 ( .A(n20500), .B(n20501), .Z(n20461) );
  AND U20480 ( .A(n20502), .B(n20503), .Z(n20501) );
  XNOR U20481 ( .A(n20504), .B(n20505), .Z(n20502) );
  IV U20482 ( .A(n20500), .Z(n20504) );
  XNOR U20483 ( .A(n20506), .B(n20507), .Z(n20499) );
  NOR U20484 ( .A(n20508), .B(n20509), .Z(n20507) );
  XNOR U20485 ( .A(n20506), .B(n20510), .Z(n20508) );
  XOR U20486 ( .A(n20511), .B(n20512), .Z(n20465) );
  NOR U20487 ( .A(n20513), .B(n20514), .Z(n20512) );
  XNOR U20488 ( .A(n20511), .B(n20515), .Z(n20513) );
  XNOR U20489 ( .A(n20403), .B(n20470), .Z(n20472) );
  XNOR U20490 ( .A(n20516), .B(n20517), .Z(n20403) );
  AND U20491 ( .A(n506), .B(n20518), .Z(n20517) );
  XNOR U20492 ( .A(n20519), .B(n20516), .Z(n20518) );
  AND U20493 ( .A(n20416), .B(n20419), .Z(n20470) );
  XOR U20494 ( .A(n20520), .B(n20498), .Z(n20419) );
  XNOR U20495 ( .A(p_input[2000]), .B(p_input[2048]), .Z(n20498) );
  XNOR U20496 ( .A(n20485), .B(n20484), .Z(n20520) );
  XNOR U20497 ( .A(n20521), .B(n20492), .Z(n20484) );
  XNOR U20498 ( .A(n20480), .B(n20479), .Z(n20492) );
  XNOR U20499 ( .A(n20522), .B(n20476), .Z(n20479) );
  XNOR U20500 ( .A(p_input[2010]), .B(p_input[2058]), .Z(n20476) );
  XOR U20501 ( .A(p_input[2011]), .B(n6319), .Z(n20522) );
  XOR U20502 ( .A(p_input[2012]), .B(p_input[2060]), .Z(n20480) );
  XOR U20503 ( .A(n20490), .B(n20523), .Z(n20521) );
  IV U20504 ( .A(n20481), .Z(n20523) );
  XOR U20505 ( .A(p_input[2001]), .B(p_input[2049]), .Z(n20481) );
  XNOR U20506 ( .A(n20524), .B(n20497), .Z(n20490) );
  XNOR U20507 ( .A(p_input[2015]), .B(n6322), .Z(n20497) );
  XOR U20508 ( .A(n20487), .B(n20496), .Z(n20524) );
  XOR U20509 ( .A(n20525), .B(n20493), .Z(n20496) );
  XOR U20510 ( .A(p_input[2013]), .B(p_input[2061]), .Z(n20493) );
  XOR U20511 ( .A(p_input[2014]), .B(n6324), .Z(n20525) );
  XOR U20512 ( .A(p_input[2009]), .B(p_input[2057]), .Z(n20487) );
  XOR U20513 ( .A(n20505), .B(n20503), .Z(n20485) );
  XNOR U20514 ( .A(n20526), .B(n20510), .Z(n20503) );
  XOR U20515 ( .A(p_input[2008]), .B(p_input[2056]), .Z(n20510) );
  XOR U20516 ( .A(n20500), .B(n20509), .Z(n20526) );
  XOR U20517 ( .A(n20527), .B(n20506), .Z(n20509) );
  XOR U20518 ( .A(p_input[2006]), .B(p_input[2054]), .Z(n20506) );
  XOR U20519 ( .A(p_input[2007]), .B(n7007), .Z(n20527) );
  XOR U20520 ( .A(p_input[2002]), .B(p_input[2050]), .Z(n20500) );
  XNOR U20521 ( .A(n20515), .B(n20514), .Z(n20505) );
  XOR U20522 ( .A(n20528), .B(n20511), .Z(n20514) );
  XOR U20523 ( .A(p_input[2003]), .B(p_input[2051]), .Z(n20511) );
  XOR U20524 ( .A(p_input[2004]), .B(n7009), .Z(n20528) );
  XOR U20525 ( .A(p_input[2005]), .B(p_input[2053]), .Z(n20515) );
  XOR U20526 ( .A(n20529), .B(n20530), .Z(n20416) );
  AND U20527 ( .A(n506), .B(n20531), .Z(n20530) );
  XNOR U20528 ( .A(n20532), .B(n20529), .Z(n20531) );
  XNOR U20529 ( .A(n20533), .B(n20534), .Z(n506) );
  NOR U20530 ( .A(n20535), .B(n20536), .Z(n20534) );
  XOR U20531 ( .A(n20425), .B(n20533), .Z(n20536) );
  AND U20532 ( .A(n20439), .B(n20537), .Z(n20425) );
  NOR U20533 ( .A(n20533), .B(n20424), .Z(n20535) );
  AND U20534 ( .A(n20538), .B(n20539), .Z(n20424) );
  XOR U20535 ( .A(n20540), .B(n20541), .Z(n20533) );
  AND U20536 ( .A(n20542), .B(n20543), .Z(n20541) );
  XNOR U20537 ( .A(n20540), .B(n20538), .Z(n20543) );
  IV U20538 ( .A(n20442), .Z(n20538) );
  XOR U20539 ( .A(n20544), .B(n20545), .Z(n20442) );
  XOR U20540 ( .A(n20546), .B(n20539), .Z(n20545) );
  AND U20541 ( .A(n20469), .B(n20547), .Z(n20539) );
  AND U20542 ( .A(n20548), .B(n20549), .Z(n20546) );
  XOR U20543 ( .A(n20550), .B(n20544), .Z(n20548) );
  XNOR U20544 ( .A(n20551), .B(n20540), .Z(n20542) );
  IV U20545 ( .A(n20439), .Z(n20551) );
  XNOR U20546 ( .A(n20552), .B(n20553), .Z(n20439) );
  XOR U20547 ( .A(n20554), .B(n20537), .Z(n20553) );
  AND U20548 ( .A(n20466), .B(n20555), .Z(n20537) );
  AND U20549 ( .A(n20556), .B(n20557), .Z(n20554) );
  XNOR U20550 ( .A(n20552), .B(n20558), .Z(n20556) );
  XOR U20551 ( .A(n20559), .B(n20560), .Z(n20540) );
  AND U20552 ( .A(n20561), .B(n20562), .Z(n20560) );
  XNOR U20553 ( .A(n20559), .B(n20469), .Z(n20562) );
  XOR U20554 ( .A(n20563), .B(n20549), .Z(n20469) );
  XNOR U20555 ( .A(n20564), .B(n20544), .Z(n20549) );
  XOR U20556 ( .A(n20565), .B(n20566), .Z(n20544) );
  AND U20557 ( .A(n20567), .B(n20568), .Z(n20566) );
  XOR U20558 ( .A(n20569), .B(n20565), .Z(n20567) );
  XNOR U20559 ( .A(n20570), .B(n20571), .Z(n20564) );
  AND U20560 ( .A(n20572), .B(n20573), .Z(n20571) );
  XOR U20561 ( .A(n20570), .B(n20574), .Z(n20572) );
  XNOR U20562 ( .A(n20550), .B(n20547), .Z(n20563) );
  AND U20563 ( .A(n20575), .B(n20576), .Z(n20547) );
  XOR U20564 ( .A(n20577), .B(n20578), .Z(n20550) );
  AND U20565 ( .A(n20579), .B(n20580), .Z(n20578) );
  XOR U20566 ( .A(n20577), .B(n20581), .Z(n20579) );
  XOR U20567 ( .A(n20466), .B(n20559), .Z(n20561) );
  XNOR U20568 ( .A(n20582), .B(n20558), .Z(n20466) );
  XNOR U20569 ( .A(n20583), .B(n20584), .Z(n20558) );
  AND U20570 ( .A(n20585), .B(n20586), .Z(n20584) );
  XOR U20571 ( .A(n20583), .B(n20587), .Z(n20585) );
  XNOR U20572 ( .A(n20557), .B(n20555), .Z(n20582) );
  AND U20573 ( .A(n20516), .B(n20588), .Z(n20555) );
  XNOR U20574 ( .A(n20589), .B(n20552), .Z(n20557) );
  XOR U20575 ( .A(n20590), .B(n20591), .Z(n20552) );
  AND U20576 ( .A(n20592), .B(n20593), .Z(n20591) );
  XOR U20577 ( .A(n20590), .B(n20594), .Z(n20592) );
  XNOR U20578 ( .A(n20595), .B(n20596), .Z(n20589) );
  AND U20579 ( .A(n20597), .B(n20598), .Z(n20596) );
  XNOR U20580 ( .A(n20595), .B(n20599), .Z(n20597) );
  XOR U20581 ( .A(n20600), .B(n20601), .Z(n20559) );
  AND U20582 ( .A(n20602), .B(n20603), .Z(n20601) );
  XNOR U20583 ( .A(n20600), .B(n20575), .Z(n20603) );
  IV U20584 ( .A(n20519), .Z(n20575) );
  XNOR U20585 ( .A(n20604), .B(n20568), .Z(n20519) );
  XNOR U20586 ( .A(n20605), .B(n20574), .Z(n20568) );
  XNOR U20587 ( .A(n20606), .B(n20607), .Z(n20574) );
  NOR U20588 ( .A(n20608), .B(n20609), .Z(n20607) );
  XOR U20589 ( .A(n20606), .B(n20610), .Z(n20608) );
  XNOR U20590 ( .A(n20573), .B(n20565), .Z(n20605) );
  XOR U20591 ( .A(n20611), .B(n20612), .Z(n20565) );
  AND U20592 ( .A(n20613), .B(n20614), .Z(n20612) );
  XOR U20593 ( .A(n20611), .B(n20615), .Z(n20613) );
  XNOR U20594 ( .A(n20616), .B(n20570), .Z(n20573) );
  XOR U20595 ( .A(n20617), .B(n20618), .Z(n20570) );
  AND U20596 ( .A(n20619), .B(n20620), .Z(n20618) );
  XNOR U20597 ( .A(n20621), .B(n20622), .Z(n20619) );
  IV U20598 ( .A(n20617), .Z(n20621) );
  XNOR U20599 ( .A(n20623), .B(n20624), .Z(n20616) );
  NOR U20600 ( .A(n20625), .B(n20626), .Z(n20624) );
  XNOR U20601 ( .A(n20623), .B(n20627), .Z(n20625) );
  XNOR U20602 ( .A(n20569), .B(n20576), .Z(n20604) );
  NOR U20603 ( .A(n20532), .B(n20628), .Z(n20576) );
  XOR U20604 ( .A(n20581), .B(n20580), .Z(n20569) );
  XNOR U20605 ( .A(n20629), .B(n20577), .Z(n20580) );
  XOR U20606 ( .A(n20630), .B(n20631), .Z(n20577) );
  AND U20607 ( .A(n20632), .B(n20633), .Z(n20631) );
  XNOR U20608 ( .A(n20634), .B(n20635), .Z(n20632) );
  IV U20609 ( .A(n20630), .Z(n20634) );
  XNOR U20610 ( .A(n20636), .B(n20637), .Z(n20629) );
  NOR U20611 ( .A(n20638), .B(n20639), .Z(n20637) );
  XNOR U20612 ( .A(n20636), .B(n20640), .Z(n20638) );
  XOR U20613 ( .A(n20641), .B(n20642), .Z(n20581) );
  NOR U20614 ( .A(n20643), .B(n20644), .Z(n20642) );
  XNOR U20615 ( .A(n20641), .B(n20645), .Z(n20643) );
  XNOR U20616 ( .A(n20646), .B(n20600), .Z(n20602) );
  IV U20617 ( .A(n20516), .Z(n20646) );
  XOR U20618 ( .A(n20647), .B(n20594), .Z(n20516) );
  XOR U20619 ( .A(n20587), .B(n20586), .Z(n20594) );
  XNOR U20620 ( .A(n20648), .B(n20583), .Z(n20586) );
  XOR U20621 ( .A(n20649), .B(n20650), .Z(n20583) );
  AND U20622 ( .A(n20651), .B(n20652), .Z(n20650) );
  XOR U20623 ( .A(n20649), .B(n20653), .Z(n20651) );
  XNOR U20624 ( .A(n20654), .B(n20655), .Z(n20648) );
  NOR U20625 ( .A(n20656), .B(n20657), .Z(n20655) );
  XNOR U20626 ( .A(n20654), .B(n20658), .Z(n20656) );
  XOR U20627 ( .A(n20659), .B(n20660), .Z(n20587) );
  NOR U20628 ( .A(n20661), .B(n20662), .Z(n20660) );
  XNOR U20629 ( .A(n20659), .B(n20663), .Z(n20661) );
  XNOR U20630 ( .A(n20593), .B(n20588), .Z(n20647) );
  AND U20631 ( .A(n20529), .B(n20664), .Z(n20588) );
  XOR U20632 ( .A(n20665), .B(n20599), .Z(n20593) );
  XNOR U20633 ( .A(n20666), .B(n20667), .Z(n20599) );
  NOR U20634 ( .A(n20668), .B(n20669), .Z(n20667) );
  XNOR U20635 ( .A(n20666), .B(n20670), .Z(n20668) );
  XNOR U20636 ( .A(n20598), .B(n20590), .Z(n20665) );
  XOR U20637 ( .A(n20671), .B(n20672), .Z(n20590) );
  AND U20638 ( .A(n20673), .B(n20674), .Z(n20672) );
  XOR U20639 ( .A(n20671), .B(n20675), .Z(n20673) );
  XNOR U20640 ( .A(n20676), .B(n20595), .Z(n20598) );
  XOR U20641 ( .A(n20677), .B(n20678), .Z(n20595) );
  AND U20642 ( .A(n20679), .B(n20680), .Z(n20678) );
  XOR U20643 ( .A(n20677), .B(n20681), .Z(n20679) );
  XNOR U20644 ( .A(n20682), .B(n20683), .Z(n20676) );
  NOR U20645 ( .A(n20684), .B(n20685), .Z(n20683) );
  XOR U20646 ( .A(n20682), .B(n20686), .Z(n20684) );
  AND U20647 ( .A(n20529), .B(n20532), .Z(n20600) );
  XOR U20648 ( .A(n20687), .B(n20628), .Z(n20532) );
  XNOR U20649 ( .A(p_input[2016]), .B(p_input[2048]), .Z(n20628) );
  XNOR U20650 ( .A(n20615), .B(n20614), .Z(n20687) );
  XNOR U20651 ( .A(n20688), .B(n20622), .Z(n20614) );
  XNOR U20652 ( .A(n20610), .B(n20609), .Z(n20622) );
  XNOR U20653 ( .A(n20689), .B(n20606), .Z(n20609) );
  XNOR U20654 ( .A(p_input[2026]), .B(p_input[2058]), .Z(n20606) );
  XOR U20655 ( .A(p_input[2027]), .B(n6319), .Z(n20689) );
  XOR U20656 ( .A(p_input[2028]), .B(p_input[2060]), .Z(n20610) );
  XOR U20657 ( .A(n20620), .B(n20690), .Z(n20688) );
  IV U20658 ( .A(n20611), .Z(n20690) );
  XOR U20659 ( .A(p_input[2017]), .B(p_input[2049]), .Z(n20611) );
  XNOR U20660 ( .A(n20691), .B(n20627), .Z(n20620) );
  XNOR U20661 ( .A(p_input[2031]), .B(n6322), .Z(n20627) );
  IV U20662 ( .A(p_input[2063]), .Z(n6322) );
  XOR U20663 ( .A(n20617), .B(n20626), .Z(n20691) );
  XOR U20664 ( .A(n20692), .B(n20623), .Z(n20626) );
  XOR U20665 ( .A(p_input[2029]), .B(p_input[2061]), .Z(n20623) );
  XOR U20666 ( .A(p_input[2030]), .B(n6324), .Z(n20692) );
  XOR U20667 ( .A(p_input[2025]), .B(p_input[2057]), .Z(n20617) );
  XOR U20668 ( .A(n20635), .B(n20633), .Z(n20615) );
  XNOR U20669 ( .A(n20693), .B(n20640), .Z(n20633) );
  XOR U20670 ( .A(p_input[2024]), .B(p_input[2056]), .Z(n20640) );
  XOR U20671 ( .A(n20630), .B(n20639), .Z(n20693) );
  XOR U20672 ( .A(n20694), .B(n20636), .Z(n20639) );
  XOR U20673 ( .A(p_input[2022]), .B(p_input[2054]), .Z(n20636) );
  XOR U20674 ( .A(p_input[2023]), .B(n7007), .Z(n20694) );
  XOR U20675 ( .A(p_input[2018]), .B(p_input[2050]), .Z(n20630) );
  XNOR U20676 ( .A(n20645), .B(n20644), .Z(n20635) );
  XOR U20677 ( .A(n20695), .B(n20641), .Z(n20644) );
  XOR U20678 ( .A(p_input[2019]), .B(p_input[2051]), .Z(n20641) );
  XOR U20679 ( .A(p_input[2020]), .B(n7009), .Z(n20695) );
  XOR U20680 ( .A(p_input[2021]), .B(p_input[2053]), .Z(n20645) );
  XOR U20681 ( .A(n20696), .B(n20675), .Z(n20529) );
  XOR U20682 ( .A(n20653), .B(n20652), .Z(n20675) );
  XNOR U20683 ( .A(n20697), .B(n20658), .Z(n20652) );
  XOR U20684 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[2056]), .Z(n20658) );
  XOR U20685 ( .A(n20649), .B(n20657), .Z(n20697) );
  XOR U20686 ( .A(n20698), .B(n20654), .Z(n20657) );
  XOR U20687 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[2054]), .Z(n20654) );
  XOR U20688 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n7007), .Z(n20698) );
  IV U20689 ( .A(p_input[2055]), .Z(n7007) );
  XNOR U20690 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n6328), .Z(n20649) );
  IV U20691 ( .A(p_input[2050]), .Z(n6328) );
  XNOR U20692 ( .A(n20663), .B(n20662), .Z(n20653) );
  XOR U20693 ( .A(n20699), .B(n20659), .Z(n20662) );
  XOR U20694 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[2051]), .Z(n20659) );
  XOR U20695 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n7009), .Z(n20699) );
  IV U20696 ( .A(p_input[2052]), .Z(n7009) );
  XOR U20697 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[2053]), .Z(n20663) );
  XNOR U20698 ( .A(n20674), .B(n20664), .Z(n20696) );
  XOR U20699 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[2048]), .Z(n20664) );
  XNOR U20700 ( .A(n20700), .B(n20681), .Z(n20674) );
  XNOR U20701 ( .A(n20670), .B(n20669), .Z(n20681) );
  XOR U20702 ( .A(n20701), .B(n20666), .Z(n20669) );
  XNOR U20703 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n6439), .Z(n20666) );
  IV U20704 ( .A(p_input[2058]), .Z(n6439) );
  XOR U20705 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n6319), .Z(n20701) );
  IV U20706 ( .A(p_input[2059]), .Z(n6319) );
  XOR U20707 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[2060]), .Z(
        n20670) );
  XNOR U20708 ( .A(n20680), .B(n20671), .Z(n20700) );
  XNOR U20709 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n6553), .Z(n20671) );
  IV U20710 ( .A(p_input[2049]), .Z(n6553) );
  XOR U20711 ( .A(n20702), .B(n20686), .Z(n20680) );
  XNOR U20712 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[2063]), .Z(
        n20686) );
  XOR U20713 ( .A(n20677), .B(n20685), .Z(n20702) );
  XOR U20714 ( .A(n20703), .B(n20682), .Z(n20685) );
  XOR U20715 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[2061]), .Z(
        n20682) );
  XOR U20716 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n6324), .Z(n20703) );
  IV U20717 ( .A(p_input[2062]), .Z(n6324) );
  XNOR U20718 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n6325), .Z(n20677) );
  IV U20719 ( .A(p_input[2057]), .Z(n6325) );
endmodule

