
module auction_BMR_N8_W32 ( p_input, o );
  input [8191:0] p_input;
  output [39:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
         n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
         n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041,
         n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
         n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057,
         n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
         n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
         n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081,
         n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
         n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097,
         n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
         n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
         n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
         n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129,
         n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
         n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
         n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153,
         n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
         n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
         n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177,
         n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185,
         n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
         n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201,
         n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
         n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217,
         n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
         n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233,
         n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241,
         n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249,
         n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257,
         n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
         n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273,
         n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
         n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289,
         n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297,
         n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305,
         n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313,
         n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321,
         n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329,
         n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337,
         n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345,
         n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353,
         n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361,
         n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369,
         n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377,
         n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385,
         n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393,
         n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401,
         n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409,
         n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417,
         n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
         n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433,
         n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441,
         n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449,
         n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457,
         n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465,
         n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473,
         n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481,
         n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489,
         n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497,
         n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505,
         n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513,
         n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521,
         n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529,
         n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537,
         n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545,
         n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553,
         n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561,
         n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569,
         n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577,
         n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585,
         n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593,
         n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601,
         n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609,
         n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617,
         n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625,
         n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633,
         n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641,
         n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649,
         n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657,
         n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665,
         n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673,
         n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681,
         n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689,
         n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697,
         n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705,
         n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713,
         n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721,
         n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729,
         n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737,
         n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745,
         n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753,
         n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761,
         n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769,
         n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777,
         n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
         n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793,
         n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801,
         n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809,
         n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817,
         n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825,
         n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833,
         n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
         n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849,
         n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
         n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865,
         n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873,
         n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
         n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889,
         n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897,
         n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905,
         n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
         n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921,
         n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929,
         n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937,
         n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945,
         n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953,
         n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961,
         n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969,
         n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977,
         n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985,
         n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993,
         n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
         n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
         n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017,
         n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025,
         n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033,
         n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041,
         n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049,
         n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057,
         n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065,
         n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073,
         n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081,
         n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089,
         n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097,
         n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105,
         n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113,
         n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121,
         n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
         n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137,
         n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145,
         n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153,
         n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161,
         n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169,
         n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177,
         n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185,
         n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193,
         n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201,
         n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209,
         n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217,
         n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225,
         n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233,
         n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241,
         n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249,
         n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257,
         n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265,
         n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273,
         n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281,
         n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289,
         n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297,
         n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305,
         n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313,
         n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321,
         n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329,
         n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337,
         n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
         n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353,
         n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
         n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369,
         n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377,
         n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385,
         n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393,
         n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401,
         n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409,
         n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
         n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425,
         n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
         n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441,
         n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449,
         n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457,
         n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465,
         n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473,
         n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481,
         n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
         n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497,
         n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
         n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513,
         n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521,
         n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529,
         n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537,
         n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545,
         n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553,
         n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
         n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569,
         n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577,
         n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585,
         n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593,
         n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601,
         n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609,
         n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617,
         n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625,
         n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
         n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641,
         n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649,
         n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657,
         n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665,
         n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673,
         n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681,
         n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689,
         n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697,
         n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
         n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713,
         n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721,
         n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729,
         n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737,
         n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745,
         n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753,
         n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761,
         n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769,
         n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
         n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785,
         n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
         n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801,
         n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809,
         n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817,
         n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825,
         n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833,
         n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841,
         n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
         n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857,
         n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865,
         n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873,
         n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881,
         n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889,
         n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897,
         n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905,
         n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913,
         n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
         n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929,
         n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
         n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945,
         n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953,
         n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961,
         n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969,
         n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977,
         n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985,
         n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993,
         n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001,
         n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009,
         n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017,
         n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025,
         n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033,
         n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041,
         n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049,
         n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057,
         n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065,
         n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073,
         n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
         n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089,
         n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097,
         n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105,
         n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113,
         n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121,
         n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129,
         n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137,
         n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145,
         n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153,
         n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161,
         n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169,
         n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177,
         n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185,
         n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193,
         n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201,
         n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209,
         n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217,
         n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225,
         n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233,
         n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241,
         n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
         n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257,
         n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265,
         n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273,
         n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281,
         n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289,
         n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297,
         n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305,
         n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313,
         n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
         n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329,
         n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337,
         n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345,
         n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353,
         n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361,
         n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369,
         n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377,
         n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385,
         n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393,
         n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401,
         n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409,
         n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417,
         n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425,
         n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433,
         n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
         n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449,
         n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457,
         n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465,
         n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473,
         n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481,
         n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489,
         n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497,
         n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505,
         n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
         n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521,
         n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529,
         n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
         n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545,
         n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553,
         n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561,
         n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
         n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577,
         n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
         n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593,
         n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601,
         n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
         n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
         n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625,
         n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633,
         n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
         n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649,
         n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657,
         n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665,
         n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673,
         n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681,
         n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689,
         n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697,
         n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705,
         n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713,
         n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721,
         n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729,
         n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737,
         n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745,
         n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753,
         n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761,
         n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769,
         n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777,
         n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785,
         n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793,
         n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801,
         n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809,
         n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817,
         n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825,
         n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833,
         n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841,
         n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849,
         n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857,
         n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865,
         n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873,
         n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881,
         n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889,
         n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897,
         n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905,
         n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913,
         n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921,
         n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929,
         n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937,
         n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945,
         n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953,
         n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961,
         n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969,
         n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977,
         n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985,
         n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993,
         n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
         n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009,
         n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017,
         n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025,
         n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033,
         n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041,
         n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049,
         n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057,
         n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065,
         n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073,
         n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081,
         n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089,
         n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097,
         n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105,
         n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113,
         n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121,
         n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129,
         n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137,
         n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145,
         n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153,
         n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161,
         n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169,
         n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177,
         n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185,
         n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193,
         n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201,
         n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209,
         n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217,
         n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225,
         n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233,
         n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241,
         n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249,
         n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257,
         n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265,
         n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273,
         n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281,
         n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289,
         n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297,
         n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305,
         n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313,
         n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321,
         n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329,
         n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337,
         n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345,
         n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353,
         n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361,
         n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369,
         n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377,
         n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385,
         n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393,
         n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401,
         n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409,
         n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417,
         n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425,
         n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
         n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441,
         n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449,
         n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457,
         n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465,
         n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473,
         n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481,
         n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489,
         n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497,
         n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505,
         n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513,
         n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521,
         n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529,
         n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537,
         n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545,
         n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553,
         n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561,
         n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569,
         n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577,
         n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585,
         n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593,
         n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601,
         n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609,
         n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617,
         n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625,
         n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633,
         n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641,
         n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649,
         n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657,
         n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665,
         n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673,
         n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681,
         n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689,
         n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697,
         n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705,
         n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713,
         n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721,
         n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729,
         n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737,
         n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745,
         n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753,
         n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761,
         n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769,
         n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777,
         n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785,
         n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793,
         n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801,
         n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809,
         n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817,
         n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825,
         n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833,
         n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841,
         n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849,
         n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857,
         n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865,
         n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873,
         n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
         n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889,
         n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897,
         n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905,
         n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913,
         n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921,
         n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929,
         n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
         n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945,
         n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953,
         n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961,
         n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969,
         n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977,
         n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985,
         n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993,
         n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001,
         n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009,
         n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017,
         n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025,
         n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033,
         n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041,
         n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049,
         n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057,
         n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065,
         n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073,
         n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081,
         n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089,
         n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097,
         n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105,
         n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113,
         n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121,
         n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129,
         n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137,
         n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145,
         n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153,
         n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161,
         n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169,
         n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177,
         n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185,
         n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193,
         n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201,
         n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209,
         n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217,
         n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225,
         n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233,
         n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
         n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249,
         n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257,
         n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265,
         n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273,
         n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281,
         n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289,
         n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297,
         n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305,
         n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
         n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321,
         n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329,
         n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337,
         n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345,
         n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353,
         n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361,
         n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369,
         n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377,
         n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
         n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393,
         n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401,
         n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409,
         n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417,
         n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425,
         n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433,
         n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441,
         n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449,
         n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
         n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465,
         n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473,
         n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481,
         n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489,
         n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497,
         n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505,
         n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513,
         n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521,
         n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
         n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537,
         n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545,
         n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
         n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561,
         n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569,
         n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577,
         n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585,
         n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593,
         n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
         n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609,
         n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617,
         n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625,
         n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633,
         n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641,
         n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649,
         n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657,
         n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665,
         n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
         n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681,
         n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689,
         n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697,
         n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705,
         n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713,
         n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721,
         n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729,
         n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737,
         n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
         n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753,
         n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761,
         n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769,
         n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777,
         n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785,
         n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793,
         n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801,
         n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809,
         n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817,
         n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825,
         n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833,
         n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841,
         n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849,
         n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857,
         n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865,
         n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873,
         n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881,
         n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889,
         n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897,
         n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905,
         n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913,
         n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921,
         n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929,
         n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937,
         n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945,
         n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953,
         n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961,
         n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969,
         n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977,
         n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985,
         n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993,
         n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001,
         n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009,
         n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017,
         n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025,
         n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033,
         n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041,
         n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049,
         n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
         n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065,
         n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073,
         n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081,
         n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
         n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097,
         n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
         n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113,
         n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121,
         n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
         n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137,
         n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145,
         n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153,
         n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
         n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169,
         n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
         n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185,
         n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193,
         n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
         n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209,
         n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217,
         n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225,
         n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233,
         n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241,
         n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249,
         n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257,
         n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265,
         n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273,
         n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281,
         n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289,
         n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297,
         n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305,
         n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313,
         n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
         n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329,
         n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337,
         n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345,
         n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353,
         n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361,
         n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369,
         n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
         n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385,
         n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
         n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401,
         n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409,
         n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417,
         n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425,
         n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433,
         n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441,
         n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449,
         n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457,
         n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465,
         n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473,
         n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481,
         n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489,
         n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497,
         n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505,
         n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513,
         n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521,
         n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529,
         n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537,
         n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545,
         n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553,
         n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561,
         n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569,
         n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577,
         n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585,
         n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593,
         n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601,
         n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609,
         n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617,
         n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625,
         n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633,
         n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641,
         n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649,
         n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657,
         n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
         n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673,
         n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
         n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689,
         n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697,
         n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705,
         n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713,
         n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721,
         n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729,
         n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737,
         n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745,
         n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753,
         n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761,
         n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769,
         n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777,
         n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785,
         n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793,
         n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801,
         n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809,
         n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817,
         n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825,
         n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833,
         n47834, n47835, n47836, n47837, n47838, n47839, n47840, n47841,
         n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849,
         n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857,
         n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865,
         n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873,
         n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881,
         n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889,
         n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897,
         n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905,
         n47906, n47907, n47908, n47909, n47910, n47911, n47912, n47913,
         n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921,
         n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929,
         n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937,
         n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945,
         n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953,
         n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961,
         n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969,
         n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977,
         n47978, n47979, n47980, n47981, n47982, n47983, n47984, n47985,
         n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993,
         n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001,
         n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009,
         n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017,
         n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025,
         n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033,
         n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041,
         n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049,
         n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48057,
         n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065,
         n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073,
         n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081,
         n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089,
         n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097,
         n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105,
         n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113,
         n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121,
         n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129,
         n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137,
         n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145,
         n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153,
         n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161,
         n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169,
         n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177,
         n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185,
         n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193,
         n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201,
         n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209,
         n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217,
         n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225,
         n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233,
         n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241,
         n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249,
         n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257,
         n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265,
         n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273,
         n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281,
         n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289,
         n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297,
         n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305,
         n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313,
         n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321,
         n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329,
         n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337,
         n48338, n48339, n48340, n48341, n48342, n48343, n48344, n48345,
         n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353,
         n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361,
         n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369,
         n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377,
         n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385,
         n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393,
         n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401,
         n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409,
         n48410, n48411, n48412, n48413, n48414, n48415, n48416, n48417,
         n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425,
         n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433,
         n48434, n48435, n48436, n48437, n48438, n48439, n48440, n48441,
         n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449,
         n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457,
         n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465,
         n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473,
         n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481,
         n48482, n48483, n48484, n48485, n48486, n48487, n48488, n48489,
         n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497,
         n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505,
         n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513,
         n48514, n48515, n48516, n48517, n48518, n48519, n48520, n48521,
         n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529,
         n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537,
         n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545,
         n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553,
         n48554, n48555, n48556, n48557, n48558, n48559, n48560, n48561,
         n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569,
         n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577,
         n48578, n48579, n48580, n48581, n48582, n48583, n48584, n48585,
         n48586, n48587, n48588, n48589, n48590, n48591, n48592, n48593,
         n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601,
         n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609,
         n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617,
         n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625,
         n48626, n48627, n48628, n48629, n48630, n48631, n48632, n48633,
         n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641,
         n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649,
         n48650, n48651, n48652, n48653, n48654, n48655, n48656, n48657,
         n48658, n48659, n48660, n48661, n48662, n48663, n48664, n48665,
         n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673,
         n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681,
         n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689,
         n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697,
         n48698, n48699, n48700, n48701, n48702, n48703, n48704, n48705,
         n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713,
         n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721,
         n48722, n48723, n48724, n48725, n48726, n48727, n48728, n48729,
         n48730, n48731, n48732, n48733, n48734, n48735, n48736, n48737,
         n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745,
         n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753,
         n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761,
         n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769,
         n48770, n48771, n48772, n48773, n48774, n48775, n48776, n48777,
         n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785,
         n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793,
         n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801,
         n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809,
         n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817,
         n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825,
         n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833,
         n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841,
         n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849,
         n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857,
         n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865,
         n48866, n48867, n48868, n48869, n48870, n48871, n48872, n48873,
         n48874, n48875, n48876, n48877, n48878, n48879, n48880, n48881,
         n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889,
         n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897,
         n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905,
         n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913,
         n48914, n48915, n48916, n48917, n48918, n48919, n48920, n48921,
         n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929,
         n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937,
         n48938, n48939, n48940, n48941, n48942, n48943, n48944, n48945,
         n48946, n48947, n48948, n48949, n48950, n48951, n48952, n48953,
         n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961,
         n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969,
         n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977,
         n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985,
         n48986, n48987, n48988, n48989, n48990, n48991, n48992, n48993,
         n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001,
         n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009,
         n49010, n49011, n49012, n49013, n49014, n49015, n49016, n49017,
         n49018, n49019, n49020, n49021, n49022, n49023, n49024, n49025,
         n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033,
         n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041,
         n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049,
         n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057,
         n49058, n49059, n49060, n49061, n49062, n49063, n49064, n49065,
         n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073,
         n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081,
         n49082, n49083, n49084, n49085, n49086, n49087, n49088, n49089,
         n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097,
         n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105,
         n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113,
         n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121,
         n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129,
         n49130, n49131, n49132, n49133, n49134, n49135, n49136, n49137,
         n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145,
         n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153,
         n49154, n49155, n49156, n49157, n49158, n49159, n49160, n49161,
         n49162, n49163, n49164, n49165, n49166, n49167, n49168, n49169,
         n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177,
         n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185,
         n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193,
         n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201,
         n49202, n49203, n49204, n49205, n49206, n49207, n49208, n49209,
         n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217,
         n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225,
         n49226, n49227, n49228, n49229, n49230, n49231, n49232, n49233,
         n49234, n49235, n49236, n49237, n49238, n49239, n49240, n49241,
         n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249,
         n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257,
         n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265,
         n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273,
         n49274, n49275, n49276, n49277, n49278, n49279, n49280, n49281,
         n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289,
         n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297,
         n49298, n49299, n49300, n49301, n49302, n49303, n49304, n49305,
         n49306, n49307, n49308, n49309, n49310, n49311, n49312, n49313,
         n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321,
         n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329,
         n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337,
         n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345,
         n49346, n49347, n49348, n49349, n49350, n49351, n49352, n49353,
         n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361,
         n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369,
         n49370, n49371, n49372, n49373, n49374, n49375, n49376, n49377,
         n49378, n49379, n49380, n49381, n49382, n49383, n49384, n49385,
         n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393,
         n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401,
         n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409,
         n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417,
         n49418, n49419, n49420, n49421, n49422, n49423, n49424, n49425,
         n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433,
         n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441,
         n49442, n49443, n49444, n49445, n49446, n49447, n49448, n49449,
         n49450, n49451, n49452, n49453, n49454, n49455, n49456, n49457,
         n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465,
         n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473,
         n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481,
         n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489,
         n49490, n49491, n49492, n49493, n49494, n49495, n49496, n49497,
         n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505,
         n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513,
         n49514, n49515, n49516, n49517, n49518, n49519, n49520, n49521,
         n49522, n49523, n49524, n49525, n49526, n49527, n49528, n49529,
         n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537,
         n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545,
         n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553,
         n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561,
         n49562, n49563, n49564, n49565, n49566, n49567, n49568, n49569,
         n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577,
         n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585,
         n49586, n49587, n49588, n49589, n49590, n49591, n49592, n49593,
         n49594, n49595, n49596, n49597, n49598, n49599, n49600, n49601,
         n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609,
         n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617,
         n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625,
         n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633,
         n49634, n49635, n49636, n49637, n49638, n49639, n49640, n49641,
         n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649,
         n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657,
         n49658, n49659, n49660, n49661, n49662, n49663, n49664, n49665,
         n49666, n49667, n49668, n49669, n49670, n49671, n49672, n49673,
         n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681,
         n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689,
         n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697,
         n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705,
         n49706, n49707, n49708, n49709, n49710, n49711, n49712, n49713,
         n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721,
         n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729,
         n49730, n49731, n49732, n49733, n49734, n49735, n49736, n49737,
         n49738, n49739, n49740, n49741, n49742, n49743, n49744, n49745,
         n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753,
         n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761,
         n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769,
         n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777,
         n49778, n49779, n49780, n49781, n49782, n49783, n49784, n49785,
         n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793,
         n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801,
         n49802, n49803, n49804, n49805, n49806, n49807, n49808, n49809,
         n49810, n49811, n49812, n49813, n49814, n49815, n49816, n49817,
         n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825,
         n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833,
         n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841,
         n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849,
         n49850, n49851, n49852, n49853, n49854, n49855, n49856, n49857,
         n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865,
         n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873,
         n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881,
         n49882, n49883, n49884, n49885, n49886, n49887, n49888, n49889,
         n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897,
         n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905,
         n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913,
         n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921,
         n49922, n49923, n49924, n49925, n49926, n49927, n49928, n49929,
         n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937,
         n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945,
         n49946, n49947, n49948, n49949, n49950, n49951, n49952, n49953,
         n49954, n49955, n49956, n49957, n49958, n49959, n49960, n49961,
         n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969,
         n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977,
         n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985,
         n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993,
         n49994, n49995, n49996, n49997, n49998, n49999, n50000, n50001,
         n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009,
         n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017,
         n50018, n50019, n50020, n50021, n50022, n50023, n50024, n50025,
         n50026, n50027, n50028, n50029, n50030, n50031, n50032, n50033,
         n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041,
         n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049,
         n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057,
         n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065,
         n50066, n50067, n50068, n50069, n50070, n50071, n50072, n50073,
         n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081,
         n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089,
         n50090, n50091, n50092, n50093, n50094, n50095, n50096, n50097,
         n50098, n50099, n50100, n50101, n50102, n50103, n50104, n50105,
         n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113,
         n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121,
         n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129,
         n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137,
         n50138, n50139, n50140, n50141, n50142, n50143, n50144, n50145,
         n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153,
         n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161,
         n50162, n50163, n50164, n50165, n50166, n50167, n50168, n50169,
         n50170, n50171, n50172, n50173, n50174, n50175, n50176, n50177,
         n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185,
         n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193,
         n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201,
         n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209,
         n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50217,
         n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225,
         n50226, n50227, n50228, n50229, n50230, n50231, n50232, n50233,
         n50234, n50235, n50236, n50237, n50238, n50239, n50240, n50241,
         n50242, n50243, n50244, n50245, n50246, n50247, n50248, n50249,
         n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257,
         n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265,
         n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273,
         n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281,
         n50282, n50283, n50284, n50285, n50286, n50287, n50288, n50289,
         n50290, n50291, n50292, n50293, n50294, n50295, n50296, n50297,
         n50298, n50299, n50300, n50301, n50302, n50303, n50304, n50305,
         n50306, n50307, n50308, n50309, n50310, n50311, n50312, n50313,
         n50314, n50315, n50316, n50317, n50318, n50319, n50320, n50321,
         n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329,
         n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337,
         n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345,
         n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353,
         n50354, n50355, n50356, n50357, n50358, n50359, n50360, n50361,
         n50362, n50363, n50364, n50365, n50366, n50367, n50368, n50369,
         n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377,
         n50378, n50379, n50380, n50381, n50382, n50383, n50384, n50385,
         n50386, n50387, n50388, n50389, n50390, n50391, n50392, n50393,
         n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401,
         n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409,
         n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417,
         n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425,
         n50426, n50427, n50428, n50429, n50430, n50431, n50432, n50433,
         n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441,
         n50442, n50443, n50444, n50445, n50446, n50447, n50448, n50449,
         n50450, n50451, n50452, n50453, n50454, n50455, n50456, n50457,
         n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465,
         n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473,
         n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481,
         n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489,
         n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497,
         n50498, n50499, n50500, n50501, n50502, n50503, n50504, n50505,
         n50506, n50507, n50508, n50509, n50510, n50511, n50512, n50513,
         n50514, n50515, n50516, n50517, n50518, n50519, n50520, n50521,
         n50522, n50523, n50524, n50525, n50526, n50527, n50528, n50529,
         n50530, n50531, n50532, n50533, n50534, n50535, n50536, n50537,
         n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545,
         n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553,
         n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561,
         n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569,
         n50570, n50571, n50572, n50573, n50574, n50575, n50576, n50577,
         n50578, n50579, n50580, n50581, n50582, n50583, n50584, n50585,
         n50586, n50587, n50588, n50589, n50590, n50591, n50592, n50593,
         n50594, n50595, n50596, n50597, n50598, n50599, n50600, n50601,
         n50602, n50603, n50604, n50605, n50606, n50607, n50608, n50609,
         n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617,
         n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625,
         n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633,
         n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641,
         n50642, n50643, n50644, n50645, n50646, n50647, n50648, n50649,
         n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657,
         n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665,
         n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673,
         n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681,
         n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689,
         n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697,
         n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705,
         n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713,
         n50714, n50715, n50716, n50717, n50718, n50719, n50720, n50721,
         n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729,
         n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737,
         n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745,
         n50746, n50747, n50748, n50749, n50750, n50751, n50752, n50753,
         n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761,
         n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769,
         n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777,
         n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785,
         n50786, n50787, n50788, n50789, n50790, n50791, n50792, n50793,
         n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801,
         n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809,
         n50810, n50811, n50812, n50813, n50814, n50815, n50816, n50817,
         n50818, n50819, n50820, n50821, n50822, n50823, n50824, n50825,
         n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833,
         n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841,
         n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849,
         n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857,
         n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865,
         n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873,
         n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881,
         n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889,
         n50890, n50891, n50892, n50893, n50894, n50895, n50896, n50897,
         n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905,
         n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913,
         n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921,
         n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929,
         n50930, n50931, n50932, n50933, n50934, n50935, n50936, n50937,
         n50938, n50939, n50940, n50941, n50942, n50943, n50944, n50945,
         n50946, n50947, n50948, n50949, n50950, n50951, n50952, n50953,
         n50954, n50955, n50956, n50957, n50958, n50959, n50960, n50961,
         n50962, n50963, n50964, n50965, n50966, n50967, n50968, n50969,
         n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977,
         n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985,
         n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993,
         n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001,
         n51002, n51003, n51004, n51005, n51006, n51007, n51008, n51009,
         n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51017,
         n51018, n51019, n51020, n51021, n51022, n51023, n51024, n51025,
         n51026, n51027, n51028, n51029, n51030, n51031, n51032, n51033,
         n51034, n51035, n51036, n51037, n51038, n51039, n51040, n51041,
         n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049,
         n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057,
         n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065,
         n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073,
         n51074, n51075, n51076, n51077, n51078, n51079, n51080, n51081,
         n51082, n51083, n51084, n51085, n51086, n51087, n51088, n51089,
         n51090, n51091, n51092, n51093, n51094, n51095, n51096, n51097,
         n51098, n51099, n51100, n51101, n51102, n51103, n51104, n51105,
         n51106, n51107, n51108, n51109, n51110, n51111, n51112, n51113,
         n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121,
         n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129,
         n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137,
         n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145,
         n51146, n51147, n51148, n51149, n51150, n51151, n51152, n51153,
         n51154, n51155, n51156, n51157, n51158, n51159, n51160, n51161,
         n51162, n51163, n51164, n51165, n51166, n51167, n51168, n51169,
         n51170, n51171, n51172, n51173, n51174, n51175, n51176, n51177,
         n51178, n51179, n51180, n51181, n51182, n51183, n51184, n51185,
         n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193,
         n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201,
         n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209,
         n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217,
         n51218, n51219, n51220, n51221, n51222, n51223, n51224, n51225,
         n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233,
         n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241,
         n51242, n51243, n51244, n51245, n51246, n51247, n51248, n51249,
         n51250, n51251, n51252, n51253, n51254, n51255, n51256, n51257,
         n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265,
         n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273,
         n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281,
         n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289,
         n51290, n51291, n51292, n51293, n51294, n51295, n51296, n51297,
         n51298, n51299, n51300, n51301, n51302, n51303, n51304, n51305,
         n51306, n51307, n51308, n51309, n51310, n51311, n51312, n51313,
         n51314, n51315, n51316, n51317, n51318, n51319, n51320, n51321,
         n51322, n51323, n51324, n51325, n51326, n51327, n51328, n51329,
         n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337,
         n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345,
         n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353,
         n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361,
         n51362, n51363, n51364, n51365, n51366, n51367, n51368, n51369,
         n51370, n51371, n51372, n51373, n51374, n51375, n51376, n51377,
         n51378, n51379, n51380, n51381, n51382, n51383, n51384, n51385,
         n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393,
         n51394, n51395, n51396, n51397, n51398, n51399, n51400, n51401,
         n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409,
         n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417,
         n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425,
         n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433,
         n51434, n51435, n51436, n51437, n51438, n51439, n51440, n51441,
         n51442, n51443, n51444, n51445, n51446, n51447, n51448, n51449,
         n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457,
         n51458, n51459, n51460, n51461, n51462, n51463, n51464, n51465,
         n51466, n51467, n51468, n51469, n51470, n51471, n51472, n51473,
         n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481,
         n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489,
         n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497,
         n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505,
         n51506, n51507, n51508, n51509, n51510, n51511, n51512, n51513,
         n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521,
         n51522, n51523, n51524, n51525, n51526, n51527, n51528, n51529,
         n51530, n51531, n51532, n51533, n51534, n51535, n51536, n51537,
         n51538, n51539, n51540, n51541, n51542, n51543, n51544, n51545,
         n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553,
         n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561,
         n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569,
         n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577,
         n51578, n51579, n51580, n51581, n51582, n51583, n51584, n51585,
         n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593,
         n51594, n51595, n51596, n51597, n51598, n51599, n51600, n51601,
         n51602, n51603, n51604, n51605, n51606, n51607, n51608, n51609,
         n51610, n51611, n51612, n51613, n51614, n51615, n51616, n51617,
         n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625,
         n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633,
         n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641,
         n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649,
         n51650, n51651, n51652, n51653, n51654, n51655, n51656, n51657,
         n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665,
         n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673,
         n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681,
         n51682, n51683, n51684, n51685, n51686, n51687, n51688, n51689,
         n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697,
         n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705,
         n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713,
         n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721,
         n51722, n51723, n51724, n51725, n51726, n51727, n51728, n51729,
         n51730, n51731, n51732, n51733, n51734, n51735, n51736, n51737,
         n51738, n51739, n51740, n51741, n51742, n51743, n51744, n51745,
         n51746, n51747, n51748, n51749, n51750, n51751, n51752, n51753,
         n51754, n51755, n51756, n51757, n51758, n51759, n51760, n51761,
         n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769,
         n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777,
         n51778, n51779, n51780, n51781, n51782, n51783, n51784, n51785,
         n51786, n51787, n51788, n51789, n51790, n51791, n51792, n51793,
         n51794, n51795, n51796, n51797, n51798, n51799, n51800, n51801,
         n51802, n51803, n51804, n51805, n51806, n51807, n51808, n51809,
         n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817,
         n51818, n51819, n51820, n51821, n51822, n51823, n51824, n51825,
         n51826, n51827, n51828, n51829, n51830, n51831, n51832, n51833,
         n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841,
         n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849,
         n51850, n51851, n51852, n51853, n51854, n51855, n51856, n51857,
         n51858, n51859, n51860, n51861, n51862, n51863, n51864, n51865,
         n51866, n51867, n51868, n51869, n51870, n51871, n51872, n51873,
         n51874, n51875, n51876, n51877, n51878, n51879, n51880, n51881,
         n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889,
         n51890, n51891, n51892, n51893, n51894, n51895, n51896, n51897,
         n51898, n51899, n51900, n51901, n51902, n51903, n51904, n51905,
         n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913,
         n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921,
         n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929,
         n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937,
         n51938, n51939, n51940, n51941, n51942, n51943, n51944, n51945,
         n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953,
         n51954, n51955, n51956, n51957, n51958, n51959, n51960, n51961,
         n51962, n51963, n51964, n51965, n51966, n51967, n51968, n51969,
         n51970, n51971, n51972, n51973, n51974, n51975, n51976, n51977,
         n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985,
         n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993,
         n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001,
         n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009,
         n52010, n52011, n52012, n52013, n52014, n52015, n52016, n52017,
         n52018, n52019, n52020, n52021, n52022, n52023, n52024, n52025,
         n52026, n52027, n52028, n52029, n52030, n52031, n52032, n52033,
         n52034, n52035, n52036, n52037, n52038, n52039, n52040, n52041,
         n52042, n52043, n52044, n52045, n52046, n52047, n52048, n52049,
         n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057,
         n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065,
         n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073,
         n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081,
         n52082, n52083, n52084, n52085, n52086, n52087, n52088, n52089,
         n52090, n52091, n52092, n52093, n52094, n52095, n52096, n52097,
         n52098, n52099, n52100, n52101, n52102, n52103, n52104, n52105,
         n52106, n52107, n52108, n52109, n52110, n52111, n52112, n52113,
         n52114, n52115, n52116, n52117, n52118, n52119, n52120, n52121,
         n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129,
         n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137,
         n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145,
         n52146, n52147, n52148, n52149, n52150, n52151, n52152, n52153,
         n52154, n52155, n52156, n52157, n52158, n52159, n52160, n52161,
         n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169,
         n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177,
         n52178, n52179, n52180, n52181, n52182, n52183, n52184, n52185,
         n52186, n52187, n52188, n52189, n52190, n52191, n52192, n52193,
         n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201,
         n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209,
         n52210, n52211, n52212, n52213, n52214, n52215, n52216, n52217,
         n52218, n52219, n52220, n52221, n52222, n52223, n52224, n52225,
         n52226, n52227, n52228, n52229, n52230, n52231, n52232, n52233,
         n52234, n52235, n52236, n52237, n52238, n52239, n52240, n52241,
         n52242, n52243, n52244, n52245, n52246, n52247, n52248, n52249,
         n52250, n52251, n52252, n52253, n52254, n52255, n52256, n52257,
         n52258, n52259, n52260, n52261, n52262, n52263, n52264, n52265,
         n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273,
         n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281,
         n52282, n52283, n52284, n52285, n52286, n52287, n52288, n52289,
         n52290, n52291, n52292, n52293, n52294, n52295, n52296, n52297,
         n52298, n52299, n52300, n52301, n52302, n52303, n52304, n52305,
         n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313,
         n52314, n52315, n52316, n52317, n52318, n52319, n52320, n52321,
         n52322, n52323, n52324, n52325, n52326, n52327, n52328, n52329,
         n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337,
         n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345,
         n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353,
         n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361,
         n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369,
         n52370, n52371, n52372, n52373, n52374, n52375, n52376, n52377,
         n52378, n52379, n52380, n52381, n52382, n52383, n52384, n52385,
         n52386, n52387, n52388, n52389, n52390, n52391, n52392, n52393,
         n52394, n52395, n52396, n52397, n52398, n52399, n52400, n52401,
         n52402, n52403, n52404, n52405, n52406, n52407, n52408, n52409,
         n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417,
         n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425,
         n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433,
         n52434, n52435, n52436, n52437, n52438, n52439, n52440, n52441,
         n52442, n52443, n52444, n52445, n52446, n52447, n52448, n52449,
         n52450, n52451, n52452, n52453, n52454, n52455, n52456, n52457,
         n52458, n52459, n52460, n52461, n52462, n52463, n52464, n52465,
         n52466, n52467, n52468, n52469, n52470, n52471, n52472, n52473,
         n52474, n52475, n52476, n52477, n52478, n52479, n52480, n52481,
         n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489,
         n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497,
         n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505,
         n52506, n52507, n52508, n52509, n52510, n52511, n52512, n52513,
         n52514, n52515, n52516, n52517, n52518, n52519, n52520, n52521,
         n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529,
         n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537,
         n52538, n52539, n52540, n52541, n52542, n52543, n52544, n52545,
         n52546, n52547, n52548, n52549, n52550, n52551, n52552, n52553,
         n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561,
         n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569,
         n52570, n52571, n52572, n52573, n52574, n52575, n52576, n52577,
         n52578, n52579, n52580, n52581, n52582, n52583, n52584, n52585,
         n52586, n52587, n52588, n52589, n52590, n52591, n52592, n52593,
         n52594, n52595, n52596, n52597, n52598, n52599, n52600, n52601,
         n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609,
         n52610, n52611, n52612, n52613, n52614, n52615, n52616, n52617,
         n52618, n52619, n52620, n52621, n52622, n52623, n52624, n52625,
         n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633,
         n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641,
         n52642, n52643, n52644, n52645, n52646, n52647, n52648, n52649,
         n52650, n52651, n52652, n52653, n52654, n52655, n52656, n52657,
         n52658, n52659, n52660, n52661, n52662, n52663, n52664, n52665,
         n52666, n52667, n52668, n52669, n52670, n52671, n52672, n52673,
         n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681,
         n52682, n52683, n52684, n52685, n52686, n52687, n52688, n52689,
         n52690, n52691, n52692, n52693, n52694, n52695, n52696, n52697,
         n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705,
         n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713,
         n52714, n52715, n52716, n52717, n52718, n52719, n52720, n52721,
         n52722, n52723, n52724, n52725, n52726, n52727, n52728, n52729,
         n52730, n52731, n52732, n52733, n52734, n52735, n52736, n52737,
         n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745,
         n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753,
         n52754, n52755, n52756, n52757, n52758, n52759, n52760, n52761,
         n52762, n52763, n52764, n52765, n52766, n52767, n52768, n52769,
         n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777,
         n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785,
         n52786, n52787, n52788, n52789, n52790, n52791, n52792, n52793,
         n52794, n52795, n52796, n52797, n52798, n52799, n52800, n52801,
         n52802, n52803, n52804, n52805, n52806, n52807, n52808, n52809,
         n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817,
         n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825,
         n52826, n52827, n52828, n52829, n52830, n52831, n52832, n52833,
         n52834, n52835, n52836, n52837, n52838, n52839, n52840, n52841,
         n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849,
         n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857,
         n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865,
         n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873,
         n52874, n52875, n52876, n52877, n52878, n52879, n52880, n52881,
         n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889,
         n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897,
         n52898, n52899, n52900, n52901, n52902, n52903, n52904, n52905,
         n52906, n52907, n52908, n52909, n52910, n52911, n52912, n52913,
         n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921,
         n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929,
         n52930, n52931, n52932, n52933, n52934, n52935, n52936, n52937,
         n52938, n52939, n52940, n52941, n52942, n52943, n52944, n52945,
         n52946, n52947, n52948, n52949, n52950, n52951, n52952, n52953,
         n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961,
         n52962, n52963, n52964, n52965, n52966, n52967, n52968, n52969,
         n52970, n52971, n52972, n52973, n52974, n52975, n52976, n52977,
         n52978, n52979, n52980, n52981, n52982, n52983, n52984, n52985,
         n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993,
         n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001,
         n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009,
         n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017,
         n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025,
         n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033,
         n53034, n53035, n53036, n53037, n53038, n53039, n53040, n53041,
         n53042, n53043, n53044, n53045, n53046, n53047, n53048, n53049,
         n53050, n53051, n53052, n53053, n53054, n53055, n53056, n53057,
         n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065,
         n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073,
         n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081,
         n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089,
         n53090, n53091, n53092, n53093, n53094, n53095, n53096, n53097,
         n53098, n53099, n53100, n53101, n53102, n53103, n53104, n53105,
         n53106, n53107, n53108, n53109, n53110, n53111, n53112, n53113,
         n53114, n53115, n53116, n53117, n53118, n53119, n53120, n53121,
         n53122, n53123, n53124, n53125, n53126, n53127, n53128, n53129,
         n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137,
         n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145,
         n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153,
         n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161,
         n53162, n53163, n53164, n53165, n53166, n53167, n53168, n53169,
         n53170, n53171, n53172, n53173, n53174, n53175, n53176, n53177,
         n53178, n53179, n53180, n53181, n53182, n53183, n53184, n53185,
         n53186, n53187, n53188, n53189, n53190, n53191, n53192, n53193,
         n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201,
         n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
         n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217,
         n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225,
         n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233,
         n53234, n53235, n53236, n53237, n53238, n53239, n53240, n53241,
         n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249,
         n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257,
         n53258, n53259, n53260, n53261, n53262, n53263, n53264, n53265,
         n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273,
         n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281,
         n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289,
         n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297,
         n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305,
         n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313,
         n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321,
         n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329,
         n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337,
         n53338, n53339, n53340, n53341, n53342, n53343, n53344, n53345,
         n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353,
         n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361,
         n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369,
         n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377,
         n53378, n53379, n53380, n53381, n53382, n53383, n53384, n53385,
         n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393,
         n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401,
         n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409,
         n53410, n53411, n53412, n53413, n53414, n53415, n53416, n53417,
         n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425,
         n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433,
         n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441,
         n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449,
         n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457,
         n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465,
         n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473,
         n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481,
         n53482, n53483, n53484, n53485, n53486, n53487, n53488, n53489,
         n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497,
         n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505,
         n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513,
         n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521,
         n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529,
         n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537,
         n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545,
         n53546, n53547, n53548, n53549, n53550, n53551, n53552, n53553,
         n53554, n53555, n53556, n53557, n53558, n53559, n53560, n53561,
         n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569,
         n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577,
         n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585,
         n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593,
         n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601,
         n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609,
         n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617,
         n53618, n53619, n53620, n53621, n53622, n53623, n53624, n53625,
         n53626, n53627, n53628, n53629, n53630, n53631, n53632, n53633,
         n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641,
         n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649,
         n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657,
         n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665,
         n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673,
         n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681,
         n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689,
         n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697,
         n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705,
         n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713,
         n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721,
         n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729,
         n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737,
         n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745,
         n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753,
         n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761,
         n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769,
         n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777,
         n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785,
         n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793,
         n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801,
         n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809,
         n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817,
         n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825,
         n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833,
         n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841,
         n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849,
         n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857,
         n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865,
         n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873,
         n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881,
         n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889,
         n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897,
         n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905,
         n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913,
         n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921,
         n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929,
         n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937,
         n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945,
         n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953,
         n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961,
         n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969,
         n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977,
         n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985,
         n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993,
         n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001,
         n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009,
         n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017,
         n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025,
         n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033,
         n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041,
         n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049,
         n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057,
         n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065,
         n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073,
         n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081,
         n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089,
         n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097,
         n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105,
         n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113,
         n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121,
         n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129,
         n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137,
         n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145,
         n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153,
         n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161,
         n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169,
         n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177,
         n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185,
         n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193,
         n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201,
         n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209,
         n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217,
         n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225,
         n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233,
         n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241,
         n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249,
         n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257,
         n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265,
         n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273,
         n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281,
         n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289,
         n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297,
         n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305,
         n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313,
         n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321,
         n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329,
         n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337,
         n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345,
         n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353,
         n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361,
         n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369,
         n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377,
         n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385,
         n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393,
         n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401,
         n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409,
         n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417,
         n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425,
         n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433,
         n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441,
         n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449,
         n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457,
         n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465,
         n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473,
         n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481,
         n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489,
         n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497,
         n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505,
         n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513,
         n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521,
         n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529,
         n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537,
         n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545,
         n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553,
         n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561,
         n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569,
         n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
         n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585,
         n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593,
         n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601,
         n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609,
         n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617,
         n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625,
         n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633,
         n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641,
         n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649,
         n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657,
         n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665,
         n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673,
         n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681,
         n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689,
         n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697,
         n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705,
         n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713,
         n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721,
         n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729,
         n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737,
         n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745,
         n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753,
         n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761,
         n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769,
         n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777,
         n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785,
         n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793,
         n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801,
         n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809,
         n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817,
         n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825,
         n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833,
         n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841,
         n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849,
         n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857,
         n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865,
         n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873,
         n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881,
         n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889,
         n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897,
         n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905,
         n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913,
         n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921,
         n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929,
         n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937,
         n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945,
         n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953,
         n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961,
         n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969,
         n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977,
         n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985,
         n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993,
         n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001,
         n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009,
         n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017,
         n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025,
         n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033,
         n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041,
         n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049,
         n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057,
         n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065,
         n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073,
         n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081,
         n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089,
         n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097,
         n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105,
         n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113,
         n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121,
         n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129,
         n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137,
         n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145,
         n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153,
         n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161,
         n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169,
         n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177,
         n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185,
         n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193,
         n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201,
         n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209,
         n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217,
         n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225,
         n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233,
         n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241,
         n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249,
         n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257,
         n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265,
         n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273,
         n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281,
         n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289,
         n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297,
         n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305,
         n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313,
         n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321,
         n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329,
         n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337,
         n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345,
         n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353,
         n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361,
         n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369,
         n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377,
         n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385,
         n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393,
         n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401,
         n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409,
         n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417,
         n55418, n55419, n55420, n55421, n55422, n55423, n55424, n55425,
         n55426, n55427, n55428, n55429, n55430, n55431, n55432, n55433,
         n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441,
         n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449,
         n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457,
         n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465,
         n55466, n55467, n55468, n55469, n55470, n55471, n55472, n55473,
         n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481,
         n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489,
         n55490, n55491, n55492, n55493, n55494, n55495, n55496, n55497,
         n55498, n55499, n55500, n55501, n55502, n55503, n55504, n55505,
         n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513,
         n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521,
         n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529,
         n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537,
         n55538, n55539, n55540, n55541, n55542, n55543, n55544, n55545,
         n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553,
         n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561,
         n55562, n55563, n55564, n55565, n55566, n55567, n55568, n55569,
         n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577,
         n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585,
         n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593,
         n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601,
         n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609,
         n55610, n55611, n55612, n55613, n55614, n55615, n55616, n55617,
         n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625,
         n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633,
         n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641,
         n55642, n55643, n55644, n55645, n55646, n55647, n55648, n55649,
         n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657,
         n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665,
         n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673,
         n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681,
         n55682, n55683, n55684, n55685, n55686, n55687, n55688, n55689,
         n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697,
         n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705,
         n55706, n55707, n55708, n55709, n55710, n55711, n55712, n55713,
         n55714, n55715, n55716, n55717, n55718, n55719, n55720, n55721,
         n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729,
         n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737,
         n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745,
         n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753,
         n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761,
         n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769,
         n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777,
         n55778, n55779, n55780, n55781, n55782, n55783, n55784, n55785,
         n55786, n55787, n55788, n55789, n55790, n55791, n55792, n55793,
         n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801,
         n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809,
         n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817,
         n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825,
         n55826, n55827, n55828, n55829, n55830, n55831, n55832, n55833,
         n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841,
         n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849,
         n55850, n55851, n55852, n55853, n55854, n55855, n55856, n55857,
         n55858, n55859, n55860, n55861, n55862, n55863, n55864, n55865,
         n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873,
         n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881,
         n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889,
         n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897,
         n55898, n55899, n55900, n55901, n55902, n55903, n55904, n55905,
         n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913,
         n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921,
         n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929,
         n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937,
         n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945,
         n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953,
         n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961,
         n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969,
         n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977,
         n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985,
         n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993,
         n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001,
         n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009,
         n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017,
         n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025,
         n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033,
         n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041,
         n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049,
         n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057,
         n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065,
         n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073,
         n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081,
         n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089,
         n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097,
         n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105,
         n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113,
         n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121,
         n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129,
         n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137,
         n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145,
         n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153,
         n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161,
         n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169,
         n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177,
         n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185,
         n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193,
         n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201,
         n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209,
         n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217,
         n56218, n56219, n56220, n56221, n56222, n56223, n56224, n56225,
         n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233,
         n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241,
         n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249,
         n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257,
         n56258, n56259, n56260, n56261, n56262, n56263, n56264, n56265,
         n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273,
         n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281,
         n56282, n56283, n56284, n56285, n56286, n56287, n56288, n56289,
         n56290, n56291, n56292, n56293, n56294, n56295, n56296, n56297,
         n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305,
         n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313,
         n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321,
         n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329,
         n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337,
         n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345,
         n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353,
         n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361,
         n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369,
         n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377,
         n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385,
         n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393,
         n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401,
         n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409,
         n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417,
         n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425,
         n56426, n56427, n56428, n56429, n56430, n56431, n56432, n56433,
         n56434, n56435, n56436, n56437, n56438, n56439, n56440, n56441,
         n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449,
         n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457,
         n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465,
         n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473,
         n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481,
         n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489,
         n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497,
         n56498, n56499, n56500, n56501, n56502, n56503, n56504, n56505,
         n56506, n56507, n56508, n56509, n56510, n56511, n56512, n56513,
         n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521,
         n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529,
         n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537,
         n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545,
         n56546, n56547, n56548, n56549, n56550, n56551, n56552, n56553,
         n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561,
         n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569,
         n56570, n56571, n56572, n56573, n56574, n56575, n56576, n56577,
         n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585,
         n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593,
         n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601,
         n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609,
         n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617,
         n56618, n56619, n56620, n56621, n56622, n56623, n56624, n56625,
         n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633,
         n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641,
         n56642, n56643, n56644, n56645, n56646, n56647, n56648, n56649,
         n56650, n56651, n56652, n56653, n56654, n56655, n56656, n56657,
         n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665,
         n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673,
         n56674, n56675, n56676, n56677, n56678, n56679, n56680, n56681,
         n56682, n56683, n56684, n56685, n56686, n56687, n56688, n56689,
         n56690, n56691, n56692, n56693, n56694, n56695, n56696, n56697,
         n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705,
         n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713,
         n56714, n56715, n56716, n56717, n56718, n56719, n56720, n56721,
         n56722, n56723, n56724, n56725, n56726, n56727, n56728, n56729,
         n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737,
         n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745,
         n56746, n56747, n56748, n56749, n56750, n56751, n56752, n56753,
         n56754, n56755, n56756, n56757, n56758, n56759, n56760, n56761,
         n56762, n56763, n56764, n56765, n56766, n56767, n56768, n56769,
         n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777,
         n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785,
         n56786, n56787, n56788, n56789, n56790, n56791, n56792, n56793,
         n56794, n56795, n56796, n56797, n56798, n56799, n56800, n56801,
         n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809,
         n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817,
         n56818, n56819, n56820, n56821, n56822, n56823, n56824, n56825,
         n56826, n56827, n56828, n56829, n56830, n56831, n56832, n56833,
         n56834, n56835, n56836, n56837, n56838, n56839, n56840, n56841,
         n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849,
         n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857,
         n56858, n56859, n56860, n56861, n56862, n56863, n56864, n56865,
         n56866, n56867, n56868, n56869, n56870, n56871, n56872, n56873,
         n56874, n56875, n56876, n56877, n56878, n56879, n56880, n56881,
         n56882, n56883, n56884, n56885, n56886, n56887, n56888, n56889,
         n56890, n56891, n56892, n56893, n56894, n56895, n56896, n56897,
         n56898, n56899, n56900, n56901, n56902, n56903, n56904, n56905,
         n56906, n56907, n56908, n56909, n56910, n56911, n56912, n56913,
         n56914, n56915, n56916, n56917, n56918, n56919, n56920, n56921,
         n56922, n56923, n56924, n56925, n56926, n56927, n56928, n56929,
         n56930, n56931, n56932, n56933, n56934, n56935, n56936, n56937,
         n56938, n56939, n56940, n56941, n56942, n56943, n56944, n56945,
         n56946, n56947, n56948, n56949, n56950, n56951, n56952, n56953,
         n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961,
         n56962, n56963, n56964, n56965, n56966, n56967, n56968, n56969,
         n56970, n56971, n56972, n56973, n56974, n56975, n56976, n56977,
         n56978, n56979, n56980, n56981, n56982, n56983, n56984, n56985,
         n56986, n56987, n56988, n56989, n56990, n56991, n56992, n56993,
         n56994, n56995, n56996, n56997, n56998, n56999, n57000, n57001,
         n57002, n57003, n57004, n57005, n57006, n57007, n57008, n57009,
         n57010, n57011, n57012, n57013, n57014, n57015, n57016, n57017,
         n57018, n57019, n57020, n57021, n57022, n57023, n57024, n57025,
         n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033,
         n57034, n57035, n57036, n57037, n57038, n57039, n57040, n57041,
         n57042, n57043, n57044, n57045, n57046, n57047, n57048, n57049,
         n57050, n57051, n57052, n57053, n57054, n57055, n57056, n57057,
         n57058, n57059, n57060, n57061, n57062, n57063, n57064, n57065,
         n57066, n57067, n57068, n57069, n57070, n57071, n57072, n57073,
         n57074, n57075, n57076, n57077, n57078, n57079, n57080, n57081,
         n57082, n57083, n57084, n57085, n57086, n57087, n57088, n57089,
         n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097,
         n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105,
         n57106, n57107, n57108, n57109, n57110, n57111, n57112, n57113,
         n57114, n57115, n57116, n57117, n57118, n57119, n57120, n57121,
         n57122, n57123, n57124, n57125, n57126, n57127, n57128, n57129,
         n57130, n57131, n57132, n57133, n57134, n57135, n57136, n57137,
         n57138, n57139, n57140, n57141, n57142, n57143, n57144, n57145,
         n57146, n57147, n57148, n57149, n57150, n57151, n57152, n57153,
         n57154, n57155, n57156, n57157, n57158, n57159, n57160, n57161,
         n57162, n57163, n57164, n57165, n57166, n57167, n57168, n57169,
         n57170, n57171, n57172, n57173, n57174, n57175, n57176, n57177,
         n57178, n57179, n57180, n57181, n57182, n57183, n57184, n57185,
         n57186, n57187, n57188, n57189, n57190, n57191, n57192, n57193,
         n57194, n57195, n57196, n57197, n57198, n57199, n57200, n57201,
         n57202, n57203, n57204, n57205, n57206, n57207, n57208, n57209,
         n57210, n57211, n57212, n57213, n57214, n57215, n57216, n57217,
         n57218, n57219, n57220, n57221, n57222, n57223, n57224, n57225,
         n57226, n57227, n57228, n57229, n57230, n57231, n57232, n57233,
         n57234, n57235, n57236, n57237, n57238, n57239, n57240, n57241,
         n57242, n57243, n57244, n57245, n57246, n57247, n57248, n57249,
         n57250, n57251, n57252, n57253, n57254, n57255, n57256, n57257,
         n57258, n57259, n57260, n57261, n57262, n57263, n57264, n57265,
         n57266, n57267, n57268, n57269, n57270, n57271, n57272, n57273,
         n57274, n57275, n57276, n57277, n57278, n57279, n57280, n57281,
         n57282, n57283, n57284, n57285, n57286, n57287, n57288, n57289,
         n57290, n57291, n57292, n57293, n57294, n57295, n57296, n57297,
         n57298, n57299, n57300, n57301, n57302, n57303, n57304, n57305,
         n57306, n57307, n57308, n57309, n57310, n57311, n57312, n57313,
         n57314, n57315, n57316, n57317, n57318, n57319, n57320, n57321,
         n57322, n57323, n57324, n57325, n57326, n57327, n57328, n57329,
         n57330, n57331, n57332, n57333, n57334, n57335, n57336, n57337,
         n57338, n57339, n57340, n57341, n57342, n57343, n57344, n57345,
         n57346, n57347, n57348, n57349, n57350, n57351, n57352, n57353,
         n57354, n57355, n57356, n57357, n57358, n57359, n57360, n57361,
         n57362, n57363, n57364, n57365, n57366, n57367, n57368, n57369,
         n57370, n57371, n57372, n57373, n57374, n57375, n57376, n57377,
         n57378, n57379, n57380, n57381, n57382, n57383, n57384, n57385,
         n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393,
         n57394, n57395, n57396, n57397, n57398, n57399, n57400, n57401,
         n57402, n57403, n57404, n57405, n57406, n57407, n57408, n57409,
         n57410, n57411, n57412, n57413, n57414, n57415, n57416, n57417,
         n57418, n57419, n57420, n57421, n57422, n57423, n57424, n57425,
         n57426, n57427, n57428, n57429, n57430, n57431, n57432, n57433,
         n57434, n57435, n57436, n57437, n57438, n57439, n57440, n57441,
         n57442, n57443, n57444, n57445, n57446, n57447, n57448, n57449,
         n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457,
         n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465,
         n57466, n57467, n57468, n57469, n57470, n57471, n57472, n57473,
         n57474, n57475, n57476, n57477, n57478, n57479, n57480, n57481,
         n57482, n57483, n57484, n57485, n57486, n57487, n57488, n57489,
         n57490, n57491, n57492, n57493, n57494, n57495, n57496, n57497,
         n57498, n57499, n57500, n57501, n57502, n57503, n57504, n57505,
         n57506, n57507, n57508, n57509, n57510, n57511, n57512, n57513,
         n57514, n57515, n57516, n57517, n57518, n57519, n57520, n57521,
         n57522, n57523, n57524, n57525, n57526, n57527, n57528, n57529,
         n57530, n57531, n57532, n57533, n57534, n57535, n57536, n57537,
         n57538, n57539, n57540, n57541, n57542, n57543, n57544, n57545,
         n57546, n57547, n57548, n57549, n57550, n57551, n57552, n57553,
         n57554, n57555, n57556, n57557, n57558, n57559, n57560, n57561,
         n57562, n57563, n57564, n57565, n57566, n57567, n57568, n57569,
         n57570, n57571, n57572, n57573, n57574, n57575, n57576, n57577,
         n57578, n57579, n57580, n57581, n57582, n57583, n57584, n57585,
         n57586, n57587, n57588, n57589, n57590, n57591, n57592, n57593,
         n57594, n57595, n57596, n57597, n57598, n57599, n57600, n57601,
         n57602, n57603, n57604, n57605, n57606, n57607, n57608, n57609,
         n57610, n57611, n57612, n57613, n57614, n57615, n57616, n57617,
         n57618, n57619, n57620, n57621, n57622, n57623, n57624, n57625,
         n57626, n57627, n57628, n57629, n57630, n57631, n57632, n57633,
         n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641,
         n57642, n57643, n57644, n57645, n57646, n57647, n57648, n57649,
         n57650, n57651, n57652, n57653, n57654, n57655, n57656, n57657,
         n57658, n57659, n57660, n57661, n57662, n57663, n57664, n57665,
         n57666, n57667, n57668, n57669, n57670, n57671, n57672, n57673,
         n57674, n57675, n57676, n57677, n57678, n57679, n57680, n57681,
         n57682, n57683, n57684, n57685, n57686, n57687, n57688, n57689,
         n57690, n57691, n57692, n57693, n57694, n57695, n57696, n57697,
         n57698, n57699, n57700, n57701, n57702, n57703, n57704, n57705,
         n57706, n57707, n57708, n57709, n57710, n57711, n57712, n57713,
         n57714, n57715, n57716, n57717, n57718, n57719, n57720, n57721,
         n57722, n57723, n57724, n57725, n57726, n57727, n57728, n57729,
         n57730, n57731, n57732, n57733, n57734, n57735, n57736, n57737,
         n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745,
         n57746, n57747, n57748, n57749, n57750, n57751, n57752, n57753,
         n57754, n57755, n57756, n57757, n57758, n57759, n57760, n57761,
         n57762, n57763, n57764, n57765, n57766, n57767, n57768, n57769,
         n57770, n57771, n57772, n57773, n57774, n57775, n57776, n57777,
         n57778, n57779, n57780, n57781, n57782, n57783, n57784, n57785,
         n57786, n57787, n57788, n57789, n57790, n57791, n57792, n57793,
         n57794, n57795, n57796, n57797, n57798, n57799, n57800, n57801,
         n57802, n57803, n57804, n57805, n57806, n57807, n57808, n57809,
         n57810, n57811, n57812, n57813, n57814, n57815, n57816, n57817,
         n57818, n57819, n57820, n57821, n57822, n57823, n57824, n57825,
         n57826, n57827, n57828, n57829, n57830, n57831, n57832, n57833,
         n57834, n57835, n57836, n57837, n57838, n57839, n57840, n57841,
         n57842, n57843, n57844, n57845, n57846, n57847, n57848, n57849,
         n57850, n57851, n57852, n57853, n57854, n57855, n57856, n57857,
         n57858, n57859, n57860, n57861, n57862, n57863, n57864, n57865,
         n57866, n57867, n57868, n57869, n57870, n57871, n57872, n57873,
         n57874, n57875, n57876, n57877, n57878, n57879, n57880, n57881,
         n57882, n57883, n57884, n57885, n57886, n57887, n57888, n57889,
         n57890, n57891, n57892, n57893, n57894, n57895, n57896, n57897,
         n57898, n57899, n57900, n57901, n57902, n57903, n57904, n57905,
         n57906, n57907, n57908, n57909, n57910, n57911, n57912, n57913,
         n57914, n57915, n57916, n57917, n57918, n57919, n57920, n57921,
         n57922, n57923, n57924, n57925, n57926, n57927, n57928, n57929,
         n57930, n57931, n57932, n57933, n57934, n57935, n57936, n57937,
         n57938, n57939, n57940, n57941, n57942, n57943, n57944, n57945,
         n57946, n57947, n57948, n57949, n57950, n57951, n57952, n57953,
         n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961,
         n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969,
         n57970, n57971, n57972, n57973, n57974, n57975, n57976, n57977,
         n57978, n57979, n57980, n57981, n57982, n57983, n57984, n57985,
         n57986, n57987, n57988, n57989, n57990, n57991, n57992, n57993,
         n57994, n57995, n57996, n57997, n57998, n57999, n58000, n58001,
         n58002, n58003, n58004, n58005, n58006, n58007, n58008, n58009,
         n58010, n58011, n58012, n58013, n58014, n58015, n58016, n58017,
         n58018, n58019, n58020, n58021, n58022, n58023, n58024, n58025,
         n58026, n58027, n58028, n58029, n58030, n58031, n58032, n58033,
         n58034, n58035, n58036, n58037, n58038, n58039, n58040, n58041,
         n58042, n58043, n58044, n58045, n58046, n58047, n58048, n58049,
         n58050, n58051, n58052, n58053, n58054, n58055, n58056, n58057,
         n58058, n58059, n58060, n58061, n58062, n58063, n58064, n58065,
         n58066, n58067, n58068, n58069, n58070, n58071, n58072, n58073,
         n58074, n58075, n58076, n58077, n58078, n58079, n58080, n58081,
         n58082, n58083, n58084, n58085, n58086, n58087, n58088, n58089,
         n58090, n58091, n58092, n58093, n58094, n58095, n58096, n58097,
         n58098, n58099, n58100, n58101, n58102, n58103, n58104, n58105,
         n58106, n58107, n58108, n58109, n58110, n58111, n58112, n58113,
         n58114, n58115, n58116, n58117, n58118, n58119, n58120, n58121,
         n58122, n58123, n58124, n58125, n58126, n58127, n58128, n58129,
         n58130, n58131, n58132, n58133, n58134, n58135, n58136, n58137,
         n58138, n58139, n58140, n58141, n58142, n58143, n58144, n58145,
         n58146, n58147, n58148, n58149, n58150, n58151, n58152, n58153,
         n58154, n58155, n58156, n58157, n58158, n58159, n58160, n58161,
         n58162, n58163, n58164, n58165, n58166, n58167, n58168, n58169,
         n58170, n58171, n58172, n58173, n58174, n58175, n58176, n58177,
         n58178, n58179, n58180, n58181, n58182, n58183, n58184, n58185,
         n58186, n58187, n58188, n58189, n58190, n58191, n58192, n58193,
         n58194, n58195, n58196, n58197, n58198, n58199, n58200, n58201,
         n58202, n58203, n58204, n58205, n58206, n58207, n58208, n58209,
         n58210, n58211, n58212, n58213, n58214, n58215, n58216, n58217,
         n58218, n58219, n58220, n58221, n58222, n58223, n58224, n58225,
         n58226, n58227, n58228, n58229, n58230, n58231, n58232, n58233,
         n58234, n58235, n58236, n58237, n58238, n58239, n58240, n58241,
         n58242, n58243, n58244, n58245, n58246, n58247, n58248, n58249,
         n58250, n58251, n58252, n58253, n58254, n58255, n58256, n58257,
         n58258, n58259, n58260, n58261, n58262, n58263, n58264, n58265,
         n58266, n58267, n58268, n58269, n58270, n58271, n58272, n58273,
         n58274, n58275, n58276, n58277, n58278, n58279, n58280, n58281,
         n58282, n58283, n58284, n58285, n58286, n58287, n58288, n58289,
         n58290, n58291, n58292, n58293, n58294, n58295, n58296, n58297,
         n58298, n58299, n58300, n58301, n58302, n58303, n58304, n58305,
         n58306, n58307, n58308, n58309, n58310, n58311, n58312, n58313,
         n58314, n58315, n58316, n58317, n58318, n58319, n58320, n58321,
         n58322, n58323, n58324, n58325, n58326, n58327, n58328, n58329,
         n58330, n58331, n58332, n58333, n58334, n58335, n58336, n58337,
         n58338, n58339, n58340, n58341, n58342, n58343, n58344, n58345,
         n58346, n58347, n58348, n58349, n58350, n58351, n58352, n58353,
         n58354, n58355, n58356, n58357, n58358, n58359, n58360, n58361,
         n58362, n58363, n58364, n58365, n58366, n58367, n58368, n58369,
         n58370, n58371, n58372, n58373, n58374, n58375, n58376, n58377,
         n58378, n58379, n58380, n58381, n58382, n58383, n58384, n58385,
         n58386, n58387, n58388, n58389, n58390, n58391, n58392, n58393,
         n58394, n58395, n58396, n58397, n58398, n58399, n58400, n58401,
         n58402, n58403, n58404, n58405, n58406, n58407, n58408, n58409,
         n58410, n58411, n58412, n58413, n58414, n58415, n58416, n58417,
         n58418, n58419, n58420, n58421, n58422, n58423, n58424, n58425,
         n58426, n58427, n58428, n58429, n58430, n58431, n58432, n58433,
         n58434, n58435, n58436, n58437, n58438, n58439, n58440, n58441,
         n58442, n58443, n58444, n58445, n58446, n58447, n58448, n58449,
         n58450, n58451, n58452, n58453, n58454, n58455, n58456, n58457,
         n58458, n58459, n58460, n58461, n58462, n58463, n58464, n58465,
         n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473,
         n58474, n58475, n58476, n58477, n58478, n58479, n58480, n58481,
         n58482, n58483, n58484, n58485, n58486, n58487, n58488, n58489,
         n58490, n58491, n58492, n58493, n58494, n58495, n58496, n58497,
         n58498, n58499, n58500, n58501, n58502, n58503, n58504, n58505,
         n58506, n58507, n58508, n58509, n58510, n58511, n58512, n58513,
         n58514, n58515, n58516, n58517, n58518, n58519, n58520, n58521,
         n58522, n58523, n58524, n58525, n58526, n58527, n58528, n58529,
         n58530, n58531, n58532, n58533, n58534, n58535, n58536, n58537,
         n58538, n58539, n58540, n58541, n58542, n58543, n58544, n58545,
         n58546, n58547, n58548, n58549, n58550, n58551, n58552, n58553,
         n58554, n58555, n58556, n58557, n58558, n58559, n58560, n58561,
         n58562, n58563, n58564, n58565, n58566, n58567, n58568, n58569,
         n58570, n58571, n58572, n58573, n58574, n58575, n58576, n58577,
         n58578, n58579, n58580, n58581, n58582, n58583, n58584, n58585,
         n58586, n58587, n58588, n58589, n58590, n58591, n58592, n58593,
         n58594, n58595, n58596, n58597, n58598, n58599, n58600, n58601,
         n58602, n58603, n58604, n58605, n58606, n58607, n58608, n58609,
         n58610, n58611, n58612, n58613, n58614, n58615, n58616, n58617,
         n58618, n58619, n58620, n58621, n58622, n58623, n58624, n58625,
         n58626, n58627, n58628, n58629, n58630, n58631, n58632, n58633,
         n58634, n58635, n58636, n58637, n58638, n58639, n58640, n58641,
         n58642, n58643, n58644, n58645, n58646, n58647, n58648, n58649,
         n58650, n58651, n58652, n58653, n58654, n58655, n58656, n58657,
         n58658, n58659, n58660, n58661, n58662, n58663, n58664, n58665,
         n58666, n58667, n58668, n58669, n58670, n58671, n58672, n58673,
         n58674, n58675, n58676, n58677, n58678, n58679, n58680, n58681,
         n58682, n58683, n58684, n58685, n58686, n58687, n58688, n58689,
         n58690, n58691, n58692, n58693, n58694, n58695, n58696, n58697,
         n58698, n58699, n58700, n58701, n58702, n58703, n58704, n58705,
         n58706, n58707, n58708, n58709, n58710, n58711, n58712, n58713,
         n58714, n58715, n58716, n58717, n58718, n58719, n58720, n58721,
         n58722, n58723, n58724, n58725, n58726, n58727, n58728, n58729,
         n58730, n58731, n58732, n58733, n58734, n58735, n58736, n58737,
         n58738, n58739, n58740, n58741, n58742, n58743, n58744, n58745,
         n58746, n58747, n58748, n58749, n58750, n58751, n58752, n58753,
         n58754, n58755, n58756, n58757, n58758, n58759, n58760, n58761,
         n58762, n58763, n58764, n58765, n58766, n58767, n58768, n58769,
         n58770, n58771, n58772, n58773, n58774, n58775, n58776, n58777,
         n58778, n58779, n58780, n58781, n58782, n58783, n58784, n58785,
         n58786, n58787, n58788, n58789, n58790, n58791, n58792, n58793,
         n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58801,
         n58802, n58803, n58804, n58805, n58806, n58807, n58808, n58809,
         n58810, n58811, n58812, n58813, n58814, n58815, n58816, n58817,
         n58818, n58819, n58820, n58821, n58822, n58823, n58824, n58825,
         n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833,
         n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841,
         n58842, n58843, n58844, n58845, n58846, n58847, n58848, n58849,
         n58850, n58851, n58852, n58853, n58854, n58855, n58856, n58857,
         n58858, n58859, n58860, n58861, n58862, n58863, n58864, n58865,
         n58866, n58867, n58868, n58869, n58870, n58871, n58872, n58873,
         n58874, n58875, n58876, n58877, n58878, n58879, n58880, n58881,
         n58882, n58883, n58884, n58885, n58886, n58887, n58888, n58889,
         n58890, n58891, n58892, n58893, n58894, n58895, n58896, n58897,
         n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905,
         n58906, n58907, n58908, n58909, n58910, n58911, n58912, n58913,
         n58914, n58915, n58916, n58917, n58918, n58919, n58920, n58921,
         n58922, n58923, n58924, n58925, n58926, n58927, n58928, n58929,
         n58930, n58931, n58932, n58933, n58934, n58935, n58936, n58937,
         n58938, n58939, n58940, n58941, n58942, n58943, n58944, n58945,
         n58946, n58947, n58948, n58949, n58950, n58951, n58952, n58953,
         n58954, n58955, n58956, n58957, n58958, n58959, n58960, n58961,
         n58962, n58963, n58964, n58965, n58966, n58967, n58968, n58969,
         n58970, n58971, n58972, n58973, n58974, n58975, n58976, n58977,
         n58978, n58979, n58980, n58981, n58982, n58983, n58984, n58985,
         n58986, n58987, n58988, n58989, n58990, n58991, n58992, n58993,
         n58994, n58995, n58996, n58997, n58998, n58999, n59000, n59001,
         n59002, n59003, n59004, n59005, n59006, n59007, n59008, n59009,
         n59010, n59011, n59012, n59013, n59014, n59015, n59016, n59017,
         n59018, n59019, n59020, n59021, n59022, n59023, n59024, n59025,
         n59026, n59027, n59028, n59029, n59030, n59031, n59032, n59033,
         n59034, n59035, n59036, n59037, n59038, n59039, n59040, n59041,
         n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049,
         n59050, n59051, n59052, n59053, n59054, n59055, n59056, n59057,
         n59058, n59059, n59060, n59061, n59062, n59063, n59064, n59065,
         n59066, n59067, n59068, n59069;

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[7]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n4), .B(n5), .Z(n3) );
  XNOR U4 ( .A(n6), .B(n7), .Z(o[8]) );
  AND U5 ( .A(o[7]), .B(n8), .Z(n6) );
  XNOR U6 ( .A(n9), .B(n7), .Z(n8) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[39]) );
  AND U8 ( .A(o[7]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[38]) );
  AND U11 ( .A(o[7]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[37]) );
  AND U14 ( .A(o[7]), .B(n22), .Z(n20) );
  XOR U15 ( .A(n23), .B(n24), .Z(n22) );
  XOR U16 ( .A(n25), .B(n26), .Z(o[36]) );
  AND U17 ( .A(o[7]), .B(n27), .Z(n25) );
  XOR U18 ( .A(n28), .B(n29), .Z(n27) );
  XOR U19 ( .A(n30), .B(n31), .Z(o[35]) );
  AND U20 ( .A(o[7]), .B(n32), .Z(n30) );
  XOR U21 ( .A(n33), .B(n34), .Z(n32) );
  XOR U22 ( .A(n35), .B(n36), .Z(o[34]) );
  AND U23 ( .A(o[7]), .B(n37), .Z(n35) );
  XOR U24 ( .A(n38), .B(n39), .Z(n37) );
  XOR U25 ( .A(n40), .B(n41), .Z(o[33]) );
  AND U26 ( .A(o[7]), .B(n42), .Z(n40) );
  XOR U27 ( .A(n43), .B(n44), .Z(n42) );
  XOR U28 ( .A(n45), .B(n46), .Z(o[32]) );
  AND U29 ( .A(o[7]), .B(n47), .Z(n45) );
  XOR U30 ( .A(n48), .B(n49), .Z(n47) );
  XOR U31 ( .A(n50), .B(n51), .Z(o[31]) );
  AND U32 ( .A(o[7]), .B(n52), .Z(n50) );
  XOR U33 ( .A(n53), .B(n54), .Z(n52) );
  XOR U34 ( .A(n55), .B(n56), .Z(o[30]) );
  AND U35 ( .A(o[7]), .B(n57), .Z(n55) );
  XOR U36 ( .A(n58), .B(n59), .Z(n57) );
  XOR U37 ( .A(n60), .B(n61), .Z(o[29]) );
  AND U38 ( .A(o[7]), .B(n62), .Z(n60) );
  XOR U39 ( .A(n63), .B(n64), .Z(n62) );
  XOR U40 ( .A(n65), .B(n66), .Z(o[28]) );
  AND U41 ( .A(o[7]), .B(n67), .Z(n65) );
  XOR U42 ( .A(n68), .B(n69), .Z(n67) );
  XOR U43 ( .A(n70), .B(n71), .Z(o[27]) );
  AND U44 ( .A(o[7]), .B(n72), .Z(n70) );
  XOR U45 ( .A(n73), .B(n74), .Z(n72) );
  XOR U46 ( .A(n75), .B(n76), .Z(o[26]) );
  AND U47 ( .A(o[7]), .B(n77), .Z(n75) );
  XOR U48 ( .A(n78), .B(n79), .Z(n77) );
  XOR U49 ( .A(n80), .B(n81), .Z(o[25]) );
  AND U50 ( .A(o[7]), .B(n82), .Z(n80) );
  XOR U51 ( .A(n83), .B(n84), .Z(n82) );
  XOR U52 ( .A(n85), .B(n86), .Z(o[24]) );
  AND U53 ( .A(o[7]), .B(n87), .Z(n85) );
  XOR U54 ( .A(n88), .B(n89), .Z(n87) );
  XOR U55 ( .A(n90), .B(n91), .Z(o[23]) );
  AND U56 ( .A(o[7]), .B(n92), .Z(n90) );
  XOR U57 ( .A(n93), .B(n94), .Z(n92) );
  XOR U58 ( .A(n95), .B(n96), .Z(o[22]) );
  AND U59 ( .A(o[7]), .B(n97), .Z(n95) );
  XOR U60 ( .A(n98), .B(n99), .Z(n97) );
  XOR U61 ( .A(n100), .B(n101), .Z(o[21]) );
  AND U62 ( .A(o[7]), .B(n102), .Z(n100) );
  XOR U63 ( .A(n103), .B(n104), .Z(n102) );
  XOR U64 ( .A(n105), .B(n106), .Z(o[20]) );
  AND U65 ( .A(o[7]), .B(n107), .Z(n105) );
  XOR U66 ( .A(n108), .B(n109), .Z(n107) );
  XOR U67 ( .A(n110), .B(n111), .Z(o[19]) );
  AND U68 ( .A(o[7]), .B(n112), .Z(n110) );
  XOR U69 ( .A(n113), .B(n114), .Z(n112) );
  XOR U70 ( .A(n115), .B(n116), .Z(o[18]) );
  AND U71 ( .A(o[7]), .B(n117), .Z(n115) );
  XOR U72 ( .A(n118), .B(n119), .Z(n117) );
  XOR U73 ( .A(n120), .B(n121), .Z(o[17]) );
  AND U74 ( .A(o[7]), .B(n122), .Z(n120) );
  XOR U75 ( .A(n123), .B(n124), .Z(n122) );
  XOR U76 ( .A(n125), .B(n126), .Z(o[16]) );
  AND U77 ( .A(o[7]), .B(n127), .Z(n125) );
  XOR U78 ( .A(n128), .B(n129), .Z(n127) );
  XOR U79 ( .A(n130), .B(n131), .Z(o[15]) );
  AND U80 ( .A(o[7]), .B(n132), .Z(n130) );
  XOR U81 ( .A(n133), .B(n134), .Z(n132) );
  XOR U82 ( .A(n135), .B(n136), .Z(o[14]) );
  AND U83 ( .A(o[7]), .B(n137), .Z(n135) );
  XOR U84 ( .A(n138), .B(n139), .Z(n137) );
  XOR U85 ( .A(n140), .B(n141), .Z(o[13]) );
  AND U86 ( .A(o[7]), .B(n142), .Z(n140) );
  XOR U87 ( .A(n143), .B(n144), .Z(n142) );
  XOR U88 ( .A(n145), .B(n146), .Z(o[12]) );
  AND U89 ( .A(o[7]), .B(n147), .Z(n145) );
  XOR U90 ( .A(n148), .B(n149), .Z(n147) );
  XOR U91 ( .A(n150), .B(n151), .Z(o[11]) );
  AND U92 ( .A(o[7]), .B(n152), .Z(n150) );
  XOR U93 ( .A(n153), .B(n154), .Z(n152) );
  XOR U94 ( .A(n155), .B(n156), .Z(o[10]) );
  AND U95 ( .A(o[7]), .B(n157), .Z(n155) );
  XOR U96 ( .A(n158), .B(n159), .Z(n157) );
  XOR U97 ( .A(n160), .B(n161), .Z(o[0]) );
  AND U98 ( .A(o[1]), .B(n162), .Z(n161) );
  XNOR U99 ( .A(n163), .B(n164), .Z(n162) );
  XNOR U100 ( .A(n165), .B(n160), .Z(n164) );
  AND U101 ( .A(o[2]), .B(n166), .Z(n165) );
  XNOR U102 ( .A(n167), .B(n168), .Z(n166) );
  XNOR U103 ( .A(n169), .B(n163), .Z(n168) );
  AND U104 ( .A(o[3]), .B(n170), .Z(n169) );
  XNOR U105 ( .A(n171), .B(n172), .Z(n170) );
  XNOR U106 ( .A(n173), .B(n167), .Z(n172) );
  AND U107 ( .A(o[4]), .B(n174), .Z(n173) );
  XNOR U108 ( .A(n175), .B(n176), .Z(n174) );
  XNOR U109 ( .A(n177), .B(n171), .Z(n176) );
  AND U110 ( .A(o[5]), .B(n178), .Z(n177) );
  XNOR U111 ( .A(n179), .B(n180), .Z(n178) );
  XNOR U112 ( .A(n181), .B(n175), .Z(n180) );
  AND U113 ( .A(o[6]), .B(n182), .Z(n181) );
  XNOR U114 ( .A(n179), .B(n183), .Z(n182) );
  XNOR U115 ( .A(n184), .B(n185), .Z(n183) );
  AND U116 ( .A(o[7]), .B(n186), .Z(n184) );
  XOR U117 ( .A(n185), .B(n187), .Z(n186) );
  XOR U118 ( .A(n188), .B(n189), .Z(n179) );
  AND U119 ( .A(o[7]), .B(n190), .Z(n189) );
  XOR U120 ( .A(n188), .B(n191), .Z(n190) );
  XOR U121 ( .A(n192), .B(n193), .Z(n175) );
  AND U122 ( .A(o[6]), .B(n194), .Z(n193) );
  XNOR U123 ( .A(n192), .B(n195), .Z(n194) );
  XNOR U124 ( .A(n196), .B(n197), .Z(n195) );
  AND U125 ( .A(o[7]), .B(n198), .Z(n196) );
  XOR U126 ( .A(n197), .B(n199), .Z(n198) );
  XOR U127 ( .A(n200), .B(n201), .Z(n192) );
  AND U128 ( .A(o[7]), .B(n202), .Z(n201) );
  XOR U129 ( .A(n200), .B(n203), .Z(n202) );
  XOR U130 ( .A(n204), .B(n205), .Z(n171) );
  AND U131 ( .A(o[5]), .B(n206), .Z(n205) );
  XNOR U132 ( .A(n207), .B(n208), .Z(n206) );
  XNOR U133 ( .A(n209), .B(n204), .Z(n208) );
  AND U134 ( .A(o[6]), .B(n210), .Z(n209) );
  XNOR U135 ( .A(n207), .B(n211), .Z(n210) );
  XNOR U136 ( .A(n212), .B(n213), .Z(n211) );
  AND U137 ( .A(o[7]), .B(n214), .Z(n212) );
  XOR U138 ( .A(n213), .B(n215), .Z(n214) );
  XOR U139 ( .A(n216), .B(n217), .Z(n207) );
  AND U140 ( .A(o[7]), .B(n218), .Z(n217) );
  XOR U141 ( .A(n216), .B(n219), .Z(n218) );
  XOR U142 ( .A(n220), .B(n221), .Z(n204) );
  AND U143 ( .A(o[6]), .B(n222), .Z(n221) );
  XNOR U144 ( .A(n220), .B(n223), .Z(n222) );
  XNOR U145 ( .A(n224), .B(n225), .Z(n223) );
  AND U146 ( .A(o[7]), .B(n226), .Z(n224) );
  XOR U147 ( .A(n225), .B(n227), .Z(n226) );
  XOR U148 ( .A(n228), .B(n229), .Z(n220) );
  AND U149 ( .A(o[7]), .B(n230), .Z(n229) );
  XOR U150 ( .A(n228), .B(n231), .Z(n230) );
  XOR U151 ( .A(n232), .B(n233), .Z(n167) );
  AND U152 ( .A(o[4]), .B(n234), .Z(n233) );
  XNOR U153 ( .A(n235), .B(n236), .Z(n234) );
  XNOR U154 ( .A(n237), .B(n232), .Z(n236) );
  AND U155 ( .A(o[5]), .B(n238), .Z(n237) );
  XNOR U156 ( .A(n239), .B(n240), .Z(n238) );
  XNOR U157 ( .A(n241), .B(n235), .Z(n240) );
  AND U158 ( .A(o[6]), .B(n242), .Z(n241) );
  XNOR U159 ( .A(n239), .B(n243), .Z(n242) );
  XNOR U160 ( .A(n244), .B(n245), .Z(n243) );
  AND U161 ( .A(o[7]), .B(n246), .Z(n244) );
  XOR U162 ( .A(n245), .B(n247), .Z(n246) );
  XOR U163 ( .A(n248), .B(n249), .Z(n239) );
  AND U164 ( .A(o[7]), .B(n250), .Z(n249) );
  XOR U165 ( .A(n248), .B(n251), .Z(n250) );
  XOR U166 ( .A(n252), .B(n253), .Z(n235) );
  AND U167 ( .A(o[6]), .B(n254), .Z(n253) );
  XNOR U168 ( .A(n252), .B(n255), .Z(n254) );
  XNOR U169 ( .A(n256), .B(n257), .Z(n255) );
  AND U170 ( .A(o[7]), .B(n258), .Z(n256) );
  XOR U171 ( .A(n257), .B(n259), .Z(n258) );
  XOR U172 ( .A(n260), .B(n261), .Z(n252) );
  AND U173 ( .A(o[7]), .B(n262), .Z(n261) );
  XOR U174 ( .A(n260), .B(n263), .Z(n262) );
  XOR U175 ( .A(n264), .B(n265), .Z(n232) );
  AND U176 ( .A(o[5]), .B(n266), .Z(n265) );
  XNOR U177 ( .A(n267), .B(n268), .Z(n266) );
  XNOR U178 ( .A(n269), .B(n264), .Z(n268) );
  AND U179 ( .A(o[6]), .B(n270), .Z(n269) );
  XNOR U180 ( .A(n267), .B(n271), .Z(n270) );
  XNOR U181 ( .A(n272), .B(n273), .Z(n271) );
  AND U182 ( .A(o[7]), .B(n274), .Z(n272) );
  XOR U183 ( .A(n273), .B(n275), .Z(n274) );
  XOR U184 ( .A(n276), .B(n277), .Z(n267) );
  AND U185 ( .A(o[7]), .B(n278), .Z(n277) );
  XOR U186 ( .A(n276), .B(n279), .Z(n278) );
  XOR U187 ( .A(n280), .B(n281), .Z(n264) );
  AND U188 ( .A(o[6]), .B(n282), .Z(n281) );
  XNOR U189 ( .A(n280), .B(n283), .Z(n282) );
  XNOR U190 ( .A(n284), .B(n285), .Z(n283) );
  AND U191 ( .A(o[7]), .B(n286), .Z(n284) );
  XOR U192 ( .A(n285), .B(n287), .Z(n286) );
  XOR U193 ( .A(n288), .B(n289), .Z(n280) );
  AND U194 ( .A(o[7]), .B(n290), .Z(n289) );
  XOR U195 ( .A(n288), .B(n291), .Z(n290) );
  XOR U196 ( .A(n292), .B(n293), .Z(n163) );
  AND U197 ( .A(o[3]), .B(n294), .Z(n293) );
  XNOR U198 ( .A(n295), .B(n296), .Z(n294) );
  XNOR U199 ( .A(n297), .B(n292), .Z(n296) );
  AND U200 ( .A(o[4]), .B(n298), .Z(n297) );
  XNOR U201 ( .A(n299), .B(n300), .Z(n298) );
  XNOR U202 ( .A(n301), .B(n295), .Z(n300) );
  AND U203 ( .A(o[5]), .B(n302), .Z(n301) );
  XNOR U204 ( .A(n303), .B(n304), .Z(n302) );
  XNOR U205 ( .A(n305), .B(n299), .Z(n304) );
  AND U206 ( .A(o[6]), .B(n306), .Z(n305) );
  XNOR U207 ( .A(n303), .B(n307), .Z(n306) );
  XNOR U208 ( .A(n308), .B(n309), .Z(n307) );
  AND U209 ( .A(o[7]), .B(n310), .Z(n308) );
  XOR U210 ( .A(n309), .B(n311), .Z(n310) );
  XOR U211 ( .A(n312), .B(n313), .Z(n303) );
  AND U212 ( .A(o[7]), .B(n314), .Z(n313) );
  XOR U213 ( .A(n312), .B(n315), .Z(n314) );
  XOR U214 ( .A(n316), .B(n317), .Z(n299) );
  AND U215 ( .A(o[6]), .B(n318), .Z(n317) );
  XNOR U216 ( .A(n316), .B(n319), .Z(n318) );
  XNOR U217 ( .A(n320), .B(n321), .Z(n319) );
  AND U218 ( .A(o[7]), .B(n322), .Z(n320) );
  XOR U219 ( .A(n321), .B(n323), .Z(n322) );
  XOR U220 ( .A(n324), .B(n325), .Z(n316) );
  AND U221 ( .A(o[7]), .B(n326), .Z(n325) );
  XOR U222 ( .A(n324), .B(n327), .Z(n326) );
  XOR U223 ( .A(n328), .B(n329), .Z(n295) );
  AND U224 ( .A(o[5]), .B(n330), .Z(n329) );
  XNOR U225 ( .A(n331), .B(n332), .Z(n330) );
  XNOR U226 ( .A(n333), .B(n328), .Z(n332) );
  AND U227 ( .A(o[6]), .B(n334), .Z(n333) );
  XNOR U228 ( .A(n331), .B(n335), .Z(n334) );
  XNOR U229 ( .A(n336), .B(n337), .Z(n335) );
  AND U230 ( .A(o[7]), .B(n338), .Z(n336) );
  XOR U231 ( .A(n337), .B(n339), .Z(n338) );
  XOR U232 ( .A(n340), .B(n341), .Z(n331) );
  AND U233 ( .A(o[7]), .B(n342), .Z(n341) );
  XOR U234 ( .A(n340), .B(n343), .Z(n342) );
  XOR U235 ( .A(n344), .B(n345), .Z(n328) );
  AND U236 ( .A(o[6]), .B(n346), .Z(n345) );
  XNOR U237 ( .A(n344), .B(n347), .Z(n346) );
  XNOR U238 ( .A(n348), .B(n349), .Z(n347) );
  AND U239 ( .A(o[7]), .B(n350), .Z(n348) );
  XOR U240 ( .A(n349), .B(n351), .Z(n350) );
  XOR U241 ( .A(n352), .B(n353), .Z(n344) );
  AND U242 ( .A(o[7]), .B(n354), .Z(n353) );
  XOR U243 ( .A(n352), .B(n355), .Z(n354) );
  XOR U244 ( .A(n356), .B(n357), .Z(n292) );
  AND U245 ( .A(o[4]), .B(n358), .Z(n357) );
  XNOR U246 ( .A(n359), .B(n360), .Z(n358) );
  XNOR U247 ( .A(n361), .B(n356), .Z(n360) );
  AND U248 ( .A(o[5]), .B(n362), .Z(n361) );
  XNOR U249 ( .A(n363), .B(n364), .Z(n362) );
  XNOR U250 ( .A(n365), .B(n359), .Z(n364) );
  AND U251 ( .A(o[6]), .B(n366), .Z(n365) );
  XNOR U252 ( .A(n363), .B(n367), .Z(n366) );
  XNOR U253 ( .A(n368), .B(n369), .Z(n367) );
  AND U254 ( .A(o[7]), .B(n370), .Z(n368) );
  XOR U255 ( .A(n369), .B(n371), .Z(n370) );
  XOR U256 ( .A(n372), .B(n373), .Z(n363) );
  AND U257 ( .A(o[7]), .B(n374), .Z(n373) );
  XOR U258 ( .A(n372), .B(n375), .Z(n374) );
  XOR U259 ( .A(n376), .B(n377), .Z(n359) );
  AND U260 ( .A(o[6]), .B(n378), .Z(n377) );
  XNOR U261 ( .A(n376), .B(n379), .Z(n378) );
  XNOR U262 ( .A(n380), .B(n381), .Z(n379) );
  AND U263 ( .A(o[7]), .B(n382), .Z(n380) );
  XOR U264 ( .A(n381), .B(n383), .Z(n382) );
  XOR U265 ( .A(n384), .B(n385), .Z(n376) );
  AND U266 ( .A(o[7]), .B(n386), .Z(n385) );
  XOR U267 ( .A(n384), .B(n387), .Z(n386) );
  XOR U268 ( .A(n388), .B(n389), .Z(n356) );
  AND U269 ( .A(o[5]), .B(n390), .Z(n389) );
  XNOR U270 ( .A(n391), .B(n392), .Z(n390) );
  XNOR U271 ( .A(n393), .B(n388), .Z(n392) );
  AND U272 ( .A(o[6]), .B(n394), .Z(n393) );
  XNOR U273 ( .A(n391), .B(n395), .Z(n394) );
  XNOR U274 ( .A(n396), .B(n397), .Z(n395) );
  AND U275 ( .A(o[7]), .B(n398), .Z(n396) );
  XOR U276 ( .A(n397), .B(n399), .Z(n398) );
  XOR U277 ( .A(n400), .B(n401), .Z(n391) );
  AND U278 ( .A(o[7]), .B(n402), .Z(n401) );
  XOR U279 ( .A(n400), .B(n403), .Z(n402) );
  XOR U280 ( .A(n404), .B(n405), .Z(n388) );
  AND U281 ( .A(o[6]), .B(n406), .Z(n405) );
  XNOR U282 ( .A(n404), .B(n407), .Z(n406) );
  XNOR U283 ( .A(n408), .B(n409), .Z(n407) );
  AND U284 ( .A(o[7]), .B(n410), .Z(n408) );
  XOR U285 ( .A(n409), .B(n411), .Z(n410) );
  XOR U286 ( .A(n412), .B(n413), .Z(n404) );
  AND U287 ( .A(o[7]), .B(n414), .Z(n413) );
  XOR U288 ( .A(n412), .B(n415), .Z(n414) );
  XOR U289 ( .A(n416), .B(n417), .Z(o[1]) );
  AND U290 ( .A(o[2]), .B(n418), .Z(n417) );
  XNOR U291 ( .A(n419), .B(n420), .Z(n418) );
  XNOR U292 ( .A(n421), .B(n416), .Z(n420) );
  AND U293 ( .A(o[3]), .B(n422), .Z(n421) );
  XNOR U294 ( .A(n423), .B(n424), .Z(n422) );
  XNOR U295 ( .A(n425), .B(n419), .Z(n424) );
  AND U296 ( .A(o[4]), .B(n426), .Z(n425) );
  XNOR U297 ( .A(n427), .B(n428), .Z(n426) );
  XNOR U298 ( .A(n429), .B(n423), .Z(n428) );
  AND U299 ( .A(o[5]), .B(n430), .Z(n429) );
  XNOR U300 ( .A(n431), .B(n432), .Z(n430) );
  XNOR U301 ( .A(n433), .B(n427), .Z(n432) );
  AND U302 ( .A(o[6]), .B(n434), .Z(n433) );
  XNOR U303 ( .A(n431), .B(n435), .Z(n434) );
  XNOR U304 ( .A(n436), .B(n437), .Z(n435) );
  AND U305 ( .A(o[7]), .B(n438), .Z(n436) );
  XOR U306 ( .A(n437), .B(n439), .Z(n438) );
  XOR U307 ( .A(n440), .B(n441), .Z(n431) );
  AND U308 ( .A(o[7]), .B(n442), .Z(n441) );
  XOR U309 ( .A(n440), .B(n443), .Z(n442) );
  XOR U310 ( .A(n444), .B(n445), .Z(n427) );
  AND U311 ( .A(o[6]), .B(n446), .Z(n445) );
  XNOR U312 ( .A(n444), .B(n447), .Z(n446) );
  XNOR U313 ( .A(n448), .B(n449), .Z(n447) );
  AND U314 ( .A(o[7]), .B(n450), .Z(n448) );
  XOR U315 ( .A(n449), .B(n451), .Z(n450) );
  XOR U316 ( .A(n452), .B(n453), .Z(n444) );
  AND U317 ( .A(o[7]), .B(n454), .Z(n453) );
  XOR U318 ( .A(n452), .B(n455), .Z(n454) );
  XOR U319 ( .A(n456), .B(n457), .Z(n423) );
  AND U320 ( .A(o[5]), .B(n458), .Z(n457) );
  XNOR U321 ( .A(n459), .B(n460), .Z(n458) );
  XNOR U322 ( .A(n461), .B(n456), .Z(n460) );
  AND U323 ( .A(o[6]), .B(n462), .Z(n461) );
  XNOR U324 ( .A(n459), .B(n463), .Z(n462) );
  XNOR U325 ( .A(n464), .B(n465), .Z(n463) );
  AND U326 ( .A(o[7]), .B(n466), .Z(n464) );
  XOR U327 ( .A(n465), .B(n467), .Z(n466) );
  XOR U328 ( .A(n468), .B(n469), .Z(n459) );
  AND U329 ( .A(o[7]), .B(n470), .Z(n469) );
  XOR U330 ( .A(n468), .B(n471), .Z(n470) );
  XOR U331 ( .A(n472), .B(n473), .Z(n456) );
  AND U332 ( .A(o[6]), .B(n474), .Z(n473) );
  XNOR U333 ( .A(n472), .B(n475), .Z(n474) );
  XNOR U334 ( .A(n476), .B(n477), .Z(n475) );
  AND U335 ( .A(o[7]), .B(n478), .Z(n476) );
  XOR U336 ( .A(n477), .B(n479), .Z(n478) );
  XOR U337 ( .A(n480), .B(n481), .Z(n472) );
  AND U338 ( .A(o[7]), .B(n482), .Z(n481) );
  XOR U339 ( .A(n480), .B(n483), .Z(n482) );
  XOR U340 ( .A(n484), .B(n485), .Z(n419) );
  AND U341 ( .A(o[4]), .B(n486), .Z(n485) );
  XNOR U342 ( .A(n487), .B(n488), .Z(n486) );
  XNOR U343 ( .A(n489), .B(n484), .Z(n488) );
  AND U344 ( .A(o[5]), .B(n490), .Z(n489) );
  XNOR U345 ( .A(n491), .B(n492), .Z(n490) );
  XNOR U346 ( .A(n493), .B(n487), .Z(n492) );
  AND U347 ( .A(o[6]), .B(n494), .Z(n493) );
  XNOR U348 ( .A(n491), .B(n495), .Z(n494) );
  XNOR U349 ( .A(n496), .B(n497), .Z(n495) );
  AND U350 ( .A(o[7]), .B(n498), .Z(n496) );
  XOR U351 ( .A(n497), .B(n499), .Z(n498) );
  XOR U352 ( .A(n500), .B(n501), .Z(n491) );
  AND U353 ( .A(o[7]), .B(n502), .Z(n501) );
  XOR U354 ( .A(n500), .B(n503), .Z(n502) );
  XOR U355 ( .A(n504), .B(n505), .Z(n487) );
  AND U356 ( .A(o[6]), .B(n506), .Z(n505) );
  XNOR U357 ( .A(n504), .B(n507), .Z(n506) );
  XNOR U358 ( .A(n508), .B(n509), .Z(n507) );
  AND U359 ( .A(o[7]), .B(n510), .Z(n508) );
  XOR U360 ( .A(n509), .B(n511), .Z(n510) );
  XOR U361 ( .A(n512), .B(n513), .Z(n504) );
  AND U362 ( .A(o[7]), .B(n514), .Z(n513) );
  XOR U363 ( .A(n512), .B(n515), .Z(n514) );
  XOR U364 ( .A(n516), .B(n517), .Z(n484) );
  AND U365 ( .A(o[5]), .B(n518), .Z(n517) );
  XNOR U366 ( .A(n519), .B(n520), .Z(n518) );
  XNOR U367 ( .A(n521), .B(n516), .Z(n520) );
  AND U368 ( .A(o[6]), .B(n522), .Z(n521) );
  XNOR U369 ( .A(n519), .B(n523), .Z(n522) );
  XNOR U370 ( .A(n524), .B(n525), .Z(n523) );
  AND U371 ( .A(o[7]), .B(n526), .Z(n524) );
  XOR U372 ( .A(n525), .B(n527), .Z(n526) );
  XOR U373 ( .A(n528), .B(n529), .Z(n519) );
  AND U374 ( .A(o[7]), .B(n530), .Z(n529) );
  XOR U375 ( .A(n528), .B(n531), .Z(n530) );
  XOR U376 ( .A(n532), .B(n533), .Z(n516) );
  AND U377 ( .A(o[6]), .B(n534), .Z(n533) );
  XNOR U378 ( .A(n532), .B(n535), .Z(n534) );
  XNOR U379 ( .A(n536), .B(n537), .Z(n535) );
  AND U380 ( .A(o[7]), .B(n538), .Z(n536) );
  XOR U381 ( .A(n537), .B(n539), .Z(n538) );
  XOR U382 ( .A(n540), .B(n541), .Z(n532) );
  AND U383 ( .A(o[7]), .B(n542), .Z(n541) );
  XOR U384 ( .A(n540), .B(n543), .Z(n542) );
  XOR U385 ( .A(n544), .B(n545), .Z(n416) );
  AND U386 ( .A(o[3]), .B(n546), .Z(n545) );
  XNOR U387 ( .A(n547), .B(n548), .Z(n546) );
  XNOR U388 ( .A(n549), .B(n544), .Z(n548) );
  AND U389 ( .A(o[4]), .B(n550), .Z(n549) );
  XNOR U390 ( .A(n551), .B(n552), .Z(n550) );
  XNOR U391 ( .A(n553), .B(n547), .Z(n552) );
  AND U392 ( .A(o[5]), .B(n554), .Z(n553) );
  XNOR U393 ( .A(n555), .B(n556), .Z(n554) );
  XNOR U394 ( .A(n557), .B(n551), .Z(n556) );
  AND U395 ( .A(o[6]), .B(n558), .Z(n557) );
  XNOR U396 ( .A(n555), .B(n559), .Z(n558) );
  XNOR U397 ( .A(n560), .B(n561), .Z(n559) );
  AND U398 ( .A(o[7]), .B(n562), .Z(n560) );
  XOR U399 ( .A(n561), .B(n563), .Z(n562) );
  XOR U400 ( .A(n564), .B(n565), .Z(n555) );
  AND U401 ( .A(o[7]), .B(n566), .Z(n565) );
  XOR U402 ( .A(n564), .B(n567), .Z(n566) );
  XOR U403 ( .A(n568), .B(n569), .Z(n551) );
  AND U404 ( .A(o[6]), .B(n570), .Z(n569) );
  XNOR U405 ( .A(n568), .B(n571), .Z(n570) );
  XNOR U406 ( .A(n572), .B(n573), .Z(n571) );
  AND U407 ( .A(o[7]), .B(n574), .Z(n572) );
  XOR U408 ( .A(n573), .B(n575), .Z(n574) );
  XOR U409 ( .A(n576), .B(n577), .Z(n568) );
  AND U410 ( .A(o[7]), .B(n578), .Z(n577) );
  XOR U411 ( .A(n576), .B(n579), .Z(n578) );
  XOR U412 ( .A(n580), .B(n581), .Z(n547) );
  AND U413 ( .A(o[5]), .B(n582), .Z(n581) );
  XNOR U414 ( .A(n583), .B(n584), .Z(n582) );
  XNOR U415 ( .A(n585), .B(n580), .Z(n584) );
  AND U416 ( .A(o[6]), .B(n586), .Z(n585) );
  XNOR U417 ( .A(n583), .B(n587), .Z(n586) );
  XNOR U418 ( .A(n588), .B(n589), .Z(n587) );
  AND U419 ( .A(o[7]), .B(n590), .Z(n588) );
  XOR U420 ( .A(n589), .B(n591), .Z(n590) );
  XOR U421 ( .A(n592), .B(n593), .Z(n583) );
  AND U422 ( .A(o[7]), .B(n594), .Z(n593) );
  XOR U423 ( .A(n592), .B(n595), .Z(n594) );
  XOR U424 ( .A(n596), .B(n597), .Z(n580) );
  AND U425 ( .A(o[6]), .B(n598), .Z(n597) );
  XNOR U426 ( .A(n596), .B(n599), .Z(n598) );
  XNOR U427 ( .A(n600), .B(n601), .Z(n599) );
  AND U428 ( .A(o[7]), .B(n602), .Z(n600) );
  XOR U429 ( .A(n601), .B(n603), .Z(n602) );
  XOR U430 ( .A(n604), .B(n605), .Z(n596) );
  AND U431 ( .A(o[7]), .B(n606), .Z(n605) );
  XOR U432 ( .A(n604), .B(n607), .Z(n606) );
  XOR U433 ( .A(n608), .B(n609), .Z(n544) );
  AND U434 ( .A(o[4]), .B(n610), .Z(n609) );
  XNOR U435 ( .A(n611), .B(n612), .Z(n610) );
  XNOR U436 ( .A(n613), .B(n608), .Z(n612) );
  AND U437 ( .A(o[5]), .B(n614), .Z(n613) );
  XNOR U438 ( .A(n615), .B(n616), .Z(n614) );
  XNOR U439 ( .A(n617), .B(n611), .Z(n616) );
  AND U440 ( .A(o[6]), .B(n618), .Z(n617) );
  XNOR U441 ( .A(n615), .B(n619), .Z(n618) );
  XNOR U442 ( .A(n620), .B(n621), .Z(n619) );
  AND U443 ( .A(o[7]), .B(n622), .Z(n620) );
  XOR U444 ( .A(n621), .B(n623), .Z(n622) );
  XOR U445 ( .A(n624), .B(n625), .Z(n615) );
  AND U446 ( .A(o[7]), .B(n626), .Z(n625) );
  XOR U447 ( .A(n624), .B(n627), .Z(n626) );
  XOR U448 ( .A(n628), .B(n629), .Z(n611) );
  AND U449 ( .A(o[6]), .B(n630), .Z(n629) );
  XNOR U450 ( .A(n628), .B(n631), .Z(n630) );
  XNOR U451 ( .A(n632), .B(n633), .Z(n631) );
  AND U452 ( .A(o[7]), .B(n634), .Z(n632) );
  XOR U453 ( .A(n633), .B(n635), .Z(n634) );
  XOR U454 ( .A(n636), .B(n637), .Z(n628) );
  AND U455 ( .A(o[7]), .B(n638), .Z(n637) );
  XOR U456 ( .A(n636), .B(n639), .Z(n638) );
  XOR U457 ( .A(n640), .B(n641), .Z(n608) );
  AND U458 ( .A(o[5]), .B(n642), .Z(n641) );
  XNOR U459 ( .A(n643), .B(n644), .Z(n642) );
  XNOR U460 ( .A(n645), .B(n640), .Z(n644) );
  AND U461 ( .A(o[6]), .B(n646), .Z(n645) );
  XNOR U462 ( .A(n643), .B(n647), .Z(n646) );
  XNOR U463 ( .A(n648), .B(n649), .Z(n647) );
  AND U464 ( .A(o[7]), .B(n650), .Z(n648) );
  XOR U465 ( .A(n649), .B(n651), .Z(n650) );
  XOR U466 ( .A(n652), .B(n653), .Z(n643) );
  AND U467 ( .A(o[7]), .B(n654), .Z(n653) );
  XOR U468 ( .A(n652), .B(n655), .Z(n654) );
  XOR U469 ( .A(n656), .B(n657), .Z(n640) );
  AND U470 ( .A(o[6]), .B(n658), .Z(n657) );
  XNOR U471 ( .A(n656), .B(n659), .Z(n658) );
  XNOR U472 ( .A(n660), .B(n661), .Z(n659) );
  AND U473 ( .A(o[7]), .B(n662), .Z(n660) );
  XOR U474 ( .A(n661), .B(n663), .Z(n662) );
  XOR U475 ( .A(n664), .B(n665), .Z(n656) );
  AND U476 ( .A(o[7]), .B(n666), .Z(n665) );
  XOR U477 ( .A(n664), .B(n667), .Z(n666) );
  XOR U478 ( .A(n668), .B(n669), .Z(n160) );
  AND U479 ( .A(o[2]), .B(n670), .Z(n669) );
  XNOR U480 ( .A(n671), .B(n672), .Z(n670) );
  XNOR U481 ( .A(n673), .B(n668), .Z(n672) );
  AND U482 ( .A(o[3]), .B(n674), .Z(n673) );
  XNOR U483 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U484 ( .A(n677), .B(n671), .Z(n676) );
  AND U485 ( .A(o[4]), .B(n678), .Z(n677) );
  XNOR U486 ( .A(n679), .B(n680), .Z(n678) );
  XNOR U487 ( .A(n681), .B(n675), .Z(n680) );
  AND U488 ( .A(o[5]), .B(n682), .Z(n681) );
  XNOR U489 ( .A(n683), .B(n684), .Z(n682) );
  XNOR U490 ( .A(n685), .B(n679), .Z(n684) );
  AND U491 ( .A(o[6]), .B(n686), .Z(n685) );
  XNOR U492 ( .A(n683), .B(n687), .Z(n686) );
  XNOR U493 ( .A(n688), .B(n689), .Z(n687) );
  AND U494 ( .A(o[7]), .B(n690), .Z(n688) );
  XOR U495 ( .A(n689), .B(n691), .Z(n690) );
  XOR U496 ( .A(n692), .B(n693), .Z(n683) );
  AND U497 ( .A(o[7]), .B(n694), .Z(n693) );
  XOR U498 ( .A(n692), .B(n695), .Z(n694) );
  XOR U499 ( .A(n696), .B(n697), .Z(n679) );
  AND U500 ( .A(o[6]), .B(n698), .Z(n697) );
  XNOR U501 ( .A(n696), .B(n699), .Z(n698) );
  XNOR U502 ( .A(n700), .B(n701), .Z(n699) );
  AND U503 ( .A(o[7]), .B(n702), .Z(n700) );
  XOR U504 ( .A(n701), .B(n703), .Z(n702) );
  XOR U505 ( .A(n704), .B(n705), .Z(n696) );
  AND U506 ( .A(o[7]), .B(n706), .Z(n705) );
  XOR U507 ( .A(n704), .B(n707), .Z(n706) );
  XOR U508 ( .A(n708), .B(n709), .Z(n675) );
  AND U509 ( .A(o[5]), .B(n710), .Z(n709) );
  XNOR U510 ( .A(n711), .B(n712), .Z(n710) );
  XNOR U511 ( .A(n713), .B(n708), .Z(n712) );
  AND U512 ( .A(o[6]), .B(n714), .Z(n713) );
  XNOR U513 ( .A(n711), .B(n715), .Z(n714) );
  XNOR U514 ( .A(n716), .B(n717), .Z(n715) );
  AND U515 ( .A(o[7]), .B(n718), .Z(n716) );
  XOR U516 ( .A(n717), .B(n719), .Z(n718) );
  XOR U517 ( .A(n720), .B(n721), .Z(n711) );
  AND U518 ( .A(o[7]), .B(n722), .Z(n721) );
  XOR U519 ( .A(n720), .B(n723), .Z(n722) );
  XOR U520 ( .A(n724), .B(n725), .Z(n708) );
  AND U521 ( .A(o[6]), .B(n726), .Z(n725) );
  XNOR U522 ( .A(n724), .B(n727), .Z(n726) );
  XNOR U523 ( .A(n728), .B(n729), .Z(n727) );
  AND U524 ( .A(o[7]), .B(n730), .Z(n728) );
  XOR U525 ( .A(n729), .B(n731), .Z(n730) );
  XOR U526 ( .A(n732), .B(n733), .Z(n724) );
  AND U527 ( .A(o[7]), .B(n734), .Z(n733) );
  XOR U528 ( .A(n732), .B(n735), .Z(n734) );
  XOR U529 ( .A(n736), .B(n737), .Z(n671) );
  AND U530 ( .A(o[4]), .B(n738), .Z(n737) );
  XNOR U531 ( .A(n739), .B(n740), .Z(n738) );
  XNOR U532 ( .A(n741), .B(n736), .Z(n740) );
  AND U533 ( .A(o[5]), .B(n742), .Z(n741) );
  XNOR U534 ( .A(n743), .B(n744), .Z(n742) );
  XNOR U535 ( .A(n745), .B(n739), .Z(n744) );
  AND U536 ( .A(o[6]), .B(n746), .Z(n745) );
  XNOR U537 ( .A(n743), .B(n747), .Z(n746) );
  XNOR U538 ( .A(n748), .B(n749), .Z(n747) );
  AND U539 ( .A(o[7]), .B(n750), .Z(n748) );
  XOR U540 ( .A(n749), .B(n751), .Z(n750) );
  XOR U541 ( .A(n752), .B(n753), .Z(n743) );
  AND U542 ( .A(o[7]), .B(n754), .Z(n753) );
  XOR U543 ( .A(n752), .B(n755), .Z(n754) );
  XOR U544 ( .A(n756), .B(n757), .Z(n739) );
  AND U545 ( .A(o[6]), .B(n758), .Z(n757) );
  XNOR U546 ( .A(n756), .B(n759), .Z(n758) );
  XNOR U547 ( .A(n760), .B(n761), .Z(n759) );
  AND U548 ( .A(o[7]), .B(n762), .Z(n760) );
  XOR U549 ( .A(n761), .B(n763), .Z(n762) );
  XOR U550 ( .A(n764), .B(n765), .Z(n756) );
  AND U551 ( .A(o[7]), .B(n766), .Z(n765) );
  XOR U552 ( .A(n764), .B(n767), .Z(n766) );
  XOR U553 ( .A(n768), .B(n769), .Z(n736) );
  AND U554 ( .A(o[5]), .B(n770), .Z(n769) );
  XNOR U555 ( .A(n771), .B(n772), .Z(n770) );
  XNOR U556 ( .A(n773), .B(n768), .Z(n772) );
  AND U557 ( .A(o[6]), .B(n774), .Z(n773) );
  XNOR U558 ( .A(n771), .B(n775), .Z(n774) );
  XNOR U559 ( .A(n776), .B(n777), .Z(n775) );
  AND U560 ( .A(o[7]), .B(n778), .Z(n776) );
  XOR U561 ( .A(n777), .B(n779), .Z(n778) );
  XOR U562 ( .A(n780), .B(n781), .Z(n771) );
  AND U563 ( .A(o[7]), .B(n782), .Z(n781) );
  XOR U564 ( .A(n780), .B(n783), .Z(n782) );
  XOR U565 ( .A(n784), .B(n785), .Z(n768) );
  AND U566 ( .A(o[6]), .B(n786), .Z(n785) );
  XNOR U567 ( .A(n784), .B(n787), .Z(n786) );
  XNOR U568 ( .A(n788), .B(n789), .Z(n787) );
  AND U569 ( .A(o[7]), .B(n790), .Z(n788) );
  XOR U570 ( .A(n789), .B(n791), .Z(n790) );
  XOR U571 ( .A(n792), .B(n793), .Z(n784) );
  AND U572 ( .A(o[7]), .B(n794), .Z(n793) );
  XOR U573 ( .A(n792), .B(n795), .Z(n794) );
  XOR U574 ( .A(n796), .B(n797), .Z(o[2]) );
  AND U575 ( .A(o[3]), .B(n798), .Z(n797) );
  XNOR U576 ( .A(n799), .B(n800), .Z(n798) );
  XNOR U577 ( .A(n801), .B(n796), .Z(n800) );
  AND U578 ( .A(o[4]), .B(n802), .Z(n801) );
  XNOR U579 ( .A(n803), .B(n804), .Z(n802) );
  XNOR U580 ( .A(n805), .B(n799), .Z(n804) );
  AND U581 ( .A(o[5]), .B(n806), .Z(n805) );
  XNOR U582 ( .A(n807), .B(n808), .Z(n806) );
  XNOR U583 ( .A(n809), .B(n803), .Z(n808) );
  AND U584 ( .A(o[6]), .B(n810), .Z(n809) );
  XNOR U585 ( .A(n807), .B(n811), .Z(n810) );
  XNOR U586 ( .A(n812), .B(n813), .Z(n811) );
  AND U587 ( .A(o[7]), .B(n814), .Z(n812) );
  XOR U588 ( .A(n813), .B(n815), .Z(n814) );
  XOR U589 ( .A(n816), .B(n817), .Z(n807) );
  AND U590 ( .A(o[7]), .B(n818), .Z(n817) );
  XOR U591 ( .A(n816), .B(n819), .Z(n818) );
  XOR U592 ( .A(n820), .B(n821), .Z(n803) );
  AND U593 ( .A(o[6]), .B(n822), .Z(n821) );
  XNOR U594 ( .A(n820), .B(n823), .Z(n822) );
  XNOR U595 ( .A(n824), .B(n825), .Z(n823) );
  AND U596 ( .A(o[7]), .B(n826), .Z(n824) );
  XOR U597 ( .A(n825), .B(n827), .Z(n826) );
  XOR U598 ( .A(n828), .B(n829), .Z(n820) );
  AND U599 ( .A(o[7]), .B(n830), .Z(n829) );
  XOR U600 ( .A(n828), .B(n831), .Z(n830) );
  XOR U601 ( .A(n832), .B(n833), .Z(n799) );
  AND U602 ( .A(o[5]), .B(n834), .Z(n833) );
  XNOR U603 ( .A(n835), .B(n836), .Z(n834) );
  XNOR U604 ( .A(n837), .B(n832), .Z(n836) );
  AND U605 ( .A(o[6]), .B(n838), .Z(n837) );
  XNOR U606 ( .A(n835), .B(n839), .Z(n838) );
  XNOR U607 ( .A(n840), .B(n841), .Z(n839) );
  AND U608 ( .A(o[7]), .B(n842), .Z(n840) );
  XOR U609 ( .A(n841), .B(n843), .Z(n842) );
  XOR U610 ( .A(n844), .B(n845), .Z(n835) );
  AND U611 ( .A(o[7]), .B(n846), .Z(n845) );
  XOR U612 ( .A(n844), .B(n847), .Z(n846) );
  XOR U613 ( .A(n848), .B(n849), .Z(n832) );
  AND U614 ( .A(o[6]), .B(n850), .Z(n849) );
  XNOR U615 ( .A(n848), .B(n851), .Z(n850) );
  XNOR U616 ( .A(n852), .B(n853), .Z(n851) );
  AND U617 ( .A(o[7]), .B(n854), .Z(n852) );
  XOR U618 ( .A(n853), .B(n855), .Z(n854) );
  XOR U619 ( .A(n856), .B(n857), .Z(n848) );
  AND U620 ( .A(o[7]), .B(n858), .Z(n857) );
  XOR U621 ( .A(n856), .B(n859), .Z(n858) );
  XOR U622 ( .A(n860), .B(n861), .Z(n796) );
  AND U623 ( .A(o[4]), .B(n862), .Z(n861) );
  XNOR U624 ( .A(n863), .B(n864), .Z(n862) );
  XNOR U625 ( .A(n865), .B(n860), .Z(n864) );
  AND U626 ( .A(o[5]), .B(n866), .Z(n865) );
  XNOR U627 ( .A(n867), .B(n868), .Z(n866) );
  XNOR U628 ( .A(n869), .B(n863), .Z(n868) );
  AND U629 ( .A(o[6]), .B(n870), .Z(n869) );
  XNOR U630 ( .A(n867), .B(n871), .Z(n870) );
  XNOR U631 ( .A(n872), .B(n873), .Z(n871) );
  AND U632 ( .A(o[7]), .B(n874), .Z(n872) );
  XOR U633 ( .A(n873), .B(n875), .Z(n874) );
  XOR U634 ( .A(n876), .B(n877), .Z(n867) );
  AND U635 ( .A(o[7]), .B(n878), .Z(n877) );
  XOR U636 ( .A(n876), .B(n879), .Z(n878) );
  XOR U637 ( .A(n880), .B(n881), .Z(n863) );
  AND U638 ( .A(o[6]), .B(n882), .Z(n881) );
  XNOR U639 ( .A(n880), .B(n883), .Z(n882) );
  XNOR U640 ( .A(n884), .B(n885), .Z(n883) );
  AND U641 ( .A(o[7]), .B(n886), .Z(n884) );
  XOR U642 ( .A(n885), .B(n887), .Z(n886) );
  XOR U643 ( .A(n888), .B(n889), .Z(n880) );
  AND U644 ( .A(o[7]), .B(n890), .Z(n889) );
  XOR U645 ( .A(n888), .B(n891), .Z(n890) );
  XOR U646 ( .A(n892), .B(n893), .Z(n860) );
  AND U647 ( .A(o[5]), .B(n894), .Z(n893) );
  XNOR U648 ( .A(n895), .B(n896), .Z(n894) );
  XNOR U649 ( .A(n897), .B(n892), .Z(n896) );
  AND U650 ( .A(o[6]), .B(n898), .Z(n897) );
  XNOR U651 ( .A(n895), .B(n899), .Z(n898) );
  XNOR U652 ( .A(n900), .B(n901), .Z(n899) );
  AND U653 ( .A(o[7]), .B(n902), .Z(n900) );
  XOR U654 ( .A(n901), .B(n903), .Z(n902) );
  XOR U655 ( .A(n904), .B(n905), .Z(n895) );
  AND U656 ( .A(o[7]), .B(n906), .Z(n905) );
  XOR U657 ( .A(n904), .B(n907), .Z(n906) );
  XOR U658 ( .A(n908), .B(n909), .Z(n892) );
  AND U659 ( .A(o[6]), .B(n910), .Z(n909) );
  XNOR U660 ( .A(n908), .B(n911), .Z(n910) );
  XNOR U661 ( .A(n912), .B(n913), .Z(n911) );
  AND U662 ( .A(o[7]), .B(n914), .Z(n912) );
  XOR U663 ( .A(n913), .B(n915), .Z(n914) );
  XOR U664 ( .A(n916), .B(n917), .Z(n908) );
  AND U665 ( .A(o[7]), .B(n918), .Z(n917) );
  XOR U666 ( .A(n916), .B(n919), .Z(n918) );
  XOR U667 ( .A(n920), .B(n921), .Z(n668) );
  AND U668 ( .A(o[3]), .B(n922), .Z(n921) );
  XNOR U669 ( .A(n923), .B(n924), .Z(n922) );
  XNOR U670 ( .A(n925), .B(n920), .Z(n924) );
  AND U671 ( .A(o[4]), .B(n926), .Z(n925) );
  XNOR U672 ( .A(n927), .B(n928), .Z(n926) );
  XNOR U673 ( .A(n929), .B(n923), .Z(n928) );
  AND U674 ( .A(o[5]), .B(n930), .Z(n929) );
  XNOR U675 ( .A(n931), .B(n932), .Z(n930) );
  XNOR U676 ( .A(n933), .B(n927), .Z(n932) );
  AND U677 ( .A(o[6]), .B(n934), .Z(n933) );
  XNOR U678 ( .A(n931), .B(n935), .Z(n934) );
  XNOR U679 ( .A(n936), .B(n937), .Z(n935) );
  AND U680 ( .A(o[7]), .B(n938), .Z(n936) );
  XOR U681 ( .A(n937), .B(n939), .Z(n938) );
  XOR U682 ( .A(n940), .B(n941), .Z(n931) );
  AND U683 ( .A(o[7]), .B(n942), .Z(n941) );
  XOR U684 ( .A(n940), .B(n943), .Z(n942) );
  XOR U685 ( .A(n944), .B(n945), .Z(n927) );
  AND U686 ( .A(o[6]), .B(n946), .Z(n945) );
  XNOR U687 ( .A(n944), .B(n947), .Z(n946) );
  XNOR U688 ( .A(n948), .B(n949), .Z(n947) );
  AND U689 ( .A(o[7]), .B(n950), .Z(n948) );
  XOR U690 ( .A(n949), .B(n951), .Z(n950) );
  XOR U691 ( .A(n952), .B(n953), .Z(n944) );
  AND U692 ( .A(o[7]), .B(n954), .Z(n953) );
  XOR U693 ( .A(n952), .B(n955), .Z(n954) );
  XOR U694 ( .A(n956), .B(n957), .Z(n923) );
  AND U695 ( .A(o[5]), .B(n958), .Z(n957) );
  XNOR U696 ( .A(n959), .B(n960), .Z(n958) );
  XNOR U697 ( .A(n961), .B(n956), .Z(n960) );
  AND U698 ( .A(o[6]), .B(n962), .Z(n961) );
  XNOR U699 ( .A(n959), .B(n963), .Z(n962) );
  XNOR U700 ( .A(n964), .B(n965), .Z(n963) );
  AND U701 ( .A(o[7]), .B(n966), .Z(n964) );
  XOR U702 ( .A(n965), .B(n967), .Z(n966) );
  XOR U703 ( .A(n968), .B(n969), .Z(n959) );
  AND U704 ( .A(o[7]), .B(n970), .Z(n969) );
  XOR U705 ( .A(n968), .B(n971), .Z(n970) );
  XOR U706 ( .A(n972), .B(n973), .Z(n956) );
  AND U707 ( .A(o[6]), .B(n974), .Z(n973) );
  XNOR U708 ( .A(n972), .B(n975), .Z(n974) );
  XNOR U709 ( .A(n976), .B(n977), .Z(n975) );
  AND U710 ( .A(o[7]), .B(n978), .Z(n976) );
  XOR U711 ( .A(n977), .B(n979), .Z(n978) );
  XOR U712 ( .A(n980), .B(n981), .Z(n972) );
  AND U713 ( .A(o[7]), .B(n982), .Z(n981) );
  XOR U714 ( .A(n980), .B(n983), .Z(n982) );
  XOR U715 ( .A(n984), .B(n985), .Z(o[3]) );
  AND U716 ( .A(o[4]), .B(n986), .Z(n985) );
  XNOR U717 ( .A(n987), .B(n988), .Z(n986) );
  XNOR U718 ( .A(n989), .B(n984), .Z(n988) );
  AND U719 ( .A(o[5]), .B(n990), .Z(n989) );
  XNOR U720 ( .A(n991), .B(n992), .Z(n990) );
  XNOR U721 ( .A(n993), .B(n987), .Z(n992) );
  AND U722 ( .A(o[6]), .B(n994), .Z(n993) );
  XNOR U723 ( .A(n991), .B(n995), .Z(n994) );
  XNOR U724 ( .A(n996), .B(n997), .Z(n995) );
  AND U725 ( .A(o[7]), .B(n998), .Z(n996) );
  XOR U726 ( .A(n997), .B(n999), .Z(n998) );
  XOR U727 ( .A(n1000), .B(n1001), .Z(n991) );
  AND U728 ( .A(o[7]), .B(n1002), .Z(n1001) );
  XOR U729 ( .A(n1000), .B(n1003), .Z(n1002) );
  XOR U730 ( .A(n1004), .B(n1005), .Z(n987) );
  AND U731 ( .A(o[6]), .B(n1006), .Z(n1005) );
  XNOR U732 ( .A(n1004), .B(n1007), .Z(n1006) );
  XNOR U733 ( .A(n1008), .B(n1009), .Z(n1007) );
  AND U734 ( .A(o[7]), .B(n1010), .Z(n1008) );
  XOR U735 ( .A(n1009), .B(n1011), .Z(n1010) );
  XOR U736 ( .A(n1012), .B(n1013), .Z(n1004) );
  AND U737 ( .A(o[7]), .B(n1014), .Z(n1013) );
  XOR U738 ( .A(n1012), .B(n1015), .Z(n1014) );
  XOR U739 ( .A(n1016), .B(n1017), .Z(n984) );
  AND U740 ( .A(o[5]), .B(n1018), .Z(n1017) );
  XNOR U741 ( .A(n1019), .B(n1020), .Z(n1018) );
  XNOR U742 ( .A(n1021), .B(n1016), .Z(n1020) );
  AND U743 ( .A(o[6]), .B(n1022), .Z(n1021) );
  XNOR U744 ( .A(n1019), .B(n1023), .Z(n1022) );
  XNOR U745 ( .A(n1024), .B(n1025), .Z(n1023) );
  AND U746 ( .A(o[7]), .B(n1026), .Z(n1024) );
  XOR U747 ( .A(n1025), .B(n1027), .Z(n1026) );
  XOR U748 ( .A(n1028), .B(n1029), .Z(n1019) );
  AND U749 ( .A(o[7]), .B(n1030), .Z(n1029) );
  XOR U750 ( .A(n1028), .B(n1031), .Z(n1030) );
  XOR U751 ( .A(n1032), .B(n1033), .Z(n1016) );
  AND U752 ( .A(o[6]), .B(n1034), .Z(n1033) );
  XNOR U753 ( .A(n1032), .B(n1035), .Z(n1034) );
  XNOR U754 ( .A(n1036), .B(n1037), .Z(n1035) );
  AND U755 ( .A(o[7]), .B(n1038), .Z(n1036) );
  XOR U756 ( .A(n1037), .B(n1039), .Z(n1038) );
  XOR U757 ( .A(n1040), .B(n1041), .Z(n1032) );
  AND U758 ( .A(o[7]), .B(n1042), .Z(n1041) );
  XOR U759 ( .A(n1040), .B(n1043), .Z(n1042) );
  XOR U760 ( .A(n1044), .B(n1045), .Z(n920) );
  AND U761 ( .A(o[4]), .B(n1046), .Z(n1045) );
  XNOR U762 ( .A(n1047), .B(n1048), .Z(n1046) );
  XNOR U763 ( .A(n1049), .B(n1044), .Z(n1048) );
  AND U764 ( .A(o[5]), .B(n1050), .Z(n1049) );
  XNOR U765 ( .A(n1051), .B(n1052), .Z(n1050) );
  XNOR U766 ( .A(n1053), .B(n1047), .Z(n1052) );
  AND U767 ( .A(o[6]), .B(n1054), .Z(n1053) );
  XNOR U768 ( .A(n1051), .B(n1055), .Z(n1054) );
  XNOR U769 ( .A(n1056), .B(n1057), .Z(n1055) );
  AND U770 ( .A(o[7]), .B(n1058), .Z(n1056) );
  XOR U771 ( .A(n1057), .B(n1059), .Z(n1058) );
  XOR U772 ( .A(n1060), .B(n1061), .Z(n1051) );
  AND U773 ( .A(o[7]), .B(n1062), .Z(n1061) );
  XOR U774 ( .A(n1060), .B(n1063), .Z(n1062) );
  XOR U775 ( .A(n1064), .B(n1065), .Z(n1047) );
  AND U776 ( .A(o[6]), .B(n1066), .Z(n1065) );
  XNOR U777 ( .A(n1064), .B(n1067), .Z(n1066) );
  XNOR U778 ( .A(n1068), .B(n1069), .Z(n1067) );
  AND U779 ( .A(o[7]), .B(n1070), .Z(n1068) );
  XOR U780 ( .A(n1069), .B(n1071), .Z(n1070) );
  XOR U781 ( .A(n1072), .B(n1073), .Z(n1064) );
  AND U782 ( .A(o[7]), .B(n1074), .Z(n1073) );
  XOR U783 ( .A(n1072), .B(n1075), .Z(n1074) );
  XOR U784 ( .A(n1076), .B(n1077), .Z(o[4]) );
  AND U785 ( .A(o[5]), .B(n1078), .Z(n1077) );
  XNOR U786 ( .A(n1079), .B(n1080), .Z(n1078) );
  XNOR U787 ( .A(n1081), .B(n1076), .Z(n1080) );
  AND U788 ( .A(o[6]), .B(n1082), .Z(n1081) );
  XNOR U789 ( .A(n1079), .B(n1083), .Z(n1082) );
  XNOR U790 ( .A(n1084), .B(n1085), .Z(n1083) );
  AND U791 ( .A(o[7]), .B(n1086), .Z(n1084) );
  XOR U792 ( .A(n1085), .B(n1087), .Z(n1086) );
  XOR U793 ( .A(n1088), .B(n1089), .Z(n1079) );
  AND U794 ( .A(o[7]), .B(n1090), .Z(n1089) );
  XOR U795 ( .A(n1088), .B(n1091), .Z(n1090) );
  XOR U796 ( .A(n1092), .B(n1093), .Z(n1076) );
  AND U797 ( .A(o[6]), .B(n1094), .Z(n1093) );
  XNOR U798 ( .A(n1092), .B(n1095), .Z(n1094) );
  XNOR U799 ( .A(n1096), .B(n1097), .Z(n1095) );
  AND U800 ( .A(o[7]), .B(n1098), .Z(n1096) );
  XOR U801 ( .A(n1097), .B(n1099), .Z(n1098) );
  XOR U802 ( .A(n1100), .B(n1101), .Z(n1092) );
  AND U803 ( .A(o[7]), .B(n1102), .Z(n1101) );
  XOR U804 ( .A(n1100), .B(n1103), .Z(n1102) );
  XOR U805 ( .A(n1104), .B(n1105), .Z(n1044) );
  AND U806 ( .A(o[5]), .B(n1106), .Z(n1105) );
  XNOR U807 ( .A(n1107), .B(n1108), .Z(n1106) );
  XNOR U808 ( .A(n1109), .B(n1104), .Z(n1108) );
  AND U809 ( .A(o[6]), .B(n1110), .Z(n1109) );
  XNOR U810 ( .A(n1107), .B(n1111), .Z(n1110) );
  XNOR U811 ( .A(n1112), .B(n1113), .Z(n1111) );
  AND U812 ( .A(o[7]), .B(n1114), .Z(n1112) );
  XOR U813 ( .A(n1113), .B(n1115), .Z(n1114) );
  XOR U814 ( .A(n1116), .B(n1117), .Z(n1107) );
  AND U815 ( .A(o[7]), .B(n1118), .Z(n1117) );
  XOR U816 ( .A(n1116), .B(n1119), .Z(n1118) );
  XOR U817 ( .A(n1120), .B(n1121), .Z(o[5]) );
  AND U818 ( .A(o[6]), .B(n1122), .Z(n1121) );
  XNOR U819 ( .A(n1120), .B(n1123), .Z(n1122) );
  XNOR U820 ( .A(n1124), .B(n1125), .Z(n1123) );
  AND U821 ( .A(o[7]), .B(n1126), .Z(n1124) );
  XOR U822 ( .A(n1125), .B(n1127), .Z(n1126) );
  XOR U823 ( .A(n1128), .B(n1129), .Z(n1120) );
  AND U824 ( .A(o[7]), .B(n1130), .Z(n1129) );
  XOR U825 ( .A(n1128), .B(n1131), .Z(n1130) );
  XOR U826 ( .A(n1132), .B(n1133), .Z(n1104) );
  AND U827 ( .A(o[6]), .B(n1134), .Z(n1133) );
  XNOR U828 ( .A(n1132), .B(n1135), .Z(n1134) );
  XNOR U829 ( .A(n1136), .B(n1137), .Z(n1135) );
  AND U830 ( .A(o[7]), .B(n1138), .Z(n1136) );
  XOR U831 ( .A(n1137), .B(n1139), .Z(n1138) );
  XOR U832 ( .A(n1140), .B(n1141), .Z(o[6]) );
  AND U833 ( .A(o[7]), .B(n1142), .Z(n1141) );
  XOR U834 ( .A(n1140), .B(n1143), .Z(n1142) );
  XOR U835 ( .A(n1144), .B(n1145), .Z(n1132) );
  AND U836 ( .A(o[7]), .B(n1146), .Z(n1145) );
  XOR U837 ( .A(n1144), .B(n1147), .Z(n1146) );
  XOR U838 ( .A(n1148), .B(n1149), .Z(o[7]) );
  AND U839 ( .A(n1150), .B(n1151), .Z(n1149) );
  XOR U840 ( .A(n1148), .B(n13), .Z(n1151) );
  XOR U841 ( .A(n1152), .B(n1153), .Z(n13) );
  AND U842 ( .A(n1143), .B(n1154), .Z(n1153) );
  XOR U843 ( .A(n1155), .B(n1152), .Z(n1154) );
  XNOR U844 ( .A(n14), .B(n1148), .Z(n1150) );
  IV U845 ( .A(n11), .Z(n14) );
  XNOR U846 ( .A(n1156), .B(n1157), .Z(n11) );
  AND U847 ( .A(n1140), .B(n1158), .Z(n1157) );
  XOR U848 ( .A(n1159), .B(n1156), .Z(n1158) );
  XOR U849 ( .A(n1160), .B(n1161), .Z(n1148) );
  AND U850 ( .A(n1162), .B(n1163), .Z(n1161) );
  XOR U851 ( .A(n1160), .B(n18), .Z(n1163) );
  XOR U852 ( .A(n1164), .B(n1165), .Z(n18) );
  AND U853 ( .A(n1143), .B(n1166), .Z(n1165) );
  XOR U854 ( .A(n1167), .B(n1164), .Z(n1166) );
  XNOR U855 ( .A(n19), .B(n1160), .Z(n1162) );
  IV U856 ( .A(n16), .Z(n19) );
  XNOR U857 ( .A(n1168), .B(n1169), .Z(n16) );
  AND U858 ( .A(n1140), .B(n1170), .Z(n1169) );
  XOR U859 ( .A(n1171), .B(n1168), .Z(n1170) );
  XOR U860 ( .A(n1172), .B(n1173), .Z(n1160) );
  AND U861 ( .A(n1174), .B(n1175), .Z(n1173) );
  XOR U862 ( .A(n1172), .B(n23), .Z(n1175) );
  XOR U863 ( .A(n1176), .B(n1177), .Z(n23) );
  AND U864 ( .A(n1143), .B(n1178), .Z(n1177) );
  XOR U865 ( .A(n1179), .B(n1176), .Z(n1178) );
  XNOR U866 ( .A(n24), .B(n1172), .Z(n1174) );
  IV U867 ( .A(n21), .Z(n24) );
  XNOR U868 ( .A(n1180), .B(n1181), .Z(n21) );
  AND U869 ( .A(n1140), .B(n1182), .Z(n1181) );
  XOR U870 ( .A(n1183), .B(n1180), .Z(n1182) );
  XOR U871 ( .A(n1184), .B(n1185), .Z(n1172) );
  AND U872 ( .A(n1186), .B(n1187), .Z(n1185) );
  XOR U873 ( .A(n1184), .B(n28), .Z(n1187) );
  XOR U874 ( .A(n1188), .B(n1189), .Z(n28) );
  AND U875 ( .A(n1143), .B(n1190), .Z(n1189) );
  XOR U876 ( .A(n1191), .B(n1188), .Z(n1190) );
  XNOR U877 ( .A(n29), .B(n1184), .Z(n1186) );
  IV U878 ( .A(n26), .Z(n29) );
  XNOR U879 ( .A(n1192), .B(n1193), .Z(n26) );
  AND U880 ( .A(n1140), .B(n1194), .Z(n1193) );
  XOR U881 ( .A(n1195), .B(n1192), .Z(n1194) );
  XOR U882 ( .A(n1196), .B(n1197), .Z(n1184) );
  AND U883 ( .A(n1198), .B(n1199), .Z(n1197) );
  XOR U884 ( .A(n1196), .B(n33), .Z(n1199) );
  XOR U885 ( .A(n1200), .B(n1201), .Z(n33) );
  AND U886 ( .A(n1143), .B(n1202), .Z(n1201) );
  XOR U887 ( .A(n1203), .B(n1200), .Z(n1202) );
  XNOR U888 ( .A(n34), .B(n1196), .Z(n1198) );
  IV U889 ( .A(n31), .Z(n34) );
  XNOR U890 ( .A(n1204), .B(n1205), .Z(n31) );
  AND U891 ( .A(n1140), .B(n1206), .Z(n1205) );
  XOR U892 ( .A(n1207), .B(n1204), .Z(n1206) );
  XOR U893 ( .A(n1208), .B(n1209), .Z(n1196) );
  AND U894 ( .A(n1210), .B(n1211), .Z(n1209) );
  XOR U895 ( .A(n1208), .B(n38), .Z(n1211) );
  XOR U896 ( .A(n1212), .B(n1213), .Z(n38) );
  AND U897 ( .A(n1143), .B(n1214), .Z(n1213) );
  XOR U898 ( .A(n1215), .B(n1212), .Z(n1214) );
  XNOR U899 ( .A(n39), .B(n1208), .Z(n1210) );
  IV U900 ( .A(n36), .Z(n39) );
  XNOR U901 ( .A(n1216), .B(n1217), .Z(n36) );
  AND U902 ( .A(n1140), .B(n1218), .Z(n1217) );
  XOR U903 ( .A(n1219), .B(n1216), .Z(n1218) );
  XOR U904 ( .A(n1220), .B(n1221), .Z(n1208) );
  AND U905 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U906 ( .A(n1220), .B(n43), .Z(n1223) );
  XOR U907 ( .A(n1224), .B(n1225), .Z(n43) );
  AND U908 ( .A(n1143), .B(n1226), .Z(n1225) );
  XOR U909 ( .A(n1227), .B(n1224), .Z(n1226) );
  XNOR U910 ( .A(n44), .B(n1220), .Z(n1222) );
  IV U911 ( .A(n41), .Z(n44) );
  XNOR U912 ( .A(n1228), .B(n1229), .Z(n41) );
  AND U913 ( .A(n1140), .B(n1230), .Z(n1229) );
  XOR U914 ( .A(n1231), .B(n1228), .Z(n1230) );
  XOR U915 ( .A(n1232), .B(n1233), .Z(n1220) );
  AND U916 ( .A(n1234), .B(n1235), .Z(n1233) );
  XOR U917 ( .A(n1232), .B(n48), .Z(n1235) );
  XOR U918 ( .A(n1236), .B(n1237), .Z(n48) );
  AND U919 ( .A(n1143), .B(n1238), .Z(n1237) );
  XOR U920 ( .A(n1239), .B(n1236), .Z(n1238) );
  XNOR U921 ( .A(n49), .B(n1232), .Z(n1234) );
  IV U922 ( .A(n46), .Z(n49) );
  XNOR U923 ( .A(n1240), .B(n1241), .Z(n46) );
  AND U924 ( .A(n1140), .B(n1242), .Z(n1241) );
  XOR U925 ( .A(n1243), .B(n1240), .Z(n1242) );
  XOR U926 ( .A(n1244), .B(n1245), .Z(n1232) );
  AND U927 ( .A(n1246), .B(n1247), .Z(n1245) );
  XOR U928 ( .A(n1244), .B(n53), .Z(n1247) );
  XOR U929 ( .A(n1248), .B(n1249), .Z(n53) );
  AND U930 ( .A(n1143), .B(n1250), .Z(n1249) );
  XOR U931 ( .A(n1251), .B(n1248), .Z(n1250) );
  XNOR U932 ( .A(n54), .B(n1244), .Z(n1246) );
  IV U933 ( .A(n51), .Z(n54) );
  XNOR U934 ( .A(n1252), .B(n1253), .Z(n51) );
  AND U935 ( .A(n1140), .B(n1254), .Z(n1253) );
  XOR U936 ( .A(n1255), .B(n1252), .Z(n1254) );
  XOR U937 ( .A(n1256), .B(n1257), .Z(n1244) );
  AND U938 ( .A(n1258), .B(n1259), .Z(n1257) );
  XOR U939 ( .A(n1256), .B(n58), .Z(n1259) );
  XOR U940 ( .A(n1260), .B(n1261), .Z(n58) );
  AND U941 ( .A(n1143), .B(n1262), .Z(n1261) );
  XOR U942 ( .A(n1263), .B(n1260), .Z(n1262) );
  XNOR U943 ( .A(n59), .B(n1256), .Z(n1258) );
  IV U944 ( .A(n56), .Z(n59) );
  XNOR U945 ( .A(n1264), .B(n1265), .Z(n56) );
  AND U946 ( .A(n1140), .B(n1266), .Z(n1265) );
  XOR U947 ( .A(n1267), .B(n1264), .Z(n1266) );
  XOR U948 ( .A(n1268), .B(n1269), .Z(n1256) );
  AND U949 ( .A(n1270), .B(n1271), .Z(n1269) );
  XOR U950 ( .A(n1268), .B(n63), .Z(n1271) );
  XOR U951 ( .A(n1272), .B(n1273), .Z(n63) );
  AND U952 ( .A(n1143), .B(n1274), .Z(n1273) );
  XOR U953 ( .A(n1275), .B(n1272), .Z(n1274) );
  XNOR U954 ( .A(n64), .B(n1268), .Z(n1270) );
  IV U955 ( .A(n61), .Z(n64) );
  XNOR U956 ( .A(n1276), .B(n1277), .Z(n61) );
  AND U957 ( .A(n1140), .B(n1278), .Z(n1277) );
  XOR U958 ( .A(n1279), .B(n1276), .Z(n1278) );
  XOR U959 ( .A(n1280), .B(n1281), .Z(n1268) );
  AND U960 ( .A(n1282), .B(n1283), .Z(n1281) );
  XOR U961 ( .A(n1280), .B(n68), .Z(n1283) );
  XOR U962 ( .A(n1284), .B(n1285), .Z(n68) );
  AND U963 ( .A(n1143), .B(n1286), .Z(n1285) );
  XOR U964 ( .A(n1287), .B(n1284), .Z(n1286) );
  XNOR U965 ( .A(n69), .B(n1280), .Z(n1282) );
  IV U966 ( .A(n66), .Z(n69) );
  XNOR U967 ( .A(n1288), .B(n1289), .Z(n66) );
  AND U968 ( .A(n1140), .B(n1290), .Z(n1289) );
  XOR U969 ( .A(n1291), .B(n1288), .Z(n1290) );
  XOR U970 ( .A(n1292), .B(n1293), .Z(n1280) );
  AND U971 ( .A(n1294), .B(n1295), .Z(n1293) );
  XOR U972 ( .A(n1292), .B(n73), .Z(n1295) );
  XOR U973 ( .A(n1296), .B(n1297), .Z(n73) );
  AND U974 ( .A(n1143), .B(n1298), .Z(n1297) );
  XOR U975 ( .A(n1299), .B(n1296), .Z(n1298) );
  XNOR U976 ( .A(n74), .B(n1292), .Z(n1294) );
  IV U977 ( .A(n71), .Z(n74) );
  XNOR U978 ( .A(n1300), .B(n1301), .Z(n71) );
  AND U979 ( .A(n1140), .B(n1302), .Z(n1301) );
  XOR U980 ( .A(n1303), .B(n1300), .Z(n1302) );
  XOR U981 ( .A(n1304), .B(n1305), .Z(n1292) );
  AND U982 ( .A(n1306), .B(n1307), .Z(n1305) );
  XOR U983 ( .A(n1304), .B(n78), .Z(n1307) );
  XOR U984 ( .A(n1308), .B(n1309), .Z(n78) );
  AND U985 ( .A(n1143), .B(n1310), .Z(n1309) );
  XOR U986 ( .A(n1311), .B(n1308), .Z(n1310) );
  XNOR U987 ( .A(n79), .B(n1304), .Z(n1306) );
  IV U988 ( .A(n76), .Z(n79) );
  XNOR U989 ( .A(n1312), .B(n1313), .Z(n76) );
  AND U990 ( .A(n1140), .B(n1314), .Z(n1313) );
  XOR U991 ( .A(n1315), .B(n1312), .Z(n1314) );
  XOR U992 ( .A(n1316), .B(n1317), .Z(n1304) );
  AND U993 ( .A(n1318), .B(n1319), .Z(n1317) );
  XOR U994 ( .A(n1316), .B(n83), .Z(n1319) );
  XOR U995 ( .A(n1320), .B(n1321), .Z(n83) );
  AND U996 ( .A(n1143), .B(n1322), .Z(n1321) );
  XOR U997 ( .A(n1323), .B(n1320), .Z(n1322) );
  XNOR U998 ( .A(n84), .B(n1316), .Z(n1318) );
  IV U999 ( .A(n81), .Z(n84) );
  XNOR U1000 ( .A(n1324), .B(n1325), .Z(n81) );
  AND U1001 ( .A(n1140), .B(n1326), .Z(n1325) );
  XOR U1002 ( .A(n1327), .B(n1324), .Z(n1326) );
  XOR U1003 ( .A(n1328), .B(n1329), .Z(n1316) );
  AND U1004 ( .A(n1330), .B(n1331), .Z(n1329) );
  XOR U1005 ( .A(n1328), .B(n88), .Z(n1331) );
  XOR U1006 ( .A(n1332), .B(n1333), .Z(n88) );
  AND U1007 ( .A(n1143), .B(n1334), .Z(n1333) );
  XOR U1008 ( .A(n1335), .B(n1332), .Z(n1334) );
  XNOR U1009 ( .A(n89), .B(n1328), .Z(n1330) );
  IV U1010 ( .A(n86), .Z(n89) );
  XNOR U1011 ( .A(n1336), .B(n1337), .Z(n86) );
  AND U1012 ( .A(n1140), .B(n1338), .Z(n1337) );
  XOR U1013 ( .A(n1339), .B(n1336), .Z(n1338) );
  XOR U1014 ( .A(n1340), .B(n1341), .Z(n1328) );
  AND U1015 ( .A(n1342), .B(n1343), .Z(n1341) );
  XOR U1016 ( .A(n1340), .B(n93), .Z(n1343) );
  XOR U1017 ( .A(n1344), .B(n1345), .Z(n93) );
  AND U1018 ( .A(n1143), .B(n1346), .Z(n1345) );
  XOR U1019 ( .A(n1347), .B(n1344), .Z(n1346) );
  XNOR U1020 ( .A(n94), .B(n1340), .Z(n1342) );
  IV U1021 ( .A(n91), .Z(n94) );
  XNOR U1022 ( .A(n1348), .B(n1349), .Z(n91) );
  AND U1023 ( .A(n1140), .B(n1350), .Z(n1349) );
  XOR U1024 ( .A(n1351), .B(n1348), .Z(n1350) );
  XOR U1025 ( .A(n1352), .B(n1353), .Z(n1340) );
  AND U1026 ( .A(n1354), .B(n1355), .Z(n1353) );
  XOR U1027 ( .A(n1352), .B(n98), .Z(n1355) );
  XOR U1028 ( .A(n1356), .B(n1357), .Z(n98) );
  AND U1029 ( .A(n1143), .B(n1358), .Z(n1357) );
  XOR U1030 ( .A(n1359), .B(n1356), .Z(n1358) );
  XNOR U1031 ( .A(n99), .B(n1352), .Z(n1354) );
  IV U1032 ( .A(n96), .Z(n99) );
  XNOR U1033 ( .A(n1360), .B(n1361), .Z(n96) );
  AND U1034 ( .A(n1140), .B(n1362), .Z(n1361) );
  XOR U1035 ( .A(n1363), .B(n1360), .Z(n1362) );
  XOR U1036 ( .A(n1364), .B(n1365), .Z(n1352) );
  AND U1037 ( .A(n1366), .B(n1367), .Z(n1365) );
  XOR U1038 ( .A(n1364), .B(n103), .Z(n1367) );
  XOR U1039 ( .A(n1368), .B(n1369), .Z(n103) );
  AND U1040 ( .A(n1143), .B(n1370), .Z(n1369) );
  XOR U1041 ( .A(n1371), .B(n1368), .Z(n1370) );
  XNOR U1042 ( .A(n104), .B(n1364), .Z(n1366) );
  IV U1043 ( .A(n101), .Z(n104) );
  XNOR U1044 ( .A(n1372), .B(n1373), .Z(n101) );
  AND U1045 ( .A(n1140), .B(n1374), .Z(n1373) );
  XOR U1046 ( .A(n1375), .B(n1372), .Z(n1374) );
  XOR U1047 ( .A(n1376), .B(n1377), .Z(n1364) );
  AND U1048 ( .A(n1378), .B(n1379), .Z(n1377) );
  XOR U1049 ( .A(n1376), .B(n108), .Z(n1379) );
  XOR U1050 ( .A(n1380), .B(n1381), .Z(n108) );
  AND U1051 ( .A(n1143), .B(n1382), .Z(n1381) );
  XOR U1052 ( .A(n1383), .B(n1380), .Z(n1382) );
  XNOR U1053 ( .A(n109), .B(n1376), .Z(n1378) );
  IV U1054 ( .A(n106), .Z(n109) );
  XNOR U1055 ( .A(n1384), .B(n1385), .Z(n106) );
  AND U1056 ( .A(n1140), .B(n1386), .Z(n1385) );
  XOR U1057 ( .A(n1387), .B(n1384), .Z(n1386) );
  XOR U1058 ( .A(n1388), .B(n1389), .Z(n1376) );
  AND U1059 ( .A(n1390), .B(n1391), .Z(n1389) );
  XOR U1060 ( .A(n1388), .B(n113), .Z(n1391) );
  XOR U1061 ( .A(n1392), .B(n1393), .Z(n113) );
  AND U1062 ( .A(n1143), .B(n1394), .Z(n1393) );
  XOR U1063 ( .A(n1395), .B(n1392), .Z(n1394) );
  XNOR U1064 ( .A(n114), .B(n1388), .Z(n1390) );
  IV U1065 ( .A(n111), .Z(n114) );
  XNOR U1066 ( .A(n1396), .B(n1397), .Z(n111) );
  AND U1067 ( .A(n1140), .B(n1398), .Z(n1397) );
  XOR U1068 ( .A(n1399), .B(n1396), .Z(n1398) );
  XOR U1069 ( .A(n1400), .B(n1401), .Z(n1388) );
  AND U1070 ( .A(n1402), .B(n1403), .Z(n1401) );
  XOR U1071 ( .A(n1400), .B(n118), .Z(n1403) );
  XOR U1072 ( .A(n1404), .B(n1405), .Z(n118) );
  AND U1073 ( .A(n1143), .B(n1406), .Z(n1405) );
  XOR U1074 ( .A(n1407), .B(n1404), .Z(n1406) );
  XNOR U1075 ( .A(n119), .B(n1400), .Z(n1402) );
  IV U1076 ( .A(n116), .Z(n119) );
  XNOR U1077 ( .A(n1408), .B(n1409), .Z(n116) );
  AND U1078 ( .A(n1140), .B(n1410), .Z(n1409) );
  XOR U1079 ( .A(n1411), .B(n1408), .Z(n1410) );
  XOR U1080 ( .A(n1412), .B(n1413), .Z(n1400) );
  AND U1081 ( .A(n1414), .B(n1415), .Z(n1413) );
  XOR U1082 ( .A(n1412), .B(n123), .Z(n1415) );
  XOR U1083 ( .A(n1416), .B(n1417), .Z(n123) );
  AND U1084 ( .A(n1143), .B(n1418), .Z(n1417) );
  XOR U1085 ( .A(n1419), .B(n1416), .Z(n1418) );
  XNOR U1086 ( .A(n124), .B(n1412), .Z(n1414) );
  IV U1087 ( .A(n121), .Z(n124) );
  XNOR U1088 ( .A(n1420), .B(n1421), .Z(n121) );
  AND U1089 ( .A(n1140), .B(n1422), .Z(n1421) );
  XOR U1090 ( .A(n1423), .B(n1420), .Z(n1422) );
  XOR U1091 ( .A(n1424), .B(n1425), .Z(n1412) );
  AND U1092 ( .A(n1426), .B(n1427), .Z(n1425) );
  XOR U1093 ( .A(n1424), .B(n128), .Z(n1427) );
  XOR U1094 ( .A(n1428), .B(n1429), .Z(n128) );
  AND U1095 ( .A(n1143), .B(n1430), .Z(n1429) );
  XOR U1096 ( .A(n1431), .B(n1428), .Z(n1430) );
  XNOR U1097 ( .A(n129), .B(n1424), .Z(n1426) );
  IV U1098 ( .A(n126), .Z(n129) );
  XNOR U1099 ( .A(n1432), .B(n1433), .Z(n126) );
  AND U1100 ( .A(n1140), .B(n1434), .Z(n1433) );
  XOR U1101 ( .A(n1435), .B(n1432), .Z(n1434) );
  XOR U1102 ( .A(n1436), .B(n1437), .Z(n1424) );
  AND U1103 ( .A(n1438), .B(n1439), .Z(n1437) );
  XOR U1104 ( .A(n1436), .B(n133), .Z(n1439) );
  XOR U1105 ( .A(n1440), .B(n1441), .Z(n133) );
  AND U1106 ( .A(n1143), .B(n1442), .Z(n1441) );
  XOR U1107 ( .A(n1443), .B(n1440), .Z(n1442) );
  XNOR U1108 ( .A(n134), .B(n1436), .Z(n1438) );
  IV U1109 ( .A(n131), .Z(n134) );
  XNOR U1110 ( .A(n1444), .B(n1445), .Z(n131) );
  AND U1111 ( .A(n1140), .B(n1446), .Z(n1445) );
  XOR U1112 ( .A(n1447), .B(n1444), .Z(n1446) );
  XOR U1113 ( .A(n1448), .B(n1449), .Z(n1436) );
  AND U1114 ( .A(n1450), .B(n1451), .Z(n1449) );
  XOR U1115 ( .A(n1448), .B(n138), .Z(n1451) );
  XOR U1116 ( .A(n1452), .B(n1453), .Z(n138) );
  AND U1117 ( .A(n1143), .B(n1454), .Z(n1453) );
  XOR U1118 ( .A(n1455), .B(n1452), .Z(n1454) );
  XNOR U1119 ( .A(n139), .B(n1448), .Z(n1450) );
  IV U1120 ( .A(n136), .Z(n139) );
  XNOR U1121 ( .A(n1456), .B(n1457), .Z(n136) );
  AND U1122 ( .A(n1140), .B(n1458), .Z(n1457) );
  XOR U1123 ( .A(n1459), .B(n1456), .Z(n1458) );
  XOR U1124 ( .A(n1460), .B(n1461), .Z(n1448) );
  AND U1125 ( .A(n1462), .B(n1463), .Z(n1461) );
  XOR U1126 ( .A(n1460), .B(n143), .Z(n1463) );
  XOR U1127 ( .A(n1464), .B(n1465), .Z(n143) );
  AND U1128 ( .A(n1143), .B(n1466), .Z(n1465) );
  XOR U1129 ( .A(n1467), .B(n1464), .Z(n1466) );
  XNOR U1130 ( .A(n144), .B(n1460), .Z(n1462) );
  IV U1131 ( .A(n141), .Z(n144) );
  XNOR U1132 ( .A(n1468), .B(n1469), .Z(n141) );
  AND U1133 ( .A(n1140), .B(n1470), .Z(n1469) );
  XOR U1134 ( .A(n1471), .B(n1468), .Z(n1470) );
  XOR U1135 ( .A(n1472), .B(n1473), .Z(n1460) );
  AND U1136 ( .A(n1474), .B(n1475), .Z(n1473) );
  XOR U1137 ( .A(n1472), .B(n148), .Z(n1475) );
  XOR U1138 ( .A(n1476), .B(n1477), .Z(n148) );
  AND U1139 ( .A(n1143), .B(n1478), .Z(n1477) );
  XOR U1140 ( .A(n1479), .B(n1476), .Z(n1478) );
  XNOR U1141 ( .A(n149), .B(n1472), .Z(n1474) );
  IV U1142 ( .A(n146), .Z(n149) );
  XNOR U1143 ( .A(n1480), .B(n1481), .Z(n146) );
  AND U1144 ( .A(n1140), .B(n1482), .Z(n1481) );
  XOR U1145 ( .A(n1483), .B(n1480), .Z(n1482) );
  XOR U1146 ( .A(n1484), .B(n1485), .Z(n1472) );
  AND U1147 ( .A(n1486), .B(n1487), .Z(n1485) );
  XOR U1148 ( .A(n1484), .B(n153), .Z(n1487) );
  XOR U1149 ( .A(n1488), .B(n1489), .Z(n153) );
  AND U1150 ( .A(n1143), .B(n1490), .Z(n1489) );
  XOR U1151 ( .A(n1491), .B(n1488), .Z(n1490) );
  XNOR U1152 ( .A(n154), .B(n1484), .Z(n1486) );
  IV U1153 ( .A(n151), .Z(n154) );
  XNOR U1154 ( .A(n1492), .B(n1493), .Z(n151) );
  AND U1155 ( .A(n1140), .B(n1494), .Z(n1493) );
  XOR U1156 ( .A(n1495), .B(n1492), .Z(n1494) );
  XOR U1157 ( .A(n1496), .B(n1497), .Z(n1484) );
  AND U1158 ( .A(n1498), .B(n1499), .Z(n1497) );
  XOR U1159 ( .A(n1496), .B(n158), .Z(n1499) );
  XOR U1160 ( .A(n1500), .B(n1501), .Z(n158) );
  AND U1161 ( .A(n1143), .B(n1502), .Z(n1501) );
  XOR U1162 ( .A(n1503), .B(n1500), .Z(n1502) );
  XNOR U1163 ( .A(n159), .B(n1496), .Z(n1498) );
  IV U1164 ( .A(n156), .Z(n159) );
  XNOR U1165 ( .A(n1504), .B(n1505), .Z(n156) );
  AND U1166 ( .A(n1140), .B(n1506), .Z(n1505) );
  XOR U1167 ( .A(n1507), .B(n1504), .Z(n1506) );
  XNOR U1168 ( .A(n1508), .B(n1509), .Z(n1496) );
  AND U1169 ( .A(n1510), .B(n1511), .Z(n1509) );
  XNOR U1170 ( .A(n1508), .B(n5), .Z(n1511) );
  XOR U1171 ( .A(n1512), .B(n1513), .Z(n5) );
  AND U1172 ( .A(n1143), .B(n1514), .Z(n1513) );
  XOR U1173 ( .A(n1512), .B(n1515), .Z(n1514) );
  XOR U1174 ( .A(n4), .B(n1508), .Z(n1510) );
  IV U1175 ( .A(n2), .Z(n4) );
  XNOR U1176 ( .A(n1516), .B(n1517), .Z(n2) );
  AND U1177 ( .A(n1140), .B(n1518), .Z(n1517) );
  XOR U1178 ( .A(n1516), .B(n1519), .Z(n1518) );
  AND U1179 ( .A(n7), .B(n9), .Z(n1508) );
  XNOR U1180 ( .A(n1520), .B(n1521), .Z(n9) );
  AND U1181 ( .A(n1143), .B(n1522), .Z(n1521) );
  XNOR U1182 ( .A(n1523), .B(n1520), .Z(n1522) );
  XOR U1183 ( .A(n1524), .B(n1525), .Z(n1143) );
  AND U1184 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U1185 ( .A(n1524), .B(n1155), .Z(n1527) );
  XOR U1186 ( .A(n1528), .B(n1529), .Z(n1155) );
  AND U1187 ( .A(n1127), .B(n1530), .Z(n1529) );
  XOR U1188 ( .A(n1531), .B(n1528), .Z(n1530) );
  XNOR U1189 ( .A(n1152), .B(n1524), .Z(n1526) );
  XOR U1190 ( .A(n1532), .B(n1533), .Z(n1152) );
  AND U1191 ( .A(n1125), .B(n1534), .Z(n1533) );
  XOR U1192 ( .A(n1535), .B(n1532), .Z(n1534) );
  XOR U1193 ( .A(n1536), .B(n1537), .Z(n1524) );
  AND U1194 ( .A(n1538), .B(n1539), .Z(n1537) );
  XOR U1195 ( .A(n1536), .B(n1167), .Z(n1539) );
  XOR U1196 ( .A(n1540), .B(n1541), .Z(n1167) );
  AND U1197 ( .A(n1127), .B(n1542), .Z(n1541) );
  XOR U1198 ( .A(n1543), .B(n1540), .Z(n1542) );
  XNOR U1199 ( .A(n1164), .B(n1536), .Z(n1538) );
  XOR U1200 ( .A(n1544), .B(n1545), .Z(n1164) );
  AND U1201 ( .A(n1125), .B(n1546), .Z(n1545) );
  XOR U1202 ( .A(n1547), .B(n1544), .Z(n1546) );
  XOR U1203 ( .A(n1548), .B(n1549), .Z(n1536) );
  AND U1204 ( .A(n1550), .B(n1551), .Z(n1549) );
  XOR U1205 ( .A(n1548), .B(n1179), .Z(n1551) );
  XOR U1206 ( .A(n1552), .B(n1553), .Z(n1179) );
  AND U1207 ( .A(n1127), .B(n1554), .Z(n1553) );
  XOR U1208 ( .A(n1555), .B(n1552), .Z(n1554) );
  XNOR U1209 ( .A(n1176), .B(n1548), .Z(n1550) );
  XOR U1210 ( .A(n1556), .B(n1557), .Z(n1176) );
  AND U1211 ( .A(n1125), .B(n1558), .Z(n1557) );
  XOR U1212 ( .A(n1559), .B(n1556), .Z(n1558) );
  XOR U1213 ( .A(n1560), .B(n1561), .Z(n1548) );
  AND U1214 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U1215 ( .A(n1560), .B(n1191), .Z(n1563) );
  XOR U1216 ( .A(n1564), .B(n1565), .Z(n1191) );
  AND U1217 ( .A(n1127), .B(n1566), .Z(n1565) );
  XOR U1218 ( .A(n1567), .B(n1564), .Z(n1566) );
  XNOR U1219 ( .A(n1188), .B(n1560), .Z(n1562) );
  XOR U1220 ( .A(n1568), .B(n1569), .Z(n1188) );
  AND U1221 ( .A(n1125), .B(n1570), .Z(n1569) );
  XOR U1222 ( .A(n1571), .B(n1568), .Z(n1570) );
  XOR U1223 ( .A(n1572), .B(n1573), .Z(n1560) );
  AND U1224 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U1225 ( .A(n1572), .B(n1203), .Z(n1575) );
  XOR U1226 ( .A(n1576), .B(n1577), .Z(n1203) );
  AND U1227 ( .A(n1127), .B(n1578), .Z(n1577) );
  XOR U1228 ( .A(n1579), .B(n1576), .Z(n1578) );
  XNOR U1229 ( .A(n1200), .B(n1572), .Z(n1574) );
  XOR U1230 ( .A(n1580), .B(n1581), .Z(n1200) );
  AND U1231 ( .A(n1125), .B(n1582), .Z(n1581) );
  XOR U1232 ( .A(n1583), .B(n1580), .Z(n1582) );
  XOR U1233 ( .A(n1584), .B(n1585), .Z(n1572) );
  AND U1234 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U1235 ( .A(n1584), .B(n1215), .Z(n1587) );
  XOR U1236 ( .A(n1588), .B(n1589), .Z(n1215) );
  AND U1237 ( .A(n1127), .B(n1590), .Z(n1589) );
  XOR U1238 ( .A(n1591), .B(n1588), .Z(n1590) );
  XNOR U1239 ( .A(n1212), .B(n1584), .Z(n1586) );
  XOR U1240 ( .A(n1592), .B(n1593), .Z(n1212) );
  AND U1241 ( .A(n1125), .B(n1594), .Z(n1593) );
  XOR U1242 ( .A(n1595), .B(n1592), .Z(n1594) );
  XOR U1243 ( .A(n1596), .B(n1597), .Z(n1584) );
  AND U1244 ( .A(n1598), .B(n1599), .Z(n1597) );
  XOR U1245 ( .A(n1596), .B(n1227), .Z(n1599) );
  XOR U1246 ( .A(n1600), .B(n1601), .Z(n1227) );
  AND U1247 ( .A(n1127), .B(n1602), .Z(n1601) );
  XOR U1248 ( .A(n1603), .B(n1600), .Z(n1602) );
  XNOR U1249 ( .A(n1224), .B(n1596), .Z(n1598) );
  XOR U1250 ( .A(n1604), .B(n1605), .Z(n1224) );
  AND U1251 ( .A(n1125), .B(n1606), .Z(n1605) );
  XOR U1252 ( .A(n1607), .B(n1604), .Z(n1606) );
  XOR U1253 ( .A(n1608), .B(n1609), .Z(n1596) );
  AND U1254 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U1255 ( .A(n1608), .B(n1239), .Z(n1611) );
  XOR U1256 ( .A(n1612), .B(n1613), .Z(n1239) );
  AND U1257 ( .A(n1127), .B(n1614), .Z(n1613) );
  XOR U1258 ( .A(n1615), .B(n1612), .Z(n1614) );
  XNOR U1259 ( .A(n1236), .B(n1608), .Z(n1610) );
  XOR U1260 ( .A(n1616), .B(n1617), .Z(n1236) );
  AND U1261 ( .A(n1125), .B(n1618), .Z(n1617) );
  XOR U1262 ( .A(n1619), .B(n1616), .Z(n1618) );
  XOR U1263 ( .A(n1620), .B(n1621), .Z(n1608) );
  AND U1264 ( .A(n1622), .B(n1623), .Z(n1621) );
  XOR U1265 ( .A(n1620), .B(n1251), .Z(n1623) );
  XOR U1266 ( .A(n1624), .B(n1625), .Z(n1251) );
  AND U1267 ( .A(n1127), .B(n1626), .Z(n1625) );
  XOR U1268 ( .A(n1627), .B(n1624), .Z(n1626) );
  XNOR U1269 ( .A(n1248), .B(n1620), .Z(n1622) );
  XOR U1270 ( .A(n1628), .B(n1629), .Z(n1248) );
  AND U1271 ( .A(n1125), .B(n1630), .Z(n1629) );
  XOR U1272 ( .A(n1631), .B(n1628), .Z(n1630) );
  XOR U1273 ( .A(n1632), .B(n1633), .Z(n1620) );
  AND U1274 ( .A(n1634), .B(n1635), .Z(n1633) );
  XOR U1275 ( .A(n1632), .B(n1263), .Z(n1635) );
  XOR U1276 ( .A(n1636), .B(n1637), .Z(n1263) );
  AND U1277 ( .A(n1127), .B(n1638), .Z(n1637) );
  XOR U1278 ( .A(n1639), .B(n1636), .Z(n1638) );
  XNOR U1279 ( .A(n1260), .B(n1632), .Z(n1634) );
  XOR U1280 ( .A(n1640), .B(n1641), .Z(n1260) );
  AND U1281 ( .A(n1125), .B(n1642), .Z(n1641) );
  XOR U1282 ( .A(n1643), .B(n1640), .Z(n1642) );
  XOR U1283 ( .A(n1644), .B(n1645), .Z(n1632) );
  AND U1284 ( .A(n1646), .B(n1647), .Z(n1645) );
  XOR U1285 ( .A(n1644), .B(n1275), .Z(n1647) );
  XOR U1286 ( .A(n1648), .B(n1649), .Z(n1275) );
  AND U1287 ( .A(n1127), .B(n1650), .Z(n1649) );
  XOR U1288 ( .A(n1651), .B(n1648), .Z(n1650) );
  XNOR U1289 ( .A(n1272), .B(n1644), .Z(n1646) );
  XOR U1290 ( .A(n1652), .B(n1653), .Z(n1272) );
  AND U1291 ( .A(n1125), .B(n1654), .Z(n1653) );
  XOR U1292 ( .A(n1655), .B(n1652), .Z(n1654) );
  XOR U1293 ( .A(n1656), .B(n1657), .Z(n1644) );
  AND U1294 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U1295 ( .A(n1656), .B(n1287), .Z(n1659) );
  XOR U1296 ( .A(n1660), .B(n1661), .Z(n1287) );
  AND U1297 ( .A(n1127), .B(n1662), .Z(n1661) );
  XOR U1298 ( .A(n1663), .B(n1660), .Z(n1662) );
  XNOR U1299 ( .A(n1284), .B(n1656), .Z(n1658) );
  XOR U1300 ( .A(n1664), .B(n1665), .Z(n1284) );
  AND U1301 ( .A(n1125), .B(n1666), .Z(n1665) );
  XOR U1302 ( .A(n1667), .B(n1664), .Z(n1666) );
  XOR U1303 ( .A(n1668), .B(n1669), .Z(n1656) );
  AND U1304 ( .A(n1670), .B(n1671), .Z(n1669) );
  XOR U1305 ( .A(n1668), .B(n1299), .Z(n1671) );
  XOR U1306 ( .A(n1672), .B(n1673), .Z(n1299) );
  AND U1307 ( .A(n1127), .B(n1674), .Z(n1673) );
  XOR U1308 ( .A(n1675), .B(n1672), .Z(n1674) );
  XNOR U1309 ( .A(n1296), .B(n1668), .Z(n1670) );
  XOR U1310 ( .A(n1676), .B(n1677), .Z(n1296) );
  AND U1311 ( .A(n1125), .B(n1678), .Z(n1677) );
  XOR U1312 ( .A(n1679), .B(n1676), .Z(n1678) );
  XOR U1313 ( .A(n1680), .B(n1681), .Z(n1668) );
  AND U1314 ( .A(n1682), .B(n1683), .Z(n1681) );
  XOR U1315 ( .A(n1680), .B(n1311), .Z(n1683) );
  XOR U1316 ( .A(n1684), .B(n1685), .Z(n1311) );
  AND U1317 ( .A(n1127), .B(n1686), .Z(n1685) );
  XOR U1318 ( .A(n1687), .B(n1684), .Z(n1686) );
  XNOR U1319 ( .A(n1308), .B(n1680), .Z(n1682) );
  XOR U1320 ( .A(n1688), .B(n1689), .Z(n1308) );
  AND U1321 ( .A(n1125), .B(n1690), .Z(n1689) );
  XOR U1322 ( .A(n1691), .B(n1688), .Z(n1690) );
  XOR U1323 ( .A(n1692), .B(n1693), .Z(n1680) );
  AND U1324 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U1325 ( .A(n1692), .B(n1323), .Z(n1695) );
  XOR U1326 ( .A(n1696), .B(n1697), .Z(n1323) );
  AND U1327 ( .A(n1127), .B(n1698), .Z(n1697) );
  XOR U1328 ( .A(n1699), .B(n1696), .Z(n1698) );
  XNOR U1329 ( .A(n1320), .B(n1692), .Z(n1694) );
  XOR U1330 ( .A(n1700), .B(n1701), .Z(n1320) );
  AND U1331 ( .A(n1125), .B(n1702), .Z(n1701) );
  XOR U1332 ( .A(n1703), .B(n1700), .Z(n1702) );
  XOR U1333 ( .A(n1704), .B(n1705), .Z(n1692) );
  AND U1334 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U1335 ( .A(n1704), .B(n1335), .Z(n1707) );
  XOR U1336 ( .A(n1708), .B(n1709), .Z(n1335) );
  AND U1337 ( .A(n1127), .B(n1710), .Z(n1709) );
  XOR U1338 ( .A(n1711), .B(n1708), .Z(n1710) );
  XNOR U1339 ( .A(n1332), .B(n1704), .Z(n1706) );
  XOR U1340 ( .A(n1712), .B(n1713), .Z(n1332) );
  AND U1341 ( .A(n1125), .B(n1714), .Z(n1713) );
  XOR U1342 ( .A(n1715), .B(n1712), .Z(n1714) );
  XOR U1343 ( .A(n1716), .B(n1717), .Z(n1704) );
  AND U1344 ( .A(n1718), .B(n1719), .Z(n1717) );
  XOR U1345 ( .A(n1716), .B(n1347), .Z(n1719) );
  XOR U1346 ( .A(n1720), .B(n1721), .Z(n1347) );
  AND U1347 ( .A(n1127), .B(n1722), .Z(n1721) );
  XOR U1348 ( .A(n1723), .B(n1720), .Z(n1722) );
  XNOR U1349 ( .A(n1344), .B(n1716), .Z(n1718) );
  XOR U1350 ( .A(n1724), .B(n1725), .Z(n1344) );
  AND U1351 ( .A(n1125), .B(n1726), .Z(n1725) );
  XOR U1352 ( .A(n1727), .B(n1724), .Z(n1726) );
  XOR U1353 ( .A(n1728), .B(n1729), .Z(n1716) );
  AND U1354 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U1355 ( .A(n1728), .B(n1359), .Z(n1731) );
  XOR U1356 ( .A(n1732), .B(n1733), .Z(n1359) );
  AND U1357 ( .A(n1127), .B(n1734), .Z(n1733) );
  XOR U1358 ( .A(n1735), .B(n1732), .Z(n1734) );
  XNOR U1359 ( .A(n1356), .B(n1728), .Z(n1730) );
  XOR U1360 ( .A(n1736), .B(n1737), .Z(n1356) );
  AND U1361 ( .A(n1125), .B(n1738), .Z(n1737) );
  XOR U1362 ( .A(n1739), .B(n1736), .Z(n1738) );
  XOR U1363 ( .A(n1740), .B(n1741), .Z(n1728) );
  AND U1364 ( .A(n1742), .B(n1743), .Z(n1741) );
  XOR U1365 ( .A(n1740), .B(n1371), .Z(n1743) );
  XOR U1366 ( .A(n1744), .B(n1745), .Z(n1371) );
  AND U1367 ( .A(n1127), .B(n1746), .Z(n1745) );
  XOR U1368 ( .A(n1747), .B(n1744), .Z(n1746) );
  XNOR U1369 ( .A(n1368), .B(n1740), .Z(n1742) );
  XOR U1370 ( .A(n1748), .B(n1749), .Z(n1368) );
  AND U1371 ( .A(n1125), .B(n1750), .Z(n1749) );
  XOR U1372 ( .A(n1751), .B(n1748), .Z(n1750) );
  XOR U1373 ( .A(n1752), .B(n1753), .Z(n1740) );
  AND U1374 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U1375 ( .A(n1752), .B(n1383), .Z(n1755) );
  XOR U1376 ( .A(n1756), .B(n1757), .Z(n1383) );
  AND U1377 ( .A(n1127), .B(n1758), .Z(n1757) );
  XOR U1378 ( .A(n1759), .B(n1756), .Z(n1758) );
  XNOR U1379 ( .A(n1380), .B(n1752), .Z(n1754) );
  XOR U1380 ( .A(n1760), .B(n1761), .Z(n1380) );
  AND U1381 ( .A(n1125), .B(n1762), .Z(n1761) );
  XOR U1382 ( .A(n1763), .B(n1760), .Z(n1762) );
  XOR U1383 ( .A(n1764), .B(n1765), .Z(n1752) );
  AND U1384 ( .A(n1766), .B(n1767), .Z(n1765) );
  XOR U1385 ( .A(n1764), .B(n1395), .Z(n1767) );
  XOR U1386 ( .A(n1768), .B(n1769), .Z(n1395) );
  AND U1387 ( .A(n1127), .B(n1770), .Z(n1769) );
  XOR U1388 ( .A(n1771), .B(n1768), .Z(n1770) );
  XNOR U1389 ( .A(n1392), .B(n1764), .Z(n1766) );
  XOR U1390 ( .A(n1772), .B(n1773), .Z(n1392) );
  AND U1391 ( .A(n1125), .B(n1774), .Z(n1773) );
  XOR U1392 ( .A(n1775), .B(n1772), .Z(n1774) );
  XOR U1393 ( .A(n1776), .B(n1777), .Z(n1764) );
  AND U1394 ( .A(n1778), .B(n1779), .Z(n1777) );
  XOR U1395 ( .A(n1776), .B(n1407), .Z(n1779) );
  XOR U1396 ( .A(n1780), .B(n1781), .Z(n1407) );
  AND U1397 ( .A(n1127), .B(n1782), .Z(n1781) );
  XOR U1398 ( .A(n1783), .B(n1780), .Z(n1782) );
  XNOR U1399 ( .A(n1404), .B(n1776), .Z(n1778) );
  XOR U1400 ( .A(n1784), .B(n1785), .Z(n1404) );
  AND U1401 ( .A(n1125), .B(n1786), .Z(n1785) );
  XOR U1402 ( .A(n1787), .B(n1784), .Z(n1786) );
  XOR U1403 ( .A(n1788), .B(n1789), .Z(n1776) );
  AND U1404 ( .A(n1790), .B(n1791), .Z(n1789) );
  XOR U1405 ( .A(n1788), .B(n1419), .Z(n1791) );
  XOR U1406 ( .A(n1792), .B(n1793), .Z(n1419) );
  AND U1407 ( .A(n1127), .B(n1794), .Z(n1793) );
  XOR U1408 ( .A(n1795), .B(n1792), .Z(n1794) );
  XNOR U1409 ( .A(n1416), .B(n1788), .Z(n1790) );
  XOR U1410 ( .A(n1796), .B(n1797), .Z(n1416) );
  AND U1411 ( .A(n1125), .B(n1798), .Z(n1797) );
  XOR U1412 ( .A(n1799), .B(n1796), .Z(n1798) );
  XOR U1413 ( .A(n1800), .B(n1801), .Z(n1788) );
  AND U1414 ( .A(n1802), .B(n1803), .Z(n1801) );
  XOR U1415 ( .A(n1800), .B(n1431), .Z(n1803) );
  XOR U1416 ( .A(n1804), .B(n1805), .Z(n1431) );
  AND U1417 ( .A(n1127), .B(n1806), .Z(n1805) );
  XOR U1418 ( .A(n1807), .B(n1804), .Z(n1806) );
  XNOR U1419 ( .A(n1428), .B(n1800), .Z(n1802) );
  XOR U1420 ( .A(n1808), .B(n1809), .Z(n1428) );
  AND U1421 ( .A(n1125), .B(n1810), .Z(n1809) );
  XOR U1422 ( .A(n1811), .B(n1808), .Z(n1810) );
  XOR U1423 ( .A(n1812), .B(n1813), .Z(n1800) );
  AND U1424 ( .A(n1814), .B(n1815), .Z(n1813) );
  XOR U1425 ( .A(n1812), .B(n1443), .Z(n1815) );
  XOR U1426 ( .A(n1816), .B(n1817), .Z(n1443) );
  AND U1427 ( .A(n1127), .B(n1818), .Z(n1817) );
  XOR U1428 ( .A(n1819), .B(n1816), .Z(n1818) );
  XNOR U1429 ( .A(n1440), .B(n1812), .Z(n1814) );
  XOR U1430 ( .A(n1820), .B(n1821), .Z(n1440) );
  AND U1431 ( .A(n1125), .B(n1822), .Z(n1821) );
  XOR U1432 ( .A(n1823), .B(n1820), .Z(n1822) );
  XOR U1433 ( .A(n1824), .B(n1825), .Z(n1812) );
  AND U1434 ( .A(n1826), .B(n1827), .Z(n1825) );
  XOR U1435 ( .A(n1824), .B(n1455), .Z(n1827) );
  XOR U1436 ( .A(n1828), .B(n1829), .Z(n1455) );
  AND U1437 ( .A(n1127), .B(n1830), .Z(n1829) );
  XOR U1438 ( .A(n1831), .B(n1828), .Z(n1830) );
  XNOR U1439 ( .A(n1452), .B(n1824), .Z(n1826) );
  XOR U1440 ( .A(n1832), .B(n1833), .Z(n1452) );
  AND U1441 ( .A(n1125), .B(n1834), .Z(n1833) );
  XOR U1442 ( .A(n1835), .B(n1832), .Z(n1834) );
  XOR U1443 ( .A(n1836), .B(n1837), .Z(n1824) );
  AND U1444 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U1445 ( .A(n1836), .B(n1467), .Z(n1839) );
  XOR U1446 ( .A(n1840), .B(n1841), .Z(n1467) );
  AND U1447 ( .A(n1127), .B(n1842), .Z(n1841) );
  XOR U1448 ( .A(n1843), .B(n1840), .Z(n1842) );
  XNOR U1449 ( .A(n1464), .B(n1836), .Z(n1838) );
  XOR U1450 ( .A(n1844), .B(n1845), .Z(n1464) );
  AND U1451 ( .A(n1125), .B(n1846), .Z(n1845) );
  XOR U1452 ( .A(n1847), .B(n1844), .Z(n1846) );
  XOR U1453 ( .A(n1848), .B(n1849), .Z(n1836) );
  AND U1454 ( .A(n1850), .B(n1851), .Z(n1849) );
  XOR U1455 ( .A(n1848), .B(n1479), .Z(n1851) );
  XOR U1456 ( .A(n1852), .B(n1853), .Z(n1479) );
  AND U1457 ( .A(n1127), .B(n1854), .Z(n1853) );
  XOR U1458 ( .A(n1855), .B(n1852), .Z(n1854) );
  XNOR U1459 ( .A(n1476), .B(n1848), .Z(n1850) );
  XOR U1460 ( .A(n1856), .B(n1857), .Z(n1476) );
  AND U1461 ( .A(n1125), .B(n1858), .Z(n1857) );
  XOR U1462 ( .A(n1859), .B(n1856), .Z(n1858) );
  XOR U1463 ( .A(n1860), .B(n1861), .Z(n1848) );
  AND U1464 ( .A(n1862), .B(n1863), .Z(n1861) );
  XOR U1465 ( .A(n1860), .B(n1491), .Z(n1863) );
  XOR U1466 ( .A(n1864), .B(n1865), .Z(n1491) );
  AND U1467 ( .A(n1127), .B(n1866), .Z(n1865) );
  XOR U1468 ( .A(n1867), .B(n1864), .Z(n1866) );
  XNOR U1469 ( .A(n1488), .B(n1860), .Z(n1862) );
  XOR U1470 ( .A(n1868), .B(n1869), .Z(n1488) );
  AND U1471 ( .A(n1125), .B(n1870), .Z(n1869) );
  XOR U1472 ( .A(n1871), .B(n1868), .Z(n1870) );
  XOR U1473 ( .A(n1872), .B(n1873), .Z(n1860) );
  AND U1474 ( .A(n1874), .B(n1875), .Z(n1873) );
  XOR U1475 ( .A(n1872), .B(n1503), .Z(n1875) );
  XOR U1476 ( .A(n1876), .B(n1877), .Z(n1503) );
  AND U1477 ( .A(n1127), .B(n1878), .Z(n1877) );
  XOR U1478 ( .A(n1879), .B(n1876), .Z(n1878) );
  XNOR U1479 ( .A(n1500), .B(n1872), .Z(n1874) );
  XOR U1480 ( .A(n1880), .B(n1881), .Z(n1500) );
  AND U1481 ( .A(n1125), .B(n1882), .Z(n1881) );
  XOR U1482 ( .A(n1883), .B(n1880), .Z(n1882) );
  XOR U1483 ( .A(n1884), .B(n1885), .Z(n1872) );
  AND U1484 ( .A(n1886), .B(n1887), .Z(n1885) );
  XNOR U1485 ( .A(n1888), .B(n1515), .Z(n1887) );
  XOR U1486 ( .A(n1889), .B(n1890), .Z(n1515) );
  AND U1487 ( .A(n1127), .B(n1891), .Z(n1890) );
  XOR U1488 ( .A(n1889), .B(n1892), .Z(n1891) );
  XNOR U1489 ( .A(n1512), .B(n1884), .Z(n1886) );
  XOR U1490 ( .A(n1893), .B(n1894), .Z(n1512) );
  AND U1491 ( .A(n1125), .B(n1895), .Z(n1894) );
  XOR U1492 ( .A(n1893), .B(n1896), .Z(n1895) );
  IV U1493 ( .A(n1888), .Z(n1884) );
  AND U1494 ( .A(n1520), .B(n1523), .Z(n1888) );
  XNOR U1495 ( .A(n1897), .B(n1898), .Z(n1523) );
  AND U1496 ( .A(n1127), .B(n1899), .Z(n1898) );
  XNOR U1497 ( .A(n1900), .B(n1897), .Z(n1899) );
  XOR U1498 ( .A(n1901), .B(n1902), .Z(n1127) );
  AND U1499 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U1500 ( .A(n1901), .B(n1531), .Z(n1904) );
  XOR U1501 ( .A(n1905), .B(n1906), .Z(n1531) );
  AND U1502 ( .A(n1087), .B(n1907), .Z(n1906) );
  XOR U1503 ( .A(n1908), .B(n1905), .Z(n1907) );
  XNOR U1504 ( .A(n1528), .B(n1901), .Z(n1903) );
  XOR U1505 ( .A(n1909), .B(n1910), .Z(n1528) );
  AND U1506 ( .A(n1085), .B(n1911), .Z(n1910) );
  XOR U1507 ( .A(n1912), .B(n1909), .Z(n1911) );
  XOR U1508 ( .A(n1913), .B(n1914), .Z(n1901) );
  AND U1509 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR U1510 ( .A(n1913), .B(n1543), .Z(n1916) );
  XOR U1511 ( .A(n1917), .B(n1918), .Z(n1543) );
  AND U1512 ( .A(n1087), .B(n1919), .Z(n1918) );
  XOR U1513 ( .A(n1920), .B(n1917), .Z(n1919) );
  XNOR U1514 ( .A(n1540), .B(n1913), .Z(n1915) );
  XOR U1515 ( .A(n1921), .B(n1922), .Z(n1540) );
  AND U1516 ( .A(n1085), .B(n1923), .Z(n1922) );
  XOR U1517 ( .A(n1924), .B(n1921), .Z(n1923) );
  XOR U1518 ( .A(n1925), .B(n1926), .Z(n1913) );
  AND U1519 ( .A(n1927), .B(n1928), .Z(n1926) );
  XOR U1520 ( .A(n1925), .B(n1555), .Z(n1928) );
  XOR U1521 ( .A(n1929), .B(n1930), .Z(n1555) );
  AND U1522 ( .A(n1087), .B(n1931), .Z(n1930) );
  XOR U1523 ( .A(n1932), .B(n1929), .Z(n1931) );
  XNOR U1524 ( .A(n1552), .B(n1925), .Z(n1927) );
  XOR U1525 ( .A(n1933), .B(n1934), .Z(n1552) );
  AND U1526 ( .A(n1085), .B(n1935), .Z(n1934) );
  XOR U1527 ( .A(n1936), .B(n1933), .Z(n1935) );
  XOR U1528 ( .A(n1937), .B(n1938), .Z(n1925) );
  AND U1529 ( .A(n1939), .B(n1940), .Z(n1938) );
  XOR U1530 ( .A(n1937), .B(n1567), .Z(n1940) );
  XOR U1531 ( .A(n1941), .B(n1942), .Z(n1567) );
  AND U1532 ( .A(n1087), .B(n1943), .Z(n1942) );
  XOR U1533 ( .A(n1944), .B(n1941), .Z(n1943) );
  XNOR U1534 ( .A(n1564), .B(n1937), .Z(n1939) );
  XOR U1535 ( .A(n1945), .B(n1946), .Z(n1564) );
  AND U1536 ( .A(n1085), .B(n1947), .Z(n1946) );
  XOR U1537 ( .A(n1948), .B(n1945), .Z(n1947) );
  XOR U1538 ( .A(n1949), .B(n1950), .Z(n1937) );
  AND U1539 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U1540 ( .A(n1949), .B(n1579), .Z(n1952) );
  XOR U1541 ( .A(n1953), .B(n1954), .Z(n1579) );
  AND U1542 ( .A(n1087), .B(n1955), .Z(n1954) );
  XOR U1543 ( .A(n1956), .B(n1953), .Z(n1955) );
  XNOR U1544 ( .A(n1576), .B(n1949), .Z(n1951) );
  XOR U1545 ( .A(n1957), .B(n1958), .Z(n1576) );
  AND U1546 ( .A(n1085), .B(n1959), .Z(n1958) );
  XOR U1547 ( .A(n1960), .B(n1957), .Z(n1959) );
  XOR U1548 ( .A(n1961), .B(n1962), .Z(n1949) );
  AND U1549 ( .A(n1963), .B(n1964), .Z(n1962) );
  XOR U1550 ( .A(n1961), .B(n1591), .Z(n1964) );
  XOR U1551 ( .A(n1965), .B(n1966), .Z(n1591) );
  AND U1552 ( .A(n1087), .B(n1967), .Z(n1966) );
  XOR U1553 ( .A(n1968), .B(n1965), .Z(n1967) );
  XNOR U1554 ( .A(n1588), .B(n1961), .Z(n1963) );
  XOR U1555 ( .A(n1969), .B(n1970), .Z(n1588) );
  AND U1556 ( .A(n1085), .B(n1971), .Z(n1970) );
  XOR U1557 ( .A(n1972), .B(n1969), .Z(n1971) );
  XOR U1558 ( .A(n1973), .B(n1974), .Z(n1961) );
  AND U1559 ( .A(n1975), .B(n1976), .Z(n1974) );
  XOR U1560 ( .A(n1973), .B(n1603), .Z(n1976) );
  XOR U1561 ( .A(n1977), .B(n1978), .Z(n1603) );
  AND U1562 ( .A(n1087), .B(n1979), .Z(n1978) );
  XOR U1563 ( .A(n1980), .B(n1977), .Z(n1979) );
  XNOR U1564 ( .A(n1600), .B(n1973), .Z(n1975) );
  XOR U1565 ( .A(n1981), .B(n1982), .Z(n1600) );
  AND U1566 ( .A(n1085), .B(n1983), .Z(n1982) );
  XOR U1567 ( .A(n1984), .B(n1981), .Z(n1983) );
  XOR U1568 ( .A(n1985), .B(n1986), .Z(n1973) );
  AND U1569 ( .A(n1987), .B(n1988), .Z(n1986) );
  XOR U1570 ( .A(n1985), .B(n1615), .Z(n1988) );
  XOR U1571 ( .A(n1989), .B(n1990), .Z(n1615) );
  AND U1572 ( .A(n1087), .B(n1991), .Z(n1990) );
  XOR U1573 ( .A(n1992), .B(n1989), .Z(n1991) );
  XNOR U1574 ( .A(n1612), .B(n1985), .Z(n1987) );
  XOR U1575 ( .A(n1993), .B(n1994), .Z(n1612) );
  AND U1576 ( .A(n1085), .B(n1995), .Z(n1994) );
  XOR U1577 ( .A(n1996), .B(n1993), .Z(n1995) );
  XOR U1578 ( .A(n1997), .B(n1998), .Z(n1985) );
  AND U1579 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR U1580 ( .A(n1997), .B(n1627), .Z(n2000) );
  XOR U1581 ( .A(n2001), .B(n2002), .Z(n1627) );
  AND U1582 ( .A(n1087), .B(n2003), .Z(n2002) );
  XOR U1583 ( .A(n2004), .B(n2001), .Z(n2003) );
  XNOR U1584 ( .A(n1624), .B(n1997), .Z(n1999) );
  XOR U1585 ( .A(n2005), .B(n2006), .Z(n1624) );
  AND U1586 ( .A(n1085), .B(n2007), .Z(n2006) );
  XOR U1587 ( .A(n2008), .B(n2005), .Z(n2007) );
  XOR U1588 ( .A(n2009), .B(n2010), .Z(n1997) );
  AND U1589 ( .A(n2011), .B(n2012), .Z(n2010) );
  XOR U1590 ( .A(n2009), .B(n1639), .Z(n2012) );
  XOR U1591 ( .A(n2013), .B(n2014), .Z(n1639) );
  AND U1592 ( .A(n1087), .B(n2015), .Z(n2014) );
  XOR U1593 ( .A(n2016), .B(n2013), .Z(n2015) );
  XNOR U1594 ( .A(n1636), .B(n2009), .Z(n2011) );
  XOR U1595 ( .A(n2017), .B(n2018), .Z(n1636) );
  AND U1596 ( .A(n1085), .B(n2019), .Z(n2018) );
  XOR U1597 ( .A(n2020), .B(n2017), .Z(n2019) );
  XOR U1598 ( .A(n2021), .B(n2022), .Z(n2009) );
  AND U1599 ( .A(n2023), .B(n2024), .Z(n2022) );
  XOR U1600 ( .A(n2021), .B(n1651), .Z(n2024) );
  XOR U1601 ( .A(n2025), .B(n2026), .Z(n1651) );
  AND U1602 ( .A(n1087), .B(n2027), .Z(n2026) );
  XOR U1603 ( .A(n2028), .B(n2025), .Z(n2027) );
  XNOR U1604 ( .A(n1648), .B(n2021), .Z(n2023) );
  XOR U1605 ( .A(n2029), .B(n2030), .Z(n1648) );
  AND U1606 ( .A(n1085), .B(n2031), .Z(n2030) );
  XOR U1607 ( .A(n2032), .B(n2029), .Z(n2031) );
  XOR U1608 ( .A(n2033), .B(n2034), .Z(n2021) );
  AND U1609 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U1610 ( .A(n2033), .B(n1663), .Z(n2036) );
  XOR U1611 ( .A(n2037), .B(n2038), .Z(n1663) );
  AND U1612 ( .A(n1087), .B(n2039), .Z(n2038) );
  XOR U1613 ( .A(n2040), .B(n2037), .Z(n2039) );
  XNOR U1614 ( .A(n1660), .B(n2033), .Z(n2035) );
  XOR U1615 ( .A(n2041), .B(n2042), .Z(n1660) );
  AND U1616 ( .A(n1085), .B(n2043), .Z(n2042) );
  XOR U1617 ( .A(n2044), .B(n2041), .Z(n2043) );
  XOR U1618 ( .A(n2045), .B(n2046), .Z(n2033) );
  AND U1619 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U1620 ( .A(n2045), .B(n1675), .Z(n2048) );
  XOR U1621 ( .A(n2049), .B(n2050), .Z(n1675) );
  AND U1622 ( .A(n1087), .B(n2051), .Z(n2050) );
  XOR U1623 ( .A(n2052), .B(n2049), .Z(n2051) );
  XNOR U1624 ( .A(n1672), .B(n2045), .Z(n2047) );
  XOR U1625 ( .A(n2053), .B(n2054), .Z(n1672) );
  AND U1626 ( .A(n1085), .B(n2055), .Z(n2054) );
  XOR U1627 ( .A(n2056), .B(n2053), .Z(n2055) );
  XOR U1628 ( .A(n2057), .B(n2058), .Z(n2045) );
  AND U1629 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U1630 ( .A(n2057), .B(n1687), .Z(n2060) );
  XOR U1631 ( .A(n2061), .B(n2062), .Z(n1687) );
  AND U1632 ( .A(n1087), .B(n2063), .Z(n2062) );
  XOR U1633 ( .A(n2064), .B(n2061), .Z(n2063) );
  XNOR U1634 ( .A(n1684), .B(n2057), .Z(n2059) );
  XOR U1635 ( .A(n2065), .B(n2066), .Z(n1684) );
  AND U1636 ( .A(n1085), .B(n2067), .Z(n2066) );
  XOR U1637 ( .A(n2068), .B(n2065), .Z(n2067) );
  XOR U1638 ( .A(n2069), .B(n2070), .Z(n2057) );
  AND U1639 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U1640 ( .A(n2069), .B(n1699), .Z(n2072) );
  XOR U1641 ( .A(n2073), .B(n2074), .Z(n1699) );
  AND U1642 ( .A(n1087), .B(n2075), .Z(n2074) );
  XOR U1643 ( .A(n2076), .B(n2073), .Z(n2075) );
  XNOR U1644 ( .A(n1696), .B(n2069), .Z(n2071) );
  XOR U1645 ( .A(n2077), .B(n2078), .Z(n1696) );
  AND U1646 ( .A(n1085), .B(n2079), .Z(n2078) );
  XOR U1647 ( .A(n2080), .B(n2077), .Z(n2079) );
  XOR U1648 ( .A(n2081), .B(n2082), .Z(n2069) );
  AND U1649 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U1650 ( .A(n2081), .B(n1711), .Z(n2084) );
  XOR U1651 ( .A(n2085), .B(n2086), .Z(n1711) );
  AND U1652 ( .A(n1087), .B(n2087), .Z(n2086) );
  XOR U1653 ( .A(n2088), .B(n2085), .Z(n2087) );
  XNOR U1654 ( .A(n1708), .B(n2081), .Z(n2083) );
  XOR U1655 ( .A(n2089), .B(n2090), .Z(n1708) );
  AND U1656 ( .A(n1085), .B(n2091), .Z(n2090) );
  XOR U1657 ( .A(n2092), .B(n2089), .Z(n2091) );
  XOR U1658 ( .A(n2093), .B(n2094), .Z(n2081) );
  AND U1659 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U1660 ( .A(n2093), .B(n1723), .Z(n2096) );
  XOR U1661 ( .A(n2097), .B(n2098), .Z(n1723) );
  AND U1662 ( .A(n1087), .B(n2099), .Z(n2098) );
  XOR U1663 ( .A(n2100), .B(n2097), .Z(n2099) );
  XNOR U1664 ( .A(n1720), .B(n2093), .Z(n2095) );
  XOR U1665 ( .A(n2101), .B(n2102), .Z(n1720) );
  AND U1666 ( .A(n1085), .B(n2103), .Z(n2102) );
  XOR U1667 ( .A(n2104), .B(n2101), .Z(n2103) );
  XOR U1668 ( .A(n2105), .B(n2106), .Z(n2093) );
  AND U1669 ( .A(n2107), .B(n2108), .Z(n2106) );
  XOR U1670 ( .A(n2105), .B(n1735), .Z(n2108) );
  XOR U1671 ( .A(n2109), .B(n2110), .Z(n1735) );
  AND U1672 ( .A(n1087), .B(n2111), .Z(n2110) );
  XOR U1673 ( .A(n2112), .B(n2109), .Z(n2111) );
  XNOR U1674 ( .A(n1732), .B(n2105), .Z(n2107) );
  XOR U1675 ( .A(n2113), .B(n2114), .Z(n1732) );
  AND U1676 ( .A(n1085), .B(n2115), .Z(n2114) );
  XOR U1677 ( .A(n2116), .B(n2113), .Z(n2115) );
  XOR U1678 ( .A(n2117), .B(n2118), .Z(n2105) );
  AND U1679 ( .A(n2119), .B(n2120), .Z(n2118) );
  XOR U1680 ( .A(n2117), .B(n1747), .Z(n2120) );
  XOR U1681 ( .A(n2121), .B(n2122), .Z(n1747) );
  AND U1682 ( .A(n1087), .B(n2123), .Z(n2122) );
  XOR U1683 ( .A(n2124), .B(n2121), .Z(n2123) );
  XNOR U1684 ( .A(n1744), .B(n2117), .Z(n2119) );
  XOR U1685 ( .A(n2125), .B(n2126), .Z(n1744) );
  AND U1686 ( .A(n1085), .B(n2127), .Z(n2126) );
  XOR U1687 ( .A(n2128), .B(n2125), .Z(n2127) );
  XOR U1688 ( .A(n2129), .B(n2130), .Z(n2117) );
  AND U1689 ( .A(n2131), .B(n2132), .Z(n2130) );
  XOR U1690 ( .A(n2129), .B(n1759), .Z(n2132) );
  XOR U1691 ( .A(n2133), .B(n2134), .Z(n1759) );
  AND U1692 ( .A(n1087), .B(n2135), .Z(n2134) );
  XOR U1693 ( .A(n2136), .B(n2133), .Z(n2135) );
  XNOR U1694 ( .A(n1756), .B(n2129), .Z(n2131) );
  XOR U1695 ( .A(n2137), .B(n2138), .Z(n1756) );
  AND U1696 ( .A(n1085), .B(n2139), .Z(n2138) );
  XOR U1697 ( .A(n2140), .B(n2137), .Z(n2139) );
  XOR U1698 ( .A(n2141), .B(n2142), .Z(n2129) );
  AND U1699 ( .A(n2143), .B(n2144), .Z(n2142) );
  XOR U1700 ( .A(n2141), .B(n1771), .Z(n2144) );
  XOR U1701 ( .A(n2145), .B(n2146), .Z(n1771) );
  AND U1702 ( .A(n1087), .B(n2147), .Z(n2146) );
  XOR U1703 ( .A(n2148), .B(n2145), .Z(n2147) );
  XNOR U1704 ( .A(n1768), .B(n2141), .Z(n2143) );
  XOR U1705 ( .A(n2149), .B(n2150), .Z(n1768) );
  AND U1706 ( .A(n1085), .B(n2151), .Z(n2150) );
  XOR U1707 ( .A(n2152), .B(n2149), .Z(n2151) );
  XOR U1708 ( .A(n2153), .B(n2154), .Z(n2141) );
  AND U1709 ( .A(n2155), .B(n2156), .Z(n2154) );
  XOR U1710 ( .A(n2153), .B(n1783), .Z(n2156) );
  XOR U1711 ( .A(n2157), .B(n2158), .Z(n1783) );
  AND U1712 ( .A(n1087), .B(n2159), .Z(n2158) );
  XOR U1713 ( .A(n2160), .B(n2157), .Z(n2159) );
  XNOR U1714 ( .A(n1780), .B(n2153), .Z(n2155) );
  XOR U1715 ( .A(n2161), .B(n2162), .Z(n1780) );
  AND U1716 ( .A(n1085), .B(n2163), .Z(n2162) );
  XOR U1717 ( .A(n2164), .B(n2161), .Z(n2163) );
  XOR U1718 ( .A(n2165), .B(n2166), .Z(n2153) );
  AND U1719 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U1720 ( .A(n2165), .B(n1795), .Z(n2168) );
  XOR U1721 ( .A(n2169), .B(n2170), .Z(n1795) );
  AND U1722 ( .A(n1087), .B(n2171), .Z(n2170) );
  XOR U1723 ( .A(n2172), .B(n2169), .Z(n2171) );
  XNOR U1724 ( .A(n1792), .B(n2165), .Z(n2167) );
  XOR U1725 ( .A(n2173), .B(n2174), .Z(n1792) );
  AND U1726 ( .A(n1085), .B(n2175), .Z(n2174) );
  XOR U1727 ( .A(n2176), .B(n2173), .Z(n2175) );
  XOR U1728 ( .A(n2177), .B(n2178), .Z(n2165) );
  AND U1729 ( .A(n2179), .B(n2180), .Z(n2178) );
  XOR U1730 ( .A(n2177), .B(n1807), .Z(n2180) );
  XOR U1731 ( .A(n2181), .B(n2182), .Z(n1807) );
  AND U1732 ( .A(n1087), .B(n2183), .Z(n2182) );
  XOR U1733 ( .A(n2184), .B(n2181), .Z(n2183) );
  XNOR U1734 ( .A(n1804), .B(n2177), .Z(n2179) );
  XOR U1735 ( .A(n2185), .B(n2186), .Z(n1804) );
  AND U1736 ( .A(n1085), .B(n2187), .Z(n2186) );
  XOR U1737 ( .A(n2188), .B(n2185), .Z(n2187) );
  XOR U1738 ( .A(n2189), .B(n2190), .Z(n2177) );
  AND U1739 ( .A(n2191), .B(n2192), .Z(n2190) );
  XOR U1740 ( .A(n2189), .B(n1819), .Z(n2192) );
  XOR U1741 ( .A(n2193), .B(n2194), .Z(n1819) );
  AND U1742 ( .A(n1087), .B(n2195), .Z(n2194) );
  XOR U1743 ( .A(n2196), .B(n2193), .Z(n2195) );
  XNOR U1744 ( .A(n1816), .B(n2189), .Z(n2191) );
  XOR U1745 ( .A(n2197), .B(n2198), .Z(n1816) );
  AND U1746 ( .A(n1085), .B(n2199), .Z(n2198) );
  XOR U1747 ( .A(n2200), .B(n2197), .Z(n2199) );
  XOR U1748 ( .A(n2201), .B(n2202), .Z(n2189) );
  AND U1749 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR U1750 ( .A(n2201), .B(n1831), .Z(n2204) );
  XOR U1751 ( .A(n2205), .B(n2206), .Z(n1831) );
  AND U1752 ( .A(n1087), .B(n2207), .Z(n2206) );
  XOR U1753 ( .A(n2208), .B(n2205), .Z(n2207) );
  XNOR U1754 ( .A(n1828), .B(n2201), .Z(n2203) );
  XOR U1755 ( .A(n2209), .B(n2210), .Z(n1828) );
  AND U1756 ( .A(n1085), .B(n2211), .Z(n2210) );
  XOR U1757 ( .A(n2212), .B(n2209), .Z(n2211) );
  XOR U1758 ( .A(n2213), .B(n2214), .Z(n2201) );
  AND U1759 ( .A(n2215), .B(n2216), .Z(n2214) );
  XOR U1760 ( .A(n2213), .B(n1843), .Z(n2216) );
  XOR U1761 ( .A(n2217), .B(n2218), .Z(n1843) );
  AND U1762 ( .A(n1087), .B(n2219), .Z(n2218) );
  XOR U1763 ( .A(n2220), .B(n2217), .Z(n2219) );
  XNOR U1764 ( .A(n1840), .B(n2213), .Z(n2215) );
  XOR U1765 ( .A(n2221), .B(n2222), .Z(n1840) );
  AND U1766 ( .A(n1085), .B(n2223), .Z(n2222) );
  XOR U1767 ( .A(n2224), .B(n2221), .Z(n2223) );
  XOR U1768 ( .A(n2225), .B(n2226), .Z(n2213) );
  AND U1769 ( .A(n2227), .B(n2228), .Z(n2226) );
  XOR U1770 ( .A(n2225), .B(n1855), .Z(n2228) );
  XOR U1771 ( .A(n2229), .B(n2230), .Z(n1855) );
  AND U1772 ( .A(n1087), .B(n2231), .Z(n2230) );
  XOR U1773 ( .A(n2232), .B(n2229), .Z(n2231) );
  XNOR U1774 ( .A(n1852), .B(n2225), .Z(n2227) );
  XOR U1775 ( .A(n2233), .B(n2234), .Z(n1852) );
  AND U1776 ( .A(n1085), .B(n2235), .Z(n2234) );
  XOR U1777 ( .A(n2236), .B(n2233), .Z(n2235) );
  XOR U1778 ( .A(n2237), .B(n2238), .Z(n2225) );
  AND U1779 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U1780 ( .A(n2237), .B(n1867), .Z(n2240) );
  XOR U1781 ( .A(n2241), .B(n2242), .Z(n1867) );
  AND U1782 ( .A(n1087), .B(n2243), .Z(n2242) );
  XOR U1783 ( .A(n2244), .B(n2241), .Z(n2243) );
  XNOR U1784 ( .A(n1864), .B(n2237), .Z(n2239) );
  XOR U1785 ( .A(n2245), .B(n2246), .Z(n1864) );
  AND U1786 ( .A(n1085), .B(n2247), .Z(n2246) );
  XOR U1787 ( .A(n2248), .B(n2245), .Z(n2247) );
  XOR U1788 ( .A(n2249), .B(n2250), .Z(n2237) );
  AND U1789 ( .A(n2251), .B(n2252), .Z(n2250) );
  XOR U1790 ( .A(n2249), .B(n1879), .Z(n2252) );
  XOR U1791 ( .A(n2253), .B(n2254), .Z(n1879) );
  AND U1792 ( .A(n1087), .B(n2255), .Z(n2254) );
  XOR U1793 ( .A(n2256), .B(n2253), .Z(n2255) );
  XNOR U1794 ( .A(n1876), .B(n2249), .Z(n2251) );
  XOR U1795 ( .A(n2257), .B(n2258), .Z(n1876) );
  AND U1796 ( .A(n1085), .B(n2259), .Z(n2258) );
  XOR U1797 ( .A(n2260), .B(n2257), .Z(n2259) );
  XOR U1798 ( .A(n2261), .B(n2262), .Z(n2249) );
  AND U1799 ( .A(n2263), .B(n2264), .Z(n2262) );
  XNOR U1800 ( .A(n2265), .B(n1892), .Z(n2264) );
  XOR U1801 ( .A(n2266), .B(n2267), .Z(n1892) );
  AND U1802 ( .A(n1087), .B(n2268), .Z(n2267) );
  XOR U1803 ( .A(n2266), .B(n2269), .Z(n2268) );
  XNOR U1804 ( .A(n1889), .B(n2261), .Z(n2263) );
  XOR U1805 ( .A(n2270), .B(n2271), .Z(n1889) );
  AND U1806 ( .A(n1085), .B(n2272), .Z(n2271) );
  XOR U1807 ( .A(n2270), .B(n2273), .Z(n2272) );
  IV U1808 ( .A(n2265), .Z(n2261) );
  AND U1809 ( .A(n1897), .B(n1900), .Z(n2265) );
  XNOR U1810 ( .A(n2274), .B(n2275), .Z(n1900) );
  AND U1811 ( .A(n1087), .B(n2276), .Z(n2275) );
  XNOR U1812 ( .A(n2277), .B(n2274), .Z(n2276) );
  XOR U1813 ( .A(n2278), .B(n2279), .Z(n1087) );
  AND U1814 ( .A(n2280), .B(n2281), .Z(n2279) );
  XOR U1815 ( .A(n2278), .B(n1908), .Z(n2281) );
  XOR U1816 ( .A(n2282), .B(n2283), .Z(n1908) );
  AND U1817 ( .A(n999), .B(n2284), .Z(n2283) );
  XOR U1818 ( .A(n2285), .B(n2282), .Z(n2284) );
  XNOR U1819 ( .A(n1905), .B(n2278), .Z(n2280) );
  XOR U1820 ( .A(n2286), .B(n2287), .Z(n1905) );
  AND U1821 ( .A(n997), .B(n2288), .Z(n2287) );
  XOR U1822 ( .A(n2289), .B(n2286), .Z(n2288) );
  XOR U1823 ( .A(n2290), .B(n2291), .Z(n2278) );
  AND U1824 ( .A(n2292), .B(n2293), .Z(n2291) );
  XOR U1825 ( .A(n2290), .B(n1920), .Z(n2293) );
  XOR U1826 ( .A(n2294), .B(n2295), .Z(n1920) );
  AND U1827 ( .A(n999), .B(n2296), .Z(n2295) );
  XOR U1828 ( .A(n2297), .B(n2294), .Z(n2296) );
  XNOR U1829 ( .A(n1917), .B(n2290), .Z(n2292) );
  XOR U1830 ( .A(n2298), .B(n2299), .Z(n1917) );
  AND U1831 ( .A(n997), .B(n2300), .Z(n2299) );
  XOR U1832 ( .A(n2301), .B(n2298), .Z(n2300) );
  XOR U1833 ( .A(n2302), .B(n2303), .Z(n2290) );
  AND U1834 ( .A(n2304), .B(n2305), .Z(n2303) );
  XOR U1835 ( .A(n2302), .B(n1932), .Z(n2305) );
  XOR U1836 ( .A(n2306), .B(n2307), .Z(n1932) );
  AND U1837 ( .A(n999), .B(n2308), .Z(n2307) );
  XOR U1838 ( .A(n2309), .B(n2306), .Z(n2308) );
  XNOR U1839 ( .A(n1929), .B(n2302), .Z(n2304) );
  XOR U1840 ( .A(n2310), .B(n2311), .Z(n1929) );
  AND U1841 ( .A(n997), .B(n2312), .Z(n2311) );
  XOR U1842 ( .A(n2313), .B(n2310), .Z(n2312) );
  XOR U1843 ( .A(n2314), .B(n2315), .Z(n2302) );
  AND U1844 ( .A(n2316), .B(n2317), .Z(n2315) );
  XOR U1845 ( .A(n2314), .B(n1944), .Z(n2317) );
  XOR U1846 ( .A(n2318), .B(n2319), .Z(n1944) );
  AND U1847 ( .A(n999), .B(n2320), .Z(n2319) );
  XOR U1848 ( .A(n2321), .B(n2318), .Z(n2320) );
  XNOR U1849 ( .A(n1941), .B(n2314), .Z(n2316) );
  XOR U1850 ( .A(n2322), .B(n2323), .Z(n1941) );
  AND U1851 ( .A(n997), .B(n2324), .Z(n2323) );
  XOR U1852 ( .A(n2325), .B(n2322), .Z(n2324) );
  XOR U1853 ( .A(n2326), .B(n2327), .Z(n2314) );
  AND U1854 ( .A(n2328), .B(n2329), .Z(n2327) );
  XOR U1855 ( .A(n2326), .B(n1956), .Z(n2329) );
  XOR U1856 ( .A(n2330), .B(n2331), .Z(n1956) );
  AND U1857 ( .A(n999), .B(n2332), .Z(n2331) );
  XOR U1858 ( .A(n2333), .B(n2330), .Z(n2332) );
  XNOR U1859 ( .A(n1953), .B(n2326), .Z(n2328) );
  XOR U1860 ( .A(n2334), .B(n2335), .Z(n1953) );
  AND U1861 ( .A(n997), .B(n2336), .Z(n2335) );
  XOR U1862 ( .A(n2337), .B(n2334), .Z(n2336) );
  XOR U1863 ( .A(n2338), .B(n2339), .Z(n2326) );
  AND U1864 ( .A(n2340), .B(n2341), .Z(n2339) );
  XOR U1865 ( .A(n2338), .B(n1968), .Z(n2341) );
  XOR U1866 ( .A(n2342), .B(n2343), .Z(n1968) );
  AND U1867 ( .A(n999), .B(n2344), .Z(n2343) );
  XOR U1868 ( .A(n2345), .B(n2342), .Z(n2344) );
  XNOR U1869 ( .A(n1965), .B(n2338), .Z(n2340) );
  XOR U1870 ( .A(n2346), .B(n2347), .Z(n1965) );
  AND U1871 ( .A(n997), .B(n2348), .Z(n2347) );
  XOR U1872 ( .A(n2349), .B(n2346), .Z(n2348) );
  XOR U1873 ( .A(n2350), .B(n2351), .Z(n2338) );
  AND U1874 ( .A(n2352), .B(n2353), .Z(n2351) );
  XOR U1875 ( .A(n2350), .B(n1980), .Z(n2353) );
  XOR U1876 ( .A(n2354), .B(n2355), .Z(n1980) );
  AND U1877 ( .A(n999), .B(n2356), .Z(n2355) );
  XOR U1878 ( .A(n2357), .B(n2354), .Z(n2356) );
  XNOR U1879 ( .A(n1977), .B(n2350), .Z(n2352) );
  XOR U1880 ( .A(n2358), .B(n2359), .Z(n1977) );
  AND U1881 ( .A(n997), .B(n2360), .Z(n2359) );
  XOR U1882 ( .A(n2361), .B(n2358), .Z(n2360) );
  XOR U1883 ( .A(n2362), .B(n2363), .Z(n2350) );
  AND U1884 ( .A(n2364), .B(n2365), .Z(n2363) );
  XOR U1885 ( .A(n2362), .B(n1992), .Z(n2365) );
  XOR U1886 ( .A(n2366), .B(n2367), .Z(n1992) );
  AND U1887 ( .A(n999), .B(n2368), .Z(n2367) );
  XOR U1888 ( .A(n2369), .B(n2366), .Z(n2368) );
  XNOR U1889 ( .A(n1989), .B(n2362), .Z(n2364) );
  XOR U1890 ( .A(n2370), .B(n2371), .Z(n1989) );
  AND U1891 ( .A(n997), .B(n2372), .Z(n2371) );
  XOR U1892 ( .A(n2373), .B(n2370), .Z(n2372) );
  XOR U1893 ( .A(n2374), .B(n2375), .Z(n2362) );
  AND U1894 ( .A(n2376), .B(n2377), .Z(n2375) );
  XOR U1895 ( .A(n2374), .B(n2004), .Z(n2377) );
  XOR U1896 ( .A(n2378), .B(n2379), .Z(n2004) );
  AND U1897 ( .A(n999), .B(n2380), .Z(n2379) );
  XOR U1898 ( .A(n2381), .B(n2378), .Z(n2380) );
  XNOR U1899 ( .A(n2001), .B(n2374), .Z(n2376) );
  XOR U1900 ( .A(n2382), .B(n2383), .Z(n2001) );
  AND U1901 ( .A(n997), .B(n2384), .Z(n2383) );
  XOR U1902 ( .A(n2385), .B(n2382), .Z(n2384) );
  XOR U1903 ( .A(n2386), .B(n2387), .Z(n2374) );
  AND U1904 ( .A(n2388), .B(n2389), .Z(n2387) );
  XOR U1905 ( .A(n2386), .B(n2016), .Z(n2389) );
  XOR U1906 ( .A(n2390), .B(n2391), .Z(n2016) );
  AND U1907 ( .A(n999), .B(n2392), .Z(n2391) );
  XOR U1908 ( .A(n2393), .B(n2390), .Z(n2392) );
  XNOR U1909 ( .A(n2013), .B(n2386), .Z(n2388) );
  XOR U1910 ( .A(n2394), .B(n2395), .Z(n2013) );
  AND U1911 ( .A(n997), .B(n2396), .Z(n2395) );
  XOR U1912 ( .A(n2397), .B(n2394), .Z(n2396) );
  XOR U1913 ( .A(n2398), .B(n2399), .Z(n2386) );
  AND U1914 ( .A(n2400), .B(n2401), .Z(n2399) );
  XOR U1915 ( .A(n2398), .B(n2028), .Z(n2401) );
  XOR U1916 ( .A(n2402), .B(n2403), .Z(n2028) );
  AND U1917 ( .A(n999), .B(n2404), .Z(n2403) );
  XOR U1918 ( .A(n2405), .B(n2402), .Z(n2404) );
  XNOR U1919 ( .A(n2025), .B(n2398), .Z(n2400) );
  XOR U1920 ( .A(n2406), .B(n2407), .Z(n2025) );
  AND U1921 ( .A(n997), .B(n2408), .Z(n2407) );
  XOR U1922 ( .A(n2409), .B(n2406), .Z(n2408) );
  XOR U1923 ( .A(n2410), .B(n2411), .Z(n2398) );
  AND U1924 ( .A(n2412), .B(n2413), .Z(n2411) );
  XOR U1925 ( .A(n2410), .B(n2040), .Z(n2413) );
  XOR U1926 ( .A(n2414), .B(n2415), .Z(n2040) );
  AND U1927 ( .A(n999), .B(n2416), .Z(n2415) );
  XOR U1928 ( .A(n2417), .B(n2414), .Z(n2416) );
  XNOR U1929 ( .A(n2037), .B(n2410), .Z(n2412) );
  XOR U1930 ( .A(n2418), .B(n2419), .Z(n2037) );
  AND U1931 ( .A(n997), .B(n2420), .Z(n2419) );
  XOR U1932 ( .A(n2421), .B(n2418), .Z(n2420) );
  XOR U1933 ( .A(n2422), .B(n2423), .Z(n2410) );
  AND U1934 ( .A(n2424), .B(n2425), .Z(n2423) );
  XOR U1935 ( .A(n2422), .B(n2052), .Z(n2425) );
  XOR U1936 ( .A(n2426), .B(n2427), .Z(n2052) );
  AND U1937 ( .A(n999), .B(n2428), .Z(n2427) );
  XOR U1938 ( .A(n2429), .B(n2426), .Z(n2428) );
  XNOR U1939 ( .A(n2049), .B(n2422), .Z(n2424) );
  XOR U1940 ( .A(n2430), .B(n2431), .Z(n2049) );
  AND U1941 ( .A(n997), .B(n2432), .Z(n2431) );
  XOR U1942 ( .A(n2433), .B(n2430), .Z(n2432) );
  XOR U1943 ( .A(n2434), .B(n2435), .Z(n2422) );
  AND U1944 ( .A(n2436), .B(n2437), .Z(n2435) );
  XOR U1945 ( .A(n2434), .B(n2064), .Z(n2437) );
  XOR U1946 ( .A(n2438), .B(n2439), .Z(n2064) );
  AND U1947 ( .A(n999), .B(n2440), .Z(n2439) );
  XOR U1948 ( .A(n2441), .B(n2438), .Z(n2440) );
  XNOR U1949 ( .A(n2061), .B(n2434), .Z(n2436) );
  XOR U1950 ( .A(n2442), .B(n2443), .Z(n2061) );
  AND U1951 ( .A(n997), .B(n2444), .Z(n2443) );
  XOR U1952 ( .A(n2445), .B(n2442), .Z(n2444) );
  XOR U1953 ( .A(n2446), .B(n2447), .Z(n2434) );
  AND U1954 ( .A(n2448), .B(n2449), .Z(n2447) );
  XOR U1955 ( .A(n2446), .B(n2076), .Z(n2449) );
  XOR U1956 ( .A(n2450), .B(n2451), .Z(n2076) );
  AND U1957 ( .A(n999), .B(n2452), .Z(n2451) );
  XOR U1958 ( .A(n2453), .B(n2450), .Z(n2452) );
  XNOR U1959 ( .A(n2073), .B(n2446), .Z(n2448) );
  XOR U1960 ( .A(n2454), .B(n2455), .Z(n2073) );
  AND U1961 ( .A(n997), .B(n2456), .Z(n2455) );
  XOR U1962 ( .A(n2457), .B(n2454), .Z(n2456) );
  XOR U1963 ( .A(n2458), .B(n2459), .Z(n2446) );
  AND U1964 ( .A(n2460), .B(n2461), .Z(n2459) );
  XOR U1965 ( .A(n2458), .B(n2088), .Z(n2461) );
  XOR U1966 ( .A(n2462), .B(n2463), .Z(n2088) );
  AND U1967 ( .A(n999), .B(n2464), .Z(n2463) );
  XOR U1968 ( .A(n2465), .B(n2462), .Z(n2464) );
  XNOR U1969 ( .A(n2085), .B(n2458), .Z(n2460) );
  XOR U1970 ( .A(n2466), .B(n2467), .Z(n2085) );
  AND U1971 ( .A(n997), .B(n2468), .Z(n2467) );
  XOR U1972 ( .A(n2469), .B(n2466), .Z(n2468) );
  XOR U1973 ( .A(n2470), .B(n2471), .Z(n2458) );
  AND U1974 ( .A(n2472), .B(n2473), .Z(n2471) );
  XOR U1975 ( .A(n2470), .B(n2100), .Z(n2473) );
  XOR U1976 ( .A(n2474), .B(n2475), .Z(n2100) );
  AND U1977 ( .A(n999), .B(n2476), .Z(n2475) );
  XOR U1978 ( .A(n2477), .B(n2474), .Z(n2476) );
  XNOR U1979 ( .A(n2097), .B(n2470), .Z(n2472) );
  XOR U1980 ( .A(n2478), .B(n2479), .Z(n2097) );
  AND U1981 ( .A(n997), .B(n2480), .Z(n2479) );
  XOR U1982 ( .A(n2481), .B(n2478), .Z(n2480) );
  XOR U1983 ( .A(n2482), .B(n2483), .Z(n2470) );
  AND U1984 ( .A(n2484), .B(n2485), .Z(n2483) );
  XOR U1985 ( .A(n2482), .B(n2112), .Z(n2485) );
  XOR U1986 ( .A(n2486), .B(n2487), .Z(n2112) );
  AND U1987 ( .A(n999), .B(n2488), .Z(n2487) );
  XOR U1988 ( .A(n2489), .B(n2486), .Z(n2488) );
  XNOR U1989 ( .A(n2109), .B(n2482), .Z(n2484) );
  XOR U1990 ( .A(n2490), .B(n2491), .Z(n2109) );
  AND U1991 ( .A(n997), .B(n2492), .Z(n2491) );
  XOR U1992 ( .A(n2493), .B(n2490), .Z(n2492) );
  XOR U1993 ( .A(n2494), .B(n2495), .Z(n2482) );
  AND U1994 ( .A(n2496), .B(n2497), .Z(n2495) );
  XOR U1995 ( .A(n2494), .B(n2124), .Z(n2497) );
  XOR U1996 ( .A(n2498), .B(n2499), .Z(n2124) );
  AND U1997 ( .A(n999), .B(n2500), .Z(n2499) );
  XOR U1998 ( .A(n2501), .B(n2498), .Z(n2500) );
  XNOR U1999 ( .A(n2121), .B(n2494), .Z(n2496) );
  XOR U2000 ( .A(n2502), .B(n2503), .Z(n2121) );
  AND U2001 ( .A(n997), .B(n2504), .Z(n2503) );
  XOR U2002 ( .A(n2505), .B(n2502), .Z(n2504) );
  XOR U2003 ( .A(n2506), .B(n2507), .Z(n2494) );
  AND U2004 ( .A(n2508), .B(n2509), .Z(n2507) );
  XOR U2005 ( .A(n2506), .B(n2136), .Z(n2509) );
  XOR U2006 ( .A(n2510), .B(n2511), .Z(n2136) );
  AND U2007 ( .A(n999), .B(n2512), .Z(n2511) );
  XOR U2008 ( .A(n2513), .B(n2510), .Z(n2512) );
  XNOR U2009 ( .A(n2133), .B(n2506), .Z(n2508) );
  XOR U2010 ( .A(n2514), .B(n2515), .Z(n2133) );
  AND U2011 ( .A(n997), .B(n2516), .Z(n2515) );
  XOR U2012 ( .A(n2517), .B(n2514), .Z(n2516) );
  XOR U2013 ( .A(n2518), .B(n2519), .Z(n2506) );
  AND U2014 ( .A(n2520), .B(n2521), .Z(n2519) );
  XOR U2015 ( .A(n2518), .B(n2148), .Z(n2521) );
  XOR U2016 ( .A(n2522), .B(n2523), .Z(n2148) );
  AND U2017 ( .A(n999), .B(n2524), .Z(n2523) );
  XOR U2018 ( .A(n2525), .B(n2522), .Z(n2524) );
  XNOR U2019 ( .A(n2145), .B(n2518), .Z(n2520) );
  XOR U2020 ( .A(n2526), .B(n2527), .Z(n2145) );
  AND U2021 ( .A(n997), .B(n2528), .Z(n2527) );
  XOR U2022 ( .A(n2529), .B(n2526), .Z(n2528) );
  XOR U2023 ( .A(n2530), .B(n2531), .Z(n2518) );
  AND U2024 ( .A(n2532), .B(n2533), .Z(n2531) );
  XOR U2025 ( .A(n2530), .B(n2160), .Z(n2533) );
  XOR U2026 ( .A(n2534), .B(n2535), .Z(n2160) );
  AND U2027 ( .A(n999), .B(n2536), .Z(n2535) );
  XOR U2028 ( .A(n2537), .B(n2534), .Z(n2536) );
  XNOR U2029 ( .A(n2157), .B(n2530), .Z(n2532) );
  XOR U2030 ( .A(n2538), .B(n2539), .Z(n2157) );
  AND U2031 ( .A(n997), .B(n2540), .Z(n2539) );
  XOR U2032 ( .A(n2541), .B(n2538), .Z(n2540) );
  XOR U2033 ( .A(n2542), .B(n2543), .Z(n2530) );
  AND U2034 ( .A(n2544), .B(n2545), .Z(n2543) );
  XOR U2035 ( .A(n2542), .B(n2172), .Z(n2545) );
  XOR U2036 ( .A(n2546), .B(n2547), .Z(n2172) );
  AND U2037 ( .A(n999), .B(n2548), .Z(n2547) );
  XOR U2038 ( .A(n2549), .B(n2546), .Z(n2548) );
  XNOR U2039 ( .A(n2169), .B(n2542), .Z(n2544) );
  XOR U2040 ( .A(n2550), .B(n2551), .Z(n2169) );
  AND U2041 ( .A(n997), .B(n2552), .Z(n2551) );
  XOR U2042 ( .A(n2553), .B(n2550), .Z(n2552) );
  XOR U2043 ( .A(n2554), .B(n2555), .Z(n2542) );
  AND U2044 ( .A(n2556), .B(n2557), .Z(n2555) );
  XOR U2045 ( .A(n2554), .B(n2184), .Z(n2557) );
  XOR U2046 ( .A(n2558), .B(n2559), .Z(n2184) );
  AND U2047 ( .A(n999), .B(n2560), .Z(n2559) );
  XOR U2048 ( .A(n2561), .B(n2558), .Z(n2560) );
  XNOR U2049 ( .A(n2181), .B(n2554), .Z(n2556) );
  XOR U2050 ( .A(n2562), .B(n2563), .Z(n2181) );
  AND U2051 ( .A(n997), .B(n2564), .Z(n2563) );
  XOR U2052 ( .A(n2565), .B(n2562), .Z(n2564) );
  XOR U2053 ( .A(n2566), .B(n2567), .Z(n2554) );
  AND U2054 ( .A(n2568), .B(n2569), .Z(n2567) );
  XOR U2055 ( .A(n2566), .B(n2196), .Z(n2569) );
  XOR U2056 ( .A(n2570), .B(n2571), .Z(n2196) );
  AND U2057 ( .A(n999), .B(n2572), .Z(n2571) );
  XOR U2058 ( .A(n2573), .B(n2570), .Z(n2572) );
  XNOR U2059 ( .A(n2193), .B(n2566), .Z(n2568) );
  XOR U2060 ( .A(n2574), .B(n2575), .Z(n2193) );
  AND U2061 ( .A(n997), .B(n2576), .Z(n2575) );
  XOR U2062 ( .A(n2577), .B(n2574), .Z(n2576) );
  XOR U2063 ( .A(n2578), .B(n2579), .Z(n2566) );
  AND U2064 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U2065 ( .A(n2578), .B(n2208), .Z(n2581) );
  XOR U2066 ( .A(n2582), .B(n2583), .Z(n2208) );
  AND U2067 ( .A(n999), .B(n2584), .Z(n2583) );
  XOR U2068 ( .A(n2585), .B(n2582), .Z(n2584) );
  XNOR U2069 ( .A(n2205), .B(n2578), .Z(n2580) );
  XOR U2070 ( .A(n2586), .B(n2587), .Z(n2205) );
  AND U2071 ( .A(n997), .B(n2588), .Z(n2587) );
  XOR U2072 ( .A(n2589), .B(n2586), .Z(n2588) );
  XOR U2073 ( .A(n2590), .B(n2591), .Z(n2578) );
  AND U2074 ( .A(n2592), .B(n2593), .Z(n2591) );
  XOR U2075 ( .A(n2590), .B(n2220), .Z(n2593) );
  XOR U2076 ( .A(n2594), .B(n2595), .Z(n2220) );
  AND U2077 ( .A(n999), .B(n2596), .Z(n2595) );
  XOR U2078 ( .A(n2597), .B(n2594), .Z(n2596) );
  XNOR U2079 ( .A(n2217), .B(n2590), .Z(n2592) );
  XOR U2080 ( .A(n2598), .B(n2599), .Z(n2217) );
  AND U2081 ( .A(n997), .B(n2600), .Z(n2599) );
  XOR U2082 ( .A(n2601), .B(n2598), .Z(n2600) );
  XOR U2083 ( .A(n2602), .B(n2603), .Z(n2590) );
  AND U2084 ( .A(n2604), .B(n2605), .Z(n2603) );
  XOR U2085 ( .A(n2602), .B(n2232), .Z(n2605) );
  XOR U2086 ( .A(n2606), .B(n2607), .Z(n2232) );
  AND U2087 ( .A(n999), .B(n2608), .Z(n2607) );
  XOR U2088 ( .A(n2609), .B(n2606), .Z(n2608) );
  XNOR U2089 ( .A(n2229), .B(n2602), .Z(n2604) );
  XOR U2090 ( .A(n2610), .B(n2611), .Z(n2229) );
  AND U2091 ( .A(n997), .B(n2612), .Z(n2611) );
  XOR U2092 ( .A(n2613), .B(n2610), .Z(n2612) );
  XOR U2093 ( .A(n2614), .B(n2615), .Z(n2602) );
  AND U2094 ( .A(n2616), .B(n2617), .Z(n2615) );
  XOR U2095 ( .A(n2614), .B(n2244), .Z(n2617) );
  XOR U2096 ( .A(n2618), .B(n2619), .Z(n2244) );
  AND U2097 ( .A(n999), .B(n2620), .Z(n2619) );
  XOR U2098 ( .A(n2621), .B(n2618), .Z(n2620) );
  XNOR U2099 ( .A(n2241), .B(n2614), .Z(n2616) );
  XOR U2100 ( .A(n2622), .B(n2623), .Z(n2241) );
  AND U2101 ( .A(n997), .B(n2624), .Z(n2623) );
  XOR U2102 ( .A(n2625), .B(n2622), .Z(n2624) );
  XOR U2103 ( .A(n2626), .B(n2627), .Z(n2614) );
  AND U2104 ( .A(n2628), .B(n2629), .Z(n2627) );
  XOR U2105 ( .A(n2626), .B(n2256), .Z(n2629) );
  XOR U2106 ( .A(n2630), .B(n2631), .Z(n2256) );
  AND U2107 ( .A(n999), .B(n2632), .Z(n2631) );
  XOR U2108 ( .A(n2633), .B(n2630), .Z(n2632) );
  XNOR U2109 ( .A(n2253), .B(n2626), .Z(n2628) );
  XOR U2110 ( .A(n2634), .B(n2635), .Z(n2253) );
  AND U2111 ( .A(n997), .B(n2636), .Z(n2635) );
  XOR U2112 ( .A(n2637), .B(n2634), .Z(n2636) );
  XOR U2113 ( .A(n2638), .B(n2639), .Z(n2626) );
  AND U2114 ( .A(n2640), .B(n2641), .Z(n2639) );
  XNOR U2115 ( .A(n2642), .B(n2269), .Z(n2641) );
  XOR U2116 ( .A(n2643), .B(n2644), .Z(n2269) );
  AND U2117 ( .A(n999), .B(n2645), .Z(n2644) );
  XOR U2118 ( .A(n2643), .B(n2646), .Z(n2645) );
  XNOR U2119 ( .A(n2266), .B(n2638), .Z(n2640) );
  XOR U2120 ( .A(n2647), .B(n2648), .Z(n2266) );
  AND U2121 ( .A(n997), .B(n2649), .Z(n2648) );
  XOR U2122 ( .A(n2647), .B(n2650), .Z(n2649) );
  IV U2123 ( .A(n2642), .Z(n2638) );
  AND U2124 ( .A(n2274), .B(n2277), .Z(n2642) );
  XNOR U2125 ( .A(n2651), .B(n2652), .Z(n2277) );
  AND U2126 ( .A(n999), .B(n2653), .Z(n2652) );
  XNOR U2127 ( .A(n2654), .B(n2651), .Z(n2653) );
  XOR U2128 ( .A(n2655), .B(n2656), .Z(n999) );
  AND U2129 ( .A(n2657), .B(n2658), .Z(n2656) );
  XOR U2130 ( .A(n2655), .B(n2285), .Z(n2658) );
  XOR U2131 ( .A(n2659), .B(n2660), .Z(n2285) );
  AND U2132 ( .A(n815), .B(n2661), .Z(n2660) );
  XOR U2133 ( .A(n2662), .B(n2659), .Z(n2661) );
  XNOR U2134 ( .A(n2282), .B(n2655), .Z(n2657) );
  XOR U2135 ( .A(n2663), .B(n2664), .Z(n2282) );
  AND U2136 ( .A(n813), .B(n2665), .Z(n2664) );
  XOR U2137 ( .A(n2666), .B(n2663), .Z(n2665) );
  XOR U2138 ( .A(n2667), .B(n2668), .Z(n2655) );
  AND U2139 ( .A(n2669), .B(n2670), .Z(n2668) );
  XOR U2140 ( .A(n2667), .B(n2297), .Z(n2670) );
  XOR U2141 ( .A(n2671), .B(n2672), .Z(n2297) );
  AND U2142 ( .A(n815), .B(n2673), .Z(n2672) );
  XOR U2143 ( .A(n2674), .B(n2671), .Z(n2673) );
  XNOR U2144 ( .A(n2294), .B(n2667), .Z(n2669) );
  XOR U2145 ( .A(n2675), .B(n2676), .Z(n2294) );
  AND U2146 ( .A(n813), .B(n2677), .Z(n2676) );
  XOR U2147 ( .A(n2678), .B(n2675), .Z(n2677) );
  XOR U2148 ( .A(n2679), .B(n2680), .Z(n2667) );
  AND U2149 ( .A(n2681), .B(n2682), .Z(n2680) );
  XOR U2150 ( .A(n2679), .B(n2309), .Z(n2682) );
  XOR U2151 ( .A(n2683), .B(n2684), .Z(n2309) );
  AND U2152 ( .A(n815), .B(n2685), .Z(n2684) );
  XOR U2153 ( .A(n2686), .B(n2683), .Z(n2685) );
  XNOR U2154 ( .A(n2306), .B(n2679), .Z(n2681) );
  XOR U2155 ( .A(n2687), .B(n2688), .Z(n2306) );
  AND U2156 ( .A(n813), .B(n2689), .Z(n2688) );
  XOR U2157 ( .A(n2690), .B(n2687), .Z(n2689) );
  XOR U2158 ( .A(n2691), .B(n2692), .Z(n2679) );
  AND U2159 ( .A(n2693), .B(n2694), .Z(n2692) );
  XOR U2160 ( .A(n2691), .B(n2321), .Z(n2694) );
  XOR U2161 ( .A(n2695), .B(n2696), .Z(n2321) );
  AND U2162 ( .A(n815), .B(n2697), .Z(n2696) );
  XOR U2163 ( .A(n2698), .B(n2695), .Z(n2697) );
  XNOR U2164 ( .A(n2318), .B(n2691), .Z(n2693) );
  XOR U2165 ( .A(n2699), .B(n2700), .Z(n2318) );
  AND U2166 ( .A(n813), .B(n2701), .Z(n2700) );
  XOR U2167 ( .A(n2702), .B(n2699), .Z(n2701) );
  XOR U2168 ( .A(n2703), .B(n2704), .Z(n2691) );
  AND U2169 ( .A(n2705), .B(n2706), .Z(n2704) );
  XOR U2170 ( .A(n2703), .B(n2333), .Z(n2706) );
  XOR U2171 ( .A(n2707), .B(n2708), .Z(n2333) );
  AND U2172 ( .A(n815), .B(n2709), .Z(n2708) );
  XOR U2173 ( .A(n2710), .B(n2707), .Z(n2709) );
  XNOR U2174 ( .A(n2330), .B(n2703), .Z(n2705) );
  XOR U2175 ( .A(n2711), .B(n2712), .Z(n2330) );
  AND U2176 ( .A(n813), .B(n2713), .Z(n2712) );
  XOR U2177 ( .A(n2714), .B(n2711), .Z(n2713) );
  XOR U2178 ( .A(n2715), .B(n2716), .Z(n2703) );
  AND U2179 ( .A(n2717), .B(n2718), .Z(n2716) );
  XOR U2180 ( .A(n2715), .B(n2345), .Z(n2718) );
  XOR U2181 ( .A(n2719), .B(n2720), .Z(n2345) );
  AND U2182 ( .A(n815), .B(n2721), .Z(n2720) );
  XOR U2183 ( .A(n2722), .B(n2719), .Z(n2721) );
  XNOR U2184 ( .A(n2342), .B(n2715), .Z(n2717) );
  XOR U2185 ( .A(n2723), .B(n2724), .Z(n2342) );
  AND U2186 ( .A(n813), .B(n2725), .Z(n2724) );
  XOR U2187 ( .A(n2726), .B(n2723), .Z(n2725) );
  XOR U2188 ( .A(n2727), .B(n2728), .Z(n2715) );
  AND U2189 ( .A(n2729), .B(n2730), .Z(n2728) );
  XOR U2190 ( .A(n2727), .B(n2357), .Z(n2730) );
  XOR U2191 ( .A(n2731), .B(n2732), .Z(n2357) );
  AND U2192 ( .A(n815), .B(n2733), .Z(n2732) );
  XOR U2193 ( .A(n2734), .B(n2731), .Z(n2733) );
  XNOR U2194 ( .A(n2354), .B(n2727), .Z(n2729) );
  XOR U2195 ( .A(n2735), .B(n2736), .Z(n2354) );
  AND U2196 ( .A(n813), .B(n2737), .Z(n2736) );
  XOR U2197 ( .A(n2738), .B(n2735), .Z(n2737) );
  XOR U2198 ( .A(n2739), .B(n2740), .Z(n2727) );
  AND U2199 ( .A(n2741), .B(n2742), .Z(n2740) );
  XOR U2200 ( .A(n2739), .B(n2369), .Z(n2742) );
  XOR U2201 ( .A(n2743), .B(n2744), .Z(n2369) );
  AND U2202 ( .A(n815), .B(n2745), .Z(n2744) );
  XOR U2203 ( .A(n2746), .B(n2743), .Z(n2745) );
  XNOR U2204 ( .A(n2366), .B(n2739), .Z(n2741) );
  XOR U2205 ( .A(n2747), .B(n2748), .Z(n2366) );
  AND U2206 ( .A(n813), .B(n2749), .Z(n2748) );
  XOR U2207 ( .A(n2750), .B(n2747), .Z(n2749) );
  XOR U2208 ( .A(n2751), .B(n2752), .Z(n2739) );
  AND U2209 ( .A(n2753), .B(n2754), .Z(n2752) );
  XOR U2210 ( .A(n2751), .B(n2381), .Z(n2754) );
  XOR U2211 ( .A(n2755), .B(n2756), .Z(n2381) );
  AND U2212 ( .A(n815), .B(n2757), .Z(n2756) );
  XOR U2213 ( .A(n2758), .B(n2755), .Z(n2757) );
  XNOR U2214 ( .A(n2378), .B(n2751), .Z(n2753) );
  XOR U2215 ( .A(n2759), .B(n2760), .Z(n2378) );
  AND U2216 ( .A(n813), .B(n2761), .Z(n2760) );
  XOR U2217 ( .A(n2762), .B(n2759), .Z(n2761) );
  XOR U2218 ( .A(n2763), .B(n2764), .Z(n2751) );
  AND U2219 ( .A(n2765), .B(n2766), .Z(n2764) );
  XOR U2220 ( .A(n2763), .B(n2393), .Z(n2766) );
  XOR U2221 ( .A(n2767), .B(n2768), .Z(n2393) );
  AND U2222 ( .A(n815), .B(n2769), .Z(n2768) );
  XOR U2223 ( .A(n2770), .B(n2767), .Z(n2769) );
  XNOR U2224 ( .A(n2390), .B(n2763), .Z(n2765) );
  XOR U2225 ( .A(n2771), .B(n2772), .Z(n2390) );
  AND U2226 ( .A(n813), .B(n2773), .Z(n2772) );
  XOR U2227 ( .A(n2774), .B(n2771), .Z(n2773) );
  XOR U2228 ( .A(n2775), .B(n2776), .Z(n2763) );
  AND U2229 ( .A(n2777), .B(n2778), .Z(n2776) );
  XOR U2230 ( .A(n2775), .B(n2405), .Z(n2778) );
  XOR U2231 ( .A(n2779), .B(n2780), .Z(n2405) );
  AND U2232 ( .A(n815), .B(n2781), .Z(n2780) );
  XOR U2233 ( .A(n2782), .B(n2779), .Z(n2781) );
  XNOR U2234 ( .A(n2402), .B(n2775), .Z(n2777) );
  XOR U2235 ( .A(n2783), .B(n2784), .Z(n2402) );
  AND U2236 ( .A(n813), .B(n2785), .Z(n2784) );
  XOR U2237 ( .A(n2786), .B(n2783), .Z(n2785) );
  XOR U2238 ( .A(n2787), .B(n2788), .Z(n2775) );
  AND U2239 ( .A(n2789), .B(n2790), .Z(n2788) );
  XOR U2240 ( .A(n2787), .B(n2417), .Z(n2790) );
  XOR U2241 ( .A(n2791), .B(n2792), .Z(n2417) );
  AND U2242 ( .A(n815), .B(n2793), .Z(n2792) );
  XOR U2243 ( .A(n2794), .B(n2791), .Z(n2793) );
  XNOR U2244 ( .A(n2414), .B(n2787), .Z(n2789) );
  XOR U2245 ( .A(n2795), .B(n2796), .Z(n2414) );
  AND U2246 ( .A(n813), .B(n2797), .Z(n2796) );
  XOR U2247 ( .A(n2798), .B(n2795), .Z(n2797) );
  XOR U2248 ( .A(n2799), .B(n2800), .Z(n2787) );
  AND U2249 ( .A(n2801), .B(n2802), .Z(n2800) );
  XOR U2250 ( .A(n2799), .B(n2429), .Z(n2802) );
  XOR U2251 ( .A(n2803), .B(n2804), .Z(n2429) );
  AND U2252 ( .A(n815), .B(n2805), .Z(n2804) );
  XOR U2253 ( .A(n2806), .B(n2803), .Z(n2805) );
  XNOR U2254 ( .A(n2426), .B(n2799), .Z(n2801) );
  XOR U2255 ( .A(n2807), .B(n2808), .Z(n2426) );
  AND U2256 ( .A(n813), .B(n2809), .Z(n2808) );
  XOR U2257 ( .A(n2810), .B(n2807), .Z(n2809) );
  XOR U2258 ( .A(n2811), .B(n2812), .Z(n2799) );
  AND U2259 ( .A(n2813), .B(n2814), .Z(n2812) );
  XOR U2260 ( .A(n2811), .B(n2441), .Z(n2814) );
  XOR U2261 ( .A(n2815), .B(n2816), .Z(n2441) );
  AND U2262 ( .A(n815), .B(n2817), .Z(n2816) );
  XOR U2263 ( .A(n2818), .B(n2815), .Z(n2817) );
  XNOR U2264 ( .A(n2438), .B(n2811), .Z(n2813) );
  XOR U2265 ( .A(n2819), .B(n2820), .Z(n2438) );
  AND U2266 ( .A(n813), .B(n2821), .Z(n2820) );
  XOR U2267 ( .A(n2822), .B(n2819), .Z(n2821) );
  XOR U2268 ( .A(n2823), .B(n2824), .Z(n2811) );
  AND U2269 ( .A(n2825), .B(n2826), .Z(n2824) );
  XOR U2270 ( .A(n2823), .B(n2453), .Z(n2826) );
  XOR U2271 ( .A(n2827), .B(n2828), .Z(n2453) );
  AND U2272 ( .A(n815), .B(n2829), .Z(n2828) );
  XOR U2273 ( .A(n2830), .B(n2827), .Z(n2829) );
  XNOR U2274 ( .A(n2450), .B(n2823), .Z(n2825) );
  XOR U2275 ( .A(n2831), .B(n2832), .Z(n2450) );
  AND U2276 ( .A(n813), .B(n2833), .Z(n2832) );
  XOR U2277 ( .A(n2834), .B(n2831), .Z(n2833) );
  XOR U2278 ( .A(n2835), .B(n2836), .Z(n2823) );
  AND U2279 ( .A(n2837), .B(n2838), .Z(n2836) );
  XOR U2280 ( .A(n2835), .B(n2465), .Z(n2838) );
  XOR U2281 ( .A(n2839), .B(n2840), .Z(n2465) );
  AND U2282 ( .A(n815), .B(n2841), .Z(n2840) );
  XOR U2283 ( .A(n2842), .B(n2839), .Z(n2841) );
  XNOR U2284 ( .A(n2462), .B(n2835), .Z(n2837) );
  XOR U2285 ( .A(n2843), .B(n2844), .Z(n2462) );
  AND U2286 ( .A(n813), .B(n2845), .Z(n2844) );
  XOR U2287 ( .A(n2846), .B(n2843), .Z(n2845) );
  XOR U2288 ( .A(n2847), .B(n2848), .Z(n2835) );
  AND U2289 ( .A(n2849), .B(n2850), .Z(n2848) );
  XOR U2290 ( .A(n2847), .B(n2477), .Z(n2850) );
  XOR U2291 ( .A(n2851), .B(n2852), .Z(n2477) );
  AND U2292 ( .A(n815), .B(n2853), .Z(n2852) );
  XOR U2293 ( .A(n2854), .B(n2851), .Z(n2853) );
  XNOR U2294 ( .A(n2474), .B(n2847), .Z(n2849) );
  XOR U2295 ( .A(n2855), .B(n2856), .Z(n2474) );
  AND U2296 ( .A(n813), .B(n2857), .Z(n2856) );
  XOR U2297 ( .A(n2858), .B(n2855), .Z(n2857) );
  XOR U2298 ( .A(n2859), .B(n2860), .Z(n2847) );
  AND U2299 ( .A(n2861), .B(n2862), .Z(n2860) );
  XOR U2300 ( .A(n2859), .B(n2489), .Z(n2862) );
  XOR U2301 ( .A(n2863), .B(n2864), .Z(n2489) );
  AND U2302 ( .A(n815), .B(n2865), .Z(n2864) );
  XOR U2303 ( .A(n2866), .B(n2863), .Z(n2865) );
  XNOR U2304 ( .A(n2486), .B(n2859), .Z(n2861) );
  XOR U2305 ( .A(n2867), .B(n2868), .Z(n2486) );
  AND U2306 ( .A(n813), .B(n2869), .Z(n2868) );
  XOR U2307 ( .A(n2870), .B(n2867), .Z(n2869) );
  XOR U2308 ( .A(n2871), .B(n2872), .Z(n2859) );
  AND U2309 ( .A(n2873), .B(n2874), .Z(n2872) );
  XOR U2310 ( .A(n2871), .B(n2501), .Z(n2874) );
  XOR U2311 ( .A(n2875), .B(n2876), .Z(n2501) );
  AND U2312 ( .A(n815), .B(n2877), .Z(n2876) );
  XOR U2313 ( .A(n2878), .B(n2875), .Z(n2877) );
  XNOR U2314 ( .A(n2498), .B(n2871), .Z(n2873) );
  XOR U2315 ( .A(n2879), .B(n2880), .Z(n2498) );
  AND U2316 ( .A(n813), .B(n2881), .Z(n2880) );
  XOR U2317 ( .A(n2882), .B(n2879), .Z(n2881) );
  XOR U2318 ( .A(n2883), .B(n2884), .Z(n2871) );
  AND U2319 ( .A(n2885), .B(n2886), .Z(n2884) );
  XOR U2320 ( .A(n2883), .B(n2513), .Z(n2886) );
  XOR U2321 ( .A(n2887), .B(n2888), .Z(n2513) );
  AND U2322 ( .A(n815), .B(n2889), .Z(n2888) );
  XOR U2323 ( .A(n2890), .B(n2887), .Z(n2889) );
  XNOR U2324 ( .A(n2510), .B(n2883), .Z(n2885) );
  XOR U2325 ( .A(n2891), .B(n2892), .Z(n2510) );
  AND U2326 ( .A(n813), .B(n2893), .Z(n2892) );
  XOR U2327 ( .A(n2894), .B(n2891), .Z(n2893) );
  XOR U2328 ( .A(n2895), .B(n2896), .Z(n2883) );
  AND U2329 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR U2330 ( .A(n2895), .B(n2525), .Z(n2898) );
  XOR U2331 ( .A(n2899), .B(n2900), .Z(n2525) );
  AND U2332 ( .A(n815), .B(n2901), .Z(n2900) );
  XOR U2333 ( .A(n2902), .B(n2899), .Z(n2901) );
  XNOR U2334 ( .A(n2522), .B(n2895), .Z(n2897) );
  XOR U2335 ( .A(n2903), .B(n2904), .Z(n2522) );
  AND U2336 ( .A(n813), .B(n2905), .Z(n2904) );
  XOR U2337 ( .A(n2906), .B(n2903), .Z(n2905) );
  XOR U2338 ( .A(n2907), .B(n2908), .Z(n2895) );
  AND U2339 ( .A(n2909), .B(n2910), .Z(n2908) );
  XOR U2340 ( .A(n2907), .B(n2537), .Z(n2910) );
  XOR U2341 ( .A(n2911), .B(n2912), .Z(n2537) );
  AND U2342 ( .A(n815), .B(n2913), .Z(n2912) );
  XOR U2343 ( .A(n2914), .B(n2911), .Z(n2913) );
  XNOR U2344 ( .A(n2534), .B(n2907), .Z(n2909) );
  XOR U2345 ( .A(n2915), .B(n2916), .Z(n2534) );
  AND U2346 ( .A(n813), .B(n2917), .Z(n2916) );
  XOR U2347 ( .A(n2918), .B(n2915), .Z(n2917) );
  XOR U2348 ( .A(n2919), .B(n2920), .Z(n2907) );
  AND U2349 ( .A(n2921), .B(n2922), .Z(n2920) );
  XOR U2350 ( .A(n2919), .B(n2549), .Z(n2922) );
  XOR U2351 ( .A(n2923), .B(n2924), .Z(n2549) );
  AND U2352 ( .A(n815), .B(n2925), .Z(n2924) );
  XOR U2353 ( .A(n2926), .B(n2923), .Z(n2925) );
  XNOR U2354 ( .A(n2546), .B(n2919), .Z(n2921) );
  XOR U2355 ( .A(n2927), .B(n2928), .Z(n2546) );
  AND U2356 ( .A(n813), .B(n2929), .Z(n2928) );
  XOR U2357 ( .A(n2930), .B(n2927), .Z(n2929) );
  XOR U2358 ( .A(n2931), .B(n2932), .Z(n2919) );
  AND U2359 ( .A(n2933), .B(n2934), .Z(n2932) );
  XOR U2360 ( .A(n2931), .B(n2561), .Z(n2934) );
  XOR U2361 ( .A(n2935), .B(n2936), .Z(n2561) );
  AND U2362 ( .A(n815), .B(n2937), .Z(n2936) );
  XOR U2363 ( .A(n2938), .B(n2935), .Z(n2937) );
  XNOR U2364 ( .A(n2558), .B(n2931), .Z(n2933) );
  XOR U2365 ( .A(n2939), .B(n2940), .Z(n2558) );
  AND U2366 ( .A(n813), .B(n2941), .Z(n2940) );
  XOR U2367 ( .A(n2942), .B(n2939), .Z(n2941) );
  XOR U2368 ( .A(n2943), .B(n2944), .Z(n2931) );
  AND U2369 ( .A(n2945), .B(n2946), .Z(n2944) );
  XOR U2370 ( .A(n2943), .B(n2573), .Z(n2946) );
  XOR U2371 ( .A(n2947), .B(n2948), .Z(n2573) );
  AND U2372 ( .A(n815), .B(n2949), .Z(n2948) );
  XOR U2373 ( .A(n2950), .B(n2947), .Z(n2949) );
  XNOR U2374 ( .A(n2570), .B(n2943), .Z(n2945) );
  XOR U2375 ( .A(n2951), .B(n2952), .Z(n2570) );
  AND U2376 ( .A(n813), .B(n2953), .Z(n2952) );
  XOR U2377 ( .A(n2954), .B(n2951), .Z(n2953) );
  XOR U2378 ( .A(n2955), .B(n2956), .Z(n2943) );
  AND U2379 ( .A(n2957), .B(n2958), .Z(n2956) );
  XOR U2380 ( .A(n2955), .B(n2585), .Z(n2958) );
  XOR U2381 ( .A(n2959), .B(n2960), .Z(n2585) );
  AND U2382 ( .A(n815), .B(n2961), .Z(n2960) );
  XOR U2383 ( .A(n2962), .B(n2959), .Z(n2961) );
  XNOR U2384 ( .A(n2582), .B(n2955), .Z(n2957) );
  XOR U2385 ( .A(n2963), .B(n2964), .Z(n2582) );
  AND U2386 ( .A(n813), .B(n2965), .Z(n2964) );
  XOR U2387 ( .A(n2966), .B(n2963), .Z(n2965) );
  XOR U2388 ( .A(n2967), .B(n2968), .Z(n2955) );
  AND U2389 ( .A(n2969), .B(n2970), .Z(n2968) );
  XOR U2390 ( .A(n2967), .B(n2597), .Z(n2970) );
  XOR U2391 ( .A(n2971), .B(n2972), .Z(n2597) );
  AND U2392 ( .A(n815), .B(n2973), .Z(n2972) );
  XOR U2393 ( .A(n2974), .B(n2971), .Z(n2973) );
  XNOR U2394 ( .A(n2594), .B(n2967), .Z(n2969) );
  XOR U2395 ( .A(n2975), .B(n2976), .Z(n2594) );
  AND U2396 ( .A(n813), .B(n2977), .Z(n2976) );
  XOR U2397 ( .A(n2978), .B(n2975), .Z(n2977) );
  XOR U2398 ( .A(n2979), .B(n2980), .Z(n2967) );
  AND U2399 ( .A(n2981), .B(n2982), .Z(n2980) );
  XOR U2400 ( .A(n2979), .B(n2609), .Z(n2982) );
  XOR U2401 ( .A(n2983), .B(n2984), .Z(n2609) );
  AND U2402 ( .A(n815), .B(n2985), .Z(n2984) );
  XOR U2403 ( .A(n2986), .B(n2983), .Z(n2985) );
  XNOR U2404 ( .A(n2606), .B(n2979), .Z(n2981) );
  XOR U2405 ( .A(n2987), .B(n2988), .Z(n2606) );
  AND U2406 ( .A(n813), .B(n2989), .Z(n2988) );
  XOR U2407 ( .A(n2990), .B(n2987), .Z(n2989) );
  XOR U2408 ( .A(n2991), .B(n2992), .Z(n2979) );
  AND U2409 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U2410 ( .A(n2991), .B(n2621), .Z(n2994) );
  XOR U2411 ( .A(n2995), .B(n2996), .Z(n2621) );
  AND U2412 ( .A(n815), .B(n2997), .Z(n2996) );
  XOR U2413 ( .A(n2998), .B(n2995), .Z(n2997) );
  XNOR U2414 ( .A(n2618), .B(n2991), .Z(n2993) );
  XOR U2415 ( .A(n2999), .B(n3000), .Z(n2618) );
  AND U2416 ( .A(n813), .B(n3001), .Z(n3000) );
  XOR U2417 ( .A(n3002), .B(n2999), .Z(n3001) );
  XOR U2418 ( .A(n3003), .B(n3004), .Z(n2991) );
  AND U2419 ( .A(n3005), .B(n3006), .Z(n3004) );
  XOR U2420 ( .A(n3003), .B(n2633), .Z(n3006) );
  XOR U2421 ( .A(n3007), .B(n3008), .Z(n2633) );
  AND U2422 ( .A(n815), .B(n3009), .Z(n3008) );
  XOR U2423 ( .A(n3010), .B(n3007), .Z(n3009) );
  XNOR U2424 ( .A(n2630), .B(n3003), .Z(n3005) );
  XOR U2425 ( .A(n3011), .B(n3012), .Z(n2630) );
  AND U2426 ( .A(n813), .B(n3013), .Z(n3012) );
  XOR U2427 ( .A(n3014), .B(n3011), .Z(n3013) );
  XOR U2428 ( .A(n3015), .B(n3016), .Z(n3003) );
  AND U2429 ( .A(n3017), .B(n3018), .Z(n3016) );
  XNOR U2430 ( .A(n3019), .B(n2646), .Z(n3018) );
  XOR U2431 ( .A(n3020), .B(n3021), .Z(n2646) );
  AND U2432 ( .A(n815), .B(n3022), .Z(n3021) );
  XOR U2433 ( .A(n3020), .B(n3023), .Z(n3022) );
  XNOR U2434 ( .A(n2643), .B(n3015), .Z(n3017) );
  XOR U2435 ( .A(n3024), .B(n3025), .Z(n2643) );
  AND U2436 ( .A(n813), .B(n3026), .Z(n3025) );
  XOR U2437 ( .A(n3024), .B(n3027), .Z(n3026) );
  IV U2438 ( .A(n3019), .Z(n3015) );
  AND U2439 ( .A(n2651), .B(n2654), .Z(n3019) );
  XNOR U2440 ( .A(n3028), .B(n3029), .Z(n2654) );
  AND U2441 ( .A(n815), .B(n3030), .Z(n3029) );
  XNOR U2442 ( .A(n3031), .B(n3028), .Z(n3030) );
  XOR U2443 ( .A(n3032), .B(n3033), .Z(n815) );
  AND U2444 ( .A(n3034), .B(n3035), .Z(n3033) );
  XOR U2445 ( .A(n3032), .B(n2662), .Z(n3035) );
  XNOR U2446 ( .A(n3036), .B(n3037), .Z(n2662) );
  AND U2447 ( .A(n3038), .B(n439), .Z(n3037) );
  AND U2448 ( .A(n3036), .B(n3039), .Z(n3038) );
  XNOR U2449 ( .A(n2659), .B(n3032), .Z(n3034) );
  XOR U2450 ( .A(n3040), .B(n3041), .Z(n2659) );
  AND U2451 ( .A(n3042), .B(n437), .Z(n3041) );
  NOR U2452 ( .A(n3040), .B(n3043), .Z(n3042) );
  XOR U2453 ( .A(n3044), .B(n3045), .Z(n3032) );
  AND U2454 ( .A(n3046), .B(n3047), .Z(n3045) );
  XOR U2455 ( .A(n3044), .B(n2674), .Z(n3047) );
  XOR U2456 ( .A(n3048), .B(n3049), .Z(n2674) );
  AND U2457 ( .A(n439), .B(n3050), .Z(n3049) );
  XOR U2458 ( .A(n3051), .B(n3048), .Z(n3050) );
  XNOR U2459 ( .A(n2671), .B(n3044), .Z(n3046) );
  XOR U2460 ( .A(n3052), .B(n3053), .Z(n2671) );
  AND U2461 ( .A(n437), .B(n3054), .Z(n3053) );
  XOR U2462 ( .A(n3055), .B(n3052), .Z(n3054) );
  XOR U2463 ( .A(n3056), .B(n3057), .Z(n3044) );
  AND U2464 ( .A(n3058), .B(n3059), .Z(n3057) );
  XOR U2465 ( .A(n3056), .B(n2686), .Z(n3059) );
  XOR U2466 ( .A(n3060), .B(n3061), .Z(n2686) );
  AND U2467 ( .A(n439), .B(n3062), .Z(n3061) );
  XOR U2468 ( .A(n3063), .B(n3060), .Z(n3062) );
  XNOR U2469 ( .A(n2683), .B(n3056), .Z(n3058) );
  XOR U2470 ( .A(n3064), .B(n3065), .Z(n2683) );
  AND U2471 ( .A(n437), .B(n3066), .Z(n3065) );
  XOR U2472 ( .A(n3067), .B(n3064), .Z(n3066) );
  XOR U2473 ( .A(n3068), .B(n3069), .Z(n3056) );
  AND U2474 ( .A(n3070), .B(n3071), .Z(n3069) );
  XOR U2475 ( .A(n3068), .B(n2698), .Z(n3071) );
  XOR U2476 ( .A(n3072), .B(n3073), .Z(n2698) );
  AND U2477 ( .A(n439), .B(n3074), .Z(n3073) );
  XOR U2478 ( .A(n3075), .B(n3072), .Z(n3074) );
  XNOR U2479 ( .A(n2695), .B(n3068), .Z(n3070) );
  XOR U2480 ( .A(n3076), .B(n3077), .Z(n2695) );
  AND U2481 ( .A(n437), .B(n3078), .Z(n3077) );
  XOR U2482 ( .A(n3079), .B(n3076), .Z(n3078) );
  XOR U2483 ( .A(n3080), .B(n3081), .Z(n3068) );
  AND U2484 ( .A(n3082), .B(n3083), .Z(n3081) );
  XOR U2485 ( .A(n3080), .B(n2710), .Z(n3083) );
  XOR U2486 ( .A(n3084), .B(n3085), .Z(n2710) );
  AND U2487 ( .A(n439), .B(n3086), .Z(n3085) );
  XOR U2488 ( .A(n3087), .B(n3084), .Z(n3086) );
  XNOR U2489 ( .A(n2707), .B(n3080), .Z(n3082) );
  XOR U2490 ( .A(n3088), .B(n3089), .Z(n2707) );
  AND U2491 ( .A(n437), .B(n3090), .Z(n3089) );
  XOR U2492 ( .A(n3091), .B(n3088), .Z(n3090) );
  XOR U2493 ( .A(n3092), .B(n3093), .Z(n3080) );
  AND U2494 ( .A(n3094), .B(n3095), .Z(n3093) );
  XOR U2495 ( .A(n3092), .B(n2722), .Z(n3095) );
  XOR U2496 ( .A(n3096), .B(n3097), .Z(n2722) );
  AND U2497 ( .A(n439), .B(n3098), .Z(n3097) );
  XOR U2498 ( .A(n3099), .B(n3096), .Z(n3098) );
  XNOR U2499 ( .A(n2719), .B(n3092), .Z(n3094) );
  XOR U2500 ( .A(n3100), .B(n3101), .Z(n2719) );
  AND U2501 ( .A(n437), .B(n3102), .Z(n3101) );
  XOR U2502 ( .A(n3103), .B(n3100), .Z(n3102) );
  XOR U2503 ( .A(n3104), .B(n3105), .Z(n3092) );
  AND U2504 ( .A(n3106), .B(n3107), .Z(n3105) );
  XOR U2505 ( .A(n3104), .B(n2734), .Z(n3107) );
  XOR U2506 ( .A(n3108), .B(n3109), .Z(n2734) );
  AND U2507 ( .A(n439), .B(n3110), .Z(n3109) );
  XOR U2508 ( .A(n3111), .B(n3108), .Z(n3110) );
  XNOR U2509 ( .A(n2731), .B(n3104), .Z(n3106) );
  XOR U2510 ( .A(n3112), .B(n3113), .Z(n2731) );
  AND U2511 ( .A(n437), .B(n3114), .Z(n3113) );
  XOR U2512 ( .A(n3115), .B(n3112), .Z(n3114) );
  XOR U2513 ( .A(n3116), .B(n3117), .Z(n3104) );
  AND U2514 ( .A(n3118), .B(n3119), .Z(n3117) );
  XOR U2515 ( .A(n3116), .B(n2746), .Z(n3119) );
  XOR U2516 ( .A(n3120), .B(n3121), .Z(n2746) );
  AND U2517 ( .A(n439), .B(n3122), .Z(n3121) );
  XOR U2518 ( .A(n3123), .B(n3120), .Z(n3122) );
  XNOR U2519 ( .A(n2743), .B(n3116), .Z(n3118) );
  XOR U2520 ( .A(n3124), .B(n3125), .Z(n2743) );
  AND U2521 ( .A(n437), .B(n3126), .Z(n3125) );
  XOR U2522 ( .A(n3127), .B(n3124), .Z(n3126) );
  XOR U2523 ( .A(n3128), .B(n3129), .Z(n3116) );
  AND U2524 ( .A(n3130), .B(n3131), .Z(n3129) );
  XOR U2525 ( .A(n3128), .B(n2758), .Z(n3131) );
  XOR U2526 ( .A(n3132), .B(n3133), .Z(n2758) );
  AND U2527 ( .A(n439), .B(n3134), .Z(n3133) );
  XOR U2528 ( .A(n3135), .B(n3132), .Z(n3134) );
  XNOR U2529 ( .A(n2755), .B(n3128), .Z(n3130) );
  XOR U2530 ( .A(n3136), .B(n3137), .Z(n2755) );
  AND U2531 ( .A(n437), .B(n3138), .Z(n3137) );
  XOR U2532 ( .A(n3139), .B(n3136), .Z(n3138) );
  XOR U2533 ( .A(n3140), .B(n3141), .Z(n3128) );
  AND U2534 ( .A(n3142), .B(n3143), .Z(n3141) );
  XOR U2535 ( .A(n3140), .B(n2770), .Z(n3143) );
  XOR U2536 ( .A(n3144), .B(n3145), .Z(n2770) );
  AND U2537 ( .A(n439), .B(n3146), .Z(n3145) );
  XOR U2538 ( .A(n3147), .B(n3144), .Z(n3146) );
  XNOR U2539 ( .A(n2767), .B(n3140), .Z(n3142) );
  XOR U2540 ( .A(n3148), .B(n3149), .Z(n2767) );
  AND U2541 ( .A(n437), .B(n3150), .Z(n3149) );
  XOR U2542 ( .A(n3151), .B(n3148), .Z(n3150) );
  XOR U2543 ( .A(n3152), .B(n3153), .Z(n3140) );
  AND U2544 ( .A(n3154), .B(n3155), .Z(n3153) );
  XOR U2545 ( .A(n3152), .B(n2782), .Z(n3155) );
  XOR U2546 ( .A(n3156), .B(n3157), .Z(n2782) );
  AND U2547 ( .A(n439), .B(n3158), .Z(n3157) );
  XOR U2548 ( .A(n3159), .B(n3156), .Z(n3158) );
  XNOR U2549 ( .A(n2779), .B(n3152), .Z(n3154) );
  XOR U2550 ( .A(n3160), .B(n3161), .Z(n2779) );
  AND U2551 ( .A(n437), .B(n3162), .Z(n3161) );
  XOR U2552 ( .A(n3163), .B(n3160), .Z(n3162) );
  XOR U2553 ( .A(n3164), .B(n3165), .Z(n3152) );
  AND U2554 ( .A(n3166), .B(n3167), .Z(n3165) );
  XOR U2555 ( .A(n3164), .B(n2794), .Z(n3167) );
  XOR U2556 ( .A(n3168), .B(n3169), .Z(n2794) );
  AND U2557 ( .A(n439), .B(n3170), .Z(n3169) );
  XOR U2558 ( .A(n3171), .B(n3168), .Z(n3170) );
  XNOR U2559 ( .A(n2791), .B(n3164), .Z(n3166) );
  XOR U2560 ( .A(n3172), .B(n3173), .Z(n2791) );
  AND U2561 ( .A(n437), .B(n3174), .Z(n3173) );
  XOR U2562 ( .A(n3175), .B(n3172), .Z(n3174) );
  XOR U2563 ( .A(n3176), .B(n3177), .Z(n3164) );
  AND U2564 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U2565 ( .A(n3176), .B(n2806), .Z(n3179) );
  XOR U2566 ( .A(n3180), .B(n3181), .Z(n2806) );
  AND U2567 ( .A(n439), .B(n3182), .Z(n3181) );
  XOR U2568 ( .A(n3183), .B(n3180), .Z(n3182) );
  XNOR U2569 ( .A(n2803), .B(n3176), .Z(n3178) );
  XOR U2570 ( .A(n3184), .B(n3185), .Z(n2803) );
  AND U2571 ( .A(n437), .B(n3186), .Z(n3185) );
  XOR U2572 ( .A(n3187), .B(n3184), .Z(n3186) );
  XOR U2573 ( .A(n3188), .B(n3189), .Z(n3176) );
  AND U2574 ( .A(n3190), .B(n3191), .Z(n3189) );
  XOR U2575 ( .A(n3188), .B(n2818), .Z(n3191) );
  XOR U2576 ( .A(n3192), .B(n3193), .Z(n2818) );
  AND U2577 ( .A(n439), .B(n3194), .Z(n3193) );
  XOR U2578 ( .A(n3195), .B(n3192), .Z(n3194) );
  XNOR U2579 ( .A(n2815), .B(n3188), .Z(n3190) );
  XOR U2580 ( .A(n3196), .B(n3197), .Z(n2815) );
  AND U2581 ( .A(n437), .B(n3198), .Z(n3197) );
  XOR U2582 ( .A(n3199), .B(n3196), .Z(n3198) );
  XOR U2583 ( .A(n3200), .B(n3201), .Z(n3188) );
  AND U2584 ( .A(n3202), .B(n3203), .Z(n3201) );
  XOR U2585 ( .A(n3200), .B(n2830), .Z(n3203) );
  XOR U2586 ( .A(n3204), .B(n3205), .Z(n2830) );
  AND U2587 ( .A(n439), .B(n3206), .Z(n3205) );
  XOR U2588 ( .A(n3207), .B(n3204), .Z(n3206) );
  XNOR U2589 ( .A(n2827), .B(n3200), .Z(n3202) );
  XOR U2590 ( .A(n3208), .B(n3209), .Z(n2827) );
  AND U2591 ( .A(n437), .B(n3210), .Z(n3209) );
  XOR U2592 ( .A(n3211), .B(n3208), .Z(n3210) );
  XOR U2593 ( .A(n3212), .B(n3213), .Z(n3200) );
  AND U2594 ( .A(n3214), .B(n3215), .Z(n3213) );
  XOR U2595 ( .A(n3212), .B(n2842), .Z(n3215) );
  XOR U2596 ( .A(n3216), .B(n3217), .Z(n2842) );
  AND U2597 ( .A(n439), .B(n3218), .Z(n3217) );
  XOR U2598 ( .A(n3219), .B(n3216), .Z(n3218) );
  XNOR U2599 ( .A(n2839), .B(n3212), .Z(n3214) );
  XOR U2600 ( .A(n3220), .B(n3221), .Z(n2839) );
  AND U2601 ( .A(n437), .B(n3222), .Z(n3221) );
  XOR U2602 ( .A(n3223), .B(n3220), .Z(n3222) );
  XOR U2603 ( .A(n3224), .B(n3225), .Z(n3212) );
  AND U2604 ( .A(n3226), .B(n3227), .Z(n3225) );
  XOR U2605 ( .A(n3224), .B(n2854), .Z(n3227) );
  XOR U2606 ( .A(n3228), .B(n3229), .Z(n2854) );
  AND U2607 ( .A(n439), .B(n3230), .Z(n3229) );
  XOR U2608 ( .A(n3231), .B(n3228), .Z(n3230) );
  XNOR U2609 ( .A(n2851), .B(n3224), .Z(n3226) );
  XOR U2610 ( .A(n3232), .B(n3233), .Z(n2851) );
  AND U2611 ( .A(n437), .B(n3234), .Z(n3233) );
  XOR U2612 ( .A(n3235), .B(n3232), .Z(n3234) );
  XOR U2613 ( .A(n3236), .B(n3237), .Z(n3224) );
  AND U2614 ( .A(n3238), .B(n3239), .Z(n3237) );
  XOR U2615 ( .A(n3236), .B(n2866), .Z(n3239) );
  XOR U2616 ( .A(n3240), .B(n3241), .Z(n2866) );
  AND U2617 ( .A(n439), .B(n3242), .Z(n3241) );
  XOR U2618 ( .A(n3243), .B(n3240), .Z(n3242) );
  XNOR U2619 ( .A(n2863), .B(n3236), .Z(n3238) );
  XOR U2620 ( .A(n3244), .B(n3245), .Z(n2863) );
  AND U2621 ( .A(n437), .B(n3246), .Z(n3245) );
  XOR U2622 ( .A(n3247), .B(n3244), .Z(n3246) );
  XOR U2623 ( .A(n3248), .B(n3249), .Z(n3236) );
  AND U2624 ( .A(n3250), .B(n3251), .Z(n3249) );
  XOR U2625 ( .A(n3248), .B(n2878), .Z(n3251) );
  XOR U2626 ( .A(n3252), .B(n3253), .Z(n2878) );
  AND U2627 ( .A(n439), .B(n3254), .Z(n3253) );
  XOR U2628 ( .A(n3255), .B(n3252), .Z(n3254) );
  XNOR U2629 ( .A(n2875), .B(n3248), .Z(n3250) );
  XOR U2630 ( .A(n3256), .B(n3257), .Z(n2875) );
  AND U2631 ( .A(n437), .B(n3258), .Z(n3257) );
  XOR U2632 ( .A(n3259), .B(n3256), .Z(n3258) );
  XOR U2633 ( .A(n3260), .B(n3261), .Z(n3248) );
  AND U2634 ( .A(n3262), .B(n3263), .Z(n3261) );
  XOR U2635 ( .A(n3260), .B(n2890), .Z(n3263) );
  XOR U2636 ( .A(n3264), .B(n3265), .Z(n2890) );
  AND U2637 ( .A(n439), .B(n3266), .Z(n3265) );
  XOR U2638 ( .A(n3267), .B(n3264), .Z(n3266) );
  XNOR U2639 ( .A(n2887), .B(n3260), .Z(n3262) );
  XOR U2640 ( .A(n3268), .B(n3269), .Z(n2887) );
  AND U2641 ( .A(n437), .B(n3270), .Z(n3269) );
  XOR U2642 ( .A(n3271), .B(n3268), .Z(n3270) );
  XOR U2643 ( .A(n3272), .B(n3273), .Z(n3260) );
  AND U2644 ( .A(n3274), .B(n3275), .Z(n3273) );
  XOR U2645 ( .A(n3272), .B(n2902), .Z(n3275) );
  XOR U2646 ( .A(n3276), .B(n3277), .Z(n2902) );
  AND U2647 ( .A(n439), .B(n3278), .Z(n3277) );
  XOR U2648 ( .A(n3279), .B(n3276), .Z(n3278) );
  XNOR U2649 ( .A(n2899), .B(n3272), .Z(n3274) );
  XOR U2650 ( .A(n3280), .B(n3281), .Z(n2899) );
  AND U2651 ( .A(n437), .B(n3282), .Z(n3281) );
  XOR U2652 ( .A(n3283), .B(n3280), .Z(n3282) );
  XOR U2653 ( .A(n3284), .B(n3285), .Z(n3272) );
  AND U2654 ( .A(n3286), .B(n3287), .Z(n3285) );
  XOR U2655 ( .A(n3284), .B(n2914), .Z(n3287) );
  XOR U2656 ( .A(n3288), .B(n3289), .Z(n2914) );
  AND U2657 ( .A(n439), .B(n3290), .Z(n3289) );
  XOR U2658 ( .A(n3291), .B(n3288), .Z(n3290) );
  XNOR U2659 ( .A(n2911), .B(n3284), .Z(n3286) );
  XOR U2660 ( .A(n3292), .B(n3293), .Z(n2911) );
  AND U2661 ( .A(n437), .B(n3294), .Z(n3293) );
  XOR U2662 ( .A(n3295), .B(n3292), .Z(n3294) );
  XOR U2663 ( .A(n3296), .B(n3297), .Z(n3284) );
  AND U2664 ( .A(n3298), .B(n3299), .Z(n3297) );
  XOR U2665 ( .A(n3296), .B(n2926), .Z(n3299) );
  XOR U2666 ( .A(n3300), .B(n3301), .Z(n2926) );
  AND U2667 ( .A(n439), .B(n3302), .Z(n3301) );
  XOR U2668 ( .A(n3303), .B(n3300), .Z(n3302) );
  XNOR U2669 ( .A(n2923), .B(n3296), .Z(n3298) );
  XOR U2670 ( .A(n3304), .B(n3305), .Z(n2923) );
  AND U2671 ( .A(n437), .B(n3306), .Z(n3305) );
  XOR U2672 ( .A(n3307), .B(n3304), .Z(n3306) );
  XOR U2673 ( .A(n3308), .B(n3309), .Z(n3296) );
  AND U2674 ( .A(n3310), .B(n3311), .Z(n3309) );
  XOR U2675 ( .A(n3308), .B(n2938), .Z(n3311) );
  XOR U2676 ( .A(n3312), .B(n3313), .Z(n2938) );
  AND U2677 ( .A(n439), .B(n3314), .Z(n3313) );
  XOR U2678 ( .A(n3315), .B(n3312), .Z(n3314) );
  XNOR U2679 ( .A(n2935), .B(n3308), .Z(n3310) );
  XOR U2680 ( .A(n3316), .B(n3317), .Z(n2935) );
  AND U2681 ( .A(n437), .B(n3318), .Z(n3317) );
  XOR U2682 ( .A(n3319), .B(n3316), .Z(n3318) );
  XOR U2683 ( .A(n3320), .B(n3321), .Z(n3308) );
  AND U2684 ( .A(n3322), .B(n3323), .Z(n3321) );
  XOR U2685 ( .A(n3320), .B(n2950), .Z(n3323) );
  XOR U2686 ( .A(n3324), .B(n3325), .Z(n2950) );
  AND U2687 ( .A(n439), .B(n3326), .Z(n3325) );
  XOR U2688 ( .A(n3327), .B(n3324), .Z(n3326) );
  XNOR U2689 ( .A(n2947), .B(n3320), .Z(n3322) );
  XOR U2690 ( .A(n3328), .B(n3329), .Z(n2947) );
  AND U2691 ( .A(n437), .B(n3330), .Z(n3329) );
  XOR U2692 ( .A(n3331), .B(n3328), .Z(n3330) );
  XOR U2693 ( .A(n3332), .B(n3333), .Z(n3320) );
  AND U2694 ( .A(n3334), .B(n3335), .Z(n3333) );
  XOR U2695 ( .A(n3332), .B(n2962), .Z(n3335) );
  XOR U2696 ( .A(n3336), .B(n3337), .Z(n2962) );
  AND U2697 ( .A(n439), .B(n3338), .Z(n3337) );
  XOR U2698 ( .A(n3339), .B(n3336), .Z(n3338) );
  XNOR U2699 ( .A(n2959), .B(n3332), .Z(n3334) );
  XOR U2700 ( .A(n3340), .B(n3341), .Z(n2959) );
  AND U2701 ( .A(n437), .B(n3342), .Z(n3341) );
  XOR U2702 ( .A(n3343), .B(n3340), .Z(n3342) );
  XOR U2703 ( .A(n3344), .B(n3345), .Z(n3332) );
  AND U2704 ( .A(n3346), .B(n3347), .Z(n3345) );
  XOR U2705 ( .A(n3344), .B(n2974), .Z(n3347) );
  XOR U2706 ( .A(n3348), .B(n3349), .Z(n2974) );
  AND U2707 ( .A(n439), .B(n3350), .Z(n3349) );
  XOR U2708 ( .A(n3351), .B(n3348), .Z(n3350) );
  XNOR U2709 ( .A(n2971), .B(n3344), .Z(n3346) );
  XOR U2710 ( .A(n3352), .B(n3353), .Z(n2971) );
  AND U2711 ( .A(n437), .B(n3354), .Z(n3353) );
  XOR U2712 ( .A(n3355), .B(n3352), .Z(n3354) );
  XOR U2713 ( .A(n3356), .B(n3357), .Z(n3344) );
  AND U2714 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR U2715 ( .A(n3356), .B(n2986), .Z(n3359) );
  XOR U2716 ( .A(n3360), .B(n3361), .Z(n2986) );
  AND U2717 ( .A(n439), .B(n3362), .Z(n3361) );
  XOR U2718 ( .A(n3363), .B(n3360), .Z(n3362) );
  XNOR U2719 ( .A(n2983), .B(n3356), .Z(n3358) );
  XOR U2720 ( .A(n3364), .B(n3365), .Z(n2983) );
  AND U2721 ( .A(n437), .B(n3366), .Z(n3365) );
  XOR U2722 ( .A(n3367), .B(n3364), .Z(n3366) );
  XOR U2723 ( .A(n3368), .B(n3369), .Z(n3356) );
  AND U2724 ( .A(n3370), .B(n3371), .Z(n3369) );
  XOR U2725 ( .A(n3368), .B(n2998), .Z(n3371) );
  XOR U2726 ( .A(n3372), .B(n3373), .Z(n2998) );
  AND U2727 ( .A(n439), .B(n3374), .Z(n3373) );
  XOR U2728 ( .A(n3375), .B(n3372), .Z(n3374) );
  XNOR U2729 ( .A(n2995), .B(n3368), .Z(n3370) );
  XOR U2730 ( .A(n3376), .B(n3377), .Z(n2995) );
  AND U2731 ( .A(n437), .B(n3378), .Z(n3377) );
  XOR U2732 ( .A(n3379), .B(n3376), .Z(n3378) );
  XOR U2733 ( .A(n3380), .B(n3381), .Z(n3368) );
  AND U2734 ( .A(n3382), .B(n3383), .Z(n3381) );
  XOR U2735 ( .A(n3380), .B(n3010), .Z(n3383) );
  XOR U2736 ( .A(n3384), .B(n3385), .Z(n3010) );
  AND U2737 ( .A(n439), .B(n3386), .Z(n3385) );
  XOR U2738 ( .A(n3387), .B(n3384), .Z(n3386) );
  XNOR U2739 ( .A(n3007), .B(n3380), .Z(n3382) );
  XOR U2740 ( .A(n3388), .B(n3389), .Z(n3007) );
  AND U2741 ( .A(n437), .B(n3390), .Z(n3389) );
  XOR U2742 ( .A(n3391), .B(n3388), .Z(n3390) );
  XOR U2743 ( .A(n3392), .B(n3393), .Z(n3380) );
  AND U2744 ( .A(n3394), .B(n3395), .Z(n3393) );
  XNOR U2745 ( .A(n3396), .B(n3023), .Z(n3395) );
  XOR U2746 ( .A(n3397), .B(n3398), .Z(n3023) );
  AND U2747 ( .A(n439), .B(n3399), .Z(n3398) );
  XOR U2748 ( .A(n3397), .B(n3400), .Z(n3399) );
  XNOR U2749 ( .A(n3020), .B(n3392), .Z(n3394) );
  XOR U2750 ( .A(n3401), .B(n3402), .Z(n3020) );
  AND U2751 ( .A(n437), .B(n3403), .Z(n3402) );
  XOR U2752 ( .A(n3401), .B(n3404), .Z(n3403) );
  IV U2753 ( .A(n3396), .Z(n3392) );
  AND U2754 ( .A(n3028), .B(n3031), .Z(n3396) );
  XNOR U2755 ( .A(n3405), .B(n3406), .Z(n3031) );
  AND U2756 ( .A(n439), .B(n3407), .Z(n3406) );
  XNOR U2757 ( .A(n3408), .B(n3405), .Z(n3407) );
  XOR U2758 ( .A(n3409), .B(n3410), .Z(n439) );
  AND U2759 ( .A(n3411), .B(n3412), .Z(n3410) );
  XOR U2760 ( .A(n3039), .B(n3409), .Z(n3412) );
  IV U2761 ( .A(n3413), .Z(n3039) );
  AND U2762 ( .A(p_input[8191]), .B(p_input[8159]), .Z(n3413) );
  XOR U2763 ( .A(n3409), .B(n3036), .Z(n3411) );
  AND U2764 ( .A(p_input[8095]), .B(p_input[8127]), .Z(n3036) );
  XOR U2765 ( .A(n3414), .B(n3415), .Z(n3409) );
  AND U2766 ( .A(n3416), .B(n3417), .Z(n3415) );
  XOR U2767 ( .A(n3414), .B(n3051), .Z(n3417) );
  XNOR U2768 ( .A(p_input[8158]), .B(n3418), .Z(n3051) );
  AND U2769 ( .A(n187), .B(n3419), .Z(n3418) );
  XOR U2770 ( .A(p_input[8190]), .B(p_input[8158]), .Z(n3419) );
  XNOR U2771 ( .A(n3048), .B(n3414), .Z(n3416) );
  XOR U2772 ( .A(n3420), .B(n3421), .Z(n3048) );
  AND U2773 ( .A(n185), .B(n3422), .Z(n3421) );
  XOR U2774 ( .A(p_input[8126]), .B(p_input[8094]), .Z(n3422) );
  XOR U2775 ( .A(n3423), .B(n3424), .Z(n3414) );
  AND U2776 ( .A(n3425), .B(n3426), .Z(n3424) );
  XOR U2777 ( .A(n3423), .B(n3063), .Z(n3426) );
  XNOR U2778 ( .A(p_input[8157]), .B(n3427), .Z(n3063) );
  AND U2779 ( .A(n187), .B(n3428), .Z(n3427) );
  XOR U2780 ( .A(p_input[8189]), .B(p_input[8157]), .Z(n3428) );
  XNOR U2781 ( .A(n3060), .B(n3423), .Z(n3425) );
  XOR U2782 ( .A(n3429), .B(n3430), .Z(n3060) );
  AND U2783 ( .A(n185), .B(n3431), .Z(n3430) );
  XOR U2784 ( .A(p_input[8125]), .B(p_input[8093]), .Z(n3431) );
  XOR U2785 ( .A(n3432), .B(n3433), .Z(n3423) );
  AND U2786 ( .A(n3434), .B(n3435), .Z(n3433) );
  XOR U2787 ( .A(n3432), .B(n3075), .Z(n3435) );
  XNOR U2788 ( .A(p_input[8156]), .B(n3436), .Z(n3075) );
  AND U2789 ( .A(n187), .B(n3437), .Z(n3436) );
  XOR U2790 ( .A(p_input[8188]), .B(p_input[8156]), .Z(n3437) );
  XNOR U2791 ( .A(n3072), .B(n3432), .Z(n3434) );
  XOR U2792 ( .A(n3438), .B(n3439), .Z(n3072) );
  AND U2793 ( .A(n185), .B(n3440), .Z(n3439) );
  XOR U2794 ( .A(p_input[8124]), .B(p_input[8092]), .Z(n3440) );
  XOR U2795 ( .A(n3441), .B(n3442), .Z(n3432) );
  AND U2796 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U2797 ( .A(n3441), .B(n3087), .Z(n3444) );
  XNOR U2798 ( .A(p_input[8155]), .B(n3445), .Z(n3087) );
  AND U2799 ( .A(n187), .B(n3446), .Z(n3445) );
  XOR U2800 ( .A(p_input[8187]), .B(p_input[8155]), .Z(n3446) );
  XNOR U2801 ( .A(n3084), .B(n3441), .Z(n3443) );
  XOR U2802 ( .A(n3447), .B(n3448), .Z(n3084) );
  AND U2803 ( .A(n185), .B(n3449), .Z(n3448) );
  XOR U2804 ( .A(p_input[8123]), .B(p_input[8091]), .Z(n3449) );
  XOR U2805 ( .A(n3450), .B(n3451), .Z(n3441) );
  AND U2806 ( .A(n3452), .B(n3453), .Z(n3451) );
  XOR U2807 ( .A(n3450), .B(n3099), .Z(n3453) );
  XNOR U2808 ( .A(p_input[8154]), .B(n3454), .Z(n3099) );
  AND U2809 ( .A(n187), .B(n3455), .Z(n3454) );
  XOR U2810 ( .A(p_input[8186]), .B(p_input[8154]), .Z(n3455) );
  XNOR U2811 ( .A(n3096), .B(n3450), .Z(n3452) );
  XOR U2812 ( .A(n3456), .B(n3457), .Z(n3096) );
  AND U2813 ( .A(n185), .B(n3458), .Z(n3457) );
  XOR U2814 ( .A(p_input[8122]), .B(p_input[8090]), .Z(n3458) );
  XOR U2815 ( .A(n3459), .B(n3460), .Z(n3450) );
  AND U2816 ( .A(n3461), .B(n3462), .Z(n3460) );
  XOR U2817 ( .A(n3459), .B(n3111), .Z(n3462) );
  XNOR U2818 ( .A(p_input[8153]), .B(n3463), .Z(n3111) );
  AND U2819 ( .A(n187), .B(n3464), .Z(n3463) );
  XOR U2820 ( .A(p_input[8185]), .B(p_input[8153]), .Z(n3464) );
  XNOR U2821 ( .A(n3108), .B(n3459), .Z(n3461) );
  XOR U2822 ( .A(n3465), .B(n3466), .Z(n3108) );
  AND U2823 ( .A(n185), .B(n3467), .Z(n3466) );
  XOR U2824 ( .A(p_input[8121]), .B(p_input[8089]), .Z(n3467) );
  XOR U2825 ( .A(n3468), .B(n3469), .Z(n3459) );
  AND U2826 ( .A(n3470), .B(n3471), .Z(n3469) );
  XOR U2827 ( .A(n3468), .B(n3123), .Z(n3471) );
  XNOR U2828 ( .A(p_input[8152]), .B(n3472), .Z(n3123) );
  AND U2829 ( .A(n187), .B(n3473), .Z(n3472) );
  XOR U2830 ( .A(p_input[8184]), .B(p_input[8152]), .Z(n3473) );
  XNOR U2831 ( .A(n3120), .B(n3468), .Z(n3470) );
  XOR U2832 ( .A(n3474), .B(n3475), .Z(n3120) );
  AND U2833 ( .A(n185), .B(n3476), .Z(n3475) );
  XOR U2834 ( .A(p_input[8120]), .B(p_input[8088]), .Z(n3476) );
  XOR U2835 ( .A(n3477), .B(n3478), .Z(n3468) );
  AND U2836 ( .A(n3479), .B(n3480), .Z(n3478) );
  XOR U2837 ( .A(n3477), .B(n3135), .Z(n3480) );
  XNOR U2838 ( .A(p_input[8151]), .B(n3481), .Z(n3135) );
  AND U2839 ( .A(n187), .B(n3482), .Z(n3481) );
  XOR U2840 ( .A(p_input[8183]), .B(p_input[8151]), .Z(n3482) );
  XNOR U2841 ( .A(n3132), .B(n3477), .Z(n3479) );
  XOR U2842 ( .A(n3483), .B(n3484), .Z(n3132) );
  AND U2843 ( .A(n185), .B(n3485), .Z(n3484) );
  XOR U2844 ( .A(p_input[8119]), .B(p_input[8087]), .Z(n3485) );
  XOR U2845 ( .A(n3486), .B(n3487), .Z(n3477) );
  AND U2846 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR U2847 ( .A(n3486), .B(n3147), .Z(n3489) );
  XNOR U2848 ( .A(p_input[8150]), .B(n3490), .Z(n3147) );
  AND U2849 ( .A(n187), .B(n3491), .Z(n3490) );
  XOR U2850 ( .A(p_input[8182]), .B(p_input[8150]), .Z(n3491) );
  XNOR U2851 ( .A(n3144), .B(n3486), .Z(n3488) );
  XOR U2852 ( .A(n3492), .B(n3493), .Z(n3144) );
  AND U2853 ( .A(n185), .B(n3494), .Z(n3493) );
  XOR U2854 ( .A(p_input[8118]), .B(p_input[8086]), .Z(n3494) );
  XOR U2855 ( .A(n3495), .B(n3496), .Z(n3486) );
  AND U2856 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR U2857 ( .A(n3495), .B(n3159), .Z(n3498) );
  XNOR U2858 ( .A(p_input[8149]), .B(n3499), .Z(n3159) );
  AND U2859 ( .A(n187), .B(n3500), .Z(n3499) );
  XOR U2860 ( .A(p_input[8181]), .B(p_input[8149]), .Z(n3500) );
  XNOR U2861 ( .A(n3156), .B(n3495), .Z(n3497) );
  XOR U2862 ( .A(n3501), .B(n3502), .Z(n3156) );
  AND U2863 ( .A(n185), .B(n3503), .Z(n3502) );
  XOR U2864 ( .A(p_input[8117]), .B(p_input[8085]), .Z(n3503) );
  XOR U2865 ( .A(n3504), .B(n3505), .Z(n3495) );
  AND U2866 ( .A(n3506), .B(n3507), .Z(n3505) );
  XOR U2867 ( .A(n3504), .B(n3171), .Z(n3507) );
  XNOR U2868 ( .A(p_input[8148]), .B(n3508), .Z(n3171) );
  AND U2869 ( .A(n187), .B(n3509), .Z(n3508) );
  XOR U2870 ( .A(p_input[8180]), .B(p_input[8148]), .Z(n3509) );
  XNOR U2871 ( .A(n3168), .B(n3504), .Z(n3506) );
  XOR U2872 ( .A(n3510), .B(n3511), .Z(n3168) );
  AND U2873 ( .A(n185), .B(n3512), .Z(n3511) );
  XOR U2874 ( .A(p_input[8116]), .B(p_input[8084]), .Z(n3512) );
  XOR U2875 ( .A(n3513), .B(n3514), .Z(n3504) );
  AND U2876 ( .A(n3515), .B(n3516), .Z(n3514) );
  XOR U2877 ( .A(n3513), .B(n3183), .Z(n3516) );
  XNOR U2878 ( .A(p_input[8147]), .B(n3517), .Z(n3183) );
  AND U2879 ( .A(n187), .B(n3518), .Z(n3517) );
  XOR U2880 ( .A(p_input[8179]), .B(p_input[8147]), .Z(n3518) );
  XNOR U2881 ( .A(n3180), .B(n3513), .Z(n3515) );
  XOR U2882 ( .A(n3519), .B(n3520), .Z(n3180) );
  AND U2883 ( .A(n185), .B(n3521), .Z(n3520) );
  XOR U2884 ( .A(p_input[8115]), .B(p_input[8083]), .Z(n3521) );
  XOR U2885 ( .A(n3522), .B(n3523), .Z(n3513) );
  AND U2886 ( .A(n3524), .B(n3525), .Z(n3523) );
  XOR U2887 ( .A(n3522), .B(n3195), .Z(n3525) );
  XNOR U2888 ( .A(p_input[8146]), .B(n3526), .Z(n3195) );
  AND U2889 ( .A(n187), .B(n3527), .Z(n3526) );
  XOR U2890 ( .A(p_input[8178]), .B(p_input[8146]), .Z(n3527) );
  XNOR U2891 ( .A(n3192), .B(n3522), .Z(n3524) );
  XOR U2892 ( .A(n3528), .B(n3529), .Z(n3192) );
  AND U2893 ( .A(n185), .B(n3530), .Z(n3529) );
  XOR U2894 ( .A(p_input[8114]), .B(p_input[8082]), .Z(n3530) );
  XOR U2895 ( .A(n3531), .B(n3532), .Z(n3522) );
  AND U2896 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR U2897 ( .A(n3531), .B(n3207), .Z(n3534) );
  XNOR U2898 ( .A(p_input[8145]), .B(n3535), .Z(n3207) );
  AND U2899 ( .A(n187), .B(n3536), .Z(n3535) );
  XOR U2900 ( .A(p_input[8177]), .B(p_input[8145]), .Z(n3536) );
  XNOR U2901 ( .A(n3204), .B(n3531), .Z(n3533) );
  XOR U2902 ( .A(n3537), .B(n3538), .Z(n3204) );
  AND U2903 ( .A(n185), .B(n3539), .Z(n3538) );
  XOR U2904 ( .A(p_input[8113]), .B(p_input[8081]), .Z(n3539) );
  XOR U2905 ( .A(n3540), .B(n3541), .Z(n3531) );
  AND U2906 ( .A(n3542), .B(n3543), .Z(n3541) );
  XOR U2907 ( .A(n3540), .B(n3219), .Z(n3543) );
  XNOR U2908 ( .A(p_input[8144]), .B(n3544), .Z(n3219) );
  AND U2909 ( .A(n187), .B(n3545), .Z(n3544) );
  XOR U2910 ( .A(p_input[8176]), .B(p_input[8144]), .Z(n3545) );
  XNOR U2911 ( .A(n3216), .B(n3540), .Z(n3542) );
  XOR U2912 ( .A(n3546), .B(n3547), .Z(n3216) );
  AND U2913 ( .A(n185), .B(n3548), .Z(n3547) );
  XOR U2914 ( .A(p_input[8112]), .B(p_input[8080]), .Z(n3548) );
  XOR U2915 ( .A(n3549), .B(n3550), .Z(n3540) );
  AND U2916 ( .A(n3551), .B(n3552), .Z(n3550) );
  XOR U2917 ( .A(n3549), .B(n3231), .Z(n3552) );
  XNOR U2918 ( .A(p_input[8143]), .B(n3553), .Z(n3231) );
  AND U2919 ( .A(n187), .B(n3554), .Z(n3553) );
  XOR U2920 ( .A(p_input[8175]), .B(p_input[8143]), .Z(n3554) );
  XNOR U2921 ( .A(n3228), .B(n3549), .Z(n3551) );
  XOR U2922 ( .A(n3555), .B(n3556), .Z(n3228) );
  AND U2923 ( .A(n185), .B(n3557), .Z(n3556) );
  XOR U2924 ( .A(p_input[8111]), .B(p_input[8079]), .Z(n3557) );
  XOR U2925 ( .A(n3558), .B(n3559), .Z(n3549) );
  AND U2926 ( .A(n3560), .B(n3561), .Z(n3559) );
  XOR U2927 ( .A(n3558), .B(n3243), .Z(n3561) );
  XNOR U2928 ( .A(p_input[8142]), .B(n3562), .Z(n3243) );
  AND U2929 ( .A(n187), .B(n3563), .Z(n3562) );
  XOR U2930 ( .A(p_input[8174]), .B(p_input[8142]), .Z(n3563) );
  XNOR U2931 ( .A(n3240), .B(n3558), .Z(n3560) );
  XOR U2932 ( .A(n3564), .B(n3565), .Z(n3240) );
  AND U2933 ( .A(n185), .B(n3566), .Z(n3565) );
  XOR U2934 ( .A(p_input[8110]), .B(p_input[8078]), .Z(n3566) );
  XOR U2935 ( .A(n3567), .B(n3568), .Z(n3558) );
  AND U2936 ( .A(n3569), .B(n3570), .Z(n3568) );
  XOR U2937 ( .A(n3567), .B(n3255), .Z(n3570) );
  XNOR U2938 ( .A(p_input[8141]), .B(n3571), .Z(n3255) );
  AND U2939 ( .A(n187), .B(n3572), .Z(n3571) );
  XOR U2940 ( .A(p_input[8173]), .B(p_input[8141]), .Z(n3572) );
  XNOR U2941 ( .A(n3252), .B(n3567), .Z(n3569) );
  XOR U2942 ( .A(n3573), .B(n3574), .Z(n3252) );
  AND U2943 ( .A(n185), .B(n3575), .Z(n3574) );
  XOR U2944 ( .A(p_input[8109]), .B(p_input[8077]), .Z(n3575) );
  XOR U2945 ( .A(n3576), .B(n3577), .Z(n3567) );
  AND U2946 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U2947 ( .A(n3576), .B(n3267), .Z(n3579) );
  XNOR U2948 ( .A(p_input[8140]), .B(n3580), .Z(n3267) );
  AND U2949 ( .A(n187), .B(n3581), .Z(n3580) );
  XOR U2950 ( .A(p_input[8172]), .B(p_input[8140]), .Z(n3581) );
  XNOR U2951 ( .A(n3264), .B(n3576), .Z(n3578) );
  XOR U2952 ( .A(n3582), .B(n3583), .Z(n3264) );
  AND U2953 ( .A(n185), .B(n3584), .Z(n3583) );
  XOR U2954 ( .A(p_input[8108]), .B(p_input[8076]), .Z(n3584) );
  XOR U2955 ( .A(n3585), .B(n3586), .Z(n3576) );
  AND U2956 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR U2957 ( .A(n3585), .B(n3279), .Z(n3588) );
  XNOR U2958 ( .A(p_input[8139]), .B(n3589), .Z(n3279) );
  AND U2959 ( .A(n187), .B(n3590), .Z(n3589) );
  XOR U2960 ( .A(p_input[8171]), .B(p_input[8139]), .Z(n3590) );
  XNOR U2961 ( .A(n3276), .B(n3585), .Z(n3587) );
  XOR U2962 ( .A(n3591), .B(n3592), .Z(n3276) );
  AND U2963 ( .A(n185), .B(n3593), .Z(n3592) );
  XOR U2964 ( .A(p_input[8107]), .B(p_input[8075]), .Z(n3593) );
  XOR U2965 ( .A(n3594), .B(n3595), .Z(n3585) );
  AND U2966 ( .A(n3596), .B(n3597), .Z(n3595) );
  XOR U2967 ( .A(n3594), .B(n3291), .Z(n3597) );
  XNOR U2968 ( .A(p_input[8138]), .B(n3598), .Z(n3291) );
  AND U2969 ( .A(n187), .B(n3599), .Z(n3598) );
  XOR U2970 ( .A(p_input[8170]), .B(p_input[8138]), .Z(n3599) );
  XNOR U2971 ( .A(n3288), .B(n3594), .Z(n3596) );
  XOR U2972 ( .A(n3600), .B(n3601), .Z(n3288) );
  AND U2973 ( .A(n185), .B(n3602), .Z(n3601) );
  XOR U2974 ( .A(p_input[8106]), .B(p_input[8074]), .Z(n3602) );
  XOR U2975 ( .A(n3603), .B(n3604), .Z(n3594) );
  AND U2976 ( .A(n3605), .B(n3606), .Z(n3604) );
  XOR U2977 ( .A(n3603), .B(n3303), .Z(n3606) );
  XNOR U2978 ( .A(p_input[8137]), .B(n3607), .Z(n3303) );
  AND U2979 ( .A(n187), .B(n3608), .Z(n3607) );
  XOR U2980 ( .A(p_input[8169]), .B(p_input[8137]), .Z(n3608) );
  XNOR U2981 ( .A(n3300), .B(n3603), .Z(n3605) );
  XOR U2982 ( .A(n3609), .B(n3610), .Z(n3300) );
  AND U2983 ( .A(n185), .B(n3611), .Z(n3610) );
  XOR U2984 ( .A(p_input[8105]), .B(p_input[8073]), .Z(n3611) );
  XOR U2985 ( .A(n3612), .B(n3613), .Z(n3603) );
  AND U2986 ( .A(n3614), .B(n3615), .Z(n3613) );
  XOR U2987 ( .A(n3612), .B(n3315), .Z(n3615) );
  XNOR U2988 ( .A(p_input[8136]), .B(n3616), .Z(n3315) );
  AND U2989 ( .A(n187), .B(n3617), .Z(n3616) );
  XOR U2990 ( .A(p_input[8168]), .B(p_input[8136]), .Z(n3617) );
  XNOR U2991 ( .A(n3312), .B(n3612), .Z(n3614) );
  XOR U2992 ( .A(n3618), .B(n3619), .Z(n3312) );
  AND U2993 ( .A(n185), .B(n3620), .Z(n3619) );
  XOR U2994 ( .A(p_input[8104]), .B(p_input[8072]), .Z(n3620) );
  XOR U2995 ( .A(n3621), .B(n3622), .Z(n3612) );
  AND U2996 ( .A(n3623), .B(n3624), .Z(n3622) );
  XOR U2997 ( .A(n3621), .B(n3327), .Z(n3624) );
  XNOR U2998 ( .A(p_input[8135]), .B(n3625), .Z(n3327) );
  AND U2999 ( .A(n187), .B(n3626), .Z(n3625) );
  XOR U3000 ( .A(p_input[8167]), .B(p_input[8135]), .Z(n3626) );
  XNOR U3001 ( .A(n3324), .B(n3621), .Z(n3623) );
  XOR U3002 ( .A(n3627), .B(n3628), .Z(n3324) );
  AND U3003 ( .A(n185), .B(n3629), .Z(n3628) );
  XOR U3004 ( .A(p_input[8103]), .B(p_input[8071]), .Z(n3629) );
  XOR U3005 ( .A(n3630), .B(n3631), .Z(n3621) );
  AND U3006 ( .A(n3632), .B(n3633), .Z(n3631) );
  XOR U3007 ( .A(n3630), .B(n3339), .Z(n3633) );
  XNOR U3008 ( .A(p_input[8134]), .B(n3634), .Z(n3339) );
  AND U3009 ( .A(n187), .B(n3635), .Z(n3634) );
  XOR U3010 ( .A(p_input[8166]), .B(p_input[8134]), .Z(n3635) );
  XNOR U3011 ( .A(n3336), .B(n3630), .Z(n3632) );
  XOR U3012 ( .A(n3636), .B(n3637), .Z(n3336) );
  AND U3013 ( .A(n185), .B(n3638), .Z(n3637) );
  XOR U3014 ( .A(p_input[8102]), .B(p_input[8070]), .Z(n3638) );
  XOR U3015 ( .A(n3639), .B(n3640), .Z(n3630) );
  AND U3016 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U3017 ( .A(n3639), .B(n3351), .Z(n3642) );
  XNOR U3018 ( .A(p_input[8133]), .B(n3643), .Z(n3351) );
  AND U3019 ( .A(n187), .B(n3644), .Z(n3643) );
  XOR U3020 ( .A(p_input[8165]), .B(p_input[8133]), .Z(n3644) );
  XNOR U3021 ( .A(n3348), .B(n3639), .Z(n3641) );
  XOR U3022 ( .A(n3645), .B(n3646), .Z(n3348) );
  AND U3023 ( .A(n185), .B(n3647), .Z(n3646) );
  XOR U3024 ( .A(p_input[8101]), .B(p_input[8069]), .Z(n3647) );
  XOR U3025 ( .A(n3648), .B(n3649), .Z(n3639) );
  AND U3026 ( .A(n3650), .B(n3651), .Z(n3649) );
  XOR U3027 ( .A(n3648), .B(n3363), .Z(n3651) );
  XNOR U3028 ( .A(p_input[8132]), .B(n3652), .Z(n3363) );
  AND U3029 ( .A(n187), .B(n3653), .Z(n3652) );
  XOR U3030 ( .A(p_input[8164]), .B(p_input[8132]), .Z(n3653) );
  XNOR U3031 ( .A(n3360), .B(n3648), .Z(n3650) );
  XOR U3032 ( .A(n3654), .B(n3655), .Z(n3360) );
  AND U3033 ( .A(n185), .B(n3656), .Z(n3655) );
  XOR U3034 ( .A(p_input[8100]), .B(p_input[8068]), .Z(n3656) );
  XOR U3035 ( .A(n3657), .B(n3658), .Z(n3648) );
  AND U3036 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U3037 ( .A(n3657), .B(n3375), .Z(n3660) );
  XNOR U3038 ( .A(p_input[8131]), .B(n3661), .Z(n3375) );
  AND U3039 ( .A(n187), .B(n3662), .Z(n3661) );
  XOR U3040 ( .A(p_input[8163]), .B(p_input[8131]), .Z(n3662) );
  XNOR U3041 ( .A(n3372), .B(n3657), .Z(n3659) );
  XOR U3042 ( .A(n3663), .B(n3664), .Z(n3372) );
  AND U3043 ( .A(n185), .B(n3665), .Z(n3664) );
  XOR U3044 ( .A(p_input[8099]), .B(p_input[8067]), .Z(n3665) );
  XOR U3045 ( .A(n3666), .B(n3667), .Z(n3657) );
  AND U3046 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U3047 ( .A(n3666), .B(n3387), .Z(n3669) );
  XNOR U3048 ( .A(p_input[8130]), .B(n3670), .Z(n3387) );
  AND U3049 ( .A(n187), .B(n3671), .Z(n3670) );
  XOR U3050 ( .A(p_input[8162]), .B(p_input[8130]), .Z(n3671) );
  XNOR U3051 ( .A(n3384), .B(n3666), .Z(n3668) );
  XOR U3052 ( .A(n3672), .B(n3673), .Z(n3384) );
  AND U3053 ( .A(n185), .B(n3674), .Z(n3673) );
  XOR U3054 ( .A(p_input[8098]), .B(p_input[8066]), .Z(n3674) );
  XOR U3055 ( .A(n3675), .B(n3676), .Z(n3666) );
  AND U3056 ( .A(n3677), .B(n3678), .Z(n3676) );
  XNOR U3057 ( .A(n3679), .B(n3400), .Z(n3678) );
  XNOR U3058 ( .A(p_input[8129]), .B(n3680), .Z(n3400) );
  AND U3059 ( .A(n187), .B(n3681), .Z(n3680) );
  XNOR U3060 ( .A(p_input[8161]), .B(n3682), .Z(n3681) );
  IV U3061 ( .A(p_input[8129]), .Z(n3682) );
  XNOR U3062 ( .A(n3397), .B(n3675), .Z(n3677) );
  XNOR U3063 ( .A(p_input[8065]), .B(n3683), .Z(n3397) );
  AND U3064 ( .A(n185), .B(n3684), .Z(n3683) );
  XOR U3065 ( .A(p_input[8097]), .B(p_input[8065]), .Z(n3684) );
  IV U3066 ( .A(n3679), .Z(n3675) );
  AND U3067 ( .A(n3405), .B(n3408), .Z(n3679) );
  XOR U3068 ( .A(p_input[8128]), .B(n3685), .Z(n3408) );
  AND U3069 ( .A(n187), .B(n3686), .Z(n3685) );
  XOR U3070 ( .A(p_input[8160]), .B(p_input[8128]), .Z(n3686) );
  XOR U3071 ( .A(n3687), .B(n3688), .Z(n187) );
  AND U3072 ( .A(n3689), .B(n3690), .Z(n3688) );
  XNOR U3073 ( .A(p_input[8191]), .B(n3687), .Z(n3690) );
  XOR U3074 ( .A(n3687), .B(p_input[8159]), .Z(n3689) );
  XOR U3075 ( .A(n3691), .B(n3692), .Z(n3687) );
  AND U3076 ( .A(n3693), .B(n3694), .Z(n3692) );
  XNOR U3077 ( .A(p_input[8190]), .B(n3691), .Z(n3694) );
  XOR U3078 ( .A(n3691), .B(p_input[8158]), .Z(n3693) );
  XOR U3079 ( .A(n3695), .B(n3696), .Z(n3691) );
  AND U3080 ( .A(n3697), .B(n3698), .Z(n3696) );
  XNOR U3081 ( .A(p_input[8189]), .B(n3695), .Z(n3698) );
  XOR U3082 ( .A(n3695), .B(p_input[8157]), .Z(n3697) );
  XOR U3083 ( .A(n3699), .B(n3700), .Z(n3695) );
  AND U3084 ( .A(n3701), .B(n3702), .Z(n3700) );
  XNOR U3085 ( .A(p_input[8188]), .B(n3699), .Z(n3702) );
  XOR U3086 ( .A(n3699), .B(p_input[8156]), .Z(n3701) );
  XOR U3087 ( .A(n3703), .B(n3704), .Z(n3699) );
  AND U3088 ( .A(n3705), .B(n3706), .Z(n3704) );
  XNOR U3089 ( .A(p_input[8187]), .B(n3703), .Z(n3706) );
  XOR U3090 ( .A(n3703), .B(p_input[8155]), .Z(n3705) );
  XOR U3091 ( .A(n3707), .B(n3708), .Z(n3703) );
  AND U3092 ( .A(n3709), .B(n3710), .Z(n3708) );
  XNOR U3093 ( .A(p_input[8186]), .B(n3707), .Z(n3710) );
  XOR U3094 ( .A(n3707), .B(p_input[8154]), .Z(n3709) );
  XOR U3095 ( .A(n3711), .B(n3712), .Z(n3707) );
  AND U3096 ( .A(n3713), .B(n3714), .Z(n3712) );
  XNOR U3097 ( .A(p_input[8185]), .B(n3711), .Z(n3714) );
  XOR U3098 ( .A(n3711), .B(p_input[8153]), .Z(n3713) );
  XOR U3099 ( .A(n3715), .B(n3716), .Z(n3711) );
  AND U3100 ( .A(n3717), .B(n3718), .Z(n3716) );
  XNOR U3101 ( .A(p_input[8184]), .B(n3715), .Z(n3718) );
  XOR U3102 ( .A(n3715), .B(p_input[8152]), .Z(n3717) );
  XOR U3103 ( .A(n3719), .B(n3720), .Z(n3715) );
  AND U3104 ( .A(n3721), .B(n3722), .Z(n3720) );
  XNOR U3105 ( .A(p_input[8183]), .B(n3719), .Z(n3722) );
  XOR U3106 ( .A(n3719), .B(p_input[8151]), .Z(n3721) );
  XOR U3107 ( .A(n3723), .B(n3724), .Z(n3719) );
  AND U3108 ( .A(n3725), .B(n3726), .Z(n3724) );
  XNOR U3109 ( .A(p_input[8182]), .B(n3723), .Z(n3726) );
  XOR U3110 ( .A(n3723), .B(p_input[8150]), .Z(n3725) );
  XOR U3111 ( .A(n3727), .B(n3728), .Z(n3723) );
  AND U3112 ( .A(n3729), .B(n3730), .Z(n3728) );
  XNOR U3113 ( .A(p_input[8181]), .B(n3727), .Z(n3730) );
  XOR U3114 ( .A(n3727), .B(p_input[8149]), .Z(n3729) );
  XOR U3115 ( .A(n3731), .B(n3732), .Z(n3727) );
  AND U3116 ( .A(n3733), .B(n3734), .Z(n3732) );
  XNOR U3117 ( .A(p_input[8180]), .B(n3731), .Z(n3734) );
  XOR U3118 ( .A(n3731), .B(p_input[8148]), .Z(n3733) );
  XOR U3119 ( .A(n3735), .B(n3736), .Z(n3731) );
  AND U3120 ( .A(n3737), .B(n3738), .Z(n3736) );
  XNOR U3121 ( .A(p_input[8179]), .B(n3735), .Z(n3738) );
  XOR U3122 ( .A(n3735), .B(p_input[8147]), .Z(n3737) );
  XOR U3123 ( .A(n3739), .B(n3740), .Z(n3735) );
  AND U3124 ( .A(n3741), .B(n3742), .Z(n3740) );
  XNOR U3125 ( .A(p_input[8178]), .B(n3739), .Z(n3742) );
  XOR U3126 ( .A(n3739), .B(p_input[8146]), .Z(n3741) );
  XOR U3127 ( .A(n3743), .B(n3744), .Z(n3739) );
  AND U3128 ( .A(n3745), .B(n3746), .Z(n3744) );
  XNOR U3129 ( .A(p_input[8177]), .B(n3743), .Z(n3746) );
  XOR U3130 ( .A(n3743), .B(p_input[8145]), .Z(n3745) );
  XOR U3131 ( .A(n3747), .B(n3748), .Z(n3743) );
  AND U3132 ( .A(n3749), .B(n3750), .Z(n3748) );
  XNOR U3133 ( .A(p_input[8176]), .B(n3747), .Z(n3750) );
  XOR U3134 ( .A(n3747), .B(p_input[8144]), .Z(n3749) );
  XOR U3135 ( .A(n3751), .B(n3752), .Z(n3747) );
  AND U3136 ( .A(n3753), .B(n3754), .Z(n3752) );
  XNOR U3137 ( .A(p_input[8175]), .B(n3751), .Z(n3754) );
  XOR U3138 ( .A(n3751), .B(p_input[8143]), .Z(n3753) );
  XOR U3139 ( .A(n3755), .B(n3756), .Z(n3751) );
  AND U3140 ( .A(n3757), .B(n3758), .Z(n3756) );
  XNOR U3141 ( .A(p_input[8174]), .B(n3755), .Z(n3758) );
  XOR U3142 ( .A(n3755), .B(p_input[8142]), .Z(n3757) );
  XOR U3143 ( .A(n3759), .B(n3760), .Z(n3755) );
  AND U3144 ( .A(n3761), .B(n3762), .Z(n3760) );
  XNOR U3145 ( .A(p_input[8173]), .B(n3759), .Z(n3762) );
  XOR U3146 ( .A(n3759), .B(p_input[8141]), .Z(n3761) );
  XOR U3147 ( .A(n3763), .B(n3764), .Z(n3759) );
  AND U3148 ( .A(n3765), .B(n3766), .Z(n3764) );
  XNOR U3149 ( .A(p_input[8172]), .B(n3763), .Z(n3766) );
  XOR U3150 ( .A(n3763), .B(p_input[8140]), .Z(n3765) );
  XOR U3151 ( .A(n3767), .B(n3768), .Z(n3763) );
  AND U3152 ( .A(n3769), .B(n3770), .Z(n3768) );
  XNOR U3153 ( .A(p_input[8171]), .B(n3767), .Z(n3770) );
  XOR U3154 ( .A(n3767), .B(p_input[8139]), .Z(n3769) );
  XOR U3155 ( .A(n3771), .B(n3772), .Z(n3767) );
  AND U3156 ( .A(n3773), .B(n3774), .Z(n3772) );
  XNOR U3157 ( .A(p_input[8170]), .B(n3771), .Z(n3774) );
  XOR U3158 ( .A(n3771), .B(p_input[8138]), .Z(n3773) );
  XOR U3159 ( .A(n3775), .B(n3776), .Z(n3771) );
  AND U3160 ( .A(n3777), .B(n3778), .Z(n3776) );
  XNOR U3161 ( .A(p_input[8169]), .B(n3775), .Z(n3778) );
  XOR U3162 ( .A(n3775), .B(p_input[8137]), .Z(n3777) );
  XOR U3163 ( .A(n3779), .B(n3780), .Z(n3775) );
  AND U3164 ( .A(n3781), .B(n3782), .Z(n3780) );
  XNOR U3165 ( .A(p_input[8168]), .B(n3779), .Z(n3782) );
  XOR U3166 ( .A(n3779), .B(p_input[8136]), .Z(n3781) );
  XOR U3167 ( .A(n3783), .B(n3784), .Z(n3779) );
  AND U3168 ( .A(n3785), .B(n3786), .Z(n3784) );
  XNOR U3169 ( .A(p_input[8167]), .B(n3783), .Z(n3786) );
  XOR U3170 ( .A(n3783), .B(p_input[8135]), .Z(n3785) );
  XOR U3171 ( .A(n3787), .B(n3788), .Z(n3783) );
  AND U3172 ( .A(n3789), .B(n3790), .Z(n3788) );
  XNOR U3173 ( .A(p_input[8166]), .B(n3787), .Z(n3790) );
  XOR U3174 ( .A(n3787), .B(p_input[8134]), .Z(n3789) );
  XOR U3175 ( .A(n3791), .B(n3792), .Z(n3787) );
  AND U3176 ( .A(n3793), .B(n3794), .Z(n3792) );
  XNOR U3177 ( .A(p_input[8165]), .B(n3791), .Z(n3794) );
  XOR U3178 ( .A(n3791), .B(p_input[8133]), .Z(n3793) );
  XOR U3179 ( .A(n3795), .B(n3796), .Z(n3791) );
  AND U3180 ( .A(n3797), .B(n3798), .Z(n3796) );
  XNOR U3181 ( .A(p_input[8164]), .B(n3795), .Z(n3798) );
  XOR U3182 ( .A(n3795), .B(p_input[8132]), .Z(n3797) );
  XOR U3183 ( .A(n3799), .B(n3800), .Z(n3795) );
  AND U3184 ( .A(n3801), .B(n3802), .Z(n3800) );
  XNOR U3185 ( .A(p_input[8163]), .B(n3799), .Z(n3802) );
  XOR U3186 ( .A(n3799), .B(p_input[8131]), .Z(n3801) );
  XOR U3187 ( .A(n3803), .B(n3804), .Z(n3799) );
  AND U3188 ( .A(n3805), .B(n3806), .Z(n3804) );
  XNOR U3189 ( .A(p_input[8162]), .B(n3803), .Z(n3806) );
  XOR U3190 ( .A(n3803), .B(p_input[8130]), .Z(n3805) );
  XNOR U3191 ( .A(n3807), .B(n3808), .Z(n3803) );
  AND U3192 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U3193 ( .A(p_input[8161]), .B(n3807), .Z(n3810) );
  XNOR U3194 ( .A(p_input[8129]), .B(n3807), .Z(n3809) );
  AND U3195 ( .A(p_input[8160]), .B(n3811), .Z(n3807) );
  IV U3196 ( .A(p_input[8128]), .Z(n3811) );
  XNOR U3197 ( .A(p_input[8064]), .B(n3812), .Z(n3405) );
  AND U3198 ( .A(n185), .B(n3813), .Z(n3812) );
  XOR U3199 ( .A(p_input[8096]), .B(p_input[8064]), .Z(n3813) );
  XOR U3200 ( .A(n3814), .B(n3815), .Z(n185) );
  AND U3201 ( .A(n3816), .B(n3817), .Z(n3815) );
  XNOR U3202 ( .A(p_input[8127]), .B(n3814), .Z(n3817) );
  XOR U3203 ( .A(n3814), .B(p_input[8095]), .Z(n3816) );
  XOR U3204 ( .A(n3818), .B(n3819), .Z(n3814) );
  AND U3205 ( .A(n3820), .B(n3821), .Z(n3819) );
  XNOR U3206 ( .A(p_input[8126]), .B(n3818), .Z(n3821) );
  XNOR U3207 ( .A(n3818), .B(n3420), .Z(n3820) );
  IV U3208 ( .A(p_input[8094]), .Z(n3420) );
  XOR U3209 ( .A(n3822), .B(n3823), .Z(n3818) );
  AND U3210 ( .A(n3824), .B(n3825), .Z(n3823) );
  XNOR U3211 ( .A(p_input[8125]), .B(n3822), .Z(n3825) );
  XNOR U3212 ( .A(n3822), .B(n3429), .Z(n3824) );
  IV U3213 ( .A(p_input[8093]), .Z(n3429) );
  XOR U3214 ( .A(n3826), .B(n3827), .Z(n3822) );
  AND U3215 ( .A(n3828), .B(n3829), .Z(n3827) );
  XNOR U3216 ( .A(p_input[8124]), .B(n3826), .Z(n3829) );
  XNOR U3217 ( .A(n3826), .B(n3438), .Z(n3828) );
  IV U3218 ( .A(p_input[8092]), .Z(n3438) );
  XOR U3219 ( .A(n3830), .B(n3831), .Z(n3826) );
  AND U3220 ( .A(n3832), .B(n3833), .Z(n3831) );
  XNOR U3221 ( .A(p_input[8123]), .B(n3830), .Z(n3833) );
  XNOR U3222 ( .A(n3830), .B(n3447), .Z(n3832) );
  IV U3223 ( .A(p_input[8091]), .Z(n3447) );
  XOR U3224 ( .A(n3834), .B(n3835), .Z(n3830) );
  AND U3225 ( .A(n3836), .B(n3837), .Z(n3835) );
  XNOR U3226 ( .A(p_input[8122]), .B(n3834), .Z(n3837) );
  XNOR U3227 ( .A(n3834), .B(n3456), .Z(n3836) );
  IV U3228 ( .A(p_input[8090]), .Z(n3456) );
  XOR U3229 ( .A(n3838), .B(n3839), .Z(n3834) );
  AND U3230 ( .A(n3840), .B(n3841), .Z(n3839) );
  XNOR U3231 ( .A(p_input[8121]), .B(n3838), .Z(n3841) );
  XNOR U3232 ( .A(n3838), .B(n3465), .Z(n3840) );
  IV U3233 ( .A(p_input[8089]), .Z(n3465) );
  XOR U3234 ( .A(n3842), .B(n3843), .Z(n3838) );
  AND U3235 ( .A(n3844), .B(n3845), .Z(n3843) );
  XNOR U3236 ( .A(p_input[8120]), .B(n3842), .Z(n3845) );
  XNOR U3237 ( .A(n3842), .B(n3474), .Z(n3844) );
  IV U3238 ( .A(p_input[8088]), .Z(n3474) );
  XOR U3239 ( .A(n3846), .B(n3847), .Z(n3842) );
  AND U3240 ( .A(n3848), .B(n3849), .Z(n3847) );
  XNOR U3241 ( .A(p_input[8119]), .B(n3846), .Z(n3849) );
  XNOR U3242 ( .A(n3846), .B(n3483), .Z(n3848) );
  IV U3243 ( .A(p_input[8087]), .Z(n3483) );
  XOR U3244 ( .A(n3850), .B(n3851), .Z(n3846) );
  AND U3245 ( .A(n3852), .B(n3853), .Z(n3851) );
  XNOR U3246 ( .A(p_input[8118]), .B(n3850), .Z(n3853) );
  XNOR U3247 ( .A(n3850), .B(n3492), .Z(n3852) );
  IV U3248 ( .A(p_input[8086]), .Z(n3492) );
  XOR U3249 ( .A(n3854), .B(n3855), .Z(n3850) );
  AND U3250 ( .A(n3856), .B(n3857), .Z(n3855) );
  XNOR U3251 ( .A(p_input[8117]), .B(n3854), .Z(n3857) );
  XNOR U3252 ( .A(n3854), .B(n3501), .Z(n3856) );
  IV U3253 ( .A(p_input[8085]), .Z(n3501) );
  XOR U3254 ( .A(n3858), .B(n3859), .Z(n3854) );
  AND U3255 ( .A(n3860), .B(n3861), .Z(n3859) );
  XNOR U3256 ( .A(p_input[8116]), .B(n3858), .Z(n3861) );
  XNOR U3257 ( .A(n3858), .B(n3510), .Z(n3860) );
  IV U3258 ( .A(p_input[8084]), .Z(n3510) );
  XOR U3259 ( .A(n3862), .B(n3863), .Z(n3858) );
  AND U3260 ( .A(n3864), .B(n3865), .Z(n3863) );
  XNOR U3261 ( .A(p_input[8115]), .B(n3862), .Z(n3865) );
  XNOR U3262 ( .A(n3862), .B(n3519), .Z(n3864) );
  IV U3263 ( .A(p_input[8083]), .Z(n3519) );
  XOR U3264 ( .A(n3866), .B(n3867), .Z(n3862) );
  AND U3265 ( .A(n3868), .B(n3869), .Z(n3867) );
  XNOR U3266 ( .A(p_input[8114]), .B(n3866), .Z(n3869) );
  XNOR U3267 ( .A(n3866), .B(n3528), .Z(n3868) );
  IV U3268 ( .A(p_input[8082]), .Z(n3528) );
  XOR U3269 ( .A(n3870), .B(n3871), .Z(n3866) );
  AND U3270 ( .A(n3872), .B(n3873), .Z(n3871) );
  XNOR U3271 ( .A(p_input[8113]), .B(n3870), .Z(n3873) );
  XNOR U3272 ( .A(n3870), .B(n3537), .Z(n3872) );
  IV U3273 ( .A(p_input[8081]), .Z(n3537) );
  XOR U3274 ( .A(n3874), .B(n3875), .Z(n3870) );
  AND U3275 ( .A(n3876), .B(n3877), .Z(n3875) );
  XNOR U3276 ( .A(p_input[8112]), .B(n3874), .Z(n3877) );
  XNOR U3277 ( .A(n3874), .B(n3546), .Z(n3876) );
  IV U3278 ( .A(p_input[8080]), .Z(n3546) );
  XOR U3279 ( .A(n3878), .B(n3879), .Z(n3874) );
  AND U3280 ( .A(n3880), .B(n3881), .Z(n3879) );
  XNOR U3281 ( .A(p_input[8111]), .B(n3878), .Z(n3881) );
  XNOR U3282 ( .A(n3878), .B(n3555), .Z(n3880) );
  IV U3283 ( .A(p_input[8079]), .Z(n3555) );
  XOR U3284 ( .A(n3882), .B(n3883), .Z(n3878) );
  AND U3285 ( .A(n3884), .B(n3885), .Z(n3883) );
  XNOR U3286 ( .A(p_input[8110]), .B(n3882), .Z(n3885) );
  XNOR U3287 ( .A(n3882), .B(n3564), .Z(n3884) );
  IV U3288 ( .A(p_input[8078]), .Z(n3564) );
  XOR U3289 ( .A(n3886), .B(n3887), .Z(n3882) );
  AND U3290 ( .A(n3888), .B(n3889), .Z(n3887) );
  XNOR U3291 ( .A(p_input[8109]), .B(n3886), .Z(n3889) );
  XNOR U3292 ( .A(n3886), .B(n3573), .Z(n3888) );
  IV U3293 ( .A(p_input[8077]), .Z(n3573) );
  XOR U3294 ( .A(n3890), .B(n3891), .Z(n3886) );
  AND U3295 ( .A(n3892), .B(n3893), .Z(n3891) );
  XNOR U3296 ( .A(p_input[8108]), .B(n3890), .Z(n3893) );
  XNOR U3297 ( .A(n3890), .B(n3582), .Z(n3892) );
  IV U3298 ( .A(p_input[8076]), .Z(n3582) );
  XOR U3299 ( .A(n3894), .B(n3895), .Z(n3890) );
  AND U3300 ( .A(n3896), .B(n3897), .Z(n3895) );
  XNOR U3301 ( .A(p_input[8107]), .B(n3894), .Z(n3897) );
  XNOR U3302 ( .A(n3894), .B(n3591), .Z(n3896) );
  IV U3303 ( .A(p_input[8075]), .Z(n3591) );
  XOR U3304 ( .A(n3898), .B(n3899), .Z(n3894) );
  AND U3305 ( .A(n3900), .B(n3901), .Z(n3899) );
  XNOR U3306 ( .A(p_input[8106]), .B(n3898), .Z(n3901) );
  XNOR U3307 ( .A(n3898), .B(n3600), .Z(n3900) );
  IV U3308 ( .A(p_input[8074]), .Z(n3600) );
  XOR U3309 ( .A(n3902), .B(n3903), .Z(n3898) );
  AND U3310 ( .A(n3904), .B(n3905), .Z(n3903) );
  XNOR U3311 ( .A(p_input[8105]), .B(n3902), .Z(n3905) );
  XNOR U3312 ( .A(n3902), .B(n3609), .Z(n3904) );
  IV U3313 ( .A(p_input[8073]), .Z(n3609) );
  XOR U3314 ( .A(n3906), .B(n3907), .Z(n3902) );
  AND U3315 ( .A(n3908), .B(n3909), .Z(n3907) );
  XNOR U3316 ( .A(p_input[8104]), .B(n3906), .Z(n3909) );
  XNOR U3317 ( .A(n3906), .B(n3618), .Z(n3908) );
  IV U3318 ( .A(p_input[8072]), .Z(n3618) );
  XOR U3319 ( .A(n3910), .B(n3911), .Z(n3906) );
  AND U3320 ( .A(n3912), .B(n3913), .Z(n3911) );
  XNOR U3321 ( .A(p_input[8103]), .B(n3910), .Z(n3913) );
  XNOR U3322 ( .A(n3910), .B(n3627), .Z(n3912) );
  IV U3323 ( .A(p_input[8071]), .Z(n3627) );
  XOR U3324 ( .A(n3914), .B(n3915), .Z(n3910) );
  AND U3325 ( .A(n3916), .B(n3917), .Z(n3915) );
  XNOR U3326 ( .A(p_input[8102]), .B(n3914), .Z(n3917) );
  XNOR U3327 ( .A(n3914), .B(n3636), .Z(n3916) );
  IV U3328 ( .A(p_input[8070]), .Z(n3636) );
  XOR U3329 ( .A(n3918), .B(n3919), .Z(n3914) );
  AND U3330 ( .A(n3920), .B(n3921), .Z(n3919) );
  XNOR U3331 ( .A(p_input[8101]), .B(n3918), .Z(n3921) );
  XNOR U3332 ( .A(n3918), .B(n3645), .Z(n3920) );
  IV U3333 ( .A(p_input[8069]), .Z(n3645) );
  XOR U3334 ( .A(n3922), .B(n3923), .Z(n3918) );
  AND U3335 ( .A(n3924), .B(n3925), .Z(n3923) );
  XNOR U3336 ( .A(p_input[8100]), .B(n3922), .Z(n3925) );
  XNOR U3337 ( .A(n3922), .B(n3654), .Z(n3924) );
  IV U3338 ( .A(p_input[8068]), .Z(n3654) );
  XOR U3339 ( .A(n3926), .B(n3927), .Z(n3922) );
  AND U3340 ( .A(n3928), .B(n3929), .Z(n3927) );
  XNOR U3341 ( .A(p_input[8099]), .B(n3926), .Z(n3929) );
  XNOR U3342 ( .A(n3926), .B(n3663), .Z(n3928) );
  IV U3343 ( .A(p_input[8067]), .Z(n3663) );
  XOR U3344 ( .A(n3930), .B(n3931), .Z(n3926) );
  AND U3345 ( .A(n3932), .B(n3933), .Z(n3931) );
  XNOR U3346 ( .A(p_input[8098]), .B(n3930), .Z(n3933) );
  XNOR U3347 ( .A(n3930), .B(n3672), .Z(n3932) );
  IV U3348 ( .A(p_input[8066]), .Z(n3672) );
  XNOR U3349 ( .A(n3934), .B(n3935), .Z(n3930) );
  AND U3350 ( .A(n3936), .B(n3937), .Z(n3935) );
  XOR U3351 ( .A(p_input[8097]), .B(n3934), .Z(n3937) );
  XNOR U3352 ( .A(p_input[8065]), .B(n3934), .Z(n3936) );
  AND U3353 ( .A(p_input[8096]), .B(n3938), .Z(n3934) );
  IV U3354 ( .A(p_input[8064]), .Z(n3938) );
  XOR U3355 ( .A(n3939), .B(n3940), .Z(n3028) );
  AND U3356 ( .A(n437), .B(n3941), .Z(n3940) );
  XNOR U3357 ( .A(n3942), .B(n3939), .Z(n3941) );
  XOR U3358 ( .A(n3943), .B(n3944), .Z(n437) );
  AND U3359 ( .A(n3945), .B(n3946), .Z(n3944) );
  XNOR U3360 ( .A(n3043), .B(n3943), .Z(n3946) );
  AND U3361 ( .A(p_input[8063]), .B(p_input[8031]), .Z(n3043) );
  XNOR U3362 ( .A(n3943), .B(n3040), .Z(n3945) );
  IV U3363 ( .A(n3947), .Z(n3040) );
  AND U3364 ( .A(p_input[7967]), .B(p_input[7999]), .Z(n3947) );
  XOR U3365 ( .A(n3948), .B(n3949), .Z(n3943) );
  AND U3366 ( .A(n3950), .B(n3951), .Z(n3949) );
  XOR U3367 ( .A(n3948), .B(n3055), .Z(n3951) );
  XNOR U3368 ( .A(p_input[8030]), .B(n3952), .Z(n3055) );
  AND U3369 ( .A(n191), .B(n3953), .Z(n3952) );
  XOR U3370 ( .A(p_input[8062]), .B(p_input[8030]), .Z(n3953) );
  XNOR U3371 ( .A(n3052), .B(n3948), .Z(n3950) );
  XOR U3372 ( .A(n3954), .B(n3955), .Z(n3052) );
  AND U3373 ( .A(n188), .B(n3956), .Z(n3955) );
  XOR U3374 ( .A(p_input[7998]), .B(p_input[7966]), .Z(n3956) );
  XOR U3375 ( .A(n3957), .B(n3958), .Z(n3948) );
  AND U3376 ( .A(n3959), .B(n3960), .Z(n3958) );
  XOR U3377 ( .A(n3957), .B(n3067), .Z(n3960) );
  XNOR U3378 ( .A(p_input[8029]), .B(n3961), .Z(n3067) );
  AND U3379 ( .A(n191), .B(n3962), .Z(n3961) );
  XOR U3380 ( .A(p_input[8061]), .B(p_input[8029]), .Z(n3962) );
  XNOR U3381 ( .A(n3064), .B(n3957), .Z(n3959) );
  XOR U3382 ( .A(n3963), .B(n3964), .Z(n3064) );
  AND U3383 ( .A(n188), .B(n3965), .Z(n3964) );
  XOR U3384 ( .A(p_input[7997]), .B(p_input[7965]), .Z(n3965) );
  XOR U3385 ( .A(n3966), .B(n3967), .Z(n3957) );
  AND U3386 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U3387 ( .A(n3966), .B(n3079), .Z(n3969) );
  XNOR U3388 ( .A(p_input[8028]), .B(n3970), .Z(n3079) );
  AND U3389 ( .A(n191), .B(n3971), .Z(n3970) );
  XOR U3390 ( .A(p_input[8060]), .B(p_input[8028]), .Z(n3971) );
  XNOR U3391 ( .A(n3076), .B(n3966), .Z(n3968) );
  XOR U3392 ( .A(n3972), .B(n3973), .Z(n3076) );
  AND U3393 ( .A(n188), .B(n3974), .Z(n3973) );
  XOR U3394 ( .A(p_input[7996]), .B(p_input[7964]), .Z(n3974) );
  XOR U3395 ( .A(n3975), .B(n3976), .Z(n3966) );
  AND U3396 ( .A(n3977), .B(n3978), .Z(n3976) );
  XOR U3397 ( .A(n3975), .B(n3091), .Z(n3978) );
  XNOR U3398 ( .A(p_input[8027]), .B(n3979), .Z(n3091) );
  AND U3399 ( .A(n191), .B(n3980), .Z(n3979) );
  XOR U3400 ( .A(p_input[8059]), .B(p_input[8027]), .Z(n3980) );
  XNOR U3401 ( .A(n3088), .B(n3975), .Z(n3977) );
  XOR U3402 ( .A(n3981), .B(n3982), .Z(n3088) );
  AND U3403 ( .A(n188), .B(n3983), .Z(n3982) );
  XOR U3404 ( .A(p_input[7995]), .B(p_input[7963]), .Z(n3983) );
  XOR U3405 ( .A(n3984), .B(n3985), .Z(n3975) );
  AND U3406 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U3407 ( .A(n3984), .B(n3103), .Z(n3987) );
  XNOR U3408 ( .A(p_input[8026]), .B(n3988), .Z(n3103) );
  AND U3409 ( .A(n191), .B(n3989), .Z(n3988) );
  XOR U3410 ( .A(p_input[8058]), .B(p_input[8026]), .Z(n3989) );
  XNOR U3411 ( .A(n3100), .B(n3984), .Z(n3986) );
  XOR U3412 ( .A(n3990), .B(n3991), .Z(n3100) );
  AND U3413 ( .A(n188), .B(n3992), .Z(n3991) );
  XOR U3414 ( .A(p_input[7994]), .B(p_input[7962]), .Z(n3992) );
  XOR U3415 ( .A(n3993), .B(n3994), .Z(n3984) );
  AND U3416 ( .A(n3995), .B(n3996), .Z(n3994) );
  XOR U3417 ( .A(n3993), .B(n3115), .Z(n3996) );
  XNOR U3418 ( .A(p_input[8025]), .B(n3997), .Z(n3115) );
  AND U3419 ( .A(n191), .B(n3998), .Z(n3997) );
  XOR U3420 ( .A(p_input[8057]), .B(p_input[8025]), .Z(n3998) );
  XNOR U3421 ( .A(n3112), .B(n3993), .Z(n3995) );
  XOR U3422 ( .A(n3999), .B(n4000), .Z(n3112) );
  AND U3423 ( .A(n188), .B(n4001), .Z(n4000) );
  XOR U3424 ( .A(p_input[7993]), .B(p_input[7961]), .Z(n4001) );
  XOR U3425 ( .A(n4002), .B(n4003), .Z(n3993) );
  AND U3426 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U3427 ( .A(n4002), .B(n3127), .Z(n4005) );
  XNOR U3428 ( .A(p_input[8024]), .B(n4006), .Z(n3127) );
  AND U3429 ( .A(n191), .B(n4007), .Z(n4006) );
  XOR U3430 ( .A(p_input[8056]), .B(p_input[8024]), .Z(n4007) );
  XNOR U3431 ( .A(n3124), .B(n4002), .Z(n4004) );
  XOR U3432 ( .A(n4008), .B(n4009), .Z(n3124) );
  AND U3433 ( .A(n188), .B(n4010), .Z(n4009) );
  XOR U3434 ( .A(p_input[7992]), .B(p_input[7960]), .Z(n4010) );
  XOR U3435 ( .A(n4011), .B(n4012), .Z(n4002) );
  AND U3436 ( .A(n4013), .B(n4014), .Z(n4012) );
  XOR U3437 ( .A(n4011), .B(n3139), .Z(n4014) );
  XNOR U3438 ( .A(p_input[8023]), .B(n4015), .Z(n3139) );
  AND U3439 ( .A(n191), .B(n4016), .Z(n4015) );
  XOR U3440 ( .A(p_input[8055]), .B(p_input[8023]), .Z(n4016) );
  XNOR U3441 ( .A(n3136), .B(n4011), .Z(n4013) );
  XOR U3442 ( .A(n4017), .B(n4018), .Z(n3136) );
  AND U3443 ( .A(n188), .B(n4019), .Z(n4018) );
  XOR U3444 ( .A(p_input[7991]), .B(p_input[7959]), .Z(n4019) );
  XOR U3445 ( .A(n4020), .B(n4021), .Z(n4011) );
  AND U3446 ( .A(n4022), .B(n4023), .Z(n4021) );
  XOR U3447 ( .A(n4020), .B(n3151), .Z(n4023) );
  XNOR U3448 ( .A(p_input[8022]), .B(n4024), .Z(n3151) );
  AND U3449 ( .A(n191), .B(n4025), .Z(n4024) );
  XOR U3450 ( .A(p_input[8054]), .B(p_input[8022]), .Z(n4025) );
  XNOR U3451 ( .A(n3148), .B(n4020), .Z(n4022) );
  XOR U3452 ( .A(n4026), .B(n4027), .Z(n3148) );
  AND U3453 ( .A(n188), .B(n4028), .Z(n4027) );
  XOR U3454 ( .A(p_input[7990]), .B(p_input[7958]), .Z(n4028) );
  XOR U3455 ( .A(n4029), .B(n4030), .Z(n4020) );
  AND U3456 ( .A(n4031), .B(n4032), .Z(n4030) );
  XOR U3457 ( .A(n4029), .B(n3163), .Z(n4032) );
  XNOR U3458 ( .A(p_input[8021]), .B(n4033), .Z(n3163) );
  AND U3459 ( .A(n191), .B(n4034), .Z(n4033) );
  XOR U3460 ( .A(p_input[8053]), .B(p_input[8021]), .Z(n4034) );
  XNOR U3461 ( .A(n3160), .B(n4029), .Z(n4031) );
  XOR U3462 ( .A(n4035), .B(n4036), .Z(n3160) );
  AND U3463 ( .A(n188), .B(n4037), .Z(n4036) );
  XOR U3464 ( .A(p_input[7989]), .B(p_input[7957]), .Z(n4037) );
  XOR U3465 ( .A(n4038), .B(n4039), .Z(n4029) );
  AND U3466 ( .A(n4040), .B(n4041), .Z(n4039) );
  XOR U3467 ( .A(n4038), .B(n3175), .Z(n4041) );
  XNOR U3468 ( .A(p_input[8020]), .B(n4042), .Z(n3175) );
  AND U3469 ( .A(n191), .B(n4043), .Z(n4042) );
  XOR U3470 ( .A(p_input[8052]), .B(p_input[8020]), .Z(n4043) );
  XNOR U3471 ( .A(n3172), .B(n4038), .Z(n4040) );
  XOR U3472 ( .A(n4044), .B(n4045), .Z(n3172) );
  AND U3473 ( .A(n188), .B(n4046), .Z(n4045) );
  XOR U3474 ( .A(p_input[7988]), .B(p_input[7956]), .Z(n4046) );
  XOR U3475 ( .A(n4047), .B(n4048), .Z(n4038) );
  AND U3476 ( .A(n4049), .B(n4050), .Z(n4048) );
  XOR U3477 ( .A(n4047), .B(n3187), .Z(n4050) );
  XNOR U3478 ( .A(p_input[8019]), .B(n4051), .Z(n3187) );
  AND U3479 ( .A(n191), .B(n4052), .Z(n4051) );
  XOR U3480 ( .A(p_input[8051]), .B(p_input[8019]), .Z(n4052) );
  XNOR U3481 ( .A(n3184), .B(n4047), .Z(n4049) );
  XOR U3482 ( .A(n4053), .B(n4054), .Z(n3184) );
  AND U3483 ( .A(n188), .B(n4055), .Z(n4054) );
  XOR U3484 ( .A(p_input[7987]), .B(p_input[7955]), .Z(n4055) );
  XOR U3485 ( .A(n4056), .B(n4057), .Z(n4047) );
  AND U3486 ( .A(n4058), .B(n4059), .Z(n4057) );
  XOR U3487 ( .A(n4056), .B(n3199), .Z(n4059) );
  XNOR U3488 ( .A(p_input[8018]), .B(n4060), .Z(n3199) );
  AND U3489 ( .A(n191), .B(n4061), .Z(n4060) );
  XOR U3490 ( .A(p_input[8050]), .B(p_input[8018]), .Z(n4061) );
  XNOR U3491 ( .A(n3196), .B(n4056), .Z(n4058) );
  XOR U3492 ( .A(n4062), .B(n4063), .Z(n3196) );
  AND U3493 ( .A(n188), .B(n4064), .Z(n4063) );
  XOR U3494 ( .A(p_input[7986]), .B(p_input[7954]), .Z(n4064) );
  XOR U3495 ( .A(n4065), .B(n4066), .Z(n4056) );
  AND U3496 ( .A(n4067), .B(n4068), .Z(n4066) );
  XOR U3497 ( .A(n4065), .B(n3211), .Z(n4068) );
  XNOR U3498 ( .A(p_input[8017]), .B(n4069), .Z(n3211) );
  AND U3499 ( .A(n191), .B(n4070), .Z(n4069) );
  XOR U3500 ( .A(p_input[8049]), .B(p_input[8017]), .Z(n4070) );
  XNOR U3501 ( .A(n3208), .B(n4065), .Z(n4067) );
  XOR U3502 ( .A(n4071), .B(n4072), .Z(n3208) );
  AND U3503 ( .A(n188), .B(n4073), .Z(n4072) );
  XOR U3504 ( .A(p_input[7985]), .B(p_input[7953]), .Z(n4073) );
  XOR U3505 ( .A(n4074), .B(n4075), .Z(n4065) );
  AND U3506 ( .A(n4076), .B(n4077), .Z(n4075) );
  XOR U3507 ( .A(n4074), .B(n3223), .Z(n4077) );
  XNOR U3508 ( .A(p_input[8016]), .B(n4078), .Z(n3223) );
  AND U3509 ( .A(n191), .B(n4079), .Z(n4078) );
  XOR U3510 ( .A(p_input[8048]), .B(p_input[8016]), .Z(n4079) );
  XNOR U3511 ( .A(n3220), .B(n4074), .Z(n4076) );
  XOR U3512 ( .A(n4080), .B(n4081), .Z(n3220) );
  AND U3513 ( .A(n188), .B(n4082), .Z(n4081) );
  XOR U3514 ( .A(p_input[7984]), .B(p_input[7952]), .Z(n4082) );
  XOR U3515 ( .A(n4083), .B(n4084), .Z(n4074) );
  AND U3516 ( .A(n4085), .B(n4086), .Z(n4084) );
  XOR U3517 ( .A(n4083), .B(n3235), .Z(n4086) );
  XNOR U3518 ( .A(p_input[8015]), .B(n4087), .Z(n3235) );
  AND U3519 ( .A(n191), .B(n4088), .Z(n4087) );
  XOR U3520 ( .A(p_input[8047]), .B(p_input[8015]), .Z(n4088) );
  XNOR U3521 ( .A(n3232), .B(n4083), .Z(n4085) );
  XOR U3522 ( .A(n4089), .B(n4090), .Z(n3232) );
  AND U3523 ( .A(n188), .B(n4091), .Z(n4090) );
  XOR U3524 ( .A(p_input[7983]), .B(p_input[7951]), .Z(n4091) );
  XOR U3525 ( .A(n4092), .B(n4093), .Z(n4083) );
  AND U3526 ( .A(n4094), .B(n4095), .Z(n4093) );
  XOR U3527 ( .A(n4092), .B(n3247), .Z(n4095) );
  XNOR U3528 ( .A(p_input[8014]), .B(n4096), .Z(n3247) );
  AND U3529 ( .A(n191), .B(n4097), .Z(n4096) );
  XOR U3530 ( .A(p_input[8046]), .B(p_input[8014]), .Z(n4097) );
  XNOR U3531 ( .A(n3244), .B(n4092), .Z(n4094) );
  XOR U3532 ( .A(n4098), .B(n4099), .Z(n3244) );
  AND U3533 ( .A(n188), .B(n4100), .Z(n4099) );
  XOR U3534 ( .A(p_input[7982]), .B(p_input[7950]), .Z(n4100) );
  XOR U3535 ( .A(n4101), .B(n4102), .Z(n4092) );
  AND U3536 ( .A(n4103), .B(n4104), .Z(n4102) );
  XOR U3537 ( .A(n4101), .B(n3259), .Z(n4104) );
  XNOR U3538 ( .A(p_input[8013]), .B(n4105), .Z(n3259) );
  AND U3539 ( .A(n191), .B(n4106), .Z(n4105) );
  XOR U3540 ( .A(p_input[8045]), .B(p_input[8013]), .Z(n4106) );
  XNOR U3541 ( .A(n3256), .B(n4101), .Z(n4103) );
  XOR U3542 ( .A(n4107), .B(n4108), .Z(n3256) );
  AND U3543 ( .A(n188), .B(n4109), .Z(n4108) );
  XOR U3544 ( .A(p_input[7981]), .B(p_input[7949]), .Z(n4109) );
  XOR U3545 ( .A(n4110), .B(n4111), .Z(n4101) );
  AND U3546 ( .A(n4112), .B(n4113), .Z(n4111) );
  XOR U3547 ( .A(n4110), .B(n3271), .Z(n4113) );
  XNOR U3548 ( .A(p_input[8012]), .B(n4114), .Z(n3271) );
  AND U3549 ( .A(n191), .B(n4115), .Z(n4114) );
  XOR U3550 ( .A(p_input[8044]), .B(p_input[8012]), .Z(n4115) );
  XNOR U3551 ( .A(n3268), .B(n4110), .Z(n4112) );
  XOR U3552 ( .A(n4116), .B(n4117), .Z(n3268) );
  AND U3553 ( .A(n188), .B(n4118), .Z(n4117) );
  XOR U3554 ( .A(p_input[7980]), .B(p_input[7948]), .Z(n4118) );
  XOR U3555 ( .A(n4119), .B(n4120), .Z(n4110) );
  AND U3556 ( .A(n4121), .B(n4122), .Z(n4120) );
  XOR U3557 ( .A(n4119), .B(n3283), .Z(n4122) );
  XNOR U3558 ( .A(p_input[8011]), .B(n4123), .Z(n3283) );
  AND U3559 ( .A(n191), .B(n4124), .Z(n4123) );
  XOR U3560 ( .A(p_input[8043]), .B(p_input[8011]), .Z(n4124) );
  XNOR U3561 ( .A(n3280), .B(n4119), .Z(n4121) );
  XOR U3562 ( .A(n4125), .B(n4126), .Z(n3280) );
  AND U3563 ( .A(n188), .B(n4127), .Z(n4126) );
  XOR U3564 ( .A(p_input[7979]), .B(p_input[7947]), .Z(n4127) );
  XOR U3565 ( .A(n4128), .B(n4129), .Z(n4119) );
  AND U3566 ( .A(n4130), .B(n4131), .Z(n4129) );
  XOR U3567 ( .A(n4128), .B(n3295), .Z(n4131) );
  XNOR U3568 ( .A(p_input[8010]), .B(n4132), .Z(n3295) );
  AND U3569 ( .A(n191), .B(n4133), .Z(n4132) );
  XOR U3570 ( .A(p_input[8042]), .B(p_input[8010]), .Z(n4133) );
  XNOR U3571 ( .A(n3292), .B(n4128), .Z(n4130) );
  XOR U3572 ( .A(n4134), .B(n4135), .Z(n3292) );
  AND U3573 ( .A(n188), .B(n4136), .Z(n4135) );
  XOR U3574 ( .A(p_input[7978]), .B(p_input[7946]), .Z(n4136) );
  XOR U3575 ( .A(n4137), .B(n4138), .Z(n4128) );
  AND U3576 ( .A(n4139), .B(n4140), .Z(n4138) );
  XOR U3577 ( .A(n4137), .B(n3307), .Z(n4140) );
  XNOR U3578 ( .A(p_input[8009]), .B(n4141), .Z(n3307) );
  AND U3579 ( .A(n191), .B(n4142), .Z(n4141) );
  XOR U3580 ( .A(p_input[8041]), .B(p_input[8009]), .Z(n4142) );
  XNOR U3581 ( .A(n3304), .B(n4137), .Z(n4139) );
  XOR U3582 ( .A(n4143), .B(n4144), .Z(n3304) );
  AND U3583 ( .A(n188), .B(n4145), .Z(n4144) );
  XOR U3584 ( .A(p_input[7977]), .B(p_input[7945]), .Z(n4145) );
  XOR U3585 ( .A(n4146), .B(n4147), .Z(n4137) );
  AND U3586 ( .A(n4148), .B(n4149), .Z(n4147) );
  XOR U3587 ( .A(n4146), .B(n3319), .Z(n4149) );
  XNOR U3588 ( .A(p_input[8008]), .B(n4150), .Z(n3319) );
  AND U3589 ( .A(n191), .B(n4151), .Z(n4150) );
  XOR U3590 ( .A(p_input[8040]), .B(p_input[8008]), .Z(n4151) );
  XNOR U3591 ( .A(n3316), .B(n4146), .Z(n4148) );
  XOR U3592 ( .A(n4152), .B(n4153), .Z(n3316) );
  AND U3593 ( .A(n188), .B(n4154), .Z(n4153) );
  XOR U3594 ( .A(p_input[7976]), .B(p_input[7944]), .Z(n4154) );
  XOR U3595 ( .A(n4155), .B(n4156), .Z(n4146) );
  AND U3596 ( .A(n4157), .B(n4158), .Z(n4156) );
  XOR U3597 ( .A(n4155), .B(n3331), .Z(n4158) );
  XNOR U3598 ( .A(p_input[8007]), .B(n4159), .Z(n3331) );
  AND U3599 ( .A(n191), .B(n4160), .Z(n4159) );
  XOR U3600 ( .A(p_input[8039]), .B(p_input[8007]), .Z(n4160) );
  XNOR U3601 ( .A(n3328), .B(n4155), .Z(n4157) );
  XOR U3602 ( .A(n4161), .B(n4162), .Z(n3328) );
  AND U3603 ( .A(n188), .B(n4163), .Z(n4162) );
  XOR U3604 ( .A(p_input[7975]), .B(p_input[7943]), .Z(n4163) );
  XOR U3605 ( .A(n4164), .B(n4165), .Z(n4155) );
  AND U3606 ( .A(n4166), .B(n4167), .Z(n4165) );
  XOR U3607 ( .A(n4164), .B(n3343), .Z(n4167) );
  XNOR U3608 ( .A(p_input[8006]), .B(n4168), .Z(n3343) );
  AND U3609 ( .A(n191), .B(n4169), .Z(n4168) );
  XOR U3610 ( .A(p_input[8038]), .B(p_input[8006]), .Z(n4169) );
  XNOR U3611 ( .A(n3340), .B(n4164), .Z(n4166) );
  XOR U3612 ( .A(n4170), .B(n4171), .Z(n3340) );
  AND U3613 ( .A(n188), .B(n4172), .Z(n4171) );
  XOR U3614 ( .A(p_input[7974]), .B(p_input[7942]), .Z(n4172) );
  XOR U3615 ( .A(n4173), .B(n4174), .Z(n4164) );
  AND U3616 ( .A(n4175), .B(n4176), .Z(n4174) );
  XOR U3617 ( .A(n4173), .B(n3355), .Z(n4176) );
  XNOR U3618 ( .A(p_input[8005]), .B(n4177), .Z(n3355) );
  AND U3619 ( .A(n191), .B(n4178), .Z(n4177) );
  XOR U3620 ( .A(p_input[8037]), .B(p_input[8005]), .Z(n4178) );
  XNOR U3621 ( .A(n3352), .B(n4173), .Z(n4175) );
  XOR U3622 ( .A(n4179), .B(n4180), .Z(n3352) );
  AND U3623 ( .A(n188), .B(n4181), .Z(n4180) );
  XOR U3624 ( .A(p_input[7973]), .B(p_input[7941]), .Z(n4181) );
  XOR U3625 ( .A(n4182), .B(n4183), .Z(n4173) );
  AND U3626 ( .A(n4184), .B(n4185), .Z(n4183) );
  XOR U3627 ( .A(n4182), .B(n3367), .Z(n4185) );
  XNOR U3628 ( .A(p_input[8004]), .B(n4186), .Z(n3367) );
  AND U3629 ( .A(n191), .B(n4187), .Z(n4186) );
  XOR U3630 ( .A(p_input[8036]), .B(p_input[8004]), .Z(n4187) );
  XNOR U3631 ( .A(n3364), .B(n4182), .Z(n4184) );
  XOR U3632 ( .A(n4188), .B(n4189), .Z(n3364) );
  AND U3633 ( .A(n188), .B(n4190), .Z(n4189) );
  XOR U3634 ( .A(p_input[7972]), .B(p_input[7940]), .Z(n4190) );
  XOR U3635 ( .A(n4191), .B(n4192), .Z(n4182) );
  AND U3636 ( .A(n4193), .B(n4194), .Z(n4192) );
  XOR U3637 ( .A(n4191), .B(n3379), .Z(n4194) );
  XNOR U3638 ( .A(p_input[8003]), .B(n4195), .Z(n3379) );
  AND U3639 ( .A(n191), .B(n4196), .Z(n4195) );
  XOR U3640 ( .A(p_input[8035]), .B(p_input[8003]), .Z(n4196) );
  XNOR U3641 ( .A(n3376), .B(n4191), .Z(n4193) );
  XOR U3642 ( .A(n4197), .B(n4198), .Z(n3376) );
  AND U3643 ( .A(n188), .B(n4199), .Z(n4198) );
  XOR U3644 ( .A(p_input[7971]), .B(p_input[7939]), .Z(n4199) );
  XOR U3645 ( .A(n4200), .B(n4201), .Z(n4191) );
  AND U3646 ( .A(n4202), .B(n4203), .Z(n4201) );
  XOR U3647 ( .A(n4200), .B(n3391), .Z(n4203) );
  XNOR U3648 ( .A(p_input[8002]), .B(n4204), .Z(n3391) );
  AND U3649 ( .A(n191), .B(n4205), .Z(n4204) );
  XOR U3650 ( .A(p_input[8034]), .B(p_input[8002]), .Z(n4205) );
  XNOR U3651 ( .A(n3388), .B(n4200), .Z(n4202) );
  XOR U3652 ( .A(n4206), .B(n4207), .Z(n3388) );
  AND U3653 ( .A(n188), .B(n4208), .Z(n4207) );
  XOR U3654 ( .A(p_input[7970]), .B(p_input[7938]), .Z(n4208) );
  XOR U3655 ( .A(n4209), .B(n4210), .Z(n4200) );
  AND U3656 ( .A(n4211), .B(n4212), .Z(n4210) );
  XNOR U3657 ( .A(n4213), .B(n3404), .Z(n4212) );
  XNOR U3658 ( .A(p_input[8001]), .B(n4214), .Z(n3404) );
  AND U3659 ( .A(n191), .B(n4215), .Z(n4214) );
  XNOR U3660 ( .A(p_input[8033]), .B(n4216), .Z(n4215) );
  IV U3661 ( .A(p_input[8001]), .Z(n4216) );
  XNOR U3662 ( .A(n3401), .B(n4209), .Z(n4211) );
  XNOR U3663 ( .A(p_input[7937]), .B(n4217), .Z(n3401) );
  AND U3664 ( .A(n188), .B(n4218), .Z(n4217) );
  XOR U3665 ( .A(p_input[7969]), .B(p_input[7937]), .Z(n4218) );
  IV U3666 ( .A(n4213), .Z(n4209) );
  AND U3667 ( .A(n3939), .B(n3942), .Z(n4213) );
  XOR U3668 ( .A(p_input[8000]), .B(n4219), .Z(n3942) );
  AND U3669 ( .A(n191), .B(n4220), .Z(n4219) );
  XOR U3670 ( .A(p_input[8032]), .B(p_input[8000]), .Z(n4220) );
  XOR U3671 ( .A(n4221), .B(n4222), .Z(n191) );
  AND U3672 ( .A(n4223), .B(n4224), .Z(n4222) );
  XNOR U3673 ( .A(p_input[8063]), .B(n4221), .Z(n4224) );
  XOR U3674 ( .A(n4221), .B(p_input[8031]), .Z(n4223) );
  XOR U3675 ( .A(n4225), .B(n4226), .Z(n4221) );
  AND U3676 ( .A(n4227), .B(n4228), .Z(n4226) );
  XNOR U3677 ( .A(p_input[8062]), .B(n4225), .Z(n4228) );
  XOR U3678 ( .A(n4225), .B(p_input[8030]), .Z(n4227) );
  XOR U3679 ( .A(n4229), .B(n4230), .Z(n4225) );
  AND U3680 ( .A(n4231), .B(n4232), .Z(n4230) );
  XNOR U3681 ( .A(p_input[8061]), .B(n4229), .Z(n4232) );
  XOR U3682 ( .A(n4229), .B(p_input[8029]), .Z(n4231) );
  XOR U3683 ( .A(n4233), .B(n4234), .Z(n4229) );
  AND U3684 ( .A(n4235), .B(n4236), .Z(n4234) );
  XNOR U3685 ( .A(p_input[8060]), .B(n4233), .Z(n4236) );
  XOR U3686 ( .A(n4233), .B(p_input[8028]), .Z(n4235) );
  XOR U3687 ( .A(n4237), .B(n4238), .Z(n4233) );
  AND U3688 ( .A(n4239), .B(n4240), .Z(n4238) );
  XNOR U3689 ( .A(p_input[8059]), .B(n4237), .Z(n4240) );
  XOR U3690 ( .A(n4237), .B(p_input[8027]), .Z(n4239) );
  XOR U3691 ( .A(n4241), .B(n4242), .Z(n4237) );
  AND U3692 ( .A(n4243), .B(n4244), .Z(n4242) );
  XNOR U3693 ( .A(p_input[8058]), .B(n4241), .Z(n4244) );
  XOR U3694 ( .A(n4241), .B(p_input[8026]), .Z(n4243) );
  XOR U3695 ( .A(n4245), .B(n4246), .Z(n4241) );
  AND U3696 ( .A(n4247), .B(n4248), .Z(n4246) );
  XNOR U3697 ( .A(p_input[8057]), .B(n4245), .Z(n4248) );
  XOR U3698 ( .A(n4245), .B(p_input[8025]), .Z(n4247) );
  XOR U3699 ( .A(n4249), .B(n4250), .Z(n4245) );
  AND U3700 ( .A(n4251), .B(n4252), .Z(n4250) );
  XNOR U3701 ( .A(p_input[8056]), .B(n4249), .Z(n4252) );
  XOR U3702 ( .A(n4249), .B(p_input[8024]), .Z(n4251) );
  XOR U3703 ( .A(n4253), .B(n4254), .Z(n4249) );
  AND U3704 ( .A(n4255), .B(n4256), .Z(n4254) );
  XNOR U3705 ( .A(p_input[8055]), .B(n4253), .Z(n4256) );
  XOR U3706 ( .A(n4253), .B(p_input[8023]), .Z(n4255) );
  XOR U3707 ( .A(n4257), .B(n4258), .Z(n4253) );
  AND U3708 ( .A(n4259), .B(n4260), .Z(n4258) );
  XNOR U3709 ( .A(p_input[8054]), .B(n4257), .Z(n4260) );
  XOR U3710 ( .A(n4257), .B(p_input[8022]), .Z(n4259) );
  XOR U3711 ( .A(n4261), .B(n4262), .Z(n4257) );
  AND U3712 ( .A(n4263), .B(n4264), .Z(n4262) );
  XNOR U3713 ( .A(p_input[8053]), .B(n4261), .Z(n4264) );
  XOR U3714 ( .A(n4261), .B(p_input[8021]), .Z(n4263) );
  XOR U3715 ( .A(n4265), .B(n4266), .Z(n4261) );
  AND U3716 ( .A(n4267), .B(n4268), .Z(n4266) );
  XNOR U3717 ( .A(p_input[8052]), .B(n4265), .Z(n4268) );
  XOR U3718 ( .A(n4265), .B(p_input[8020]), .Z(n4267) );
  XOR U3719 ( .A(n4269), .B(n4270), .Z(n4265) );
  AND U3720 ( .A(n4271), .B(n4272), .Z(n4270) );
  XNOR U3721 ( .A(p_input[8051]), .B(n4269), .Z(n4272) );
  XOR U3722 ( .A(n4269), .B(p_input[8019]), .Z(n4271) );
  XOR U3723 ( .A(n4273), .B(n4274), .Z(n4269) );
  AND U3724 ( .A(n4275), .B(n4276), .Z(n4274) );
  XNOR U3725 ( .A(p_input[8050]), .B(n4273), .Z(n4276) );
  XOR U3726 ( .A(n4273), .B(p_input[8018]), .Z(n4275) );
  XOR U3727 ( .A(n4277), .B(n4278), .Z(n4273) );
  AND U3728 ( .A(n4279), .B(n4280), .Z(n4278) );
  XNOR U3729 ( .A(p_input[8049]), .B(n4277), .Z(n4280) );
  XOR U3730 ( .A(n4277), .B(p_input[8017]), .Z(n4279) );
  XOR U3731 ( .A(n4281), .B(n4282), .Z(n4277) );
  AND U3732 ( .A(n4283), .B(n4284), .Z(n4282) );
  XNOR U3733 ( .A(p_input[8048]), .B(n4281), .Z(n4284) );
  XOR U3734 ( .A(n4281), .B(p_input[8016]), .Z(n4283) );
  XOR U3735 ( .A(n4285), .B(n4286), .Z(n4281) );
  AND U3736 ( .A(n4287), .B(n4288), .Z(n4286) );
  XNOR U3737 ( .A(p_input[8047]), .B(n4285), .Z(n4288) );
  XOR U3738 ( .A(n4285), .B(p_input[8015]), .Z(n4287) );
  XOR U3739 ( .A(n4289), .B(n4290), .Z(n4285) );
  AND U3740 ( .A(n4291), .B(n4292), .Z(n4290) );
  XNOR U3741 ( .A(p_input[8046]), .B(n4289), .Z(n4292) );
  XOR U3742 ( .A(n4289), .B(p_input[8014]), .Z(n4291) );
  XOR U3743 ( .A(n4293), .B(n4294), .Z(n4289) );
  AND U3744 ( .A(n4295), .B(n4296), .Z(n4294) );
  XNOR U3745 ( .A(p_input[8045]), .B(n4293), .Z(n4296) );
  XOR U3746 ( .A(n4293), .B(p_input[8013]), .Z(n4295) );
  XOR U3747 ( .A(n4297), .B(n4298), .Z(n4293) );
  AND U3748 ( .A(n4299), .B(n4300), .Z(n4298) );
  XNOR U3749 ( .A(p_input[8044]), .B(n4297), .Z(n4300) );
  XOR U3750 ( .A(n4297), .B(p_input[8012]), .Z(n4299) );
  XOR U3751 ( .A(n4301), .B(n4302), .Z(n4297) );
  AND U3752 ( .A(n4303), .B(n4304), .Z(n4302) );
  XNOR U3753 ( .A(p_input[8043]), .B(n4301), .Z(n4304) );
  XOR U3754 ( .A(n4301), .B(p_input[8011]), .Z(n4303) );
  XOR U3755 ( .A(n4305), .B(n4306), .Z(n4301) );
  AND U3756 ( .A(n4307), .B(n4308), .Z(n4306) );
  XNOR U3757 ( .A(p_input[8042]), .B(n4305), .Z(n4308) );
  XOR U3758 ( .A(n4305), .B(p_input[8010]), .Z(n4307) );
  XOR U3759 ( .A(n4309), .B(n4310), .Z(n4305) );
  AND U3760 ( .A(n4311), .B(n4312), .Z(n4310) );
  XNOR U3761 ( .A(p_input[8041]), .B(n4309), .Z(n4312) );
  XOR U3762 ( .A(n4309), .B(p_input[8009]), .Z(n4311) );
  XOR U3763 ( .A(n4313), .B(n4314), .Z(n4309) );
  AND U3764 ( .A(n4315), .B(n4316), .Z(n4314) );
  XNOR U3765 ( .A(p_input[8040]), .B(n4313), .Z(n4316) );
  XOR U3766 ( .A(n4313), .B(p_input[8008]), .Z(n4315) );
  XOR U3767 ( .A(n4317), .B(n4318), .Z(n4313) );
  AND U3768 ( .A(n4319), .B(n4320), .Z(n4318) );
  XNOR U3769 ( .A(p_input[8039]), .B(n4317), .Z(n4320) );
  XOR U3770 ( .A(n4317), .B(p_input[8007]), .Z(n4319) );
  XOR U3771 ( .A(n4321), .B(n4322), .Z(n4317) );
  AND U3772 ( .A(n4323), .B(n4324), .Z(n4322) );
  XNOR U3773 ( .A(p_input[8038]), .B(n4321), .Z(n4324) );
  XOR U3774 ( .A(n4321), .B(p_input[8006]), .Z(n4323) );
  XOR U3775 ( .A(n4325), .B(n4326), .Z(n4321) );
  AND U3776 ( .A(n4327), .B(n4328), .Z(n4326) );
  XNOR U3777 ( .A(p_input[8037]), .B(n4325), .Z(n4328) );
  XOR U3778 ( .A(n4325), .B(p_input[8005]), .Z(n4327) );
  XOR U3779 ( .A(n4329), .B(n4330), .Z(n4325) );
  AND U3780 ( .A(n4331), .B(n4332), .Z(n4330) );
  XNOR U3781 ( .A(p_input[8036]), .B(n4329), .Z(n4332) );
  XOR U3782 ( .A(n4329), .B(p_input[8004]), .Z(n4331) );
  XOR U3783 ( .A(n4333), .B(n4334), .Z(n4329) );
  AND U3784 ( .A(n4335), .B(n4336), .Z(n4334) );
  XNOR U3785 ( .A(p_input[8035]), .B(n4333), .Z(n4336) );
  XOR U3786 ( .A(n4333), .B(p_input[8003]), .Z(n4335) );
  XOR U3787 ( .A(n4337), .B(n4338), .Z(n4333) );
  AND U3788 ( .A(n4339), .B(n4340), .Z(n4338) );
  XNOR U3789 ( .A(p_input[8034]), .B(n4337), .Z(n4340) );
  XOR U3790 ( .A(n4337), .B(p_input[8002]), .Z(n4339) );
  XNOR U3791 ( .A(n4341), .B(n4342), .Z(n4337) );
  AND U3792 ( .A(n4343), .B(n4344), .Z(n4342) );
  XOR U3793 ( .A(p_input[8033]), .B(n4341), .Z(n4344) );
  XNOR U3794 ( .A(p_input[8001]), .B(n4341), .Z(n4343) );
  AND U3795 ( .A(p_input[8032]), .B(n4345), .Z(n4341) );
  IV U3796 ( .A(p_input[8000]), .Z(n4345) );
  XNOR U3797 ( .A(p_input[7936]), .B(n4346), .Z(n3939) );
  AND U3798 ( .A(n188), .B(n4347), .Z(n4346) );
  XOR U3799 ( .A(p_input[7968]), .B(p_input[7936]), .Z(n4347) );
  XOR U3800 ( .A(n4348), .B(n4349), .Z(n188) );
  AND U3801 ( .A(n4350), .B(n4351), .Z(n4349) );
  XNOR U3802 ( .A(p_input[7999]), .B(n4348), .Z(n4351) );
  XOR U3803 ( .A(n4348), .B(p_input[7967]), .Z(n4350) );
  XOR U3804 ( .A(n4352), .B(n4353), .Z(n4348) );
  AND U3805 ( .A(n4354), .B(n4355), .Z(n4353) );
  XNOR U3806 ( .A(p_input[7998]), .B(n4352), .Z(n4355) );
  XNOR U3807 ( .A(n4352), .B(n3954), .Z(n4354) );
  IV U3808 ( .A(p_input[7966]), .Z(n3954) );
  XOR U3809 ( .A(n4356), .B(n4357), .Z(n4352) );
  AND U3810 ( .A(n4358), .B(n4359), .Z(n4357) );
  XNOR U3811 ( .A(p_input[7997]), .B(n4356), .Z(n4359) );
  XNOR U3812 ( .A(n4356), .B(n3963), .Z(n4358) );
  IV U3813 ( .A(p_input[7965]), .Z(n3963) );
  XOR U3814 ( .A(n4360), .B(n4361), .Z(n4356) );
  AND U3815 ( .A(n4362), .B(n4363), .Z(n4361) );
  XNOR U3816 ( .A(p_input[7996]), .B(n4360), .Z(n4363) );
  XNOR U3817 ( .A(n4360), .B(n3972), .Z(n4362) );
  IV U3818 ( .A(p_input[7964]), .Z(n3972) );
  XOR U3819 ( .A(n4364), .B(n4365), .Z(n4360) );
  AND U3820 ( .A(n4366), .B(n4367), .Z(n4365) );
  XNOR U3821 ( .A(p_input[7995]), .B(n4364), .Z(n4367) );
  XNOR U3822 ( .A(n4364), .B(n3981), .Z(n4366) );
  IV U3823 ( .A(p_input[7963]), .Z(n3981) );
  XOR U3824 ( .A(n4368), .B(n4369), .Z(n4364) );
  AND U3825 ( .A(n4370), .B(n4371), .Z(n4369) );
  XNOR U3826 ( .A(p_input[7994]), .B(n4368), .Z(n4371) );
  XNOR U3827 ( .A(n4368), .B(n3990), .Z(n4370) );
  IV U3828 ( .A(p_input[7962]), .Z(n3990) );
  XOR U3829 ( .A(n4372), .B(n4373), .Z(n4368) );
  AND U3830 ( .A(n4374), .B(n4375), .Z(n4373) );
  XNOR U3831 ( .A(p_input[7993]), .B(n4372), .Z(n4375) );
  XNOR U3832 ( .A(n4372), .B(n3999), .Z(n4374) );
  IV U3833 ( .A(p_input[7961]), .Z(n3999) );
  XOR U3834 ( .A(n4376), .B(n4377), .Z(n4372) );
  AND U3835 ( .A(n4378), .B(n4379), .Z(n4377) );
  XNOR U3836 ( .A(p_input[7992]), .B(n4376), .Z(n4379) );
  XNOR U3837 ( .A(n4376), .B(n4008), .Z(n4378) );
  IV U3838 ( .A(p_input[7960]), .Z(n4008) );
  XOR U3839 ( .A(n4380), .B(n4381), .Z(n4376) );
  AND U3840 ( .A(n4382), .B(n4383), .Z(n4381) );
  XNOR U3841 ( .A(p_input[7991]), .B(n4380), .Z(n4383) );
  XNOR U3842 ( .A(n4380), .B(n4017), .Z(n4382) );
  IV U3843 ( .A(p_input[7959]), .Z(n4017) );
  XOR U3844 ( .A(n4384), .B(n4385), .Z(n4380) );
  AND U3845 ( .A(n4386), .B(n4387), .Z(n4385) );
  XNOR U3846 ( .A(p_input[7990]), .B(n4384), .Z(n4387) );
  XNOR U3847 ( .A(n4384), .B(n4026), .Z(n4386) );
  IV U3848 ( .A(p_input[7958]), .Z(n4026) );
  XOR U3849 ( .A(n4388), .B(n4389), .Z(n4384) );
  AND U3850 ( .A(n4390), .B(n4391), .Z(n4389) );
  XNOR U3851 ( .A(p_input[7989]), .B(n4388), .Z(n4391) );
  XNOR U3852 ( .A(n4388), .B(n4035), .Z(n4390) );
  IV U3853 ( .A(p_input[7957]), .Z(n4035) );
  XOR U3854 ( .A(n4392), .B(n4393), .Z(n4388) );
  AND U3855 ( .A(n4394), .B(n4395), .Z(n4393) );
  XNOR U3856 ( .A(p_input[7988]), .B(n4392), .Z(n4395) );
  XNOR U3857 ( .A(n4392), .B(n4044), .Z(n4394) );
  IV U3858 ( .A(p_input[7956]), .Z(n4044) );
  XOR U3859 ( .A(n4396), .B(n4397), .Z(n4392) );
  AND U3860 ( .A(n4398), .B(n4399), .Z(n4397) );
  XNOR U3861 ( .A(p_input[7987]), .B(n4396), .Z(n4399) );
  XNOR U3862 ( .A(n4396), .B(n4053), .Z(n4398) );
  IV U3863 ( .A(p_input[7955]), .Z(n4053) );
  XOR U3864 ( .A(n4400), .B(n4401), .Z(n4396) );
  AND U3865 ( .A(n4402), .B(n4403), .Z(n4401) );
  XNOR U3866 ( .A(p_input[7986]), .B(n4400), .Z(n4403) );
  XNOR U3867 ( .A(n4400), .B(n4062), .Z(n4402) );
  IV U3868 ( .A(p_input[7954]), .Z(n4062) );
  XOR U3869 ( .A(n4404), .B(n4405), .Z(n4400) );
  AND U3870 ( .A(n4406), .B(n4407), .Z(n4405) );
  XNOR U3871 ( .A(p_input[7985]), .B(n4404), .Z(n4407) );
  XNOR U3872 ( .A(n4404), .B(n4071), .Z(n4406) );
  IV U3873 ( .A(p_input[7953]), .Z(n4071) );
  XOR U3874 ( .A(n4408), .B(n4409), .Z(n4404) );
  AND U3875 ( .A(n4410), .B(n4411), .Z(n4409) );
  XNOR U3876 ( .A(p_input[7984]), .B(n4408), .Z(n4411) );
  XNOR U3877 ( .A(n4408), .B(n4080), .Z(n4410) );
  IV U3878 ( .A(p_input[7952]), .Z(n4080) );
  XOR U3879 ( .A(n4412), .B(n4413), .Z(n4408) );
  AND U3880 ( .A(n4414), .B(n4415), .Z(n4413) );
  XNOR U3881 ( .A(p_input[7983]), .B(n4412), .Z(n4415) );
  XNOR U3882 ( .A(n4412), .B(n4089), .Z(n4414) );
  IV U3883 ( .A(p_input[7951]), .Z(n4089) );
  XOR U3884 ( .A(n4416), .B(n4417), .Z(n4412) );
  AND U3885 ( .A(n4418), .B(n4419), .Z(n4417) );
  XNOR U3886 ( .A(p_input[7982]), .B(n4416), .Z(n4419) );
  XNOR U3887 ( .A(n4416), .B(n4098), .Z(n4418) );
  IV U3888 ( .A(p_input[7950]), .Z(n4098) );
  XOR U3889 ( .A(n4420), .B(n4421), .Z(n4416) );
  AND U3890 ( .A(n4422), .B(n4423), .Z(n4421) );
  XNOR U3891 ( .A(p_input[7981]), .B(n4420), .Z(n4423) );
  XNOR U3892 ( .A(n4420), .B(n4107), .Z(n4422) );
  IV U3893 ( .A(p_input[7949]), .Z(n4107) );
  XOR U3894 ( .A(n4424), .B(n4425), .Z(n4420) );
  AND U3895 ( .A(n4426), .B(n4427), .Z(n4425) );
  XNOR U3896 ( .A(p_input[7980]), .B(n4424), .Z(n4427) );
  XNOR U3897 ( .A(n4424), .B(n4116), .Z(n4426) );
  IV U3898 ( .A(p_input[7948]), .Z(n4116) );
  XOR U3899 ( .A(n4428), .B(n4429), .Z(n4424) );
  AND U3900 ( .A(n4430), .B(n4431), .Z(n4429) );
  XNOR U3901 ( .A(p_input[7979]), .B(n4428), .Z(n4431) );
  XNOR U3902 ( .A(n4428), .B(n4125), .Z(n4430) );
  IV U3903 ( .A(p_input[7947]), .Z(n4125) );
  XOR U3904 ( .A(n4432), .B(n4433), .Z(n4428) );
  AND U3905 ( .A(n4434), .B(n4435), .Z(n4433) );
  XNOR U3906 ( .A(p_input[7978]), .B(n4432), .Z(n4435) );
  XNOR U3907 ( .A(n4432), .B(n4134), .Z(n4434) );
  IV U3908 ( .A(p_input[7946]), .Z(n4134) );
  XOR U3909 ( .A(n4436), .B(n4437), .Z(n4432) );
  AND U3910 ( .A(n4438), .B(n4439), .Z(n4437) );
  XNOR U3911 ( .A(p_input[7977]), .B(n4436), .Z(n4439) );
  XNOR U3912 ( .A(n4436), .B(n4143), .Z(n4438) );
  IV U3913 ( .A(p_input[7945]), .Z(n4143) );
  XOR U3914 ( .A(n4440), .B(n4441), .Z(n4436) );
  AND U3915 ( .A(n4442), .B(n4443), .Z(n4441) );
  XNOR U3916 ( .A(p_input[7976]), .B(n4440), .Z(n4443) );
  XNOR U3917 ( .A(n4440), .B(n4152), .Z(n4442) );
  IV U3918 ( .A(p_input[7944]), .Z(n4152) );
  XOR U3919 ( .A(n4444), .B(n4445), .Z(n4440) );
  AND U3920 ( .A(n4446), .B(n4447), .Z(n4445) );
  XNOR U3921 ( .A(p_input[7975]), .B(n4444), .Z(n4447) );
  XNOR U3922 ( .A(n4444), .B(n4161), .Z(n4446) );
  IV U3923 ( .A(p_input[7943]), .Z(n4161) );
  XOR U3924 ( .A(n4448), .B(n4449), .Z(n4444) );
  AND U3925 ( .A(n4450), .B(n4451), .Z(n4449) );
  XNOR U3926 ( .A(p_input[7974]), .B(n4448), .Z(n4451) );
  XNOR U3927 ( .A(n4448), .B(n4170), .Z(n4450) );
  IV U3928 ( .A(p_input[7942]), .Z(n4170) );
  XOR U3929 ( .A(n4452), .B(n4453), .Z(n4448) );
  AND U3930 ( .A(n4454), .B(n4455), .Z(n4453) );
  XNOR U3931 ( .A(p_input[7973]), .B(n4452), .Z(n4455) );
  XNOR U3932 ( .A(n4452), .B(n4179), .Z(n4454) );
  IV U3933 ( .A(p_input[7941]), .Z(n4179) );
  XOR U3934 ( .A(n4456), .B(n4457), .Z(n4452) );
  AND U3935 ( .A(n4458), .B(n4459), .Z(n4457) );
  XNOR U3936 ( .A(p_input[7972]), .B(n4456), .Z(n4459) );
  XNOR U3937 ( .A(n4456), .B(n4188), .Z(n4458) );
  IV U3938 ( .A(p_input[7940]), .Z(n4188) );
  XOR U3939 ( .A(n4460), .B(n4461), .Z(n4456) );
  AND U3940 ( .A(n4462), .B(n4463), .Z(n4461) );
  XNOR U3941 ( .A(p_input[7971]), .B(n4460), .Z(n4463) );
  XNOR U3942 ( .A(n4460), .B(n4197), .Z(n4462) );
  IV U3943 ( .A(p_input[7939]), .Z(n4197) );
  XOR U3944 ( .A(n4464), .B(n4465), .Z(n4460) );
  AND U3945 ( .A(n4466), .B(n4467), .Z(n4465) );
  XNOR U3946 ( .A(p_input[7970]), .B(n4464), .Z(n4467) );
  XNOR U3947 ( .A(n4464), .B(n4206), .Z(n4466) );
  IV U3948 ( .A(p_input[7938]), .Z(n4206) );
  XNOR U3949 ( .A(n4468), .B(n4469), .Z(n4464) );
  AND U3950 ( .A(n4470), .B(n4471), .Z(n4469) );
  XOR U3951 ( .A(p_input[7969]), .B(n4468), .Z(n4471) );
  XNOR U3952 ( .A(p_input[7937]), .B(n4468), .Z(n4470) );
  AND U3953 ( .A(p_input[7968]), .B(n4472), .Z(n4468) );
  IV U3954 ( .A(p_input[7936]), .Z(n4472) );
  XOR U3955 ( .A(n4473), .B(n4474), .Z(n2651) );
  AND U3956 ( .A(n813), .B(n4475), .Z(n4474) );
  XNOR U3957 ( .A(n4476), .B(n4473), .Z(n4475) );
  XOR U3958 ( .A(n4477), .B(n4478), .Z(n813) );
  AND U3959 ( .A(n4479), .B(n4480), .Z(n4478) );
  XOR U3960 ( .A(n4477), .B(n2666), .Z(n4480) );
  XNOR U3961 ( .A(n4481), .B(n4482), .Z(n2666) );
  AND U3962 ( .A(n4483), .B(n443), .Z(n4482) );
  AND U3963 ( .A(n4481), .B(n4484), .Z(n4483) );
  XNOR U3964 ( .A(n2663), .B(n4477), .Z(n4479) );
  XOR U3965 ( .A(n4485), .B(n4486), .Z(n2663) );
  AND U3966 ( .A(n4487), .B(n440), .Z(n4486) );
  NOR U3967 ( .A(n4485), .B(n4488), .Z(n4487) );
  XOR U3968 ( .A(n4489), .B(n4490), .Z(n4477) );
  AND U3969 ( .A(n4491), .B(n4492), .Z(n4490) );
  XOR U3970 ( .A(n4489), .B(n2678), .Z(n4492) );
  XOR U3971 ( .A(n4493), .B(n4494), .Z(n2678) );
  AND U3972 ( .A(n443), .B(n4495), .Z(n4494) );
  XOR U3973 ( .A(n4496), .B(n4493), .Z(n4495) );
  XNOR U3974 ( .A(n2675), .B(n4489), .Z(n4491) );
  XOR U3975 ( .A(n4497), .B(n4498), .Z(n2675) );
  AND U3976 ( .A(n440), .B(n4499), .Z(n4498) );
  XOR U3977 ( .A(n4500), .B(n4497), .Z(n4499) );
  XOR U3978 ( .A(n4501), .B(n4502), .Z(n4489) );
  AND U3979 ( .A(n4503), .B(n4504), .Z(n4502) );
  XOR U3980 ( .A(n4501), .B(n2690), .Z(n4504) );
  XOR U3981 ( .A(n4505), .B(n4506), .Z(n2690) );
  AND U3982 ( .A(n443), .B(n4507), .Z(n4506) );
  XOR U3983 ( .A(n4508), .B(n4505), .Z(n4507) );
  XNOR U3984 ( .A(n2687), .B(n4501), .Z(n4503) );
  XOR U3985 ( .A(n4509), .B(n4510), .Z(n2687) );
  AND U3986 ( .A(n440), .B(n4511), .Z(n4510) );
  XOR U3987 ( .A(n4512), .B(n4509), .Z(n4511) );
  XOR U3988 ( .A(n4513), .B(n4514), .Z(n4501) );
  AND U3989 ( .A(n4515), .B(n4516), .Z(n4514) );
  XOR U3990 ( .A(n4513), .B(n2702), .Z(n4516) );
  XOR U3991 ( .A(n4517), .B(n4518), .Z(n2702) );
  AND U3992 ( .A(n443), .B(n4519), .Z(n4518) );
  XOR U3993 ( .A(n4520), .B(n4517), .Z(n4519) );
  XNOR U3994 ( .A(n2699), .B(n4513), .Z(n4515) );
  XOR U3995 ( .A(n4521), .B(n4522), .Z(n2699) );
  AND U3996 ( .A(n440), .B(n4523), .Z(n4522) );
  XOR U3997 ( .A(n4524), .B(n4521), .Z(n4523) );
  XOR U3998 ( .A(n4525), .B(n4526), .Z(n4513) );
  AND U3999 ( .A(n4527), .B(n4528), .Z(n4526) );
  XOR U4000 ( .A(n4525), .B(n2714), .Z(n4528) );
  XOR U4001 ( .A(n4529), .B(n4530), .Z(n2714) );
  AND U4002 ( .A(n443), .B(n4531), .Z(n4530) );
  XOR U4003 ( .A(n4532), .B(n4529), .Z(n4531) );
  XNOR U4004 ( .A(n2711), .B(n4525), .Z(n4527) );
  XOR U4005 ( .A(n4533), .B(n4534), .Z(n2711) );
  AND U4006 ( .A(n440), .B(n4535), .Z(n4534) );
  XOR U4007 ( .A(n4536), .B(n4533), .Z(n4535) );
  XOR U4008 ( .A(n4537), .B(n4538), .Z(n4525) );
  AND U4009 ( .A(n4539), .B(n4540), .Z(n4538) );
  XOR U4010 ( .A(n4537), .B(n2726), .Z(n4540) );
  XOR U4011 ( .A(n4541), .B(n4542), .Z(n2726) );
  AND U4012 ( .A(n443), .B(n4543), .Z(n4542) );
  XOR U4013 ( .A(n4544), .B(n4541), .Z(n4543) );
  XNOR U4014 ( .A(n2723), .B(n4537), .Z(n4539) );
  XOR U4015 ( .A(n4545), .B(n4546), .Z(n2723) );
  AND U4016 ( .A(n440), .B(n4547), .Z(n4546) );
  XOR U4017 ( .A(n4548), .B(n4545), .Z(n4547) );
  XOR U4018 ( .A(n4549), .B(n4550), .Z(n4537) );
  AND U4019 ( .A(n4551), .B(n4552), .Z(n4550) );
  XOR U4020 ( .A(n4549), .B(n2738), .Z(n4552) );
  XOR U4021 ( .A(n4553), .B(n4554), .Z(n2738) );
  AND U4022 ( .A(n443), .B(n4555), .Z(n4554) );
  XOR U4023 ( .A(n4556), .B(n4553), .Z(n4555) );
  XNOR U4024 ( .A(n2735), .B(n4549), .Z(n4551) );
  XOR U4025 ( .A(n4557), .B(n4558), .Z(n2735) );
  AND U4026 ( .A(n440), .B(n4559), .Z(n4558) );
  XOR U4027 ( .A(n4560), .B(n4557), .Z(n4559) );
  XOR U4028 ( .A(n4561), .B(n4562), .Z(n4549) );
  AND U4029 ( .A(n4563), .B(n4564), .Z(n4562) );
  XOR U4030 ( .A(n4561), .B(n2750), .Z(n4564) );
  XOR U4031 ( .A(n4565), .B(n4566), .Z(n2750) );
  AND U4032 ( .A(n443), .B(n4567), .Z(n4566) );
  XOR U4033 ( .A(n4568), .B(n4565), .Z(n4567) );
  XNOR U4034 ( .A(n2747), .B(n4561), .Z(n4563) );
  XOR U4035 ( .A(n4569), .B(n4570), .Z(n2747) );
  AND U4036 ( .A(n440), .B(n4571), .Z(n4570) );
  XOR U4037 ( .A(n4572), .B(n4569), .Z(n4571) );
  XOR U4038 ( .A(n4573), .B(n4574), .Z(n4561) );
  AND U4039 ( .A(n4575), .B(n4576), .Z(n4574) );
  XOR U4040 ( .A(n4573), .B(n2762), .Z(n4576) );
  XOR U4041 ( .A(n4577), .B(n4578), .Z(n2762) );
  AND U4042 ( .A(n443), .B(n4579), .Z(n4578) );
  XOR U4043 ( .A(n4580), .B(n4577), .Z(n4579) );
  XNOR U4044 ( .A(n2759), .B(n4573), .Z(n4575) );
  XOR U4045 ( .A(n4581), .B(n4582), .Z(n2759) );
  AND U4046 ( .A(n440), .B(n4583), .Z(n4582) );
  XOR U4047 ( .A(n4584), .B(n4581), .Z(n4583) );
  XOR U4048 ( .A(n4585), .B(n4586), .Z(n4573) );
  AND U4049 ( .A(n4587), .B(n4588), .Z(n4586) );
  XOR U4050 ( .A(n4585), .B(n2774), .Z(n4588) );
  XOR U4051 ( .A(n4589), .B(n4590), .Z(n2774) );
  AND U4052 ( .A(n443), .B(n4591), .Z(n4590) );
  XOR U4053 ( .A(n4592), .B(n4589), .Z(n4591) );
  XNOR U4054 ( .A(n2771), .B(n4585), .Z(n4587) );
  XOR U4055 ( .A(n4593), .B(n4594), .Z(n2771) );
  AND U4056 ( .A(n440), .B(n4595), .Z(n4594) );
  XOR U4057 ( .A(n4596), .B(n4593), .Z(n4595) );
  XOR U4058 ( .A(n4597), .B(n4598), .Z(n4585) );
  AND U4059 ( .A(n4599), .B(n4600), .Z(n4598) );
  XOR U4060 ( .A(n4597), .B(n2786), .Z(n4600) );
  XOR U4061 ( .A(n4601), .B(n4602), .Z(n2786) );
  AND U4062 ( .A(n443), .B(n4603), .Z(n4602) );
  XOR U4063 ( .A(n4604), .B(n4601), .Z(n4603) );
  XNOR U4064 ( .A(n2783), .B(n4597), .Z(n4599) );
  XOR U4065 ( .A(n4605), .B(n4606), .Z(n2783) );
  AND U4066 ( .A(n440), .B(n4607), .Z(n4606) );
  XOR U4067 ( .A(n4608), .B(n4605), .Z(n4607) );
  XOR U4068 ( .A(n4609), .B(n4610), .Z(n4597) );
  AND U4069 ( .A(n4611), .B(n4612), .Z(n4610) );
  XOR U4070 ( .A(n4609), .B(n2798), .Z(n4612) );
  XOR U4071 ( .A(n4613), .B(n4614), .Z(n2798) );
  AND U4072 ( .A(n443), .B(n4615), .Z(n4614) );
  XOR U4073 ( .A(n4616), .B(n4613), .Z(n4615) );
  XNOR U4074 ( .A(n2795), .B(n4609), .Z(n4611) );
  XOR U4075 ( .A(n4617), .B(n4618), .Z(n2795) );
  AND U4076 ( .A(n440), .B(n4619), .Z(n4618) );
  XOR U4077 ( .A(n4620), .B(n4617), .Z(n4619) );
  XOR U4078 ( .A(n4621), .B(n4622), .Z(n4609) );
  AND U4079 ( .A(n4623), .B(n4624), .Z(n4622) );
  XOR U4080 ( .A(n4621), .B(n2810), .Z(n4624) );
  XOR U4081 ( .A(n4625), .B(n4626), .Z(n2810) );
  AND U4082 ( .A(n443), .B(n4627), .Z(n4626) );
  XOR U4083 ( .A(n4628), .B(n4625), .Z(n4627) );
  XNOR U4084 ( .A(n2807), .B(n4621), .Z(n4623) );
  XOR U4085 ( .A(n4629), .B(n4630), .Z(n2807) );
  AND U4086 ( .A(n440), .B(n4631), .Z(n4630) );
  XOR U4087 ( .A(n4632), .B(n4629), .Z(n4631) );
  XOR U4088 ( .A(n4633), .B(n4634), .Z(n4621) );
  AND U4089 ( .A(n4635), .B(n4636), .Z(n4634) );
  XOR U4090 ( .A(n4633), .B(n2822), .Z(n4636) );
  XOR U4091 ( .A(n4637), .B(n4638), .Z(n2822) );
  AND U4092 ( .A(n443), .B(n4639), .Z(n4638) );
  XOR U4093 ( .A(n4640), .B(n4637), .Z(n4639) );
  XNOR U4094 ( .A(n2819), .B(n4633), .Z(n4635) );
  XOR U4095 ( .A(n4641), .B(n4642), .Z(n2819) );
  AND U4096 ( .A(n440), .B(n4643), .Z(n4642) );
  XOR U4097 ( .A(n4644), .B(n4641), .Z(n4643) );
  XOR U4098 ( .A(n4645), .B(n4646), .Z(n4633) );
  AND U4099 ( .A(n4647), .B(n4648), .Z(n4646) );
  XOR U4100 ( .A(n4645), .B(n2834), .Z(n4648) );
  XOR U4101 ( .A(n4649), .B(n4650), .Z(n2834) );
  AND U4102 ( .A(n443), .B(n4651), .Z(n4650) );
  XOR U4103 ( .A(n4652), .B(n4649), .Z(n4651) );
  XNOR U4104 ( .A(n2831), .B(n4645), .Z(n4647) );
  XOR U4105 ( .A(n4653), .B(n4654), .Z(n2831) );
  AND U4106 ( .A(n440), .B(n4655), .Z(n4654) );
  XOR U4107 ( .A(n4656), .B(n4653), .Z(n4655) );
  XOR U4108 ( .A(n4657), .B(n4658), .Z(n4645) );
  AND U4109 ( .A(n4659), .B(n4660), .Z(n4658) );
  XOR U4110 ( .A(n4657), .B(n2846), .Z(n4660) );
  XOR U4111 ( .A(n4661), .B(n4662), .Z(n2846) );
  AND U4112 ( .A(n443), .B(n4663), .Z(n4662) );
  XOR U4113 ( .A(n4664), .B(n4661), .Z(n4663) );
  XNOR U4114 ( .A(n2843), .B(n4657), .Z(n4659) );
  XOR U4115 ( .A(n4665), .B(n4666), .Z(n2843) );
  AND U4116 ( .A(n440), .B(n4667), .Z(n4666) );
  XOR U4117 ( .A(n4668), .B(n4665), .Z(n4667) );
  XOR U4118 ( .A(n4669), .B(n4670), .Z(n4657) );
  AND U4119 ( .A(n4671), .B(n4672), .Z(n4670) );
  XOR U4120 ( .A(n4669), .B(n2858), .Z(n4672) );
  XOR U4121 ( .A(n4673), .B(n4674), .Z(n2858) );
  AND U4122 ( .A(n443), .B(n4675), .Z(n4674) );
  XOR U4123 ( .A(n4676), .B(n4673), .Z(n4675) );
  XNOR U4124 ( .A(n2855), .B(n4669), .Z(n4671) );
  XOR U4125 ( .A(n4677), .B(n4678), .Z(n2855) );
  AND U4126 ( .A(n440), .B(n4679), .Z(n4678) );
  XOR U4127 ( .A(n4680), .B(n4677), .Z(n4679) );
  XOR U4128 ( .A(n4681), .B(n4682), .Z(n4669) );
  AND U4129 ( .A(n4683), .B(n4684), .Z(n4682) );
  XOR U4130 ( .A(n4681), .B(n2870), .Z(n4684) );
  XOR U4131 ( .A(n4685), .B(n4686), .Z(n2870) );
  AND U4132 ( .A(n443), .B(n4687), .Z(n4686) );
  XOR U4133 ( .A(n4688), .B(n4685), .Z(n4687) );
  XNOR U4134 ( .A(n2867), .B(n4681), .Z(n4683) );
  XOR U4135 ( .A(n4689), .B(n4690), .Z(n2867) );
  AND U4136 ( .A(n440), .B(n4691), .Z(n4690) );
  XOR U4137 ( .A(n4692), .B(n4689), .Z(n4691) );
  XOR U4138 ( .A(n4693), .B(n4694), .Z(n4681) );
  AND U4139 ( .A(n4695), .B(n4696), .Z(n4694) );
  XOR U4140 ( .A(n4693), .B(n2882), .Z(n4696) );
  XOR U4141 ( .A(n4697), .B(n4698), .Z(n2882) );
  AND U4142 ( .A(n443), .B(n4699), .Z(n4698) );
  XOR U4143 ( .A(n4700), .B(n4697), .Z(n4699) );
  XNOR U4144 ( .A(n2879), .B(n4693), .Z(n4695) );
  XOR U4145 ( .A(n4701), .B(n4702), .Z(n2879) );
  AND U4146 ( .A(n440), .B(n4703), .Z(n4702) );
  XOR U4147 ( .A(n4704), .B(n4701), .Z(n4703) );
  XOR U4148 ( .A(n4705), .B(n4706), .Z(n4693) );
  AND U4149 ( .A(n4707), .B(n4708), .Z(n4706) );
  XOR U4150 ( .A(n4705), .B(n2894), .Z(n4708) );
  XOR U4151 ( .A(n4709), .B(n4710), .Z(n2894) );
  AND U4152 ( .A(n443), .B(n4711), .Z(n4710) );
  XOR U4153 ( .A(n4712), .B(n4709), .Z(n4711) );
  XNOR U4154 ( .A(n2891), .B(n4705), .Z(n4707) );
  XOR U4155 ( .A(n4713), .B(n4714), .Z(n2891) );
  AND U4156 ( .A(n440), .B(n4715), .Z(n4714) );
  XOR U4157 ( .A(n4716), .B(n4713), .Z(n4715) );
  XOR U4158 ( .A(n4717), .B(n4718), .Z(n4705) );
  AND U4159 ( .A(n4719), .B(n4720), .Z(n4718) );
  XOR U4160 ( .A(n4717), .B(n2906), .Z(n4720) );
  XOR U4161 ( .A(n4721), .B(n4722), .Z(n2906) );
  AND U4162 ( .A(n443), .B(n4723), .Z(n4722) );
  XOR U4163 ( .A(n4724), .B(n4721), .Z(n4723) );
  XNOR U4164 ( .A(n2903), .B(n4717), .Z(n4719) );
  XOR U4165 ( .A(n4725), .B(n4726), .Z(n2903) );
  AND U4166 ( .A(n440), .B(n4727), .Z(n4726) );
  XOR U4167 ( .A(n4728), .B(n4725), .Z(n4727) );
  XOR U4168 ( .A(n4729), .B(n4730), .Z(n4717) );
  AND U4169 ( .A(n4731), .B(n4732), .Z(n4730) );
  XOR U4170 ( .A(n4729), .B(n2918), .Z(n4732) );
  XOR U4171 ( .A(n4733), .B(n4734), .Z(n2918) );
  AND U4172 ( .A(n443), .B(n4735), .Z(n4734) );
  XOR U4173 ( .A(n4736), .B(n4733), .Z(n4735) );
  XNOR U4174 ( .A(n2915), .B(n4729), .Z(n4731) );
  XOR U4175 ( .A(n4737), .B(n4738), .Z(n2915) );
  AND U4176 ( .A(n440), .B(n4739), .Z(n4738) );
  XOR U4177 ( .A(n4740), .B(n4737), .Z(n4739) );
  XOR U4178 ( .A(n4741), .B(n4742), .Z(n4729) );
  AND U4179 ( .A(n4743), .B(n4744), .Z(n4742) );
  XOR U4180 ( .A(n4741), .B(n2930), .Z(n4744) );
  XOR U4181 ( .A(n4745), .B(n4746), .Z(n2930) );
  AND U4182 ( .A(n443), .B(n4747), .Z(n4746) );
  XOR U4183 ( .A(n4748), .B(n4745), .Z(n4747) );
  XNOR U4184 ( .A(n2927), .B(n4741), .Z(n4743) );
  XOR U4185 ( .A(n4749), .B(n4750), .Z(n2927) );
  AND U4186 ( .A(n440), .B(n4751), .Z(n4750) );
  XOR U4187 ( .A(n4752), .B(n4749), .Z(n4751) );
  XOR U4188 ( .A(n4753), .B(n4754), .Z(n4741) );
  AND U4189 ( .A(n4755), .B(n4756), .Z(n4754) );
  XOR U4190 ( .A(n4753), .B(n2942), .Z(n4756) );
  XOR U4191 ( .A(n4757), .B(n4758), .Z(n2942) );
  AND U4192 ( .A(n443), .B(n4759), .Z(n4758) );
  XOR U4193 ( .A(n4760), .B(n4757), .Z(n4759) );
  XNOR U4194 ( .A(n2939), .B(n4753), .Z(n4755) );
  XOR U4195 ( .A(n4761), .B(n4762), .Z(n2939) );
  AND U4196 ( .A(n440), .B(n4763), .Z(n4762) );
  XOR U4197 ( .A(n4764), .B(n4761), .Z(n4763) );
  XOR U4198 ( .A(n4765), .B(n4766), .Z(n4753) );
  AND U4199 ( .A(n4767), .B(n4768), .Z(n4766) );
  XOR U4200 ( .A(n4765), .B(n2954), .Z(n4768) );
  XOR U4201 ( .A(n4769), .B(n4770), .Z(n2954) );
  AND U4202 ( .A(n443), .B(n4771), .Z(n4770) );
  XOR U4203 ( .A(n4772), .B(n4769), .Z(n4771) );
  XNOR U4204 ( .A(n2951), .B(n4765), .Z(n4767) );
  XOR U4205 ( .A(n4773), .B(n4774), .Z(n2951) );
  AND U4206 ( .A(n440), .B(n4775), .Z(n4774) );
  XOR U4207 ( .A(n4776), .B(n4773), .Z(n4775) );
  XOR U4208 ( .A(n4777), .B(n4778), .Z(n4765) );
  AND U4209 ( .A(n4779), .B(n4780), .Z(n4778) );
  XOR U4210 ( .A(n4777), .B(n2966), .Z(n4780) );
  XOR U4211 ( .A(n4781), .B(n4782), .Z(n2966) );
  AND U4212 ( .A(n443), .B(n4783), .Z(n4782) );
  XOR U4213 ( .A(n4784), .B(n4781), .Z(n4783) );
  XNOR U4214 ( .A(n2963), .B(n4777), .Z(n4779) );
  XOR U4215 ( .A(n4785), .B(n4786), .Z(n2963) );
  AND U4216 ( .A(n440), .B(n4787), .Z(n4786) );
  XOR U4217 ( .A(n4788), .B(n4785), .Z(n4787) );
  XOR U4218 ( .A(n4789), .B(n4790), .Z(n4777) );
  AND U4219 ( .A(n4791), .B(n4792), .Z(n4790) );
  XOR U4220 ( .A(n4789), .B(n2978), .Z(n4792) );
  XOR U4221 ( .A(n4793), .B(n4794), .Z(n2978) );
  AND U4222 ( .A(n443), .B(n4795), .Z(n4794) );
  XOR U4223 ( .A(n4796), .B(n4793), .Z(n4795) );
  XNOR U4224 ( .A(n2975), .B(n4789), .Z(n4791) );
  XOR U4225 ( .A(n4797), .B(n4798), .Z(n2975) );
  AND U4226 ( .A(n440), .B(n4799), .Z(n4798) );
  XOR U4227 ( .A(n4800), .B(n4797), .Z(n4799) );
  XOR U4228 ( .A(n4801), .B(n4802), .Z(n4789) );
  AND U4229 ( .A(n4803), .B(n4804), .Z(n4802) );
  XOR U4230 ( .A(n4801), .B(n2990), .Z(n4804) );
  XOR U4231 ( .A(n4805), .B(n4806), .Z(n2990) );
  AND U4232 ( .A(n443), .B(n4807), .Z(n4806) );
  XOR U4233 ( .A(n4808), .B(n4805), .Z(n4807) );
  XNOR U4234 ( .A(n2987), .B(n4801), .Z(n4803) );
  XOR U4235 ( .A(n4809), .B(n4810), .Z(n2987) );
  AND U4236 ( .A(n440), .B(n4811), .Z(n4810) );
  XOR U4237 ( .A(n4812), .B(n4809), .Z(n4811) );
  XOR U4238 ( .A(n4813), .B(n4814), .Z(n4801) );
  AND U4239 ( .A(n4815), .B(n4816), .Z(n4814) );
  XOR U4240 ( .A(n4813), .B(n3002), .Z(n4816) );
  XOR U4241 ( .A(n4817), .B(n4818), .Z(n3002) );
  AND U4242 ( .A(n443), .B(n4819), .Z(n4818) );
  XOR U4243 ( .A(n4820), .B(n4817), .Z(n4819) );
  XNOR U4244 ( .A(n2999), .B(n4813), .Z(n4815) );
  XOR U4245 ( .A(n4821), .B(n4822), .Z(n2999) );
  AND U4246 ( .A(n440), .B(n4823), .Z(n4822) );
  XOR U4247 ( .A(n4824), .B(n4821), .Z(n4823) );
  XOR U4248 ( .A(n4825), .B(n4826), .Z(n4813) );
  AND U4249 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4250 ( .A(n4825), .B(n3014), .Z(n4828) );
  XOR U4251 ( .A(n4829), .B(n4830), .Z(n3014) );
  AND U4252 ( .A(n443), .B(n4831), .Z(n4830) );
  XOR U4253 ( .A(n4832), .B(n4829), .Z(n4831) );
  XNOR U4254 ( .A(n3011), .B(n4825), .Z(n4827) );
  XOR U4255 ( .A(n4833), .B(n4834), .Z(n3011) );
  AND U4256 ( .A(n440), .B(n4835), .Z(n4834) );
  XOR U4257 ( .A(n4836), .B(n4833), .Z(n4835) );
  XOR U4258 ( .A(n4837), .B(n4838), .Z(n4825) );
  AND U4259 ( .A(n4839), .B(n4840), .Z(n4838) );
  XNOR U4260 ( .A(n4841), .B(n3027), .Z(n4840) );
  XOR U4261 ( .A(n4842), .B(n4843), .Z(n3027) );
  AND U4262 ( .A(n443), .B(n4844), .Z(n4843) );
  XOR U4263 ( .A(n4842), .B(n4845), .Z(n4844) );
  XNOR U4264 ( .A(n3024), .B(n4837), .Z(n4839) );
  XOR U4265 ( .A(n4846), .B(n4847), .Z(n3024) );
  AND U4266 ( .A(n440), .B(n4848), .Z(n4847) );
  XOR U4267 ( .A(n4846), .B(n4849), .Z(n4848) );
  IV U4268 ( .A(n4841), .Z(n4837) );
  AND U4269 ( .A(n4473), .B(n4476), .Z(n4841) );
  XNOR U4270 ( .A(n4850), .B(n4851), .Z(n4476) );
  AND U4271 ( .A(n443), .B(n4852), .Z(n4851) );
  XNOR U4272 ( .A(n4853), .B(n4850), .Z(n4852) );
  XOR U4273 ( .A(n4854), .B(n4855), .Z(n443) );
  AND U4274 ( .A(n4856), .B(n4857), .Z(n4855) );
  XOR U4275 ( .A(n4484), .B(n4854), .Z(n4857) );
  IV U4276 ( .A(n4858), .Z(n4484) );
  AND U4277 ( .A(p_input[7935]), .B(p_input[7903]), .Z(n4858) );
  XOR U4278 ( .A(n4854), .B(n4481), .Z(n4856) );
  AND U4279 ( .A(p_input[7839]), .B(p_input[7871]), .Z(n4481) );
  XOR U4280 ( .A(n4859), .B(n4860), .Z(n4854) );
  AND U4281 ( .A(n4861), .B(n4862), .Z(n4860) );
  XOR U4282 ( .A(n4859), .B(n4496), .Z(n4862) );
  XNOR U4283 ( .A(p_input[7902]), .B(n4863), .Z(n4496) );
  AND U4284 ( .A(n199), .B(n4864), .Z(n4863) );
  XOR U4285 ( .A(p_input[7934]), .B(p_input[7902]), .Z(n4864) );
  XNOR U4286 ( .A(n4493), .B(n4859), .Z(n4861) );
  XOR U4287 ( .A(n4865), .B(n4866), .Z(n4493) );
  AND U4288 ( .A(n197), .B(n4867), .Z(n4866) );
  XOR U4289 ( .A(p_input[7870]), .B(p_input[7838]), .Z(n4867) );
  XOR U4290 ( .A(n4868), .B(n4869), .Z(n4859) );
  AND U4291 ( .A(n4870), .B(n4871), .Z(n4869) );
  XOR U4292 ( .A(n4868), .B(n4508), .Z(n4871) );
  XNOR U4293 ( .A(p_input[7901]), .B(n4872), .Z(n4508) );
  AND U4294 ( .A(n199), .B(n4873), .Z(n4872) );
  XOR U4295 ( .A(p_input[7933]), .B(p_input[7901]), .Z(n4873) );
  XNOR U4296 ( .A(n4505), .B(n4868), .Z(n4870) );
  XOR U4297 ( .A(n4874), .B(n4875), .Z(n4505) );
  AND U4298 ( .A(n197), .B(n4876), .Z(n4875) );
  XOR U4299 ( .A(p_input[7869]), .B(p_input[7837]), .Z(n4876) );
  XOR U4300 ( .A(n4877), .B(n4878), .Z(n4868) );
  AND U4301 ( .A(n4879), .B(n4880), .Z(n4878) );
  XOR U4302 ( .A(n4877), .B(n4520), .Z(n4880) );
  XNOR U4303 ( .A(p_input[7900]), .B(n4881), .Z(n4520) );
  AND U4304 ( .A(n199), .B(n4882), .Z(n4881) );
  XOR U4305 ( .A(p_input[7932]), .B(p_input[7900]), .Z(n4882) );
  XNOR U4306 ( .A(n4517), .B(n4877), .Z(n4879) );
  XOR U4307 ( .A(n4883), .B(n4884), .Z(n4517) );
  AND U4308 ( .A(n197), .B(n4885), .Z(n4884) );
  XOR U4309 ( .A(p_input[7868]), .B(p_input[7836]), .Z(n4885) );
  XOR U4310 ( .A(n4886), .B(n4887), .Z(n4877) );
  AND U4311 ( .A(n4888), .B(n4889), .Z(n4887) );
  XOR U4312 ( .A(n4886), .B(n4532), .Z(n4889) );
  XNOR U4313 ( .A(p_input[7899]), .B(n4890), .Z(n4532) );
  AND U4314 ( .A(n199), .B(n4891), .Z(n4890) );
  XOR U4315 ( .A(p_input[7931]), .B(p_input[7899]), .Z(n4891) );
  XNOR U4316 ( .A(n4529), .B(n4886), .Z(n4888) );
  XOR U4317 ( .A(n4892), .B(n4893), .Z(n4529) );
  AND U4318 ( .A(n197), .B(n4894), .Z(n4893) );
  XOR U4319 ( .A(p_input[7867]), .B(p_input[7835]), .Z(n4894) );
  XOR U4320 ( .A(n4895), .B(n4896), .Z(n4886) );
  AND U4321 ( .A(n4897), .B(n4898), .Z(n4896) );
  XOR U4322 ( .A(n4895), .B(n4544), .Z(n4898) );
  XNOR U4323 ( .A(p_input[7898]), .B(n4899), .Z(n4544) );
  AND U4324 ( .A(n199), .B(n4900), .Z(n4899) );
  XOR U4325 ( .A(p_input[7930]), .B(p_input[7898]), .Z(n4900) );
  XNOR U4326 ( .A(n4541), .B(n4895), .Z(n4897) );
  XOR U4327 ( .A(n4901), .B(n4902), .Z(n4541) );
  AND U4328 ( .A(n197), .B(n4903), .Z(n4902) );
  XOR U4329 ( .A(p_input[7866]), .B(p_input[7834]), .Z(n4903) );
  XOR U4330 ( .A(n4904), .B(n4905), .Z(n4895) );
  AND U4331 ( .A(n4906), .B(n4907), .Z(n4905) );
  XOR U4332 ( .A(n4904), .B(n4556), .Z(n4907) );
  XNOR U4333 ( .A(p_input[7897]), .B(n4908), .Z(n4556) );
  AND U4334 ( .A(n199), .B(n4909), .Z(n4908) );
  XOR U4335 ( .A(p_input[7929]), .B(p_input[7897]), .Z(n4909) );
  XNOR U4336 ( .A(n4553), .B(n4904), .Z(n4906) );
  XOR U4337 ( .A(n4910), .B(n4911), .Z(n4553) );
  AND U4338 ( .A(n197), .B(n4912), .Z(n4911) );
  XOR U4339 ( .A(p_input[7865]), .B(p_input[7833]), .Z(n4912) );
  XOR U4340 ( .A(n4913), .B(n4914), .Z(n4904) );
  AND U4341 ( .A(n4915), .B(n4916), .Z(n4914) );
  XOR U4342 ( .A(n4913), .B(n4568), .Z(n4916) );
  XNOR U4343 ( .A(p_input[7896]), .B(n4917), .Z(n4568) );
  AND U4344 ( .A(n199), .B(n4918), .Z(n4917) );
  XOR U4345 ( .A(p_input[7928]), .B(p_input[7896]), .Z(n4918) );
  XNOR U4346 ( .A(n4565), .B(n4913), .Z(n4915) );
  XOR U4347 ( .A(n4919), .B(n4920), .Z(n4565) );
  AND U4348 ( .A(n197), .B(n4921), .Z(n4920) );
  XOR U4349 ( .A(p_input[7864]), .B(p_input[7832]), .Z(n4921) );
  XOR U4350 ( .A(n4922), .B(n4923), .Z(n4913) );
  AND U4351 ( .A(n4924), .B(n4925), .Z(n4923) );
  XOR U4352 ( .A(n4922), .B(n4580), .Z(n4925) );
  XNOR U4353 ( .A(p_input[7895]), .B(n4926), .Z(n4580) );
  AND U4354 ( .A(n199), .B(n4927), .Z(n4926) );
  XOR U4355 ( .A(p_input[7927]), .B(p_input[7895]), .Z(n4927) );
  XNOR U4356 ( .A(n4577), .B(n4922), .Z(n4924) );
  XOR U4357 ( .A(n4928), .B(n4929), .Z(n4577) );
  AND U4358 ( .A(n197), .B(n4930), .Z(n4929) );
  XOR U4359 ( .A(p_input[7863]), .B(p_input[7831]), .Z(n4930) );
  XOR U4360 ( .A(n4931), .B(n4932), .Z(n4922) );
  AND U4361 ( .A(n4933), .B(n4934), .Z(n4932) );
  XOR U4362 ( .A(n4931), .B(n4592), .Z(n4934) );
  XNOR U4363 ( .A(p_input[7894]), .B(n4935), .Z(n4592) );
  AND U4364 ( .A(n199), .B(n4936), .Z(n4935) );
  XOR U4365 ( .A(p_input[7926]), .B(p_input[7894]), .Z(n4936) );
  XNOR U4366 ( .A(n4589), .B(n4931), .Z(n4933) );
  XOR U4367 ( .A(n4937), .B(n4938), .Z(n4589) );
  AND U4368 ( .A(n197), .B(n4939), .Z(n4938) );
  XOR U4369 ( .A(p_input[7862]), .B(p_input[7830]), .Z(n4939) );
  XOR U4370 ( .A(n4940), .B(n4941), .Z(n4931) );
  AND U4371 ( .A(n4942), .B(n4943), .Z(n4941) );
  XOR U4372 ( .A(n4940), .B(n4604), .Z(n4943) );
  XNOR U4373 ( .A(p_input[7893]), .B(n4944), .Z(n4604) );
  AND U4374 ( .A(n199), .B(n4945), .Z(n4944) );
  XOR U4375 ( .A(p_input[7925]), .B(p_input[7893]), .Z(n4945) );
  XNOR U4376 ( .A(n4601), .B(n4940), .Z(n4942) );
  XOR U4377 ( .A(n4946), .B(n4947), .Z(n4601) );
  AND U4378 ( .A(n197), .B(n4948), .Z(n4947) );
  XOR U4379 ( .A(p_input[7861]), .B(p_input[7829]), .Z(n4948) );
  XOR U4380 ( .A(n4949), .B(n4950), .Z(n4940) );
  AND U4381 ( .A(n4951), .B(n4952), .Z(n4950) );
  XOR U4382 ( .A(n4949), .B(n4616), .Z(n4952) );
  XNOR U4383 ( .A(p_input[7892]), .B(n4953), .Z(n4616) );
  AND U4384 ( .A(n199), .B(n4954), .Z(n4953) );
  XOR U4385 ( .A(p_input[7924]), .B(p_input[7892]), .Z(n4954) );
  XNOR U4386 ( .A(n4613), .B(n4949), .Z(n4951) );
  XOR U4387 ( .A(n4955), .B(n4956), .Z(n4613) );
  AND U4388 ( .A(n197), .B(n4957), .Z(n4956) );
  XOR U4389 ( .A(p_input[7860]), .B(p_input[7828]), .Z(n4957) );
  XOR U4390 ( .A(n4958), .B(n4959), .Z(n4949) );
  AND U4391 ( .A(n4960), .B(n4961), .Z(n4959) );
  XOR U4392 ( .A(n4958), .B(n4628), .Z(n4961) );
  XNOR U4393 ( .A(p_input[7891]), .B(n4962), .Z(n4628) );
  AND U4394 ( .A(n199), .B(n4963), .Z(n4962) );
  XOR U4395 ( .A(p_input[7923]), .B(p_input[7891]), .Z(n4963) );
  XNOR U4396 ( .A(n4625), .B(n4958), .Z(n4960) );
  XOR U4397 ( .A(n4964), .B(n4965), .Z(n4625) );
  AND U4398 ( .A(n197), .B(n4966), .Z(n4965) );
  XOR U4399 ( .A(p_input[7859]), .B(p_input[7827]), .Z(n4966) );
  XOR U4400 ( .A(n4967), .B(n4968), .Z(n4958) );
  AND U4401 ( .A(n4969), .B(n4970), .Z(n4968) );
  XOR U4402 ( .A(n4967), .B(n4640), .Z(n4970) );
  XNOR U4403 ( .A(p_input[7890]), .B(n4971), .Z(n4640) );
  AND U4404 ( .A(n199), .B(n4972), .Z(n4971) );
  XOR U4405 ( .A(p_input[7922]), .B(p_input[7890]), .Z(n4972) );
  XNOR U4406 ( .A(n4637), .B(n4967), .Z(n4969) );
  XOR U4407 ( .A(n4973), .B(n4974), .Z(n4637) );
  AND U4408 ( .A(n197), .B(n4975), .Z(n4974) );
  XOR U4409 ( .A(p_input[7858]), .B(p_input[7826]), .Z(n4975) );
  XOR U4410 ( .A(n4976), .B(n4977), .Z(n4967) );
  AND U4411 ( .A(n4978), .B(n4979), .Z(n4977) );
  XOR U4412 ( .A(n4976), .B(n4652), .Z(n4979) );
  XNOR U4413 ( .A(p_input[7889]), .B(n4980), .Z(n4652) );
  AND U4414 ( .A(n199), .B(n4981), .Z(n4980) );
  XOR U4415 ( .A(p_input[7921]), .B(p_input[7889]), .Z(n4981) );
  XNOR U4416 ( .A(n4649), .B(n4976), .Z(n4978) );
  XOR U4417 ( .A(n4982), .B(n4983), .Z(n4649) );
  AND U4418 ( .A(n197), .B(n4984), .Z(n4983) );
  XOR U4419 ( .A(p_input[7857]), .B(p_input[7825]), .Z(n4984) );
  XOR U4420 ( .A(n4985), .B(n4986), .Z(n4976) );
  AND U4421 ( .A(n4987), .B(n4988), .Z(n4986) );
  XOR U4422 ( .A(n4985), .B(n4664), .Z(n4988) );
  XNOR U4423 ( .A(p_input[7888]), .B(n4989), .Z(n4664) );
  AND U4424 ( .A(n199), .B(n4990), .Z(n4989) );
  XOR U4425 ( .A(p_input[7920]), .B(p_input[7888]), .Z(n4990) );
  XNOR U4426 ( .A(n4661), .B(n4985), .Z(n4987) );
  XOR U4427 ( .A(n4991), .B(n4992), .Z(n4661) );
  AND U4428 ( .A(n197), .B(n4993), .Z(n4992) );
  XOR U4429 ( .A(p_input[7856]), .B(p_input[7824]), .Z(n4993) );
  XOR U4430 ( .A(n4994), .B(n4995), .Z(n4985) );
  AND U4431 ( .A(n4996), .B(n4997), .Z(n4995) );
  XOR U4432 ( .A(n4994), .B(n4676), .Z(n4997) );
  XNOR U4433 ( .A(p_input[7887]), .B(n4998), .Z(n4676) );
  AND U4434 ( .A(n199), .B(n4999), .Z(n4998) );
  XOR U4435 ( .A(p_input[7919]), .B(p_input[7887]), .Z(n4999) );
  XNOR U4436 ( .A(n4673), .B(n4994), .Z(n4996) );
  XOR U4437 ( .A(n5000), .B(n5001), .Z(n4673) );
  AND U4438 ( .A(n197), .B(n5002), .Z(n5001) );
  XOR U4439 ( .A(p_input[7855]), .B(p_input[7823]), .Z(n5002) );
  XOR U4440 ( .A(n5003), .B(n5004), .Z(n4994) );
  AND U4441 ( .A(n5005), .B(n5006), .Z(n5004) );
  XOR U4442 ( .A(n5003), .B(n4688), .Z(n5006) );
  XNOR U4443 ( .A(p_input[7886]), .B(n5007), .Z(n4688) );
  AND U4444 ( .A(n199), .B(n5008), .Z(n5007) );
  XOR U4445 ( .A(p_input[7918]), .B(p_input[7886]), .Z(n5008) );
  XNOR U4446 ( .A(n4685), .B(n5003), .Z(n5005) );
  XOR U4447 ( .A(n5009), .B(n5010), .Z(n4685) );
  AND U4448 ( .A(n197), .B(n5011), .Z(n5010) );
  XOR U4449 ( .A(p_input[7854]), .B(p_input[7822]), .Z(n5011) );
  XOR U4450 ( .A(n5012), .B(n5013), .Z(n5003) );
  AND U4451 ( .A(n5014), .B(n5015), .Z(n5013) );
  XOR U4452 ( .A(n5012), .B(n4700), .Z(n5015) );
  XNOR U4453 ( .A(p_input[7885]), .B(n5016), .Z(n4700) );
  AND U4454 ( .A(n199), .B(n5017), .Z(n5016) );
  XOR U4455 ( .A(p_input[7917]), .B(p_input[7885]), .Z(n5017) );
  XNOR U4456 ( .A(n4697), .B(n5012), .Z(n5014) );
  XOR U4457 ( .A(n5018), .B(n5019), .Z(n4697) );
  AND U4458 ( .A(n197), .B(n5020), .Z(n5019) );
  XOR U4459 ( .A(p_input[7853]), .B(p_input[7821]), .Z(n5020) );
  XOR U4460 ( .A(n5021), .B(n5022), .Z(n5012) );
  AND U4461 ( .A(n5023), .B(n5024), .Z(n5022) );
  XOR U4462 ( .A(n5021), .B(n4712), .Z(n5024) );
  XNOR U4463 ( .A(p_input[7884]), .B(n5025), .Z(n4712) );
  AND U4464 ( .A(n199), .B(n5026), .Z(n5025) );
  XOR U4465 ( .A(p_input[7916]), .B(p_input[7884]), .Z(n5026) );
  XNOR U4466 ( .A(n4709), .B(n5021), .Z(n5023) );
  XOR U4467 ( .A(n5027), .B(n5028), .Z(n4709) );
  AND U4468 ( .A(n197), .B(n5029), .Z(n5028) );
  XOR U4469 ( .A(p_input[7852]), .B(p_input[7820]), .Z(n5029) );
  XOR U4470 ( .A(n5030), .B(n5031), .Z(n5021) );
  AND U4471 ( .A(n5032), .B(n5033), .Z(n5031) );
  XOR U4472 ( .A(n5030), .B(n4724), .Z(n5033) );
  XNOR U4473 ( .A(p_input[7883]), .B(n5034), .Z(n4724) );
  AND U4474 ( .A(n199), .B(n5035), .Z(n5034) );
  XOR U4475 ( .A(p_input[7915]), .B(p_input[7883]), .Z(n5035) );
  XNOR U4476 ( .A(n4721), .B(n5030), .Z(n5032) );
  XOR U4477 ( .A(n5036), .B(n5037), .Z(n4721) );
  AND U4478 ( .A(n197), .B(n5038), .Z(n5037) );
  XOR U4479 ( .A(p_input[7851]), .B(p_input[7819]), .Z(n5038) );
  XOR U4480 ( .A(n5039), .B(n5040), .Z(n5030) );
  AND U4481 ( .A(n5041), .B(n5042), .Z(n5040) );
  XOR U4482 ( .A(n5039), .B(n4736), .Z(n5042) );
  XNOR U4483 ( .A(p_input[7882]), .B(n5043), .Z(n4736) );
  AND U4484 ( .A(n199), .B(n5044), .Z(n5043) );
  XOR U4485 ( .A(p_input[7914]), .B(p_input[7882]), .Z(n5044) );
  XNOR U4486 ( .A(n4733), .B(n5039), .Z(n5041) );
  XOR U4487 ( .A(n5045), .B(n5046), .Z(n4733) );
  AND U4488 ( .A(n197), .B(n5047), .Z(n5046) );
  XOR U4489 ( .A(p_input[7850]), .B(p_input[7818]), .Z(n5047) );
  XOR U4490 ( .A(n5048), .B(n5049), .Z(n5039) );
  AND U4491 ( .A(n5050), .B(n5051), .Z(n5049) );
  XOR U4492 ( .A(n5048), .B(n4748), .Z(n5051) );
  XNOR U4493 ( .A(p_input[7881]), .B(n5052), .Z(n4748) );
  AND U4494 ( .A(n199), .B(n5053), .Z(n5052) );
  XOR U4495 ( .A(p_input[7913]), .B(p_input[7881]), .Z(n5053) );
  XNOR U4496 ( .A(n4745), .B(n5048), .Z(n5050) );
  XOR U4497 ( .A(n5054), .B(n5055), .Z(n4745) );
  AND U4498 ( .A(n197), .B(n5056), .Z(n5055) );
  XOR U4499 ( .A(p_input[7849]), .B(p_input[7817]), .Z(n5056) );
  XOR U4500 ( .A(n5057), .B(n5058), .Z(n5048) );
  AND U4501 ( .A(n5059), .B(n5060), .Z(n5058) );
  XOR U4502 ( .A(n5057), .B(n4760), .Z(n5060) );
  XNOR U4503 ( .A(p_input[7880]), .B(n5061), .Z(n4760) );
  AND U4504 ( .A(n199), .B(n5062), .Z(n5061) );
  XOR U4505 ( .A(p_input[7912]), .B(p_input[7880]), .Z(n5062) );
  XNOR U4506 ( .A(n4757), .B(n5057), .Z(n5059) );
  XOR U4507 ( .A(n5063), .B(n5064), .Z(n4757) );
  AND U4508 ( .A(n197), .B(n5065), .Z(n5064) );
  XOR U4509 ( .A(p_input[7848]), .B(p_input[7816]), .Z(n5065) );
  XOR U4510 ( .A(n5066), .B(n5067), .Z(n5057) );
  AND U4511 ( .A(n5068), .B(n5069), .Z(n5067) );
  XOR U4512 ( .A(n5066), .B(n4772), .Z(n5069) );
  XNOR U4513 ( .A(p_input[7879]), .B(n5070), .Z(n4772) );
  AND U4514 ( .A(n199), .B(n5071), .Z(n5070) );
  XOR U4515 ( .A(p_input[7911]), .B(p_input[7879]), .Z(n5071) );
  XNOR U4516 ( .A(n4769), .B(n5066), .Z(n5068) );
  XOR U4517 ( .A(n5072), .B(n5073), .Z(n4769) );
  AND U4518 ( .A(n197), .B(n5074), .Z(n5073) );
  XOR U4519 ( .A(p_input[7847]), .B(p_input[7815]), .Z(n5074) );
  XOR U4520 ( .A(n5075), .B(n5076), .Z(n5066) );
  AND U4521 ( .A(n5077), .B(n5078), .Z(n5076) );
  XOR U4522 ( .A(n5075), .B(n4784), .Z(n5078) );
  XNOR U4523 ( .A(p_input[7878]), .B(n5079), .Z(n4784) );
  AND U4524 ( .A(n199), .B(n5080), .Z(n5079) );
  XOR U4525 ( .A(p_input[7910]), .B(p_input[7878]), .Z(n5080) );
  XNOR U4526 ( .A(n4781), .B(n5075), .Z(n5077) );
  XOR U4527 ( .A(n5081), .B(n5082), .Z(n4781) );
  AND U4528 ( .A(n197), .B(n5083), .Z(n5082) );
  XOR U4529 ( .A(p_input[7846]), .B(p_input[7814]), .Z(n5083) );
  XOR U4530 ( .A(n5084), .B(n5085), .Z(n5075) );
  AND U4531 ( .A(n5086), .B(n5087), .Z(n5085) );
  XOR U4532 ( .A(n5084), .B(n4796), .Z(n5087) );
  XNOR U4533 ( .A(p_input[7877]), .B(n5088), .Z(n4796) );
  AND U4534 ( .A(n199), .B(n5089), .Z(n5088) );
  XOR U4535 ( .A(p_input[7909]), .B(p_input[7877]), .Z(n5089) );
  XNOR U4536 ( .A(n4793), .B(n5084), .Z(n5086) );
  XOR U4537 ( .A(n5090), .B(n5091), .Z(n4793) );
  AND U4538 ( .A(n197), .B(n5092), .Z(n5091) );
  XOR U4539 ( .A(p_input[7845]), .B(p_input[7813]), .Z(n5092) );
  XOR U4540 ( .A(n5093), .B(n5094), .Z(n5084) );
  AND U4541 ( .A(n5095), .B(n5096), .Z(n5094) );
  XOR U4542 ( .A(n5093), .B(n4808), .Z(n5096) );
  XNOR U4543 ( .A(p_input[7876]), .B(n5097), .Z(n4808) );
  AND U4544 ( .A(n199), .B(n5098), .Z(n5097) );
  XOR U4545 ( .A(p_input[7908]), .B(p_input[7876]), .Z(n5098) );
  XNOR U4546 ( .A(n4805), .B(n5093), .Z(n5095) );
  XOR U4547 ( .A(n5099), .B(n5100), .Z(n4805) );
  AND U4548 ( .A(n197), .B(n5101), .Z(n5100) );
  XOR U4549 ( .A(p_input[7844]), .B(p_input[7812]), .Z(n5101) );
  XOR U4550 ( .A(n5102), .B(n5103), .Z(n5093) );
  AND U4551 ( .A(n5104), .B(n5105), .Z(n5103) );
  XOR U4552 ( .A(n5102), .B(n4820), .Z(n5105) );
  XNOR U4553 ( .A(p_input[7875]), .B(n5106), .Z(n4820) );
  AND U4554 ( .A(n199), .B(n5107), .Z(n5106) );
  XOR U4555 ( .A(p_input[7907]), .B(p_input[7875]), .Z(n5107) );
  XNOR U4556 ( .A(n4817), .B(n5102), .Z(n5104) );
  XOR U4557 ( .A(n5108), .B(n5109), .Z(n4817) );
  AND U4558 ( .A(n197), .B(n5110), .Z(n5109) );
  XOR U4559 ( .A(p_input[7843]), .B(p_input[7811]), .Z(n5110) );
  XOR U4560 ( .A(n5111), .B(n5112), .Z(n5102) );
  AND U4561 ( .A(n5113), .B(n5114), .Z(n5112) );
  XOR U4562 ( .A(n5111), .B(n4832), .Z(n5114) );
  XNOR U4563 ( .A(p_input[7874]), .B(n5115), .Z(n4832) );
  AND U4564 ( .A(n199), .B(n5116), .Z(n5115) );
  XOR U4565 ( .A(p_input[7906]), .B(p_input[7874]), .Z(n5116) );
  XNOR U4566 ( .A(n4829), .B(n5111), .Z(n5113) );
  XOR U4567 ( .A(n5117), .B(n5118), .Z(n4829) );
  AND U4568 ( .A(n197), .B(n5119), .Z(n5118) );
  XOR U4569 ( .A(p_input[7842]), .B(p_input[7810]), .Z(n5119) );
  XOR U4570 ( .A(n5120), .B(n5121), .Z(n5111) );
  AND U4571 ( .A(n5122), .B(n5123), .Z(n5121) );
  XNOR U4572 ( .A(n5124), .B(n4845), .Z(n5123) );
  XNOR U4573 ( .A(p_input[7873]), .B(n5125), .Z(n4845) );
  AND U4574 ( .A(n199), .B(n5126), .Z(n5125) );
  XNOR U4575 ( .A(p_input[7905]), .B(n5127), .Z(n5126) );
  IV U4576 ( .A(p_input[7873]), .Z(n5127) );
  XNOR U4577 ( .A(n4842), .B(n5120), .Z(n5122) );
  XNOR U4578 ( .A(p_input[7809]), .B(n5128), .Z(n4842) );
  AND U4579 ( .A(n197), .B(n5129), .Z(n5128) );
  XOR U4580 ( .A(p_input[7841]), .B(p_input[7809]), .Z(n5129) );
  IV U4581 ( .A(n5124), .Z(n5120) );
  AND U4582 ( .A(n4850), .B(n4853), .Z(n5124) );
  XOR U4583 ( .A(p_input[7872]), .B(n5130), .Z(n4853) );
  AND U4584 ( .A(n199), .B(n5131), .Z(n5130) );
  XOR U4585 ( .A(p_input[7904]), .B(p_input[7872]), .Z(n5131) );
  XOR U4586 ( .A(n5132), .B(n5133), .Z(n199) );
  AND U4587 ( .A(n5134), .B(n5135), .Z(n5133) );
  XNOR U4588 ( .A(p_input[7935]), .B(n5132), .Z(n5135) );
  XOR U4589 ( .A(n5132), .B(p_input[7903]), .Z(n5134) );
  XOR U4590 ( .A(n5136), .B(n5137), .Z(n5132) );
  AND U4591 ( .A(n5138), .B(n5139), .Z(n5137) );
  XNOR U4592 ( .A(p_input[7934]), .B(n5136), .Z(n5139) );
  XOR U4593 ( .A(n5136), .B(p_input[7902]), .Z(n5138) );
  XOR U4594 ( .A(n5140), .B(n5141), .Z(n5136) );
  AND U4595 ( .A(n5142), .B(n5143), .Z(n5141) );
  XNOR U4596 ( .A(p_input[7933]), .B(n5140), .Z(n5143) );
  XOR U4597 ( .A(n5140), .B(p_input[7901]), .Z(n5142) );
  XOR U4598 ( .A(n5144), .B(n5145), .Z(n5140) );
  AND U4599 ( .A(n5146), .B(n5147), .Z(n5145) );
  XNOR U4600 ( .A(p_input[7932]), .B(n5144), .Z(n5147) );
  XOR U4601 ( .A(n5144), .B(p_input[7900]), .Z(n5146) );
  XOR U4602 ( .A(n5148), .B(n5149), .Z(n5144) );
  AND U4603 ( .A(n5150), .B(n5151), .Z(n5149) );
  XNOR U4604 ( .A(p_input[7931]), .B(n5148), .Z(n5151) );
  XOR U4605 ( .A(n5148), .B(p_input[7899]), .Z(n5150) );
  XOR U4606 ( .A(n5152), .B(n5153), .Z(n5148) );
  AND U4607 ( .A(n5154), .B(n5155), .Z(n5153) );
  XNOR U4608 ( .A(p_input[7930]), .B(n5152), .Z(n5155) );
  XOR U4609 ( .A(n5152), .B(p_input[7898]), .Z(n5154) );
  XOR U4610 ( .A(n5156), .B(n5157), .Z(n5152) );
  AND U4611 ( .A(n5158), .B(n5159), .Z(n5157) );
  XNOR U4612 ( .A(p_input[7929]), .B(n5156), .Z(n5159) );
  XOR U4613 ( .A(n5156), .B(p_input[7897]), .Z(n5158) );
  XOR U4614 ( .A(n5160), .B(n5161), .Z(n5156) );
  AND U4615 ( .A(n5162), .B(n5163), .Z(n5161) );
  XNOR U4616 ( .A(p_input[7928]), .B(n5160), .Z(n5163) );
  XOR U4617 ( .A(n5160), .B(p_input[7896]), .Z(n5162) );
  XOR U4618 ( .A(n5164), .B(n5165), .Z(n5160) );
  AND U4619 ( .A(n5166), .B(n5167), .Z(n5165) );
  XNOR U4620 ( .A(p_input[7927]), .B(n5164), .Z(n5167) );
  XOR U4621 ( .A(n5164), .B(p_input[7895]), .Z(n5166) );
  XOR U4622 ( .A(n5168), .B(n5169), .Z(n5164) );
  AND U4623 ( .A(n5170), .B(n5171), .Z(n5169) );
  XNOR U4624 ( .A(p_input[7926]), .B(n5168), .Z(n5171) );
  XOR U4625 ( .A(n5168), .B(p_input[7894]), .Z(n5170) );
  XOR U4626 ( .A(n5172), .B(n5173), .Z(n5168) );
  AND U4627 ( .A(n5174), .B(n5175), .Z(n5173) );
  XNOR U4628 ( .A(p_input[7925]), .B(n5172), .Z(n5175) );
  XOR U4629 ( .A(n5172), .B(p_input[7893]), .Z(n5174) );
  XOR U4630 ( .A(n5176), .B(n5177), .Z(n5172) );
  AND U4631 ( .A(n5178), .B(n5179), .Z(n5177) );
  XNOR U4632 ( .A(p_input[7924]), .B(n5176), .Z(n5179) );
  XOR U4633 ( .A(n5176), .B(p_input[7892]), .Z(n5178) );
  XOR U4634 ( .A(n5180), .B(n5181), .Z(n5176) );
  AND U4635 ( .A(n5182), .B(n5183), .Z(n5181) );
  XNOR U4636 ( .A(p_input[7923]), .B(n5180), .Z(n5183) );
  XOR U4637 ( .A(n5180), .B(p_input[7891]), .Z(n5182) );
  XOR U4638 ( .A(n5184), .B(n5185), .Z(n5180) );
  AND U4639 ( .A(n5186), .B(n5187), .Z(n5185) );
  XNOR U4640 ( .A(p_input[7922]), .B(n5184), .Z(n5187) );
  XOR U4641 ( .A(n5184), .B(p_input[7890]), .Z(n5186) );
  XOR U4642 ( .A(n5188), .B(n5189), .Z(n5184) );
  AND U4643 ( .A(n5190), .B(n5191), .Z(n5189) );
  XNOR U4644 ( .A(p_input[7921]), .B(n5188), .Z(n5191) );
  XOR U4645 ( .A(n5188), .B(p_input[7889]), .Z(n5190) );
  XOR U4646 ( .A(n5192), .B(n5193), .Z(n5188) );
  AND U4647 ( .A(n5194), .B(n5195), .Z(n5193) );
  XNOR U4648 ( .A(p_input[7920]), .B(n5192), .Z(n5195) );
  XOR U4649 ( .A(n5192), .B(p_input[7888]), .Z(n5194) );
  XOR U4650 ( .A(n5196), .B(n5197), .Z(n5192) );
  AND U4651 ( .A(n5198), .B(n5199), .Z(n5197) );
  XNOR U4652 ( .A(p_input[7919]), .B(n5196), .Z(n5199) );
  XOR U4653 ( .A(n5196), .B(p_input[7887]), .Z(n5198) );
  XOR U4654 ( .A(n5200), .B(n5201), .Z(n5196) );
  AND U4655 ( .A(n5202), .B(n5203), .Z(n5201) );
  XNOR U4656 ( .A(p_input[7918]), .B(n5200), .Z(n5203) );
  XOR U4657 ( .A(n5200), .B(p_input[7886]), .Z(n5202) );
  XOR U4658 ( .A(n5204), .B(n5205), .Z(n5200) );
  AND U4659 ( .A(n5206), .B(n5207), .Z(n5205) );
  XNOR U4660 ( .A(p_input[7917]), .B(n5204), .Z(n5207) );
  XOR U4661 ( .A(n5204), .B(p_input[7885]), .Z(n5206) );
  XOR U4662 ( .A(n5208), .B(n5209), .Z(n5204) );
  AND U4663 ( .A(n5210), .B(n5211), .Z(n5209) );
  XNOR U4664 ( .A(p_input[7916]), .B(n5208), .Z(n5211) );
  XOR U4665 ( .A(n5208), .B(p_input[7884]), .Z(n5210) );
  XOR U4666 ( .A(n5212), .B(n5213), .Z(n5208) );
  AND U4667 ( .A(n5214), .B(n5215), .Z(n5213) );
  XNOR U4668 ( .A(p_input[7915]), .B(n5212), .Z(n5215) );
  XOR U4669 ( .A(n5212), .B(p_input[7883]), .Z(n5214) );
  XOR U4670 ( .A(n5216), .B(n5217), .Z(n5212) );
  AND U4671 ( .A(n5218), .B(n5219), .Z(n5217) );
  XNOR U4672 ( .A(p_input[7914]), .B(n5216), .Z(n5219) );
  XOR U4673 ( .A(n5216), .B(p_input[7882]), .Z(n5218) );
  XOR U4674 ( .A(n5220), .B(n5221), .Z(n5216) );
  AND U4675 ( .A(n5222), .B(n5223), .Z(n5221) );
  XNOR U4676 ( .A(p_input[7913]), .B(n5220), .Z(n5223) );
  XOR U4677 ( .A(n5220), .B(p_input[7881]), .Z(n5222) );
  XOR U4678 ( .A(n5224), .B(n5225), .Z(n5220) );
  AND U4679 ( .A(n5226), .B(n5227), .Z(n5225) );
  XNOR U4680 ( .A(p_input[7912]), .B(n5224), .Z(n5227) );
  XOR U4681 ( .A(n5224), .B(p_input[7880]), .Z(n5226) );
  XOR U4682 ( .A(n5228), .B(n5229), .Z(n5224) );
  AND U4683 ( .A(n5230), .B(n5231), .Z(n5229) );
  XNOR U4684 ( .A(p_input[7911]), .B(n5228), .Z(n5231) );
  XOR U4685 ( .A(n5228), .B(p_input[7879]), .Z(n5230) );
  XOR U4686 ( .A(n5232), .B(n5233), .Z(n5228) );
  AND U4687 ( .A(n5234), .B(n5235), .Z(n5233) );
  XNOR U4688 ( .A(p_input[7910]), .B(n5232), .Z(n5235) );
  XOR U4689 ( .A(n5232), .B(p_input[7878]), .Z(n5234) );
  XOR U4690 ( .A(n5236), .B(n5237), .Z(n5232) );
  AND U4691 ( .A(n5238), .B(n5239), .Z(n5237) );
  XNOR U4692 ( .A(p_input[7909]), .B(n5236), .Z(n5239) );
  XOR U4693 ( .A(n5236), .B(p_input[7877]), .Z(n5238) );
  XOR U4694 ( .A(n5240), .B(n5241), .Z(n5236) );
  AND U4695 ( .A(n5242), .B(n5243), .Z(n5241) );
  XNOR U4696 ( .A(p_input[7908]), .B(n5240), .Z(n5243) );
  XOR U4697 ( .A(n5240), .B(p_input[7876]), .Z(n5242) );
  XOR U4698 ( .A(n5244), .B(n5245), .Z(n5240) );
  AND U4699 ( .A(n5246), .B(n5247), .Z(n5245) );
  XNOR U4700 ( .A(p_input[7907]), .B(n5244), .Z(n5247) );
  XOR U4701 ( .A(n5244), .B(p_input[7875]), .Z(n5246) );
  XOR U4702 ( .A(n5248), .B(n5249), .Z(n5244) );
  AND U4703 ( .A(n5250), .B(n5251), .Z(n5249) );
  XNOR U4704 ( .A(p_input[7906]), .B(n5248), .Z(n5251) );
  XOR U4705 ( .A(n5248), .B(p_input[7874]), .Z(n5250) );
  XNOR U4706 ( .A(n5252), .B(n5253), .Z(n5248) );
  AND U4707 ( .A(n5254), .B(n5255), .Z(n5253) );
  XOR U4708 ( .A(p_input[7905]), .B(n5252), .Z(n5255) );
  XNOR U4709 ( .A(p_input[7873]), .B(n5252), .Z(n5254) );
  AND U4710 ( .A(p_input[7904]), .B(n5256), .Z(n5252) );
  IV U4711 ( .A(p_input[7872]), .Z(n5256) );
  XNOR U4712 ( .A(p_input[7808]), .B(n5257), .Z(n4850) );
  AND U4713 ( .A(n197), .B(n5258), .Z(n5257) );
  XOR U4714 ( .A(p_input[7840]), .B(p_input[7808]), .Z(n5258) );
  XOR U4715 ( .A(n5259), .B(n5260), .Z(n197) );
  AND U4716 ( .A(n5261), .B(n5262), .Z(n5260) );
  XNOR U4717 ( .A(p_input[7871]), .B(n5259), .Z(n5262) );
  XOR U4718 ( .A(n5259), .B(p_input[7839]), .Z(n5261) );
  XOR U4719 ( .A(n5263), .B(n5264), .Z(n5259) );
  AND U4720 ( .A(n5265), .B(n5266), .Z(n5264) );
  XNOR U4721 ( .A(p_input[7870]), .B(n5263), .Z(n5266) );
  XNOR U4722 ( .A(n5263), .B(n4865), .Z(n5265) );
  IV U4723 ( .A(p_input[7838]), .Z(n4865) );
  XOR U4724 ( .A(n5267), .B(n5268), .Z(n5263) );
  AND U4725 ( .A(n5269), .B(n5270), .Z(n5268) );
  XNOR U4726 ( .A(p_input[7869]), .B(n5267), .Z(n5270) );
  XNOR U4727 ( .A(n5267), .B(n4874), .Z(n5269) );
  IV U4728 ( .A(p_input[7837]), .Z(n4874) );
  XOR U4729 ( .A(n5271), .B(n5272), .Z(n5267) );
  AND U4730 ( .A(n5273), .B(n5274), .Z(n5272) );
  XNOR U4731 ( .A(p_input[7868]), .B(n5271), .Z(n5274) );
  XNOR U4732 ( .A(n5271), .B(n4883), .Z(n5273) );
  IV U4733 ( .A(p_input[7836]), .Z(n4883) );
  XOR U4734 ( .A(n5275), .B(n5276), .Z(n5271) );
  AND U4735 ( .A(n5277), .B(n5278), .Z(n5276) );
  XNOR U4736 ( .A(p_input[7867]), .B(n5275), .Z(n5278) );
  XNOR U4737 ( .A(n5275), .B(n4892), .Z(n5277) );
  IV U4738 ( .A(p_input[7835]), .Z(n4892) );
  XOR U4739 ( .A(n5279), .B(n5280), .Z(n5275) );
  AND U4740 ( .A(n5281), .B(n5282), .Z(n5280) );
  XNOR U4741 ( .A(p_input[7866]), .B(n5279), .Z(n5282) );
  XNOR U4742 ( .A(n5279), .B(n4901), .Z(n5281) );
  IV U4743 ( .A(p_input[7834]), .Z(n4901) );
  XOR U4744 ( .A(n5283), .B(n5284), .Z(n5279) );
  AND U4745 ( .A(n5285), .B(n5286), .Z(n5284) );
  XNOR U4746 ( .A(p_input[7865]), .B(n5283), .Z(n5286) );
  XNOR U4747 ( .A(n5283), .B(n4910), .Z(n5285) );
  IV U4748 ( .A(p_input[7833]), .Z(n4910) );
  XOR U4749 ( .A(n5287), .B(n5288), .Z(n5283) );
  AND U4750 ( .A(n5289), .B(n5290), .Z(n5288) );
  XNOR U4751 ( .A(p_input[7864]), .B(n5287), .Z(n5290) );
  XNOR U4752 ( .A(n5287), .B(n4919), .Z(n5289) );
  IV U4753 ( .A(p_input[7832]), .Z(n4919) );
  XOR U4754 ( .A(n5291), .B(n5292), .Z(n5287) );
  AND U4755 ( .A(n5293), .B(n5294), .Z(n5292) );
  XNOR U4756 ( .A(p_input[7863]), .B(n5291), .Z(n5294) );
  XNOR U4757 ( .A(n5291), .B(n4928), .Z(n5293) );
  IV U4758 ( .A(p_input[7831]), .Z(n4928) );
  XOR U4759 ( .A(n5295), .B(n5296), .Z(n5291) );
  AND U4760 ( .A(n5297), .B(n5298), .Z(n5296) );
  XNOR U4761 ( .A(p_input[7862]), .B(n5295), .Z(n5298) );
  XNOR U4762 ( .A(n5295), .B(n4937), .Z(n5297) );
  IV U4763 ( .A(p_input[7830]), .Z(n4937) );
  XOR U4764 ( .A(n5299), .B(n5300), .Z(n5295) );
  AND U4765 ( .A(n5301), .B(n5302), .Z(n5300) );
  XNOR U4766 ( .A(p_input[7861]), .B(n5299), .Z(n5302) );
  XNOR U4767 ( .A(n5299), .B(n4946), .Z(n5301) );
  IV U4768 ( .A(p_input[7829]), .Z(n4946) );
  XOR U4769 ( .A(n5303), .B(n5304), .Z(n5299) );
  AND U4770 ( .A(n5305), .B(n5306), .Z(n5304) );
  XNOR U4771 ( .A(p_input[7860]), .B(n5303), .Z(n5306) );
  XNOR U4772 ( .A(n5303), .B(n4955), .Z(n5305) );
  IV U4773 ( .A(p_input[7828]), .Z(n4955) );
  XOR U4774 ( .A(n5307), .B(n5308), .Z(n5303) );
  AND U4775 ( .A(n5309), .B(n5310), .Z(n5308) );
  XNOR U4776 ( .A(p_input[7859]), .B(n5307), .Z(n5310) );
  XNOR U4777 ( .A(n5307), .B(n4964), .Z(n5309) );
  IV U4778 ( .A(p_input[7827]), .Z(n4964) );
  XOR U4779 ( .A(n5311), .B(n5312), .Z(n5307) );
  AND U4780 ( .A(n5313), .B(n5314), .Z(n5312) );
  XNOR U4781 ( .A(p_input[7858]), .B(n5311), .Z(n5314) );
  XNOR U4782 ( .A(n5311), .B(n4973), .Z(n5313) );
  IV U4783 ( .A(p_input[7826]), .Z(n4973) );
  XOR U4784 ( .A(n5315), .B(n5316), .Z(n5311) );
  AND U4785 ( .A(n5317), .B(n5318), .Z(n5316) );
  XNOR U4786 ( .A(p_input[7857]), .B(n5315), .Z(n5318) );
  XNOR U4787 ( .A(n5315), .B(n4982), .Z(n5317) );
  IV U4788 ( .A(p_input[7825]), .Z(n4982) );
  XOR U4789 ( .A(n5319), .B(n5320), .Z(n5315) );
  AND U4790 ( .A(n5321), .B(n5322), .Z(n5320) );
  XNOR U4791 ( .A(p_input[7856]), .B(n5319), .Z(n5322) );
  XNOR U4792 ( .A(n5319), .B(n4991), .Z(n5321) );
  IV U4793 ( .A(p_input[7824]), .Z(n4991) );
  XOR U4794 ( .A(n5323), .B(n5324), .Z(n5319) );
  AND U4795 ( .A(n5325), .B(n5326), .Z(n5324) );
  XNOR U4796 ( .A(p_input[7855]), .B(n5323), .Z(n5326) );
  XNOR U4797 ( .A(n5323), .B(n5000), .Z(n5325) );
  IV U4798 ( .A(p_input[7823]), .Z(n5000) );
  XOR U4799 ( .A(n5327), .B(n5328), .Z(n5323) );
  AND U4800 ( .A(n5329), .B(n5330), .Z(n5328) );
  XNOR U4801 ( .A(p_input[7854]), .B(n5327), .Z(n5330) );
  XNOR U4802 ( .A(n5327), .B(n5009), .Z(n5329) );
  IV U4803 ( .A(p_input[7822]), .Z(n5009) );
  XOR U4804 ( .A(n5331), .B(n5332), .Z(n5327) );
  AND U4805 ( .A(n5333), .B(n5334), .Z(n5332) );
  XNOR U4806 ( .A(p_input[7853]), .B(n5331), .Z(n5334) );
  XNOR U4807 ( .A(n5331), .B(n5018), .Z(n5333) );
  IV U4808 ( .A(p_input[7821]), .Z(n5018) );
  XOR U4809 ( .A(n5335), .B(n5336), .Z(n5331) );
  AND U4810 ( .A(n5337), .B(n5338), .Z(n5336) );
  XNOR U4811 ( .A(p_input[7852]), .B(n5335), .Z(n5338) );
  XNOR U4812 ( .A(n5335), .B(n5027), .Z(n5337) );
  IV U4813 ( .A(p_input[7820]), .Z(n5027) );
  XOR U4814 ( .A(n5339), .B(n5340), .Z(n5335) );
  AND U4815 ( .A(n5341), .B(n5342), .Z(n5340) );
  XNOR U4816 ( .A(p_input[7851]), .B(n5339), .Z(n5342) );
  XNOR U4817 ( .A(n5339), .B(n5036), .Z(n5341) );
  IV U4818 ( .A(p_input[7819]), .Z(n5036) );
  XOR U4819 ( .A(n5343), .B(n5344), .Z(n5339) );
  AND U4820 ( .A(n5345), .B(n5346), .Z(n5344) );
  XNOR U4821 ( .A(p_input[7850]), .B(n5343), .Z(n5346) );
  XNOR U4822 ( .A(n5343), .B(n5045), .Z(n5345) );
  IV U4823 ( .A(p_input[7818]), .Z(n5045) );
  XOR U4824 ( .A(n5347), .B(n5348), .Z(n5343) );
  AND U4825 ( .A(n5349), .B(n5350), .Z(n5348) );
  XNOR U4826 ( .A(p_input[7849]), .B(n5347), .Z(n5350) );
  XNOR U4827 ( .A(n5347), .B(n5054), .Z(n5349) );
  IV U4828 ( .A(p_input[7817]), .Z(n5054) );
  XOR U4829 ( .A(n5351), .B(n5352), .Z(n5347) );
  AND U4830 ( .A(n5353), .B(n5354), .Z(n5352) );
  XNOR U4831 ( .A(p_input[7848]), .B(n5351), .Z(n5354) );
  XNOR U4832 ( .A(n5351), .B(n5063), .Z(n5353) );
  IV U4833 ( .A(p_input[7816]), .Z(n5063) );
  XOR U4834 ( .A(n5355), .B(n5356), .Z(n5351) );
  AND U4835 ( .A(n5357), .B(n5358), .Z(n5356) );
  XNOR U4836 ( .A(p_input[7847]), .B(n5355), .Z(n5358) );
  XNOR U4837 ( .A(n5355), .B(n5072), .Z(n5357) );
  IV U4838 ( .A(p_input[7815]), .Z(n5072) );
  XOR U4839 ( .A(n5359), .B(n5360), .Z(n5355) );
  AND U4840 ( .A(n5361), .B(n5362), .Z(n5360) );
  XNOR U4841 ( .A(p_input[7846]), .B(n5359), .Z(n5362) );
  XNOR U4842 ( .A(n5359), .B(n5081), .Z(n5361) );
  IV U4843 ( .A(p_input[7814]), .Z(n5081) );
  XOR U4844 ( .A(n5363), .B(n5364), .Z(n5359) );
  AND U4845 ( .A(n5365), .B(n5366), .Z(n5364) );
  XNOR U4846 ( .A(p_input[7845]), .B(n5363), .Z(n5366) );
  XNOR U4847 ( .A(n5363), .B(n5090), .Z(n5365) );
  IV U4848 ( .A(p_input[7813]), .Z(n5090) );
  XOR U4849 ( .A(n5367), .B(n5368), .Z(n5363) );
  AND U4850 ( .A(n5369), .B(n5370), .Z(n5368) );
  XNOR U4851 ( .A(p_input[7844]), .B(n5367), .Z(n5370) );
  XNOR U4852 ( .A(n5367), .B(n5099), .Z(n5369) );
  IV U4853 ( .A(p_input[7812]), .Z(n5099) );
  XOR U4854 ( .A(n5371), .B(n5372), .Z(n5367) );
  AND U4855 ( .A(n5373), .B(n5374), .Z(n5372) );
  XNOR U4856 ( .A(p_input[7843]), .B(n5371), .Z(n5374) );
  XNOR U4857 ( .A(n5371), .B(n5108), .Z(n5373) );
  IV U4858 ( .A(p_input[7811]), .Z(n5108) );
  XOR U4859 ( .A(n5375), .B(n5376), .Z(n5371) );
  AND U4860 ( .A(n5377), .B(n5378), .Z(n5376) );
  XNOR U4861 ( .A(p_input[7842]), .B(n5375), .Z(n5378) );
  XNOR U4862 ( .A(n5375), .B(n5117), .Z(n5377) );
  IV U4863 ( .A(p_input[7810]), .Z(n5117) );
  XNOR U4864 ( .A(n5379), .B(n5380), .Z(n5375) );
  AND U4865 ( .A(n5381), .B(n5382), .Z(n5380) );
  XOR U4866 ( .A(p_input[7841]), .B(n5379), .Z(n5382) );
  XNOR U4867 ( .A(p_input[7809]), .B(n5379), .Z(n5381) );
  AND U4868 ( .A(p_input[7840]), .B(n5383), .Z(n5379) );
  IV U4869 ( .A(p_input[7808]), .Z(n5383) );
  XOR U4870 ( .A(n5384), .B(n5385), .Z(n4473) );
  AND U4871 ( .A(n440), .B(n5386), .Z(n5385) );
  XNOR U4872 ( .A(n5387), .B(n5384), .Z(n5386) );
  XOR U4873 ( .A(n5388), .B(n5389), .Z(n440) );
  AND U4874 ( .A(n5390), .B(n5391), .Z(n5389) );
  XNOR U4875 ( .A(n4488), .B(n5388), .Z(n5391) );
  AND U4876 ( .A(p_input[7807]), .B(p_input[7775]), .Z(n4488) );
  XNOR U4877 ( .A(n5388), .B(n4485), .Z(n5390) );
  IV U4878 ( .A(n5392), .Z(n4485) );
  AND U4879 ( .A(p_input[7711]), .B(p_input[7743]), .Z(n5392) );
  XOR U4880 ( .A(n5393), .B(n5394), .Z(n5388) );
  AND U4881 ( .A(n5395), .B(n5396), .Z(n5394) );
  XOR U4882 ( .A(n5393), .B(n4500), .Z(n5396) );
  XNOR U4883 ( .A(p_input[7774]), .B(n5397), .Z(n4500) );
  AND U4884 ( .A(n203), .B(n5398), .Z(n5397) );
  XOR U4885 ( .A(p_input[7806]), .B(p_input[7774]), .Z(n5398) );
  XNOR U4886 ( .A(n4497), .B(n5393), .Z(n5395) );
  XOR U4887 ( .A(n5399), .B(n5400), .Z(n4497) );
  AND U4888 ( .A(n200), .B(n5401), .Z(n5400) );
  XOR U4889 ( .A(p_input[7742]), .B(p_input[7710]), .Z(n5401) );
  XOR U4890 ( .A(n5402), .B(n5403), .Z(n5393) );
  AND U4891 ( .A(n5404), .B(n5405), .Z(n5403) );
  XOR U4892 ( .A(n5402), .B(n4512), .Z(n5405) );
  XNOR U4893 ( .A(p_input[7773]), .B(n5406), .Z(n4512) );
  AND U4894 ( .A(n203), .B(n5407), .Z(n5406) );
  XOR U4895 ( .A(p_input[7805]), .B(p_input[7773]), .Z(n5407) );
  XNOR U4896 ( .A(n4509), .B(n5402), .Z(n5404) );
  XOR U4897 ( .A(n5408), .B(n5409), .Z(n4509) );
  AND U4898 ( .A(n200), .B(n5410), .Z(n5409) );
  XOR U4899 ( .A(p_input[7741]), .B(p_input[7709]), .Z(n5410) );
  XOR U4900 ( .A(n5411), .B(n5412), .Z(n5402) );
  AND U4901 ( .A(n5413), .B(n5414), .Z(n5412) );
  XOR U4902 ( .A(n5411), .B(n4524), .Z(n5414) );
  XNOR U4903 ( .A(p_input[7772]), .B(n5415), .Z(n4524) );
  AND U4904 ( .A(n203), .B(n5416), .Z(n5415) );
  XOR U4905 ( .A(p_input[7804]), .B(p_input[7772]), .Z(n5416) );
  XNOR U4906 ( .A(n4521), .B(n5411), .Z(n5413) );
  XOR U4907 ( .A(n5417), .B(n5418), .Z(n4521) );
  AND U4908 ( .A(n200), .B(n5419), .Z(n5418) );
  XOR U4909 ( .A(p_input[7740]), .B(p_input[7708]), .Z(n5419) );
  XOR U4910 ( .A(n5420), .B(n5421), .Z(n5411) );
  AND U4911 ( .A(n5422), .B(n5423), .Z(n5421) );
  XOR U4912 ( .A(n5420), .B(n4536), .Z(n5423) );
  XNOR U4913 ( .A(p_input[7771]), .B(n5424), .Z(n4536) );
  AND U4914 ( .A(n203), .B(n5425), .Z(n5424) );
  XOR U4915 ( .A(p_input[7803]), .B(p_input[7771]), .Z(n5425) );
  XNOR U4916 ( .A(n4533), .B(n5420), .Z(n5422) );
  XOR U4917 ( .A(n5426), .B(n5427), .Z(n4533) );
  AND U4918 ( .A(n200), .B(n5428), .Z(n5427) );
  XOR U4919 ( .A(p_input[7739]), .B(p_input[7707]), .Z(n5428) );
  XOR U4920 ( .A(n5429), .B(n5430), .Z(n5420) );
  AND U4921 ( .A(n5431), .B(n5432), .Z(n5430) );
  XOR U4922 ( .A(n5429), .B(n4548), .Z(n5432) );
  XNOR U4923 ( .A(p_input[7770]), .B(n5433), .Z(n4548) );
  AND U4924 ( .A(n203), .B(n5434), .Z(n5433) );
  XOR U4925 ( .A(p_input[7802]), .B(p_input[7770]), .Z(n5434) );
  XNOR U4926 ( .A(n4545), .B(n5429), .Z(n5431) );
  XOR U4927 ( .A(n5435), .B(n5436), .Z(n4545) );
  AND U4928 ( .A(n200), .B(n5437), .Z(n5436) );
  XOR U4929 ( .A(p_input[7738]), .B(p_input[7706]), .Z(n5437) );
  XOR U4930 ( .A(n5438), .B(n5439), .Z(n5429) );
  AND U4931 ( .A(n5440), .B(n5441), .Z(n5439) );
  XOR U4932 ( .A(n5438), .B(n4560), .Z(n5441) );
  XNOR U4933 ( .A(p_input[7769]), .B(n5442), .Z(n4560) );
  AND U4934 ( .A(n203), .B(n5443), .Z(n5442) );
  XOR U4935 ( .A(p_input[7801]), .B(p_input[7769]), .Z(n5443) );
  XNOR U4936 ( .A(n4557), .B(n5438), .Z(n5440) );
  XOR U4937 ( .A(n5444), .B(n5445), .Z(n4557) );
  AND U4938 ( .A(n200), .B(n5446), .Z(n5445) );
  XOR U4939 ( .A(p_input[7737]), .B(p_input[7705]), .Z(n5446) );
  XOR U4940 ( .A(n5447), .B(n5448), .Z(n5438) );
  AND U4941 ( .A(n5449), .B(n5450), .Z(n5448) );
  XOR U4942 ( .A(n5447), .B(n4572), .Z(n5450) );
  XNOR U4943 ( .A(p_input[7768]), .B(n5451), .Z(n4572) );
  AND U4944 ( .A(n203), .B(n5452), .Z(n5451) );
  XOR U4945 ( .A(p_input[7800]), .B(p_input[7768]), .Z(n5452) );
  XNOR U4946 ( .A(n4569), .B(n5447), .Z(n5449) );
  XOR U4947 ( .A(n5453), .B(n5454), .Z(n4569) );
  AND U4948 ( .A(n200), .B(n5455), .Z(n5454) );
  XOR U4949 ( .A(p_input[7736]), .B(p_input[7704]), .Z(n5455) );
  XOR U4950 ( .A(n5456), .B(n5457), .Z(n5447) );
  AND U4951 ( .A(n5458), .B(n5459), .Z(n5457) );
  XOR U4952 ( .A(n5456), .B(n4584), .Z(n5459) );
  XNOR U4953 ( .A(p_input[7767]), .B(n5460), .Z(n4584) );
  AND U4954 ( .A(n203), .B(n5461), .Z(n5460) );
  XOR U4955 ( .A(p_input[7799]), .B(p_input[7767]), .Z(n5461) );
  XNOR U4956 ( .A(n4581), .B(n5456), .Z(n5458) );
  XOR U4957 ( .A(n5462), .B(n5463), .Z(n4581) );
  AND U4958 ( .A(n200), .B(n5464), .Z(n5463) );
  XOR U4959 ( .A(p_input[7735]), .B(p_input[7703]), .Z(n5464) );
  XOR U4960 ( .A(n5465), .B(n5466), .Z(n5456) );
  AND U4961 ( .A(n5467), .B(n5468), .Z(n5466) );
  XOR U4962 ( .A(n5465), .B(n4596), .Z(n5468) );
  XNOR U4963 ( .A(p_input[7766]), .B(n5469), .Z(n4596) );
  AND U4964 ( .A(n203), .B(n5470), .Z(n5469) );
  XOR U4965 ( .A(p_input[7798]), .B(p_input[7766]), .Z(n5470) );
  XNOR U4966 ( .A(n4593), .B(n5465), .Z(n5467) );
  XOR U4967 ( .A(n5471), .B(n5472), .Z(n4593) );
  AND U4968 ( .A(n200), .B(n5473), .Z(n5472) );
  XOR U4969 ( .A(p_input[7734]), .B(p_input[7702]), .Z(n5473) );
  XOR U4970 ( .A(n5474), .B(n5475), .Z(n5465) );
  AND U4971 ( .A(n5476), .B(n5477), .Z(n5475) );
  XOR U4972 ( .A(n5474), .B(n4608), .Z(n5477) );
  XNOR U4973 ( .A(p_input[7765]), .B(n5478), .Z(n4608) );
  AND U4974 ( .A(n203), .B(n5479), .Z(n5478) );
  XOR U4975 ( .A(p_input[7797]), .B(p_input[7765]), .Z(n5479) );
  XNOR U4976 ( .A(n4605), .B(n5474), .Z(n5476) );
  XOR U4977 ( .A(n5480), .B(n5481), .Z(n4605) );
  AND U4978 ( .A(n200), .B(n5482), .Z(n5481) );
  XOR U4979 ( .A(p_input[7733]), .B(p_input[7701]), .Z(n5482) );
  XOR U4980 ( .A(n5483), .B(n5484), .Z(n5474) );
  AND U4981 ( .A(n5485), .B(n5486), .Z(n5484) );
  XOR U4982 ( .A(n5483), .B(n4620), .Z(n5486) );
  XNOR U4983 ( .A(p_input[7764]), .B(n5487), .Z(n4620) );
  AND U4984 ( .A(n203), .B(n5488), .Z(n5487) );
  XOR U4985 ( .A(p_input[7796]), .B(p_input[7764]), .Z(n5488) );
  XNOR U4986 ( .A(n4617), .B(n5483), .Z(n5485) );
  XOR U4987 ( .A(n5489), .B(n5490), .Z(n4617) );
  AND U4988 ( .A(n200), .B(n5491), .Z(n5490) );
  XOR U4989 ( .A(p_input[7732]), .B(p_input[7700]), .Z(n5491) );
  XOR U4990 ( .A(n5492), .B(n5493), .Z(n5483) );
  AND U4991 ( .A(n5494), .B(n5495), .Z(n5493) );
  XOR U4992 ( .A(n5492), .B(n4632), .Z(n5495) );
  XNOR U4993 ( .A(p_input[7763]), .B(n5496), .Z(n4632) );
  AND U4994 ( .A(n203), .B(n5497), .Z(n5496) );
  XOR U4995 ( .A(p_input[7795]), .B(p_input[7763]), .Z(n5497) );
  XNOR U4996 ( .A(n4629), .B(n5492), .Z(n5494) );
  XOR U4997 ( .A(n5498), .B(n5499), .Z(n4629) );
  AND U4998 ( .A(n200), .B(n5500), .Z(n5499) );
  XOR U4999 ( .A(p_input[7731]), .B(p_input[7699]), .Z(n5500) );
  XOR U5000 ( .A(n5501), .B(n5502), .Z(n5492) );
  AND U5001 ( .A(n5503), .B(n5504), .Z(n5502) );
  XOR U5002 ( .A(n5501), .B(n4644), .Z(n5504) );
  XNOR U5003 ( .A(p_input[7762]), .B(n5505), .Z(n4644) );
  AND U5004 ( .A(n203), .B(n5506), .Z(n5505) );
  XOR U5005 ( .A(p_input[7794]), .B(p_input[7762]), .Z(n5506) );
  XNOR U5006 ( .A(n4641), .B(n5501), .Z(n5503) );
  XOR U5007 ( .A(n5507), .B(n5508), .Z(n4641) );
  AND U5008 ( .A(n200), .B(n5509), .Z(n5508) );
  XOR U5009 ( .A(p_input[7730]), .B(p_input[7698]), .Z(n5509) );
  XOR U5010 ( .A(n5510), .B(n5511), .Z(n5501) );
  AND U5011 ( .A(n5512), .B(n5513), .Z(n5511) );
  XOR U5012 ( .A(n5510), .B(n4656), .Z(n5513) );
  XNOR U5013 ( .A(p_input[7761]), .B(n5514), .Z(n4656) );
  AND U5014 ( .A(n203), .B(n5515), .Z(n5514) );
  XOR U5015 ( .A(p_input[7793]), .B(p_input[7761]), .Z(n5515) );
  XNOR U5016 ( .A(n4653), .B(n5510), .Z(n5512) );
  XOR U5017 ( .A(n5516), .B(n5517), .Z(n4653) );
  AND U5018 ( .A(n200), .B(n5518), .Z(n5517) );
  XOR U5019 ( .A(p_input[7729]), .B(p_input[7697]), .Z(n5518) );
  XOR U5020 ( .A(n5519), .B(n5520), .Z(n5510) );
  AND U5021 ( .A(n5521), .B(n5522), .Z(n5520) );
  XOR U5022 ( .A(n5519), .B(n4668), .Z(n5522) );
  XNOR U5023 ( .A(p_input[7760]), .B(n5523), .Z(n4668) );
  AND U5024 ( .A(n203), .B(n5524), .Z(n5523) );
  XOR U5025 ( .A(p_input[7792]), .B(p_input[7760]), .Z(n5524) );
  XNOR U5026 ( .A(n4665), .B(n5519), .Z(n5521) );
  XOR U5027 ( .A(n5525), .B(n5526), .Z(n4665) );
  AND U5028 ( .A(n200), .B(n5527), .Z(n5526) );
  XOR U5029 ( .A(p_input[7728]), .B(p_input[7696]), .Z(n5527) );
  XOR U5030 ( .A(n5528), .B(n5529), .Z(n5519) );
  AND U5031 ( .A(n5530), .B(n5531), .Z(n5529) );
  XOR U5032 ( .A(n5528), .B(n4680), .Z(n5531) );
  XNOR U5033 ( .A(p_input[7759]), .B(n5532), .Z(n4680) );
  AND U5034 ( .A(n203), .B(n5533), .Z(n5532) );
  XOR U5035 ( .A(p_input[7791]), .B(p_input[7759]), .Z(n5533) );
  XNOR U5036 ( .A(n4677), .B(n5528), .Z(n5530) );
  XOR U5037 ( .A(n5534), .B(n5535), .Z(n4677) );
  AND U5038 ( .A(n200), .B(n5536), .Z(n5535) );
  XOR U5039 ( .A(p_input[7727]), .B(p_input[7695]), .Z(n5536) );
  XOR U5040 ( .A(n5537), .B(n5538), .Z(n5528) );
  AND U5041 ( .A(n5539), .B(n5540), .Z(n5538) );
  XOR U5042 ( .A(n5537), .B(n4692), .Z(n5540) );
  XNOR U5043 ( .A(p_input[7758]), .B(n5541), .Z(n4692) );
  AND U5044 ( .A(n203), .B(n5542), .Z(n5541) );
  XOR U5045 ( .A(p_input[7790]), .B(p_input[7758]), .Z(n5542) );
  XNOR U5046 ( .A(n4689), .B(n5537), .Z(n5539) );
  XOR U5047 ( .A(n5543), .B(n5544), .Z(n4689) );
  AND U5048 ( .A(n200), .B(n5545), .Z(n5544) );
  XOR U5049 ( .A(p_input[7726]), .B(p_input[7694]), .Z(n5545) );
  XOR U5050 ( .A(n5546), .B(n5547), .Z(n5537) );
  AND U5051 ( .A(n5548), .B(n5549), .Z(n5547) );
  XOR U5052 ( .A(n5546), .B(n4704), .Z(n5549) );
  XNOR U5053 ( .A(p_input[7757]), .B(n5550), .Z(n4704) );
  AND U5054 ( .A(n203), .B(n5551), .Z(n5550) );
  XOR U5055 ( .A(p_input[7789]), .B(p_input[7757]), .Z(n5551) );
  XNOR U5056 ( .A(n4701), .B(n5546), .Z(n5548) );
  XOR U5057 ( .A(n5552), .B(n5553), .Z(n4701) );
  AND U5058 ( .A(n200), .B(n5554), .Z(n5553) );
  XOR U5059 ( .A(p_input[7725]), .B(p_input[7693]), .Z(n5554) );
  XOR U5060 ( .A(n5555), .B(n5556), .Z(n5546) );
  AND U5061 ( .A(n5557), .B(n5558), .Z(n5556) );
  XOR U5062 ( .A(n5555), .B(n4716), .Z(n5558) );
  XNOR U5063 ( .A(p_input[7756]), .B(n5559), .Z(n4716) );
  AND U5064 ( .A(n203), .B(n5560), .Z(n5559) );
  XOR U5065 ( .A(p_input[7788]), .B(p_input[7756]), .Z(n5560) );
  XNOR U5066 ( .A(n4713), .B(n5555), .Z(n5557) );
  XOR U5067 ( .A(n5561), .B(n5562), .Z(n4713) );
  AND U5068 ( .A(n200), .B(n5563), .Z(n5562) );
  XOR U5069 ( .A(p_input[7724]), .B(p_input[7692]), .Z(n5563) );
  XOR U5070 ( .A(n5564), .B(n5565), .Z(n5555) );
  AND U5071 ( .A(n5566), .B(n5567), .Z(n5565) );
  XOR U5072 ( .A(n5564), .B(n4728), .Z(n5567) );
  XNOR U5073 ( .A(p_input[7755]), .B(n5568), .Z(n4728) );
  AND U5074 ( .A(n203), .B(n5569), .Z(n5568) );
  XOR U5075 ( .A(p_input[7787]), .B(p_input[7755]), .Z(n5569) );
  XNOR U5076 ( .A(n4725), .B(n5564), .Z(n5566) );
  XOR U5077 ( .A(n5570), .B(n5571), .Z(n4725) );
  AND U5078 ( .A(n200), .B(n5572), .Z(n5571) );
  XOR U5079 ( .A(p_input[7723]), .B(p_input[7691]), .Z(n5572) );
  XOR U5080 ( .A(n5573), .B(n5574), .Z(n5564) );
  AND U5081 ( .A(n5575), .B(n5576), .Z(n5574) );
  XOR U5082 ( .A(n5573), .B(n4740), .Z(n5576) );
  XNOR U5083 ( .A(p_input[7754]), .B(n5577), .Z(n4740) );
  AND U5084 ( .A(n203), .B(n5578), .Z(n5577) );
  XOR U5085 ( .A(p_input[7786]), .B(p_input[7754]), .Z(n5578) );
  XNOR U5086 ( .A(n4737), .B(n5573), .Z(n5575) );
  XOR U5087 ( .A(n5579), .B(n5580), .Z(n4737) );
  AND U5088 ( .A(n200), .B(n5581), .Z(n5580) );
  XOR U5089 ( .A(p_input[7722]), .B(p_input[7690]), .Z(n5581) );
  XOR U5090 ( .A(n5582), .B(n5583), .Z(n5573) );
  AND U5091 ( .A(n5584), .B(n5585), .Z(n5583) );
  XOR U5092 ( .A(n5582), .B(n4752), .Z(n5585) );
  XNOR U5093 ( .A(p_input[7753]), .B(n5586), .Z(n4752) );
  AND U5094 ( .A(n203), .B(n5587), .Z(n5586) );
  XOR U5095 ( .A(p_input[7785]), .B(p_input[7753]), .Z(n5587) );
  XNOR U5096 ( .A(n4749), .B(n5582), .Z(n5584) );
  XOR U5097 ( .A(n5588), .B(n5589), .Z(n4749) );
  AND U5098 ( .A(n200), .B(n5590), .Z(n5589) );
  XOR U5099 ( .A(p_input[7721]), .B(p_input[7689]), .Z(n5590) );
  XOR U5100 ( .A(n5591), .B(n5592), .Z(n5582) );
  AND U5101 ( .A(n5593), .B(n5594), .Z(n5592) );
  XOR U5102 ( .A(n5591), .B(n4764), .Z(n5594) );
  XNOR U5103 ( .A(p_input[7752]), .B(n5595), .Z(n4764) );
  AND U5104 ( .A(n203), .B(n5596), .Z(n5595) );
  XOR U5105 ( .A(p_input[7784]), .B(p_input[7752]), .Z(n5596) );
  XNOR U5106 ( .A(n4761), .B(n5591), .Z(n5593) );
  XOR U5107 ( .A(n5597), .B(n5598), .Z(n4761) );
  AND U5108 ( .A(n200), .B(n5599), .Z(n5598) );
  XOR U5109 ( .A(p_input[7720]), .B(p_input[7688]), .Z(n5599) );
  XOR U5110 ( .A(n5600), .B(n5601), .Z(n5591) );
  AND U5111 ( .A(n5602), .B(n5603), .Z(n5601) );
  XOR U5112 ( .A(n5600), .B(n4776), .Z(n5603) );
  XNOR U5113 ( .A(p_input[7751]), .B(n5604), .Z(n4776) );
  AND U5114 ( .A(n203), .B(n5605), .Z(n5604) );
  XOR U5115 ( .A(p_input[7783]), .B(p_input[7751]), .Z(n5605) );
  XNOR U5116 ( .A(n4773), .B(n5600), .Z(n5602) );
  XOR U5117 ( .A(n5606), .B(n5607), .Z(n4773) );
  AND U5118 ( .A(n200), .B(n5608), .Z(n5607) );
  XOR U5119 ( .A(p_input[7719]), .B(p_input[7687]), .Z(n5608) );
  XOR U5120 ( .A(n5609), .B(n5610), .Z(n5600) );
  AND U5121 ( .A(n5611), .B(n5612), .Z(n5610) );
  XOR U5122 ( .A(n5609), .B(n4788), .Z(n5612) );
  XNOR U5123 ( .A(p_input[7750]), .B(n5613), .Z(n4788) );
  AND U5124 ( .A(n203), .B(n5614), .Z(n5613) );
  XOR U5125 ( .A(p_input[7782]), .B(p_input[7750]), .Z(n5614) );
  XNOR U5126 ( .A(n4785), .B(n5609), .Z(n5611) );
  XOR U5127 ( .A(n5615), .B(n5616), .Z(n4785) );
  AND U5128 ( .A(n200), .B(n5617), .Z(n5616) );
  XOR U5129 ( .A(p_input[7718]), .B(p_input[7686]), .Z(n5617) );
  XOR U5130 ( .A(n5618), .B(n5619), .Z(n5609) );
  AND U5131 ( .A(n5620), .B(n5621), .Z(n5619) );
  XOR U5132 ( .A(n5618), .B(n4800), .Z(n5621) );
  XNOR U5133 ( .A(p_input[7749]), .B(n5622), .Z(n4800) );
  AND U5134 ( .A(n203), .B(n5623), .Z(n5622) );
  XOR U5135 ( .A(p_input[7781]), .B(p_input[7749]), .Z(n5623) );
  XNOR U5136 ( .A(n4797), .B(n5618), .Z(n5620) );
  XOR U5137 ( .A(n5624), .B(n5625), .Z(n4797) );
  AND U5138 ( .A(n200), .B(n5626), .Z(n5625) );
  XOR U5139 ( .A(p_input[7717]), .B(p_input[7685]), .Z(n5626) );
  XOR U5140 ( .A(n5627), .B(n5628), .Z(n5618) );
  AND U5141 ( .A(n5629), .B(n5630), .Z(n5628) );
  XOR U5142 ( .A(n5627), .B(n4812), .Z(n5630) );
  XNOR U5143 ( .A(p_input[7748]), .B(n5631), .Z(n4812) );
  AND U5144 ( .A(n203), .B(n5632), .Z(n5631) );
  XOR U5145 ( .A(p_input[7780]), .B(p_input[7748]), .Z(n5632) );
  XNOR U5146 ( .A(n4809), .B(n5627), .Z(n5629) );
  XOR U5147 ( .A(n5633), .B(n5634), .Z(n4809) );
  AND U5148 ( .A(n200), .B(n5635), .Z(n5634) );
  XOR U5149 ( .A(p_input[7716]), .B(p_input[7684]), .Z(n5635) );
  XOR U5150 ( .A(n5636), .B(n5637), .Z(n5627) );
  AND U5151 ( .A(n5638), .B(n5639), .Z(n5637) );
  XOR U5152 ( .A(n5636), .B(n4824), .Z(n5639) );
  XNOR U5153 ( .A(p_input[7747]), .B(n5640), .Z(n4824) );
  AND U5154 ( .A(n203), .B(n5641), .Z(n5640) );
  XOR U5155 ( .A(p_input[7779]), .B(p_input[7747]), .Z(n5641) );
  XNOR U5156 ( .A(n4821), .B(n5636), .Z(n5638) );
  XOR U5157 ( .A(n5642), .B(n5643), .Z(n4821) );
  AND U5158 ( .A(n200), .B(n5644), .Z(n5643) );
  XOR U5159 ( .A(p_input[7715]), .B(p_input[7683]), .Z(n5644) );
  XOR U5160 ( .A(n5645), .B(n5646), .Z(n5636) );
  AND U5161 ( .A(n5647), .B(n5648), .Z(n5646) );
  XOR U5162 ( .A(n5645), .B(n4836), .Z(n5648) );
  XNOR U5163 ( .A(p_input[7746]), .B(n5649), .Z(n4836) );
  AND U5164 ( .A(n203), .B(n5650), .Z(n5649) );
  XOR U5165 ( .A(p_input[7778]), .B(p_input[7746]), .Z(n5650) );
  XNOR U5166 ( .A(n4833), .B(n5645), .Z(n5647) );
  XOR U5167 ( .A(n5651), .B(n5652), .Z(n4833) );
  AND U5168 ( .A(n200), .B(n5653), .Z(n5652) );
  XOR U5169 ( .A(p_input[7714]), .B(p_input[7682]), .Z(n5653) );
  XOR U5170 ( .A(n5654), .B(n5655), .Z(n5645) );
  AND U5171 ( .A(n5656), .B(n5657), .Z(n5655) );
  XNOR U5172 ( .A(n5658), .B(n4849), .Z(n5657) );
  XNOR U5173 ( .A(p_input[7745]), .B(n5659), .Z(n4849) );
  AND U5174 ( .A(n203), .B(n5660), .Z(n5659) );
  XNOR U5175 ( .A(p_input[7777]), .B(n5661), .Z(n5660) );
  IV U5176 ( .A(p_input[7745]), .Z(n5661) );
  XNOR U5177 ( .A(n4846), .B(n5654), .Z(n5656) );
  XNOR U5178 ( .A(p_input[7681]), .B(n5662), .Z(n4846) );
  AND U5179 ( .A(n200), .B(n5663), .Z(n5662) );
  XOR U5180 ( .A(p_input[7713]), .B(p_input[7681]), .Z(n5663) );
  IV U5181 ( .A(n5658), .Z(n5654) );
  AND U5182 ( .A(n5384), .B(n5387), .Z(n5658) );
  XOR U5183 ( .A(p_input[7744]), .B(n5664), .Z(n5387) );
  AND U5184 ( .A(n203), .B(n5665), .Z(n5664) );
  XOR U5185 ( .A(p_input[7776]), .B(p_input[7744]), .Z(n5665) );
  XOR U5186 ( .A(n5666), .B(n5667), .Z(n203) );
  AND U5187 ( .A(n5668), .B(n5669), .Z(n5667) );
  XNOR U5188 ( .A(p_input[7807]), .B(n5666), .Z(n5669) );
  XOR U5189 ( .A(n5666), .B(p_input[7775]), .Z(n5668) );
  XOR U5190 ( .A(n5670), .B(n5671), .Z(n5666) );
  AND U5191 ( .A(n5672), .B(n5673), .Z(n5671) );
  XNOR U5192 ( .A(p_input[7806]), .B(n5670), .Z(n5673) );
  XOR U5193 ( .A(n5670), .B(p_input[7774]), .Z(n5672) );
  XOR U5194 ( .A(n5674), .B(n5675), .Z(n5670) );
  AND U5195 ( .A(n5676), .B(n5677), .Z(n5675) );
  XNOR U5196 ( .A(p_input[7805]), .B(n5674), .Z(n5677) );
  XOR U5197 ( .A(n5674), .B(p_input[7773]), .Z(n5676) );
  XOR U5198 ( .A(n5678), .B(n5679), .Z(n5674) );
  AND U5199 ( .A(n5680), .B(n5681), .Z(n5679) );
  XNOR U5200 ( .A(p_input[7804]), .B(n5678), .Z(n5681) );
  XOR U5201 ( .A(n5678), .B(p_input[7772]), .Z(n5680) );
  XOR U5202 ( .A(n5682), .B(n5683), .Z(n5678) );
  AND U5203 ( .A(n5684), .B(n5685), .Z(n5683) );
  XNOR U5204 ( .A(p_input[7803]), .B(n5682), .Z(n5685) );
  XOR U5205 ( .A(n5682), .B(p_input[7771]), .Z(n5684) );
  XOR U5206 ( .A(n5686), .B(n5687), .Z(n5682) );
  AND U5207 ( .A(n5688), .B(n5689), .Z(n5687) );
  XNOR U5208 ( .A(p_input[7802]), .B(n5686), .Z(n5689) );
  XOR U5209 ( .A(n5686), .B(p_input[7770]), .Z(n5688) );
  XOR U5210 ( .A(n5690), .B(n5691), .Z(n5686) );
  AND U5211 ( .A(n5692), .B(n5693), .Z(n5691) );
  XNOR U5212 ( .A(p_input[7801]), .B(n5690), .Z(n5693) );
  XOR U5213 ( .A(n5690), .B(p_input[7769]), .Z(n5692) );
  XOR U5214 ( .A(n5694), .B(n5695), .Z(n5690) );
  AND U5215 ( .A(n5696), .B(n5697), .Z(n5695) );
  XNOR U5216 ( .A(p_input[7800]), .B(n5694), .Z(n5697) );
  XOR U5217 ( .A(n5694), .B(p_input[7768]), .Z(n5696) );
  XOR U5218 ( .A(n5698), .B(n5699), .Z(n5694) );
  AND U5219 ( .A(n5700), .B(n5701), .Z(n5699) );
  XNOR U5220 ( .A(p_input[7799]), .B(n5698), .Z(n5701) );
  XOR U5221 ( .A(n5698), .B(p_input[7767]), .Z(n5700) );
  XOR U5222 ( .A(n5702), .B(n5703), .Z(n5698) );
  AND U5223 ( .A(n5704), .B(n5705), .Z(n5703) );
  XNOR U5224 ( .A(p_input[7798]), .B(n5702), .Z(n5705) );
  XOR U5225 ( .A(n5702), .B(p_input[7766]), .Z(n5704) );
  XOR U5226 ( .A(n5706), .B(n5707), .Z(n5702) );
  AND U5227 ( .A(n5708), .B(n5709), .Z(n5707) );
  XNOR U5228 ( .A(p_input[7797]), .B(n5706), .Z(n5709) );
  XOR U5229 ( .A(n5706), .B(p_input[7765]), .Z(n5708) );
  XOR U5230 ( .A(n5710), .B(n5711), .Z(n5706) );
  AND U5231 ( .A(n5712), .B(n5713), .Z(n5711) );
  XNOR U5232 ( .A(p_input[7796]), .B(n5710), .Z(n5713) );
  XOR U5233 ( .A(n5710), .B(p_input[7764]), .Z(n5712) );
  XOR U5234 ( .A(n5714), .B(n5715), .Z(n5710) );
  AND U5235 ( .A(n5716), .B(n5717), .Z(n5715) );
  XNOR U5236 ( .A(p_input[7795]), .B(n5714), .Z(n5717) );
  XOR U5237 ( .A(n5714), .B(p_input[7763]), .Z(n5716) );
  XOR U5238 ( .A(n5718), .B(n5719), .Z(n5714) );
  AND U5239 ( .A(n5720), .B(n5721), .Z(n5719) );
  XNOR U5240 ( .A(p_input[7794]), .B(n5718), .Z(n5721) );
  XOR U5241 ( .A(n5718), .B(p_input[7762]), .Z(n5720) );
  XOR U5242 ( .A(n5722), .B(n5723), .Z(n5718) );
  AND U5243 ( .A(n5724), .B(n5725), .Z(n5723) );
  XNOR U5244 ( .A(p_input[7793]), .B(n5722), .Z(n5725) );
  XOR U5245 ( .A(n5722), .B(p_input[7761]), .Z(n5724) );
  XOR U5246 ( .A(n5726), .B(n5727), .Z(n5722) );
  AND U5247 ( .A(n5728), .B(n5729), .Z(n5727) );
  XNOR U5248 ( .A(p_input[7792]), .B(n5726), .Z(n5729) );
  XOR U5249 ( .A(n5726), .B(p_input[7760]), .Z(n5728) );
  XOR U5250 ( .A(n5730), .B(n5731), .Z(n5726) );
  AND U5251 ( .A(n5732), .B(n5733), .Z(n5731) );
  XNOR U5252 ( .A(p_input[7791]), .B(n5730), .Z(n5733) );
  XOR U5253 ( .A(n5730), .B(p_input[7759]), .Z(n5732) );
  XOR U5254 ( .A(n5734), .B(n5735), .Z(n5730) );
  AND U5255 ( .A(n5736), .B(n5737), .Z(n5735) );
  XNOR U5256 ( .A(p_input[7790]), .B(n5734), .Z(n5737) );
  XOR U5257 ( .A(n5734), .B(p_input[7758]), .Z(n5736) );
  XOR U5258 ( .A(n5738), .B(n5739), .Z(n5734) );
  AND U5259 ( .A(n5740), .B(n5741), .Z(n5739) );
  XNOR U5260 ( .A(p_input[7789]), .B(n5738), .Z(n5741) );
  XOR U5261 ( .A(n5738), .B(p_input[7757]), .Z(n5740) );
  XOR U5262 ( .A(n5742), .B(n5743), .Z(n5738) );
  AND U5263 ( .A(n5744), .B(n5745), .Z(n5743) );
  XNOR U5264 ( .A(p_input[7788]), .B(n5742), .Z(n5745) );
  XOR U5265 ( .A(n5742), .B(p_input[7756]), .Z(n5744) );
  XOR U5266 ( .A(n5746), .B(n5747), .Z(n5742) );
  AND U5267 ( .A(n5748), .B(n5749), .Z(n5747) );
  XNOR U5268 ( .A(p_input[7787]), .B(n5746), .Z(n5749) );
  XOR U5269 ( .A(n5746), .B(p_input[7755]), .Z(n5748) );
  XOR U5270 ( .A(n5750), .B(n5751), .Z(n5746) );
  AND U5271 ( .A(n5752), .B(n5753), .Z(n5751) );
  XNOR U5272 ( .A(p_input[7786]), .B(n5750), .Z(n5753) );
  XOR U5273 ( .A(n5750), .B(p_input[7754]), .Z(n5752) );
  XOR U5274 ( .A(n5754), .B(n5755), .Z(n5750) );
  AND U5275 ( .A(n5756), .B(n5757), .Z(n5755) );
  XNOR U5276 ( .A(p_input[7785]), .B(n5754), .Z(n5757) );
  XOR U5277 ( .A(n5754), .B(p_input[7753]), .Z(n5756) );
  XOR U5278 ( .A(n5758), .B(n5759), .Z(n5754) );
  AND U5279 ( .A(n5760), .B(n5761), .Z(n5759) );
  XNOR U5280 ( .A(p_input[7784]), .B(n5758), .Z(n5761) );
  XOR U5281 ( .A(n5758), .B(p_input[7752]), .Z(n5760) );
  XOR U5282 ( .A(n5762), .B(n5763), .Z(n5758) );
  AND U5283 ( .A(n5764), .B(n5765), .Z(n5763) );
  XNOR U5284 ( .A(p_input[7783]), .B(n5762), .Z(n5765) );
  XOR U5285 ( .A(n5762), .B(p_input[7751]), .Z(n5764) );
  XOR U5286 ( .A(n5766), .B(n5767), .Z(n5762) );
  AND U5287 ( .A(n5768), .B(n5769), .Z(n5767) );
  XNOR U5288 ( .A(p_input[7782]), .B(n5766), .Z(n5769) );
  XOR U5289 ( .A(n5766), .B(p_input[7750]), .Z(n5768) );
  XOR U5290 ( .A(n5770), .B(n5771), .Z(n5766) );
  AND U5291 ( .A(n5772), .B(n5773), .Z(n5771) );
  XNOR U5292 ( .A(p_input[7781]), .B(n5770), .Z(n5773) );
  XOR U5293 ( .A(n5770), .B(p_input[7749]), .Z(n5772) );
  XOR U5294 ( .A(n5774), .B(n5775), .Z(n5770) );
  AND U5295 ( .A(n5776), .B(n5777), .Z(n5775) );
  XNOR U5296 ( .A(p_input[7780]), .B(n5774), .Z(n5777) );
  XOR U5297 ( .A(n5774), .B(p_input[7748]), .Z(n5776) );
  XOR U5298 ( .A(n5778), .B(n5779), .Z(n5774) );
  AND U5299 ( .A(n5780), .B(n5781), .Z(n5779) );
  XNOR U5300 ( .A(p_input[7779]), .B(n5778), .Z(n5781) );
  XOR U5301 ( .A(n5778), .B(p_input[7747]), .Z(n5780) );
  XOR U5302 ( .A(n5782), .B(n5783), .Z(n5778) );
  AND U5303 ( .A(n5784), .B(n5785), .Z(n5783) );
  XNOR U5304 ( .A(p_input[7778]), .B(n5782), .Z(n5785) );
  XOR U5305 ( .A(n5782), .B(p_input[7746]), .Z(n5784) );
  XNOR U5306 ( .A(n5786), .B(n5787), .Z(n5782) );
  AND U5307 ( .A(n5788), .B(n5789), .Z(n5787) );
  XOR U5308 ( .A(p_input[7777]), .B(n5786), .Z(n5789) );
  XNOR U5309 ( .A(p_input[7745]), .B(n5786), .Z(n5788) );
  AND U5310 ( .A(p_input[7776]), .B(n5790), .Z(n5786) );
  IV U5311 ( .A(p_input[7744]), .Z(n5790) );
  XNOR U5312 ( .A(p_input[7680]), .B(n5791), .Z(n5384) );
  AND U5313 ( .A(n200), .B(n5792), .Z(n5791) );
  XOR U5314 ( .A(p_input[7712]), .B(p_input[7680]), .Z(n5792) );
  XOR U5315 ( .A(n5793), .B(n5794), .Z(n200) );
  AND U5316 ( .A(n5795), .B(n5796), .Z(n5794) );
  XNOR U5317 ( .A(p_input[7743]), .B(n5793), .Z(n5796) );
  XOR U5318 ( .A(n5793), .B(p_input[7711]), .Z(n5795) );
  XOR U5319 ( .A(n5797), .B(n5798), .Z(n5793) );
  AND U5320 ( .A(n5799), .B(n5800), .Z(n5798) );
  XNOR U5321 ( .A(p_input[7742]), .B(n5797), .Z(n5800) );
  XNOR U5322 ( .A(n5797), .B(n5399), .Z(n5799) );
  IV U5323 ( .A(p_input[7710]), .Z(n5399) );
  XOR U5324 ( .A(n5801), .B(n5802), .Z(n5797) );
  AND U5325 ( .A(n5803), .B(n5804), .Z(n5802) );
  XNOR U5326 ( .A(p_input[7741]), .B(n5801), .Z(n5804) );
  XNOR U5327 ( .A(n5801), .B(n5408), .Z(n5803) );
  IV U5328 ( .A(p_input[7709]), .Z(n5408) );
  XOR U5329 ( .A(n5805), .B(n5806), .Z(n5801) );
  AND U5330 ( .A(n5807), .B(n5808), .Z(n5806) );
  XNOR U5331 ( .A(p_input[7740]), .B(n5805), .Z(n5808) );
  XNOR U5332 ( .A(n5805), .B(n5417), .Z(n5807) );
  IV U5333 ( .A(p_input[7708]), .Z(n5417) );
  XOR U5334 ( .A(n5809), .B(n5810), .Z(n5805) );
  AND U5335 ( .A(n5811), .B(n5812), .Z(n5810) );
  XNOR U5336 ( .A(p_input[7739]), .B(n5809), .Z(n5812) );
  XNOR U5337 ( .A(n5809), .B(n5426), .Z(n5811) );
  IV U5338 ( .A(p_input[7707]), .Z(n5426) );
  XOR U5339 ( .A(n5813), .B(n5814), .Z(n5809) );
  AND U5340 ( .A(n5815), .B(n5816), .Z(n5814) );
  XNOR U5341 ( .A(p_input[7738]), .B(n5813), .Z(n5816) );
  XNOR U5342 ( .A(n5813), .B(n5435), .Z(n5815) );
  IV U5343 ( .A(p_input[7706]), .Z(n5435) );
  XOR U5344 ( .A(n5817), .B(n5818), .Z(n5813) );
  AND U5345 ( .A(n5819), .B(n5820), .Z(n5818) );
  XNOR U5346 ( .A(p_input[7737]), .B(n5817), .Z(n5820) );
  XNOR U5347 ( .A(n5817), .B(n5444), .Z(n5819) );
  IV U5348 ( .A(p_input[7705]), .Z(n5444) );
  XOR U5349 ( .A(n5821), .B(n5822), .Z(n5817) );
  AND U5350 ( .A(n5823), .B(n5824), .Z(n5822) );
  XNOR U5351 ( .A(p_input[7736]), .B(n5821), .Z(n5824) );
  XNOR U5352 ( .A(n5821), .B(n5453), .Z(n5823) );
  IV U5353 ( .A(p_input[7704]), .Z(n5453) );
  XOR U5354 ( .A(n5825), .B(n5826), .Z(n5821) );
  AND U5355 ( .A(n5827), .B(n5828), .Z(n5826) );
  XNOR U5356 ( .A(p_input[7735]), .B(n5825), .Z(n5828) );
  XNOR U5357 ( .A(n5825), .B(n5462), .Z(n5827) );
  IV U5358 ( .A(p_input[7703]), .Z(n5462) );
  XOR U5359 ( .A(n5829), .B(n5830), .Z(n5825) );
  AND U5360 ( .A(n5831), .B(n5832), .Z(n5830) );
  XNOR U5361 ( .A(p_input[7734]), .B(n5829), .Z(n5832) );
  XNOR U5362 ( .A(n5829), .B(n5471), .Z(n5831) );
  IV U5363 ( .A(p_input[7702]), .Z(n5471) );
  XOR U5364 ( .A(n5833), .B(n5834), .Z(n5829) );
  AND U5365 ( .A(n5835), .B(n5836), .Z(n5834) );
  XNOR U5366 ( .A(p_input[7733]), .B(n5833), .Z(n5836) );
  XNOR U5367 ( .A(n5833), .B(n5480), .Z(n5835) );
  IV U5368 ( .A(p_input[7701]), .Z(n5480) );
  XOR U5369 ( .A(n5837), .B(n5838), .Z(n5833) );
  AND U5370 ( .A(n5839), .B(n5840), .Z(n5838) );
  XNOR U5371 ( .A(p_input[7732]), .B(n5837), .Z(n5840) );
  XNOR U5372 ( .A(n5837), .B(n5489), .Z(n5839) );
  IV U5373 ( .A(p_input[7700]), .Z(n5489) );
  XOR U5374 ( .A(n5841), .B(n5842), .Z(n5837) );
  AND U5375 ( .A(n5843), .B(n5844), .Z(n5842) );
  XNOR U5376 ( .A(p_input[7731]), .B(n5841), .Z(n5844) );
  XNOR U5377 ( .A(n5841), .B(n5498), .Z(n5843) );
  IV U5378 ( .A(p_input[7699]), .Z(n5498) );
  XOR U5379 ( .A(n5845), .B(n5846), .Z(n5841) );
  AND U5380 ( .A(n5847), .B(n5848), .Z(n5846) );
  XNOR U5381 ( .A(p_input[7730]), .B(n5845), .Z(n5848) );
  XNOR U5382 ( .A(n5845), .B(n5507), .Z(n5847) );
  IV U5383 ( .A(p_input[7698]), .Z(n5507) );
  XOR U5384 ( .A(n5849), .B(n5850), .Z(n5845) );
  AND U5385 ( .A(n5851), .B(n5852), .Z(n5850) );
  XNOR U5386 ( .A(p_input[7729]), .B(n5849), .Z(n5852) );
  XNOR U5387 ( .A(n5849), .B(n5516), .Z(n5851) );
  IV U5388 ( .A(p_input[7697]), .Z(n5516) );
  XOR U5389 ( .A(n5853), .B(n5854), .Z(n5849) );
  AND U5390 ( .A(n5855), .B(n5856), .Z(n5854) );
  XNOR U5391 ( .A(p_input[7728]), .B(n5853), .Z(n5856) );
  XNOR U5392 ( .A(n5853), .B(n5525), .Z(n5855) );
  IV U5393 ( .A(p_input[7696]), .Z(n5525) );
  XOR U5394 ( .A(n5857), .B(n5858), .Z(n5853) );
  AND U5395 ( .A(n5859), .B(n5860), .Z(n5858) );
  XNOR U5396 ( .A(p_input[7727]), .B(n5857), .Z(n5860) );
  XNOR U5397 ( .A(n5857), .B(n5534), .Z(n5859) );
  IV U5398 ( .A(p_input[7695]), .Z(n5534) );
  XOR U5399 ( .A(n5861), .B(n5862), .Z(n5857) );
  AND U5400 ( .A(n5863), .B(n5864), .Z(n5862) );
  XNOR U5401 ( .A(p_input[7726]), .B(n5861), .Z(n5864) );
  XNOR U5402 ( .A(n5861), .B(n5543), .Z(n5863) );
  IV U5403 ( .A(p_input[7694]), .Z(n5543) );
  XOR U5404 ( .A(n5865), .B(n5866), .Z(n5861) );
  AND U5405 ( .A(n5867), .B(n5868), .Z(n5866) );
  XNOR U5406 ( .A(p_input[7725]), .B(n5865), .Z(n5868) );
  XNOR U5407 ( .A(n5865), .B(n5552), .Z(n5867) );
  IV U5408 ( .A(p_input[7693]), .Z(n5552) );
  XOR U5409 ( .A(n5869), .B(n5870), .Z(n5865) );
  AND U5410 ( .A(n5871), .B(n5872), .Z(n5870) );
  XNOR U5411 ( .A(p_input[7724]), .B(n5869), .Z(n5872) );
  XNOR U5412 ( .A(n5869), .B(n5561), .Z(n5871) );
  IV U5413 ( .A(p_input[7692]), .Z(n5561) );
  XOR U5414 ( .A(n5873), .B(n5874), .Z(n5869) );
  AND U5415 ( .A(n5875), .B(n5876), .Z(n5874) );
  XNOR U5416 ( .A(p_input[7723]), .B(n5873), .Z(n5876) );
  XNOR U5417 ( .A(n5873), .B(n5570), .Z(n5875) );
  IV U5418 ( .A(p_input[7691]), .Z(n5570) );
  XOR U5419 ( .A(n5877), .B(n5878), .Z(n5873) );
  AND U5420 ( .A(n5879), .B(n5880), .Z(n5878) );
  XNOR U5421 ( .A(p_input[7722]), .B(n5877), .Z(n5880) );
  XNOR U5422 ( .A(n5877), .B(n5579), .Z(n5879) );
  IV U5423 ( .A(p_input[7690]), .Z(n5579) );
  XOR U5424 ( .A(n5881), .B(n5882), .Z(n5877) );
  AND U5425 ( .A(n5883), .B(n5884), .Z(n5882) );
  XNOR U5426 ( .A(p_input[7721]), .B(n5881), .Z(n5884) );
  XNOR U5427 ( .A(n5881), .B(n5588), .Z(n5883) );
  IV U5428 ( .A(p_input[7689]), .Z(n5588) );
  XOR U5429 ( .A(n5885), .B(n5886), .Z(n5881) );
  AND U5430 ( .A(n5887), .B(n5888), .Z(n5886) );
  XNOR U5431 ( .A(p_input[7720]), .B(n5885), .Z(n5888) );
  XNOR U5432 ( .A(n5885), .B(n5597), .Z(n5887) );
  IV U5433 ( .A(p_input[7688]), .Z(n5597) );
  XOR U5434 ( .A(n5889), .B(n5890), .Z(n5885) );
  AND U5435 ( .A(n5891), .B(n5892), .Z(n5890) );
  XNOR U5436 ( .A(p_input[7719]), .B(n5889), .Z(n5892) );
  XNOR U5437 ( .A(n5889), .B(n5606), .Z(n5891) );
  IV U5438 ( .A(p_input[7687]), .Z(n5606) );
  XOR U5439 ( .A(n5893), .B(n5894), .Z(n5889) );
  AND U5440 ( .A(n5895), .B(n5896), .Z(n5894) );
  XNOR U5441 ( .A(p_input[7718]), .B(n5893), .Z(n5896) );
  XNOR U5442 ( .A(n5893), .B(n5615), .Z(n5895) );
  IV U5443 ( .A(p_input[7686]), .Z(n5615) );
  XOR U5444 ( .A(n5897), .B(n5898), .Z(n5893) );
  AND U5445 ( .A(n5899), .B(n5900), .Z(n5898) );
  XNOR U5446 ( .A(p_input[7717]), .B(n5897), .Z(n5900) );
  XNOR U5447 ( .A(n5897), .B(n5624), .Z(n5899) );
  IV U5448 ( .A(p_input[7685]), .Z(n5624) );
  XOR U5449 ( .A(n5901), .B(n5902), .Z(n5897) );
  AND U5450 ( .A(n5903), .B(n5904), .Z(n5902) );
  XNOR U5451 ( .A(p_input[7716]), .B(n5901), .Z(n5904) );
  XNOR U5452 ( .A(n5901), .B(n5633), .Z(n5903) );
  IV U5453 ( .A(p_input[7684]), .Z(n5633) );
  XOR U5454 ( .A(n5905), .B(n5906), .Z(n5901) );
  AND U5455 ( .A(n5907), .B(n5908), .Z(n5906) );
  XNOR U5456 ( .A(p_input[7715]), .B(n5905), .Z(n5908) );
  XNOR U5457 ( .A(n5905), .B(n5642), .Z(n5907) );
  IV U5458 ( .A(p_input[7683]), .Z(n5642) );
  XOR U5459 ( .A(n5909), .B(n5910), .Z(n5905) );
  AND U5460 ( .A(n5911), .B(n5912), .Z(n5910) );
  XNOR U5461 ( .A(p_input[7714]), .B(n5909), .Z(n5912) );
  XNOR U5462 ( .A(n5909), .B(n5651), .Z(n5911) );
  IV U5463 ( .A(p_input[7682]), .Z(n5651) );
  XNOR U5464 ( .A(n5913), .B(n5914), .Z(n5909) );
  AND U5465 ( .A(n5915), .B(n5916), .Z(n5914) );
  XOR U5466 ( .A(p_input[7713]), .B(n5913), .Z(n5916) );
  XNOR U5467 ( .A(p_input[7681]), .B(n5913), .Z(n5915) );
  AND U5468 ( .A(p_input[7712]), .B(n5917), .Z(n5913) );
  IV U5469 ( .A(p_input[7680]), .Z(n5917) );
  XOR U5470 ( .A(n5918), .B(n5919), .Z(n2274) );
  AND U5471 ( .A(n997), .B(n5920), .Z(n5919) );
  XNOR U5472 ( .A(n5921), .B(n5918), .Z(n5920) );
  XOR U5473 ( .A(n5922), .B(n5923), .Z(n997) );
  AND U5474 ( .A(n5924), .B(n5925), .Z(n5923) );
  XOR U5475 ( .A(n5922), .B(n2289), .Z(n5925) );
  XOR U5476 ( .A(n5926), .B(n5927), .Z(n2289) );
  AND U5477 ( .A(n819), .B(n5928), .Z(n5927) );
  XOR U5478 ( .A(n5929), .B(n5926), .Z(n5928) );
  XNOR U5479 ( .A(n2286), .B(n5922), .Z(n5924) );
  XOR U5480 ( .A(n5930), .B(n5931), .Z(n2286) );
  AND U5481 ( .A(n816), .B(n5932), .Z(n5931) );
  XOR U5482 ( .A(n5933), .B(n5930), .Z(n5932) );
  XOR U5483 ( .A(n5934), .B(n5935), .Z(n5922) );
  AND U5484 ( .A(n5936), .B(n5937), .Z(n5935) );
  XOR U5485 ( .A(n5934), .B(n2301), .Z(n5937) );
  XOR U5486 ( .A(n5938), .B(n5939), .Z(n2301) );
  AND U5487 ( .A(n819), .B(n5940), .Z(n5939) );
  XOR U5488 ( .A(n5941), .B(n5938), .Z(n5940) );
  XNOR U5489 ( .A(n2298), .B(n5934), .Z(n5936) );
  XOR U5490 ( .A(n5942), .B(n5943), .Z(n2298) );
  AND U5491 ( .A(n816), .B(n5944), .Z(n5943) );
  XOR U5492 ( .A(n5945), .B(n5942), .Z(n5944) );
  XOR U5493 ( .A(n5946), .B(n5947), .Z(n5934) );
  AND U5494 ( .A(n5948), .B(n5949), .Z(n5947) );
  XOR U5495 ( .A(n5946), .B(n2313), .Z(n5949) );
  XOR U5496 ( .A(n5950), .B(n5951), .Z(n2313) );
  AND U5497 ( .A(n819), .B(n5952), .Z(n5951) );
  XOR U5498 ( .A(n5953), .B(n5950), .Z(n5952) );
  XNOR U5499 ( .A(n2310), .B(n5946), .Z(n5948) );
  XOR U5500 ( .A(n5954), .B(n5955), .Z(n2310) );
  AND U5501 ( .A(n816), .B(n5956), .Z(n5955) );
  XOR U5502 ( .A(n5957), .B(n5954), .Z(n5956) );
  XOR U5503 ( .A(n5958), .B(n5959), .Z(n5946) );
  AND U5504 ( .A(n5960), .B(n5961), .Z(n5959) );
  XOR U5505 ( .A(n5958), .B(n2325), .Z(n5961) );
  XOR U5506 ( .A(n5962), .B(n5963), .Z(n2325) );
  AND U5507 ( .A(n819), .B(n5964), .Z(n5963) );
  XOR U5508 ( .A(n5965), .B(n5962), .Z(n5964) );
  XNOR U5509 ( .A(n2322), .B(n5958), .Z(n5960) );
  XOR U5510 ( .A(n5966), .B(n5967), .Z(n2322) );
  AND U5511 ( .A(n816), .B(n5968), .Z(n5967) );
  XOR U5512 ( .A(n5969), .B(n5966), .Z(n5968) );
  XOR U5513 ( .A(n5970), .B(n5971), .Z(n5958) );
  AND U5514 ( .A(n5972), .B(n5973), .Z(n5971) );
  XOR U5515 ( .A(n5970), .B(n2337), .Z(n5973) );
  XOR U5516 ( .A(n5974), .B(n5975), .Z(n2337) );
  AND U5517 ( .A(n819), .B(n5976), .Z(n5975) );
  XOR U5518 ( .A(n5977), .B(n5974), .Z(n5976) );
  XNOR U5519 ( .A(n2334), .B(n5970), .Z(n5972) );
  XOR U5520 ( .A(n5978), .B(n5979), .Z(n2334) );
  AND U5521 ( .A(n816), .B(n5980), .Z(n5979) );
  XOR U5522 ( .A(n5981), .B(n5978), .Z(n5980) );
  XOR U5523 ( .A(n5982), .B(n5983), .Z(n5970) );
  AND U5524 ( .A(n5984), .B(n5985), .Z(n5983) );
  XOR U5525 ( .A(n5982), .B(n2349), .Z(n5985) );
  XOR U5526 ( .A(n5986), .B(n5987), .Z(n2349) );
  AND U5527 ( .A(n819), .B(n5988), .Z(n5987) );
  XOR U5528 ( .A(n5989), .B(n5986), .Z(n5988) );
  XNOR U5529 ( .A(n2346), .B(n5982), .Z(n5984) );
  XOR U5530 ( .A(n5990), .B(n5991), .Z(n2346) );
  AND U5531 ( .A(n816), .B(n5992), .Z(n5991) );
  XOR U5532 ( .A(n5993), .B(n5990), .Z(n5992) );
  XOR U5533 ( .A(n5994), .B(n5995), .Z(n5982) );
  AND U5534 ( .A(n5996), .B(n5997), .Z(n5995) );
  XOR U5535 ( .A(n5994), .B(n2361), .Z(n5997) );
  XOR U5536 ( .A(n5998), .B(n5999), .Z(n2361) );
  AND U5537 ( .A(n819), .B(n6000), .Z(n5999) );
  XOR U5538 ( .A(n6001), .B(n5998), .Z(n6000) );
  XNOR U5539 ( .A(n2358), .B(n5994), .Z(n5996) );
  XOR U5540 ( .A(n6002), .B(n6003), .Z(n2358) );
  AND U5541 ( .A(n816), .B(n6004), .Z(n6003) );
  XOR U5542 ( .A(n6005), .B(n6002), .Z(n6004) );
  XOR U5543 ( .A(n6006), .B(n6007), .Z(n5994) );
  AND U5544 ( .A(n6008), .B(n6009), .Z(n6007) );
  XOR U5545 ( .A(n6006), .B(n2373), .Z(n6009) );
  XOR U5546 ( .A(n6010), .B(n6011), .Z(n2373) );
  AND U5547 ( .A(n819), .B(n6012), .Z(n6011) );
  XOR U5548 ( .A(n6013), .B(n6010), .Z(n6012) );
  XNOR U5549 ( .A(n2370), .B(n6006), .Z(n6008) );
  XOR U5550 ( .A(n6014), .B(n6015), .Z(n2370) );
  AND U5551 ( .A(n816), .B(n6016), .Z(n6015) );
  XOR U5552 ( .A(n6017), .B(n6014), .Z(n6016) );
  XOR U5553 ( .A(n6018), .B(n6019), .Z(n6006) );
  AND U5554 ( .A(n6020), .B(n6021), .Z(n6019) );
  XOR U5555 ( .A(n6018), .B(n2385), .Z(n6021) );
  XOR U5556 ( .A(n6022), .B(n6023), .Z(n2385) );
  AND U5557 ( .A(n819), .B(n6024), .Z(n6023) );
  XOR U5558 ( .A(n6025), .B(n6022), .Z(n6024) );
  XNOR U5559 ( .A(n2382), .B(n6018), .Z(n6020) );
  XOR U5560 ( .A(n6026), .B(n6027), .Z(n2382) );
  AND U5561 ( .A(n816), .B(n6028), .Z(n6027) );
  XOR U5562 ( .A(n6029), .B(n6026), .Z(n6028) );
  XOR U5563 ( .A(n6030), .B(n6031), .Z(n6018) );
  AND U5564 ( .A(n6032), .B(n6033), .Z(n6031) );
  XOR U5565 ( .A(n6030), .B(n2397), .Z(n6033) );
  XOR U5566 ( .A(n6034), .B(n6035), .Z(n2397) );
  AND U5567 ( .A(n819), .B(n6036), .Z(n6035) );
  XOR U5568 ( .A(n6037), .B(n6034), .Z(n6036) );
  XNOR U5569 ( .A(n2394), .B(n6030), .Z(n6032) );
  XOR U5570 ( .A(n6038), .B(n6039), .Z(n2394) );
  AND U5571 ( .A(n816), .B(n6040), .Z(n6039) );
  XOR U5572 ( .A(n6041), .B(n6038), .Z(n6040) );
  XOR U5573 ( .A(n6042), .B(n6043), .Z(n6030) );
  AND U5574 ( .A(n6044), .B(n6045), .Z(n6043) );
  XOR U5575 ( .A(n6042), .B(n2409), .Z(n6045) );
  XOR U5576 ( .A(n6046), .B(n6047), .Z(n2409) );
  AND U5577 ( .A(n819), .B(n6048), .Z(n6047) );
  XOR U5578 ( .A(n6049), .B(n6046), .Z(n6048) );
  XNOR U5579 ( .A(n2406), .B(n6042), .Z(n6044) );
  XOR U5580 ( .A(n6050), .B(n6051), .Z(n2406) );
  AND U5581 ( .A(n816), .B(n6052), .Z(n6051) );
  XOR U5582 ( .A(n6053), .B(n6050), .Z(n6052) );
  XOR U5583 ( .A(n6054), .B(n6055), .Z(n6042) );
  AND U5584 ( .A(n6056), .B(n6057), .Z(n6055) );
  XOR U5585 ( .A(n6054), .B(n2421), .Z(n6057) );
  XOR U5586 ( .A(n6058), .B(n6059), .Z(n2421) );
  AND U5587 ( .A(n819), .B(n6060), .Z(n6059) );
  XOR U5588 ( .A(n6061), .B(n6058), .Z(n6060) );
  XNOR U5589 ( .A(n2418), .B(n6054), .Z(n6056) );
  XOR U5590 ( .A(n6062), .B(n6063), .Z(n2418) );
  AND U5591 ( .A(n816), .B(n6064), .Z(n6063) );
  XOR U5592 ( .A(n6065), .B(n6062), .Z(n6064) );
  XOR U5593 ( .A(n6066), .B(n6067), .Z(n6054) );
  AND U5594 ( .A(n6068), .B(n6069), .Z(n6067) );
  XOR U5595 ( .A(n6066), .B(n2433), .Z(n6069) );
  XOR U5596 ( .A(n6070), .B(n6071), .Z(n2433) );
  AND U5597 ( .A(n819), .B(n6072), .Z(n6071) );
  XOR U5598 ( .A(n6073), .B(n6070), .Z(n6072) );
  XNOR U5599 ( .A(n2430), .B(n6066), .Z(n6068) );
  XOR U5600 ( .A(n6074), .B(n6075), .Z(n2430) );
  AND U5601 ( .A(n816), .B(n6076), .Z(n6075) );
  XOR U5602 ( .A(n6077), .B(n6074), .Z(n6076) );
  XOR U5603 ( .A(n6078), .B(n6079), .Z(n6066) );
  AND U5604 ( .A(n6080), .B(n6081), .Z(n6079) );
  XOR U5605 ( .A(n6078), .B(n2445), .Z(n6081) );
  XOR U5606 ( .A(n6082), .B(n6083), .Z(n2445) );
  AND U5607 ( .A(n819), .B(n6084), .Z(n6083) );
  XOR U5608 ( .A(n6085), .B(n6082), .Z(n6084) );
  XNOR U5609 ( .A(n2442), .B(n6078), .Z(n6080) );
  XOR U5610 ( .A(n6086), .B(n6087), .Z(n2442) );
  AND U5611 ( .A(n816), .B(n6088), .Z(n6087) );
  XOR U5612 ( .A(n6089), .B(n6086), .Z(n6088) );
  XOR U5613 ( .A(n6090), .B(n6091), .Z(n6078) );
  AND U5614 ( .A(n6092), .B(n6093), .Z(n6091) );
  XOR U5615 ( .A(n6090), .B(n2457), .Z(n6093) );
  XOR U5616 ( .A(n6094), .B(n6095), .Z(n2457) );
  AND U5617 ( .A(n819), .B(n6096), .Z(n6095) );
  XOR U5618 ( .A(n6097), .B(n6094), .Z(n6096) );
  XNOR U5619 ( .A(n2454), .B(n6090), .Z(n6092) );
  XOR U5620 ( .A(n6098), .B(n6099), .Z(n2454) );
  AND U5621 ( .A(n816), .B(n6100), .Z(n6099) );
  XOR U5622 ( .A(n6101), .B(n6098), .Z(n6100) );
  XOR U5623 ( .A(n6102), .B(n6103), .Z(n6090) );
  AND U5624 ( .A(n6104), .B(n6105), .Z(n6103) );
  XOR U5625 ( .A(n6102), .B(n2469), .Z(n6105) );
  XOR U5626 ( .A(n6106), .B(n6107), .Z(n2469) );
  AND U5627 ( .A(n819), .B(n6108), .Z(n6107) );
  XOR U5628 ( .A(n6109), .B(n6106), .Z(n6108) );
  XNOR U5629 ( .A(n2466), .B(n6102), .Z(n6104) );
  XOR U5630 ( .A(n6110), .B(n6111), .Z(n2466) );
  AND U5631 ( .A(n816), .B(n6112), .Z(n6111) );
  XOR U5632 ( .A(n6113), .B(n6110), .Z(n6112) );
  XOR U5633 ( .A(n6114), .B(n6115), .Z(n6102) );
  AND U5634 ( .A(n6116), .B(n6117), .Z(n6115) );
  XOR U5635 ( .A(n6114), .B(n2481), .Z(n6117) );
  XOR U5636 ( .A(n6118), .B(n6119), .Z(n2481) );
  AND U5637 ( .A(n819), .B(n6120), .Z(n6119) );
  XOR U5638 ( .A(n6121), .B(n6118), .Z(n6120) );
  XNOR U5639 ( .A(n2478), .B(n6114), .Z(n6116) );
  XOR U5640 ( .A(n6122), .B(n6123), .Z(n2478) );
  AND U5641 ( .A(n816), .B(n6124), .Z(n6123) );
  XOR U5642 ( .A(n6125), .B(n6122), .Z(n6124) );
  XOR U5643 ( .A(n6126), .B(n6127), .Z(n6114) );
  AND U5644 ( .A(n6128), .B(n6129), .Z(n6127) );
  XOR U5645 ( .A(n6126), .B(n2493), .Z(n6129) );
  XOR U5646 ( .A(n6130), .B(n6131), .Z(n2493) );
  AND U5647 ( .A(n819), .B(n6132), .Z(n6131) );
  XOR U5648 ( .A(n6133), .B(n6130), .Z(n6132) );
  XNOR U5649 ( .A(n2490), .B(n6126), .Z(n6128) );
  XOR U5650 ( .A(n6134), .B(n6135), .Z(n2490) );
  AND U5651 ( .A(n816), .B(n6136), .Z(n6135) );
  XOR U5652 ( .A(n6137), .B(n6134), .Z(n6136) );
  XOR U5653 ( .A(n6138), .B(n6139), .Z(n6126) );
  AND U5654 ( .A(n6140), .B(n6141), .Z(n6139) );
  XOR U5655 ( .A(n6138), .B(n2505), .Z(n6141) );
  XOR U5656 ( .A(n6142), .B(n6143), .Z(n2505) );
  AND U5657 ( .A(n819), .B(n6144), .Z(n6143) );
  XOR U5658 ( .A(n6145), .B(n6142), .Z(n6144) );
  XNOR U5659 ( .A(n2502), .B(n6138), .Z(n6140) );
  XOR U5660 ( .A(n6146), .B(n6147), .Z(n2502) );
  AND U5661 ( .A(n816), .B(n6148), .Z(n6147) );
  XOR U5662 ( .A(n6149), .B(n6146), .Z(n6148) );
  XOR U5663 ( .A(n6150), .B(n6151), .Z(n6138) );
  AND U5664 ( .A(n6152), .B(n6153), .Z(n6151) );
  XOR U5665 ( .A(n6150), .B(n2517), .Z(n6153) );
  XOR U5666 ( .A(n6154), .B(n6155), .Z(n2517) );
  AND U5667 ( .A(n819), .B(n6156), .Z(n6155) );
  XOR U5668 ( .A(n6157), .B(n6154), .Z(n6156) );
  XNOR U5669 ( .A(n2514), .B(n6150), .Z(n6152) );
  XOR U5670 ( .A(n6158), .B(n6159), .Z(n2514) );
  AND U5671 ( .A(n816), .B(n6160), .Z(n6159) );
  XOR U5672 ( .A(n6161), .B(n6158), .Z(n6160) );
  XOR U5673 ( .A(n6162), .B(n6163), .Z(n6150) );
  AND U5674 ( .A(n6164), .B(n6165), .Z(n6163) );
  XOR U5675 ( .A(n6162), .B(n2529), .Z(n6165) );
  XOR U5676 ( .A(n6166), .B(n6167), .Z(n2529) );
  AND U5677 ( .A(n819), .B(n6168), .Z(n6167) );
  XOR U5678 ( .A(n6169), .B(n6166), .Z(n6168) );
  XNOR U5679 ( .A(n2526), .B(n6162), .Z(n6164) );
  XOR U5680 ( .A(n6170), .B(n6171), .Z(n2526) );
  AND U5681 ( .A(n816), .B(n6172), .Z(n6171) );
  XOR U5682 ( .A(n6173), .B(n6170), .Z(n6172) );
  XOR U5683 ( .A(n6174), .B(n6175), .Z(n6162) );
  AND U5684 ( .A(n6176), .B(n6177), .Z(n6175) );
  XOR U5685 ( .A(n6174), .B(n2541), .Z(n6177) );
  XOR U5686 ( .A(n6178), .B(n6179), .Z(n2541) );
  AND U5687 ( .A(n819), .B(n6180), .Z(n6179) );
  XOR U5688 ( .A(n6181), .B(n6178), .Z(n6180) );
  XNOR U5689 ( .A(n2538), .B(n6174), .Z(n6176) );
  XOR U5690 ( .A(n6182), .B(n6183), .Z(n2538) );
  AND U5691 ( .A(n816), .B(n6184), .Z(n6183) );
  XOR U5692 ( .A(n6185), .B(n6182), .Z(n6184) );
  XOR U5693 ( .A(n6186), .B(n6187), .Z(n6174) );
  AND U5694 ( .A(n6188), .B(n6189), .Z(n6187) );
  XOR U5695 ( .A(n6186), .B(n2553), .Z(n6189) );
  XOR U5696 ( .A(n6190), .B(n6191), .Z(n2553) );
  AND U5697 ( .A(n819), .B(n6192), .Z(n6191) );
  XOR U5698 ( .A(n6193), .B(n6190), .Z(n6192) );
  XNOR U5699 ( .A(n2550), .B(n6186), .Z(n6188) );
  XOR U5700 ( .A(n6194), .B(n6195), .Z(n2550) );
  AND U5701 ( .A(n816), .B(n6196), .Z(n6195) );
  XOR U5702 ( .A(n6197), .B(n6194), .Z(n6196) );
  XOR U5703 ( .A(n6198), .B(n6199), .Z(n6186) );
  AND U5704 ( .A(n6200), .B(n6201), .Z(n6199) );
  XOR U5705 ( .A(n6198), .B(n2565), .Z(n6201) );
  XOR U5706 ( .A(n6202), .B(n6203), .Z(n2565) );
  AND U5707 ( .A(n819), .B(n6204), .Z(n6203) );
  XOR U5708 ( .A(n6205), .B(n6202), .Z(n6204) );
  XNOR U5709 ( .A(n2562), .B(n6198), .Z(n6200) );
  XOR U5710 ( .A(n6206), .B(n6207), .Z(n2562) );
  AND U5711 ( .A(n816), .B(n6208), .Z(n6207) );
  XOR U5712 ( .A(n6209), .B(n6206), .Z(n6208) );
  XOR U5713 ( .A(n6210), .B(n6211), .Z(n6198) );
  AND U5714 ( .A(n6212), .B(n6213), .Z(n6211) );
  XOR U5715 ( .A(n6210), .B(n2577), .Z(n6213) );
  XOR U5716 ( .A(n6214), .B(n6215), .Z(n2577) );
  AND U5717 ( .A(n819), .B(n6216), .Z(n6215) );
  XOR U5718 ( .A(n6217), .B(n6214), .Z(n6216) );
  XNOR U5719 ( .A(n2574), .B(n6210), .Z(n6212) );
  XOR U5720 ( .A(n6218), .B(n6219), .Z(n2574) );
  AND U5721 ( .A(n816), .B(n6220), .Z(n6219) );
  XOR U5722 ( .A(n6221), .B(n6218), .Z(n6220) );
  XOR U5723 ( .A(n6222), .B(n6223), .Z(n6210) );
  AND U5724 ( .A(n6224), .B(n6225), .Z(n6223) );
  XOR U5725 ( .A(n6222), .B(n2589), .Z(n6225) );
  XOR U5726 ( .A(n6226), .B(n6227), .Z(n2589) );
  AND U5727 ( .A(n819), .B(n6228), .Z(n6227) );
  XOR U5728 ( .A(n6229), .B(n6226), .Z(n6228) );
  XNOR U5729 ( .A(n2586), .B(n6222), .Z(n6224) );
  XOR U5730 ( .A(n6230), .B(n6231), .Z(n2586) );
  AND U5731 ( .A(n816), .B(n6232), .Z(n6231) );
  XOR U5732 ( .A(n6233), .B(n6230), .Z(n6232) );
  XOR U5733 ( .A(n6234), .B(n6235), .Z(n6222) );
  AND U5734 ( .A(n6236), .B(n6237), .Z(n6235) );
  XOR U5735 ( .A(n6234), .B(n2601), .Z(n6237) );
  XOR U5736 ( .A(n6238), .B(n6239), .Z(n2601) );
  AND U5737 ( .A(n819), .B(n6240), .Z(n6239) );
  XOR U5738 ( .A(n6241), .B(n6238), .Z(n6240) );
  XNOR U5739 ( .A(n2598), .B(n6234), .Z(n6236) );
  XOR U5740 ( .A(n6242), .B(n6243), .Z(n2598) );
  AND U5741 ( .A(n816), .B(n6244), .Z(n6243) );
  XOR U5742 ( .A(n6245), .B(n6242), .Z(n6244) );
  XOR U5743 ( .A(n6246), .B(n6247), .Z(n6234) );
  AND U5744 ( .A(n6248), .B(n6249), .Z(n6247) );
  XOR U5745 ( .A(n6246), .B(n2613), .Z(n6249) );
  XOR U5746 ( .A(n6250), .B(n6251), .Z(n2613) );
  AND U5747 ( .A(n819), .B(n6252), .Z(n6251) );
  XOR U5748 ( .A(n6253), .B(n6250), .Z(n6252) );
  XNOR U5749 ( .A(n2610), .B(n6246), .Z(n6248) );
  XOR U5750 ( .A(n6254), .B(n6255), .Z(n2610) );
  AND U5751 ( .A(n816), .B(n6256), .Z(n6255) );
  XOR U5752 ( .A(n6257), .B(n6254), .Z(n6256) );
  XOR U5753 ( .A(n6258), .B(n6259), .Z(n6246) );
  AND U5754 ( .A(n6260), .B(n6261), .Z(n6259) );
  XOR U5755 ( .A(n6258), .B(n2625), .Z(n6261) );
  XOR U5756 ( .A(n6262), .B(n6263), .Z(n2625) );
  AND U5757 ( .A(n819), .B(n6264), .Z(n6263) );
  XOR U5758 ( .A(n6265), .B(n6262), .Z(n6264) );
  XNOR U5759 ( .A(n2622), .B(n6258), .Z(n6260) );
  XOR U5760 ( .A(n6266), .B(n6267), .Z(n2622) );
  AND U5761 ( .A(n816), .B(n6268), .Z(n6267) );
  XOR U5762 ( .A(n6269), .B(n6266), .Z(n6268) );
  XOR U5763 ( .A(n6270), .B(n6271), .Z(n6258) );
  AND U5764 ( .A(n6272), .B(n6273), .Z(n6271) );
  XOR U5765 ( .A(n6270), .B(n2637), .Z(n6273) );
  XOR U5766 ( .A(n6274), .B(n6275), .Z(n2637) );
  AND U5767 ( .A(n819), .B(n6276), .Z(n6275) );
  XOR U5768 ( .A(n6277), .B(n6274), .Z(n6276) );
  XNOR U5769 ( .A(n2634), .B(n6270), .Z(n6272) );
  XOR U5770 ( .A(n6278), .B(n6279), .Z(n2634) );
  AND U5771 ( .A(n816), .B(n6280), .Z(n6279) );
  XOR U5772 ( .A(n6281), .B(n6278), .Z(n6280) );
  XOR U5773 ( .A(n6282), .B(n6283), .Z(n6270) );
  AND U5774 ( .A(n6284), .B(n6285), .Z(n6283) );
  XNOR U5775 ( .A(n6286), .B(n2650), .Z(n6285) );
  XOR U5776 ( .A(n6287), .B(n6288), .Z(n2650) );
  AND U5777 ( .A(n819), .B(n6289), .Z(n6288) );
  XOR U5778 ( .A(n6287), .B(n6290), .Z(n6289) );
  XNOR U5779 ( .A(n2647), .B(n6282), .Z(n6284) );
  XOR U5780 ( .A(n6291), .B(n6292), .Z(n2647) );
  AND U5781 ( .A(n816), .B(n6293), .Z(n6292) );
  XOR U5782 ( .A(n6291), .B(n6294), .Z(n6293) );
  IV U5783 ( .A(n6286), .Z(n6282) );
  AND U5784 ( .A(n5918), .B(n5921), .Z(n6286) );
  XNOR U5785 ( .A(n6295), .B(n6296), .Z(n5921) );
  AND U5786 ( .A(n819), .B(n6297), .Z(n6296) );
  XNOR U5787 ( .A(n6298), .B(n6295), .Z(n6297) );
  XOR U5788 ( .A(n6299), .B(n6300), .Z(n819) );
  AND U5789 ( .A(n6301), .B(n6302), .Z(n6300) );
  XOR U5790 ( .A(n6299), .B(n5929), .Z(n6302) );
  XNOR U5791 ( .A(n6303), .B(n6304), .Z(n5929) );
  AND U5792 ( .A(n6305), .B(n451), .Z(n6304) );
  AND U5793 ( .A(n6303), .B(n6306), .Z(n6305) );
  XNOR U5794 ( .A(n5926), .B(n6299), .Z(n6301) );
  XOR U5795 ( .A(n6307), .B(n6308), .Z(n5926) );
  AND U5796 ( .A(n6309), .B(n449), .Z(n6308) );
  NOR U5797 ( .A(n6307), .B(n6310), .Z(n6309) );
  XOR U5798 ( .A(n6311), .B(n6312), .Z(n6299) );
  AND U5799 ( .A(n6313), .B(n6314), .Z(n6312) );
  XOR U5800 ( .A(n6311), .B(n5941), .Z(n6314) );
  XOR U5801 ( .A(n6315), .B(n6316), .Z(n5941) );
  AND U5802 ( .A(n451), .B(n6317), .Z(n6316) );
  XOR U5803 ( .A(n6318), .B(n6315), .Z(n6317) );
  XNOR U5804 ( .A(n5938), .B(n6311), .Z(n6313) );
  XOR U5805 ( .A(n6319), .B(n6320), .Z(n5938) );
  AND U5806 ( .A(n449), .B(n6321), .Z(n6320) );
  XOR U5807 ( .A(n6322), .B(n6319), .Z(n6321) );
  XOR U5808 ( .A(n6323), .B(n6324), .Z(n6311) );
  AND U5809 ( .A(n6325), .B(n6326), .Z(n6324) );
  XOR U5810 ( .A(n6323), .B(n5953), .Z(n6326) );
  XOR U5811 ( .A(n6327), .B(n6328), .Z(n5953) );
  AND U5812 ( .A(n451), .B(n6329), .Z(n6328) );
  XOR U5813 ( .A(n6330), .B(n6327), .Z(n6329) );
  XNOR U5814 ( .A(n5950), .B(n6323), .Z(n6325) );
  XOR U5815 ( .A(n6331), .B(n6332), .Z(n5950) );
  AND U5816 ( .A(n449), .B(n6333), .Z(n6332) );
  XOR U5817 ( .A(n6334), .B(n6331), .Z(n6333) );
  XOR U5818 ( .A(n6335), .B(n6336), .Z(n6323) );
  AND U5819 ( .A(n6337), .B(n6338), .Z(n6336) );
  XOR U5820 ( .A(n6335), .B(n5965), .Z(n6338) );
  XOR U5821 ( .A(n6339), .B(n6340), .Z(n5965) );
  AND U5822 ( .A(n451), .B(n6341), .Z(n6340) );
  XOR U5823 ( .A(n6342), .B(n6339), .Z(n6341) );
  XNOR U5824 ( .A(n5962), .B(n6335), .Z(n6337) );
  XOR U5825 ( .A(n6343), .B(n6344), .Z(n5962) );
  AND U5826 ( .A(n449), .B(n6345), .Z(n6344) );
  XOR U5827 ( .A(n6346), .B(n6343), .Z(n6345) );
  XOR U5828 ( .A(n6347), .B(n6348), .Z(n6335) );
  AND U5829 ( .A(n6349), .B(n6350), .Z(n6348) );
  XOR U5830 ( .A(n6347), .B(n5977), .Z(n6350) );
  XOR U5831 ( .A(n6351), .B(n6352), .Z(n5977) );
  AND U5832 ( .A(n451), .B(n6353), .Z(n6352) );
  XOR U5833 ( .A(n6354), .B(n6351), .Z(n6353) );
  XNOR U5834 ( .A(n5974), .B(n6347), .Z(n6349) );
  XOR U5835 ( .A(n6355), .B(n6356), .Z(n5974) );
  AND U5836 ( .A(n449), .B(n6357), .Z(n6356) );
  XOR U5837 ( .A(n6358), .B(n6355), .Z(n6357) );
  XOR U5838 ( .A(n6359), .B(n6360), .Z(n6347) );
  AND U5839 ( .A(n6361), .B(n6362), .Z(n6360) );
  XOR U5840 ( .A(n6359), .B(n5989), .Z(n6362) );
  XOR U5841 ( .A(n6363), .B(n6364), .Z(n5989) );
  AND U5842 ( .A(n451), .B(n6365), .Z(n6364) );
  XOR U5843 ( .A(n6366), .B(n6363), .Z(n6365) );
  XNOR U5844 ( .A(n5986), .B(n6359), .Z(n6361) );
  XOR U5845 ( .A(n6367), .B(n6368), .Z(n5986) );
  AND U5846 ( .A(n449), .B(n6369), .Z(n6368) );
  XOR U5847 ( .A(n6370), .B(n6367), .Z(n6369) );
  XOR U5848 ( .A(n6371), .B(n6372), .Z(n6359) );
  AND U5849 ( .A(n6373), .B(n6374), .Z(n6372) );
  XOR U5850 ( .A(n6371), .B(n6001), .Z(n6374) );
  XOR U5851 ( .A(n6375), .B(n6376), .Z(n6001) );
  AND U5852 ( .A(n451), .B(n6377), .Z(n6376) );
  XOR U5853 ( .A(n6378), .B(n6375), .Z(n6377) );
  XNOR U5854 ( .A(n5998), .B(n6371), .Z(n6373) );
  XOR U5855 ( .A(n6379), .B(n6380), .Z(n5998) );
  AND U5856 ( .A(n449), .B(n6381), .Z(n6380) );
  XOR U5857 ( .A(n6382), .B(n6379), .Z(n6381) );
  XOR U5858 ( .A(n6383), .B(n6384), .Z(n6371) );
  AND U5859 ( .A(n6385), .B(n6386), .Z(n6384) );
  XOR U5860 ( .A(n6383), .B(n6013), .Z(n6386) );
  XOR U5861 ( .A(n6387), .B(n6388), .Z(n6013) );
  AND U5862 ( .A(n451), .B(n6389), .Z(n6388) );
  XOR U5863 ( .A(n6390), .B(n6387), .Z(n6389) );
  XNOR U5864 ( .A(n6010), .B(n6383), .Z(n6385) );
  XOR U5865 ( .A(n6391), .B(n6392), .Z(n6010) );
  AND U5866 ( .A(n449), .B(n6393), .Z(n6392) );
  XOR U5867 ( .A(n6394), .B(n6391), .Z(n6393) );
  XOR U5868 ( .A(n6395), .B(n6396), .Z(n6383) );
  AND U5869 ( .A(n6397), .B(n6398), .Z(n6396) );
  XOR U5870 ( .A(n6395), .B(n6025), .Z(n6398) );
  XOR U5871 ( .A(n6399), .B(n6400), .Z(n6025) );
  AND U5872 ( .A(n451), .B(n6401), .Z(n6400) );
  XOR U5873 ( .A(n6402), .B(n6399), .Z(n6401) );
  XNOR U5874 ( .A(n6022), .B(n6395), .Z(n6397) );
  XOR U5875 ( .A(n6403), .B(n6404), .Z(n6022) );
  AND U5876 ( .A(n449), .B(n6405), .Z(n6404) );
  XOR U5877 ( .A(n6406), .B(n6403), .Z(n6405) );
  XOR U5878 ( .A(n6407), .B(n6408), .Z(n6395) );
  AND U5879 ( .A(n6409), .B(n6410), .Z(n6408) );
  XOR U5880 ( .A(n6407), .B(n6037), .Z(n6410) );
  XOR U5881 ( .A(n6411), .B(n6412), .Z(n6037) );
  AND U5882 ( .A(n451), .B(n6413), .Z(n6412) );
  XOR U5883 ( .A(n6414), .B(n6411), .Z(n6413) );
  XNOR U5884 ( .A(n6034), .B(n6407), .Z(n6409) );
  XOR U5885 ( .A(n6415), .B(n6416), .Z(n6034) );
  AND U5886 ( .A(n449), .B(n6417), .Z(n6416) );
  XOR U5887 ( .A(n6418), .B(n6415), .Z(n6417) );
  XOR U5888 ( .A(n6419), .B(n6420), .Z(n6407) );
  AND U5889 ( .A(n6421), .B(n6422), .Z(n6420) );
  XOR U5890 ( .A(n6419), .B(n6049), .Z(n6422) );
  XOR U5891 ( .A(n6423), .B(n6424), .Z(n6049) );
  AND U5892 ( .A(n451), .B(n6425), .Z(n6424) );
  XOR U5893 ( .A(n6426), .B(n6423), .Z(n6425) );
  XNOR U5894 ( .A(n6046), .B(n6419), .Z(n6421) );
  XOR U5895 ( .A(n6427), .B(n6428), .Z(n6046) );
  AND U5896 ( .A(n449), .B(n6429), .Z(n6428) );
  XOR U5897 ( .A(n6430), .B(n6427), .Z(n6429) );
  XOR U5898 ( .A(n6431), .B(n6432), .Z(n6419) );
  AND U5899 ( .A(n6433), .B(n6434), .Z(n6432) );
  XOR U5900 ( .A(n6431), .B(n6061), .Z(n6434) );
  XOR U5901 ( .A(n6435), .B(n6436), .Z(n6061) );
  AND U5902 ( .A(n451), .B(n6437), .Z(n6436) );
  XOR U5903 ( .A(n6438), .B(n6435), .Z(n6437) );
  XNOR U5904 ( .A(n6058), .B(n6431), .Z(n6433) );
  XOR U5905 ( .A(n6439), .B(n6440), .Z(n6058) );
  AND U5906 ( .A(n449), .B(n6441), .Z(n6440) );
  XOR U5907 ( .A(n6442), .B(n6439), .Z(n6441) );
  XOR U5908 ( .A(n6443), .B(n6444), .Z(n6431) );
  AND U5909 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U5910 ( .A(n6443), .B(n6073), .Z(n6446) );
  XOR U5911 ( .A(n6447), .B(n6448), .Z(n6073) );
  AND U5912 ( .A(n451), .B(n6449), .Z(n6448) );
  XOR U5913 ( .A(n6450), .B(n6447), .Z(n6449) );
  XNOR U5914 ( .A(n6070), .B(n6443), .Z(n6445) );
  XOR U5915 ( .A(n6451), .B(n6452), .Z(n6070) );
  AND U5916 ( .A(n449), .B(n6453), .Z(n6452) );
  XOR U5917 ( .A(n6454), .B(n6451), .Z(n6453) );
  XOR U5918 ( .A(n6455), .B(n6456), .Z(n6443) );
  AND U5919 ( .A(n6457), .B(n6458), .Z(n6456) );
  XOR U5920 ( .A(n6455), .B(n6085), .Z(n6458) );
  XOR U5921 ( .A(n6459), .B(n6460), .Z(n6085) );
  AND U5922 ( .A(n451), .B(n6461), .Z(n6460) );
  XOR U5923 ( .A(n6462), .B(n6459), .Z(n6461) );
  XNOR U5924 ( .A(n6082), .B(n6455), .Z(n6457) );
  XOR U5925 ( .A(n6463), .B(n6464), .Z(n6082) );
  AND U5926 ( .A(n449), .B(n6465), .Z(n6464) );
  XOR U5927 ( .A(n6466), .B(n6463), .Z(n6465) );
  XOR U5928 ( .A(n6467), .B(n6468), .Z(n6455) );
  AND U5929 ( .A(n6469), .B(n6470), .Z(n6468) );
  XOR U5930 ( .A(n6467), .B(n6097), .Z(n6470) );
  XOR U5931 ( .A(n6471), .B(n6472), .Z(n6097) );
  AND U5932 ( .A(n451), .B(n6473), .Z(n6472) );
  XOR U5933 ( .A(n6474), .B(n6471), .Z(n6473) );
  XNOR U5934 ( .A(n6094), .B(n6467), .Z(n6469) );
  XOR U5935 ( .A(n6475), .B(n6476), .Z(n6094) );
  AND U5936 ( .A(n449), .B(n6477), .Z(n6476) );
  XOR U5937 ( .A(n6478), .B(n6475), .Z(n6477) );
  XOR U5938 ( .A(n6479), .B(n6480), .Z(n6467) );
  AND U5939 ( .A(n6481), .B(n6482), .Z(n6480) );
  XOR U5940 ( .A(n6479), .B(n6109), .Z(n6482) );
  XOR U5941 ( .A(n6483), .B(n6484), .Z(n6109) );
  AND U5942 ( .A(n451), .B(n6485), .Z(n6484) );
  XOR U5943 ( .A(n6486), .B(n6483), .Z(n6485) );
  XNOR U5944 ( .A(n6106), .B(n6479), .Z(n6481) );
  XOR U5945 ( .A(n6487), .B(n6488), .Z(n6106) );
  AND U5946 ( .A(n449), .B(n6489), .Z(n6488) );
  XOR U5947 ( .A(n6490), .B(n6487), .Z(n6489) );
  XOR U5948 ( .A(n6491), .B(n6492), .Z(n6479) );
  AND U5949 ( .A(n6493), .B(n6494), .Z(n6492) );
  XOR U5950 ( .A(n6491), .B(n6121), .Z(n6494) );
  XOR U5951 ( .A(n6495), .B(n6496), .Z(n6121) );
  AND U5952 ( .A(n451), .B(n6497), .Z(n6496) );
  XOR U5953 ( .A(n6498), .B(n6495), .Z(n6497) );
  XNOR U5954 ( .A(n6118), .B(n6491), .Z(n6493) );
  XOR U5955 ( .A(n6499), .B(n6500), .Z(n6118) );
  AND U5956 ( .A(n449), .B(n6501), .Z(n6500) );
  XOR U5957 ( .A(n6502), .B(n6499), .Z(n6501) );
  XOR U5958 ( .A(n6503), .B(n6504), .Z(n6491) );
  AND U5959 ( .A(n6505), .B(n6506), .Z(n6504) );
  XOR U5960 ( .A(n6503), .B(n6133), .Z(n6506) );
  XOR U5961 ( .A(n6507), .B(n6508), .Z(n6133) );
  AND U5962 ( .A(n451), .B(n6509), .Z(n6508) );
  XOR U5963 ( .A(n6510), .B(n6507), .Z(n6509) );
  XNOR U5964 ( .A(n6130), .B(n6503), .Z(n6505) );
  XOR U5965 ( .A(n6511), .B(n6512), .Z(n6130) );
  AND U5966 ( .A(n449), .B(n6513), .Z(n6512) );
  XOR U5967 ( .A(n6514), .B(n6511), .Z(n6513) );
  XOR U5968 ( .A(n6515), .B(n6516), .Z(n6503) );
  AND U5969 ( .A(n6517), .B(n6518), .Z(n6516) );
  XOR U5970 ( .A(n6515), .B(n6145), .Z(n6518) );
  XOR U5971 ( .A(n6519), .B(n6520), .Z(n6145) );
  AND U5972 ( .A(n451), .B(n6521), .Z(n6520) );
  XOR U5973 ( .A(n6522), .B(n6519), .Z(n6521) );
  XNOR U5974 ( .A(n6142), .B(n6515), .Z(n6517) );
  XOR U5975 ( .A(n6523), .B(n6524), .Z(n6142) );
  AND U5976 ( .A(n449), .B(n6525), .Z(n6524) );
  XOR U5977 ( .A(n6526), .B(n6523), .Z(n6525) );
  XOR U5978 ( .A(n6527), .B(n6528), .Z(n6515) );
  AND U5979 ( .A(n6529), .B(n6530), .Z(n6528) );
  XOR U5980 ( .A(n6527), .B(n6157), .Z(n6530) );
  XOR U5981 ( .A(n6531), .B(n6532), .Z(n6157) );
  AND U5982 ( .A(n451), .B(n6533), .Z(n6532) );
  XOR U5983 ( .A(n6534), .B(n6531), .Z(n6533) );
  XNOR U5984 ( .A(n6154), .B(n6527), .Z(n6529) );
  XOR U5985 ( .A(n6535), .B(n6536), .Z(n6154) );
  AND U5986 ( .A(n449), .B(n6537), .Z(n6536) );
  XOR U5987 ( .A(n6538), .B(n6535), .Z(n6537) );
  XOR U5988 ( .A(n6539), .B(n6540), .Z(n6527) );
  AND U5989 ( .A(n6541), .B(n6542), .Z(n6540) );
  XOR U5990 ( .A(n6539), .B(n6169), .Z(n6542) );
  XOR U5991 ( .A(n6543), .B(n6544), .Z(n6169) );
  AND U5992 ( .A(n451), .B(n6545), .Z(n6544) );
  XOR U5993 ( .A(n6546), .B(n6543), .Z(n6545) );
  XNOR U5994 ( .A(n6166), .B(n6539), .Z(n6541) );
  XOR U5995 ( .A(n6547), .B(n6548), .Z(n6166) );
  AND U5996 ( .A(n449), .B(n6549), .Z(n6548) );
  XOR U5997 ( .A(n6550), .B(n6547), .Z(n6549) );
  XOR U5998 ( .A(n6551), .B(n6552), .Z(n6539) );
  AND U5999 ( .A(n6553), .B(n6554), .Z(n6552) );
  XOR U6000 ( .A(n6551), .B(n6181), .Z(n6554) );
  XOR U6001 ( .A(n6555), .B(n6556), .Z(n6181) );
  AND U6002 ( .A(n451), .B(n6557), .Z(n6556) );
  XOR U6003 ( .A(n6558), .B(n6555), .Z(n6557) );
  XNOR U6004 ( .A(n6178), .B(n6551), .Z(n6553) );
  XOR U6005 ( .A(n6559), .B(n6560), .Z(n6178) );
  AND U6006 ( .A(n449), .B(n6561), .Z(n6560) );
  XOR U6007 ( .A(n6562), .B(n6559), .Z(n6561) );
  XOR U6008 ( .A(n6563), .B(n6564), .Z(n6551) );
  AND U6009 ( .A(n6565), .B(n6566), .Z(n6564) );
  XOR U6010 ( .A(n6563), .B(n6193), .Z(n6566) );
  XOR U6011 ( .A(n6567), .B(n6568), .Z(n6193) );
  AND U6012 ( .A(n451), .B(n6569), .Z(n6568) );
  XOR U6013 ( .A(n6570), .B(n6567), .Z(n6569) );
  XNOR U6014 ( .A(n6190), .B(n6563), .Z(n6565) );
  XOR U6015 ( .A(n6571), .B(n6572), .Z(n6190) );
  AND U6016 ( .A(n449), .B(n6573), .Z(n6572) );
  XOR U6017 ( .A(n6574), .B(n6571), .Z(n6573) );
  XOR U6018 ( .A(n6575), .B(n6576), .Z(n6563) );
  AND U6019 ( .A(n6577), .B(n6578), .Z(n6576) );
  XOR U6020 ( .A(n6575), .B(n6205), .Z(n6578) );
  XOR U6021 ( .A(n6579), .B(n6580), .Z(n6205) );
  AND U6022 ( .A(n451), .B(n6581), .Z(n6580) );
  XOR U6023 ( .A(n6582), .B(n6579), .Z(n6581) );
  XNOR U6024 ( .A(n6202), .B(n6575), .Z(n6577) );
  XOR U6025 ( .A(n6583), .B(n6584), .Z(n6202) );
  AND U6026 ( .A(n449), .B(n6585), .Z(n6584) );
  XOR U6027 ( .A(n6586), .B(n6583), .Z(n6585) );
  XOR U6028 ( .A(n6587), .B(n6588), .Z(n6575) );
  AND U6029 ( .A(n6589), .B(n6590), .Z(n6588) );
  XOR U6030 ( .A(n6587), .B(n6217), .Z(n6590) );
  XOR U6031 ( .A(n6591), .B(n6592), .Z(n6217) );
  AND U6032 ( .A(n451), .B(n6593), .Z(n6592) );
  XOR U6033 ( .A(n6594), .B(n6591), .Z(n6593) );
  XNOR U6034 ( .A(n6214), .B(n6587), .Z(n6589) );
  XOR U6035 ( .A(n6595), .B(n6596), .Z(n6214) );
  AND U6036 ( .A(n449), .B(n6597), .Z(n6596) );
  XOR U6037 ( .A(n6598), .B(n6595), .Z(n6597) );
  XOR U6038 ( .A(n6599), .B(n6600), .Z(n6587) );
  AND U6039 ( .A(n6601), .B(n6602), .Z(n6600) );
  XOR U6040 ( .A(n6599), .B(n6229), .Z(n6602) );
  XOR U6041 ( .A(n6603), .B(n6604), .Z(n6229) );
  AND U6042 ( .A(n451), .B(n6605), .Z(n6604) );
  XOR U6043 ( .A(n6606), .B(n6603), .Z(n6605) );
  XNOR U6044 ( .A(n6226), .B(n6599), .Z(n6601) );
  XOR U6045 ( .A(n6607), .B(n6608), .Z(n6226) );
  AND U6046 ( .A(n449), .B(n6609), .Z(n6608) );
  XOR U6047 ( .A(n6610), .B(n6607), .Z(n6609) );
  XOR U6048 ( .A(n6611), .B(n6612), .Z(n6599) );
  AND U6049 ( .A(n6613), .B(n6614), .Z(n6612) );
  XOR U6050 ( .A(n6611), .B(n6241), .Z(n6614) );
  XOR U6051 ( .A(n6615), .B(n6616), .Z(n6241) );
  AND U6052 ( .A(n451), .B(n6617), .Z(n6616) );
  XOR U6053 ( .A(n6618), .B(n6615), .Z(n6617) );
  XNOR U6054 ( .A(n6238), .B(n6611), .Z(n6613) );
  XOR U6055 ( .A(n6619), .B(n6620), .Z(n6238) );
  AND U6056 ( .A(n449), .B(n6621), .Z(n6620) );
  XOR U6057 ( .A(n6622), .B(n6619), .Z(n6621) );
  XOR U6058 ( .A(n6623), .B(n6624), .Z(n6611) );
  AND U6059 ( .A(n6625), .B(n6626), .Z(n6624) );
  XOR U6060 ( .A(n6623), .B(n6253), .Z(n6626) );
  XOR U6061 ( .A(n6627), .B(n6628), .Z(n6253) );
  AND U6062 ( .A(n451), .B(n6629), .Z(n6628) );
  XOR U6063 ( .A(n6630), .B(n6627), .Z(n6629) );
  XNOR U6064 ( .A(n6250), .B(n6623), .Z(n6625) );
  XOR U6065 ( .A(n6631), .B(n6632), .Z(n6250) );
  AND U6066 ( .A(n449), .B(n6633), .Z(n6632) );
  XOR U6067 ( .A(n6634), .B(n6631), .Z(n6633) );
  XOR U6068 ( .A(n6635), .B(n6636), .Z(n6623) );
  AND U6069 ( .A(n6637), .B(n6638), .Z(n6636) );
  XOR U6070 ( .A(n6635), .B(n6265), .Z(n6638) );
  XOR U6071 ( .A(n6639), .B(n6640), .Z(n6265) );
  AND U6072 ( .A(n451), .B(n6641), .Z(n6640) );
  XOR U6073 ( .A(n6642), .B(n6639), .Z(n6641) );
  XNOR U6074 ( .A(n6262), .B(n6635), .Z(n6637) );
  XOR U6075 ( .A(n6643), .B(n6644), .Z(n6262) );
  AND U6076 ( .A(n449), .B(n6645), .Z(n6644) );
  XOR U6077 ( .A(n6646), .B(n6643), .Z(n6645) );
  XOR U6078 ( .A(n6647), .B(n6648), .Z(n6635) );
  AND U6079 ( .A(n6649), .B(n6650), .Z(n6648) );
  XOR U6080 ( .A(n6647), .B(n6277), .Z(n6650) );
  XOR U6081 ( .A(n6651), .B(n6652), .Z(n6277) );
  AND U6082 ( .A(n451), .B(n6653), .Z(n6652) );
  XOR U6083 ( .A(n6654), .B(n6651), .Z(n6653) );
  XNOR U6084 ( .A(n6274), .B(n6647), .Z(n6649) );
  XOR U6085 ( .A(n6655), .B(n6656), .Z(n6274) );
  AND U6086 ( .A(n449), .B(n6657), .Z(n6656) );
  XOR U6087 ( .A(n6658), .B(n6655), .Z(n6657) );
  XOR U6088 ( .A(n6659), .B(n6660), .Z(n6647) );
  AND U6089 ( .A(n6661), .B(n6662), .Z(n6660) );
  XNOR U6090 ( .A(n6663), .B(n6290), .Z(n6662) );
  XOR U6091 ( .A(n6664), .B(n6665), .Z(n6290) );
  AND U6092 ( .A(n451), .B(n6666), .Z(n6665) );
  XOR U6093 ( .A(n6664), .B(n6667), .Z(n6666) );
  XNOR U6094 ( .A(n6287), .B(n6659), .Z(n6661) );
  XOR U6095 ( .A(n6668), .B(n6669), .Z(n6287) );
  AND U6096 ( .A(n449), .B(n6670), .Z(n6669) );
  XOR U6097 ( .A(n6668), .B(n6671), .Z(n6670) );
  IV U6098 ( .A(n6663), .Z(n6659) );
  AND U6099 ( .A(n6295), .B(n6298), .Z(n6663) );
  XNOR U6100 ( .A(n6672), .B(n6673), .Z(n6298) );
  AND U6101 ( .A(n451), .B(n6674), .Z(n6673) );
  XNOR U6102 ( .A(n6675), .B(n6672), .Z(n6674) );
  XOR U6103 ( .A(n6676), .B(n6677), .Z(n451) );
  AND U6104 ( .A(n6678), .B(n6679), .Z(n6677) );
  XOR U6105 ( .A(n6306), .B(n6676), .Z(n6679) );
  IV U6106 ( .A(n6680), .Z(n6306) );
  AND U6107 ( .A(p_input[7679]), .B(p_input[7647]), .Z(n6680) );
  XOR U6108 ( .A(n6676), .B(n6303), .Z(n6678) );
  AND U6109 ( .A(p_input[7583]), .B(p_input[7615]), .Z(n6303) );
  XOR U6110 ( .A(n6681), .B(n6682), .Z(n6676) );
  AND U6111 ( .A(n6683), .B(n6684), .Z(n6682) );
  XOR U6112 ( .A(n6681), .B(n6318), .Z(n6684) );
  XNOR U6113 ( .A(p_input[7646]), .B(n6685), .Z(n6318) );
  AND U6114 ( .A(n215), .B(n6686), .Z(n6685) );
  XOR U6115 ( .A(p_input[7678]), .B(p_input[7646]), .Z(n6686) );
  XNOR U6116 ( .A(n6315), .B(n6681), .Z(n6683) );
  XOR U6117 ( .A(n6687), .B(n6688), .Z(n6315) );
  AND U6118 ( .A(n213), .B(n6689), .Z(n6688) );
  XOR U6119 ( .A(p_input[7614]), .B(p_input[7582]), .Z(n6689) );
  XOR U6120 ( .A(n6690), .B(n6691), .Z(n6681) );
  AND U6121 ( .A(n6692), .B(n6693), .Z(n6691) );
  XOR U6122 ( .A(n6690), .B(n6330), .Z(n6693) );
  XNOR U6123 ( .A(p_input[7645]), .B(n6694), .Z(n6330) );
  AND U6124 ( .A(n215), .B(n6695), .Z(n6694) );
  XOR U6125 ( .A(p_input[7677]), .B(p_input[7645]), .Z(n6695) );
  XNOR U6126 ( .A(n6327), .B(n6690), .Z(n6692) );
  XOR U6127 ( .A(n6696), .B(n6697), .Z(n6327) );
  AND U6128 ( .A(n213), .B(n6698), .Z(n6697) );
  XOR U6129 ( .A(p_input[7613]), .B(p_input[7581]), .Z(n6698) );
  XOR U6130 ( .A(n6699), .B(n6700), .Z(n6690) );
  AND U6131 ( .A(n6701), .B(n6702), .Z(n6700) );
  XOR U6132 ( .A(n6699), .B(n6342), .Z(n6702) );
  XNOR U6133 ( .A(p_input[7644]), .B(n6703), .Z(n6342) );
  AND U6134 ( .A(n215), .B(n6704), .Z(n6703) );
  XOR U6135 ( .A(p_input[7676]), .B(p_input[7644]), .Z(n6704) );
  XNOR U6136 ( .A(n6339), .B(n6699), .Z(n6701) );
  XOR U6137 ( .A(n6705), .B(n6706), .Z(n6339) );
  AND U6138 ( .A(n213), .B(n6707), .Z(n6706) );
  XOR U6139 ( .A(p_input[7612]), .B(p_input[7580]), .Z(n6707) );
  XOR U6140 ( .A(n6708), .B(n6709), .Z(n6699) );
  AND U6141 ( .A(n6710), .B(n6711), .Z(n6709) );
  XOR U6142 ( .A(n6708), .B(n6354), .Z(n6711) );
  XNOR U6143 ( .A(p_input[7643]), .B(n6712), .Z(n6354) );
  AND U6144 ( .A(n215), .B(n6713), .Z(n6712) );
  XOR U6145 ( .A(p_input[7675]), .B(p_input[7643]), .Z(n6713) );
  XNOR U6146 ( .A(n6351), .B(n6708), .Z(n6710) );
  XOR U6147 ( .A(n6714), .B(n6715), .Z(n6351) );
  AND U6148 ( .A(n213), .B(n6716), .Z(n6715) );
  XOR U6149 ( .A(p_input[7611]), .B(p_input[7579]), .Z(n6716) );
  XOR U6150 ( .A(n6717), .B(n6718), .Z(n6708) );
  AND U6151 ( .A(n6719), .B(n6720), .Z(n6718) );
  XOR U6152 ( .A(n6717), .B(n6366), .Z(n6720) );
  XNOR U6153 ( .A(p_input[7642]), .B(n6721), .Z(n6366) );
  AND U6154 ( .A(n215), .B(n6722), .Z(n6721) );
  XOR U6155 ( .A(p_input[7674]), .B(p_input[7642]), .Z(n6722) );
  XNOR U6156 ( .A(n6363), .B(n6717), .Z(n6719) );
  XOR U6157 ( .A(n6723), .B(n6724), .Z(n6363) );
  AND U6158 ( .A(n213), .B(n6725), .Z(n6724) );
  XOR U6159 ( .A(p_input[7610]), .B(p_input[7578]), .Z(n6725) );
  XOR U6160 ( .A(n6726), .B(n6727), .Z(n6717) );
  AND U6161 ( .A(n6728), .B(n6729), .Z(n6727) );
  XOR U6162 ( .A(n6726), .B(n6378), .Z(n6729) );
  XNOR U6163 ( .A(p_input[7641]), .B(n6730), .Z(n6378) );
  AND U6164 ( .A(n215), .B(n6731), .Z(n6730) );
  XOR U6165 ( .A(p_input[7673]), .B(p_input[7641]), .Z(n6731) );
  XNOR U6166 ( .A(n6375), .B(n6726), .Z(n6728) );
  XOR U6167 ( .A(n6732), .B(n6733), .Z(n6375) );
  AND U6168 ( .A(n213), .B(n6734), .Z(n6733) );
  XOR U6169 ( .A(p_input[7609]), .B(p_input[7577]), .Z(n6734) );
  XOR U6170 ( .A(n6735), .B(n6736), .Z(n6726) );
  AND U6171 ( .A(n6737), .B(n6738), .Z(n6736) );
  XOR U6172 ( .A(n6735), .B(n6390), .Z(n6738) );
  XNOR U6173 ( .A(p_input[7640]), .B(n6739), .Z(n6390) );
  AND U6174 ( .A(n215), .B(n6740), .Z(n6739) );
  XOR U6175 ( .A(p_input[7672]), .B(p_input[7640]), .Z(n6740) );
  XNOR U6176 ( .A(n6387), .B(n6735), .Z(n6737) );
  XOR U6177 ( .A(n6741), .B(n6742), .Z(n6387) );
  AND U6178 ( .A(n213), .B(n6743), .Z(n6742) );
  XOR U6179 ( .A(p_input[7608]), .B(p_input[7576]), .Z(n6743) );
  XOR U6180 ( .A(n6744), .B(n6745), .Z(n6735) );
  AND U6181 ( .A(n6746), .B(n6747), .Z(n6745) );
  XOR U6182 ( .A(n6744), .B(n6402), .Z(n6747) );
  XNOR U6183 ( .A(p_input[7639]), .B(n6748), .Z(n6402) );
  AND U6184 ( .A(n215), .B(n6749), .Z(n6748) );
  XOR U6185 ( .A(p_input[7671]), .B(p_input[7639]), .Z(n6749) );
  XNOR U6186 ( .A(n6399), .B(n6744), .Z(n6746) );
  XOR U6187 ( .A(n6750), .B(n6751), .Z(n6399) );
  AND U6188 ( .A(n213), .B(n6752), .Z(n6751) );
  XOR U6189 ( .A(p_input[7607]), .B(p_input[7575]), .Z(n6752) );
  XOR U6190 ( .A(n6753), .B(n6754), .Z(n6744) );
  AND U6191 ( .A(n6755), .B(n6756), .Z(n6754) );
  XOR U6192 ( .A(n6753), .B(n6414), .Z(n6756) );
  XNOR U6193 ( .A(p_input[7638]), .B(n6757), .Z(n6414) );
  AND U6194 ( .A(n215), .B(n6758), .Z(n6757) );
  XOR U6195 ( .A(p_input[7670]), .B(p_input[7638]), .Z(n6758) );
  XNOR U6196 ( .A(n6411), .B(n6753), .Z(n6755) );
  XOR U6197 ( .A(n6759), .B(n6760), .Z(n6411) );
  AND U6198 ( .A(n213), .B(n6761), .Z(n6760) );
  XOR U6199 ( .A(p_input[7606]), .B(p_input[7574]), .Z(n6761) );
  XOR U6200 ( .A(n6762), .B(n6763), .Z(n6753) );
  AND U6201 ( .A(n6764), .B(n6765), .Z(n6763) );
  XOR U6202 ( .A(n6762), .B(n6426), .Z(n6765) );
  XNOR U6203 ( .A(p_input[7637]), .B(n6766), .Z(n6426) );
  AND U6204 ( .A(n215), .B(n6767), .Z(n6766) );
  XOR U6205 ( .A(p_input[7669]), .B(p_input[7637]), .Z(n6767) );
  XNOR U6206 ( .A(n6423), .B(n6762), .Z(n6764) );
  XOR U6207 ( .A(n6768), .B(n6769), .Z(n6423) );
  AND U6208 ( .A(n213), .B(n6770), .Z(n6769) );
  XOR U6209 ( .A(p_input[7605]), .B(p_input[7573]), .Z(n6770) );
  XOR U6210 ( .A(n6771), .B(n6772), .Z(n6762) );
  AND U6211 ( .A(n6773), .B(n6774), .Z(n6772) );
  XOR U6212 ( .A(n6771), .B(n6438), .Z(n6774) );
  XNOR U6213 ( .A(p_input[7636]), .B(n6775), .Z(n6438) );
  AND U6214 ( .A(n215), .B(n6776), .Z(n6775) );
  XOR U6215 ( .A(p_input[7668]), .B(p_input[7636]), .Z(n6776) );
  XNOR U6216 ( .A(n6435), .B(n6771), .Z(n6773) );
  XOR U6217 ( .A(n6777), .B(n6778), .Z(n6435) );
  AND U6218 ( .A(n213), .B(n6779), .Z(n6778) );
  XOR U6219 ( .A(p_input[7604]), .B(p_input[7572]), .Z(n6779) );
  XOR U6220 ( .A(n6780), .B(n6781), .Z(n6771) );
  AND U6221 ( .A(n6782), .B(n6783), .Z(n6781) );
  XOR U6222 ( .A(n6780), .B(n6450), .Z(n6783) );
  XNOR U6223 ( .A(p_input[7635]), .B(n6784), .Z(n6450) );
  AND U6224 ( .A(n215), .B(n6785), .Z(n6784) );
  XOR U6225 ( .A(p_input[7667]), .B(p_input[7635]), .Z(n6785) );
  XNOR U6226 ( .A(n6447), .B(n6780), .Z(n6782) );
  XOR U6227 ( .A(n6786), .B(n6787), .Z(n6447) );
  AND U6228 ( .A(n213), .B(n6788), .Z(n6787) );
  XOR U6229 ( .A(p_input[7603]), .B(p_input[7571]), .Z(n6788) );
  XOR U6230 ( .A(n6789), .B(n6790), .Z(n6780) );
  AND U6231 ( .A(n6791), .B(n6792), .Z(n6790) );
  XOR U6232 ( .A(n6789), .B(n6462), .Z(n6792) );
  XNOR U6233 ( .A(p_input[7634]), .B(n6793), .Z(n6462) );
  AND U6234 ( .A(n215), .B(n6794), .Z(n6793) );
  XOR U6235 ( .A(p_input[7666]), .B(p_input[7634]), .Z(n6794) );
  XNOR U6236 ( .A(n6459), .B(n6789), .Z(n6791) );
  XOR U6237 ( .A(n6795), .B(n6796), .Z(n6459) );
  AND U6238 ( .A(n213), .B(n6797), .Z(n6796) );
  XOR U6239 ( .A(p_input[7602]), .B(p_input[7570]), .Z(n6797) );
  XOR U6240 ( .A(n6798), .B(n6799), .Z(n6789) );
  AND U6241 ( .A(n6800), .B(n6801), .Z(n6799) );
  XOR U6242 ( .A(n6798), .B(n6474), .Z(n6801) );
  XNOR U6243 ( .A(p_input[7633]), .B(n6802), .Z(n6474) );
  AND U6244 ( .A(n215), .B(n6803), .Z(n6802) );
  XOR U6245 ( .A(p_input[7665]), .B(p_input[7633]), .Z(n6803) );
  XNOR U6246 ( .A(n6471), .B(n6798), .Z(n6800) );
  XOR U6247 ( .A(n6804), .B(n6805), .Z(n6471) );
  AND U6248 ( .A(n213), .B(n6806), .Z(n6805) );
  XOR U6249 ( .A(p_input[7601]), .B(p_input[7569]), .Z(n6806) );
  XOR U6250 ( .A(n6807), .B(n6808), .Z(n6798) );
  AND U6251 ( .A(n6809), .B(n6810), .Z(n6808) );
  XOR U6252 ( .A(n6807), .B(n6486), .Z(n6810) );
  XNOR U6253 ( .A(p_input[7632]), .B(n6811), .Z(n6486) );
  AND U6254 ( .A(n215), .B(n6812), .Z(n6811) );
  XOR U6255 ( .A(p_input[7664]), .B(p_input[7632]), .Z(n6812) );
  XNOR U6256 ( .A(n6483), .B(n6807), .Z(n6809) );
  XOR U6257 ( .A(n6813), .B(n6814), .Z(n6483) );
  AND U6258 ( .A(n213), .B(n6815), .Z(n6814) );
  XOR U6259 ( .A(p_input[7600]), .B(p_input[7568]), .Z(n6815) );
  XOR U6260 ( .A(n6816), .B(n6817), .Z(n6807) );
  AND U6261 ( .A(n6818), .B(n6819), .Z(n6817) );
  XOR U6262 ( .A(n6816), .B(n6498), .Z(n6819) );
  XNOR U6263 ( .A(p_input[7631]), .B(n6820), .Z(n6498) );
  AND U6264 ( .A(n215), .B(n6821), .Z(n6820) );
  XOR U6265 ( .A(p_input[7663]), .B(p_input[7631]), .Z(n6821) );
  XNOR U6266 ( .A(n6495), .B(n6816), .Z(n6818) );
  XOR U6267 ( .A(n6822), .B(n6823), .Z(n6495) );
  AND U6268 ( .A(n213), .B(n6824), .Z(n6823) );
  XOR U6269 ( .A(p_input[7599]), .B(p_input[7567]), .Z(n6824) );
  XOR U6270 ( .A(n6825), .B(n6826), .Z(n6816) );
  AND U6271 ( .A(n6827), .B(n6828), .Z(n6826) );
  XOR U6272 ( .A(n6825), .B(n6510), .Z(n6828) );
  XNOR U6273 ( .A(p_input[7630]), .B(n6829), .Z(n6510) );
  AND U6274 ( .A(n215), .B(n6830), .Z(n6829) );
  XOR U6275 ( .A(p_input[7662]), .B(p_input[7630]), .Z(n6830) );
  XNOR U6276 ( .A(n6507), .B(n6825), .Z(n6827) );
  XOR U6277 ( .A(n6831), .B(n6832), .Z(n6507) );
  AND U6278 ( .A(n213), .B(n6833), .Z(n6832) );
  XOR U6279 ( .A(p_input[7598]), .B(p_input[7566]), .Z(n6833) );
  XOR U6280 ( .A(n6834), .B(n6835), .Z(n6825) );
  AND U6281 ( .A(n6836), .B(n6837), .Z(n6835) );
  XOR U6282 ( .A(n6834), .B(n6522), .Z(n6837) );
  XNOR U6283 ( .A(p_input[7629]), .B(n6838), .Z(n6522) );
  AND U6284 ( .A(n215), .B(n6839), .Z(n6838) );
  XOR U6285 ( .A(p_input[7661]), .B(p_input[7629]), .Z(n6839) );
  XNOR U6286 ( .A(n6519), .B(n6834), .Z(n6836) );
  XOR U6287 ( .A(n6840), .B(n6841), .Z(n6519) );
  AND U6288 ( .A(n213), .B(n6842), .Z(n6841) );
  XOR U6289 ( .A(p_input[7597]), .B(p_input[7565]), .Z(n6842) );
  XOR U6290 ( .A(n6843), .B(n6844), .Z(n6834) );
  AND U6291 ( .A(n6845), .B(n6846), .Z(n6844) );
  XOR U6292 ( .A(n6843), .B(n6534), .Z(n6846) );
  XNOR U6293 ( .A(p_input[7628]), .B(n6847), .Z(n6534) );
  AND U6294 ( .A(n215), .B(n6848), .Z(n6847) );
  XOR U6295 ( .A(p_input[7660]), .B(p_input[7628]), .Z(n6848) );
  XNOR U6296 ( .A(n6531), .B(n6843), .Z(n6845) );
  XOR U6297 ( .A(n6849), .B(n6850), .Z(n6531) );
  AND U6298 ( .A(n213), .B(n6851), .Z(n6850) );
  XOR U6299 ( .A(p_input[7596]), .B(p_input[7564]), .Z(n6851) );
  XOR U6300 ( .A(n6852), .B(n6853), .Z(n6843) );
  AND U6301 ( .A(n6854), .B(n6855), .Z(n6853) );
  XOR U6302 ( .A(n6852), .B(n6546), .Z(n6855) );
  XNOR U6303 ( .A(p_input[7627]), .B(n6856), .Z(n6546) );
  AND U6304 ( .A(n215), .B(n6857), .Z(n6856) );
  XOR U6305 ( .A(p_input[7659]), .B(p_input[7627]), .Z(n6857) );
  XNOR U6306 ( .A(n6543), .B(n6852), .Z(n6854) );
  XOR U6307 ( .A(n6858), .B(n6859), .Z(n6543) );
  AND U6308 ( .A(n213), .B(n6860), .Z(n6859) );
  XOR U6309 ( .A(p_input[7595]), .B(p_input[7563]), .Z(n6860) );
  XOR U6310 ( .A(n6861), .B(n6862), .Z(n6852) );
  AND U6311 ( .A(n6863), .B(n6864), .Z(n6862) );
  XOR U6312 ( .A(n6861), .B(n6558), .Z(n6864) );
  XNOR U6313 ( .A(p_input[7626]), .B(n6865), .Z(n6558) );
  AND U6314 ( .A(n215), .B(n6866), .Z(n6865) );
  XOR U6315 ( .A(p_input[7658]), .B(p_input[7626]), .Z(n6866) );
  XNOR U6316 ( .A(n6555), .B(n6861), .Z(n6863) );
  XOR U6317 ( .A(n6867), .B(n6868), .Z(n6555) );
  AND U6318 ( .A(n213), .B(n6869), .Z(n6868) );
  XOR U6319 ( .A(p_input[7594]), .B(p_input[7562]), .Z(n6869) );
  XOR U6320 ( .A(n6870), .B(n6871), .Z(n6861) );
  AND U6321 ( .A(n6872), .B(n6873), .Z(n6871) );
  XOR U6322 ( .A(n6870), .B(n6570), .Z(n6873) );
  XNOR U6323 ( .A(p_input[7625]), .B(n6874), .Z(n6570) );
  AND U6324 ( .A(n215), .B(n6875), .Z(n6874) );
  XOR U6325 ( .A(p_input[7657]), .B(p_input[7625]), .Z(n6875) );
  XNOR U6326 ( .A(n6567), .B(n6870), .Z(n6872) );
  XOR U6327 ( .A(n6876), .B(n6877), .Z(n6567) );
  AND U6328 ( .A(n213), .B(n6878), .Z(n6877) );
  XOR U6329 ( .A(p_input[7593]), .B(p_input[7561]), .Z(n6878) );
  XOR U6330 ( .A(n6879), .B(n6880), .Z(n6870) );
  AND U6331 ( .A(n6881), .B(n6882), .Z(n6880) );
  XOR U6332 ( .A(n6879), .B(n6582), .Z(n6882) );
  XNOR U6333 ( .A(p_input[7624]), .B(n6883), .Z(n6582) );
  AND U6334 ( .A(n215), .B(n6884), .Z(n6883) );
  XOR U6335 ( .A(p_input[7656]), .B(p_input[7624]), .Z(n6884) );
  XNOR U6336 ( .A(n6579), .B(n6879), .Z(n6881) );
  XOR U6337 ( .A(n6885), .B(n6886), .Z(n6579) );
  AND U6338 ( .A(n213), .B(n6887), .Z(n6886) );
  XOR U6339 ( .A(p_input[7592]), .B(p_input[7560]), .Z(n6887) );
  XOR U6340 ( .A(n6888), .B(n6889), .Z(n6879) );
  AND U6341 ( .A(n6890), .B(n6891), .Z(n6889) );
  XOR U6342 ( .A(n6888), .B(n6594), .Z(n6891) );
  XNOR U6343 ( .A(p_input[7623]), .B(n6892), .Z(n6594) );
  AND U6344 ( .A(n215), .B(n6893), .Z(n6892) );
  XOR U6345 ( .A(p_input[7655]), .B(p_input[7623]), .Z(n6893) );
  XNOR U6346 ( .A(n6591), .B(n6888), .Z(n6890) );
  XOR U6347 ( .A(n6894), .B(n6895), .Z(n6591) );
  AND U6348 ( .A(n213), .B(n6896), .Z(n6895) );
  XOR U6349 ( .A(p_input[7591]), .B(p_input[7559]), .Z(n6896) );
  XOR U6350 ( .A(n6897), .B(n6898), .Z(n6888) );
  AND U6351 ( .A(n6899), .B(n6900), .Z(n6898) );
  XOR U6352 ( .A(n6897), .B(n6606), .Z(n6900) );
  XNOR U6353 ( .A(p_input[7622]), .B(n6901), .Z(n6606) );
  AND U6354 ( .A(n215), .B(n6902), .Z(n6901) );
  XOR U6355 ( .A(p_input[7654]), .B(p_input[7622]), .Z(n6902) );
  XNOR U6356 ( .A(n6603), .B(n6897), .Z(n6899) );
  XOR U6357 ( .A(n6903), .B(n6904), .Z(n6603) );
  AND U6358 ( .A(n213), .B(n6905), .Z(n6904) );
  XOR U6359 ( .A(p_input[7590]), .B(p_input[7558]), .Z(n6905) );
  XOR U6360 ( .A(n6906), .B(n6907), .Z(n6897) );
  AND U6361 ( .A(n6908), .B(n6909), .Z(n6907) );
  XOR U6362 ( .A(n6906), .B(n6618), .Z(n6909) );
  XNOR U6363 ( .A(p_input[7621]), .B(n6910), .Z(n6618) );
  AND U6364 ( .A(n215), .B(n6911), .Z(n6910) );
  XOR U6365 ( .A(p_input[7653]), .B(p_input[7621]), .Z(n6911) );
  XNOR U6366 ( .A(n6615), .B(n6906), .Z(n6908) );
  XOR U6367 ( .A(n6912), .B(n6913), .Z(n6615) );
  AND U6368 ( .A(n213), .B(n6914), .Z(n6913) );
  XOR U6369 ( .A(p_input[7589]), .B(p_input[7557]), .Z(n6914) );
  XOR U6370 ( .A(n6915), .B(n6916), .Z(n6906) );
  AND U6371 ( .A(n6917), .B(n6918), .Z(n6916) );
  XOR U6372 ( .A(n6915), .B(n6630), .Z(n6918) );
  XNOR U6373 ( .A(p_input[7620]), .B(n6919), .Z(n6630) );
  AND U6374 ( .A(n215), .B(n6920), .Z(n6919) );
  XOR U6375 ( .A(p_input[7652]), .B(p_input[7620]), .Z(n6920) );
  XNOR U6376 ( .A(n6627), .B(n6915), .Z(n6917) );
  XOR U6377 ( .A(n6921), .B(n6922), .Z(n6627) );
  AND U6378 ( .A(n213), .B(n6923), .Z(n6922) );
  XOR U6379 ( .A(p_input[7588]), .B(p_input[7556]), .Z(n6923) );
  XOR U6380 ( .A(n6924), .B(n6925), .Z(n6915) );
  AND U6381 ( .A(n6926), .B(n6927), .Z(n6925) );
  XOR U6382 ( .A(n6924), .B(n6642), .Z(n6927) );
  XNOR U6383 ( .A(p_input[7619]), .B(n6928), .Z(n6642) );
  AND U6384 ( .A(n215), .B(n6929), .Z(n6928) );
  XOR U6385 ( .A(p_input[7651]), .B(p_input[7619]), .Z(n6929) );
  XNOR U6386 ( .A(n6639), .B(n6924), .Z(n6926) );
  XOR U6387 ( .A(n6930), .B(n6931), .Z(n6639) );
  AND U6388 ( .A(n213), .B(n6932), .Z(n6931) );
  XOR U6389 ( .A(p_input[7587]), .B(p_input[7555]), .Z(n6932) );
  XOR U6390 ( .A(n6933), .B(n6934), .Z(n6924) );
  AND U6391 ( .A(n6935), .B(n6936), .Z(n6934) );
  XOR U6392 ( .A(n6933), .B(n6654), .Z(n6936) );
  XNOR U6393 ( .A(p_input[7618]), .B(n6937), .Z(n6654) );
  AND U6394 ( .A(n215), .B(n6938), .Z(n6937) );
  XOR U6395 ( .A(p_input[7650]), .B(p_input[7618]), .Z(n6938) );
  XNOR U6396 ( .A(n6651), .B(n6933), .Z(n6935) );
  XOR U6397 ( .A(n6939), .B(n6940), .Z(n6651) );
  AND U6398 ( .A(n213), .B(n6941), .Z(n6940) );
  XOR U6399 ( .A(p_input[7586]), .B(p_input[7554]), .Z(n6941) );
  XOR U6400 ( .A(n6942), .B(n6943), .Z(n6933) );
  AND U6401 ( .A(n6944), .B(n6945), .Z(n6943) );
  XNOR U6402 ( .A(n6946), .B(n6667), .Z(n6945) );
  XNOR U6403 ( .A(p_input[7617]), .B(n6947), .Z(n6667) );
  AND U6404 ( .A(n215), .B(n6948), .Z(n6947) );
  XNOR U6405 ( .A(p_input[7649]), .B(n6949), .Z(n6948) );
  IV U6406 ( .A(p_input[7617]), .Z(n6949) );
  XNOR U6407 ( .A(n6664), .B(n6942), .Z(n6944) );
  XNOR U6408 ( .A(p_input[7553]), .B(n6950), .Z(n6664) );
  AND U6409 ( .A(n213), .B(n6951), .Z(n6950) );
  XOR U6410 ( .A(p_input[7585]), .B(p_input[7553]), .Z(n6951) );
  IV U6411 ( .A(n6946), .Z(n6942) );
  AND U6412 ( .A(n6672), .B(n6675), .Z(n6946) );
  XOR U6413 ( .A(p_input[7616]), .B(n6952), .Z(n6675) );
  AND U6414 ( .A(n215), .B(n6953), .Z(n6952) );
  XOR U6415 ( .A(p_input[7648]), .B(p_input[7616]), .Z(n6953) );
  XOR U6416 ( .A(n6954), .B(n6955), .Z(n215) );
  AND U6417 ( .A(n6956), .B(n6957), .Z(n6955) );
  XNOR U6418 ( .A(p_input[7679]), .B(n6954), .Z(n6957) );
  XOR U6419 ( .A(n6954), .B(p_input[7647]), .Z(n6956) );
  XOR U6420 ( .A(n6958), .B(n6959), .Z(n6954) );
  AND U6421 ( .A(n6960), .B(n6961), .Z(n6959) );
  XNOR U6422 ( .A(p_input[7678]), .B(n6958), .Z(n6961) );
  XOR U6423 ( .A(n6958), .B(p_input[7646]), .Z(n6960) );
  XOR U6424 ( .A(n6962), .B(n6963), .Z(n6958) );
  AND U6425 ( .A(n6964), .B(n6965), .Z(n6963) );
  XNOR U6426 ( .A(p_input[7677]), .B(n6962), .Z(n6965) );
  XOR U6427 ( .A(n6962), .B(p_input[7645]), .Z(n6964) );
  XOR U6428 ( .A(n6966), .B(n6967), .Z(n6962) );
  AND U6429 ( .A(n6968), .B(n6969), .Z(n6967) );
  XNOR U6430 ( .A(p_input[7676]), .B(n6966), .Z(n6969) );
  XOR U6431 ( .A(n6966), .B(p_input[7644]), .Z(n6968) );
  XOR U6432 ( .A(n6970), .B(n6971), .Z(n6966) );
  AND U6433 ( .A(n6972), .B(n6973), .Z(n6971) );
  XNOR U6434 ( .A(p_input[7675]), .B(n6970), .Z(n6973) );
  XOR U6435 ( .A(n6970), .B(p_input[7643]), .Z(n6972) );
  XOR U6436 ( .A(n6974), .B(n6975), .Z(n6970) );
  AND U6437 ( .A(n6976), .B(n6977), .Z(n6975) );
  XNOR U6438 ( .A(p_input[7674]), .B(n6974), .Z(n6977) );
  XOR U6439 ( .A(n6974), .B(p_input[7642]), .Z(n6976) );
  XOR U6440 ( .A(n6978), .B(n6979), .Z(n6974) );
  AND U6441 ( .A(n6980), .B(n6981), .Z(n6979) );
  XNOR U6442 ( .A(p_input[7673]), .B(n6978), .Z(n6981) );
  XOR U6443 ( .A(n6978), .B(p_input[7641]), .Z(n6980) );
  XOR U6444 ( .A(n6982), .B(n6983), .Z(n6978) );
  AND U6445 ( .A(n6984), .B(n6985), .Z(n6983) );
  XNOR U6446 ( .A(p_input[7672]), .B(n6982), .Z(n6985) );
  XOR U6447 ( .A(n6982), .B(p_input[7640]), .Z(n6984) );
  XOR U6448 ( .A(n6986), .B(n6987), .Z(n6982) );
  AND U6449 ( .A(n6988), .B(n6989), .Z(n6987) );
  XNOR U6450 ( .A(p_input[7671]), .B(n6986), .Z(n6989) );
  XOR U6451 ( .A(n6986), .B(p_input[7639]), .Z(n6988) );
  XOR U6452 ( .A(n6990), .B(n6991), .Z(n6986) );
  AND U6453 ( .A(n6992), .B(n6993), .Z(n6991) );
  XNOR U6454 ( .A(p_input[7670]), .B(n6990), .Z(n6993) );
  XOR U6455 ( .A(n6990), .B(p_input[7638]), .Z(n6992) );
  XOR U6456 ( .A(n6994), .B(n6995), .Z(n6990) );
  AND U6457 ( .A(n6996), .B(n6997), .Z(n6995) );
  XNOR U6458 ( .A(p_input[7669]), .B(n6994), .Z(n6997) );
  XOR U6459 ( .A(n6994), .B(p_input[7637]), .Z(n6996) );
  XOR U6460 ( .A(n6998), .B(n6999), .Z(n6994) );
  AND U6461 ( .A(n7000), .B(n7001), .Z(n6999) );
  XNOR U6462 ( .A(p_input[7668]), .B(n6998), .Z(n7001) );
  XOR U6463 ( .A(n6998), .B(p_input[7636]), .Z(n7000) );
  XOR U6464 ( .A(n7002), .B(n7003), .Z(n6998) );
  AND U6465 ( .A(n7004), .B(n7005), .Z(n7003) );
  XNOR U6466 ( .A(p_input[7667]), .B(n7002), .Z(n7005) );
  XOR U6467 ( .A(n7002), .B(p_input[7635]), .Z(n7004) );
  XOR U6468 ( .A(n7006), .B(n7007), .Z(n7002) );
  AND U6469 ( .A(n7008), .B(n7009), .Z(n7007) );
  XNOR U6470 ( .A(p_input[7666]), .B(n7006), .Z(n7009) );
  XOR U6471 ( .A(n7006), .B(p_input[7634]), .Z(n7008) );
  XOR U6472 ( .A(n7010), .B(n7011), .Z(n7006) );
  AND U6473 ( .A(n7012), .B(n7013), .Z(n7011) );
  XNOR U6474 ( .A(p_input[7665]), .B(n7010), .Z(n7013) );
  XOR U6475 ( .A(n7010), .B(p_input[7633]), .Z(n7012) );
  XOR U6476 ( .A(n7014), .B(n7015), .Z(n7010) );
  AND U6477 ( .A(n7016), .B(n7017), .Z(n7015) );
  XNOR U6478 ( .A(p_input[7664]), .B(n7014), .Z(n7017) );
  XOR U6479 ( .A(n7014), .B(p_input[7632]), .Z(n7016) );
  XOR U6480 ( .A(n7018), .B(n7019), .Z(n7014) );
  AND U6481 ( .A(n7020), .B(n7021), .Z(n7019) );
  XNOR U6482 ( .A(p_input[7663]), .B(n7018), .Z(n7021) );
  XOR U6483 ( .A(n7018), .B(p_input[7631]), .Z(n7020) );
  XOR U6484 ( .A(n7022), .B(n7023), .Z(n7018) );
  AND U6485 ( .A(n7024), .B(n7025), .Z(n7023) );
  XNOR U6486 ( .A(p_input[7662]), .B(n7022), .Z(n7025) );
  XOR U6487 ( .A(n7022), .B(p_input[7630]), .Z(n7024) );
  XOR U6488 ( .A(n7026), .B(n7027), .Z(n7022) );
  AND U6489 ( .A(n7028), .B(n7029), .Z(n7027) );
  XNOR U6490 ( .A(p_input[7661]), .B(n7026), .Z(n7029) );
  XOR U6491 ( .A(n7026), .B(p_input[7629]), .Z(n7028) );
  XOR U6492 ( .A(n7030), .B(n7031), .Z(n7026) );
  AND U6493 ( .A(n7032), .B(n7033), .Z(n7031) );
  XNOR U6494 ( .A(p_input[7660]), .B(n7030), .Z(n7033) );
  XOR U6495 ( .A(n7030), .B(p_input[7628]), .Z(n7032) );
  XOR U6496 ( .A(n7034), .B(n7035), .Z(n7030) );
  AND U6497 ( .A(n7036), .B(n7037), .Z(n7035) );
  XNOR U6498 ( .A(p_input[7659]), .B(n7034), .Z(n7037) );
  XOR U6499 ( .A(n7034), .B(p_input[7627]), .Z(n7036) );
  XOR U6500 ( .A(n7038), .B(n7039), .Z(n7034) );
  AND U6501 ( .A(n7040), .B(n7041), .Z(n7039) );
  XNOR U6502 ( .A(p_input[7658]), .B(n7038), .Z(n7041) );
  XOR U6503 ( .A(n7038), .B(p_input[7626]), .Z(n7040) );
  XOR U6504 ( .A(n7042), .B(n7043), .Z(n7038) );
  AND U6505 ( .A(n7044), .B(n7045), .Z(n7043) );
  XNOR U6506 ( .A(p_input[7657]), .B(n7042), .Z(n7045) );
  XOR U6507 ( .A(n7042), .B(p_input[7625]), .Z(n7044) );
  XOR U6508 ( .A(n7046), .B(n7047), .Z(n7042) );
  AND U6509 ( .A(n7048), .B(n7049), .Z(n7047) );
  XNOR U6510 ( .A(p_input[7656]), .B(n7046), .Z(n7049) );
  XOR U6511 ( .A(n7046), .B(p_input[7624]), .Z(n7048) );
  XOR U6512 ( .A(n7050), .B(n7051), .Z(n7046) );
  AND U6513 ( .A(n7052), .B(n7053), .Z(n7051) );
  XNOR U6514 ( .A(p_input[7655]), .B(n7050), .Z(n7053) );
  XOR U6515 ( .A(n7050), .B(p_input[7623]), .Z(n7052) );
  XOR U6516 ( .A(n7054), .B(n7055), .Z(n7050) );
  AND U6517 ( .A(n7056), .B(n7057), .Z(n7055) );
  XNOR U6518 ( .A(p_input[7654]), .B(n7054), .Z(n7057) );
  XOR U6519 ( .A(n7054), .B(p_input[7622]), .Z(n7056) );
  XOR U6520 ( .A(n7058), .B(n7059), .Z(n7054) );
  AND U6521 ( .A(n7060), .B(n7061), .Z(n7059) );
  XNOR U6522 ( .A(p_input[7653]), .B(n7058), .Z(n7061) );
  XOR U6523 ( .A(n7058), .B(p_input[7621]), .Z(n7060) );
  XOR U6524 ( .A(n7062), .B(n7063), .Z(n7058) );
  AND U6525 ( .A(n7064), .B(n7065), .Z(n7063) );
  XNOR U6526 ( .A(p_input[7652]), .B(n7062), .Z(n7065) );
  XOR U6527 ( .A(n7062), .B(p_input[7620]), .Z(n7064) );
  XOR U6528 ( .A(n7066), .B(n7067), .Z(n7062) );
  AND U6529 ( .A(n7068), .B(n7069), .Z(n7067) );
  XNOR U6530 ( .A(p_input[7651]), .B(n7066), .Z(n7069) );
  XOR U6531 ( .A(n7066), .B(p_input[7619]), .Z(n7068) );
  XOR U6532 ( .A(n7070), .B(n7071), .Z(n7066) );
  AND U6533 ( .A(n7072), .B(n7073), .Z(n7071) );
  XNOR U6534 ( .A(p_input[7650]), .B(n7070), .Z(n7073) );
  XOR U6535 ( .A(n7070), .B(p_input[7618]), .Z(n7072) );
  XNOR U6536 ( .A(n7074), .B(n7075), .Z(n7070) );
  AND U6537 ( .A(n7076), .B(n7077), .Z(n7075) );
  XOR U6538 ( .A(p_input[7649]), .B(n7074), .Z(n7077) );
  XNOR U6539 ( .A(p_input[7617]), .B(n7074), .Z(n7076) );
  AND U6540 ( .A(p_input[7648]), .B(n7078), .Z(n7074) );
  IV U6541 ( .A(p_input[7616]), .Z(n7078) );
  XNOR U6542 ( .A(p_input[7552]), .B(n7079), .Z(n6672) );
  AND U6543 ( .A(n213), .B(n7080), .Z(n7079) );
  XOR U6544 ( .A(p_input[7584]), .B(p_input[7552]), .Z(n7080) );
  XOR U6545 ( .A(n7081), .B(n7082), .Z(n213) );
  AND U6546 ( .A(n7083), .B(n7084), .Z(n7082) );
  XNOR U6547 ( .A(p_input[7615]), .B(n7081), .Z(n7084) );
  XOR U6548 ( .A(n7081), .B(p_input[7583]), .Z(n7083) );
  XOR U6549 ( .A(n7085), .B(n7086), .Z(n7081) );
  AND U6550 ( .A(n7087), .B(n7088), .Z(n7086) );
  XNOR U6551 ( .A(p_input[7614]), .B(n7085), .Z(n7088) );
  XNOR U6552 ( .A(n7085), .B(n6687), .Z(n7087) );
  IV U6553 ( .A(p_input[7582]), .Z(n6687) );
  XOR U6554 ( .A(n7089), .B(n7090), .Z(n7085) );
  AND U6555 ( .A(n7091), .B(n7092), .Z(n7090) );
  XNOR U6556 ( .A(p_input[7613]), .B(n7089), .Z(n7092) );
  XNOR U6557 ( .A(n7089), .B(n6696), .Z(n7091) );
  IV U6558 ( .A(p_input[7581]), .Z(n6696) );
  XOR U6559 ( .A(n7093), .B(n7094), .Z(n7089) );
  AND U6560 ( .A(n7095), .B(n7096), .Z(n7094) );
  XNOR U6561 ( .A(p_input[7612]), .B(n7093), .Z(n7096) );
  XNOR U6562 ( .A(n7093), .B(n6705), .Z(n7095) );
  IV U6563 ( .A(p_input[7580]), .Z(n6705) );
  XOR U6564 ( .A(n7097), .B(n7098), .Z(n7093) );
  AND U6565 ( .A(n7099), .B(n7100), .Z(n7098) );
  XNOR U6566 ( .A(p_input[7611]), .B(n7097), .Z(n7100) );
  XNOR U6567 ( .A(n7097), .B(n6714), .Z(n7099) );
  IV U6568 ( .A(p_input[7579]), .Z(n6714) );
  XOR U6569 ( .A(n7101), .B(n7102), .Z(n7097) );
  AND U6570 ( .A(n7103), .B(n7104), .Z(n7102) );
  XNOR U6571 ( .A(p_input[7610]), .B(n7101), .Z(n7104) );
  XNOR U6572 ( .A(n7101), .B(n6723), .Z(n7103) );
  IV U6573 ( .A(p_input[7578]), .Z(n6723) );
  XOR U6574 ( .A(n7105), .B(n7106), .Z(n7101) );
  AND U6575 ( .A(n7107), .B(n7108), .Z(n7106) );
  XNOR U6576 ( .A(p_input[7609]), .B(n7105), .Z(n7108) );
  XNOR U6577 ( .A(n7105), .B(n6732), .Z(n7107) );
  IV U6578 ( .A(p_input[7577]), .Z(n6732) );
  XOR U6579 ( .A(n7109), .B(n7110), .Z(n7105) );
  AND U6580 ( .A(n7111), .B(n7112), .Z(n7110) );
  XNOR U6581 ( .A(p_input[7608]), .B(n7109), .Z(n7112) );
  XNOR U6582 ( .A(n7109), .B(n6741), .Z(n7111) );
  IV U6583 ( .A(p_input[7576]), .Z(n6741) );
  XOR U6584 ( .A(n7113), .B(n7114), .Z(n7109) );
  AND U6585 ( .A(n7115), .B(n7116), .Z(n7114) );
  XNOR U6586 ( .A(p_input[7607]), .B(n7113), .Z(n7116) );
  XNOR U6587 ( .A(n7113), .B(n6750), .Z(n7115) );
  IV U6588 ( .A(p_input[7575]), .Z(n6750) );
  XOR U6589 ( .A(n7117), .B(n7118), .Z(n7113) );
  AND U6590 ( .A(n7119), .B(n7120), .Z(n7118) );
  XNOR U6591 ( .A(p_input[7606]), .B(n7117), .Z(n7120) );
  XNOR U6592 ( .A(n7117), .B(n6759), .Z(n7119) );
  IV U6593 ( .A(p_input[7574]), .Z(n6759) );
  XOR U6594 ( .A(n7121), .B(n7122), .Z(n7117) );
  AND U6595 ( .A(n7123), .B(n7124), .Z(n7122) );
  XNOR U6596 ( .A(p_input[7605]), .B(n7121), .Z(n7124) );
  XNOR U6597 ( .A(n7121), .B(n6768), .Z(n7123) );
  IV U6598 ( .A(p_input[7573]), .Z(n6768) );
  XOR U6599 ( .A(n7125), .B(n7126), .Z(n7121) );
  AND U6600 ( .A(n7127), .B(n7128), .Z(n7126) );
  XNOR U6601 ( .A(p_input[7604]), .B(n7125), .Z(n7128) );
  XNOR U6602 ( .A(n7125), .B(n6777), .Z(n7127) );
  IV U6603 ( .A(p_input[7572]), .Z(n6777) );
  XOR U6604 ( .A(n7129), .B(n7130), .Z(n7125) );
  AND U6605 ( .A(n7131), .B(n7132), .Z(n7130) );
  XNOR U6606 ( .A(p_input[7603]), .B(n7129), .Z(n7132) );
  XNOR U6607 ( .A(n7129), .B(n6786), .Z(n7131) );
  IV U6608 ( .A(p_input[7571]), .Z(n6786) );
  XOR U6609 ( .A(n7133), .B(n7134), .Z(n7129) );
  AND U6610 ( .A(n7135), .B(n7136), .Z(n7134) );
  XNOR U6611 ( .A(p_input[7602]), .B(n7133), .Z(n7136) );
  XNOR U6612 ( .A(n7133), .B(n6795), .Z(n7135) );
  IV U6613 ( .A(p_input[7570]), .Z(n6795) );
  XOR U6614 ( .A(n7137), .B(n7138), .Z(n7133) );
  AND U6615 ( .A(n7139), .B(n7140), .Z(n7138) );
  XNOR U6616 ( .A(p_input[7601]), .B(n7137), .Z(n7140) );
  XNOR U6617 ( .A(n7137), .B(n6804), .Z(n7139) );
  IV U6618 ( .A(p_input[7569]), .Z(n6804) );
  XOR U6619 ( .A(n7141), .B(n7142), .Z(n7137) );
  AND U6620 ( .A(n7143), .B(n7144), .Z(n7142) );
  XNOR U6621 ( .A(p_input[7600]), .B(n7141), .Z(n7144) );
  XNOR U6622 ( .A(n7141), .B(n6813), .Z(n7143) );
  IV U6623 ( .A(p_input[7568]), .Z(n6813) );
  XOR U6624 ( .A(n7145), .B(n7146), .Z(n7141) );
  AND U6625 ( .A(n7147), .B(n7148), .Z(n7146) );
  XNOR U6626 ( .A(p_input[7599]), .B(n7145), .Z(n7148) );
  XNOR U6627 ( .A(n7145), .B(n6822), .Z(n7147) );
  IV U6628 ( .A(p_input[7567]), .Z(n6822) );
  XOR U6629 ( .A(n7149), .B(n7150), .Z(n7145) );
  AND U6630 ( .A(n7151), .B(n7152), .Z(n7150) );
  XNOR U6631 ( .A(p_input[7598]), .B(n7149), .Z(n7152) );
  XNOR U6632 ( .A(n7149), .B(n6831), .Z(n7151) );
  IV U6633 ( .A(p_input[7566]), .Z(n6831) );
  XOR U6634 ( .A(n7153), .B(n7154), .Z(n7149) );
  AND U6635 ( .A(n7155), .B(n7156), .Z(n7154) );
  XNOR U6636 ( .A(p_input[7597]), .B(n7153), .Z(n7156) );
  XNOR U6637 ( .A(n7153), .B(n6840), .Z(n7155) );
  IV U6638 ( .A(p_input[7565]), .Z(n6840) );
  XOR U6639 ( .A(n7157), .B(n7158), .Z(n7153) );
  AND U6640 ( .A(n7159), .B(n7160), .Z(n7158) );
  XNOR U6641 ( .A(p_input[7596]), .B(n7157), .Z(n7160) );
  XNOR U6642 ( .A(n7157), .B(n6849), .Z(n7159) );
  IV U6643 ( .A(p_input[7564]), .Z(n6849) );
  XOR U6644 ( .A(n7161), .B(n7162), .Z(n7157) );
  AND U6645 ( .A(n7163), .B(n7164), .Z(n7162) );
  XNOR U6646 ( .A(p_input[7595]), .B(n7161), .Z(n7164) );
  XNOR U6647 ( .A(n7161), .B(n6858), .Z(n7163) );
  IV U6648 ( .A(p_input[7563]), .Z(n6858) );
  XOR U6649 ( .A(n7165), .B(n7166), .Z(n7161) );
  AND U6650 ( .A(n7167), .B(n7168), .Z(n7166) );
  XNOR U6651 ( .A(p_input[7594]), .B(n7165), .Z(n7168) );
  XNOR U6652 ( .A(n7165), .B(n6867), .Z(n7167) );
  IV U6653 ( .A(p_input[7562]), .Z(n6867) );
  XOR U6654 ( .A(n7169), .B(n7170), .Z(n7165) );
  AND U6655 ( .A(n7171), .B(n7172), .Z(n7170) );
  XNOR U6656 ( .A(p_input[7593]), .B(n7169), .Z(n7172) );
  XNOR U6657 ( .A(n7169), .B(n6876), .Z(n7171) );
  IV U6658 ( .A(p_input[7561]), .Z(n6876) );
  XOR U6659 ( .A(n7173), .B(n7174), .Z(n7169) );
  AND U6660 ( .A(n7175), .B(n7176), .Z(n7174) );
  XNOR U6661 ( .A(p_input[7592]), .B(n7173), .Z(n7176) );
  XNOR U6662 ( .A(n7173), .B(n6885), .Z(n7175) );
  IV U6663 ( .A(p_input[7560]), .Z(n6885) );
  XOR U6664 ( .A(n7177), .B(n7178), .Z(n7173) );
  AND U6665 ( .A(n7179), .B(n7180), .Z(n7178) );
  XNOR U6666 ( .A(p_input[7591]), .B(n7177), .Z(n7180) );
  XNOR U6667 ( .A(n7177), .B(n6894), .Z(n7179) );
  IV U6668 ( .A(p_input[7559]), .Z(n6894) );
  XOR U6669 ( .A(n7181), .B(n7182), .Z(n7177) );
  AND U6670 ( .A(n7183), .B(n7184), .Z(n7182) );
  XNOR U6671 ( .A(p_input[7590]), .B(n7181), .Z(n7184) );
  XNOR U6672 ( .A(n7181), .B(n6903), .Z(n7183) );
  IV U6673 ( .A(p_input[7558]), .Z(n6903) );
  XOR U6674 ( .A(n7185), .B(n7186), .Z(n7181) );
  AND U6675 ( .A(n7187), .B(n7188), .Z(n7186) );
  XNOR U6676 ( .A(p_input[7589]), .B(n7185), .Z(n7188) );
  XNOR U6677 ( .A(n7185), .B(n6912), .Z(n7187) );
  IV U6678 ( .A(p_input[7557]), .Z(n6912) );
  XOR U6679 ( .A(n7189), .B(n7190), .Z(n7185) );
  AND U6680 ( .A(n7191), .B(n7192), .Z(n7190) );
  XNOR U6681 ( .A(p_input[7588]), .B(n7189), .Z(n7192) );
  XNOR U6682 ( .A(n7189), .B(n6921), .Z(n7191) );
  IV U6683 ( .A(p_input[7556]), .Z(n6921) );
  XOR U6684 ( .A(n7193), .B(n7194), .Z(n7189) );
  AND U6685 ( .A(n7195), .B(n7196), .Z(n7194) );
  XNOR U6686 ( .A(p_input[7587]), .B(n7193), .Z(n7196) );
  XNOR U6687 ( .A(n7193), .B(n6930), .Z(n7195) );
  IV U6688 ( .A(p_input[7555]), .Z(n6930) );
  XOR U6689 ( .A(n7197), .B(n7198), .Z(n7193) );
  AND U6690 ( .A(n7199), .B(n7200), .Z(n7198) );
  XNOR U6691 ( .A(p_input[7586]), .B(n7197), .Z(n7200) );
  XNOR U6692 ( .A(n7197), .B(n6939), .Z(n7199) );
  IV U6693 ( .A(p_input[7554]), .Z(n6939) );
  XNOR U6694 ( .A(n7201), .B(n7202), .Z(n7197) );
  AND U6695 ( .A(n7203), .B(n7204), .Z(n7202) );
  XOR U6696 ( .A(p_input[7585]), .B(n7201), .Z(n7204) );
  XNOR U6697 ( .A(p_input[7553]), .B(n7201), .Z(n7203) );
  AND U6698 ( .A(p_input[7584]), .B(n7205), .Z(n7201) );
  IV U6699 ( .A(p_input[7552]), .Z(n7205) );
  XOR U6700 ( .A(n7206), .B(n7207), .Z(n6295) );
  AND U6701 ( .A(n449), .B(n7208), .Z(n7207) );
  XNOR U6702 ( .A(n7209), .B(n7206), .Z(n7208) );
  XOR U6703 ( .A(n7210), .B(n7211), .Z(n449) );
  AND U6704 ( .A(n7212), .B(n7213), .Z(n7211) );
  XNOR U6705 ( .A(n6310), .B(n7210), .Z(n7213) );
  AND U6706 ( .A(p_input[7551]), .B(p_input[7519]), .Z(n6310) );
  XNOR U6707 ( .A(n7210), .B(n6307), .Z(n7212) );
  IV U6708 ( .A(n7214), .Z(n6307) );
  AND U6709 ( .A(p_input[7455]), .B(p_input[7487]), .Z(n7214) );
  XOR U6710 ( .A(n7215), .B(n7216), .Z(n7210) );
  AND U6711 ( .A(n7217), .B(n7218), .Z(n7216) );
  XOR U6712 ( .A(n7215), .B(n6322), .Z(n7218) );
  XNOR U6713 ( .A(p_input[7518]), .B(n7219), .Z(n6322) );
  AND U6714 ( .A(n219), .B(n7220), .Z(n7219) );
  XOR U6715 ( .A(p_input[7550]), .B(p_input[7518]), .Z(n7220) );
  XNOR U6716 ( .A(n6319), .B(n7215), .Z(n7217) );
  XOR U6717 ( .A(n7221), .B(n7222), .Z(n6319) );
  AND U6718 ( .A(n216), .B(n7223), .Z(n7222) );
  XOR U6719 ( .A(p_input[7486]), .B(p_input[7454]), .Z(n7223) );
  XOR U6720 ( .A(n7224), .B(n7225), .Z(n7215) );
  AND U6721 ( .A(n7226), .B(n7227), .Z(n7225) );
  XOR U6722 ( .A(n7224), .B(n6334), .Z(n7227) );
  XNOR U6723 ( .A(p_input[7517]), .B(n7228), .Z(n6334) );
  AND U6724 ( .A(n219), .B(n7229), .Z(n7228) );
  XOR U6725 ( .A(p_input[7549]), .B(p_input[7517]), .Z(n7229) );
  XNOR U6726 ( .A(n6331), .B(n7224), .Z(n7226) );
  XOR U6727 ( .A(n7230), .B(n7231), .Z(n6331) );
  AND U6728 ( .A(n216), .B(n7232), .Z(n7231) );
  XOR U6729 ( .A(p_input[7485]), .B(p_input[7453]), .Z(n7232) );
  XOR U6730 ( .A(n7233), .B(n7234), .Z(n7224) );
  AND U6731 ( .A(n7235), .B(n7236), .Z(n7234) );
  XOR U6732 ( .A(n7233), .B(n6346), .Z(n7236) );
  XNOR U6733 ( .A(p_input[7516]), .B(n7237), .Z(n6346) );
  AND U6734 ( .A(n219), .B(n7238), .Z(n7237) );
  XOR U6735 ( .A(p_input[7548]), .B(p_input[7516]), .Z(n7238) );
  XNOR U6736 ( .A(n6343), .B(n7233), .Z(n7235) );
  XOR U6737 ( .A(n7239), .B(n7240), .Z(n6343) );
  AND U6738 ( .A(n216), .B(n7241), .Z(n7240) );
  XOR U6739 ( .A(p_input[7484]), .B(p_input[7452]), .Z(n7241) );
  XOR U6740 ( .A(n7242), .B(n7243), .Z(n7233) );
  AND U6741 ( .A(n7244), .B(n7245), .Z(n7243) );
  XOR U6742 ( .A(n7242), .B(n6358), .Z(n7245) );
  XNOR U6743 ( .A(p_input[7515]), .B(n7246), .Z(n6358) );
  AND U6744 ( .A(n219), .B(n7247), .Z(n7246) );
  XOR U6745 ( .A(p_input[7547]), .B(p_input[7515]), .Z(n7247) );
  XNOR U6746 ( .A(n6355), .B(n7242), .Z(n7244) );
  XOR U6747 ( .A(n7248), .B(n7249), .Z(n6355) );
  AND U6748 ( .A(n216), .B(n7250), .Z(n7249) );
  XOR U6749 ( .A(p_input[7483]), .B(p_input[7451]), .Z(n7250) );
  XOR U6750 ( .A(n7251), .B(n7252), .Z(n7242) );
  AND U6751 ( .A(n7253), .B(n7254), .Z(n7252) );
  XOR U6752 ( .A(n7251), .B(n6370), .Z(n7254) );
  XNOR U6753 ( .A(p_input[7514]), .B(n7255), .Z(n6370) );
  AND U6754 ( .A(n219), .B(n7256), .Z(n7255) );
  XOR U6755 ( .A(p_input[7546]), .B(p_input[7514]), .Z(n7256) );
  XNOR U6756 ( .A(n6367), .B(n7251), .Z(n7253) );
  XOR U6757 ( .A(n7257), .B(n7258), .Z(n6367) );
  AND U6758 ( .A(n216), .B(n7259), .Z(n7258) );
  XOR U6759 ( .A(p_input[7482]), .B(p_input[7450]), .Z(n7259) );
  XOR U6760 ( .A(n7260), .B(n7261), .Z(n7251) );
  AND U6761 ( .A(n7262), .B(n7263), .Z(n7261) );
  XOR U6762 ( .A(n7260), .B(n6382), .Z(n7263) );
  XNOR U6763 ( .A(p_input[7513]), .B(n7264), .Z(n6382) );
  AND U6764 ( .A(n219), .B(n7265), .Z(n7264) );
  XOR U6765 ( .A(p_input[7545]), .B(p_input[7513]), .Z(n7265) );
  XNOR U6766 ( .A(n6379), .B(n7260), .Z(n7262) );
  XOR U6767 ( .A(n7266), .B(n7267), .Z(n6379) );
  AND U6768 ( .A(n216), .B(n7268), .Z(n7267) );
  XOR U6769 ( .A(p_input[7481]), .B(p_input[7449]), .Z(n7268) );
  XOR U6770 ( .A(n7269), .B(n7270), .Z(n7260) );
  AND U6771 ( .A(n7271), .B(n7272), .Z(n7270) );
  XOR U6772 ( .A(n7269), .B(n6394), .Z(n7272) );
  XNOR U6773 ( .A(p_input[7512]), .B(n7273), .Z(n6394) );
  AND U6774 ( .A(n219), .B(n7274), .Z(n7273) );
  XOR U6775 ( .A(p_input[7544]), .B(p_input[7512]), .Z(n7274) );
  XNOR U6776 ( .A(n6391), .B(n7269), .Z(n7271) );
  XOR U6777 ( .A(n7275), .B(n7276), .Z(n6391) );
  AND U6778 ( .A(n216), .B(n7277), .Z(n7276) );
  XOR U6779 ( .A(p_input[7480]), .B(p_input[7448]), .Z(n7277) );
  XOR U6780 ( .A(n7278), .B(n7279), .Z(n7269) );
  AND U6781 ( .A(n7280), .B(n7281), .Z(n7279) );
  XOR U6782 ( .A(n7278), .B(n6406), .Z(n7281) );
  XNOR U6783 ( .A(p_input[7511]), .B(n7282), .Z(n6406) );
  AND U6784 ( .A(n219), .B(n7283), .Z(n7282) );
  XOR U6785 ( .A(p_input[7543]), .B(p_input[7511]), .Z(n7283) );
  XNOR U6786 ( .A(n6403), .B(n7278), .Z(n7280) );
  XOR U6787 ( .A(n7284), .B(n7285), .Z(n6403) );
  AND U6788 ( .A(n216), .B(n7286), .Z(n7285) );
  XOR U6789 ( .A(p_input[7479]), .B(p_input[7447]), .Z(n7286) );
  XOR U6790 ( .A(n7287), .B(n7288), .Z(n7278) );
  AND U6791 ( .A(n7289), .B(n7290), .Z(n7288) );
  XOR U6792 ( .A(n7287), .B(n6418), .Z(n7290) );
  XNOR U6793 ( .A(p_input[7510]), .B(n7291), .Z(n6418) );
  AND U6794 ( .A(n219), .B(n7292), .Z(n7291) );
  XOR U6795 ( .A(p_input[7542]), .B(p_input[7510]), .Z(n7292) );
  XNOR U6796 ( .A(n6415), .B(n7287), .Z(n7289) );
  XOR U6797 ( .A(n7293), .B(n7294), .Z(n6415) );
  AND U6798 ( .A(n216), .B(n7295), .Z(n7294) );
  XOR U6799 ( .A(p_input[7478]), .B(p_input[7446]), .Z(n7295) );
  XOR U6800 ( .A(n7296), .B(n7297), .Z(n7287) );
  AND U6801 ( .A(n7298), .B(n7299), .Z(n7297) );
  XOR U6802 ( .A(n7296), .B(n6430), .Z(n7299) );
  XNOR U6803 ( .A(p_input[7509]), .B(n7300), .Z(n6430) );
  AND U6804 ( .A(n219), .B(n7301), .Z(n7300) );
  XOR U6805 ( .A(p_input[7541]), .B(p_input[7509]), .Z(n7301) );
  XNOR U6806 ( .A(n6427), .B(n7296), .Z(n7298) );
  XOR U6807 ( .A(n7302), .B(n7303), .Z(n6427) );
  AND U6808 ( .A(n216), .B(n7304), .Z(n7303) );
  XOR U6809 ( .A(p_input[7477]), .B(p_input[7445]), .Z(n7304) );
  XOR U6810 ( .A(n7305), .B(n7306), .Z(n7296) );
  AND U6811 ( .A(n7307), .B(n7308), .Z(n7306) );
  XOR U6812 ( .A(n7305), .B(n6442), .Z(n7308) );
  XNOR U6813 ( .A(p_input[7508]), .B(n7309), .Z(n6442) );
  AND U6814 ( .A(n219), .B(n7310), .Z(n7309) );
  XOR U6815 ( .A(p_input[7540]), .B(p_input[7508]), .Z(n7310) );
  XNOR U6816 ( .A(n6439), .B(n7305), .Z(n7307) );
  XOR U6817 ( .A(n7311), .B(n7312), .Z(n6439) );
  AND U6818 ( .A(n216), .B(n7313), .Z(n7312) );
  XOR U6819 ( .A(p_input[7476]), .B(p_input[7444]), .Z(n7313) );
  XOR U6820 ( .A(n7314), .B(n7315), .Z(n7305) );
  AND U6821 ( .A(n7316), .B(n7317), .Z(n7315) );
  XOR U6822 ( .A(n7314), .B(n6454), .Z(n7317) );
  XNOR U6823 ( .A(p_input[7507]), .B(n7318), .Z(n6454) );
  AND U6824 ( .A(n219), .B(n7319), .Z(n7318) );
  XOR U6825 ( .A(p_input[7539]), .B(p_input[7507]), .Z(n7319) );
  XNOR U6826 ( .A(n6451), .B(n7314), .Z(n7316) );
  XOR U6827 ( .A(n7320), .B(n7321), .Z(n6451) );
  AND U6828 ( .A(n216), .B(n7322), .Z(n7321) );
  XOR U6829 ( .A(p_input[7475]), .B(p_input[7443]), .Z(n7322) );
  XOR U6830 ( .A(n7323), .B(n7324), .Z(n7314) );
  AND U6831 ( .A(n7325), .B(n7326), .Z(n7324) );
  XOR U6832 ( .A(n7323), .B(n6466), .Z(n7326) );
  XNOR U6833 ( .A(p_input[7506]), .B(n7327), .Z(n6466) );
  AND U6834 ( .A(n219), .B(n7328), .Z(n7327) );
  XOR U6835 ( .A(p_input[7538]), .B(p_input[7506]), .Z(n7328) );
  XNOR U6836 ( .A(n6463), .B(n7323), .Z(n7325) );
  XOR U6837 ( .A(n7329), .B(n7330), .Z(n6463) );
  AND U6838 ( .A(n216), .B(n7331), .Z(n7330) );
  XOR U6839 ( .A(p_input[7474]), .B(p_input[7442]), .Z(n7331) );
  XOR U6840 ( .A(n7332), .B(n7333), .Z(n7323) );
  AND U6841 ( .A(n7334), .B(n7335), .Z(n7333) );
  XOR U6842 ( .A(n7332), .B(n6478), .Z(n7335) );
  XNOR U6843 ( .A(p_input[7505]), .B(n7336), .Z(n6478) );
  AND U6844 ( .A(n219), .B(n7337), .Z(n7336) );
  XOR U6845 ( .A(p_input[7537]), .B(p_input[7505]), .Z(n7337) );
  XNOR U6846 ( .A(n6475), .B(n7332), .Z(n7334) );
  XOR U6847 ( .A(n7338), .B(n7339), .Z(n6475) );
  AND U6848 ( .A(n216), .B(n7340), .Z(n7339) );
  XOR U6849 ( .A(p_input[7473]), .B(p_input[7441]), .Z(n7340) );
  XOR U6850 ( .A(n7341), .B(n7342), .Z(n7332) );
  AND U6851 ( .A(n7343), .B(n7344), .Z(n7342) );
  XOR U6852 ( .A(n7341), .B(n6490), .Z(n7344) );
  XNOR U6853 ( .A(p_input[7504]), .B(n7345), .Z(n6490) );
  AND U6854 ( .A(n219), .B(n7346), .Z(n7345) );
  XOR U6855 ( .A(p_input[7536]), .B(p_input[7504]), .Z(n7346) );
  XNOR U6856 ( .A(n6487), .B(n7341), .Z(n7343) );
  XOR U6857 ( .A(n7347), .B(n7348), .Z(n6487) );
  AND U6858 ( .A(n216), .B(n7349), .Z(n7348) );
  XOR U6859 ( .A(p_input[7472]), .B(p_input[7440]), .Z(n7349) );
  XOR U6860 ( .A(n7350), .B(n7351), .Z(n7341) );
  AND U6861 ( .A(n7352), .B(n7353), .Z(n7351) );
  XOR U6862 ( .A(n7350), .B(n6502), .Z(n7353) );
  XNOR U6863 ( .A(p_input[7503]), .B(n7354), .Z(n6502) );
  AND U6864 ( .A(n219), .B(n7355), .Z(n7354) );
  XOR U6865 ( .A(p_input[7535]), .B(p_input[7503]), .Z(n7355) );
  XNOR U6866 ( .A(n6499), .B(n7350), .Z(n7352) );
  XOR U6867 ( .A(n7356), .B(n7357), .Z(n6499) );
  AND U6868 ( .A(n216), .B(n7358), .Z(n7357) );
  XOR U6869 ( .A(p_input[7471]), .B(p_input[7439]), .Z(n7358) );
  XOR U6870 ( .A(n7359), .B(n7360), .Z(n7350) );
  AND U6871 ( .A(n7361), .B(n7362), .Z(n7360) );
  XOR U6872 ( .A(n7359), .B(n6514), .Z(n7362) );
  XNOR U6873 ( .A(p_input[7502]), .B(n7363), .Z(n6514) );
  AND U6874 ( .A(n219), .B(n7364), .Z(n7363) );
  XOR U6875 ( .A(p_input[7534]), .B(p_input[7502]), .Z(n7364) );
  XNOR U6876 ( .A(n6511), .B(n7359), .Z(n7361) );
  XOR U6877 ( .A(n7365), .B(n7366), .Z(n6511) );
  AND U6878 ( .A(n216), .B(n7367), .Z(n7366) );
  XOR U6879 ( .A(p_input[7470]), .B(p_input[7438]), .Z(n7367) );
  XOR U6880 ( .A(n7368), .B(n7369), .Z(n7359) );
  AND U6881 ( .A(n7370), .B(n7371), .Z(n7369) );
  XOR U6882 ( .A(n7368), .B(n6526), .Z(n7371) );
  XNOR U6883 ( .A(p_input[7501]), .B(n7372), .Z(n6526) );
  AND U6884 ( .A(n219), .B(n7373), .Z(n7372) );
  XOR U6885 ( .A(p_input[7533]), .B(p_input[7501]), .Z(n7373) );
  XNOR U6886 ( .A(n6523), .B(n7368), .Z(n7370) );
  XOR U6887 ( .A(n7374), .B(n7375), .Z(n6523) );
  AND U6888 ( .A(n216), .B(n7376), .Z(n7375) );
  XOR U6889 ( .A(p_input[7469]), .B(p_input[7437]), .Z(n7376) );
  XOR U6890 ( .A(n7377), .B(n7378), .Z(n7368) );
  AND U6891 ( .A(n7379), .B(n7380), .Z(n7378) );
  XOR U6892 ( .A(n7377), .B(n6538), .Z(n7380) );
  XNOR U6893 ( .A(p_input[7500]), .B(n7381), .Z(n6538) );
  AND U6894 ( .A(n219), .B(n7382), .Z(n7381) );
  XOR U6895 ( .A(p_input[7532]), .B(p_input[7500]), .Z(n7382) );
  XNOR U6896 ( .A(n6535), .B(n7377), .Z(n7379) );
  XOR U6897 ( .A(n7383), .B(n7384), .Z(n6535) );
  AND U6898 ( .A(n216), .B(n7385), .Z(n7384) );
  XOR U6899 ( .A(p_input[7468]), .B(p_input[7436]), .Z(n7385) );
  XOR U6900 ( .A(n7386), .B(n7387), .Z(n7377) );
  AND U6901 ( .A(n7388), .B(n7389), .Z(n7387) );
  XOR U6902 ( .A(n7386), .B(n6550), .Z(n7389) );
  XNOR U6903 ( .A(p_input[7499]), .B(n7390), .Z(n6550) );
  AND U6904 ( .A(n219), .B(n7391), .Z(n7390) );
  XOR U6905 ( .A(p_input[7531]), .B(p_input[7499]), .Z(n7391) );
  XNOR U6906 ( .A(n6547), .B(n7386), .Z(n7388) );
  XOR U6907 ( .A(n7392), .B(n7393), .Z(n6547) );
  AND U6908 ( .A(n216), .B(n7394), .Z(n7393) );
  XOR U6909 ( .A(p_input[7467]), .B(p_input[7435]), .Z(n7394) );
  XOR U6910 ( .A(n7395), .B(n7396), .Z(n7386) );
  AND U6911 ( .A(n7397), .B(n7398), .Z(n7396) );
  XOR U6912 ( .A(n7395), .B(n6562), .Z(n7398) );
  XNOR U6913 ( .A(p_input[7498]), .B(n7399), .Z(n6562) );
  AND U6914 ( .A(n219), .B(n7400), .Z(n7399) );
  XOR U6915 ( .A(p_input[7530]), .B(p_input[7498]), .Z(n7400) );
  XNOR U6916 ( .A(n6559), .B(n7395), .Z(n7397) );
  XOR U6917 ( .A(n7401), .B(n7402), .Z(n6559) );
  AND U6918 ( .A(n216), .B(n7403), .Z(n7402) );
  XOR U6919 ( .A(p_input[7466]), .B(p_input[7434]), .Z(n7403) );
  XOR U6920 ( .A(n7404), .B(n7405), .Z(n7395) );
  AND U6921 ( .A(n7406), .B(n7407), .Z(n7405) );
  XOR U6922 ( .A(n7404), .B(n6574), .Z(n7407) );
  XNOR U6923 ( .A(p_input[7497]), .B(n7408), .Z(n6574) );
  AND U6924 ( .A(n219), .B(n7409), .Z(n7408) );
  XOR U6925 ( .A(p_input[7529]), .B(p_input[7497]), .Z(n7409) );
  XNOR U6926 ( .A(n6571), .B(n7404), .Z(n7406) );
  XOR U6927 ( .A(n7410), .B(n7411), .Z(n6571) );
  AND U6928 ( .A(n216), .B(n7412), .Z(n7411) );
  XOR U6929 ( .A(p_input[7465]), .B(p_input[7433]), .Z(n7412) );
  XOR U6930 ( .A(n7413), .B(n7414), .Z(n7404) );
  AND U6931 ( .A(n7415), .B(n7416), .Z(n7414) );
  XOR U6932 ( .A(n7413), .B(n6586), .Z(n7416) );
  XNOR U6933 ( .A(p_input[7496]), .B(n7417), .Z(n6586) );
  AND U6934 ( .A(n219), .B(n7418), .Z(n7417) );
  XOR U6935 ( .A(p_input[7528]), .B(p_input[7496]), .Z(n7418) );
  XNOR U6936 ( .A(n6583), .B(n7413), .Z(n7415) );
  XOR U6937 ( .A(n7419), .B(n7420), .Z(n6583) );
  AND U6938 ( .A(n216), .B(n7421), .Z(n7420) );
  XOR U6939 ( .A(p_input[7464]), .B(p_input[7432]), .Z(n7421) );
  XOR U6940 ( .A(n7422), .B(n7423), .Z(n7413) );
  AND U6941 ( .A(n7424), .B(n7425), .Z(n7423) );
  XOR U6942 ( .A(n7422), .B(n6598), .Z(n7425) );
  XNOR U6943 ( .A(p_input[7495]), .B(n7426), .Z(n6598) );
  AND U6944 ( .A(n219), .B(n7427), .Z(n7426) );
  XOR U6945 ( .A(p_input[7527]), .B(p_input[7495]), .Z(n7427) );
  XNOR U6946 ( .A(n6595), .B(n7422), .Z(n7424) );
  XOR U6947 ( .A(n7428), .B(n7429), .Z(n6595) );
  AND U6948 ( .A(n216), .B(n7430), .Z(n7429) );
  XOR U6949 ( .A(p_input[7463]), .B(p_input[7431]), .Z(n7430) );
  XOR U6950 ( .A(n7431), .B(n7432), .Z(n7422) );
  AND U6951 ( .A(n7433), .B(n7434), .Z(n7432) );
  XOR U6952 ( .A(n7431), .B(n6610), .Z(n7434) );
  XNOR U6953 ( .A(p_input[7494]), .B(n7435), .Z(n6610) );
  AND U6954 ( .A(n219), .B(n7436), .Z(n7435) );
  XOR U6955 ( .A(p_input[7526]), .B(p_input[7494]), .Z(n7436) );
  XNOR U6956 ( .A(n6607), .B(n7431), .Z(n7433) );
  XOR U6957 ( .A(n7437), .B(n7438), .Z(n6607) );
  AND U6958 ( .A(n216), .B(n7439), .Z(n7438) );
  XOR U6959 ( .A(p_input[7462]), .B(p_input[7430]), .Z(n7439) );
  XOR U6960 ( .A(n7440), .B(n7441), .Z(n7431) );
  AND U6961 ( .A(n7442), .B(n7443), .Z(n7441) );
  XOR U6962 ( .A(n7440), .B(n6622), .Z(n7443) );
  XNOR U6963 ( .A(p_input[7493]), .B(n7444), .Z(n6622) );
  AND U6964 ( .A(n219), .B(n7445), .Z(n7444) );
  XOR U6965 ( .A(p_input[7525]), .B(p_input[7493]), .Z(n7445) );
  XNOR U6966 ( .A(n6619), .B(n7440), .Z(n7442) );
  XOR U6967 ( .A(n7446), .B(n7447), .Z(n6619) );
  AND U6968 ( .A(n216), .B(n7448), .Z(n7447) );
  XOR U6969 ( .A(p_input[7461]), .B(p_input[7429]), .Z(n7448) );
  XOR U6970 ( .A(n7449), .B(n7450), .Z(n7440) );
  AND U6971 ( .A(n7451), .B(n7452), .Z(n7450) );
  XOR U6972 ( .A(n7449), .B(n6634), .Z(n7452) );
  XNOR U6973 ( .A(p_input[7492]), .B(n7453), .Z(n6634) );
  AND U6974 ( .A(n219), .B(n7454), .Z(n7453) );
  XOR U6975 ( .A(p_input[7524]), .B(p_input[7492]), .Z(n7454) );
  XNOR U6976 ( .A(n6631), .B(n7449), .Z(n7451) );
  XOR U6977 ( .A(n7455), .B(n7456), .Z(n6631) );
  AND U6978 ( .A(n216), .B(n7457), .Z(n7456) );
  XOR U6979 ( .A(p_input[7460]), .B(p_input[7428]), .Z(n7457) );
  XOR U6980 ( .A(n7458), .B(n7459), .Z(n7449) );
  AND U6981 ( .A(n7460), .B(n7461), .Z(n7459) );
  XOR U6982 ( .A(n7458), .B(n6646), .Z(n7461) );
  XNOR U6983 ( .A(p_input[7491]), .B(n7462), .Z(n6646) );
  AND U6984 ( .A(n219), .B(n7463), .Z(n7462) );
  XOR U6985 ( .A(p_input[7523]), .B(p_input[7491]), .Z(n7463) );
  XNOR U6986 ( .A(n6643), .B(n7458), .Z(n7460) );
  XOR U6987 ( .A(n7464), .B(n7465), .Z(n6643) );
  AND U6988 ( .A(n216), .B(n7466), .Z(n7465) );
  XOR U6989 ( .A(p_input[7459]), .B(p_input[7427]), .Z(n7466) );
  XOR U6990 ( .A(n7467), .B(n7468), .Z(n7458) );
  AND U6991 ( .A(n7469), .B(n7470), .Z(n7468) );
  XOR U6992 ( .A(n7467), .B(n6658), .Z(n7470) );
  XNOR U6993 ( .A(p_input[7490]), .B(n7471), .Z(n6658) );
  AND U6994 ( .A(n219), .B(n7472), .Z(n7471) );
  XOR U6995 ( .A(p_input[7522]), .B(p_input[7490]), .Z(n7472) );
  XNOR U6996 ( .A(n6655), .B(n7467), .Z(n7469) );
  XOR U6997 ( .A(n7473), .B(n7474), .Z(n6655) );
  AND U6998 ( .A(n216), .B(n7475), .Z(n7474) );
  XOR U6999 ( .A(p_input[7458]), .B(p_input[7426]), .Z(n7475) );
  XOR U7000 ( .A(n7476), .B(n7477), .Z(n7467) );
  AND U7001 ( .A(n7478), .B(n7479), .Z(n7477) );
  XNOR U7002 ( .A(n7480), .B(n6671), .Z(n7479) );
  XNOR U7003 ( .A(p_input[7489]), .B(n7481), .Z(n6671) );
  AND U7004 ( .A(n219), .B(n7482), .Z(n7481) );
  XNOR U7005 ( .A(p_input[7521]), .B(n7483), .Z(n7482) );
  IV U7006 ( .A(p_input[7489]), .Z(n7483) );
  XNOR U7007 ( .A(n6668), .B(n7476), .Z(n7478) );
  XNOR U7008 ( .A(p_input[7425]), .B(n7484), .Z(n6668) );
  AND U7009 ( .A(n216), .B(n7485), .Z(n7484) );
  XOR U7010 ( .A(p_input[7457]), .B(p_input[7425]), .Z(n7485) );
  IV U7011 ( .A(n7480), .Z(n7476) );
  AND U7012 ( .A(n7206), .B(n7209), .Z(n7480) );
  XOR U7013 ( .A(p_input[7488]), .B(n7486), .Z(n7209) );
  AND U7014 ( .A(n219), .B(n7487), .Z(n7486) );
  XOR U7015 ( .A(p_input[7520]), .B(p_input[7488]), .Z(n7487) );
  XOR U7016 ( .A(n7488), .B(n7489), .Z(n219) );
  AND U7017 ( .A(n7490), .B(n7491), .Z(n7489) );
  XNOR U7018 ( .A(p_input[7551]), .B(n7488), .Z(n7491) );
  XOR U7019 ( .A(n7488), .B(p_input[7519]), .Z(n7490) );
  XOR U7020 ( .A(n7492), .B(n7493), .Z(n7488) );
  AND U7021 ( .A(n7494), .B(n7495), .Z(n7493) );
  XNOR U7022 ( .A(p_input[7550]), .B(n7492), .Z(n7495) );
  XOR U7023 ( .A(n7492), .B(p_input[7518]), .Z(n7494) );
  XOR U7024 ( .A(n7496), .B(n7497), .Z(n7492) );
  AND U7025 ( .A(n7498), .B(n7499), .Z(n7497) );
  XNOR U7026 ( .A(p_input[7549]), .B(n7496), .Z(n7499) );
  XOR U7027 ( .A(n7496), .B(p_input[7517]), .Z(n7498) );
  XOR U7028 ( .A(n7500), .B(n7501), .Z(n7496) );
  AND U7029 ( .A(n7502), .B(n7503), .Z(n7501) );
  XNOR U7030 ( .A(p_input[7548]), .B(n7500), .Z(n7503) );
  XOR U7031 ( .A(n7500), .B(p_input[7516]), .Z(n7502) );
  XOR U7032 ( .A(n7504), .B(n7505), .Z(n7500) );
  AND U7033 ( .A(n7506), .B(n7507), .Z(n7505) );
  XNOR U7034 ( .A(p_input[7547]), .B(n7504), .Z(n7507) );
  XOR U7035 ( .A(n7504), .B(p_input[7515]), .Z(n7506) );
  XOR U7036 ( .A(n7508), .B(n7509), .Z(n7504) );
  AND U7037 ( .A(n7510), .B(n7511), .Z(n7509) );
  XNOR U7038 ( .A(p_input[7546]), .B(n7508), .Z(n7511) );
  XOR U7039 ( .A(n7508), .B(p_input[7514]), .Z(n7510) );
  XOR U7040 ( .A(n7512), .B(n7513), .Z(n7508) );
  AND U7041 ( .A(n7514), .B(n7515), .Z(n7513) );
  XNOR U7042 ( .A(p_input[7545]), .B(n7512), .Z(n7515) );
  XOR U7043 ( .A(n7512), .B(p_input[7513]), .Z(n7514) );
  XOR U7044 ( .A(n7516), .B(n7517), .Z(n7512) );
  AND U7045 ( .A(n7518), .B(n7519), .Z(n7517) );
  XNOR U7046 ( .A(p_input[7544]), .B(n7516), .Z(n7519) );
  XOR U7047 ( .A(n7516), .B(p_input[7512]), .Z(n7518) );
  XOR U7048 ( .A(n7520), .B(n7521), .Z(n7516) );
  AND U7049 ( .A(n7522), .B(n7523), .Z(n7521) );
  XNOR U7050 ( .A(p_input[7543]), .B(n7520), .Z(n7523) );
  XOR U7051 ( .A(n7520), .B(p_input[7511]), .Z(n7522) );
  XOR U7052 ( .A(n7524), .B(n7525), .Z(n7520) );
  AND U7053 ( .A(n7526), .B(n7527), .Z(n7525) );
  XNOR U7054 ( .A(p_input[7542]), .B(n7524), .Z(n7527) );
  XOR U7055 ( .A(n7524), .B(p_input[7510]), .Z(n7526) );
  XOR U7056 ( .A(n7528), .B(n7529), .Z(n7524) );
  AND U7057 ( .A(n7530), .B(n7531), .Z(n7529) );
  XNOR U7058 ( .A(p_input[7541]), .B(n7528), .Z(n7531) );
  XOR U7059 ( .A(n7528), .B(p_input[7509]), .Z(n7530) );
  XOR U7060 ( .A(n7532), .B(n7533), .Z(n7528) );
  AND U7061 ( .A(n7534), .B(n7535), .Z(n7533) );
  XNOR U7062 ( .A(p_input[7540]), .B(n7532), .Z(n7535) );
  XOR U7063 ( .A(n7532), .B(p_input[7508]), .Z(n7534) );
  XOR U7064 ( .A(n7536), .B(n7537), .Z(n7532) );
  AND U7065 ( .A(n7538), .B(n7539), .Z(n7537) );
  XNOR U7066 ( .A(p_input[7539]), .B(n7536), .Z(n7539) );
  XOR U7067 ( .A(n7536), .B(p_input[7507]), .Z(n7538) );
  XOR U7068 ( .A(n7540), .B(n7541), .Z(n7536) );
  AND U7069 ( .A(n7542), .B(n7543), .Z(n7541) );
  XNOR U7070 ( .A(p_input[7538]), .B(n7540), .Z(n7543) );
  XOR U7071 ( .A(n7540), .B(p_input[7506]), .Z(n7542) );
  XOR U7072 ( .A(n7544), .B(n7545), .Z(n7540) );
  AND U7073 ( .A(n7546), .B(n7547), .Z(n7545) );
  XNOR U7074 ( .A(p_input[7537]), .B(n7544), .Z(n7547) );
  XOR U7075 ( .A(n7544), .B(p_input[7505]), .Z(n7546) );
  XOR U7076 ( .A(n7548), .B(n7549), .Z(n7544) );
  AND U7077 ( .A(n7550), .B(n7551), .Z(n7549) );
  XNOR U7078 ( .A(p_input[7536]), .B(n7548), .Z(n7551) );
  XOR U7079 ( .A(n7548), .B(p_input[7504]), .Z(n7550) );
  XOR U7080 ( .A(n7552), .B(n7553), .Z(n7548) );
  AND U7081 ( .A(n7554), .B(n7555), .Z(n7553) );
  XNOR U7082 ( .A(p_input[7535]), .B(n7552), .Z(n7555) );
  XOR U7083 ( .A(n7552), .B(p_input[7503]), .Z(n7554) );
  XOR U7084 ( .A(n7556), .B(n7557), .Z(n7552) );
  AND U7085 ( .A(n7558), .B(n7559), .Z(n7557) );
  XNOR U7086 ( .A(p_input[7534]), .B(n7556), .Z(n7559) );
  XOR U7087 ( .A(n7556), .B(p_input[7502]), .Z(n7558) );
  XOR U7088 ( .A(n7560), .B(n7561), .Z(n7556) );
  AND U7089 ( .A(n7562), .B(n7563), .Z(n7561) );
  XNOR U7090 ( .A(p_input[7533]), .B(n7560), .Z(n7563) );
  XOR U7091 ( .A(n7560), .B(p_input[7501]), .Z(n7562) );
  XOR U7092 ( .A(n7564), .B(n7565), .Z(n7560) );
  AND U7093 ( .A(n7566), .B(n7567), .Z(n7565) );
  XNOR U7094 ( .A(p_input[7532]), .B(n7564), .Z(n7567) );
  XOR U7095 ( .A(n7564), .B(p_input[7500]), .Z(n7566) );
  XOR U7096 ( .A(n7568), .B(n7569), .Z(n7564) );
  AND U7097 ( .A(n7570), .B(n7571), .Z(n7569) );
  XNOR U7098 ( .A(p_input[7531]), .B(n7568), .Z(n7571) );
  XOR U7099 ( .A(n7568), .B(p_input[7499]), .Z(n7570) );
  XOR U7100 ( .A(n7572), .B(n7573), .Z(n7568) );
  AND U7101 ( .A(n7574), .B(n7575), .Z(n7573) );
  XNOR U7102 ( .A(p_input[7530]), .B(n7572), .Z(n7575) );
  XOR U7103 ( .A(n7572), .B(p_input[7498]), .Z(n7574) );
  XOR U7104 ( .A(n7576), .B(n7577), .Z(n7572) );
  AND U7105 ( .A(n7578), .B(n7579), .Z(n7577) );
  XNOR U7106 ( .A(p_input[7529]), .B(n7576), .Z(n7579) );
  XOR U7107 ( .A(n7576), .B(p_input[7497]), .Z(n7578) );
  XOR U7108 ( .A(n7580), .B(n7581), .Z(n7576) );
  AND U7109 ( .A(n7582), .B(n7583), .Z(n7581) );
  XNOR U7110 ( .A(p_input[7528]), .B(n7580), .Z(n7583) );
  XOR U7111 ( .A(n7580), .B(p_input[7496]), .Z(n7582) );
  XOR U7112 ( .A(n7584), .B(n7585), .Z(n7580) );
  AND U7113 ( .A(n7586), .B(n7587), .Z(n7585) );
  XNOR U7114 ( .A(p_input[7527]), .B(n7584), .Z(n7587) );
  XOR U7115 ( .A(n7584), .B(p_input[7495]), .Z(n7586) );
  XOR U7116 ( .A(n7588), .B(n7589), .Z(n7584) );
  AND U7117 ( .A(n7590), .B(n7591), .Z(n7589) );
  XNOR U7118 ( .A(p_input[7526]), .B(n7588), .Z(n7591) );
  XOR U7119 ( .A(n7588), .B(p_input[7494]), .Z(n7590) );
  XOR U7120 ( .A(n7592), .B(n7593), .Z(n7588) );
  AND U7121 ( .A(n7594), .B(n7595), .Z(n7593) );
  XNOR U7122 ( .A(p_input[7525]), .B(n7592), .Z(n7595) );
  XOR U7123 ( .A(n7592), .B(p_input[7493]), .Z(n7594) );
  XOR U7124 ( .A(n7596), .B(n7597), .Z(n7592) );
  AND U7125 ( .A(n7598), .B(n7599), .Z(n7597) );
  XNOR U7126 ( .A(p_input[7524]), .B(n7596), .Z(n7599) );
  XOR U7127 ( .A(n7596), .B(p_input[7492]), .Z(n7598) );
  XOR U7128 ( .A(n7600), .B(n7601), .Z(n7596) );
  AND U7129 ( .A(n7602), .B(n7603), .Z(n7601) );
  XNOR U7130 ( .A(p_input[7523]), .B(n7600), .Z(n7603) );
  XOR U7131 ( .A(n7600), .B(p_input[7491]), .Z(n7602) );
  XOR U7132 ( .A(n7604), .B(n7605), .Z(n7600) );
  AND U7133 ( .A(n7606), .B(n7607), .Z(n7605) );
  XNOR U7134 ( .A(p_input[7522]), .B(n7604), .Z(n7607) );
  XOR U7135 ( .A(n7604), .B(p_input[7490]), .Z(n7606) );
  XNOR U7136 ( .A(n7608), .B(n7609), .Z(n7604) );
  AND U7137 ( .A(n7610), .B(n7611), .Z(n7609) );
  XOR U7138 ( .A(p_input[7521]), .B(n7608), .Z(n7611) );
  XNOR U7139 ( .A(p_input[7489]), .B(n7608), .Z(n7610) );
  AND U7140 ( .A(p_input[7520]), .B(n7612), .Z(n7608) );
  IV U7141 ( .A(p_input[7488]), .Z(n7612) );
  XNOR U7142 ( .A(p_input[7424]), .B(n7613), .Z(n7206) );
  AND U7143 ( .A(n216), .B(n7614), .Z(n7613) );
  XOR U7144 ( .A(p_input[7456]), .B(p_input[7424]), .Z(n7614) );
  XOR U7145 ( .A(n7615), .B(n7616), .Z(n216) );
  AND U7146 ( .A(n7617), .B(n7618), .Z(n7616) );
  XNOR U7147 ( .A(p_input[7487]), .B(n7615), .Z(n7618) );
  XOR U7148 ( .A(n7615), .B(p_input[7455]), .Z(n7617) );
  XOR U7149 ( .A(n7619), .B(n7620), .Z(n7615) );
  AND U7150 ( .A(n7621), .B(n7622), .Z(n7620) );
  XNOR U7151 ( .A(p_input[7486]), .B(n7619), .Z(n7622) );
  XNOR U7152 ( .A(n7619), .B(n7221), .Z(n7621) );
  IV U7153 ( .A(p_input[7454]), .Z(n7221) );
  XOR U7154 ( .A(n7623), .B(n7624), .Z(n7619) );
  AND U7155 ( .A(n7625), .B(n7626), .Z(n7624) );
  XNOR U7156 ( .A(p_input[7485]), .B(n7623), .Z(n7626) );
  XNOR U7157 ( .A(n7623), .B(n7230), .Z(n7625) );
  IV U7158 ( .A(p_input[7453]), .Z(n7230) );
  XOR U7159 ( .A(n7627), .B(n7628), .Z(n7623) );
  AND U7160 ( .A(n7629), .B(n7630), .Z(n7628) );
  XNOR U7161 ( .A(p_input[7484]), .B(n7627), .Z(n7630) );
  XNOR U7162 ( .A(n7627), .B(n7239), .Z(n7629) );
  IV U7163 ( .A(p_input[7452]), .Z(n7239) );
  XOR U7164 ( .A(n7631), .B(n7632), .Z(n7627) );
  AND U7165 ( .A(n7633), .B(n7634), .Z(n7632) );
  XNOR U7166 ( .A(p_input[7483]), .B(n7631), .Z(n7634) );
  XNOR U7167 ( .A(n7631), .B(n7248), .Z(n7633) );
  IV U7168 ( .A(p_input[7451]), .Z(n7248) );
  XOR U7169 ( .A(n7635), .B(n7636), .Z(n7631) );
  AND U7170 ( .A(n7637), .B(n7638), .Z(n7636) );
  XNOR U7171 ( .A(p_input[7482]), .B(n7635), .Z(n7638) );
  XNOR U7172 ( .A(n7635), .B(n7257), .Z(n7637) );
  IV U7173 ( .A(p_input[7450]), .Z(n7257) );
  XOR U7174 ( .A(n7639), .B(n7640), .Z(n7635) );
  AND U7175 ( .A(n7641), .B(n7642), .Z(n7640) );
  XNOR U7176 ( .A(p_input[7481]), .B(n7639), .Z(n7642) );
  XNOR U7177 ( .A(n7639), .B(n7266), .Z(n7641) );
  IV U7178 ( .A(p_input[7449]), .Z(n7266) );
  XOR U7179 ( .A(n7643), .B(n7644), .Z(n7639) );
  AND U7180 ( .A(n7645), .B(n7646), .Z(n7644) );
  XNOR U7181 ( .A(p_input[7480]), .B(n7643), .Z(n7646) );
  XNOR U7182 ( .A(n7643), .B(n7275), .Z(n7645) );
  IV U7183 ( .A(p_input[7448]), .Z(n7275) );
  XOR U7184 ( .A(n7647), .B(n7648), .Z(n7643) );
  AND U7185 ( .A(n7649), .B(n7650), .Z(n7648) );
  XNOR U7186 ( .A(p_input[7479]), .B(n7647), .Z(n7650) );
  XNOR U7187 ( .A(n7647), .B(n7284), .Z(n7649) );
  IV U7188 ( .A(p_input[7447]), .Z(n7284) );
  XOR U7189 ( .A(n7651), .B(n7652), .Z(n7647) );
  AND U7190 ( .A(n7653), .B(n7654), .Z(n7652) );
  XNOR U7191 ( .A(p_input[7478]), .B(n7651), .Z(n7654) );
  XNOR U7192 ( .A(n7651), .B(n7293), .Z(n7653) );
  IV U7193 ( .A(p_input[7446]), .Z(n7293) );
  XOR U7194 ( .A(n7655), .B(n7656), .Z(n7651) );
  AND U7195 ( .A(n7657), .B(n7658), .Z(n7656) );
  XNOR U7196 ( .A(p_input[7477]), .B(n7655), .Z(n7658) );
  XNOR U7197 ( .A(n7655), .B(n7302), .Z(n7657) );
  IV U7198 ( .A(p_input[7445]), .Z(n7302) );
  XOR U7199 ( .A(n7659), .B(n7660), .Z(n7655) );
  AND U7200 ( .A(n7661), .B(n7662), .Z(n7660) );
  XNOR U7201 ( .A(p_input[7476]), .B(n7659), .Z(n7662) );
  XNOR U7202 ( .A(n7659), .B(n7311), .Z(n7661) );
  IV U7203 ( .A(p_input[7444]), .Z(n7311) );
  XOR U7204 ( .A(n7663), .B(n7664), .Z(n7659) );
  AND U7205 ( .A(n7665), .B(n7666), .Z(n7664) );
  XNOR U7206 ( .A(p_input[7475]), .B(n7663), .Z(n7666) );
  XNOR U7207 ( .A(n7663), .B(n7320), .Z(n7665) );
  IV U7208 ( .A(p_input[7443]), .Z(n7320) );
  XOR U7209 ( .A(n7667), .B(n7668), .Z(n7663) );
  AND U7210 ( .A(n7669), .B(n7670), .Z(n7668) );
  XNOR U7211 ( .A(p_input[7474]), .B(n7667), .Z(n7670) );
  XNOR U7212 ( .A(n7667), .B(n7329), .Z(n7669) );
  IV U7213 ( .A(p_input[7442]), .Z(n7329) );
  XOR U7214 ( .A(n7671), .B(n7672), .Z(n7667) );
  AND U7215 ( .A(n7673), .B(n7674), .Z(n7672) );
  XNOR U7216 ( .A(p_input[7473]), .B(n7671), .Z(n7674) );
  XNOR U7217 ( .A(n7671), .B(n7338), .Z(n7673) );
  IV U7218 ( .A(p_input[7441]), .Z(n7338) );
  XOR U7219 ( .A(n7675), .B(n7676), .Z(n7671) );
  AND U7220 ( .A(n7677), .B(n7678), .Z(n7676) );
  XNOR U7221 ( .A(p_input[7472]), .B(n7675), .Z(n7678) );
  XNOR U7222 ( .A(n7675), .B(n7347), .Z(n7677) );
  IV U7223 ( .A(p_input[7440]), .Z(n7347) );
  XOR U7224 ( .A(n7679), .B(n7680), .Z(n7675) );
  AND U7225 ( .A(n7681), .B(n7682), .Z(n7680) );
  XNOR U7226 ( .A(p_input[7471]), .B(n7679), .Z(n7682) );
  XNOR U7227 ( .A(n7679), .B(n7356), .Z(n7681) );
  IV U7228 ( .A(p_input[7439]), .Z(n7356) );
  XOR U7229 ( .A(n7683), .B(n7684), .Z(n7679) );
  AND U7230 ( .A(n7685), .B(n7686), .Z(n7684) );
  XNOR U7231 ( .A(p_input[7470]), .B(n7683), .Z(n7686) );
  XNOR U7232 ( .A(n7683), .B(n7365), .Z(n7685) );
  IV U7233 ( .A(p_input[7438]), .Z(n7365) );
  XOR U7234 ( .A(n7687), .B(n7688), .Z(n7683) );
  AND U7235 ( .A(n7689), .B(n7690), .Z(n7688) );
  XNOR U7236 ( .A(p_input[7469]), .B(n7687), .Z(n7690) );
  XNOR U7237 ( .A(n7687), .B(n7374), .Z(n7689) );
  IV U7238 ( .A(p_input[7437]), .Z(n7374) );
  XOR U7239 ( .A(n7691), .B(n7692), .Z(n7687) );
  AND U7240 ( .A(n7693), .B(n7694), .Z(n7692) );
  XNOR U7241 ( .A(p_input[7468]), .B(n7691), .Z(n7694) );
  XNOR U7242 ( .A(n7691), .B(n7383), .Z(n7693) );
  IV U7243 ( .A(p_input[7436]), .Z(n7383) );
  XOR U7244 ( .A(n7695), .B(n7696), .Z(n7691) );
  AND U7245 ( .A(n7697), .B(n7698), .Z(n7696) );
  XNOR U7246 ( .A(p_input[7467]), .B(n7695), .Z(n7698) );
  XNOR U7247 ( .A(n7695), .B(n7392), .Z(n7697) );
  IV U7248 ( .A(p_input[7435]), .Z(n7392) );
  XOR U7249 ( .A(n7699), .B(n7700), .Z(n7695) );
  AND U7250 ( .A(n7701), .B(n7702), .Z(n7700) );
  XNOR U7251 ( .A(p_input[7466]), .B(n7699), .Z(n7702) );
  XNOR U7252 ( .A(n7699), .B(n7401), .Z(n7701) );
  IV U7253 ( .A(p_input[7434]), .Z(n7401) );
  XOR U7254 ( .A(n7703), .B(n7704), .Z(n7699) );
  AND U7255 ( .A(n7705), .B(n7706), .Z(n7704) );
  XNOR U7256 ( .A(p_input[7465]), .B(n7703), .Z(n7706) );
  XNOR U7257 ( .A(n7703), .B(n7410), .Z(n7705) );
  IV U7258 ( .A(p_input[7433]), .Z(n7410) );
  XOR U7259 ( .A(n7707), .B(n7708), .Z(n7703) );
  AND U7260 ( .A(n7709), .B(n7710), .Z(n7708) );
  XNOR U7261 ( .A(p_input[7464]), .B(n7707), .Z(n7710) );
  XNOR U7262 ( .A(n7707), .B(n7419), .Z(n7709) );
  IV U7263 ( .A(p_input[7432]), .Z(n7419) );
  XOR U7264 ( .A(n7711), .B(n7712), .Z(n7707) );
  AND U7265 ( .A(n7713), .B(n7714), .Z(n7712) );
  XNOR U7266 ( .A(p_input[7463]), .B(n7711), .Z(n7714) );
  XNOR U7267 ( .A(n7711), .B(n7428), .Z(n7713) );
  IV U7268 ( .A(p_input[7431]), .Z(n7428) );
  XOR U7269 ( .A(n7715), .B(n7716), .Z(n7711) );
  AND U7270 ( .A(n7717), .B(n7718), .Z(n7716) );
  XNOR U7271 ( .A(p_input[7462]), .B(n7715), .Z(n7718) );
  XNOR U7272 ( .A(n7715), .B(n7437), .Z(n7717) );
  IV U7273 ( .A(p_input[7430]), .Z(n7437) );
  XOR U7274 ( .A(n7719), .B(n7720), .Z(n7715) );
  AND U7275 ( .A(n7721), .B(n7722), .Z(n7720) );
  XNOR U7276 ( .A(p_input[7461]), .B(n7719), .Z(n7722) );
  XNOR U7277 ( .A(n7719), .B(n7446), .Z(n7721) );
  IV U7278 ( .A(p_input[7429]), .Z(n7446) );
  XOR U7279 ( .A(n7723), .B(n7724), .Z(n7719) );
  AND U7280 ( .A(n7725), .B(n7726), .Z(n7724) );
  XNOR U7281 ( .A(p_input[7460]), .B(n7723), .Z(n7726) );
  XNOR U7282 ( .A(n7723), .B(n7455), .Z(n7725) );
  IV U7283 ( .A(p_input[7428]), .Z(n7455) );
  XOR U7284 ( .A(n7727), .B(n7728), .Z(n7723) );
  AND U7285 ( .A(n7729), .B(n7730), .Z(n7728) );
  XNOR U7286 ( .A(p_input[7459]), .B(n7727), .Z(n7730) );
  XNOR U7287 ( .A(n7727), .B(n7464), .Z(n7729) );
  IV U7288 ( .A(p_input[7427]), .Z(n7464) );
  XOR U7289 ( .A(n7731), .B(n7732), .Z(n7727) );
  AND U7290 ( .A(n7733), .B(n7734), .Z(n7732) );
  XNOR U7291 ( .A(p_input[7458]), .B(n7731), .Z(n7734) );
  XNOR U7292 ( .A(n7731), .B(n7473), .Z(n7733) );
  IV U7293 ( .A(p_input[7426]), .Z(n7473) );
  XNOR U7294 ( .A(n7735), .B(n7736), .Z(n7731) );
  AND U7295 ( .A(n7737), .B(n7738), .Z(n7736) );
  XOR U7296 ( .A(p_input[7457]), .B(n7735), .Z(n7738) );
  XNOR U7297 ( .A(p_input[7425]), .B(n7735), .Z(n7737) );
  AND U7298 ( .A(p_input[7456]), .B(n7739), .Z(n7735) );
  IV U7299 ( .A(p_input[7424]), .Z(n7739) );
  XOR U7300 ( .A(n7740), .B(n7741), .Z(n5918) );
  AND U7301 ( .A(n816), .B(n7742), .Z(n7741) );
  XNOR U7302 ( .A(n7743), .B(n7740), .Z(n7742) );
  XOR U7303 ( .A(n7744), .B(n7745), .Z(n816) );
  AND U7304 ( .A(n7746), .B(n7747), .Z(n7745) );
  XOR U7305 ( .A(n7744), .B(n5933), .Z(n7747) );
  XNOR U7306 ( .A(n7748), .B(n7749), .Z(n5933) );
  AND U7307 ( .A(n7750), .B(n455), .Z(n7749) );
  AND U7308 ( .A(n7748), .B(n7751), .Z(n7750) );
  XNOR U7309 ( .A(n5930), .B(n7744), .Z(n7746) );
  XOR U7310 ( .A(n7752), .B(n7753), .Z(n5930) );
  AND U7311 ( .A(n7754), .B(n452), .Z(n7753) );
  NOR U7312 ( .A(n7752), .B(n7755), .Z(n7754) );
  XOR U7313 ( .A(n7756), .B(n7757), .Z(n7744) );
  AND U7314 ( .A(n7758), .B(n7759), .Z(n7757) );
  XOR U7315 ( .A(n7756), .B(n5945), .Z(n7759) );
  XOR U7316 ( .A(n7760), .B(n7761), .Z(n5945) );
  AND U7317 ( .A(n455), .B(n7762), .Z(n7761) );
  XOR U7318 ( .A(n7763), .B(n7760), .Z(n7762) );
  XNOR U7319 ( .A(n5942), .B(n7756), .Z(n7758) );
  XOR U7320 ( .A(n7764), .B(n7765), .Z(n5942) );
  AND U7321 ( .A(n452), .B(n7766), .Z(n7765) );
  XOR U7322 ( .A(n7767), .B(n7764), .Z(n7766) );
  XOR U7323 ( .A(n7768), .B(n7769), .Z(n7756) );
  AND U7324 ( .A(n7770), .B(n7771), .Z(n7769) );
  XOR U7325 ( .A(n7768), .B(n5957), .Z(n7771) );
  XOR U7326 ( .A(n7772), .B(n7773), .Z(n5957) );
  AND U7327 ( .A(n455), .B(n7774), .Z(n7773) );
  XOR U7328 ( .A(n7775), .B(n7772), .Z(n7774) );
  XNOR U7329 ( .A(n5954), .B(n7768), .Z(n7770) );
  XOR U7330 ( .A(n7776), .B(n7777), .Z(n5954) );
  AND U7331 ( .A(n452), .B(n7778), .Z(n7777) );
  XOR U7332 ( .A(n7779), .B(n7776), .Z(n7778) );
  XOR U7333 ( .A(n7780), .B(n7781), .Z(n7768) );
  AND U7334 ( .A(n7782), .B(n7783), .Z(n7781) );
  XOR U7335 ( .A(n7780), .B(n5969), .Z(n7783) );
  XOR U7336 ( .A(n7784), .B(n7785), .Z(n5969) );
  AND U7337 ( .A(n455), .B(n7786), .Z(n7785) );
  XOR U7338 ( .A(n7787), .B(n7784), .Z(n7786) );
  XNOR U7339 ( .A(n5966), .B(n7780), .Z(n7782) );
  XOR U7340 ( .A(n7788), .B(n7789), .Z(n5966) );
  AND U7341 ( .A(n452), .B(n7790), .Z(n7789) );
  XOR U7342 ( .A(n7791), .B(n7788), .Z(n7790) );
  XOR U7343 ( .A(n7792), .B(n7793), .Z(n7780) );
  AND U7344 ( .A(n7794), .B(n7795), .Z(n7793) );
  XOR U7345 ( .A(n7792), .B(n5981), .Z(n7795) );
  XOR U7346 ( .A(n7796), .B(n7797), .Z(n5981) );
  AND U7347 ( .A(n455), .B(n7798), .Z(n7797) );
  XOR U7348 ( .A(n7799), .B(n7796), .Z(n7798) );
  XNOR U7349 ( .A(n5978), .B(n7792), .Z(n7794) );
  XOR U7350 ( .A(n7800), .B(n7801), .Z(n5978) );
  AND U7351 ( .A(n452), .B(n7802), .Z(n7801) );
  XOR U7352 ( .A(n7803), .B(n7800), .Z(n7802) );
  XOR U7353 ( .A(n7804), .B(n7805), .Z(n7792) );
  AND U7354 ( .A(n7806), .B(n7807), .Z(n7805) );
  XOR U7355 ( .A(n7804), .B(n5993), .Z(n7807) );
  XOR U7356 ( .A(n7808), .B(n7809), .Z(n5993) );
  AND U7357 ( .A(n455), .B(n7810), .Z(n7809) );
  XOR U7358 ( .A(n7811), .B(n7808), .Z(n7810) );
  XNOR U7359 ( .A(n5990), .B(n7804), .Z(n7806) );
  XOR U7360 ( .A(n7812), .B(n7813), .Z(n5990) );
  AND U7361 ( .A(n452), .B(n7814), .Z(n7813) );
  XOR U7362 ( .A(n7815), .B(n7812), .Z(n7814) );
  XOR U7363 ( .A(n7816), .B(n7817), .Z(n7804) );
  AND U7364 ( .A(n7818), .B(n7819), .Z(n7817) );
  XOR U7365 ( .A(n7816), .B(n6005), .Z(n7819) );
  XOR U7366 ( .A(n7820), .B(n7821), .Z(n6005) );
  AND U7367 ( .A(n455), .B(n7822), .Z(n7821) );
  XOR U7368 ( .A(n7823), .B(n7820), .Z(n7822) );
  XNOR U7369 ( .A(n6002), .B(n7816), .Z(n7818) );
  XOR U7370 ( .A(n7824), .B(n7825), .Z(n6002) );
  AND U7371 ( .A(n452), .B(n7826), .Z(n7825) );
  XOR U7372 ( .A(n7827), .B(n7824), .Z(n7826) );
  XOR U7373 ( .A(n7828), .B(n7829), .Z(n7816) );
  AND U7374 ( .A(n7830), .B(n7831), .Z(n7829) );
  XOR U7375 ( .A(n7828), .B(n6017), .Z(n7831) );
  XOR U7376 ( .A(n7832), .B(n7833), .Z(n6017) );
  AND U7377 ( .A(n455), .B(n7834), .Z(n7833) );
  XOR U7378 ( .A(n7835), .B(n7832), .Z(n7834) );
  XNOR U7379 ( .A(n6014), .B(n7828), .Z(n7830) );
  XOR U7380 ( .A(n7836), .B(n7837), .Z(n6014) );
  AND U7381 ( .A(n452), .B(n7838), .Z(n7837) );
  XOR U7382 ( .A(n7839), .B(n7836), .Z(n7838) );
  XOR U7383 ( .A(n7840), .B(n7841), .Z(n7828) );
  AND U7384 ( .A(n7842), .B(n7843), .Z(n7841) );
  XOR U7385 ( .A(n7840), .B(n6029), .Z(n7843) );
  XOR U7386 ( .A(n7844), .B(n7845), .Z(n6029) );
  AND U7387 ( .A(n455), .B(n7846), .Z(n7845) );
  XOR U7388 ( .A(n7847), .B(n7844), .Z(n7846) );
  XNOR U7389 ( .A(n6026), .B(n7840), .Z(n7842) );
  XOR U7390 ( .A(n7848), .B(n7849), .Z(n6026) );
  AND U7391 ( .A(n452), .B(n7850), .Z(n7849) );
  XOR U7392 ( .A(n7851), .B(n7848), .Z(n7850) );
  XOR U7393 ( .A(n7852), .B(n7853), .Z(n7840) );
  AND U7394 ( .A(n7854), .B(n7855), .Z(n7853) );
  XOR U7395 ( .A(n7852), .B(n6041), .Z(n7855) );
  XOR U7396 ( .A(n7856), .B(n7857), .Z(n6041) );
  AND U7397 ( .A(n455), .B(n7858), .Z(n7857) );
  XOR U7398 ( .A(n7859), .B(n7856), .Z(n7858) );
  XNOR U7399 ( .A(n6038), .B(n7852), .Z(n7854) );
  XOR U7400 ( .A(n7860), .B(n7861), .Z(n6038) );
  AND U7401 ( .A(n452), .B(n7862), .Z(n7861) );
  XOR U7402 ( .A(n7863), .B(n7860), .Z(n7862) );
  XOR U7403 ( .A(n7864), .B(n7865), .Z(n7852) );
  AND U7404 ( .A(n7866), .B(n7867), .Z(n7865) );
  XOR U7405 ( .A(n7864), .B(n6053), .Z(n7867) );
  XOR U7406 ( .A(n7868), .B(n7869), .Z(n6053) );
  AND U7407 ( .A(n455), .B(n7870), .Z(n7869) );
  XOR U7408 ( .A(n7871), .B(n7868), .Z(n7870) );
  XNOR U7409 ( .A(n6050), .B(n7864), .Z(n7866) );
  XOR U7410 ( .A(n7872), .B(n7873), .Z(n6050) );
  AND U7411 ( .A(n452), .B(n7874), .Z(n7873) );
  XOR U7412 ( .A(n7875), .B(n7872), .Z(n7874) );
  XOR U7413 ( .A(n7876), .B(n7877), .Z(n7864) );
  AND U7414 ( .A(n7878), .B(n7879), .Z(n7877) );
  XOR U7415 ( .A(n7876), .B(n6065), .Z(n7879) );
  XOR U7416 ( .A(n7880), .B(n7881), .Z(n6065) );
  AND U7417 ( .A(n455), .B(n7882), .Z(n7881) );
  XOR U7418 ( .A(n7883), .B(n7880), .Z(n7882) );
  XNOR U7419 ( .A(n6062), .B(n7876), .Z(n7878) );
  XOR U7420 ( .A(n7884), .B(n7885), .Z(n6062) );
  AND U7421 ( .A(n452), .B(n7886), .Z(n7885) );
  XOR U7422 ( .A(n7887), .B(n7884), .Z(n7886) );
  XOR U7423 ( .A(n7888), .B(n7889), .Z(n7876) );
  AND U7424 ( .A(n7890), .B(n7891), .Z(n7889) );
  XOR U7425 ( .A(n7888), .B(n6077), .Z(n7891) );
  XOR U7426 ( .A(n7892), .B(n7893), .Z(n6077) );
  AND U7427 ( .A(n455), .B(n7894), .Z(n7893) );
  XOR U7428 ( .A(n7895), .B(n7892), .Z(n7894) );
  XNOR U7429 ( .A(n6074), .B(n7888), .Z(n7890) );
  XOR U7430 ( .A(n7896), .B(n7897), .Z(n6074) );
  AND U7431 ( .A(n452), .B(n7898), .Z(n7897) );
  XOR U7432 ( .A(n7899), .B(n7896), .Z(n7898) );
  XOR U7433 ( .A(n7900), .B(n7901), .Z(n7888) );
  AND U7434 ( .A(n7902), .B(n7903), .Z(n7901) );
  XOR U7435 ( .A(n7900), .B(n6089), .Z(n7903) );
  XOR U7436 ( .A(n7904), .B(n7905), .Z(n6089) );
  AND U7437 ( .A(n455), .B(n7906), .Z(n7905) );
  XOR U7438 ( .A(n7907), .B(n7904), .Z(n7906) );
  XNOR U7439 ( .A(n6086), .B(n7900), .Z(n7902) );
  XOR U7440 ( .A(n7908), .B(n7909), .Z(n6086) );
  AND U7441 ( .A(n452), .B(n7910), .Z(n7909) );
  XOR U7442 ( .A(n7911), .B(n7908), .Z(n7910) );
  XOR U7443 ( .A(n7912), .B(n7913), .Z(n7900) );
  AND U7444 ( .A(n7914), .B(n7915), .Z(n7913) );
  XOR U7445 ( .A(n7912), .B(n6101), .Z(n7915) );
  XOR U7446 ( .A(n7916), .B(n7917), .Z(n6101) );
  AND U7447 ( .A(n455), .B(n7918), .Z(n7917) );
  XOR U7448 ( .A(n7919), .B(n7916), .Z(n7918) );
  XNOR U7449 ( .A(n6098), .B(n7912), .Z(n7914) );
  XOR U7450 ( .A(n7920), .B(n7921), .Z(n6098) );
  AND U7451 ( .A(n452), .B(n7922), .Z(n7921) );
  XOR U7452 ( .A(n7923), .B(n7920), .Z(n7922) );
  XOR U7453 ( .A(n7924), .B(n7925), .Z(n7912) );
  AND U7454 ( .A(n7926), .B(n7927), .Z(n7925) );
  XOR U7455 ( .A(n7924), .B(n6113), .Z(n7927) );
  XOR U7456 ( .A(n7928), .B(n7929), .Z(n6113) );
  AND U7457 ( .A(n455), .B(n7930), .Z(n7929) );
  XOR U7458 ( .A(n7931), .B(n7928), .Z(n7930) );
  XNOR U7459 ( .A(n6110), .B(n7924), .Z(n7926) );
  XOR U7460 ( .A(n7932), .B(n7933), .Z(n6110) );
  AND U7461 ( .A(n452), .B(n7934), .Z(n7933) );
  XOR U7462 ( .A(n7935), .B(n7932), .Z(n7934) );
  XOR U7463 ( .A(n7936), .B(n7937), .Z(n7924) );
  AND U7464 ( .A(n7938), .B(n7939), .Z(n7937) );
  XOR U7465 ( .A(n7936), .B(n6125), .Z(n7939) );
  XOR U7466 ( .A(n7940), .B(n7941), .Z(n6125) );
  AND U7467 ( .A(n455), .B(n7942), .Z(n7941) );
  XOR U7468 ( .A(n7943), .B(n7940), .Z(n7942) );
  XNOR U7469 ( .A(n6122), .B(n7936), .Z(n7938) );
  XOR U7470 ( .A(n7944), .B(n7945), .Z(n6122) );
  AND U7471 ( .A(n452), .B(n7946), .Z(n7945) );
  XOR U7472 ( .A(n7947), .B(n7944), .Z(n7946) );
  XOR U7473 ( .A(n7948), .B(n7949), .Z(n7936) );
  AND U7474 ( .A(n7950), .B(n7951), .Z(n7949) );
  XOR U7475 ( .A(n7948), .B(n6137), .Z(n7951) );
  XOR U7476 ( .A(n7952), .B(n7953), .Z(n6137) );
  AND U7477 ( .A(n455), .B(n7954), .Z(n7953) );
  XOR U7478 ( .A(n7955), .B(n7952), .Z(n7954) );
  XNOR U7479 ( .A(n6134), .B(n7948), .Z(n7950) );
  XOR U7480 ( .A(n7956), .B(n7957), .Z(n6134) );
  AND U7481 ( .A(n452), .B(n7958), .Z(n7957) );
  XOR U7482 ( .A(n7959), .B(n7956), .Z(n7958) );
  XOR U7483 ( .A(n7960), .B(n7961), .Z(n7948) );
  AND U7484 ( .A(n7962), .B(n7963), .Z(n7961) );
  XOR U7485 ( .A(n7960), .B(n6149), .Z(n7963) );
  XOR U7486 ( .A(n7964), .B(n7965), .Z(n6149) );
  AND U7487 ( .A(n455), .B(n7966), .Z(n7965) );
  XOR U7488 ( .A(n7967), .B(n7964), .Z(n7966) );
  XNOR U7489 ( .A(n6146), .B(n7960), .Z(n7962) );
  XOR U7490 ( .A(n7968), .B(n7969), .Z(n6146) );
  AND U7491 ( .A(n452), .B(n7970), .Z(n7969) );
  XOR U7492 ( .A(n7971), .B(n7968), .Z(n7970) );
  XOR U7493 ( .A(n7972), .B(n7973), .Z(n7960) );
  AND U7494 ( .A(n7974), .B(n7975), .Z(n7973) );
  XOR U7495 ( .A(n7972), .B(n6161), .Z(n7975) );
  XOR U7496 ( .A(n7976), .B(n7977), .Z(n6161) );
  AND U7497 ( .A(n455), .B(n7978), .Z(n7977) );
  XOR U7498 ( .A(n7979), .B(n7976), .Z(n7978) );
  XNOR U7499 ( .A(n6158), .B(n7972), .Z(n7974) );
  XOR U7500 ( .A(n7980), .B(n7981), .Z(n6158) );
  AND U7501 ( .A(n452), .B(n7982), .Z(n7981) );
  XOR U7502 ( .A(n7983), .B(n7980), .Z(n7982) );
  XOR U7503 ( .A(n7984), .B(n7985), .Z(n7972) );
  AND U7504 ( .A(n7986), .B(n7987), .Z(n7985) );
  XOR U7505 ( .A(n7984), .B(n6173), .Z(n7987) );
  XOR U7506 ( .A(n7988), .B(n7989), .Z(n6173) );
  AND U7507 ( .A(n455), .B(n7990), .Z(n7989) );
  XOR U7508 ( .A(n7991), .B(n7988), .Z(n7990) );
  XNOR U7509 ( .A(n6170), .B(n7984), .Z(n7986) );
  XOR U7510 ( .A(n7992), .B(n7993), .Z(n6170) );
  AND U7511 ( .A(n452), .B(n7994), .Z(n7993) );
  XOR U7512 ( .A(n7995), .B(n7992), .Z(n7994) );
  XOR U7513 ( .A(n7996), .B(n7997), .Z(n7984) );
  AND U7514 ( .A(n7998), .B(n7999), .Z(n7997) );
  XOR U7515 ( .A(n7996), .B(n6185), .Z(n7999) );
  XOR U7516 ( .A(n8000), .B(n8001), .Z(n6185) );
  AND U7517 ( .A(n455), .B(n8002), .Z(n8001) );
  XOR U7518 ( .A(n8003), .B(n8000), .Z(n8002) );
  XNOR U7519 ( .A(n6182), .B(n7996), .Z(n7998) );
  XOR U7520 ( .A(n8004), .B(n8005), .Z(n6182) );
  AND U7521 ( .A(n452), .B(n8006), .Z(n8005) );
  XOR U7522 ( .A(n8007), .B(n8004), .Z(n8006) );
  XOR U7523 ( .A(n8008), .B(n8009), .Z(n7996) );
  AND U7524 ( .A(n8010), .B(n8011), .Z(n8009) );
  XOR U7525 ( .A(n8008), .B(n6197), .Z(n8011) );
  XOR U7526 ( .A(n8012), .B(n8013), .Z(n6197) );
  AND U7527 ( .A(n455), .B(n8014), .Z(n8013) );
  XOR U7528 ( .A(n8015), .B(n8012), .Z(n8014) );
  XNOR U7529 ( .A(n6194), .B(n8008), .Z(n8010) );
  XOR U7530 ( .A(n8016), .B(n8017), .Z(n6194) );
  AND U7531 ( .A(n452), .B(n8018), .Z(n8017) );
  XOR U7532 ( .A(n8019), .B(n8016), .Z(n8018) );
  XOR U7533 ( .A(n8020), .B(n8021), .Z(n8008) );
  AND U7534 ( .A(n8022), .B(n8023), .Z(n8021) );
  XOR U7535 ( .A(n8020), .B(n6209), .Z(n8023) );
  XOR U7536 ( .A(n8024), .B(n8025), .Z(n6209) );
  AND U7537 ( .A(n455), .B(n8026), .Z(n8025) );
  XOR U7538 ( .A(n8027), .B(n8024), .Z(n8026) );
  XNOR U7539 ( .A(n6206), .B(n8020), .Z(n8022) );
  XOR U7540 ( .A(n8028), .B(n8029), .Z(n6206) );
  AND U7541 ( .A(n452), .B(n8030), .Z(n8029) );
  XOR U7542 ( .A(n8031), .B(n8028), .Z(n8030) );
  XOR U7543 ( .A(n8032), .B(n8033), .Z(n8020) );
  AND U7544 ( .A(n8034), .B(n8035), .Z(n8033) );
  XOR U7545 ( .A(n8032), .B(n6221), .Z(n8035) );
  XOR U7546 ( .A(n8036), .B(n8037), .Z(n6221) );
  AND U7547 ( .A(n455), .B(n8038), .Z(n8037) );
  XOR U7548 ( .A(n8039), .B(n8036), .Z(n8038) );
  XNOR U7549 ( .A(n6218), .B(n8032), .Z(n8034) );
  XOR U7550 ( .A(n8040), .B(n8041), .Z(n6218) );
  AND U7551 ( .A(n452), .B(n8042), .Z(n8041) );
  XOR U7552 ( .A(n8043), .B(n8040), .Z(n8042) );
  XOR U7553 ( .A(n8044), .B(n8045), .Z(n8032) );
  AND U7554 ( .A(n8046), .B(n8047), .Z(n8045) );
  XOR U7555 ( .A(n8044), .B(n6233), .Z(n8047) );
  XOR U7556 ( .A(n8048), .B(n8049), .Z(n6233) );
  AND U7557 ( .A(n455), .B(n8050), .Z(n8049) );
  XOR U7558 ( .A(n8051), .B(n8048), .Z(n8050) );
  XNOR U7559 ( .A(n6230), .B(n8044), .Z(n8046) );
  XOR U7560 ( .A(n8052), .B(n8053), .Z(n6230) );
  AND U7561 ( .A(n452), .B(n8054), .Z(n8053) );
  XOR U7562 ( .A(n8055), .B(n8052), .Z(n8054) );
  XOR U7563 ( .A(n8056), .B(n8057), .Z(n8044) );
  AND U7564 ( .A(n8058), .B(n8059), .Z(n8057) );
  XOR U7565 ( .A(n8056), .B(n6245), .Z(n8059) );
  XOR U7566 ( .A(n8060), .B(n8061), .Z(n6245) );
  AND U7567 ( .A(n455), .B(n8062), .Z(n8061) );
  XOR U7568 ( .A(n8063), .B(n8060), .Z(n8062) );
  XNOR U7569 ( .A(n6242), .B(n8056), .Z(n8058) );
  XOR U7570 ( .A(n8064), .B(n8065), .Z(n6242) );
  AND U7571 ( .A(n452), .B(n8066), .Z(n8065) );
  XOR U7572 ( .A(n8067), .B(n8064), .Z(n8066) );
  XOR U7573 ( .A(n8068), .B(n8069), .Z(n8056) );
  AND U7574 ( .A(n8070), .B(n8071), .Z(n8069) );
  XOR U7575 ( .A(n8068), .B(n6257), .Z(n8071) );
  XOR U7576 ( .A(n8072), .B(n8073), .Z(n6257) );
  AND U7577 ( .A(n455), .B(n8074), .Z(n8073) );
  XOR U7578 ( .A(n8075), .B(n8072), .Z(n8074) );
  XNOR U7579 ( .A(n6254), .B(n8068), .Z(n8070) );
  XOR U7580 ( .A(n8076), .B(n8077), .Z(n6254) );
  AND U7581 ( .A(n452), .B(n8078), .Z(n8077) );
  XOR U7582 ( .A(n8079), .B(n8076), .Z(n8078) );
  XOR U7583 ( .A(n8080), .B(n8081), .Z(n8068) );
  AND U7584 ( .A(n8082), .B(n8083), .Z(n8081) );
  XOR U7585 ( .A(n8080), .B(n6269), .Z(n8083) );
  XOR U7586 ( .A(n8084), .B(n8085), .Z(n6269) );
  AND U7587 ( .A(n455), .B(n8086), .Z(n8085) );
  XOR U7588 ( .A(n8087), .B(n8084), .Z(n8086) );
  XNOR U7589 ( .A(n6266), .B(n8080), .Z(n8082) );
  XOR U7590 ( .A(n8088), .B(n8089), .Z(n6266) );
  AND U7591 ( .A(n452), .B(n8090), .Z(n8089) );
  XOR U7592 ( .A(n8091), .B(n8088), .Z(n8090) );
  XOR U7593 ( .A(n8092), .B(n8093), .Z(n8080) );
  AND U7594 ( .A(n8094), .B(n8095), .Z(n8093) );
  XOR U7595 ( .A(n8092), .B(n6281), .Z(n8095) );
  XOR U7596 ( .A(n8096), .B(n8097), .Z(n6281) );
  AND U7597 ( .A(n455), .B(n8098), .Z(n8097) );
  XOR U7598 ( .A(n8099), .B(n8096), .Z(n8098) );
  XNOR U7599 ( .A(n6278), .B(n8092), .Z(n8094) );
  XOR U7600 ( .A(n8100), .B(n8101), .Z(n6278) );
  AND U7601 ( .A(n452), .B(n8102), .Z(n8101) );
  XOR U7602 ( .A(n8103), .B(n8100), .Z(n8102) );
  XOR U7603 ( .A(n8104), .B(n8105), .Z(n8092) );
  AND U7604 ( .A(n8106), .B(n8107), .Z(n8105) );
  XNOR U7605 ( .A(n8108), .B(n6294), .Z(n8107) );
  XOR U7606 ( .A(n8109), .B(n8110), .Z(n6294) );
  AND U7607 ( .A(n455), .B(n8111), .Z(n8110) );
  XOR U7608 ( .A(n8109), .B(n8112), .Z(n8111) );
  XNOR U7609 ( .A(n6291), .B(n8104), .Z(n8106) );
  XOR U7610 ( .A(n8113), .B(n8114), .Z(n6291) );
  AND U7611 ( .A(n452), .B(n8115), .Z(n8114) );
  XOR U7612 ( .A(n8113), .B(n8116), .Z(n8115) );
  IV U7613 ( .A(n8108), .Z(n8104) );
  AND U7614 ( .A(n7740), .B(n7743), .Z(n8108) );
  XNOR U7615 ( .A(n8117), .B(n8118), .Z(n7743) );
  AND U7616 ( .A(n455), .B(n8119), .Z(n8118) );
  XNOR U7617 ( .A(n8120), .B(n8117), .Z(n8119) );
  XOR U7618 ( .A(n8121), .B(n8122), .Z(n455) );
  AND U7619 ( .A(n8123), .B(n8124), .Z(n8122) );
  XOR U7620 ( .A(n7751), .B(n8121), .Z(n8124) );
  IV U7621 ( .A(n8125), .Z(n7751) );
  AND U7622 ( .A(p_input[7423]), .B(p_input[7391]), .Z(n8125) );
  XOR U7623 ( .A(n8121), .B(n7748), .Z(n8123) );
  AND U7624 ( .A(p_input[7327]), .B(p_input[7359]), .Z(n7748) );
  XOR U7625 ( .A(n8126), .B(n8127), .Z(n8121) );
  AND U7626 ( .A(n8128), .B(n8129), .Z(n8127) );
  XOR U7627 ( .A(n8126), .B(n7763), .Z(n8129) );
  XNOR U7628 ( .A(p_input[7390]), .B(n8130), .Z(n7763) );
  AND U7629 ( .A(n227), .B(n8131), .Z(n8130) );
  XOR U7630 ( .A(p_input[7422]), .B(p_input[7390]), .Z(n8131) );
  XNOR U7631 ( .A(n7760), .B(n8126), .Z(n8128) );
  XOR U7632 ( .A(n8132), .B(n8133), .Z(n7760) );
  AND U7633 ( .A(n225), .B(n8134), .Z(n8133) );
  XOR U7634 ( .A(p_input[7358]), .B(p_input[7326]), .Z(n8134) );
  XOR U7635 ( .A(n8135), .B(n8136), .Z(n8126) );
  AND U7636 ( .A(n8137), .B(n8138), .Z(n8136) );
  XOR U7637 ( .A(n8135), .B(n7775), .Z(n8138) );
  XNOR U7638 ( .A(p_input[7389]), .B(n8139), .Z(n7775) );
  AND U7639 ( .A(n227), .B(n8140), .Z(n8139) );
  XOR U7640 ( .A(p_input[7421]), .B(p_input[7389]), .Z(n8140) );
  XNOR U7641 ( .A(n7772), .B(n8135), .Z(n8137) );
  XOR U7642 ( .A(n8141), .B(n8142), .Z(n7772) );
  AND U7643 ( .A(n225), .B(n8143), .Z(n8142) );
  XOR U7644 ( .A(p_input[7357]), .B(p_input[7325]), .Z(n8143) );
  XOR U7645 ( .A(n8144), .B(n8145), .Z(n8135) );
  AND U7646 ( .A(n8146), .B(n8147), .Z(n8145) );
  XOR U7647 ( .A(n8144), .B(n7787), .Z(n8147) );
  XNOR U7648 ( .A(p_input[7388]), .B(n8148), .Z(n7787) );
  AND U7649 ( .A(n227), .B(n8149), .Z(n8148) );
  XOR U7650 ( .A(p_input[7420]), .B(p_input[7388]), .Z(n8149) );
  XNOR U7651 ( .A(n7784), .B(n8144), .Z(n8146) );
  XOR U7652 ( .A(n8150), .B(n8151), .Z(n7784) );
  AND U7653 ( .A(n225), .B(n8152), .Z(n8151) );
  XOR U7654 ( .A(p_input[7356]), .B(p_input[7324]), .Z(n8152) );
  XOR U7655 ( .A(n8153), .B(n8154), .Z(n8144) );
  AND U7656 ( .A(n8155), .B(n8156), .Z(n8154) );
  XOR U7657 ( .A(n8153), .B(n7799), .Z(n8156) );
  XNOR U7658 ( .A(p_input[7387]), .B(n8157), .Z(n7799) );
  AND U7659 ( .A(n227), .B(n8158), .Z(n8157) );
  XOR U7660 ( .A(p_input[7419]), .B(p_input[7387]), .Z(n8158) );
  XNOR U7661 ( .A(n7796), .B(n8153), .Z(n8155) );
  XOR U7662 ( .A(n8159), .B(n8160), .Z(n7796) );
  AND U7663 ( .A(n225), .B(n8161), .Z(n8160) );
  XOR U7664 ( .A(p_input[7355]), .B(p_input[7323]), .Z(n8161) );
  XOR U7665 ( .A(n8162), .B(n8163), .Z(n8153) );
  AND U7666 ( .A(n8164), .B(n8165), .Z(n8163) );
  XOR U7667 ( .A(n8162), .B(n7811), .Z(n8165) );
  XNOR U7668 ( .A(p_input[7386]), .B(n8166), .Z(n7811) );
  AND U7669 ( .A(n227), .B(n8167), .Z(n8166) );
  XOR U7670 ( .A(p_input[7418]), .B(p_input[7386]), .Z(n8167) );
  XNOR U7671 ( .A(n7808), .B(n8162), .Z(n8164) );
  XOR U7672 ( .A(n8168), .B(n8169), .Z(n7808) );
  AND U7673 ( .A(n225), .B(n8170), .Z(n8169) );
  XOR U7674 ( .A(p_input[7354]), .B(p_input[7322]), .Z(n8170) );
  XOR U7675 ( .A(n8171), .B(n8172), .Z(n8162) );
  AND U7676 ( .A(n8173), .B(n8174), .Z(n8172) );
  XOR U7677 ( .A(n8171), .B(n7823), .Z(n8174) );
  XNOR U7678 ( .A(p_input[7385]), .B(n8175), .Z(n7823) );
  AND U7679 ( .A(n227), .B(n8176), .Z(n8175) );
  XOR U7680 ( .A(p_input[7417]), .B(p_input[7385]), .Z(n8176) );
  XNOR U7681 ( .A(n7820), .B(n8171), .Z(n8173) );
  XOR U7682 ( .A(n8177), .B(n8178), .Z(n7820) );
  AND U7683 ( .A(n225), .B(n8179), .Z(n8178) );
  XOR U7684 ( .A(p_input[7353]), .B(p_input[7321]), .Z(n8179) );
  XOR U7685 ( .A(n8180), .B(n8181), .Z(n8171) );
  AND U7686 ( .A(n8182), .B(n8183), .Z(n8181) );
  XOR U7687 ( .A(n8180), .B(n7835), .Z(n8183) );
  XNOR U7688 ( .A(p_input[7384]), .B(n8184), .Z(n7835) );
  AND U7689 ( .A(n227), .B(n8185), .Z(n8184) );
  XOR U7690 ( .A(p_input[7416]), .B(p_input[7384]), .Z(n8185) );
  XNOR U7691 ( .A(n7832), .B(n8180), .Z(n8182) );
  XOR U7692 ( .A(n8186), .B(n8187), .Z(n7832) );
  AND U7693 ( .A(n225), .B(n8188), .Z(n8187) );
  XOR U7694 ( .A(p_input[7352]), .B(p_input[7320]), .Z(n8188) );
  XOR U7695 ( .A(n8189), .B(n8190), .Z(n8180) );
  AND U7696 ( .A(n8191), .B(n8192), .Z(n8190) );
  XOR U7697 ( .A(n8189), .B(n7847), .Z(n8192) );
  XNOR U7698 ( .A(p_input[7383]), .B(n8193), .Z(n7847) );
  AND U7699 ( .A(n227), .B(n8194), .Z(n8193) );
  XOR U7700 ( .A(p_input[7415]), .B(p_input[7383]), .Z(n8194) );
  XNOR U7701 ( .A(n7844), .B(n8189), .Z(n8191) );
  XOR U7702 ( .A(n8195), .B(n8196), .Z(n7844) );
  AND U7703 ( .A(n225), .B(n8197), .Z(n8196) );
  XOR U7704 ( .A(p_input[7351]), .B(p_input[7319]), .Z(n8197) );
  XOR U7705 ( .A(n8198), .B(n8199), .Z(n8189) );
  AND U7706 ( .A(n8200), .B(n8201), .Z(n8199) );
  XOR U7707 ( .A(n8198), .B(n7859), .Z(n8201) );
  XNOR U7708 ( .A(p_input[7382]), .B(n8202), .Z(n7859) );
  AND U7709 ( .A(n227), .B(n8203), .Z(n8202) );
  XOR U7710 ( .A(p_input[7414]), .B(p_input[7382]), .Z(n8203) );
  XNOR U7711 ( .A(n7856), .B(n8198), .Z(n8200) );
  XOR U7712 ( .A(n8204), .B(n8205), .Z(n7856) );
  AND U7713 ( .A(n225), .B(n8206), .Z(n8205) );
  XOR U7714 ( .A(p_input[7350]), .B(p_input[7318]), .Z(n8206) );
  XOR U7715 ( .A(n8207), .B(n8208), .Z(n8198) );
  AND U7716 ( .A(n8209), .B(n8210), .Z(n8208) );
  XOR U7717 ( .A(n8207), .B(n7871), .Z(n8210) );
  XNOR U7718 ( .A(p_input[7381]), .B(n8211), .Z(n7871) );
  AND U7719 ( .A(n227), .B(n8212), .Z(n8211) );
  XOR U7720 ( .A(p_input[7413]), .B(p_input[7381]), .Z(n8212) );
  XNOR U7721 ( .A(n7868), .B(n8207), .Z(n8209) );
  XOR U7722 ( .A(n8213), .B(n8214), .Z(n7868) );
  AND U7723 ( .A(n225), .B(n8215), .Z(n8214) );
  XOR U7724 ( .A(p_input[7349]), .B(p_input[7317]), .Z(n8215) );
  XOR U7725 ( .A(n8216), .B(n8217), .Z(n8207) );
  AND U7726 ( .A(n8218), .B(n8219), .Z(n8217) );
  XOR U7727 ( .A(n8216), .B(n7883), .Z(n8219) );
  XNOR U7728 ( .A(p_input[7380]), .B(n8220), .Z(n7883) );
  AND U7729 ( .A(n227), .B(n8221), .Z(n8220) );
  XOR U7730 ( .A(p_input[7412]), .B(p_input[7380]), .Z(n8221) );
  XNOR U7731 ( .A(n7880), .B(n8216), .Z(n8218) );
  XOR U7732 ( .A(n8222), .B(n8223), .Z(n7880) );
  AND U7733 ( .A(n225), .B(n8224), .Z(n8223) );
  XOR U7734 ( .A(p_input[7348]), .B(p_input[7316]), .Z(n8224) );
  XOR U7735 ( .A(n8225), .B(n8226), .Z(n8216) );
  AND U7736 ( .A(n8227), .B(n8228), .Z(n8226) );
  XOR U7737 ( .A(n8225), .B(n7895), .Z(n8228) );
  XNOR U7738 ( .A(p_input[7379]), .B(n8229), .Z(n7895) );
  AND U7739 ( .A(n227), .B(n8230), .Z(n8229) );
  XOR U7740 ( .A(p_input[7411]), .B(p_input[7379]), .Z(n8230) );
  XNOR U7741 ( .A(n7892), .B(n8225), .Z(n8227) );
  XOR U7742 ( .A(n8231), .B(n8232), .Z(n7892) );
  AND U7743 ( .A(n225), .B(n8233), .Z(n8232) );
  XOR U7744 ( .A(p_input[7347]), .B(p_input[7315]), .Z(n8233) );
  XOR U7745 ( .A(n8234), .B(n8235), .Z(n8225) );
  AND U7746 ( .A(n8236), .B(n8237), .Z(n8235) );
  XOR U7747 ( .A(n8234), .B(n7907), .Z(n8237) );
  XNOR U7748 ( .A(p_input[7378]), .B(n8238), .Z(n7907) );
  AND U7749 ( .A(n227), .B(n8239), .Z(n8238) );
  XOR U7750 ( .A(p_input[7410]), .B(p_input[7378]), .Z(n8239) );
  XNOR U7751 ( .A(n7904), .B(n8234), .Z(n8236) );
  XOR U7752 ( .A(n8240), .B(n8241), .Z(n7904) );
  AND U7753 ( .A(n225), .B(n8242), .Z(n8241) );
  XOR U7754 ( .A(p_input[7346]), .B(p_input[7314]), .Z(n8242) );
  XOR U7755 ( .A(n8243), .B(n8244), .Z(n8234) );
  AND U7756 ( .A(n8245), .B(n8246), .Z(n8244) );
  XOR U7757 ( .A(n8243), .B(n7919), .Z(n8246) );
  XNOR U7758 ( .A(p_input[7377]), .B(n8247), .Z(n7919) );
  AND U7759 ( .A(n227), .B(n8248), .Z(n8247) );
  XOR U7760 ( .A(p_input[7409]), .B(p_input[7377]), .Z(n8248) );
  XNOR U7761 ( .A(n7916), .B(n8243), .Z(n8245) );
  XOR U7762 ( .A(n8249), .B(n8250), .Z(n7916) );
  AND U7763 ( .A(n225), .B(n8251), .Z(n8250) );
  XOR U7764 ( .A(p_input[7345]), .B(p_input[7313]), .Z(n8251) );
  XOR U7765 ( .A(n8252), .B(n8253), .Z(n8243) );
  AND U7766 ( .A(n8254), .B(n8255), .Z(n8253) );
  XOR U7767 ( .A(n8252), .B(n7931), .Z(n8255) );
  XNOR U7768 ( .A(p_input[7376]), .B(n8256), .Z(n7931) );
  AND U7769 ( .A(n227), .B(n8257), .Z(n8256) );
  XOR U7770 ( .A(p_input[7408]), .B(p_input[7376]), .Z(n8257) );
  XNOR U7771 ( .A(n7928), .B(n8252), .Z(n8254) );
  XOR U7772 ( .A(n8258), .B(n8259), .Z(n7928) );
  AND U7773 ( .A(n225), .B(n8260), .Z(n8259) );
  XOR U7774 ( .A(p_input[7344]), .B(p_input[7312]), .Z(n8260) );
  XOR U7775 ( .A(n8261), .B(n8262), .Z(n8252) );
  AND U7776 ( .A(n8263), .B(n8264), .Z(n8262) );
  XOR U7777 ( .A(n8261), .B(n7943), .Z(n8264) );
  XNOR U7778 ( .A(p_input[7375]), .B(n8265), .Z(n7943) );
  AND U7779 ( .A(n227), .B(n8266), .Z(n8265) );
  XOR U7780 ( .A(p_input[7407]), .B(p_input[7375]), .Z(n8266) );
  XNOR U7781 ( .A(n7940), .B(n8261), .Z(n8263) );
  XOR U7782 ( .A(n8267), .B(n8268), .Z(n7940) );
  AND U7783 ( .A(n225), .B(n8269), .Z(n8268) );
  XOR U7784 ( .A(p_input[7343]), .B(p_input[7311]), .Z(n8269) );
  XOR U7785 ( .A(n8270), .B(n8271), .Z(n8261) );
  AND U7786 ( .A(n8272), .B(n8273), .Z(n8271) );
  XOR U7787 ( .A(n8270), .B(n7955), .Z(n8273) );
  XNOR U7788 ( .A(p_input[7374]), .B(n8274), .Z(n7955) );
  AND U7789 ( .A(n227), .B(n8275), .Z(n8274) );
  XOR U7790 ( .A(p_input[7406]), .B(p_input[7374]), .Z(n8275) );
  XNOR U7791 ( .A(n7952), .B(n8270), .Z(n8272) );
  XOR U7792 ( .A(n8276), .B(n8277), .Z(n7952) );
  AND U7793 ( .A(n225), .B(n8278), .Z(n8277) );
  XOR U7794 ( .A(p_input[7342]), .B(p_input[7310]), .Z(n8278) );
  XOR U7795 ( .A(n8279), .B(n8280), .Z(n8270) );
  AND U7796 ( .A(n8281), .B(n8282), .Z(n8280) );
  XOR U7797 ( .A(n8279), .B(n7967), .Z(n8282) );
  XNOR U7798 ( .A(p_input[7373]), .B(n8283), .Z(n7967) );
  AND U7799 ( .A(n227), .B(n8284), .Z(n8283) );
  XOR U7800 ( .A(p_input[7405]), .B(p_input[7373]), .Z(n8284) );
  XNOR U7801 ( .A(n7964), .B(n8279), .Z(n8281) );
  XOR U7802 ( .A(n8285), .B(n8286), .Z(n7964) );
  AND U7803 ( .A(n225), .B(n8287), .Z(n8286) );
  XOR U7804 ( .A(p_input[7341]), .B(p_input[7309]), .Z(n8287) );
  XOR U7805 ( .A(n8288), .B(n8289), .Z(n8279) );
  AND U7806 ( .A(n8290), .B(n8291), .Z(n8289) );
  XOR U7807 ( .A(n8288), .B(n7979), .Z(n8291) );
  XNOR U7808 ( .A(p_input[7372]), .B(n8292), .Z(n7979) );
  AND U7809 ( .A(n227), .B(n8293), .Z(n8292) );
  XOR U7810 ( .A(p_input[7404]), .B(p_input[7372]), .Z(n8293) );
  XNOR U7811 ( .A(n7976), .B(n8288), .Z(n8290) );
  XOR U7812 ( .A(n8294), .B(n8295), .Z(n7976) );
  AND U7813 ( .A(n225), .B(n8296), .Z(n8295) );
  XOR U7814 ( .A(p_input[7340]), .B(p_input[7308]), .Z(n8296) );
  XOR U7815 ( .A(n8297), .B(n8298), .Z(n8288) );
  AND U7816 ( .A(n8299), .B(n8300), .Z(n8298) );
  XOR U7817 ( .A(n8297), .B(n7991), .Z(n8300) );
  XNOR U7818 ( .A(p_input[7371]), .B(n8301), .Z(n7991) );
  AND U7819 ( .A(n227), .B(n8302), .Z(n8301) );
  XOR U7820 ( .A(p_input[7403]), .B(p_input[7371]), .Z(n8302) );
  XNOR U7821 ( .A(n7988), .B(n8297), .Z(n8299) );
  XOR U7822 ( .A(n8303), .B(n8304), .Z(n7988) );
  AND U7823 ( .A(n225), .B(n8305), .Z(n8304) );
  XOR U7824 ( .A(p_input[7339]), .B(p_input[7307]), .Z(n8305) );
  XOR U7825 ( .A(n8306), .B(n8307), .Z(n8297) );
  AND U7826 ( .A(n8308), .B(n8309), .Z(n8307) );
  XOR U7827 ( .A(n8306), .B(n8003), .Z(n8309) );
  XNOR U7828 ( .A(p_input[7370]), .B(n8310), .Z(n8003) );
  AND U7829 ( .A(n227), .B(n8311), .Z(n8310) );
  XOR U7830 ( .A(p_input[7402]), .B(p_input[7370]), .Z(n8311) );
  XNOR U7831 ( .A(n8000), .B(n8306), .Z(n8308) );
  XOR U7832 ( .A(n8312), .B(n8313), .Z(n8000) );
  AND U7833 ( .A(n225), .B(n8314), .Z(n8313) );
  XOR U7834 ( .A(p_input[7338]), .B(p_input[7306]), .Z(n8314) );
  XOR U7835 ( .A(n8315), .B(n8316), .Z(n8306) );
  AND U7836 ( .A(n8317), .B(n8318), .Z(n8316) );
  XOR U7837 ( .A(n8315), .B(n8015), .Z(n8318) );
  XNOR U7838 ( .A(p_input[7369]), .B(n8319), .Z(n8015) );
  AND U7839 ( .A(n227), .B(n8320), .Z(n8319) );
  XOR U7840 ( .A(p_input[7401]), .B(p_input[7369]), .Z(n8320) );
  XNOR U7841 ( .A(n8012), .B(n8315), .Z(n8317) );
  XOR U7842 ( .A(n8321), .B(n8322), .Z(n8012) );
  AND U7843 ( .A(n225), .B(n8323), .Z(n8322) );
  XOR U7844 ( .A(p_input[7337]), .B(p_input[7305]), .Z(n8323) );
  XOR U7845 ( .A(n8324), .B(n8325), .Z(n8315) );
  AND U7846 ( .A(n8326), .B(n8327), .Z(n8325) );
  XOR U7847 ( .A(n8324), .B(n8027), .Z(n8327) );
  XNOR U7848 ( .A(p_input[7368]), .B(n8328), .Z(n8027) );
  AND U7849 ( .A(n227), .B(n8329), .Z(n8328) );
  XOR U7850 ( .A(p_input[7400]), .B(p_input[7368]), .Z(n8329) );
  XNOR U7851 ( .A(n8024), .B(n8324), .Z(n8326) );
  XOR U7852 ( .A(n8330), .B(n8331), .Z(n8024) );
  AND U7853 ( .A(n225), .B(n8332), .Z(n8331) );
  XOR U7854 ( .A(p_input[7336]), .B(p_input[7304]), .Z(n8332) );
  XOR U7855 ( .A(n8333), .B(n8334), .Z(n8324) );
  AND U7856 ( .A(n8335), .B(n8336), .Z(n8334) );
  XOR U7857 ( .A(n8333), .B(n8039), .Z(n8336) );
  XNOR U7858 ( .A(p_input[7367]), .B(n8337), .Z(n8039) );
  AND U7859 ( .A(n227), .B(n8338), .Z(n8337) );
  XOR U7860 ( .A(p_input[7399]), .B(p_input[7367]), .Z(n8338) );
  XNOR U7861 ( .A(n8036), .B(n8333), .Z(n8335) );
  XOR U7862 ( .A(n8339), .B(n8340), .Z(n8036) );
  AND U7863 ( .A(n225), .B(n8341), .Z(n8340) );
  XOR U7864 ( .A(p_input[7335]), .B(p_input[7303]), .Z(n8341) );
  XOR U7865 ( .A(n8342), .B(n8343), .Z(n8333) );
  AND U7866 ( .A(n8344), .B(n8345), .Z(n8343) );
  XOR U7867 ( .A(n8342), .B(n8051), .Z(n8345) );
  XNOR U7868 ( .A(p_input[7366]), .B(n8346), .Z(n8051) );
  AND U7869 ( .A(n227), .B(n8347), .Z(n8346) );
  XOR U7870 ( .A(p_input[7398]), .B(p_input[7366]), .Z(n8347) );
  XNOR U7871 ( .A(n8048), .B(n8342), .Z(n8344) );
  XOR U7872 ( .A(n8348), .B(n8349), .Z(n8048) );
  AND U7873 ( .A(n225), .B(n8350), .Z(n8349) );
  XOR U7874 ( .A(p_input[7334]), .B(p_input[7302]), .Z(n8350) );
  XOR U7875 ( .A(n8351), .B(n8352), .Z(n8342) );
  AND U7876 ( .A(n8353), .B(n8354), .Z(n8352) );
  XOR U7877 ( .A(n8351), .B(n8063), .Z(n8354) );
  XNOR U7878 ( .A(p_input[7365]), .B(n8355), .Z(n8063) );
  AND U7879 ( .A(n227), .B(n8356), .Z(n8355) );
  XOR U7880 ( .A(p_input[7397]), .B(p_input[7365]), .Z(n8356) );
  XNOR U7881 ( .A(n8060), .B(n8351), .Z(n8353) );
  XOR U7882 ( .A(n8357), .B(n8358), .Z(n8060) );
  AND U7883 ( .A(n225), .B(n8359), .Z(n8358) );
  XOR U7884 ( .A(p_input[7333]), .B(p_input[7301]), .Z(n8359) );
  XOR U7885 ( .A(n8360), .B(n8361), .Z(n8351) );
  AND U7886 ( .A(n8362), .B(n8363), .Z(n8361) );
  XOR U7887 ( .A(n8360), .B(n8075), .Z(n8363) );
  XNOR U7888 ( .A(p_input[7364]), .B(n8364), .Z(n8075) );
  AND U7889 ( .A(n227), .B(n8365), .Z(n8364) );
  XOR U7890 ( .A(p_input[7396]), .B(p_input[7364]), .Z(n8365) );
  XNOR U7891 ( .A(n8072), .B(n8360), .Z(n8362) );
  XOR U7892 ( .A(n8366), .B(n8367), .Z(n8072) );
  AND U7893 ( .A(n225), .B(n8368), .Z(n8367) );
  XOR U7894 ( .A(p_input[7332]), .B(p_input[7300]), .Z(n8368) );
  XOR U7895 ( .A(n8369), .B(n8370), .Z(n8360) );
  AND U7896 ( .A(n8371), .B(n8372), .Z(n8370) );
  XOR U7897 ( .A(n8369), .B(n8087), .Z(n8372) );
  XNOR U7898 ( .A(p_input[7363]), .B(n8373), .Z(n8087) );
  AND U7899 ( .A(n227), .B(n8374), .Z(n8373) );
  XOR U7900 ( .A(p_input[7395]), .B(p_input[7363]), .Z(n8374) );
  XNOR U7901 ( .A(n8084), .B(n8369), .Z(n8371) );
  XOR U7902 ( .A(n8375), .B(n8376), .Z(n8084) );
  AND U7903 ( .A(n225), .B(n8377), .Z(n8376) );
  XOR U7904 ( .A(p_input[7331]), .B(p_input[7299]), .Z(n8377) );
  XOR U7905 ( .A(n8378), .B(n8379), .Z(n8369) );
  AND U7906 ( .A(n8380), .B(n8381), .Z(n8379) );
  XOR U7907 ( .A(n8378), .B(n8099), .Z(n8381) );
  XNOR U7908 ( .A(p_input[7362]), .B(n8382), .Z(n8099) );
  AND U7909 ( .A(n227), .B(n8383), .Z(n8382) );
  XOR U7910 ( .A(p_input[7394]), .B(p_input[7362]), .Z(n8383) );
  XNOR U7911 ( .A(n8096), .B(n8378), .Z(n8380) );
  XOR U7912 ( .A(n8384), .B(n8385), .Z(n8096) );
  AND U7913 ( .A(n225), .B(n8386), .Z(n8385) );
  XOR U7914 ( .A(p_input[7330]), .B(p_input[7298]), .Z(n8386) );
  XOR U7915 ( .A(n8387), .B(n8388), .Z(n8378) );
  AND U7916 ( .A(n8389), .B(n8390), .Z(n8388) );
  XNOR U7917 ( .A(n8391), .B(n8112), .Z(n8390) );
  XNOR U7918 ( .A(p_input[7361]), .B(n8392), .Z(n8112) );
  AND U7919 ( .A(n227), .B(n8393), .Z(n8392) );
  XNOR U7920 ( .A(p_input[7393]), .B(n8394), .Z(n8393) );
  IV U7921 ( .A(p_input[7361]), .Z(n8394) );
  XNOR U7922 ( .A(n8109), .B(n8387), .Z(n8389) );
  XNOR U7923 ( .A(p_input[7297]), .B(n8395), .Z(n8109) );
  AND U7924 ( .A(n225), .B(n8396), .Z(n8395) );
  XOR U7925 ( .A(p_input[7329]), .B(p_input[7297]), .Z(n8396) );
  IV U7926 ( .A(n8391), .Z(n8387) );
  AND U7927 ( .A(n8117), .B(n8120), .Z(n8391) );
  XOR U7928 ( .A(p_input[7360]), .B(n8397), .Z(n8120) );
  AND U7929 ( .A(n227), .B(n8398), .Z(n8397) );
  XOR U7930 ( .A(p_input[7392]), .B(p_input[7360]), .Z(n8398) );
  XOR U7931 ( .A(n8399), .B(n8400), .Z(n227) );
  AND U7932 ( .A(n8401), .B(n8402), .Z(n8400) );
  XNOR U7933 ( .A(p_input[7423]), .B(n8399), .Z(n8402) );
  XOR U7934 ( .A(n8399), .B(p_input[7391]), .Z(n8401) );
  XOR U7935 ( .A(n8403), .B(n8404), .Z(n8399) );
  AND U7936 ( .A(n8405), .B(n8406), .Z(n8404) );
  XNOR U7937 ( .A(p_input[7422]), .B(n8403), .Z(n8406) );
  XOR U7938 ( .A(n8403), .B(p_input[7390]), .Z(n8405) );
  XOR U7939 ( .A(n8407), .B(n8408), .Z(n8403) );
  AND U7940 ( .A(n8409), .B(n8410), .Z(n8408) );
  XNOR U7941 ( .A(p_input[7421]), .B(n8407), .Z(n8410) );
  XOR U7942 ( .A(n8407), .B(p_input[7389]), .Z(n8409) );
  XOR U7943 ( .A(n8411), .B(n8412), .Z(n8407) );
  AND U7944 ( .A(n8413), .B(n8414), .Z(n8412) );
  XNOR U7945 ( .A(p_input[7420]), .B(n8411), .Z(n8414) );
  XOR U7946 ( .A(n8411), .B(p_input[7388]), .Z(n8413) );
  XOR U7947 ( .A(n8415), .B(n8416), .Z(n8411) );
  AND U7948 ( .A(n8417), .B(n8418), .Z(n8416) );
  XNOR U7949 ( .A(p_input[7419]), .B(n8415), .Z(n8418) );
  XOR U7950 ( .A(n8415), .B(p_input[7387]), .Z(n8417) );
  XOR U7951 ( .A(n8419), .B(n8420), .Z(n8415) );
  AND U7952 ( .A(n8421), .B(n8422), .Z(n8420) );
  XNOR U7953 ( .A(p_input[7418]), .B(n8419), .Z(n8422) );
  XOR U7954 ( .A(n8419), .B(p_input[7386]), .Z(n8421) );
  XOR U7955 ( .A(n8423), .B(n8424), .Z(n8419) );
  AND U7956 ( .A(n8425), .B(n8426), .Z(n8424) );
  XNOR U7957 ( .A(p_input[7417]), .B(n8423), .Z(n8426) );
  XOR U7958 ( .A(n8423), .B(p_input[7385]), .Z(n8425) );
  XOR U7959 ( .A(n8427), .B(n8428), .Z(n8423) );
  AND U7960 ( .A(n8429), .B(n8430), .Z(n8428) );
  XNOR U7961 ( .A(p_input[7416]), .B(n8427), .Z(n8430) );
  XOR U7962 ( .A(n8427), .B(p_input[7384]), .Z(n8429) );
  XOR U7963 ( .A(n8431), .B(n8432), .Z(n8427) );
  AND U7964 ( .A(n8433), .B(n8434), .Z(n8432) );
  XNOR U7965 ( .A(p_input[7415]), .B(n8431), .Z(n8434) );
  XOR U7966 ( .A(n8431), .B(p_input[7383]), .Z(n8433) );
  XOR U7967 ( .A(n8435), .B(n8436), .Z(n8431) );
  AND U7968 ( .A(n8437), .B(n8438), .Z(n8436) );
  XNOR U7969 ( .A(p_input[7414]), .B(n8435), .Z(n8438) );
  XOR U7970 ( .A(n8435), .B(p_input[7382]), .Z(n8437) );
  XOR U7971 ( .A(n8439), .B(n8440), .Z(n8435) );
  AND U7972 ( .A(n8441), .B(n8442), .Z(n8440) );
  XNOR U7973 ( .A(p_input[7413]), .B(n8439), .Z(n8442) );
  XOR U7974 ( .A(n8439), .B(p_input[7381]), .Z(n8441) );
  XOR U7975 ( .A(n8443), .B(n8444), .Z(n8439) );
  AND U7976 ( .A(n8445), .B(n8446), .Z(n8444) );
  XNOR U7977 ( .A(p_input[7412]), .B(n8443), .Z(n8446) );
  XOR U7978 ( .A(n8443), .B(p_input[7380]), .Z(n8445) );
  XOR U7979 ( .A(n8447), .B(n8448), .Z(n8443) );
  AND U7980 ( .A(n8449), .B(n8450), .Z(n8448) );
  XNOR U7981 ( .A(p_input[7411]), .B(n8447), .Z(n8450) );
  XOR U7982 ( .A(n8447), .B(p_input[7379]), .Z(n8449) );
  XOR U7983 ( .A(n8451), .B(n8452), .Z(n8447) );
  AND U7984 ( .A(n8453), .B(n8454), .Z(n8452) );
  XNOR U7985 ( .A(p_input[7410]), .B(n8451), .Z(n8454) );
  XOR U7986 ( .A(n8451), .B(p_input[7378]), .Z(n8453) );
  XOR U7987 ( .A(n8455), .B(n8456), .Z(n8451) );
  AND U7988 ( .A(n8457), .B(n8458), .Z(n8456) );
  XNOR U7989 ( .A(p_input[7409]), .B(n8455), .Z(n8458) );
  XOR U7990 ( .A(n8455), .B(p_input[7377]), .Z(n8457) );
  XOR U7991 ( .A(n8459), .B(n8460), .Z(n8455) );
  AND U7992 ( .A(n8461), .B(n8462), .Z(n8460) );
  XNOR U7993 ( .A(p_input[7408]), .B(n8459), .Z(n8462) );
  XOR U7994 ( .A(n8459), .B(p_input[7376]), .Z(n8461) );
  XOR U7995 ( .A(n8463), .B(n8464), .Z(n8459) );
  AND U7996 ( .A(n8465), .B(n8466), .Z(n8464) );
  XNOR U7997 ( .A(p_input[7407]), .B(n8463), .Z(n8466) );
  XOR U7998 ( .A(n8463), .B(p_input[7375]), .Z(n8465) );
  XOR U7999 ( .A(n8467), .B(n8468), .Z(n8463) );
  AND U8000 ( .A(n8469), .B(n8470), .Z(n8468) );
  XNOR U8001 ( .A(p_input[7406]), .B(n8467), .Z(n8470) );
  XOR U8002 ( .A(n8467), .B(p_input[7374]), .Z(n8469) );
  XOR U8003 ( .A(n8471), .B(n8472), .Z(n8467) );
  AND U8004 ( .A(n8473), .B(n8474), .Z(n8472) );
  XNOR U8005 ( .A(p_input[7405]), .B(n8471), .Z(n8474) );
  XOR U8006 ( .A(n8471), .B(p_input[7373]), .Z(n8473) );
  XOR U8007 ( .A(n8475), .B(n8476), .Z(n8471) );
  AND U8008 ( .A(n8477), .B(n8478), .Z(n8476) );
  XNOR U8009 ( .A(p_input[7404]), .B(n8475), .Z(n8478) );
  XOR U8010 ( .A(n8475), .B(p_input[7372]), .Z(n8477) );
  XOR U8011 ( .A(n8479), .B(n8480), .Z(n8475) );
  AND U8012 ( .A(n8481), .B(n8482), .Z(n8480) );
  XNOR U8013 ( .A(p_input[7403]), .B(n8479), .Z(n8482) );
  XOR U8014 ( .A(n8479), .B(p_input[7371]), .Z(n8481) );
  XOR U8015 ( .A(n8483), .B(n8484), .Z(n8479) );
  AND U8016 ( .A(n8485), .B(n8486), .Z(n8484) );
  XNOR U8017 ( .A(p_input[7402]), .B(n8483), .Z(n8486) );
  XOR U8018 ( .A(n8483), .B(p_input[7370]), .Z(n8485) );
  XOR U8019 ( .A(n8487), .B(n8488), .Z(n8483) );
  AND U8020 ( .A(n8489), .B(n8490), .Z(n8488) );
  XNOR U8021 ( .A(p_input[7401]), .B(n8487), .Z(n8490) );
  XOR U8022 ( .A(n8487), .B(p_input[7369]), .Z(n8489) );
  XOR U8023 ( .A(n8491), .B(n8492), .Z(n8487) );
  AND U8024 ( .A(n8493), .B(n8494), .Z(n8492) );
  XNOR U8025 ( .A(p_input[7400]), .B(n8491), .Z(n8494) );
  XOR U8026 ( .A(n8491), .B(p_input[7368]), .Z(n8493) );
  XOR U8027 ( .A(n8495), .B(n8496), .Z(n8491) );
  AND U8028 ( .A(n8497), .B(n8498), .Z(n8496) );
  XNOR U8029 ( .A(p_input[7399]), .B(n8495), .Z(n8498) );
  XOR U8030 ( .A(n8495), .B(p_input[7367]), .Z(n8497) );
  XOR U8031 ( .A(n8499), .B(n8500), .Z(n8495) );
  AND U8032 ( .A(n8501), .B(n8502), .Z(n8500) );
  XNOR U8033 ( .A(p_input[7398]), .B(n8499), .Z(n8502) );
  XOR U8034 ( .A(n8499), .B(p_input[7366]), .Z(n8501) );
  XOR U8035 ( .A(n8503), .B(n8504), .Z(n8499) );
  AND U8036 ( .A(n8505), .B(n8506), .Z(n8504) );
  XNOR U8037 ( .A(p_input[7397]), .B(n8503), .Z(n8506) );
  XOR U8038 ( .A(n8503), .B(p_input[7365]), .Z(n8505) );
  XOR U8039 ( .A(n8507), .B(n8508), .Z(n8503) );
  AND U8040 ( .A(n8509), .B(n8510), .Z(n8508) );
  XNOR U8041 ( .A(p_input[7396]), .B(n8507), .Z(n8510) );
  XOR U8042 ( .A(n8507), .B(p_input[7364]), .Z(n8509) );
  XOR U8043 ( .A(n8511), .B(n8512), .Z(n8507) );
  AND U8044 ( .A(n8513), .B(n8514), .Z(n8512) );
  XNOR U8045 ( .A(p_input[7395]), .B(n8511), .Z(n8514) );
  XOR U8046 ( .A(n8511), .B(p_input[7363]), .Z(n8513) );
  XOR U8047 ( .A(n8515), .B(n8516), .Z(n8511) );
  AND U8048 ( .A(n8517), .B(n8518), .Z(n8516) );
  XNOR U8049 ( .A(p_input[7394]), .B(n8515), .Z(n8518) );
  XOR U8050 ( .A(n8515), .B(p_input[7362]), .Z(n8517) );
  XNOR U8051 ( .A(n8519), .B(n8520), .Z(n8515) );
  AND U8052 ( .A(n8521), .B(n8522), .Z(n8520) );
  XOR U8053 ( .A(p_input[7393]), .B(n8519), .Z(n8522) );
  XNOR U8054 ( .A(p_input[7361]), .B(n8519), .Z(n8521) );
  AND U8055 ( .A(p_input[7392]), .B(n8523), .Z(n8519) );
  IV U8056 ( .A(p_input[7360]), .Z(n8523) );
  XNOR U8057 ( .A(p_input[7296]), .B(n8524), .Z(n8117) );
  AND U8058 ( .A(n225), .B(n8525), .Z(n8524) );
  XOR U8059 ( .A(p_input[7328]), .B(p_input[7296]), .Z(n8525) );
  XOR U8060 ( .A(n8526), .B(n8527), .Z(n225) );
  AND U8061 ( .A(n8528), .B(n8529), .Z(n8527) );
  XNOR U8062 ( .A(p_input[7359]), .B(n8526), .Z(n8529) );
  XOR U8063 ( .A(n8526), .B(p_input[7327]), .Z(n8528) );
  XOR U8064 ( .A(n8530), .B(n8531), .Z(n8526) );
  AND U8065 ( .A(n8532), .B(n8533), .Z(n8531) );
  XNOR U8066 ( .A(p_input[7358]), .B(n8530), .Z(n8533) );
  XNOR U8067 ( .A(n8530), .B(n8132), .Z(n8532) );
  IV U8068 ( .A(p_input[7326]), .Z(n8132) );
  XOR U8069 ( .A(n8534), .B(n8535), .Z(n8530) );
  AND U8070 ( .A(n8536), .B(n8537), .Z(n8535) );
  XNOR U8071 ( .A(p_input[7357]), .B(n8534), .Z(n8537) );
  XNOR U8072 ( .A(n8534), .B(n8141), .Z(n8536) );
  IV U8073 ( .A(p_input[7325]), .Z(n8141) );
  XOR U8074 ( .A(n8538), .B(n8539), .Z(n8534) );
  AND U8075 ( .A(n8540), .B(n8541), .Z(n8539) );
  XNOR U8076 ( .A(p_input[7356]), .B(n8538), .Z(n8541) );
  XNOR U8077 ( .A(n8538), .B(n8150), .Z(n8540) );
  IV U8078 ( .A(p_input[7324]), .Z(n8150) );
  XOR U8079 ( .A(n8542), .B(n8543), .Z(n8538) );
  AND U8080 ( .A(n8544), .B(n8545), .Z(n8543) );
  XNOR U8081 ( .A(p_input[7355]), .B(n8542), .Z(n8545) );
  XNOR U8082 ( .A(n8542), .B(n8159), .Z(n8544) );
  IV U8083 ( .A(p_input[7323]), .Z(n8159) );
  XOR U8084 ( .A(n8546), .B(n8547), .Z(n8542) );
  AND U8085 ( .A(n8548), .B(n8549), .Z(n8547) );
  XNOR U8086 ( .A(p_input[7354]), .B(n8546), .Z(n8549) );
  XNOR U8087 ( .A(n8546), .B(n8168), .Z(n8548) );
  IV U8088 ( .A(p_input[7322]), .Z(n8168) );
  XOR U8089 ( .A(n8550), .B(n8551), .Z(n8546) );
  AND U8090 ( .A(n8552), .B(n8553), .Z(n8551) );
  XNOR U8091 ( .A(p_input[7353]), .B(n8550), .Z(n8553) );
  XNOR U8092 ( .A(n8550), .B(n8177), .Z(n8552) );
  IV U8093 ( .A(p_input[7321]), .Z(n8177) );
  XOR U8094 ( .A(n8554), .B(n8555), .Z(n8550) );
  AND U8095 ( .A(n8556), .B(n8557), .Z(n8555) );
  XNOR U8096 ( .A(p_input[7352]), .B(n8554), .Z(n8557) );
  XNOR U8097 ( .A(n8554), .B(n8186), .Z(n8556) );
  IV U8098 ( .A(p_input[7320]), .Z(n8186) );
  XOR U8099 ( .A(n8558), .B(n8559), .Z(n8554) );
  AND U8100 ( .A(n8560), .B(n8561), .Z(n8559) );
  XNOR U8101 ( .A(p_input[7351]), .B(n8558), .Z(n8561) );
  XNOR U8102 ( .A(n8558), .B(n8195), .Z(n8560) );
  IV U8103 ( .A(p_input[7319]), .Z(n8195) );
  XOR U8104 ( .A(n8562), .B(n8563), .Z(n8558) );
  AND U8105 ( .A(n8564), .B(n8565), .Z(n8563) );
  XNOR U8106 ( .A(p_input[7350]), .B(n8562), .Z(n8565) );
  XNOR U8107 ( .A(n8562), .B(n8204), .Z(n8564) );
  IV U8108 ( .A(p_input[7318]), .Z(n8204) );
  XOR U8109 ( .A(n8566), .B(n8567), .Z(n8562) );
  AND U8110 ( .A(n8568), .B(n8569), .Z(n8567) );
  XNOR U8111 ( .A(p_input[7349]), .B(n8566), .Z(n8569) );
  XNOR U8112 ( .A(n8566), .B(n8213), .Z(n8568) );
  IV U8113 ( .A(p_input[7317]), .Z(n8213) );
  XOR U8114 ( .A(n8570), .B(n8571), .Z(n8566) );
  AND U8115 ( .A(n8572), .B(n8573), .Z(n8571) );
  XNOR U8116 ( .A(p_input[7348]), .B(n8570), .Z(n8573) );
  XNOR U8117 ( .A(n8570), .B(n8222), .Z(n8572) );
  IV U8118 ( .A(p_input[7316]), .Z(n8222) );
  XOR U8119 ( .A(n8574), .B(n8575), .Z(n8570) );
  AND U8120 ( .A(n8576), .B(n8577), .Z(n8575) );
  XNOR U8121 ( .A(p_input[7347]), .B(n8574), .Z(n8577) );
  XNOR U8122 ( .A(n8574), .B(n8231), .Z(n8576) );
  IV U8123 ( .A(p_input[7315]), .Z(n8231) );
  XOR U8124 ( .A(n8578), .B(n8579), .Z(n8574) );
  AND U8125 ( .A(n8580), .B(n8581), .Z(n8579) );
  XNOR U8126 ( .A(p_input[7346]), .B(n8578), .Z(n8581) );
  XNOR U8127 ( .A(n8578), .B(n8240), .Z(n8580) );
  IV U8128 ( .A(p_input[7314]), .Z(n8240) );
  XOR U8129 ( .A(n8582), .B(n8583), .Z(n8578) );
  AND U8130 ( .A(n8584), .B(n8585), .Z(n8583) );
  XNOR U8131 ( .A(p_input[7345]), .B(n8582), .Z(n8585) );
  XNOR U8132 ( .A(n8582), .B(n8249), .Z(n8584) );
  IV U8133 ( .A(p_input[7313]), .Z(n8249) );
  XOR U8134 ( .A(n8586), .B(n8587), .Z(n8582) );
  AND U8135 ( .A(n8588), .B(n8589), .Z(n8587) );
  XNOR U8136 ( .A(p_input[7344]), .B(n8586), .Z(n8589) );
  XNOR U8137 ( .A(n8586), .B(n8258), .Z(n8588) );
  IV U8138 ( .A(p_input[7312]), .Z(n8258) );
  XOR U8139 ( .A(n8590), .B(n8591), .Z(n8586) );
  AND U8140 ( .A(n8592), .B(n8593), .Z(n8591) );
  XNOR U8141 ( .A(p_input[7343]), .B(n8590), .Z(n8593) );
  XNOR U8142 ( .A(n8590), .B(n8267), .Z(n8592) );
  IV U8143 ( .A(p_input[7311]), .Z(n8267) );
  XOR U8144 ( .A(n8594), .B(n8595), .Z(n8590) );
  AND U8145 ( .A(n8596), .B(n8597), .Z(n8595) );
  XNOR U8146 ( .A(p_input[7342]), .B(n8594), .Z(n8597) );
  XNOR U8147 ( .A(n8594), .B(n8276), .Z(n8596) );
  IV U8148 ( .A(p_input[7310]), .Z(n8276) );
  XOR U8149 ( .A(n8598), .B(n8599), .Z(n8594) );
  AND U8150 ( .A(n8600), .B(n8601), .Z(n8599) );
  XNOR U8151 ( .A(p_input[7341]), .B(n8598), .Z(n8601) );
  XNOR U8152 ( .A(n8598), .B(n8285), .Z(n8600) );
  IV U8153 ( .A(p_input[7309]), .Z(n8285) );
  XOR U8154 ( .A(n8602), .B(n8603), .Z(n8598) );
  AND U8155 ( .A(n8604), .B(n8605), .Z(n8603) );
  XNOR U8156 ( .A(p_input[7340]), .B(n8602), .Z(n8605) );
  XNOR U8157 ( .A(n8602), .B(n8294), .Z(n8604) );
  IV U8158 ( .A(p_input[7308]), .Z(n8294) );
  XOR U8159 ( .A(n8606), .B(n8607), .Z(n8602) );
  AND U8160 ( .A(n8608), .B(n8609), .Z(n8607) );
  XNOR U8161 ( .A(p_input[7339]), .B(n8606), .Z(n8609) );
  XNOR U8162 ( .A(n8606), .B(n8303), .Z(n8608) );
  IV U8163 ( .A(p_input[7307]), .Z(n8303) );
  XOR U8164 ( .A(n8610), .B(n8611), .Z(n8606) );
  AND U8165 ( .A(n8612), .B(n8613), .Z(n8611) );
  XNOR U8166 ( .A(p_input[7338]), .B(n8610), .Z(n8613) );
  XNOR U8167 ( .A(n8610), .B(n8312), .Z(n8612) );
  IV U8168 ( .A(p_input[7306]), .Z(n8312) );
  XOR U8169 ( .A(n8614), .B(n8615), .Z(n8610) );
  AND U8170 ( .A(n8616), .B(n8617), .Z(n8615) );
  XNOR U8171 ( .A(p_input[7337]), .B(n8614), .Z(n8617) );
  XNOR U8172 ( .A(n8614), .B(n8321), .Z(n8616) );
  IV U8173 ( .A(p_input[7305]), .Z(n8321) );
  XOR U8174 ( .A(n8618), .B(n8619), .Z(n8614) );
  AND U8175 ( .A(n8620), .B(n8621), .Z(n8619) );
  XNOR U8176 ( .A(p_input[7336]), .B(n8618), .Z(n8621) );
  XNOR U8177 ( .A(n8618), .B(n8330), .Z(n8620) );
  IV U8178 ( .A(p_input[7304]), .Z(n8330) );
  XOR U8179 ( .A(n8622), .B(n8623), .Z(n8618) );
  AND U8180 ( .A(n8624), .B(n8625), .Z(n8623) );
  XNOR U8181 ( .A(p_input[7335]), .B(n8622), .Z(n8625) );
  XNOR U8182 ( .A(n8622), .B(n8339), .Z(n8624) );
  IV U8183 ( .A(p_input[7303]), .Z(n8339) );
  XOR U8184 ( .A(n8626), .B(n8627), .Z(n8622) );
  AND U8185 ( .A(n8628), .B(n8629), .Z(n8627) );
  XNOR U8186 ( .A(p_input[7334]), .B(n8626), .Z(n8629) );
  XNOR U8187 ( .A(n8626), .B(n8348), .Z(n8628) );
  IV U8188 ( .A(p_input[7302]), .Z(n8348) );
  XOR U8189 ( .A(n8630), .B(n8631), .Z(n8626) );
  AND U8190 ( .A(n8632), .B(n8633), .Z(n8631) );
  XNOR U8191 ( .A(p_input[7333]), .B(n8630), .Z(n8633) );
  XNOR U8192 ( .A(n8630), .B(n8357), .Z(n8632) );
  IV U8193 ( .A(p_input[7301]), .Z(n8357) );
  XOR U8194 ( .A(n8634), .B(n8635), .Z(n8630) );
  AND U8195 ( .A(n8636), .B(n8637), .Z(n8635) );
  XNOR U8196 ( .A(p_input[7332]), .B(n8634), .Z(n8637) );
  XNOR U8197 ( .A(n8634), .B(n8366), .Z(n8636) );
  IV U8198 ( .A(p_input[7300]), .Z(n8366) );
  XOR U8199 ( .A(n8638), .B(n8639), .Z(n8634) );
  AND U8200 ( .A(n8640), .B(n8641), .Z(n8639) );
  XNOR U8201 ( .A(p_input[7331]), .B(n8638), .Z(n8641) );
  XNOR U8202 ( .A(n8638), .B(n8375), .Z(n8640) );
  IV U8203 ( .A(p_input[7299]), .Z(n8375) );
  XOR U8204 ( .A(n8642), .B(n8643), .Z(n8638) );
  AND U8205 ( .A(n8644), .B(n8645), .Z(n8643) );
  XNOR U8206 ( .A(p_input[7330]), .B(n8642), .Z(n8645) );
  XNOR U8207 ( .A(n8642), .B(n8384), .Z(n8644) );
  IV U8208 ( .A(p_input[7298]), .Z(n8384) );
  XNOR U8209 ( .A(n8646), .B(n8647), .Z(n8642) );
  AND U8210 ( .A(n8648), .B(n8649), .Z(n8647) );
  XOR U8211 ( .A(p_input[7329]), .B(n8646), .Z(n8649) );
  XNOR U8212 ( .A(p_input[7297]), .B(n8646), .Z(n8648) );
  AND U8213 ( .A(p_input[7328]), .B(n8650), .Z(n8646) );
  IV U8214 ( .A(p_input[7296]), .Z(n8650) );
  XOR U8215 ( .A(n8651), .B(n8652), .Z(n7740) );
  AND U8216 ( .A(n452), .B(n8653), .Z(n8652) );
  XNOR U8217 ( .A(n8654), .B(n8651), .Z(n8653) );
  XOR U8218 ( .A(n8655), .B(n8656), .Z(n452) );
  AND U8219 ( .A(n8657), .B(n8658), .Z(n8656) );
  XNOR U8220 ( .A(n7755), .B(n8655), .Z(n8658) );
  AND U8221 ( .A(p_input[7295]), .B(p_input[7263]), .Z(n7755) );
  XNOR U8222 ( .A(n8655), .B(n7752), .Z(n8657) );
  IV U8223 ( .A(n8659), .Z(n7752) );
  AND U8224 ( .A(p_input[7199]), .B(p_input[7231]), .Z(n8659) );
  XOR U8225 ( .A(n8660), .B(n8661), .Z(n8655) );
  AND U8226 ( .A(n8662), .B(n8663), .Z(n8661) );
  XOR U8227 ( .A(n8660), .B(n7767), .Z(n8663) );
  XNOR U8228 ( .A(p_input[7262]), .B(n8664), .Z(n7767) );
  AND U8229 ( .A(n231), .B(n8665), .Z(n8664) );
  XOR U8230 ( .A(p_input[7294]), .B(p_input[7262]), .Z(n8665) );
  XNOR U8231 ( .A(n7764), .B(n8660), .Z(n8662) );
  XOR U8232 ( .A(n8666), .B(n8667), .Z(n7764) );
  AND U8233 ( .A(n228), .B(n8668), .Z(n8667) );
  XOR U8234 ( .A(p_input[7230]), .B(p_input[7198]), .Z(n8668) );
  XOR U8235 ( .A(n8669), .B(n8670), .Z(n8660) );
  AND U8236 ( .A(n8671), .B(n8672), .Z(n8670) );
  XOR U8237 ( .A(n8669), .B(n7779), .Z(n8672) );
  XNOR U8238 ( .A(p_input[7261]), .B(n8673), .Z(n7779) );
  AND U8239 ( .A(n231), .B(n8674), .Z(n8673) );
  XOR U8240 ( .A(p_input[7293]), .B(p_input[7261]), .Z(n8674) );
  XNOR U8241 ( .A(n7776), .B(n8669), .Z(n8671) );
  XOR U8242 ( .A(n8675), .B(n8676), .Z(n7776) );
  AND U8243 ( .A(n228), .B(n8677), .Z(n8676) );
  XOR U8244 ( .A(p_input[7229]), .B(p_input[7197]), .Z(n8677) );
  XOR U8245 ( .A(n8678), .B(n8679), .Z(n8669) );
  AND U8246 ( .A(n8680), .B(n8681), .Z(n8679) );
  XOR U8247 ( .A(n8678), .B(n7791), .Z(n8681) );
  XNOR U8248 ( .A(p_input[7260]), .B(n8682), .Z(n7791) );
  AND U8249 ( .A(n231), .B(n8683), .Z(n8682) );
  XOR U8250 ( .A(p_input[7292]), .B(p_input[7260]), .Z(n8683) );
  XNOR U8251 ( .A(n7788), .B(n8678), .Z(n8680) );
  XOR U8252 ( .A(n8684), .B(n8685), .Z(n7788) );
  AND U8253 ( .A(n228), .B(n8686), .Z(n8685) );
  XOR U8254 ( .A(p_input[7228]), .B(p_input[7196]), .Z(n8686) );
  XOR U8255 ( .A(n8687), .B(n8688), .Z(n8678) );
  AND U8256 ( .A(n8689), .B(n8690), .Z(n8688) );
  XOR U8257 ( .A(n8687), .B(n7803), .Z(n8690) );
  XNOR U8258 ( .A(p_input[7259]), .B(n8691), .Z(n7803) );
  AND U8259 ( .A(n231), .B(n8692), .Z(n8691) );
  XOR U8260 ( .A(p_input[7291]), .B(p_input[7259]), .Z(n8692) );
  XNOR U8261 ( .A(n7800), .B(n8687), .Z(n8689) );
  XOR U8262 ( .A(n8693), .B(n8694), .Z(n7800) );
  AND U8263 ( .A(n228), .B(n8695), .Z(n8694) );
  XOR U8264 ( .A(p_input[7227]), .B(p_input[7195]), .Z(n8695) );
  XOR U8265 ( .A(n8696), .B(n8697), .Z(n8687) );
  AND U8266 ( .A(n8698), .B(n8699), .Z(n8697) );
  XOR U8267 ( .A(n8696), .B(n7815), .Z(n8699) );
  XNOR U8268 ( .A(p_input[7258]), .B(n8700), .Z(n7815) );
  AND U8269 ( .A(n231), .B(n8701), .Z(n8700) );
  XOR U8270 ( .A(p_input[7290]), .B(p_input[7258]), .Z(n8701) );
  XNOR U8271 ( .A(n7812), .B(n8696), .Z(n8698) );
  XOR U8272 ( .A(n8702), .B(n8703), .Z(n7812) );
  AND U8273 ( .A(n228), .B(n8704), .Z(n8703) );
  XOR U8274 ( .A(p_input[7226]), .B(p_input[7194]), .Z(n8704) );
  XOR U8275 ( .A(n8705), .B(n8706), .Z(n8696) );
  AND U8276 ( .A(n8707), .B(n8708), .Z(n8706) );
  XOR U8277 ( .A(n8705), .B(n7827), .Z(n8708) );
  XNOR U8278 ( .A(p_input[7257]), .B(n8709), .Z(n7827) );
  AND U8279 ( .A(n231), .B(n8710), .Z(n8709) );
  XOR U8280 ( .A(p_input[7289]), .B(p_input[7257]), .Z(n8710) );
  XNOR U8281 ( .A(n7824), .B(n8705), .Z(n8707) );
  XOR U8282 ( .A(n8711), .B(n8712), .Z(n7824) );
  AND U8283 ( .A(n228), .B(n8713), .Z(n8712) );
  XOR U8284 ( .A(p_input[7225]), .B(p_input[7193]), .Z(n8713) );
  XOR U8285 ( .A(n8714), .B(n8715), .Z(n8705) );
  AND U8286 ( .A(n8716), .B(n8717), .Z(n8715) );
  XOR U8287 ( .A(n8714), .B(n7839), .Z(n8717) );
  XNOR U8288 ( .A(p_input[7256]), .B(n8718), .Z(n7839) );
  AND U8289 ( .A(n231), .B(n8719), .Z(n8718) );
  XOR U8290 ( .A(p_input[7288]), .B(p_input[7256]), .Z(n8719) );
  XNOR U8291 ( .A(n7836), .B(n8714), .Z(n8716) );
  XOR U8292 ( .A(n8720), .B(n8721), .Z(n7836) );
  AND U8293 ( .A(n228), .B(n8722), .Z(n8721) );
  XOR U8294 ( .A(p_input[7224]), .B(p_input[7192]), .Z(n8722) );
  XOR U8295 ( .A(n8723), .B(n8724), .Z(n8714) );
  AND U8296 ( .A(n8725), .B(n8726), .Z(n8724) );
  XOR U8297 ( .A(n8723), .B(n7851), .Z(n8726) );
  XNOR U8298 ( .A(p_input[7255]), .B(n8727), .Z(n7851) );
  AND U8299 ( .A(n231), .B(n8728), .Z(n8727) );
  XOR U8300 ( .A(p_input[7287]), .B(p_input[7255]), .Z(n8728) );
  XNOR U8301 ( .A(n7848), .B(n8723), .Z(n8725) );
  XOR U8302 ( .A(n8729), .B(n8730), .Z(n7848) );
  AND U8303 ( .A(n228), .B(n8731), .Z(n8730) );
  XOR U8304 ( .A(p_input[7223]), .B(p_input[7191]), .Z(n8731) );
  XOR U8305 ( .A(n8732), .B(n8733), .Z(n8723) );
  AND U8306 ( .A(n8734), .B(n8735), .Z(n8733) );
  XOR U8307 ( .A(n8732), .B(n7863), .Z(n8735) );
  XNOR U8308 ( .A(p_input[7254]), .B(n8736), .Z(n7863) );
  AND U8309 ( .A(n231), .B(n8737), .Z(n8736) );
  XOR U8310 ( .A(p_input[7286]), .B(p_input[7254]), .Z(n8737) );
  XNOR U8311 ( .A(n7860), .B(n8732), .Z(n8734) );
  XOR U8312 ( .A(n8738), .B(n8739), .Z(n7860) );
  AND U8313 ( .A(n228), .B(n8740), .Z(n8739) );
  XOR U8314 ( .A(p_input[7222]), .B(p_input[7190]), .Z(n8740) );
  XOR U8315 ( .A(n8741), .B(n8742), .Z(n8732) );
  AND U8316 ( .A(n8743), .B(n8744), .Z(n8742) );
  XOR U8317 ( .A(n8741), .B(n7875), .Z(n8744) );
  XNOR U8318 ( .A(p_input[7253]), .B(n8745), .Z(n7875) );
  AND U8319 ( .A(n231), .B(n8746), .Z(n8745) );
  XOR U8320 ( .A(p_input[7285]), .B(p_input[7253]), .Z(n8746) );
  XNOR U8321 ( .A(n7872), .B(n8741), .Z(n8743) );
  XOR U8322 ( .A(n8747), .B(n8748), .Z(n7872) );
  AND U8323 ( .A(n228), .B(n8749), .Z(n8748) );
  XOR U8324 ( .A(p_input[7221]), .B(p_input[7189]), .Z(n8749) );
  XOR U8325 ( .A(n8750), .B(n8751), .Z(n8741) );
  AND U8326 ( .A(n8752), .B(n8753), .Z(n8751) );
  XOR U8327 ( .A(n8750), .B(n7887), .Z(n8753) );
  XNOR U8328 ( .A(p_input[7252]), .B(n8754), .Z(n7887) );
  AND U8329 ( .A(n231), .B(n8755), .Z(n8754) );
  XOR U8330 ( .A(p_input[7284]), .B(p_input[7252]), .Z(n8755) );
  XNOR U8331 ( .A(n7884), .B(n8750), .Z(n8752) );
  XOR U8332 ( .A(n8756), .B(n8757), .Z(n7884) );
  AND U8333 ( .A(n228), .B(n8758), .Z(n8757) );
  XOR U8334 ( .A(p_input[7220]), .B(p_input[7188]), .Z(n8758) );
  XOR U8335 ( .A(n8759), .B(n8760), .Z(n8750) );
  AND U8336 ( .A(n8761), .B(n8762), .Z(n8760) );
  XOR U8337 ( .A(n8759), .B(n7899), .Z(n8762) );
  XNOR U8338 ( .A(p_input[7251]), .B(n8763), .Z(n7899) );
  AND U8339 ( .A(n231), .B(n8764), .Z(n8763) );
  XOR U8340 ( .A(p_input[7283]), .B(p_input[7251]), .Z(n8764) );
  XNOR U8341 ( .A(n7896), .B(n8759), .Z(n8761) );
  XOR U8342 ( .A(n8765), .B(n8766), .Z(n7896) );
  AND U8343 ( .A(n228), .B(n8767), .Z(n8766) );
  XOR U8344 ( .A(p_input[7219]), .B(p_input[7187]), .Z(n8767) );
  XOR U8345 ( .A(n8768), .B(n8769), .Z(n8759) );
  AND U8346 ( .A(n8770), .B(n8771), .Z(n8769) );
  XOR U8347 ( .A(n8768), .B(n7911), .Z(n8771) );
  XNOR U8348 ( .A(p_input[7250]), .B(n8772), .Z(n7911) );
  AND U8349 ( .A(n231), .B(n8773), .Z(n8772) );
  XOR U8350 ( .A(p_input[7282]), .B(p_input[7250]), .Z(n8773) );
  XNOR U8351 ( .A(n7908), .B(n8768), .Z(n8770) );
  XOR U8352 ( .A(n8774), .B(n8775), .Z(n7908) );
  AND U8353 ( .A(n228), .B(n8776), .Z(n8775) );
  XOR U8354 ( .A(p_input[7218]), .B(p_input[7186]), .Z(n8776) );
  XOR U8355 ( .A(n8777), .B(n8778), .Z(n8768) );
  AND U8356 ( .A(n8779), .B(n8780), .Z(n8778) );
  XOR U8357 ( .A(n8777), .B(n7923), .Z(n8780) );
  XNOR U8358 ( .A(p_input[7249]), .B(n8781), .Z(n7923) );
  AND U8359 ( .A(n231), .B(n8782), .Z(n8781) );
  XOR U8360 ( .A(p_input[7281]), .B(p_input[7249]), .Z(n8782) );
  XNOR U8361 ( .A(n7920), .B(n8777), .Z(n8779) );
  XOR U8362 ( .A(n8783), .B(n8784), .Z(n7920) );
  AND U8363 ( .A(n228), .B(n8785), .Z(n8784) );
  XOR U8364 ( .A(p_input[7217]), .B(p_input[7185]), .Z(n8785) );
  XOR U8365 ( .A(n8786), .B(n8787), .Z(n8777) );
  AND U8366 ( .A(n8788), .B(n8789), .Z(n8787) );
  XOR U8367 ( .A(n8786), .B(n7935), .Z(n8789) );
  XNOR U8368 ( .A(p_input[7248]), .B(n8790), .Z(n7935) );
  AND U8369 ( .A(n231), .B(n8791), .Z(n8790) );
  XOR U8370 ( .A(p_input[7280]), .B(p_input[7248]), .Z(n8791) );
  XNOR U8371 ( .A(n7932), .B(n8786), .Z(n8788) );
  XOR U8372 ( .A(n8792), .B(n8793), .Z(n7932) );
  AND U8373 ( .A(n228), .B(n8794), .Z(n8793) );
  XOR U8374 ( .A(p_input[7216]), .B(p_input[7184]), .Z(n8794) );
  XOR U8375 ( .A(n8795), .B(n8796), .Z(n8786) );
  AND U8376 ( .A(n8797), .B(n8798), .Z(n8796) );
  XOR U8377 ( .A(n8795), .B(n7947), .Z(n8798) );
  XNOR U8378 ( .A(p_input[7247]), .B(n8799), .Z(n7947) );
  AND U8379 ( .A(n231), .B(n8800), .Z(n8799) );
  XOR U8380 ( .A(p_input[7279]), .B(p_input[7247]), .Z(n8800) );
  XNOR U8381 ( .A(n7944), .B(n8795), .Z(n8797) );
  XOR U8382 ( .A(n8801), .B(n8802), .Z(n7944) );
  AND U8383 ( .A(n228), .B(n8803), .Z(n8802) );
  XOR U8384 ( .A(p_input[7215]), .B(p_input[7183]), .Z(n8803) );
  XOR U8385 ( .A(n8804), .B(n8805), .Z(n8795) );
  AND U8386 ( .A(n8806), .B(n8807), .Z(n8805) );
  XOR U8387 ( .A(n8804), .B(n7959), .Z(n8807) );
  XNOR U8388 ( .A(p_input[7246]), .B(n8808), .Z(n7959) );
  AND U8389 ( .A(n231), .B(n8809), .Z(n8808) );
  XOR U8390 ( .A(p_input[7278]), .B(p_input[7246]), .Z(n8809) );
  XNOR U8391 ( .A(n7956), .B(n8804), .Z(n8806) );
  XOR U8392 ( .A(n8810), .B(n8811), .Z(n7956) );
  AND U8393 ( .A(n228), .B(n8812), .Z(n8811) );
  XOR U8394 ( .A(p_input[7214]), .B(p_input[7182]), .Z(n8812) );
  XOR U8395 ( .A(n8813), .B(n8814), .Z(n8804) );
  AND U8396 ( .A(n8815), .B(n8816), .Z(n8814) );
  XOR U8397 ( .A(n8813), .B(n7971), .Z(n8816) );
  XNOR U8398 ( .A(p_input[7245]), .B(n8817), .Z(n7971) );
  AND U8399 ( .A(n231), .B(n8818), .Z(n8817) );
  XOR U8400 ( .A(p_input[7277]), .B(p_input[7245]), .Z(n8818) );
  XNOR U8401 ( .A(n7968), .B(n8813), .Z(n8815) );
  XOR U8402 ( .A(n8819), .B(n8820), .Z(n7968) );
  AND U8403 ( .A(n228), .B(n8821), .Z(n8820) );
  XOR U8404 ( .A(p_input[7213]), .B(p_input[7181]), .Z(n8821) );
  XOR U8405 ( .A(n8822), .B(n8823), .Z(n8813) );
  AND U8406 ( .A(n8824), .B(n8825), .Z(n8823) );
  XOR U8407 ( .A(n8822), .B(n7983), .Z(n8825) );
  XNOR U8408 ( .A(p_input[7244]), .B(n8826), .Z(n7983) );
  AND U8409 ( .A(n231), .B(n8827), .Z(n8826) );
  XOR U8410 ( .A(p_input[7276]), .B(p_input[7244]), .Z(n8827) );
  XNOR U8411 ( .A(n7980), .B(n8822), .Z(n8824) );
  XOR U8412 ( .A(n8828), .B(n8829), .Z(n7980) );
  AND U8413 ( .A(n228), .B(n8830), .Z(n8829) );
  XOR U8414 ( .A(p_input[7212]), .B(p_input[7180]), .Z(n8830) );
  XOR U8415 ( .A(n8831), .B(n8832), .Z(n8822) );
  AND U8416 ( .A(n8833), .B(n8834), .Z(n8832) );
  XOR U8417 ( .A(n8831), .B(n7995), .Z(n8834) );
  XNOR U8418 ( .A(p_input[7243]), .B(n8835), .Z(n7995) );
  AND U8419 ( .A(n231), .B(n8836), .Z(n8835) );
  XOR U8420 ( .A(p_input[7275]), .B(p_input[7243]), .Z(n8836) );
  XNOR U8421 ( .A(n7992), .B(n8831), .Z(n8833) );
  XOR U8422 ( .A(n8837), .B(n8838), .Z(n7992) );
  AND U8423 ( .A(n228), .B(n8839), .Z(n8838) );
  XOR U8424 ( .A(p_input[7211]), .B(p_input[7179]), .Z(n8839) );
  XOR U8425 ( .A(n8840), .B(n8841), .Z(n8831) );
  AND U8426 ( .A(n8842), .B(n8843), .Z(n8841) );
  XOR U8427 ( .A(n8840), .B(n8007), .Z(n8843) );
  XNOR U8428 ( .A(p_input[7242]), .B(n8844), .Z(n8007) );
  AND U8429 ( .A(n231), .B(n8845), .Z(n8844) );
  XOR U8430 ( .A(p_input[7274]), .B(p_input[7242]), .Z(n8845) );
  XNOR U8431 ( .A(n8004), .B(n8840), .Z(n8842) );
  XOR U8432 ( .A(n8846), .B(n8847), .Z(n8004) );
  AND U8433 ( .A(n228), .B(n8848), .Z(n8847) );
  XOR U8434 ( .A(p_input[7210]), .B(p_input[7178]), .Z(n8848) );
  XOR U8435 ( .A(n8849), .B(n8850), .Z(n8840) );
  AND U8436 ( .A(n8851), .B(n8852), .Z(n8850) );
  XOR U8437 ( .A(n8849), .B(n8019), .Z(n8852) );
  XNOR U8438 ( .A(p_input[7241]), .B(n8853), .Z(n8019) );
  AND U8439 ( .A(n231), .B(n8854), .Z(n8853) );
  XOR U8440 ( .A(p_input[7273]), .B(p_input[7241]), .Z(n8854) );
  XNOR U8441 ( .A(n8016), .B(n8849), .Z(n8851) );
  XOR U8442 ( .A(n8855), .B(n8856), .Z(n8016) );
  AND U8443 ( .A(n228), .B(n8857), .Z(n8856) );
  XOR U8444 ( .A(p_input[7209]), .B(p_input[7177]), .Z(n8857) );
  XOR U8445 ( .A(n8858), .B(n8859), .Z(n8849) );
  AND U8446 ( .A(n8860), .B(n8861), .Z(n8859) );
  XOR U8447 ( .A(n8858), .B(n8031), .Z(n8861) );
  XNOR U8448 ( .A(p_input[7240]), .B(n8862), .Z(n8031) );
  AND U8449 ( .A(n231), .B(n8863), .Z(n8862) );
  XOR U8450 ( .A(p_input[7272]), .B(p_input[7240]), .Z(n8863) );
  XNOR U8451 ( .A(n8028), .B(n8858), .Z(n8860) );
  XOR U8452 ( .A(n8864), .B(n8865), .Z(n8028) );
  AND U8453 ( .A(n228), .B(n8866), .Z(n8865) );
  XOR U8454 ( .A(p_input[7208]), .B(p_input[7176]), .Z(n8866) );
  XOR U8455 ( .A(n8867), .B(n8868), .Z(n8858) );
  AND U8456 ( .A(n8869), .B(n8870), .Z(n8868) );
  XOR U8457 ( .A(n8867), .B(n8043), .Z(n8870) );
  XNOR U8458 ( .A(p_input[7239]), .B(n8871), .Z(n8043) );
  AND U8459 ( .A(n231), .B(n8872), .Z(n8871) );
  XOR U8460 ( .A(p_input[7271]), .B(p_input[7239]), .Z(n8872) );
  XNOR U8461 ( .A(n8040), .B(n8867), .Z(n8869) );
  XOR U8462 ( .A(n8873), .B(n8874), .Z(n8040) );
  AND U8463 ( .A(n228), .B(n8875), .Z(n8874) );
  XOR U8464 ( .A(p_input[7207]), .B(p_input[7175]), .Z(n8875) );
  XOR U8465 ( .A(n8876), .B(n8877), .Z(n8867) );
  AND U8466 ( .A(n8878), .B(n8879), .Z(n8877) );
  XOR U8467 ( .A(n8876), .B(n8055), .Z(n8879) );
  XNOR U8468 ( .A(p_input[7238]), .B(n8880), .Z(n8055) );
  AND U8469 ( .A(n231), .B(n8881), .Z(n8880) );
  XOR U8470 ( .A(p_input[7270]), .B(p_input[7238]), .Z(n8881) );
  XNOR U8471 ( .A(n8052), .B(n8876), .Z(n8878) );
  XOR U8472 ( .A(n8882), .B(n8883), .Z(n8052) );
  AND U8473 ( .A(n228), .B(n8884), .Z(n8883) );
  XOR U8474 ( .A(p_input[7206]), .B(p_input[7174]), .Z(n8884) );
  XOR U8475 ( .A(n8885), .B(n8886), .Z(n8876) );
  AND U8476 ( .A(n8887), .B(n8888), .Z(n8886) );
  XOR U8477 ( .A(n8885), .B(n8067), .Z(n8888) );
  XNOR U8478 ( .A(p_input[7237]), .B(n8889), .Z(n8067) );
  AND U8479 ( .A(n231), .B(n8890), .Z(n8889) );
  XOR U8480 ( .A(p_input[7269]), .B(p_input[7237]), .Z(n8890) );
  XNOR U8481 ( .A(n8064), .B(n8885), .Z(n8887) );
  XOR U8482 ( .A(n8891), .B(n8892), .Z(n8064) );
  AND U8483 ( .A(n228), .B(n8893), .Z(n8892) );
  XOR U8484 ( .A(p_input[7205]), .B(p_input[7173]), .Z(n8893) );
  XOR U8485 ( .A(n8894), .B(n8895), .Z(n8885) );
  AND U8486 ( .A(n8896), .B(n8897), .Z(n8895) );
  XOR U8487 ( .A(n8894), .B(n8079), .Z(n8897) );
  XNOR U8488 ( .A(p_input[7236]), .B(n8898), .Z(n8079) );
  AND U8489 ( .A(n231), .B(n8899), .Z(n8898) );
  XOR U8490 ( .A(p_input[7268]), .B(p_input[7236]), .Z(n8899) );
  XNOR U8491 ( .A(n8076), .B(n8894), .Z(n8896) );
  XOR U8492 ( .A(n8900), .B(n8901), .Z(n8076) );
  AND U8493 ( .A(n228), .B(n8902), .Z(n8901) );
  XOR U8494 ( .A(p_input[7204]), .B(p_input[7172]), .Z(n8902) );
  XOR U8495 ( .A(n8903), .B(n8904), .Z(n8894) );
  AND U8496 ( .A(n8905), .B(n8906), .Z(n8904) );
  XOR U8497 ( .A(n8903), .B(n8091), .Z(n8906) );
  XNOR U8498 ( .A(p_input[7235]), .B(n8907), .Z(n8091) );
  AND U8499 ( .A(n231), .B(n8908), .Z(n8907) );
  XOR U8500 ( .A(p_input[7267]), .B(p_input[7235]), .Z(n8908) );
  XNOR U8501 ( .A(n8088), .B(n8903), .Z(n8905) );
  XOR U8502 ( .A(n8909), .B(n8910), .Z(n8088) );
  AND U8503 ( .A(n228), .B(n8911), .Z(n8910) );
  XOR U8504 ( .A(p_input[7203]), .B(p_input[7171]), .Z(n8911) );
  XOR U8505 ( .A(n8912), .B(n8913), .Z(n8903) );
  AND U8506 ( .A(n8914), .B(n8915), .Z(n8913) );
  XOR U8507 ( .A(n8912), .B(n8103), .Z(n8915) );
  XNOR U8508 ( .A(p_input[7234]), .B(n8916), .Z(n8103) );
  AND U8509 ( .A(n231), .B(n8917), .Z(n8916) );
  XOR U8510 ( .A(p_input[7266]), .B(p_input[7234]), .Z(n8917) );
  XNOR U8511 ( .A(n8100), .B(n8912), .Z(n8914) );
  XOR U8512 ( .A(n8918), .B(n8919), .Z(n8100) );
  AND U8513 ( .A(n228), .B(n8920), .Z(n8919) );
  XOR U8514 ( .A(p_input[7202]), .B(p_input[7170]), .Z(n8920) );
  XOR U8515 ( .A(n8921), .B(n8922), .Z(n8912) );
  AND U8516 ( .A(n8923), .B(n8924), .Z(n8922) );
  XNOR U8517 ( .A(n8925), .B(n8116), .Z(n8924) );
  XNOR U8518 ( .A(p_input[7233]), .B(n8926), .Z(n8116) );
  AND U8519 ( .A(n231), .B(n8927), .Z(n8926) );
  XNOR U8520 ( .A(p_input[7265]), .B(n8928), .Z(n8927) );
  IV U8521 ( .A(p_input[7233]), .Z(n8928) );
  XNOR U8522 ( .A(n8113), .B(n8921), .Z(n8923) );
  XNOR U8523 ( .A(p_input[7169]), .B(n8929), .Z(n8113) );
  AND U8524 ( .A(n228), .B(n8930), .Z(n8929) );
  XOR U8525 ( .A(p_input[7201]), .B(p_input[7169]), .Z(n8930) );
  IV U8526 ( .A(n8925), .Z(n8921) );
  AND U8527 ( .A(n8651), .B(n8654), .Z(n8925) );
  XOR U8528 ( .A(p_input[7232]), .B(n8931), .Z(n8654) );
  AND U8529 ( .A(n231), .B(n8932), .Z(n8931) );
  XOR U8530 ( .A(p_input[7264]), .B(p_input[7232]), .Z(n8932) );
  XOR U8531 ( .A(n8933), .B(n8934), .Z(n231) );
  AND U8532 ( .A(n8935), .B(n8936), .Z(n8934) );
  XNOR U8533 ( .A(p_input[7295]), .B(n8933), .Z(n8936) );
  XOR U8534 ( .A(n8933), .B(p_input[7263]), .Z(n8935) );
  XOR U8535 ( .A(n8937), .B(n8938), .Z(n8933) );
  AND U8536 ( .A(n8939), .B(n8940), .Z(n8938) );
  XNOR U8537 ( .A(p_input[7294]), .B(n8937), .Z(n8940) );
  XOR U8538 ( .A(n8937), .B(p_input[7262]), .Z(n8939) );
  XOR U8539 ( .A(n8941), .B(n8942), .Z(n8937) );
  AND U8540 ( .A(n8943), .B(n8944), .Z(n8942) );
  XNOR U8541 ( .A(p_input[7293]), .B(n8941), .Z(n8944) );
  XOR U8542 ( .A(n8941), .B(p_input[7261]), .Z(n8943) );
  XOR U8543 ( .A(n8945), .B(n8946), .Z(n8941) );
  AND U8544 ( .A(n8947), .B(n8948), .Z(n8946) );
  XNOR U8545 ( .A(p_input[7292]), .B(n8945), .Z(n8948) );
  XOR U8546 ( .A(n8945), .B(p_input[7260]), .Z(n8947) );
  XOR U8547 ( .A(n8949), .B(n8950), .Z(n8945) );
  AND U8548 ( .A(n8951), .B(n8952), .Z(n8950) );
  XNOR U8549 ( .A(p_input[7291]), .B(n8949), .Z(n8952) );
  XOR U8550 ( .A(n8949), .B(p_input[7259]), .Z(n8951) );
  XOR U8551 ( .A(n8953), .B(n8954), .Z(n8949) );
  AND U8552 ( .A(n8955), .B(n8956), .Z(n8954) );
  XNOR U8553 ( .A(p_input[7290]), .B(n8953), .Z(n8956) );
  XOR U8554 ( .A(n8953), .B(p_input[7258]), .Z(n8955) );
  XOR U8555 ( .A(n8957), .B(n8958), .Z(n8953) );
  AND U8556 ( .A(n8959), .B(n8960), .Z(n8958) );
  XNOR U8557 ( .A(p_input[7289]), .B(n8957), .Z(n8960) );
  XOR U8558 ( .A(n8957), .B(p_input[7257]), .Z(n8959) );
  XOR U8559 ( .A(n8961), .B(n8962), .Z(n8957) );
  AND U8560 ( .A(n8963), .B(n8964), .Z(n8962) );
  XNOR U8561 ( .A(p_input[7288]), .B(n8961), .Z(n8964) );
  XOR U8562 ( .A(n8961), .B(p_input[7256]), .Z(n8963) );
  XOR U8563 ( .A(n8965), .B(n8966), .Z(n8961) );
  AND U8564 ( .A(n8967), .B(n8968), .Z(n8966) );
  XNOR U8565 ( .A(p_input[7287]), .B(n8965), .Z(n8968) );
  XOR U8566 ( .A(n8965), .B(p_input[7255]), .Z(n8967) );
  XOR U8567 ( .A(n8969), .B(n8970), .Z(n8965) );
  AND U8568 ( .A(n8971), .B(n8972), .Z(n8970) );
  XNOR U8569 ( .A(p_input[7286]), .B(n8969), .Z(n8972) );
  XOR U8570 ( .A(n8969), .B(p_input[7254]), .Z(n8971) );
  XOR U8571 ( .A(n8973), .B(n8974), .Z(n8969) );
  AND U8572 ( .A(n8975), .B(n8976), .Z(n8974) );
  XNOR U8573 ( .A(p_input[7285]), .B(n8973), .Z(n8976) );
  XOR U8574 ( .A(n8973), .B(p_input[7253]), .Z(n8975) );
  XOR U8575 ( .A(n8977), .B(n8978), .Z(n8973) );
  AND U8576 ( .A(n8979), .B(n8980), .Z(n8978) );
  XNOR U8577 ( .A(p_input[7284]), .B(n8977), .Z(n8980) );
  XOR U8578 ( .A(n8977), .B(p_input[7252]), .Z(n8979) );
  XOR U8579 ( .A(n8981), .B(n8982), .Z(n8977) );
  AND U8580 ( .A(n8983), .B(n8984), .Z(n8982) );
  XNOR U8581 ( .A(p_input[7283]), .B(n8981), .Z(n8984) );
  XOR U8582 ( .A(n8981), .B(p_input[7251]), .Z(n8983) );
  XOR U8583 ( .A(n8985), .B(n8986), .Z(n8981) );
  AND U8584 ( .A(n8987), .B(n8988), .Z(n8986) );
  XNOR U8585 ( .A(p_input[7282]), .B(n8985), .Z(n8988) );
  XOR U8586 ( .A(n8985), .B(p_input[7250]), .Z(n8987) );
  XOR U8587 ( .A(n8989), .B(n8990), .Z(n8985) );
  AND U8588 ( .A(n8991), .B(n8992), .Z(n8990) );
  XNOR U8589 ( .A(p_input[7281]), .B(n8989), .Z(n8992) );
  XOR U8590 ( .A(n8989), .B(p_input[7249]), .Z(n8991) );
  XOR U8591 ( .A(n8993), .B(n8994), .Z(n8989) );
  AND U8592 ( .A(n8995), .B(n8996), .Z(n8994) );
  XNOR U8593 ( .A(p_input[7280]), .B(n8993), .Z(n8996) );
  XOR U8594 ( .A(n8993), .B(p_input[7248]), .Z(n8995) );
  XOR U8595 ( .A(n8997), .B(n8998), .Z(n8993) );
  AND U8596 ( .A(n8999), .B(n9000), .Z(n8998) );
  XNOR U8597 ( .A(p_input[7279]), .B(n8997), .Z(n9000) );
  XOR U8598 ( .A(n8997), .B(p_input[7247]), .Z(n8999) );
  XOR U8599 ( .A(n9001), .B(n9002), .Z(n8997) );
  AND U8600 ( .A(n9003), .B(n9004), .Z(n9002) );
  XNOR U8601 ( .A(p_input[7278]), .B(n9001), .Z(n9004) );
  XOR U8602 ( .A(n9001), .B(p_input[7246]), .Z(n9003) );
  XOR U8603 ( .A(n9005), .B(n9006), .Z(n9001) );
  AND U8604 ( .A(n9007), .B(n9008), .Z(n9006) );
  XNOR U8605 ( .A(p_input[7277]), .B(n9005), .Z(n9008) );
  XOR U8606 ( .A(n9005), .B(p_input[7245]), .Z(n9007) );
  XOR U8607 ( .A(n9009), .B(n9010), .Z(n9005) );
  AND U8608 ( .A(n9011), .B(n9012), .Z(n9010) );
  XNOR U8609 ( .A(p_input[7276]), .B(n9009), .Z(n9012) );
  XOR U8610 ( .A(n9009), .B(p_input[7244]), .Z(n9011) );
  XOR U8611 ( .A(n9013), .B(n9014), .Z(n9009) );
  AND U8612 ( .A(n9015), .B(n9016), .Z(n9014) );
  XNOR U8613 ( .A(p_input[7275]), .B(n9013), .Z(n9016) );
  XOR U8614 ( .A(n9013), .B(p_input[7243]), .Z(n9015) );
  XOR U8615 ( .A(n9017), .B(n9018), .Z(n9013) );
  AND U8616 ( .A(n9019), .B(n9020), .Z(n9018) );
  XNOR U8617 ( .A(p_input[7274]), .B(n9017), .Z(n9020) );
  XOR U8618 ( .A(n9017), .B(p_input[7242]), .Z(n9019) );
  XOR U8619 ( .A(n9021), .B(n9022), .Z(n9017) );
  AND U8620 ( .A(n9023), .B(n9024), .Z(n9022) );
  XNOR U8621 ( .A(p_input[7273]), .B(n9021), .Z(n9024) );
  XOR U8622 ( .A(n9021), .B(p_input[7241]), .Z(n9023) );
  XOR U8623 ( .A(n9025), .B(n9026), .Z(n9021) );
  AND U8624 ( .A(n9027), .B(n9028), .Z(n9026) );
  XNOR U8625 ( .A(p_input[7272]), .B(n9025), .Z(n9028) );
  XOR U8626 ( .A(n9025), .B(p_input[7240]), .Z(n9027) );
  XOR U8627 ( .A(n9029), .B(n9030), .Z(n9025) );
  AND U8628 ( .A(n9031), .B(n9032), .Z(n9030) );
  XNOR U8629 ( .A(p_input[7271]), .B(n9029), .Z(n9032) );
  XOR U8630 ( .A(n9029), .B(p_input[7239]), .Z(n9031) );
  XOR U8631 ( .A(n9033), .B(n9034), .Z(n9029) );
  AND U8632 ( .A(n9035), .B(n9036), .Z(n9034) );
  XNOR U8633 ( .A(p_input[7270]), .B(n9033), .Z(n9036) );
  XOR U8634 ( .A(n9033), .B(p_input[7238]), .Z(n9035) );
  XOR U8635 ( .A(n9037), .B(n9038), .Z(n9033) );
  AND U8636 ( .A(n9039), .B(n9040), .Z(n9038) );
  XNOR U8637 ( .A(p_input[7269]), .B(n9037), .Z(n9040) );
  XOR U8638 ( .A(n9037), .B(p_input[7237]), .Z(n9039) );
  XOR U8639 ( .A(n9041), .B(n9042), .Z(n9037) );
  AND U8640 ( .A(n9043), .B(n9044), .Z(n9042) );
  XNOR U8641 ( .A(p_input[7268]), .B(n9041), .Z(n9044) );
  XOR U8642 ( .A(n9041), .B(p_input[7236]), .Z(n9043) );
  XOR U8643 ( .A(n9045), .B(n9046), .Z(n9041) );
  AND U8644 ( .A(n9047), .B(n9048), .Z(n9046) );
  XNOR U8645 ( .A(p_input[7267]), .B(n9045), .Z(n9048) );
  XOR U8646 ( .A(n9045), .B(p_input[7235]), .Z(n9047) );
  XOR U8647 ( .A(n9049), .B(n9050), .Z(n9045) );
  AND U8648 ( .A(n9051), .B(n9052), .Z(n9050) );
  XNOR U8649 ( .A(p_input[7266]), .B(n9049), .Z(n9052) );
  XOR U8650 ( .A(n9049), .B(p_input[7234]), .Z(n9051) );
  XNOR U8651 ( .A(n9053), .B(n9054), .Z(n9049) );
  AND U8652 ( .A(n9055), .B(n9056), .Z(n9054) );
  XOR U8653 ( .A(p_input[7265]), .B(n9053), .Z(n9056) );
  XNOR U8654 ( .A(p_input[7233]), .B(n9053), .Z(n9055) );
  AND U8655 ( .A(p_input[7264]), .B(n9057), .Z(n9053) );
  IV U8656 ( .A(p_input[7232]), .Z(n9057) );
  XNOR U8657 ( .A(p_input[7168]), .B(n9058), .Z(n8651) );
  AND U8658 ( .A(n228), .B(n9059), .Z(n9058) );
  XOR U8659 ( .A(p_input[7200]), .B(p_input[7168]), .Z(n9059) );
  XOR U8660 ( .A(n9060), .B(n9061), .Z(n228) );
  AND U8661 ( .A(n9062), .B(n9063), .Z(n9061) );
  XNOR U8662 ( .A(p_input[7231]), .B(n9060), .Z(n9063) );
  XOR U8663 ( .A(n9060), .B(p_input[7199]), .Z(n9062) );
  XOR U8664 ( .A(n9064), .B(n9065), .Z(n9060) );
  AND U8665 ( .A(n9066), .B(n9067), .Z(n9065) );
  XNOR U8666 ( .A(p_input[7230]), .B(n9064), .Z(n9067) );
  XNOR U8667 ( .A(n9064), .B(n8666), .Z(n9066) );
  IV U8668 ( .A(p_input[7198]), .Z(n8666) );
  XOR U8669 ( .A(n9068), .B(n9069), .Z(n9064) );
  AND U8670 ( .A(n9070), .B(n9071), .Z(n9069) );
  XNOR U8671 ( .A(p_input[7229]), .B(n9068), .Z(n9071) );
  XNOR U8672 ( .A(n9068), .B(n8675), .Z(n9070) );
  IV U8673 ( .A(p_input[7197]), .Z(n8675) );
  XOR U8674 ( .A(n9072), .B(n9073), .Z(n9068) );
  AND U8675 ( .A(n9074), .B(n9075), .Z(n9073) );
  XNOR U8676 ( .A(p_input[7228]), .B(n9072), .Z(n9075) );
  XNOR U8677 ( .A(n9072), .B(n8684), .Z(n9074) );
  IV U8678 ( .A(p_input[7196]), .Z(n8684) );
  XOR U8679 ( .A(n9076), .B(n9077), .Z(n9072) );
  AND U8680 ( .A(n9078), .B(n9079), .Z(n9077) );
  XNOR U8681 ( .A(p_input[7227]), .B(n9076), .Z(n9079) );
  XNOR U8682 ( .A(n9076), .B(n8693), .Z(n9078) );
  IV U8683 ( .A(p_input[7195]), .Z(n8693) );
  XOR U8684 ( .A(n9080), .B(n9081), .Z(n9076) );
  AND U8685 ( .A(n9082), .B(n9083), .Z(n9081) );
  XNOR U8686 ( .A(p_input[7226]), .B(n9080), .Z(n9083) );
  XNOR U8687 ( .A(n9080), .B(n8702), .Z(n9082) );
  IV U8688 ( .A(p_input[7194]), .Z(n8702) );
  XOR U8689 ( .A(n9084), .B(n9085), .Z(n9080) );
  AND U8690 ( .A(n9086), .B(n9087), .Z(n9085) );
  XNOR U8691 ( .A(p_input[7225]), .B(n9084), .Z(n9087) );
  XNOR U8692 ( .A(n9084), .B(n8711), .Z(n9086) );
  IV U8693 ( .A(p_input[7193]), .Z(n8711) );
  XOR U8694 ( .A(n9088), .B(n9089), .Z(n9084) );
  AND U8695 ( .A(n9090), .B(n9091), .Z(n9089) );
  XNOR U8696 ( .A(p_input[7224]), .B(n9088), .Z(n9091) );
  XNOR U8697 ( .A(n9088), .B(n8720), .Z(n9090) );
  IV U8698 ( .A(p_input[7192]), .Z(n8720) );
  XOR U8699 ( .A(n9092), .B(n9093), .Z(n9088) );
  AND U8700 ( .A(n9094), .B(n9095), .Z(n9093) );
  XNOR U8701 ( .A(p_input[7223]), .B(n9092), .Z(n9095) );
  XNOR U8702 ( .A(n9092), .B(n8729), .Z(n9094) );
  IV U8703 ( .A(p_input[7191]), .Z(n8729) );
  XOR U8704 ( .A(n9096), .B(n9097), .Z(n9092) );
  AND U8705 ( .A(n9098), .B(n9099), .Z(n9097) );
  XNOR U8706 ( .A(p_input[7222]), .B(n9096), .Z(n9099) );
  XNOR U8707 ( .A(n9096), .B(n8738), .Z(n9098) );
  IV U8708 ( .A(p_input[7190]), .Z(n8738) );
  XOR U8709 ( .A(n9100), .B(n9101), .Z(n9096) );
  AND U8710 ( .A(n9102), .B(n9103), .Z(n9101) );
  XNOR U8711 ( .A(p_input[7221]), .B(n9100), .Z(n9103) );
  XNOR U8712 ( .A(n9100), .B(n8747), .Z(n9102) );
  IV U8713 ( .A(p_input[7189]), .Z(n8747) );
  XOR U8714 ( .A(n9104), .B(n9105), .Z(n9100) );
  AND U8715 ( .A(n9106), .B(n9107), .Z(n9105) );
  XNOR U8716 ( .A(p_input[7220]), .B(n9104), .Z(n9107) );
  XNOR U8717 ( .A(n9104), .B(n8756), .Z(n9106) );
  IV U8718 ( .A(p_input[7188]), .Z(n8756) );
  XOR U8719 ( .A(n9108), .B(n9109), .Z(n9104) );
  AND U8720 ( .A(n9110), .B(n9111), .Z(n9109) );
  XNOR U8721 ( .A(p_input[7219]), .B(n9108), .Z(n9111) );
  XNOR U8722 ( .A(n9108), .B(n8765), .Z(n9110) );
  IV U8723 ( .A(p_input[7187]), .Z(n8765) );
  XOR U8724 ( .A(n9112), .B(n9113), .Z(n9108) );
  AND U8725 ( .A(n9114), .B(n9115), .Z(n9113) );
  XNOR U8726 ( .A(p_input[7218]), .B(n9112), .Z(n9115) );
  XNOR U8727 ( .A(n9112), .B(n8774), .Z(n9114) );
  IV U8728 ( .A(p_input[7186]), .Z(n8774) );
  XOR U8729 ( .A(n9116), .B(n9117), .Z(n9112) );
  AND U8730 ( .A(n9118), .B(n9119), .Z(n9117) );
  XNOR U8731 ( .A(p_input[7217]), .B(n9116), .Z(n9119) );
  XNOR U8732 ( .A(n9116), .B(n8783), .Z(n9118) );
  IV U8733 ( .A(p_input[7185]), .Z(n8783) );
  XOR U8734 ( .A(n9120), .B(n9121), .Z(n9116) );
  AND U8735 ( .A(n9122), .B(n9123), .Z(n9121) );
  XNOR U8736 ( .A(p_input[7216]), .B(n9120), .Z(n9123) );
  XNOR U8737 ( .A(n9120), .B(n8792), .Z(n9122) );
  IV U8738 ( .A(p_input[7184]), .Z(n8792) );
  XOR U8739 ( .A(n9124), .B(n9125), .Z(n9120) );
  AND U8740 ( .A(n9126), .B(n9127), .Z(n9125) );
  XNOR U8741 ( .A(p_input[7215]), .B(n9124), .Z(n9127) );
  XNOR U8742 ( .A(n9124), .B(n8801), .Z(n9126) );
  IV U8743 ( .A(p_input[7183]), .Z(n8801) );
  XOR U8744 ( .A(n9128), .B(n9129), .Z(n9124) );
  AND U8745 ( .A(n9130), .B(n9131), .Z(n9129) );
  XNOR U8746 ( .A(p_input[7214]), .B(n9128), .Z(n9131) );
  XNOR U8747 ( .A(n9128), .B(n8810), .Z(n9130) );
  IV U8748 ( .A(p_input[7182]), .Z(n8810) );
  XOR U8749 ( .A(n9132), .B(n9133), .Z(n9128) );
  AND U8750 ( .A(n9134), .B(n9135), .Z(n9133) );
  XNOR U8751 ( .A(p_input[7213]), .B(n9132), .Z(n9135) );
  XNOR U8752 ( .A(n9132), .B(n8819), .Z(n9134) );
  IV U8753 ( .A(p_input[7181]), .Z(n8819) );
  XOR U8754 ( .A(n9136), .B(n9137), .Z(n9132) );
  AND U8755 ( .A(n9138), .B(n9139), .Z(n9137) );
  XNOR U8756 ( .A(p_input[7212]), .B(n9136), .Z(n9139) );
  XNOR U8757 ( .A(n9136), .B(n8828), .Z(n9138) );
  IV U8758 ( .A(p_input[7180]), .Z(n8828) );
  XOR U8759 ( .A(n9140), .B(n9141), .Z(n9136) );
  AND U8760 ( .A(n9142), .B(n9143), .Z(n9141) );
  XNOR U8761 ( .A(p_input[7211]), .B(n9140), .Z(n9143) );
  XNOR U8762 ( .A(n9140), .B(n8837), .Z(n9142) );
  IV U8763 ( .A(p_input[7179]), .Z(n8837) );
  XOR U8764 ( .A(n9144), .B(n9145), .Z(n9140) );
  AND U8765 ( .A(n9146), .B(n9147), .Z(n9145) );
  XNOR U8766 ( .A(p_input[7210]), .B(n9144), .Z(n9147) );
  XNOR U8767 ( .A(n9144), .B(n8846), .Z(n9146) );
  IV U8768 ( .A(p_input[7178]), .Z(n8846) );
  XOR U8769 ( .A(n9148), .B(n9149), .Z(n9144) );
  AND U8770 ( .A(n9150), .B(n9151), .Z(n9149) );
  XNOR U8771 ( .A(p_input[7209]), .B(n9148), .Z(n9151) );
  XNOR U8772 ( .A(n9148), .B(n8855), .Z(n9150) );
  IV U8773 ( .A(p_input[7177]), .Z(n8855) );
  XOR U8774 ( .A(n9152), .B(n9153), .Z(n9148) );
  AND U8775 ( .A(n9154), .B(n9155), .Z(n9153) );
  XNOR U8776 ( .A(p_input[7208]), .B(n9152), .Z(n9155) );
  XNOR U8777 ( .A(n9152), .B(n8864), .Z(n9154) );
  IV U8778 ( .A(p_input[7176]), .Z(n8864) );
  XOR U8779 ( .A(n9156), .B(n9157), .Z(n9152) );
  AND U8780 ( .A(n9158), .B(n9159), .Z(n9157) );
  XNOR U8781 ( .A(p_input[7207]), .B(n9156), .Z(n9159) );
  XNOR U8782 ( .A(n9156), .B(n8873), .Z(n9158) );
  IV U8783 ( .A(p_input[7175]), .Z(n8873) );
  XOR U8784 ( .A(n9160), .B(n9161), .Z(n9156) );
  AND U8785 ( .A(n9162), .B(n9163), .Z(n9161) );
  XNOR U8786 ( .A(p_input[7206]), .B(n9160), .Z(n9163) );
  XNOR U8787 ( .A(n9160), .B(n8882), .Z(n9162) );
  IV U8788 ( .A(p_input[7174]), .Z(n8882) );
  XOR U8789 ( .A(n9164), .B(n9165), .Z(n9160) );
  AND U8790 ( .A(n9166), .B(n9167), .Z(n9165) );
  XNOR U8791 ( .A(p_input[7205]), .B(n9164), .Z(n9167) );
  XNOR U8792 ( .A(n9164), .B(n8891), .Z(n9166) );
  IV U8793 ( .A(p_input[7173]), .Z(n8891) );
  XOR U8794 ( .A(n9168), .B(n9169), .Z(n9164) );
  AND U8795 ( .A(n9170), .B(n9171), .Z(n9169) );
  XNOR U8796 ( .A(p_input[7204]), .B(n9168), .Z(n9171) );
  XNOR U8797 ( .A(n9168), .B(n8900), .Z(n9170) );
  IV U8798 ( .A(p_input[7172]), .Z(n8900) );
  XOR U8799 ( .A(n9172), .B(n9173), .Z(n9168) );
  AND U8800 ( .A(n9174), .B(n9175), .Z(n9173) );
  XNOR U8801 ( .A(p_input[7203]), .B(n9172), .Z(n9175) );
  XNOR U8802 ( .A(n9172), .B(n8909), .Z(n9174) );
  IV U8803 ( .A(p_input[7171]), .Z(n8909) );
  XOR U8804 ( .A(n9176), .B(n9177), .Z(n9172) );
  AND U8805 ( .A(n9178), .B(n9179), .Z(n9177) );
  XNOR U8806 ( .A(p_input[7202]), .B(n9176), .Z(n9179) );
  XNOR U8807 ( .A(n9176), .B(n8918), .Z(n9178) );
  IV U8808 ( .A(p_input[7170]), .Z(n8918) );
  XNOR U8809 ( .A(n9180), .B(n9181), .Z(n9176) );
  AND U8810 ( .A(n9182), .B(n9183), .Z(n9181) );
  XOR U8811 ( .A(p_input[7201]), .B(n9180), .Z(n9183) );
  XNOR U8812 ( .A(p_input[7169]), .B(n9180), .Z(n9182) );
  AND U8813 ( .A(p_input[7200]), .B(n9184), .Z(n9180) );
  IV U8814 ( .A(p_input[7168]), .Z(n9184) );
  XOR U8815 ( .A(n9185), .B(n9186), .Z(n1897) );
  AND U8816 ( .A(n1085), .B(n9187), .Z(n9186) );
  XNOR U8817 ( .A(n9188), .B(n9185), .Z(n9187) );
  XOR U8818 ( .A(n9189), .B(n9190), .Z(n1085) );
  AND U8819 ( .A(n9191), .B(n9192), .Z(n9190) );
  XOR U8820 ( .A(n9189), .B(n1912), .Z(n9192) );
  XOR U8821 ( .A(n9193), .B(n9194), .Z(n1912) );
  AND U8822 ( .A(n1003), .B(n9195), .Z(n9194) );
  XOR U8823 ( .A(n9196), .B(n9193), .Z(n9195) );
  XNOR U8824 ( .A(n1909), .B(n9189), .Z(n9191) );
  XOR U8825 ( .A(n9197), .B(n9198), .Z(n1909) );
  AND U8826 ( .A(n1000), .B(n9199), .Z(n9198) );
  XOR U8827 ( .A(n9200), .B(n9197), .Z(n9199) );
  XOR U8828 ( .A(n9201), .B(n9202), .Z(n9189) );
  AND U8829 ( .A(n9203), .B(n9204), .Z(n9202) );
  XOR U8830 ( .A(n9201), .B(n1924), .Z(n9204) );
  XOR U8831 ( .A(n9205), .B(n9206), .Z(n1924) );
  AND U8832 ( .A(n1003), .B(n9207), .Z(n9206) );
  XOR U8833 ( .A(n9208), .B(n9205), .Z(n9207) );
  XNOR U8834 ( .A(n1921), .B(n9201), .Z(n9203) );
  XOR U8835 ( .A(n9209), .B(n9210), .Z(n1921) );
  AND U8836 ( .A(n1000), .B(n9211), .Z(n9210) );
  XOR U8837 ( .A(n9212), .B(n9209), .Z(n9211) );
  XOR U8838 ( .A(n9213), .B(n9214), .Z(n9201) );
  AND U8839 ( .A(n9215), .B(n9216), .Z(n9214) );
  XOR U8840 ( .A(n9213), .B(n1936), .Z(n9216) );
  XOR U8841 ( .A(n9217), .B(n9218), .Z(n1936) );
  AND U8842 ( .A(n1003), .B(n9219), .Z(n9218) );
  XOR U8843 ( .A(n9220), .B(n9217), .Z(n9219) );
  XNOR U8844 ( .A(n1933), .B(n9213), .Z(n9215) );
  XOR U8845 ( .A(n9221), .B(n9222), .Z(n1933) );
  AND U8846 ( .A(n1000), .B(n9223), .Z(n9222) );
  XOR U8847 ( .A(n9224), .B(n9221), .Z(n9223) );
  XOR U8848 ( .A(n9225), .B(n9226), .Z(n9213) );
  AND U8849 ( .A(n9227), .B(n9228), .Z(n9226) );
  XOR U8850 ( .A(n9225), .B(n1948), .Z(n9228) );
  XOR U8851 ( .A(n9229), .B(n9230), .Z(n1948) );
  AND U8852 ( .A(n1003), .B(n9231), .Z(n9230) );
  XOR U8853 ( .A(n9232), .B(n9229), .Z(n9231) );
  XNOR U8854 ( .A(n1945), .B(n9225), .Z(n9227) );
  XOR U8855 ( .A(n9233), .B(n9234), .Z(n1945) );
  AND U8856 ( .A(n1000), .B(n9235), .Z(n9234) );
  XOR U8857 ( .A(n9236), .B(n9233), .Z(n9235) );
  XOR U8858 ( .A(n9237), .B(n9238), .Z(n9225) );
  AND U8859 ( .A(n9239), .B(n9240), .Z(n9238) );
  XOR U8860 ( .A(n9237), .B(n1960), .Z(n9240) );
  XOR U8861 ( .A(n9241), .B(n9242), .Z(n1960) );
  AND U8862 ( .A(n1003), .B(n9243), .Z(n9242) );
  XOR U8863 ( .A(n9244), .B(n9241), .Z(n9243) );
  XNOR U8864 ( .A(n1957), .B(n9237), .Z(n9239) );
  XOR U8865 ( .A(n9245), .B(n9246), .Z(n1957) );
  AND U8866 ( .A(n1000), .B(n9247), .Z(n9246) );
  XOR U8867 ( .A(n9248), .B(n9245), .Z(n9247) );
  XOR U8868 ( .A(n9249), .B(n9250), .Z(n9237) );
  AND U8869 ( .A(n9251), .B(n9252), .Z(n9250) );
  XOR U8870 ( .A(n9249), .B(n1972), .Z(n9252) );
  XOR U8871 ( .A(n9253), .B(n9254), .Z(n1972) );
  AND U8872 ( .A(n1003), .B(n9255), .Z(n9254) );
  XOR U8873 ( .A(n9256), .B(n9253), .Z(n9255) );
  XNOR U8874 ( .A(n1969), .B(n9249), .Z(n9251) );
  XOR U8875 ( .A(n9257), .B(n9258), .Z(n1969) );
  AND U8876 ( .A(n1000), .B(n9259), .Z(n9258) );
  XOR U8877 ( .A(n9260), .B(n9257), .Z(n9259) );
  XOR U8878 ( .A(n9261), .B(n9262), .Z(n9249) );
  AND U8879 ( .A(n9263), .B(n9264), .Z(n9262) );
  XOR U8880 ( .A(n9261), .B(n1984), .Z(n9264) );
  XOR U8881 ( .A(n9265), .B(n9266), .Z(n1984) );
  AND U8882 ( .A(n1003), .B(n9267), .Z(n9266) );
  XOR U8883 ( .A(n9268), .B(n9265), .Z(n9267) );
  XNOR U8884 ( .A(n1981), .B(n9261), .Z(n9263) );
  XOR U8885 ( .A(n9269), .B(n9270), .Z(n1981) );
  AND U8886 ( .A(n1000), .B(n9271), .Z(n9270) );
  XOR U8887 ( .A(n9272), .B(n9269), .Z(n9271) );
  XOR U8888 ( .A(n9273), .B(n9274), .Z(n9261) );
  AND U8889 ( .A(n9275), .B(n9276), .Z(n9274) );
  XOR U8890 ( .A(n9273), .B(n1996), .Z(n9276) );
  XOR U8891 ( .A(n9277), .B(n9278), .Z(n1996) );
  AND U8892 ( .A(n1003), .B(n9279), .Z(n9278) );
  XOR U8893 ( .A(n9280), .B(n9277), .Z(n9279) );
  XNOR U8894 ( .A(n1993), .B(n9273), .Z(n9275) );
  XOR U8895 ( .A(n9281), .B(n9282), .Z(n1993) );
  AND U8896 ( .A(n1000), .B(n9283), .Z(n9282) );
  XOR U8897 ( .A(n9284), .B(n9281), .Z(n9283) );
  XOR U8898 ( .A(n9285), .B(n9286), .Z(n9273) );
  AND U8899 ( .A(n9287), .B(n9288), .Z(n9286) );
  XOR U8900 ( .A(n9285), .B(n2008), .Z(n9288) );
  XOR U8901 ( .A(n9289), .B(n9290), .Z(n2008) );
  AND U8902 ( .A(n1003), .B(n9291), .Z(n9290) );
  XOR U8903 ( .A(n9292), .B(n9289), .Z(n9291) );
  XNOR U8904 ( .A(n2005), .B(n9285), .Z(n9287) );
  XOR U8905 ( .A(n9293), .B(n9294), .Z(n2005) );
  AND U8906 ( .A(n1000), .B(n9295), .Z(n9294) );
  XOR U8907 ( .A(n9296), .B(n9293), .Z(n9295) );
  XOR U8908 ( .A(n9297), .B(n9298), .Z(n9285) );
  AND U8909 ( .A(n9299), .B(n9300), .Z(n9298) );
  XOR U8910 ( .A(n9297), .B(n2020), .Z(n9300) );
  XOR U8911 ( .A(n9301), .B(n9302), .Z(n2020) );
  AND U8912 ( .A(n1003), .B(n9303), .Z(n9302) );
  XOR U8913 ( .A(n9304), .B(n9301), .Z(n9303) );
  XNOR U8914 ( .A(n2017), .B(n9297), .Z(n9299) );
  XOR U8915 ( .A(n9305), .B(n9306), .Z(n2017) );
  AND U8916 ( .A(n1000), .B(n9307), .Z(n9306) );
  XOR U8917 ( .A(n9308), .B(n9305), .Z(n9307) );
  XOR U8918 ( .A(n9309), .B(n9310), .Z(n9297) );
  AND U8919 ( .A(n9311), .B(n9312), .Z(n9310) );
  XOR U8920 ( .A(n9309), .B(n2032), .Z(n9312) );
  XOR U8921 ( .A(n9313), .B(n9314), .Z(n2032) );
  AND U8922 ( .A(n1003), .B(n9315), .Z(n9314) );
  XOR U8923 ( .A(n9316), .B(n9313), .Z(n9315) );
  XNOR U8924 ( .A(n2029), .B(n9309), .Z(n9311) );
  XOR U8925 ( .A(n9317), .B(n9318), .Z(n2029) );
  AND U8926 ( .A(n1000), .B(n9319), .Z(n9318) );
  XOR U8927 ( .A(n9320), .B(n9317), .Z(n9319) );
  XOR U8928 ( .A(n9321), .B(n9322), .Z(n9309) );
  AND U8929 ( .A(n9323), .B(n9324), .Z(n9322) );
  XOR U8930 ( .A(n9321), .B(n2044), .Z(n9324) );
  XOR U8931 ( .A(n9325), .B(n9326), .Z(n2044) );
  AND U8932 ( .A(n1003), .B(n9327), .Z(n9326) );
  XOR U8933 ( .A(n9328), .B(n9325), .Z(n9327) );
  XNOR U8934 ( .A(n2041), .B(n9321), .Z(n9323) );
  XOR U8935 ( .A(n9329), .B(n9330), .Z(n2041) );
  AND U8936 ( .A(n1000), .B(n9331), .Z(n9330) );
  XOR U8937 ( .A(n9332), .B(n9329), .Z(n9331) );
  XOR U8938 ( .A(n9333), .B(n9334), .Z(n9321) );
  AND U8939 ( .A(n9335), .B(n9336), .Z(n9334) );
  XOR U8940 ( .A(n9333), .B(n2056), .Z(n9336) );
  XOR U8941 ( .A(n9337), .B(n9338), .Z(n2056) );
  AND U8942 ( .A(n1003), .B(n9339), .Z(n9338) );
  XOR U8943 ( .A(n9340), .B(n9337), .Z(n9339) );
  XNOR U8944 ( .A(n2053), .B(n9333), .Z(n9335) );
  XOR U8945 ( .A(n9341), .B(n9342), .Z(n2053) );
  AND U8946 ( .A(n1000), .B(n9343), .Z(n9342) );
  XOR U8947 ( .A(n9344), .B(n9341), .Z(n9343) );
  XOR U8948 ( .A(n9345), .B(n9346), .Z(n9333) );
  AND U8949 ( .A(n9347), .B(n9348), .Z(n9346) );
  XOR U8950 ( .A(n9345), .B(n2068), .Z(n9348) );
  XOR U8951 ( .A(n9349), .B(n9350), .Z(n2068) );
  AND U8952 ( .A(n1003), .B(n9351), .Z(n9350) );
  XOR U8953 ( .A(n9352), .B(n9349), .Z(n9351) );
  XNOR U8954 ( .A(n2065), .B(n9345), .Z(n9347) );
  XOR U8955 ( .A(n9353), .B(n9354), .Z(n2065) );
  AND U8956 ( .A(n1000), .B(n9355), .Z(n9354) );
  XOR U8957 ( .A(n9356), .B(n9353), .Z(n9355) );
  XOR U8958 ( .A(n9357), .B(n9358), .Z(n9345) );
  AND U8959 ( .A(n9359), .B(n9360), .Z(n9358) );
  XOR U8960 ( .A(n9357), .B(n2080), .Z(n9360) );
  XOR U8961 ( .A(n9361), .B(n9362), .Z(n2080) );
  AND U8962 ( .A(n1003), .B(n9363), .Z(n9362) );
  XOR U8963 ( .A(n9364), .B(n9361), .Z(n9363) );
  XNOR U8964 ( .A(n2077), .B(n9357), .Z(n9359) );
  XOR U8965 ( .A(n9365), .B(n9366), .Z(n2077) );
  AND U8966 ( .A(n1000), .B(n9367), .Z(n9366) );
  XOR U8967 ( .A(n9368), .B(n9365), .Z(n9367) );
  XOR U8968 ( .A(n9369), .B(n9370), .Z(n9357) );
  AND U8969 ( .A(n9371), .B(n9372), .Z(n9370) );
  XOR U8970 ( .A(n9369), .B(n2092), .Z(n9372) );
  XOR U8971 ( .A(n9373), .B(n9374), .Z(n2092) );
  AND U8972 ( .A(n1003), .B(n9375), .Z(n9374) );
  XOR U8973 ( .A(n9376), .B(n9373), .Z(n9375) );
  XNOR U8974 ( .A(n2089), .B(n9369), .Z(n9371) );
  XOR U8975 ( .A(n9377), .B(n9378), .Z(n2089) );
  AND U8976 ( .A(n1000), .B(n9379), .Z(n9378) );
  XOR U8977 ( .A(n9380), .B(n9377), .Z(n9379) );
  XOR U8978 ( .A(n9381), .B(n9382), .Z(n9369) );
  AND U8979 ( .A(n9383), .B(n9384), .Z(n9382) );
  XOR U8980 ( .A(n9381), .B(n2104), .Z(n9384) );
  XOR U8981 ( .A(n9385), .B(n9386), .Z(n2104) );
  AND U8982 ( .A(n1003), .B(n9387), .Z(n9386) );
  XOR U8983 ( .A(n9388), .B(n9385), .Z(n9387) );
  XNOR U8984 ( .A(n2101), .B(n9381), .Z(n9383) );
  XOR U8985 ( .A(n9389), .B(n9390), .Z(n2101) );
  AND U8986 ( .A(n1000), .B(n9391), .Z(n9390) );
  XOR U8987 ( .A(n9392), .B(n9389), .Z(n9391) );
  XOR U8988 ( .A(n9393), .B(n9394), .Z(n9381) );
  AND U8989 ( .A(n9395), .B(n9396), .Z(n9394) );
  XOR U8990 ( .A(n9393), .B(n2116), .Z(n9396) );
  XOR U8991 ( .A(n9397), .B(n9398), .Z(n2116) );
  AND U8992 ( .A(n1003), .B(n9399), .Z(n9398) );
  XOR U8993 ( .A(n9400), .B(n9397), .Z(n9399) );
  XNOR U8994 ( .A(n2113), .B(n9393), .Z(n9395) );
  XOR U8995 ( .A(n9401), .B(n9402), .Z(n2113) );
  AND U8996 ( .A(n1000), .B(n9403), .Z(n9402) );
  XOR U8997 ( .A(n9404), .B(n9401), .Z(n9403) );
  XOR U8998 ( .A(n9405), .B(n9406), .Z(n9393) );
  AND U8999 ( .A(n9407), .B(n9408), .Z(n9406) );
  XOR U9000 ( .A(n9405), .B(n2128), .Z(n9408) );
  XOR U9001 ( .A(n9409), .B(n9410), .Z(n2128) );
  AND U9002 ( .A(n1003), .B(n9411), .Z(n9410) );
  XOR U9003 ( .A(n9412), .B(n9409), .Z(n9411) );
  XNOR U9004 ( .A(n2125), .B(n9405), .Z(n9407) );
  XOR U9005 ( .A(n9413), .B(n9414), .Z(n2125) );
  AND U9006 ( .A(n1000), .B(n9415), .Z(n9414) );
  XOR U9007 ( .A(n9416), .B(n9413), .Z(n9415) );
  XOR U9008 ( .A(n9417), .B(n9418), .Z(n9405) );
  AND U9009 ( .A(n9419), .B(n9420), .Z(n9418) );
  XOR U9010 ( .A(n9417), .B(n2140), .Z(n9420) );
  XOR U9011 ( .A(n9421), .B(n9422), .Z(n2140) );
  AND U9012 ( .A(n1003), .B(n9423), .Z(n9422) );
  XOR U9013 ( .A(n9424), .B(n9421), .Z(n9423) );
  XNOR U9014 ( .A(n2137), .B(n9417), .Z(n9419) );
  XOR U9015 ( .A(n9425), .B(n9426), .Z(n2137) );
  AND U9016 ( .A(n1000), .B(n9427), .Z(n9426) );
  XOR U9017 ( .A(n9428), .B(n9425), .Z(n9427) );
  XOR U9018 ( .A(n9429), .B(n9430), .Z(n9417) );
  AND U9019 ( .A(n9431), .B(n9432), .Z(n9430) );
  XOR U9020 ( .A(n9429), .B(n2152), .Z(n9432) );
  XOR U9021 ( .A(n9433), .B(n9434), .Z(n2152) );
  AND U9022 ( .A(n1003), .B(n9435), .Z(n9434) );
  XOR U9023 ( .A(n9436), .B(n9433), .Z(n9435) );
  XNOR U9024 ( .A(n2149), .B(n9429), .Z(n9431) );
  XOR U9025 ( .A(n9437), .B(n9438), .Z(n2149) );
  AND U9026 ( .A(n1000), .B(n9439), .Z(n9438) );
  XOR U9027 ( .A(n9440), .B(n9437), .Z(n9439) );
  XOR U9028 ( .A(n9441), .B(n9442), .Z(n9429) );
  AND U9029 ( .A(n9443), .B(n9444), .Z(n9442) );
  XOR U9030 ( .A(n9441), .B(n2164), .Z(n9444) );
  XOR U9031 ( .A(n9445), .B(n9446), .Z(n2164) );
  AND U9032 ( .A(n1003), .B(n9447), .Z(n9446) );
  XOR U9033 ( .A(n9448), .B(n9445), .Z(n9447) );
  XNOR U9034 ( .A(n2161), .B(n9441), .Z(n9443) );
  XOR U9035 ( .A(n9449), .B(n9450), .Z(n2161) );
  AND U9036 ( .A(n1000), .B(n9451), .Z(n9450) );
  XOR U9037 ( .A(n9452), .B(n9449), .Z(n9451) );
  XOR U9038 ( .A(n9453), .B(n9454), .Z(n9441) );
  AND U9039 ( .A(n9455), .B(n9456), .Z(n9454) );
  XOR U9040 ( .A(n9453), .B(n2176), .Z(n9456) );
  XOR U9041 ( .A(n9457), .B(n9458), .Z(n2176) );
  AND U9042 ( .A(n1003), .B(n9459), .Z(n9458) );
  XOR U9043 ( .A(n9460), .B(n9457), .Z(n9459) );
  XNOR U9044 ( .A(n2173), .B(n9453), .Z(n9455) );
  XOR U9045 ( .A(n9461), .B(n9462), .Z(n2173) );
  AND U9046 ( .A(n1000), .B(n9463), .Z(n9462) );
  XOR U9047 ( .A(n9464), .B(n9461), .Z(n9463) );
  XOR U9048 ( .A(n9465), .B(n9466), .Z(n9453) );
  AND U9049 ( .A(n9467), .B(n9468), .Z(n9466) );
  XOR U9050 ( .A(n9465), .B(n2188), .Z(n9468) );
  XOR U9051 ( .A(n9469), .B(n9470), .Z(n2188) );
  AND U9052 ( .A(n1003), .B(n9471), .Z(n9470) );
  XOR U9053 ( .A(n9472), .B(n9469), .Z(n9471) );
  XNOR U9054 ( .A(n2185), .B(n9465), .Z(n9467) );
  XOR U9055 ( .A(n9473), .B(n9474), .Z(n2185) );
  AND U9056 ( .A(n1000), .B(n9475), .Z(n9474) );
  XOR U9057 ( .A(n9476), .B(n9473), .Z(n9475) );
  XOR U9058 ( .A(n9477), .B(n9478), .Z(n9465) );
  AND U9059 ( .A(n9479), .B(n9480), .Z(n9478) );
  XOR U9060 ( .A(n9477), .B(n2200), .Z(n9480) );
  XOR U9061 ( .A(n9481), .B(n9482), .Z(n2200) );
  AND U9062 ( .A(n1003), .B(n9483), .Z(n9482) );
  XOR U9063 ( .A(n9484), .B(n9481), .Z(n9483) );
  XNOR U9064 ( .A(n2197), .B(n9477), .Z(n9479) );
  XOR U9065 ( .A(n9485), .B(n9486), .Z(n2197) );
  AND U9066 ( .A(n1000), .B(n9487), .Z(n9486) );
  XOR U9067 ( .A(n9488), .B(n9485), .Z(n9487) );
  XOR U9068 ( .A(n9489), .B(n9490), .Z(n9477) );
  AND U9069 ( .A(n9491), .B(n9492), .Z(n9490) );
  XOR U9070 ( .A(n9489), .B(n2212), .Z(n9492) );
  XOR U9071 ( .A(n9493), .B(n9494), .Z(n2212) );
  AND U9072 ( .A(n1003), .B(n9495), .Z(n9494) );
  XOR U9073 ( .A(n9496), .B(n9493), .Z(n9495) );
  XNOR U9074 ( .A(n2209), .B(n9489), .Z(n9491) );
  XOR U9075 ( .A(n9497), .B(n9498), .Z(n2209) );
  AND U9076 ( .A(n1000), .B(n9499), .Z(n9498) );
  XOR U9077 ( .A(n9500), .B(n9497), .Z(n9499) );
  XOR U9078 ( .A(n9501), .B(n9502), .Z(n9489) );
  AND U9079 ( .A(n9503), .B(n9504), .Z(n9502) );
  XOR U9080 ( .A(n9501), .B(n2224), .Z(n9504) );
  XOR U9081 ( .A(n9505), .B(n9506), .Z(n2224) );
  AND U9082 ( .A(n1003), .B(n9507), .Z(n9506) );
  XOR U9083 ( .A(n9508), .B(n9505), .Z(n9507) );
  XNOR U9084 ( .A(n2221), .B(n9501), .Z(n9503) );
  XOR U9085 ( .A(n9509), .B(n9510), .Z(n2221) );
  AND U9086 ( .A(n1000), .B(n9511), .Z(n9510) );
  XOR U9087 ( .A(n9512), .B(n9509), .Z(n9511) );
  XOR U9088 ( .A(n9513), .B(n9514), .Z(n9501) );
  AND U9089 ( .A(n9515), .B(n9516), .Z(n9514) );
  XOR U9090 ( .A(n9513), .B(n2236), .Z(n9516) );
  XOR U9091 ( .A(n9517), .B(n9518), .Z(n2236) );
  AND U9092 ( .A(n1003), .B(n9519), .Z(n9518) );
  XOR U9093 ( .A(n9520), .B(n9517), .Z(n9519) );
  XNOR U9094 ( .A(n2233), .B(n9513), .Z(n9515) );
  XOR U9095 ( .A(n9521), .B(n9522), .Z(n2233) );
  AND U9096 ( .A(n1000), .B(n9523), .Z(n9522) );
  XOR U9097 ( .A(n9524), .B(n9521), .Z(n9523) );
  XOR U9098 ( .A(n9525), .B(n9526), .Z(n9513) );
  AND U9099 ( .A(n9527), .B(n9528), .Z(n9526) );
  XOR U9100 ( .A(n9525), .B(n2248), .Z(n9528) );
  XOR U9101 ( .A(n9529), .B(n9530), .Z(n2248) );
  AND U9102 ( .A(n1003), .B(n9531), .Z(n9530) );
  XOR U9103 ( .A(n9532), .B(n9529), .Z(n9531) );
  XNOR U9104 ( .A(n2245), .B(n9525), .Z(n9527) );
  XOR U9105 ( .A(n9533), .B(n9534), .Z(n2245) );
  AND U9106 ( .A(n1000), .B(n9535), .Z(n9534) );
  XOR U9107 ( .A(n9536), .B(n9533), .Z(n9535) );
  XOR U9108 ( .A(n9537), .B(n9538), .Z(n9525) );
  AND U9109 ( .A(n9539), .B(n9540), .Z(n9538) );
  XOR U9110 ( .A(n9537), .B(n2260), .Z(n9540) );
  XOR U9111 ( .A(n9541), .B(n9542), .Z(n2260) );
  AND U9112 ( .A(n1003), .B(n9543), .Z(n9542) );
  XOR U9113 ( .A(n9544), .B(n9541), .Z(n9543) );
  XNOR U9114 ( .A(n2257), .B(n9537), .Z(n9539) );
  XOR U9115 ( .A(n9545), .B(n9546), .Z(n2257) );
  AND U9116 ( .A(n1000), .B(n9547), .Z(n9546) );
  XOR U9117 ( .A(n9548), .B(n9545), .Z(n9547) );
  XOR U9118 ( .A(n9549), .B(n9550), .Z(n9537) );
  AND U9119 ( .A(n9551), .B(n9552), .Z(n9550) );
  XNOR U9120 ( .A(n9553), .B(n2273), .Z(n9552) );
  XOR U9121 ( .A(n9554), .B(n9555), .Z(n2273) );
  AND U9122 ( .A(n1003), .B(n9556), .Z(n9555) );
  XOR U9123 ( .A(n9554), .B(n9557), .Z(n9556) );
  XNOR U9124 ( .A(n2270), .B(n9549), .Z(n9551) );
  XOR U9125 ( .A(n9558), .B(n9559), .Z(n2270) );
  AND U9126 ( .A(n1000), .B(n9560), .Z(n9559) );
  XOR U9127 ( .A(n9558), .B(n9561), .Z(n9560) );
  IV U9128 ( .A(n9553), .Z(n9549) );
  AND U9129 ( .A(n9185), .B(n9188), .Z(n9553) );
  XNOR U9130 ( .A(n9562), .B(n9563), .Z(n9188) );
  AND U9131 ( .A(n1003), .B(n9564), .Z(n9563) );
  XNOR U9132 ( .A(n9565), .B(n9562), .Z(n9564) );
  XOR U9133 ( .A(n9566), .B(n9567), .Z(n1003) );
  AND U9134 ( .A(n9568), .B(n9569), .Z(n9567) );
  XOR U9135 ( .A(n9566), .B(n9196), .Z(n9569) );
  XOR U9136 ( .A(n9570), .B(n9571), .Z(n9196) );
  AND U9137 ( .A(n827), .B(n9572), .Z(n9571) );
  XOR U9138 ( .A(n9573), .B(n9570), .Z(n9572) );
  XNOR U9139 ( .A(n9193), .B(n9566), .Z(n9568) );
  XOR U9140 ( .A(n9574), .B(n9575), .Z(n9193) );
  AND U9141 ( .A(n825), .B(n9576), .Z(n9575) );
  XOR U9142 ( .A(n9577), .B(n9574), .Z(n9576) );
  XOR U9143 ( .A(n9578), .B(n9579), .Z(n9566) );
  AND U9144 ( .A(n9580), .B(n9581), .Z(n9579) );
  XOR U9145 ( .A(n9578), .B(n9208), .Z(n9581) );
  XOR U9146 ( .A(n9582), .B(n9583), .Z(n9208) );
  AND U9147 ( .A(n827), .B(n9584), .Z(n9583) );
  XOR U9148 ( .A(n9585), .B(n9582), .Z(n9584) );
  XNOR U9149 ( .A(n9205), .B(n9578), .Z(n9580) );
  XOR U9150 ( .A(n9586), .B(n9587), .Z(n9205) );
  AND U9151 ( .A(n825), .B(n9588), .Z(n9587) );
  XOR U9152 ( .A(n9589), .B(n9586), .Z(n9588) );
  XOR U9153 ( .A(n9590), .B(n9591), .Z(n9578) );
  AND U9154 ( .A(n9592), .B(n9593), .Z(n9591) );
  XOR U9155 ( .A(n9590), .B(n9220), .Z(n9593) );
  XOR U9156 ( .A(n9594), .B(n9595), .Z(n9220) );
  AND U9157 ( .A(n827), .B(n9596), .Z(n9595) );
  XOR U9158 ( .A(n9597), .B(n9594), .Z(n9596) );
  XNOR U9159 ( .A(n9217), .B(n9590), .Z(n9592) );
  XOR U9160 ( .A(n9598), .B(n9599), .Z(n9217) );
  AND U9161 ( .A(n825), .B(n9600), .Z(n9599) );
  XOR U9162 ( .A(n9601), .B(n9598), .Z(n9600) );
  XOR U9163 ( .A(n9602), .B(n9603), .Z(n9590) );
  AND U9164 ( .A(n9604), .B(n9605), .Z(n9603) );
  XOR U9165 ( .A(n9602), .B(n9232), .Z(n9605) );
  XOR U9166 ( .A(n9606), .B(n9607), .Z(n9232) );
  AND U9167 ( .A(n827), .B(n9608), .Z(n9607) );
  XOR U9168 ( .A(n9609), .B(n9606), .Z(n9608) );
  XNOR U9169 ( .A(n9229), .B(n9602), .Z(n9604) );
  XOR U9170 ( .A(n9610), .B(n9611), .Z(n9229) );
  AND U9171 ( .A(n825), .B(n9612), .Z(n9611) );
  XOR U9172 ( .A(n9613), .B(n9610), .Z(n9612) );
  XOR U9173 ( .A(n9614), .B(n9615), .Z(n9602) );
  AND U9174 ( .A(n9616), .B(n9617), .Z(n9615) );
  XOR U9175 ( .A(n9614), .B(n9244), .Z(n9617) );
  XOR U9176 ( .A(n9618), .B(n9619), .Z(n9244) );
  AND U9177 ( .A(n827), .B(n9620), .Z(n9619) );
  XOR U9178 ( .A(n9621), .B(n9618), .Z(n9620) );
  XNOR U9179 ( .A(n9241), .B(n9614), .Z(n9616) );
  XOR U9180 ( .A(n9622), .B(n9623), .Z(n9241) );
  AND U9181 ( .A(n825), .B(n9624), .Z(n9623) );
  XOR U9182 ( .A(n9625), .B(n9622), .Z(n9624) );
  XOR U9183 ( .A(n9626), .B(n9627), .Z(n9614) );
  AND U9184 ( .A(n9628), .B(n9629), .Z(n9627) );
  XOR U9185 ( .A(n9626), .B(n9256), .Z(n9629) );
  XOR U9186 ( .A(n9630), .B(n9631), .Z(n9256) );
  AND U9187 ( .A(n827), .B(n9632), .Z(n9631) );
  XOR U9188 ( .A(n9633), .B(n9630), .Z(n9632) );
  XNOR U9189 ( .A(n9253), .B(n9626), .Z(n9628) );
  XOR U9190 ( .A(n9634), .B(n9635), .Z(n9253) );
  AND U9191 ( .A(n825), .B(n9636), .Z(n9635) );
  XOR U9192 ( .A(n9637), .B(n9634), .Z(n9636) );
  XOR U9193 ( .A(n9638), .B(n9639), .Z(n9626) );
  AND U9194 ( .A(n9640), .B(n9641), .Z(n9639) );
  XOR U9195 ( .A(n9638), .B(n9268), .Z(n9641) );
  XOR U9196 ( .A(n9642), .B(n9643), .Z(n9268) );
  AND U9197 ( .A(n827), .B(n9644), .Z(n9643) );
  XOR U9198 ( .A(n9645), .B(n9642), .Z(n9644) );
  XNOR U9199 ( .A(n9265), .B(n9638), .Z(n9640) );
  XOR U9200 ( .A(n9646), .B(n9647), .Z(n9265) );
  AND U9201 ( .A(n825), .B(n9648), .Z(n9647) );
  XOR U9202 ( .A(n9649), .B(n9646), .Z(n9648) );
  XOR U9203 ( .A(n9650), .B(n9651), .Z(n9638) );
  AND U9204 ( .A(n9652), .B(n9653), .Z(n9651) );
  XOR U9205 ( .A(n9650), .B(n9280), .Z(n9653) );
  XOR U9206 ( .A(n9654), .B(n9655), .Z(n9280) );
  AND U9207 ( .A(n827), .B(n9656), .Z(n9655) );
  XOR U9208 ( .A(n9657), .B(n9654), .Z(n9656) );
  XNOR U9209 ( .A(n9277), .B(n9650), .Z(n9652) );
  XOR U9210 ( .A(n9658), .B(n9659), .Z(n9277) );
  AND U9211 ( .A(n825), .B(n9660), .Z(n9659) );
  XOR U9212 ( .A(n9661), .B(n9658), .Z(n9660) );
  XOR U9213 ( .A(n9662), .B(n9663), .Z(n9650) );
  AND U9214 ( .A(n9664), .B(n9665), .Z(n9663) );
  XOR U9215 ( .A(n9662), .B(n9292), .Z(n9665) );
  XOR U9216 ( .A(n9666), .B(n9667), .Z(n9292) );
  AND U9217 ( .A(n827), .B(n9668), .Z(n9667) );
  XOR U9218 ( .A(n9669), .B(n9666), .Z(n9668) );
  XNOR U9219 ( .A(n9289), .B(n9662), .Z(n9664) );
  XOR U9220 ( .A(n9670), .B(n9671), .Z(n9289) );
  AND U9221 ( .A(n825), .B(n9672), .Z(n9671) );
  XOR U9222 ( .A(n9673), .B(n9670), .Z(n9672) );
  XOR U9223 ( .A(n9674), .B(n9675), .Z(n9662) );
  AND U9224 ( .A(n9676), .B(n9677), .Z(n9675) );
  XOR U9225 ( .A(n9674), .B(n9304), .Z(n9677) );
  XOR U9226 ( .A(n9678), .B(n9679), .Z(n9304) );
  AND U9227 ( .A(n827), .B(n9680), .Z(n9679) );
  XOR U9228 ( .A(n9681), .B(n9678), .Z(n9680) );
  XNOR U9229 ( .A(n9301), .B(n9674), .Z(n9676) );
  XOR U9230 ( .A(n9682), .B(n9683), .Z(n9301) );
  AND U9231 ( .A(n825), .B(n9684), .Z(n9683) );
  XOR U9232 ( .A(n9685), .B(n9682), .Z(n9684) );
  XOR U9233 ( .A(n9686), .B(n9687), .Z(n9674) );
  AND U9234 ( .A(n9688), .B(n9689), .Z(n9687) );
  XOR U9235 ( .A(n9686), .B(n9316), .Z(n9689) );
  XOR U9236 ( .A(n9690), .B(n9691), .Z(n9316) );
  AND U9237 ( .A(n827), .B(n9692), .Z(n9691) );
  XOR U9238 ( .A(n9693), .B(n9690), .Z(n9692) );
  XNOR U9239 ( .A(n9313), .B(n9686), .Z(n9688) );
  XOR U9240 ( .A(n9694), .B(n9695), .Z(n9313) );
  AND U9241 ( .A(n825), .B(n9696), .Z(n9695) );
  XOR U9242 ( .A(n9697), .B(n9694), .Z(n9696) );
  XOR U9243 ( .A(n9698), .B(n9699), .Z(n9686) );
  AND U9244 ( .A(n9700), .B(n9701), .Z(n9699) );
  XOR U9245 ( .A(n9698), .B(n9328), .Z(n9701) );
  XOR U9246 ( .A(n9702), .B(n9703), .Z(n9328) );
  AND U9247 ( .A(n827), .B(n9704), .Z(n9703) );
  XOR U9248 ( .A(n9705), .B(n9702), .Z(n9704) );
  XNOR U9249 ( .A(n9325), .B(n9698), .Z(n9700) );
  XOR U9250 ( .A(n9706), .B(n9707), .Z(n9325) );
  AND U9251 ( .A(n825), .B(n9708), .Z(n9707) );
  XOR U9252 ( .A(n9709), .B(n9706), .Z(n9708) );
  XOR U9253 ( .A(n9710), .B(n9711), .Z(n9698) );
  AND U9254 ( .A(n9712), .B(n9713), .Z(n9711) );
  XOR U9255 ( .A(n9710), .B(n9340), .Z(n9713) );
  XOR U9256 ( .A(n9714), .B(n9715), .Z(n9340) );
  AND U9257 ( .A(n827), .B(n9716), .Z(n9715) );
  XOR U9258 ( .A(n9717), .B(n9714), .Z(n9716) );
  XNOR U9259 ( .A(n9337), .B(n9710), .Z(n9712) );
  XOR U9260 ( .A(n9718), .B(n9719), .Z(n9337) );
  AND U9261 ( .A(n825), .B(n9720), .Z(n9719) );
  XOR U9262 ( .A(n9721), .B(n9718), .Z(n9720) );
  XOR U9263 ( .A(n9722), .B(n9723), .Z(n9710) );
  AND U9264 ( .A(n9724), .B(n9725), .Z(n9723) );
  XOR U9265 ( .A(n9722), .B(n9352), .Z(n9725) );
  XOR U9266 ( .A(n9726), .B(n9727), .Z(n9352) );
  AND U9267 ( .A(n827), .B(n9728), .Z(n9727) );
  XOR U9268 ( .A(n9729), .B(n9726), .Z(n9728) );
  XNOR U9269 ( .A(n9349), .B(n9722), .Z(n9724) );
  XOR U9270 ( .A(n9730), .B(n9731), .Z(n9349) );
  AND U9271 ( .A(n825), .B(n9732), .Z(n9731) );
  XOR U9272 ( .A(n9733), .B(n9730), .Z(n9732) );
  XOR U9273 ( .A(n9734), .B(n9735), .Z(n9722) );
  AND U9274 ( .A(n9736), .B(n9737), .Z(n9735) );
  XOR U9275 ( .A(n9734), .B(n9364), .Z(n9737) );
  XOR U9276 ( .A(n9738), .B(n9739), .Z(n9364) );
  AND U9277 ( .A(n827), .B(n9740), .Z(n9739) );
  XOR U9278 ( .A(n9741), .B(n9738), .Z(n9740) );
  XNOR U9279 ( .A(n9361), .B(n9734), .Z(n9736) );
  XOR U9280 ( .A(n9742), .B(n9743), .Z(n9361) );
  AND U9281 ( .A(n825), .B(n9744), .Z(n9743) );
  XOR U9282 ( .A(n9745), .B(n9742), .Z(n9744) );
  XOR U9283 ( .A(n9746), .B(n9747), .Z(n9734) );
  AND U9284 ( .A(n9748), .B(n9749), .Z(n9747) );
  XOR U9285 ( .A(n9746), .B(n9376), .Z(n9749) );
  XOR U9286 ( .A(n9750), .B(n9751), .Z(n9376) );
  AND U9287 ( .A(n827), .B(n9752), .Z(n9751) );
  XOR U9288 ( .A(n9753), .B(n9750), .Z(n9752) );
  XNOR U9289 ( .A(n9373), .B(n9746), .Z(n9748) );
  XOR U9290 ( .A(n9754), .B(n9755), .Z(n9373) );
  AND U9291 ( .A(n825), .B(n9756), .Z(n9755) );
  XOR U9292 ( .A(n9757), .B(n9754), .Z(n9756) );
  XOR U9293 ( .A(n9758), .B(n9759), .Z(n9746) );
  AND U9294 ( .A(n9760), .B(n9761), .Z(n9759) );
  XOR U9295 ( .A(n9758), .B(n9388), .Z(n9761) );
  XOR U9296 ( .A(n9762), .B(n9763), .Z(n9388) );
  AND U9297 ( .A(n827), .B(n9764), .Z(n9763) );
  XOR U9298 ( .A(n9765), .B(n9762), .Z(n9764) );
  XNOR U9299 ( .A(n9385), .B(n9758), .Z(n9760) );
  XOR U9300 ( .A(n9766), .B(n9767), .Z(n9385) );
  AND U9301 ( .A(n825), .B(n9768), .Z(n9767) );
  XOR U9302 ( .A(n9769), .B(n9766), .Z(n9768) );
  XOR U9303 ( .A(n9770), .B(n9771), .Z(n9758) );
  AND U9304 ( .A(n9772), .B(n9773), .Z(n9771) );
  XOR U9305 ( .A(n9770), .B(n9400), .Z(n9773) );
  XOR U9306 ( .A(n9774), .B(n9775), .Z(n9400) );
  AND U9307 ( .A(n827), .B(n9776), .Z(n9775) );
  XOR U9308 ( .A(n9777), .B(n9774), .Z(n9776) );
  XNOR U9309 ( .A(n9397), .B(n9770), .Z(n9772) );
  XOR U9310 ( .A(n9778), .B(n9779), .Z(n9397) );
  AND U9311 ( .A(n825), .B(n9780), .Z(n9779) );
  XOR U9312 ( .A(n9781), .B(n9778), .Z(n9780) );
  XOR U9313 ( .A(n9782), .B(n9783), .Z(n9770) );
  AND U9314 ( .A(n9784), .B(n9785), .Z(n9783) );
  XOR U9315 ( .A(n9782), .B(n9412), .Z(n9785) );
  XOR U9316 ( .A(n9786), .B(n9787), .Z(n9412) );
  AND U9317 ( .A(n827), .B(n9788), .Z(n9787) );
  XOR U9318 ( .A(n9789), .B(n9786), .Z(n9788) );
  XNOR U9319 ( .A(n9409), .B(n9782), .Z(n9784) );
  XOR U9320 ( .A(n9790), .B(n9791), .Z(n9409) );
  AND U9321 ( .A(n825), .B(n9792), .Z(n9791) );
  XOR U9322 ( .A(n9793), .B(n9790), .Z(n9792) );
  XOR U9323 ( .A(n9794), .B(n9795), .Z(n9782) );
  AND U9324 ( .A(n9796), .B(n9797), .Z(n9795) );
  XOR U9325 ( .A(n9794), .B(n9424), .Z(n9797) );
  XOR U9326 ( .A(n9798), .B(n9799), .Z(n9424) );
  AND U9327 ( .A(n827), .B(n9800), .Z(n9799) );
  XOR U9328 ( .A(n9801), .B(n9798), .Z(n9800) );
  XNOR U9329 ( .A(n9421), .B(n9794), .Z(n9796) );
  XOR U9330 ( .A(n9802), .B(n9803), .Z(n9421) );
  AND U9331 ( .A(n825), .B(n9804), .Z(n9803) );
  XOR U9332 ( .A(n9805), .B(n9802), .Z(n9804) );
  XOR U9333 ( .A(n9806), .B(n9807), .Z(n9794) );
  AND U9334 ( .A(n9808), .B(n9809), .Z(n9807) );
  XOR U9335 ( .A(n9806), .B(n9436), .Z(n9809) );
  XOR U9336 ( .A(n9810), .B(n9811), .Z(n9436) );
  AND U9337 ( .A(n827), .B(n9812), .Z(n9811) );
  XOR U9338 ( .A(n9813), .B(n9810), .Z(n9812) );
  XNOR U9339 ( .A(n9433), .B(n9806), .Z(n9808) );
  XOR U9340 ( .A(n9814), .B(n9815), .Z(n9433) );
  AND U9341 ( .A(n825), .B(n9816), .Z(n9815) );
  XOR U9342 ( .A(n9817), .B(n9814), .Z(n9816) );
  XOR U9343 ( .A(n9818), .B(n9819), .Z(n9806) );
  AND U9344 ( .A(n9820), .B(n9821), .Z(n9819) );
  XOR U9345 ( .A(n9818), .B(n9448), .Z(n9821) );
  XOR U9346 ( .A(n9822), .B(n9823), .Z(n9448) );
  AND U9347 ( .A(n827), .B(n9824), .Z(n9823) );
  XOR U9348 ( .A(n9825), .B(n9822), .Z(n9824) );
  XNOR U9349 ( .A(n9445), .B(n9818), .Z(n9820) );
  XOR U9350 ( .A(n9826), .B(n9827), .Z(n9445) );
  AND U9351 ( .A(n825), .B(n9828), .Z(n9827) );
  XOR U9352 ( .A(n9829), .B(n9826), .Z(n9828) );
  XOR U9353 ( .A(n9830), .B(n9831), .Z(n9818) );
  AND U9354 ( .A(n9832), .B(n9833), .Z(n9831) );
  XOR U9355 ( .A(n9830), .B(n9460), .Z(n9833) );
  XOR U9356 ( .A(n9834), .B(n9835), .Z(n9460) );
  AND U9357 ( .A(n827), .B(n9836), .Z(n9835) );
  XOR U9358 ( .A(n9837), .B(n9834), .Z(n9836) );
  XNOR U9359 ( .A(n9457), .B(n9830), .Z(n9832) );
  XOR U9360 ( .A(n9838), .B(n9839), .Z(n9457) );
  AND U9361 ( .A(n825), .B(n9840), .Z(n9839) );
  XOR U9362 ( .A(n9841), .B(n9838), .Z(n9840) );
  XOR U9363 ( .A(n9842), .B(n9843), .Z(n9830) );
  AND U9364 ( .A(n9844), .B(n9845), .Z(n9843) );
  XOR U9365 ( .A(n9842), .B(n9472), .Z(n9845) );
  XOR U9366 ( .A(n9846), .B(n9847), .Z(n9472) );
  AND U9367 ( .A(n827), .B(n9848), .Z(n9847) );
  XOR U9368 ( .A(n9849), .B(n9846), .Z(n9848) );
  XNOR U9369 ( .A(n9469), .B(n9842), .Z(n9844) );
  XOR U9370 ( .A(n9850), .B(n9851), .Z(n9469) );
  AND U9371 ( .A(n825), .B(n9852), .Z(n9851) );
  XOR U9372 ( .A(n9853), .B(n9850), .Z(n9852) );
  XOR U9373 ( .A(n9854), .B(n9855), .Z(n9842) );
  AND U9374 ( .A(n9856), .B(n9857), .Z(n9855) );
  XOR U9375 ( .A(n9854), .B(n9484), .Z(n9857) );
  XOR U9376 ( .A(n9858), .B(n9859), .Z(n9484) );
  AND U9377 ( .A(n827), .B(n9860), .Z(n9859) );
  XOR U9378 ( .A(n9861), .B(n9858), .Z(n9860) );
  XNOR U9379 ( .A(n9481), .B(n9854), .Z(n9856) );
  XOR U9380 ( .A(n9862), .B(n9863), .Z(n9481) );
  AND U9381 ( .A(n825), .B(n9864), .Z(n9863) );
  XOR U9382 ( .A(n9865), .B(n9862), .Z(n9864) );
  XOR U9383 ( .A(n9866), .B(n9867), .Z(n9854) );
  AND U9384 ( .A(n9868), .B(n9869), .Z(n9867) );
  XOR U9385 ( .A(n9866), .B(n9496), .Z(n9869) );
  XOR U9386 ( .A(n9870), .B(n9871), .Z(n9496) );
  AND U9387 ( .A(n827), .B(n9872), .Z(n9871) );
  XOR U9388 ( .A(n9873), .B(n9870), .Z(n9872) );
  XNOR U9389 ( .A(n9493), .B(n9866), .Z(n9868) );
  XOR U9390 ( .A(n9874), .B(n9875), .Z(n9493) );
  AND U9391 ( .A(n825), .B(n9876), .Z(n9875) );
  XOR U9392 ( .A(n9877), .B(n9874), .Z(n9876) );
  XOR U9393 ( .A(n9878), .B(n9879), .Z(n9866) );
  AND U9394 ( .A(n9880), .B(n9881), .Z(n9879) );
  XOR U9395 ( .A(n9878), .B(n9508), .Z(n9881) );
  XOR U9396 ( .A(n9882), .B(n9883), .Z(n9508) );
  AND U9397 ( .A(n827), .B(n9884), .Z(n9883) );
  XOR U9398 ( .A(n9885), .B(n9882), .Z(n9884) );
  XNOR U9399 ( .A(n9505), .B(n9878), .Z(n9880) );
  XOR U9400 ( .A(n9886), .B(n9887), .Z(n9505) );
  AND U9401 ( .A(n825), .B(n9888), .Z(n9887) );
  XOR U9402 ( .A(n9889), .B(n9886), .Z(n9888) );
  XOR U9403 ( .A(n9890), .B(n9891), .Z(n9878) );
  AND U9404 ( .A(n9892), .B(n9893), .Z(n9891) );
  XOR U9405 ( .A(n9890), .B(n9520), .Z(n9893) );
  XOR U9406 ( .A(n9894), .B(n9895), .Z(n9520) );
  AND U9407 ( .A(n827), .B(n9896), .Z(n9895) );
  XOR U9408 ( .A(n9897), .B(n9894), .Z(n9896) );
  XNOR U9409 ( .A(n9517), .B(n9890), .Z(n9892) );
  XOR U9410 ( .A(n9898), .B(n9899), .Z(n9517) );
  AND U9411 ( .A(n825), .B(n9900), .Z(n9899) );
  XOR U9412 ( .A(n9901), .B(n9898), .Z(n9900) );
  XOR U9413 ( .A(n9902), .B(n9903), .Z(n9890) );
  AND U9414 ( .A(n9904), .B(n9905), .Z(n9903) );
  XOR U9415 ( .A(n9902), .B(n9532), .Z(n9905) );
  XOR U9416 ( .A(n9906), .B(n9907), .Z(n9532) );
  AND U9417 ( .A(n827), .B(n9908), .Z(n9907) );
  XOR U9418 ( .A(n9909), .B(n9906), .Z(n9908) );
  XNOR U9419 ( .A(n9529), .B(n9902), .Z(n9904) );
  XOR U9420 ( .A(n9910), .B(n9911), .Z(n9529) );
  AND U9421 ( .A(n825), .B(n9912), .Z(n9911) );
  XOR U9422 ( .A(n9913), .B(n9910), .Z(n9912) );
  XOR U9423 ( .A(n9914), .B(n9915), .Z(n9902) );
  AND U9424 ( .A(n9916), .B(n9917), .Z(n9915) );
  XOR U9425 ( .A(n9914), .B(n9544), .Z(n9917) );
  XOR U9426 ( .A(n9918), .B(n9919), .Z(n9544) );
  AND U9427 ( .A(n827), .B(n9920), .Z(n9919) );
  XOR U9428 ( .A(n9921), .B(n9918), .Z(n9920) );
  XNOR U9429 ( .A(n9541), .B(n9914), .Z(n9916) );
  XOR U9430 ( .A(n9922), .B(n9923), .Z(n9541) );
  AND U9431 ( .A(n825), .B(n9924), .Z(n9923) );
  XOR U9432 ( .A(n9925), .B(n9922), .Z(n9924) );
  XOR U9433 ( .A(n9926), .B(n9927), .Z(n9914) );
  AND U9434 ( .A(n9928), .B(n9929), .Z(n9927) );
  XNOR U9435 ( .A(n9930), .B(n9557), .Z(n9929) );
  XOR U9436 ( .A(n9931), .B(n9932), .Z(n9557) );
  AND U9437 ( .A(n827), .B(n9933), .Z(n9932) );
  XOR U9438 ( .A(n9931), .B(n9934), .Z(n9933) );
  XNOR U9439 ( .A(n9554), .B(n9926), .Z(n9928) );
  XOR U9440 ( .A(n9935), .B(n9936), .Z(n9554) );
  AND U9441 ( .A(n825), .B(n9937), .Z(n9936) );
  XOR U9442 ( .A(n9935), .B(n9938), .Z(n9937) );
  IV U9443 ( .A(n9930), .Z(n9926) );
  AND U9444 ( .A(n9562), .B(n9565), .Z(n9930) );
  XNOR U9445 ( .A(n9939), .B(n9940), .Z(n9565) );
  AND U9446 ( .A(n827), .B(n9941), .Z(n9940) );
  XNOR U9447 ( .A(n9942), .B(n9939), .Z(n9941) );
  XOR U9448 ( .A(n9943), .B(n9944), .Z(n827) );
  AND U9449 ( .A(n9945), .B(n9946), .Z(n9944) );
  XOR U9450 ( .A(n9943), .B(n9573), .Z(n9946) );
  XNOR U9451 ( .A(n9947), .B(n9948), .Z(n9573) );
  AND U9452 ( .A(n9949), .B(n467), .Z(n9948) );
  AND U9453 ( .A(n9947), .B(n9950), .Z(n9949) );
  XNOR U9454 ( .A(n9570), .B(n9943), .Z(n9945) );
  XOR U9455 ( .A(n9951), .B(n9952), .Z(n9570) );
  AND U9456 ( .A(n9953), .B(n465), .Z(n9952) );
  NOR U9457 ( .A(n9951), .B(n9954), .Z(n9953) );
  XOR U9458 ( .A(n9955), .B(n9956), .Z(n9943) );
  AND U9459 ( .A(n9957), .B(n9958), .Z(n9956) );
  XOR U9460 ( .A(n9955), .B(n9585), .Z(n9958) );
  XOR U9461 ( .A(n9959), .B(n9960), .Z(n9585) );
  AND U9462 ( .A(n467), .B(n9961), .Z(n9960) );
  XOR U9463 ( .A(n9962), .B(n9959), .Z(n9961) );
  XNOR U9464 ( .A(n9582), .B(n9955), .Z(n9957) );
  XOR U9465 ( .A(n9963), .B(n9964), .Z(n9582) );
  AND U9466 ( .A(n465), .B(n9965), .Z(n9964) );
  XOR U9467 ( .A(n9966), .B(n9963), .Z(n9965) );
  XOR U9468 ( .A(n9967), .B(n9968), .Z(n9955) );
  AND U9469 ( .A(n9969), .B(n9970), .Z(n9968) );
  XOR U9470 ( .A(n9967), .B(n9597), .Z(n9970) );
  XOR U9471 ( .A(n9971), .B(n9972), .Z(n9597) );
  AND U9472 ( .A(n467), .B(n9973), .Z(n9972) );
  XOR U9473 ( .A(n9974), .B(n9971), .Z(n9973) );
  XNOR U9474 ( .A(n9594), .B(n9967), .Z(n9969) );
  XOR U9475 ( .A(n9975), .B(n9976), .Z(n9594) );
  AND U9476 ( .A(n465), .B(n9977), .Z(n9976) );
  XOR U9477 ( .A(n9978), .B(n9975), .Z(n9977) );
  XOR U9478 ( .A(n9979), .B(n9980), .Z(n9967) );
  AND U9479 ( .A(n9981), .B(n9982), .Z(n9980) );
  XOR U9480 ( .A(n9979), .B(n9609), .Z(n9982) );
  XOR U9481 ( .A(n9983), .B(n9984), .Z(n9609) );
  AND U9482 ( .A(n467), .B(n9985), .Z(n9984) );
  XOR U9483 ( .A(n9986), .B(n9983), .Z(n9985) );
  XNOR U9484 ( .A(n9606), .B(n9979), .Z(n9981) );
  XOR U9485 ( .A(n9987), .B(n9988), .Z(n9606) );
  AND U9486 ( .A(n465), .B(n9989), .Z(n9988) );
  XOR U9487 ( .A(n9990), .B(n9987), .Z(n9989) );
  XOR U9488 ( .A(n9991), .B(n9992), .Z(n9979) );
  AND U9489 ( .A(n9993), .B(n9994), .Z(n9992) );
  XOR U9490 ( .A(n9991), .B(n9621), .Z(n9994) );
  XOR U9491 ( .A(n9995), .B(n9996), .Z(n9621) );
  AND U9492 ( .A(n467), .B(n9997), .Z(n9996) );
  XOR U9493 ( .A(n9998), .B(n9995), .Z(n9997) );
  XNOR U9494 ( .A(n9618), .B(n9991), .Z(n9993) );
  XOR U9495 ( .A(n9999), .B(n10000), .Z(n9618) );
  AND U9496 ( .A(n465), .B(n10001), .Z(n10000) );
  XOR U9497 ( .A(n10002), .B(n9999), .Z(n10001) );
  XOR U9498 ( .A(n10003), .B(n10004), .Z(n9991) );
  AND U9499 ( .A(n10005), .B(n10006), .Z(n10004) );
  XOR U9500 ( .A(n10003), .B(n9633), .Z(n10006) );
  XOR U9501 ( .A(n10007), .B(n10008), .Z(n9633) );
  AND U9502 ( .A(n467), .B(n10009), .Z(n10008) );
  XOR U9503 ( .A(n10010), .B(n10007), .Z(n10009) );
  XNOR U9504 ( .A(n9630), .B(n10003), .Z(n10005) );
  XOR U9505 ( .A(n10011), .B(n10012), .Z(n9630) );
  AND U9506 ( .A(n465), .B(n10013), .Z(n10012) );
  XOR U9507 ( .A(n10014), .B(n10011), .Z(n10013) );
  XOR U9508 ( .A(n10015), .B(n10016), .Z(n10003) );
  AND U9509 ( .A(n10017), .B(n10018), .Z(n10016) );
  XOR U9510 ( .A(n10015), .B(n9645), .Z(n10018) );
  XOR U9511 ( .A(n10019), .B(n10020), .Z(n9645) );
  AND U9512 ( .A(n467), .B(n10021), .Z(n10020) );
  XOR U9513 ( .A(n10022), .B(n10019), .Z(n10021) );
  XNOR U9514 ( .A(n9642), .B(n10015), .Z(n10017) );
  XOR U9515 ( .A(n10023), .B(n10024), .Z(n9642) );
  AND U9516 ( .A(n465), .B(n10025), .Z(n10024) );
  XOR U9517 ( .A(n10026), .B(n10023), .Z(n10025) );
  XOR U9518 ( .A(n10027), .B(n10028), .Z(n10015) );
  AND U9519 ( .A(n10029), .B(n10030), .Z(n10028) );
  XOR U9520 ( .A(n10027), .B(n9657), .Z(n10030) );
  XOR U9521 ( .A(n10031), .B(n10032), .Z(n9657) );
  AND U9522 ( .A(n467), .B(n10033), .Z(n10032) );
  XOR U9523 ( .A(n10034), .B(n10031), .Z(n10033) );
  XNOR U9524 ( .A(n9654), .B(n10027), .Z(n10029) );
  XOR U9525 ( .A(n10035), .B(n10036), .Z(n9654) );
  AND U9526 ( .A(n465), .B(n10037), .Z(n10036) );
  XOR U9527 ( .A(n10038), .B(n10035), .Z(n10037) );
  XOR U9528 ( .A(n10039), .B(n10040), .Z(n10027) );
  AND U9529 ( .A(n10041), .B(n10042), .Z(n10040) );
  XOR U9530 ( .A(n10039), .B(n9669), .Z(n10042) );
  XOR U9531 ( .A(n10043), .B(n10044), .Z(n9669) );
  AND U9532 ( .A(n467), .B(n10045), .Z(n10044) );
  XOR U9533 ( .A(n10046), .B(n10043), .Z(n10045) );
  XNOR U9534 ( .A(n9666), .B(n10039), .Z(n10041) );
  XOR U9535 ( .A(n10047), .B(n10048), .Z(n9666) );
  AND U9536 ( .A(n465), .B(n10049), .Z(n10048) );
  XOR U9537 ( .A(n10050), .B(n10047), .Z(n10049) );
  XOR U9538 ( .A(n10051), .B(n10052), .Z(n10039) );
  AND U9539 ( .A(n10053), .B(n10054), .Z(n10052) );
  XOR U9540 ( .A(n10051), .B(n9681), .Z(n10054) );
  XOR U9541 ( .A(n10055), .B(n10056), .Z(n9681) );
  AND U9542 ( .A(n467), .B(n10057), .Z(n10056) );
  XOR U9543 ( .A(n10058), .B(n10055), .Z(n10057) );
  XNOR U9544 ( .A(n9678), .B(n10051), .Z(n10053) );
  XOR U9545 ( .A(n10059), .B(n10060), .Z(n9678) );
  AND U9546 ( .A(n465), .B(n10061), .Z(n10060) );
  XOR U9547 ( .A(n10062), .B(n10059), .Z(n10061) );
  XOR U9548 ( .A(n10063), .B(n10064), .Z(n10051) );
  AND U9549 ( .A(n10065), .B(n10066), .Z(n10064) );
  XOR U9550 ( .A(n10063), .B(n9693), .Z(n10066) );
  XOR U9551 ( .A(n10067), .B(n10068), .Z(n9693) );
  AND U9552 ( .A(n467), .B(n10069), .Z(n10068) );
  XOR U9553 ( .A(n10070), .B(n10067), .Z(n10069) );
  XNOR U9554 ( .A(n9690), .B(n10063), .Z(n10065) );
  XOR U9555 ( .A(n10071), .B(n10072), .Z(n9690) );
  AND U9556 ( .A(n465), .B(n10073), .Z(n10072) );
  XOR U9557 ( .A(n10074), .B(n10071), .Z(n10073) );
  XOR U9558 ( .A(n10075), .B(n10076), .Z(n10063) );
  AND U9559 ( .A(n10077), .B(n10078), .Z(n10076) );
  XOR U9560 ( .A(n10075), .B(n9705), .Z(n10078) );
  XOR U9561 ( .A(n10079), .B(n10080), .Z(n9705) );
  AND U9562 ( .A(n467), .B(n10081), .Z(n10080) );
  XOR U9563 ( .A(n10082), .B(n10079), .Z(n10081) );
  XNOR U9564 ( .A(n9702), .B(n10075), .Z(n10077) );
  XOR U9565 ( .A(n10083), .B(n10084), .Z(n9702) );
  AND U9566 ( .A(n465), .B(n10085), .Z(n10084) );
  XOR U9567 ( .A(n10086), .B(n10083), .Z(n10085) );
  XOR U9568 ( .A(n10087), .B(n10088), .Z(n10075) );
  AND U9569 ( .A(n10089), .B(n10090), .Z(n10088) );
  XOR U9570 ( .A(n10087), .B(n9717), .Z(n10090) );
  XOR U9571 ( .A(n10091), .B(n10092), .Z(n9717) );
  AND U9572 ( .A(n467), .B(n10093), .Z(n10092) );
  XOR U9573 ( .A(n10094), .B(n10091), .Z(n10093) );
  XNOR U9574 ( .A(n9714), .B(n10087), .Z(n10089) );
  XOR U9575 ( .A(n10095), .B(n10096), .Z(n9714) );
  AND U9576 ( .A(n465), .B(n10097), .Z(n10096) );
  XOR U9577 ( .A(n10098), .B(n10095), .Z(n10097) );
  XOR U9578 ( .A(n10099), .B(n10100), .Z(n10087) );
  AND U9579 ( .A(n10101), .B(n10102), .Z(n10100) );
  XOR U9580 ( .A(n10099), .B(n9729), .Z(n10102) );
  XOR U9581 ( .A(n10103), .B(n10104), .Z(n9729) );
  AND U9582 ( .A(n467), .B(n10105), .Z(n10104) );
  XOR U9583 ( .A(n10106), .B(n10103), .Z(n10105) );
  XNOR U9584 ( .A(n9726), .B(n10099), .Z(n10101) );
  XOR U9585 ( .A(n10107), .B(n10108), .Z(n9726) );
  AND U9586 ( .A(n465), .B(n10109), .Z(n10108) );
  XOR U9587 ( .A(n10110), .B(n10107), .Z(n10109) );
  XOR U9588 ( .A(n10111), .B(n10112), .Z(n10099) );
  AND U9589 ( .A(n10113), .B(n10114), .Z(n10112) );
  XOR U9590 ( .A(n10111), .B(n9741), .Z(n10114) );
  XOR U9591 ( .A(n10115), .B(n10116), .Z(n9741) );
  AND U9592 ( .A(n467), .B(n10117), .Z(n10116) );
  XOR U9593 ( .A(n10118), .B(n10115), .Z(n10117) );
  XNOR U9594 ( .A(n9738), .B(n10111), .Z(n10113) );
  XOR U9595 ( .A(n10119), .B(n10120), .Z(n9738) );
  AND U9596 ( .A(n465), .B(n10121), .Z(n10120) );
  XOR U9597 ( .A(n10122), .B(n10119), .Z(n10121) );
  XOR U9598 ( .A(n10123), .B(n10124), .Z(n10111) );
  AND U9599 ( .A(n10125), .B(n10126), .Z(n10124) );
  XOR U9600 ( .A(n10123), .B(n9753), .Z(n10126) );
  XOR U9601 ( .A(n10127), .B(n10128), .Z(n9753) );
  AND U9602 ( .A(n467), .B(n10129), .Z(n10128) );
  XOR U9603 ( .A(n10130), .B(n10127), .Z(n10129) );
  XNOR U9604 ( .A(n9750), .B(n10123), .Z(n10125) );
  XOR U9605 ( .A(n10131), .B(n10132), .Z(n9750) );
  AND U9606 ( .A(n465), .B(n10133), .Z(n10132) );
  XOR U9607 ( .A(n10134), .B(n10131), .Z(n10133) );
  XOR U9608 ( .A(n10135), .B(n10136), .Z(n10123) );
  AND U9609 ( .A(n10137), .B(n10138), .Z(n10136) );
  XOR U9610 ( .A(n10135), .B(n9765), .Z(n10138) );
  XOR U9611 ( .A(n10139), .B(n10140), .Z(n9765) );
  AND U9612 ( .A(n467), .B(n10141), .Z(n10140) );
  XOR U9613 ( .A(n10142), .B(n10139), .Z(n10141) );
  XNOR U9614 ( .A(n9762), .B(n10135), .Z(n10137) );
  XOR U9615 ( .A(n10143), .B(n10144), .Z(n9762) );
  AND U9616 ( .A(n465), .B(n10145), .Z(n10144) );
  XOR U9617 ( .A(n10146), .B(n10143), .Z(n10145) );
  XOR U9618 ( .A(n10147), .B(n10148), .Z(n10135) );
  AND U9619 ( .A(n10149), .B(n10150), .Z(n10148) );
  XOR U9620 ( .A(n10147), .B(n9777), .Z(n10150) );
  XOR U9621 ( .A(n10151), .B(n10152), .Z(n9777) );
  AND U9622 ( .A(n467), .B(n10153), .Z(n10152) );
  XOR U9623 ( .A(n10154), .B(n10151), .Z(n10153) );
  XNOR U9624 ( .A(n9774), .B(n10147), .Z(n10149) );
  XOR U9625 ( .A(n10155), .B(n10156), .Z(n9774) );
  AND U9626 ( .A(n465), .B(n10157), .Z(n10156) );
  XOR U9627 ( .A(n10158), .B(n10155), .Z(n10157) );
  XOR U9628 ( .A(n10159), .B(n10160), .Z(n10147) );
  AND U9629 ( .A(n10161), .B(n10162), .Z(n10160) );
  XOR U9630 ( .A(n10159), .B(n9789), .Z(n10162) );
  XOR U9631 ( .A(n10163), .B(n10164), .Z(n9789) );
  AND U9632 ( .A(n467), .B(n10165), .Z(n10164) );
  XOR U9633 ( .A(n10166), .B(n10163), .Z(n10165) );
  XNOR U9634 ( .A(n9786), .B(n10159), .Z(n10161) );
  XOR U9635 ( .A(n10167), .B(n10168), .Z(n9786) );
  AND U9636 ( .A(n465), .B(n10169), .Z(n10168) );
  XOR U9637 ( .A(n10170), .B(n10167), .Z(n10169) );
  XOR U9638 ( .A(n10171), .B(n10172), .Z(n10159) );
  AND U9639 ( .A(n10173), .B(n10174), .Z(n10172) );
  XOR U9640 ( .A(n10171), .B(n9801), .Z(n10174) );
  XOR U9641 ( .A(n10175), .B(n10176), .Z(n9801) );
  AND U9642 ( .A(n467), .B(n10177), .Z(n10176) );
  XOR U9643 ( .A(n10178), .B(n10175), .Z(n10177) );
  XNOR U9644 ( .A(n9798), .B(n10171), .Z(n10173) );
  XOR U9645 ( .A(n10179), .B(n10180), .Z(n9798) );
  AND U9646 ( .A(n465), .B(n10181), .Z(n10180) );
  XOR U9647 ( .A(n10182), .B(n10179), .Z(n10181) );
  XOR U9648 ( .A(n10183), .B(n10184), .Z(n10171) );
  AND U9649 ( .A(n10185), .B(n10186), .Z(n10184) );
  XOR U9650 ( .A(n10183), .B(n9813), .Z(n10186) );
  XOR U9651 ( .A(n10187), .B(n10188), .Z(n9813) );
  AND U9652 ( .A(n467), .B(n10189), .Z(n10188) );
  XOR U9653 ( .A(n10190), .B(n10187), .Z(n10189) );
  XNOR U9654 ( .A(n9810), .B(n10183), .Z(n10185) );
  XOR U9655 ( .A(n10191), .B(n10192), .Z(n9810) );
  AND U9656 ( .A(n465), .B(n10193), .Z(n10192) );
  XOR U9657 ( .A(n10194), .B(n10191), .Z(n10193) );
  XOR U9658 ( .A(n10195), .B(n10196), .Z(n10183) );
  AND U9659 ( .A(n10197), .B(n10198), .Z(n10196) );
  XOR U9660 ( .A(n10195), .B(n9825), .Z(n10198) );
  XOR U9661 ( .A(n10199), .B(n10200), .Z(n9825) );
  AND U9662 ( .A(n467), .B(n10201), .Z(n10200) );
  XOR U9663 ( .A(n10202), .B(n10199), .Z(n10201) );
  XNOR U9664 ( .A(n9822), .B(n10195), .Z(n10197) );
  XOR U9665 ( .A(n10203), .B(n10204), .Z(n9822) );
  AND U9666 ( .A(n465), .B(n10205), .Z(n10204) );
  XOR U9667 ( .A(n10206), .B(n10203), .Z(n10205) );
  XOR U9668 ( .A(n10207), .B(n10208), .Z(n10195) );
  AND U9669 ( .A(n10209), .B(n10210), .Z(n10208) );
  XOR U9670 ( .A(n10207), .B(n9837), .Z(n10210) );
  XOR U9671 ( .A(n10211), .B(n10212), .Z(n9837) );
  AND U9672 ( .A(n467), .B(n10213), .Z(n10212) );
  XOR U9673 ( .A(n10214), .B(n10211), .Z(n10213) );
  XNOR U9674 ( .A(n9834), .B(n10207), .Z(n10209) );
  XOR U9675 ( .A(n10215), .B(n10216), .Z(n9834) );
  AND U9676 ( .A(n465), .B(n10217), .Z(n10216) );
  XOR U9677 ( .A(n10218), .B(n10215), .Z(n10217) );
  XOR U9678 ( .A(n10219), .B(n10220), .Z(n10207) );
  AND U9679 ( .A(n10221), .B(n10222), .Z(n10220) );
  XOR U9680 ( .A(n10219), .B(n9849), .Z(n10222) );
  XOR U9681 ( .A(n10223), .B(n10224), .Z(n9849) );
  AND U9682 ( .A(n467), .B(n10225), .Z(n10224) );
  XOR U9683 ( .A(n10226), .B(n10223), .Z(n10225) );
  XNOR U9684 ( .A(n9846), .B(n10219), .Z(n10221) );
  XOR U9685 ( .A(n10227), .B(n10228), .Z(n9846) );
  AND U9686 ( .A(n465), .B(n10229), .Z(n10228) );
  XOR U9687 ( .A(n10230), .B(n10227), .Z(n10229) );
  XOR U9688 ( .A(n10231), .B(n10232), .Z(n10219) );
  AND U9689 ( .A(n10233), .B(n10234), .Z(n10232) );
  XOR U9690 ( .A(n10231), .B(n9861), .Z(n10234) );
  XOR U9691 ( .A(n10235), .B(n10236), .Z(n9861) );
  AND U9692 ( .A(n467), .B(n10237), .Z(n10236) );
  XOR U9693 ( .A(n10238), .B(n10235), .Z(n10237) );
  XNOR U9694 ( .A(n9858), .B(n10231), .Z(n10233) );
  XOR U9695 ( .A(n10239), .B(n10240), .Z(n9858) );
  AND U9696 ( .A(n465), .B(n10241), .Z(n10240) );
  XOR U9697 ( .A(n10242), .B(n10239), .Z(n10241) );
  XOR U9698 ( .A(n10243), .B(n10244), .Z(n10231) );
  AND U9699 ( .A(n10245), .B(n10246), .Z(n10244) );
  XOR U9700 ( .A(n10243), .B(n9873), .Z(n10246) );
  XOR U9701 ( .A(n10247), .B(n10248), .Z(n9873) );
  AND U9702 ( .A(n467), .B(n10249), .Z(n10248) );
  XOR U9703 ( .A(n10250), .B(n10247), .Z(n10249) );
  XNOR U9704 ( .A(n9870), .B(n10243), .Z(n10245) );
  XOR U9705 ( .A(n10251), .B(n10252), .Z(n9870) );
  AND U9706 ( .A(n465), .B(n10253), .Z(n10252) );
  XOR U9707 ( .A(n10254), .B(n10251), .Z(n10253) );
  XOR U9708 ( .A(n10255), .B(n10256), .Z(n10243) );
  AND U9709 ( .A(n10257), .B(n10258), .Z(n10256) );
  XOR U9710 ( .A(n10255), .B(n9885), .Z(n10258) );
  XOR U9711 ( .A(n10259), .B(n10260), .Z(n9885) );
  AND U9712 ( .A(n467), .B(n10261), .Z(n10260) );
  XOR U9713 ( .A(n10262), .B(n10259), .Z(n10261) );
  XNOR U9714 ( .A(n9882), .B(n10255), .Z(n10257) );
  XOR U9715 ( .A(n10263), .B(n10264), .Z(n9882) );
  AND U9716 ( .A(n465), .B(n10265), .Z(n10264) );
  XOR U9717 ( .A(n10266), .B(n10263), .Z(n10265) );
  XOR U9718 ( .A(n10267), .B(n10268), .Z(n10255) );
  AND U9719 ( .A(n10269), .B(n10270), .Z(n10268) );
  XOR U9720 ( .A(n10267), .B(n9897), .Z(n10270) );
  XOR U9721 ( .A(n10271), .B(n10272), .Z(n9897) );
  AND U9722 ( .A(n467), .B(n10273), .Z(n10272) );
  XOR U9723 ( .A(n10274), .B(n10271), .Z(n10273) );
  XNOR U9724 ( .A(n9894), .B(n10267), .Z(n10269) );
  XOR U9725 ( .A(n10275), .B(n10276), .Z(n9894) );
  AND U9726 ( .A(n465), .B(n10277), .Z(n10276) );
  XOR U9727 ( .A(n10278), .B(n10275), .Z(n10277) );
  XOR U9728 ( .A(n10279), .B(n10280), .Z(n10267) );
  AND U9729 ( .A(n10281), .B(n10282), .Z(n10280) );
  XOR U9730 ( .A(n10279), .B(n9909), .Z(n10282) );
  XOR U9731 ( .A(n10283), .B(n10284), .Z(n9909) );
  AND U9732 ( .A(n467), .B(n10285), .Z(n10284) );
  XOR U9733 ( .A(n10286), .B(n10283), .Z(n10285) );
  XNOR U9734 ( .A(n9906), .B(n10279), .Z(n10281) );
  XOR U9735 ( .A(n10287), .B(n10288), .Z(n9906) );
  AND U9736 ( .A(n465), .B(n10289), .Z(n10288) );
  XOR U9737 ( .A(n10290), .B(n10287), .Z(n10289) );
  XOR U9738 ( .A(n10291), .B(n10292), .Z(n10279) );
  AND U9739 ( .A(n10293), .B(n10294), .Z(n10292) );
  XOR U9740 ( .A(n10291), .B(n9921), .Z(n10294) );
  XOR U9741 ( .A(n10295), .B(n10296), .Z(n9921) );
  AND U9742 ( .A(n467), .B(n10297), .Z(n10296) );
  XOR U9743 ( .A(n10298), .B(n10295), .Z(n10297) );
  XNOR U9744 ( .A(n9918), .B(n10291), .Z(n10293) );
  XOR U9745 ( .A(n10299), .B(n10300), .Z(n9918) );
  AND U9746 ( .A(n465), .B(n10301), .Z(n10300) );
  XOR U9747 ( .A(n10302), .B(n10299), .Z(n10301) );
  XOR U9748 ( .A(n10303), .B(n10304), .Z(n10291) );
  AND U9749 ( .A(n10305), .B(n10306), .Z(n10304) );
  XNOR U9750 ( .A(n10307), .B(n9934), .Z(n10306) );
  XOR U9751 ( .A(n10308), .B(n10309), .Z(n9934) );
  AND U9752 ( .A(n467), .B(n10310), .Z(n10309) );
  XOR U9753 ( .A(n10308), .B(n10311), .Z(n10310) );
  XNOR U9754 ( .A(n9931), .B(n10303), .Z(n10305) );
  XOR U9755 ( .A(n10312), .B(n10313), .Z(n9931) );
  AND U9756 ( .A(n465), .B(n10314), .Z(n10313) );
  XOR U9757 ( .A(n10312), .B(n10315), .Z(n10314) );
  IV U9758 ( .A(n10307), .Z(n10303) );
  AND U9759 ( .A(n9939), .B(n9942), .Z(n10307) );
  XNOR U9760 ( .A(n10316), .B(n10317), .Z(n9942) );
  AND U9761 ( .A(n467), .B(n10318), .Z(n10317) );
  XNOR U9762 ( .A(n10319), .B(n10316), .Z(n10318) );
  XOR U9763 ( .A(n10320), .B(n10321), .Z(n467) );
  AND U9764 ( .A(n10322), .B(n10323), .Z(n10321) );
  XOR U9765 ( .A(n9950), .B(n10320), .Z(n10323) );
  IV U9766 ( .A(n10324), .Z(n9950) );
  AND U9767 ( .A(p_input[7167]), .B(p_input[7135]), .Z(n10324) );
  XOR U9768 ( .A(n10320), .B(n9947), .Z(n10322) );
  AND U9769 ( .A(p_input[7071]), .B(p_input[7103]), .Z(n9947) );
  XOR U9770 ( .A(n10325), .B(n10326), .Z(n10320) );
  AND U9771 ( .A(n10327), .B(n10328), .Z(n10326) );
  XOR U9772 ( .A(n10325), .B(n9962), .Z(n10328) );
  XNOR U9773 ( .A(p_input[7134]), .B(n10329), .Z(n9962) );
  AND U9774 ( .A(n247), .B(n10330), .Z(n10329) );
  XOR U9775 ( .A(p_input[7166]), .B(p_input[7134]), .Z(n10330) );
  XNOR U9776 ( .A(n9959), .B(n10325), .Z(n10327) );
  XOR U9777 ( .A(n10331), .B(n10332), .Z(n9959) );
  AND U9778 ( .A(n245), .B(n10333), .Z(n10332) );
  XOR U9779 ( .A(p_input[7102]), .B(p_input[7070]), .Z(n10333) );
  XOR U9780 ( .A(n10334), .B(n10335), .Z(n10325) );
  AND U9781 ( .A(n10336), .B(n10337), .Z(n10335) );
  XOR U9782 ( .A(n10334), .B(n9974), .Z(n10337) );
  XNOR U9783 ( .A(p_input[7133]), .B(n10338), .Z(n9974) );
  AND U9784 ( .A(n247), .B(n10339), .Z(n10338) );
  XOR U9785 ( .A(p_input[7165]), .B(p_input[7133]), .Z(n10339) );
  XNOR U9786 ( .A(n9971), .B(n10334), .Z(n10336) );
  XOR U9787 ( .A(n10340), .B(n10341), .Z(n9971) );
  AND U9788 ( .A(n245), .B(n10342), .Z(n10341) );
  XOR U9789 ( .A(p_input[7101]), .B(p_input[7069]), .Z(n10342) );
  XOR U9790 ( .A(n10343), .B(n10344), .Z(n10334) );
  AND U9791 ( .A(n10345), .B(n10346), .Z(n10344) );
  XOR U9792 ( .A(n10343), .B(n9986), .Z(n10346) );
  XNOR U9793 ( .A(p_input[7132]), .B(n10347), .Z(n9986) );
  AND U9794 ( .A(n247), .B(n10348), .Z(n10347) );
  XOR U9795 ( .A(p_input[7164]), .B(p_input[7132]), .Z(n10348) );
  XNOR U9796 ( .A(n9983), .B(n10343), .Z(n10345) );
  XOR U9797 ( .A(n10349), .B(n10350), .Z(n9983) );
  AND U9798 ( .A(n245), .B(n10351), .Z(n10350) );
  XOR U9799 ( .A(p_input[7100]), .B(p_input[7068]), .Z(n10351) );
  XOR U9800 ( .A(n10352), .B(n10353), .Z(n10343) );
  AND U9801 ( .A(n10354), .B(n10355), .Z(n10353) );
  XOR U9802 ( .A(n10352), .B(n9998), .Z(n10355) );
  XNOR U9803 ( .A(p_input[7131]), .B(n10356), .Z(n9998) );
  AND U9804 ( .A(n247), .B(n10357), .Z(n10356) );
  XOR U9805 ( .A(p_input[7163]), .B(p_input[7131]), .Z(n10357) );
  XNOR U9806 ( .A(n9995), .B(n10352), .Z(n10354) );
  XOR U9807 ( .A(n10358), .B(n10359), .Z(n9995) );
  AND U9808 ( .A(n245), .B(n10360), .Z(n10359) );
  XOR U9809 ( .A(p_input[7099]), .B(p_input[7067]), .Z(n10360) );
  XOR U9810 ( .A(n10361), .B(n10362), .Z(n10352) );
  AND U9811 ( .A(n10363), .B(n10364), .Z(n10362) );
  XOR U9812 ( .A(n10361), .B(n10010), .Z(n10364) );
  XNOR U9813 ( .A(p_input[7130]), .B(n10365), .Z(n10010) );
  AND U9814 ( .A(n247), .B(n10366), .Z(n10365) );
  XOR U9815 ( .A(p_input[7162]), .B(p_input[7130]), .Z(n10366) );
  XNOR U9816 ( .A(n10007), .B(n10361), .Z(n10363) );
  XOR U9817 ( .A(n10367), .B(n10368), .Z(n10007) );
  AND U9818 ( .A(n245), .B(n10369), .Z(n10368) );
  XOR U9819 ( .A(p_input[7098]), .B(p_input[7066]), .Z(n10369) );
  XOR U9820 ( .A(n10370), .B(n10371), .Z(n10361) );
  AND U9821 ( .A(n10372), .B(n10373), .Z(n10371) );
  XOR U9822 ( .A(n10370), .B(n10022), .Z(n10373) );
  XNOR U9823 ( .A(p_input[7129]), .B(n10374), .Z(n10022) );
  AND U9824 ( .A(n247), .B(n10375), .Z(n10374) );
  XOR U9825 ( .A(p_input[7161]), .B(p_input[7129]), .Z(n10375) );
  XNOR U9826 ( .A(n10019), .B(n10370), .Z(n10372) );
  XOR U9827 ( .A(n10376), .B(n10377), .Z(n10019) );
  AND U9828 ( .A(n245), .B(n10378), .Z(n10377) );
  XOR U9829 ( .A(p_input[7097]), .B(p_input[7065]), .Z(n10378) );
  XOR U9830 ( .A(n10379), .B(n10380), .Z(n10370) );
  AND U9831 ( .A(n10381), .B(n10382), .Z(n10380) );
  XOR U9832 ( .A(n10379), .B(n10034), .Z(n10382) );
  XNOR U9833 ( .A(p_input[7128]), .B(n10383), .Z(n10034) );
  AND U9834 ( .A(n247), .B(n10384), .Z(n10383) );
  XOR U9835 ( .A(p_input[7160]), .B(p_input[7128]), .Z(n10384) );
  XNOR U9836 ( .A(n10031), .B(n10379), .Z(n10381) );
  XOR U9837 ( .A(n10385), .B(n10386), .Z(n10031) );
  AND U9838 ( .A(n245), .B(n10387), .Z(n10386) );
  XOR U9839 ( .A(p_input[7096]), .B(p_input[7064]), .Z(n10387) );
  XOR U9840 ( .A(n10388), .B(n10389), .Z(n10379) );
  AND U9841 ( .A(n10390), .B(n10391), .Z(n10389) );
  XOR U9842 ( .A(n10388), .B(n10046), .Z(n10391) );
  XNOR U9843 ( .A(p_input[7127]), .B(n10392), .Z(n10046) );
  AND U9844 ( .A(n247), .B(n10393), .Z(n10392) );
  XOR U9845 ( .A(p_input[7159]), .B(p_input[7127]), .Z(n10393) );
  XNOR U9846 ( .A(n10043), .B(n10388), .Z(n10390) );
  XOR U9847 ( .A(n10394), .B(n10395), .Z(n10043) );
  AND U9848 ( .A(n245), .B(n10396), .Z(n10395) );
  XOR U9849 ( .A(p_input[7095]), .B(p_input[7063]), .Z(n10396) );
  XOR U9850 ( .A(n10397), .B(n10398), .Z(n10388) );
  AND U9851 ( .A(n10399), .B(n10400), .Z(n10398) );
  XOR U9852 ( .A(n10397), .B(n10058), .Z(n10400) );
  XNOR U9853 ( .A(p_input[7126]), .B(n10401), .Z(n10058) );
  AND U9854 ( .A(n247), .B(n10402), .Z(n10401) );
  XOR U9855 ( .A(p_input[7158]), .B(p_input[7126]), .Z(n10402) );
  XNOR U9856 ( .A(n10055), .B(n10397), .Z(n10399) );
  XOR U9857 ( .A(n10403), .B(n10404), .Z(n10055) );
  AND U9858 ( .A(n245), .B(n10405), .Z(n10404) );
  XOR U9859 ( .A(p_input[7094]), .B(p_input[7062]), .Z(n10405) );
  XOR U9860 ( .A(n10406), .B(n10407), .Z(n10397) );
  AND U9861 ( .A(n10408), .B(n10409), .Z(n10407) );
  XOR U9862 ( .A(n10406), .B(n10070), .Z(n10409) );
  XNOR U9863 ( .A(p_input[7125]), .B(n10410), .Z(n10070) );
  AND U9864 ( .A(n247), .B(n10411), .Z(n10410) );
  XOR U9865 ( .A(p_input[7157]), .B(p_input[7125]), .Z(n10411) );
  XNOR U9866 ( .A(n10067), .B(n10406), .Z(n10408) );
  XOR U9867 ( .A(n10412), .B(n10413), .Z(n10067) );
  AND U9868 ( .A(n245), .B(n10414), .Z(n10413) );
  XOR U9869 ( .A(p_input[7093]), .B(p_input[7061]), .Z(n10414) );
  XOR U9870 ( .A(n10415), .B(n10416), .Z(n10406) );
  AND U9871 ( .A(n10417), .B(n10418), .Z(n10416) );
  XOR U9872 ( .A(n10415), .B(n10082), .Z(n10418) );
  XNOR U9873 ( .A(p_input[7124]), .B(n10419), .Z(n10082) );
  AND U9874 ( .A(n247), .B(n10420), .Z(n10419) );
  XOR U9875 ( .A(p_input[7156]), .B(p_input[7124]), .Z(n10420) );
  XNOR U9876 ( .A(n10079), .B(n10415), .Z(n10417) );
  XOR U9877 ( .A(n10421), .B(n10422), .Z(n10079) );
  AND U9878 ( .A(n245), .B(n10423), .Z(n10422) );
  XOR U9879 ( .A(p_input[7092]), .B(p_input[7060]), .Z(n10423) );
  XOR U9880 ( .A(n10424), .B(n10425), .Z(n10415) );
  AND U9881 ( .A(n10426), .B(n10427), .Z(n10425) );
  XOR U9882 ( .A(n10424), .B(n10094), .Z(n10427) );
  XNOR U9883 ( .A(p_input[7123]), .B(n10428), .Z(n10094) );
  AND U9884 ( .A(n247), .B(n10429), .Z(n10428) );
  XOR U9885 ( .A(p_input[7155]), .B(p_input[7123]), .Z(n10429) );
  XNOR U9886 ( .A(n10091), .B(n10424), .Z(n10426) );
  XOR U9887 ( .A(n10430), .B(n10431), .Z(n10091) );
  AND U9888 ( .A(n245), .B(n10432), .Z(n10431) );
  XOR U9889 ( .A(p_input[7091]), .B(p_input[7059]), .Z(n10432) );
  XOR U9890 ( .A(n10433), .B(n10434), .Z(n10424) );
  AND U9891 ( .A(n10435), .B(n10436), .Z(n10434) );
  XOR U9892 ( .A(n10433), .B(n10106), .Z(n10436) );
  XNOR U9893 ( .A(p_input[7122]), .B(n10437), .Z(n10106) );
  AND U9894 ( .A(n247), .B(n10438), .Z(n10437) );
  XOR U9895 ( .A(p_input[7154]), .B(p_input[7122]), .Z(n10438) );
  XNOR U9896 ( .A(n10103), .B(n10433), .Z(n10435) );
  XOR U9897 ( .A(n10439), .B(n10440), .Z(n10103) );
  AND U9898 ( .A(n245), .B(n10441), .Z(n10440) );
  XOR U9899 ( .A(p_input[7090]), .B(p_input[7058]), .Z(n10441) );
  XOR U9900 ( .A(n10442), .B(n10443), .Z(n10433) );
  AND U9901 ( .A(n10444), .B(n10445), .Z(n10443) );
  XOR U9902 ( .A(n10442), .B(n10118), .Z(n10445) );
  XNOR U9903 ( .A(p_input[7121]), .B(n10446), .Z(n10118) );
  AND U9904 ( .A(n247), .B(n10447), .Z(n10446) );
  XOR U9905 ( .A(p_input[7153]), .B(p_input[7121]), .Z(n10447) );
  XNOR U9906 ( .A(n10115), .B(n10442), .Z(n10444) );
  XOR U9907 ( .A(n10448), .B(n10449), .Z(n10115) );
  AND U9908 ( .A(n245), .B(n10450), .Z(n10449) );
  XOR U9909 ( .A(p_input[7089]), .B(p_input[7057]), .Z(n10450) );
  XOR U9910 ( .A(n10451), .B(n10452), .Z(n10442) );
  AND U9911 ( .A(n10453), .B(n10454), .Z(n10452) );
  XOR U9912 ( .A(n10451), .B(n10130), .Z(n10454) );
  XNOR U9913 ( .A(p_input[7120]), .B(n10455), .Z(n10130) );
  AND U9914 ( .A(n247), .B(n10456), .Z(n10455) );
  XOR U9915 ( .A(p_input[7152]), .B(p_input[7120]), .Z(n10456) );
  XNOR U9916 ( .A(n10127), .B(n10451), .Z(n10453) );
  XOR U9917 ( .A(n10457), .B(n10458), .Z(n10127) );
  AND U9918 ( .A(n245), .B(n10459), .Z(n10458) );
  XOR U9919 ( .A(p_input[7088]), .B(p_input[7056]), .Z(n10459) );
  XOR U9920 ( .A(n10460), .B(n10461), .Z(n10451) );
  AND U9921 ( .A(n10462), .B(n10463), .Z(n10461) );
  XOR U9922 ( .A(n10460), .B(n10142), .Z(n10463) );
  XNOR U9923 ( .A(p_input[7119]), .B(n10464), .Z(n10142) );
  AND U9924 ( .A(n247), .B(n10465), .Z(n10464) );
  XOR U9925 ( .A(p_input[7151]), .B(p_input[7119]), .Z(n10465) );
  XNOR U9926 ( .A(n10139), .B(n10460), .Z(n10462) );
  XOR U9927 ( .A(n10466), .B(n10467), .Z(n10139) );
  AND U9928 ( .A(n245), .B(n10468), .Z(n10467) );
  XOR U9929 ( .A(p_input[7087]), .B(p_input[7055]), .Z(n10468) );
  XOR U9930 ( .A(n10469), .B(n10470), .Z(n10460) );
  AND U9931 ( .A(n10471), .B(n10472), .Z(n10470) );
  XOR U9932 ( .A(n10469), .B(n10154), .Z(n10472) );
  XNOR U9933 ( .A(p_input[7118]), .B(n10473), .Z(n10154) );
  AND U9934 ( .A(n247), .B(n10474), .Z(n10473) );
  XOR U9935 ( .A(p_input[7150]), .B(p_input[7118]), .Z(n10474) );
  XNOR U9936 ( .A(n10151), .B(n10469), .Z(n10471) );
  XOR U9937 ( .A(n10475), .B(n10476), .Z(n10151) );
  AND U9938 ( .A(n245), .B(n10477), .Z(n10476) );
  XOR U9939 ( .A(p_input[7086]), .B(p_input[7054]), .Z(n10477) );
  XOR U9940 ( .A(n10478), .B(n10479), .Z(n10469) );
  AND U9941 ( .A(n10480), .B(n10481), .Z(n10479) );
  XOR U9942 ( .A(n10478), .B(n10166), .Z(n10481) );
  XNOR U9943 ( .A(p_input[7117]), .B(n10482), .Z(n10166) );
  AND U9944 ( .A(n247), .B(n10483), .Z(n10482) );
  XOR U9945 ( .A(p_input[7149]), .B(p_input[7117]), .Z(n10483) );
  XNOR U9946 ( .A(n10163), .B(n10478), .Z(n10480) );
  XOR U9947 ( .A(n10484), .B(n10485), .Z(n10163) );
  AND U9948 ( .A(n245), .B(n10486), .Z(n10485) );
  XOR U9949 ( .A(p_input[7085]), .B(p_input[7053]), .Z(n10486) );
  XOR U9950 ( .A(n10487), .B(n10488), .Z(n10478) );
  AND U9951 ( .A(n10489), .B(n10490), .Z(n10488) );
  XOR U9952 ( .A(n10487), .B(n10178), .Z(n10490) );
  XNOR U9953 ( .A(p_input[7116]), .B(n10491), .Z(n10178) );
  AND U9954 ( .A(n247), .B(n10492), .Z(n10491) );
  XOR U9955 ( .A(p_input[7148]), .B(p_input[7116]), .Z(n10492) );
  XNOR U9956 ( .A(n10175), .B(n10487), .Z(n10489) );
  XOR U9957 ( .A(n10493), .B(n10494), .Z(n10175) );
  AND U9958 ( .A(n245), .B(n10495), .Z(n10494) );
  XOR U9959 ( .A(p_input[7084]), .B(p_input[7052]), .Z(n10495) );
  XOR U9960 ( .A(n10496), .B(n10497), .Z(n10487) );
  AND U9961 ( .A(n10498), .B(n10499), .Z(n10497) );
  XOR U9962 ( .A(n10496), .B(n10190), .Z(n10499) );
  XNOR U9963 ( .A(p_input[7115]), .B(n10500), .Z(n10190) );
  AND U9964 ( .A(n247), .B(n10501), .Z(n10500) );
  XOR U9965 ( .A(p_input[7147]), .B(p_input[7115]), .Z(n10501) );
  XNOR U9966 ( .A(n10187), .B(n10496), .Z(n10498) );
  XOR U9967 ( .A(n10502), .B(n10503), .Z(n10187) );
  AND U9968 ( .A(n245), .B(n10504), .Z(n10503) );
  XOR U9969 ( .A(p_input[7083]), .B(p_input[7051]), .Z(n10504) );
  XOR U9970 ( .A(n10505), .B(n10506), .Z(n10496) );
  AND U9971 ( .A(n10507), .B(n10508), .Z(n10506) );
  XOR U9972 ( .A(n10505), .B(n10202), .Z(n10508) );
  XNOR U9973 ( .A(p_input[7114]), .B(n10509), .Z(n10202) );
  AND U9974 ( .A(n247), .B(n10510), .Z(n10509) );
  XOR U9975 ( .A(p_input[7146]), .B(p_input[7114]), .Z(n10510) );
  XNOR U9976 ( .A(n10199), .B(n10505), .Z(n10507) );
  XOR U9977 ( .A(n10511), .B(n10512), .Z(n10199) );
  AND U9978 ( .A(n245), .B(n10513), .Z(n10512) );
  XOR U9979 ( .A(p_input[7082]), .B(p_input[7050]), .Z(n10513) );
  XOR U9980 ( .A(n10514), .B(n10515), .Z(n10505) );
  AND U9981 ( .A(n10516), .B(n10517), .Z(n10515) );
  XOR U9982 ( .A(n10514), .B(n10214), .Z(n10517) );
  XNOR U9983 ( .A(p_input[7113]), .B(n10518), .Z(n10214) );
  AND U9984 ( .A(n247), .B(n10519), .Z(n10518) );
  XOR U9985 ( .A(p_input[7145]), .B(p_input[7113]), .Z(n10519) );
  XNOR U9986 ( .A(n10211), .B(n10514), .Z(n10516) );
  XOR U9987 ( .A(n10520), .B(n10521), .Z(n10211) );
  AND U9988 ( .A(n245), .B(n10522), .Z(n10521) );
  XOR U9989 ( .A(p_input[7081]), .B(p_input[7049]), .Z(n10522) );
  XOR U9990 ( .A(n10523), .B(n10524), .Z(n10514) );
  AND U9991 ( .A(n10525), .B(n10526), .Z(n10524) );
  XOR U9992 ( .A(n10523), .B(n10226), .Z(n10526) );
  XNOR U9993 ( .A(p_input[7112]), .B(n10527), .Z(n10226) );
  AND U9994 ( .A(n247), .B(n10528), .Z(n10527) );
  XOR U9995 ( .A(p_input[7144]), .B(p_input[7112]), .Z(n10528) );
  XNOR U9996 ( .A(n10223), .B(n10523), .Z(n10525) );
  XOR U9997 ( .A(n10529), .B(n10530), .Z(n10223) );
  AND U9998 ( .A(n245), .B(n10531), .Z(n10530) );
  XOR U9999 ( .A(p_input[7080]), .B(p_input[7048]), .Z(n10531) );
  XOR U10000 ( .A(n10532), .B(n10533), .Z(n10523) );
  AND U10001 ( .A(n10534), .B(n10535), .Z(n10533) );
  XOR U10002 ( .A(n10532), .B(n10238), .Z(n10535) );
  XNOR U10003 ( .A(p_input[7111]), .B(n10536), .Z(n10238) );
  AND U10004 ( .A(n247), .B(n10537), .Z(n10536) );
  XOR U10005 ( .A(p_input[7143]), .B(p_input[7111]), .Z(n10537) );
  XNOR U10006 ( .A(n10235), .B(n10532), .Z(n10534) );
  XOR U10007 ( .A(n10538), .B(n10539), .Z(n10235) );
  AND U10008 ( .A(n245), .B(n10540), .Z(n10539) );
  XOR U10009 ( .A(p_input[7079]), .B(p_input[7047]), .Z(n10540) );
  XOR U10010 ( .A(n10541), .B(n10542), .Z(n10532) );
  AND U10011 ( .A(n10543), .B(n10544), .Z(n10542) );
  XOR U10012 ( .A(n10541), .B(n10250), .Z(n10544) );
  XNOR U10013 ( .A(p_input[7110]), .B(n10545), .Z(n10250) );
  AND U10014 ( .A(n247), .B(n10546), .Z(n10545) );
  XOR U10015 ( .A(p_input[7142]), .B(p_input[7110]), .Z(n10546) );
  XNOR U10016 ( .A(n10247), .B(n10541), .Z(n10543) );
  XOR U10017 ( .A(n10547), .B(n10548), .Z(n10247) );
  AND U10018 ( .A(n245), .B(n10549), .Z(n10548) );
  XOR U10019 ( .A(p_input[7078]), .B(p_input[7046]), .Z(n10549) );
  XOR U10020 ( .A(n10550), .B(n10551), .Z(n10541) );
  AND U10021 ( .A(n10552), .B(n10553), .Z(n10551) );
  XOR U10022 ( .A(n10550), .B(n10262), .Z(n10553) );
  XNOR U10023 ( .A(p_input[7109]), .B(n10554), .Z(n10262) );
  AND U10024 ( .A(n247), .B(n10555), .Z(n10554) );
  XOR U10025 ( .A(p_input[7141]), .B(p_input[7109]), .Z(n10555) );
  XNOR U10026 ( .A(n10259), .B(n10550), .Z(n10552) );
  XOR U10027 ( .A(n10556), .B(n10557), .Z(n10259) );
  AND U10028 ( .A(n245), .B(n10558), .Z(n10557) );
  XOR U10029 ( .A(p_input[7077]), .B(p_input[7045]), .Z(n10558) );
  XOR U10030 ( .A(n10559), .B(n10560), .Z(n10550) );
  AND U10031 ( .A(n10561), .B(n10562), .Z(n10560) );
  XOR U10032 ( .A(n10559), .B(n10274), .Z(n10562) );
  XNOR U10033 ( .A(p_input[7108]), .B(n10563), .Z(n10274) );
  AND U10034 ( .A(n247), .B(n10564), .Z(n10563) );
  XOR U10035 ( .A(p_input[7140]), .B(p_input[7108]), .Z(n10564) );
  XNOR U10036 ( .A(n10271), .B(n10559), .Z(n10561) );
  XOR U10037 ( .A(n10565), .B(n10566), .Z(n10271) );
  AND U10038 ( .A(n245), .B(n10567), .Z(n10566) );
  XOR U10039 ( .A(p_input[7076]), .B(p_input[7044]), .Z(n10567) );
  XOR U10040 ( .A(n10568), .B(n10569), .Z(n10559) );
  AND U10041 ( .A(n10570), .B(n10571), .Z(n10569) );
  XOR U10042 ( .A(n10568), .B(n10286), .Z(n10571) );
  XNOR U10043 ( .A(p_input[7107]), .B(n10572), .Z(n10286) );
  AND U10044 ( .A(n247), .B(n10573), .Z(n10572) );
  XOR U10045 ( .A(p_input[7139]), .B(p_input[7107]), .Z(n10573) );
  XNOR U10046 ( .A(n10283), .B(n10568), .Z(n10570) );
  XOR U10047 ( .A(n10574), .B(n10575), .Z(n10283) );
  AND U10048 ( .A(n245), .B(n10576), .Z(n10575) );
  XOR U10049 ( .A(p_input[7075]), .B(p_input[7043]), .Z(n10576) );
  XOR U10050 ( .A(n10577), .B(n10578), .Z(n10568) );
  AND U10051 ( .A(n10579), .B(n10580), .Z(n10578) );
  XOR U10052 ( .A(n10577), .B(n10298), .Z(n10580) );
  XNOR U10053 ( .A(p_input[7106]), .B(n10581), .Z(n10298) );
  AND U10054 ( .A(n247), .B(n10582), .Z(n10581) );
  XOR U10055 ( .A(p_input[7138]), .B(p_input[7106]), .Z(n10582) );
  XNOR U10056 ( .A(n10295), .B(n10577), .Z(n10579) );
  XOR U10057 ( .A(n10583), .B(n10584), .Z(n10295) );
  AND U10058 ( .A(n245), .B(n10585), .Z(n10584) );
  XOR U10059 ( .A(p_input[7074]), .B(p_input[7042]), .Z(n10585) );
  XOR U10060 ( .A(n10586), .B(n10587), .Z(n10577) );
  AND U10061 ( .A(n10588), .B(n10589), .Z(n10587) );
  XNOR U10062 ( .A(n10590), .B(n10311), .Z(n10589) );
  XNOR U10063 ( .A(p_input[7105]), .B(n10591), .Z(n10311) );
  AND U10064 ( .A(n247), .B(n10592), .Z(n10591) );
  XNOR U10065 ( .A(p_input[7137]), .B(n10593), .Z(n10592) );
  IV U10066 ( .A(p_input[7105]), .Z(n10593) );
  XNOR U10067 ( .A(n10308), .B(n10586), .Z(n10588) );
  XNOR U10068 ( .A(p_input[7041]), .B(n10594), .Z(n10308) );
  AND U10069 ( .A(n245), .B(n10595), .Z(n10594) );
  XOR U10070 ( .A(p_input[7073]), .B(p_input[7041]), .Z(n10595) );
  IV U10071 ( .A(n10590), .Z(n10586) );
  AND U10072 ( .A(n10316), .B(n10319), .Z(n10590) );
  XOR U10073 ( .A(p_input[7104]), .B(n10596), .Z(n10319) );
  AND U10074 ( .A(n247), .B(n10597), .Z(n10596) );
  XOR U10075 ( .A(p_input[7136]), .B(p_input[7104]), .Z(n10597) );
  XOR U10076 ( .A(n10598), .B(n10599), .Z(n247) );
  AND U10077 ( .A(n10600), .B(n10601), .Z(n10599) );
  XNOR U10078 ( .A(p_input[7167]), .B(n10598), .Z(n10601) );
  XOR U10079 ( .A(n10598), .B(p_input[7135]), .Z(n10600) );
  XOR U10080 ( .A(n10602), .B(n10603), .Z(n10598) );
  AND U10081 ( .A(n10604), .B(n10605), .Z(n10603) );
  XNOR U10082 ( .A(p_input[7166]), .B(n10602), .Z(n10605) );
  XOR U10083 ( .A(n10602), .B(p_input[7134]), .Z(n10604) );
  XOR U10084 ( .A(n10606), .B(n10607), .Z(n10602) );
  AND U10085 ( .A(n10608), .B(n10609), .Z(n10607) );
  XNOR U10086 ( .A(p_input[7165]), .B(n10606), .Z(n10609) );
  XOR U10087 ( .A(n10606), .B(p_input[7133]), .Z(n10608) );
  XOR U10088 ( .A(n10610), .B(n10611), .Z(n10606) );
  AND U10089 ( .A(n10612), .B(n10613), .Z(n10611) );
  XNOR U10090 ( .A(p_input[7164]), .B(n10610), .Z(n10613) );
  XOR U10091 ( .A(n10610), .B(p_input[7132]), .Z(n10612) );
  XOR U10092 ( .A(n10614), .B(n10615), .Z(n10610) );
  AND U10093 ( .A(n10616), .B(n10617), .Z(n10615) );
  XNOR U10094 ( .A(p_input[7163]), .B(n10614), .Z(n10617) );
  XOR U10095 ( .A(n10614), .B(p_input[7131]), .Z(n10616) );
  XOR U10096 ( .A(n10618), .B(n10619), .Z(n10614) );
  AND U10097 ( .A(n10620), .B(n10621), .Z(n10619) );
  XNOR U10098 ( .A(p_input[7162]), .B(n10618), .Z(n10621) );
  XOR U10099 ( .A(n10618), .B(p_input[7130]), .Z(n10620) );
  XOR U10100 ( .A(n10622), .B(n10623), .Z(n10618) );
  AND U10101 ( .A(n10624), .B(n10625), .Z(n10623) );
  XNOR U10102 ( .A(p_input[7161]), .B(n10622), .Z(n10625) );
  XOR U10103 ( .A(n10622), .B(p_input[7129]), .Z(n10624) );
  XOR U10104 ( .A(n10626), .B(n10627), .Z(n10622) );
  AND U10105 ( .A(n10628), .B(n10629), .Z(n10627) );
  XNOR U10106 ( .A(p_input[7160]), .B(n10626), .Z(n10629) );
  XOR U10107 ( .A(n10626), .B(p_input[7128]), .Z(n10628) );
  XOR U10108 ( .A(n10630), .B(n10631), .Z(n10626) );
  AND U10109 ( .A(n10632), .B(n10633), .Z(n10631) );
  XNOR U10110 ( .A(p_input[7159]), .B(n10630), .Z(n10633) );
  XOR U10111 ( .A(n10630), .B(p_input[7127]), .Z(n10632) );
  XOR U10112 ( .A(n10634), .B(n10635), .Z(n10630) );
  AND U10113 ( .A(n10636), .B(n10637), .Z(n10635) );
  XNOR U10114 ( .A(p_input[7158]), .B(n10634), .Z(n10637) );
  XOR U10115 ( .A(n10634), .B(p_input[7126]), .Z(n10636) );
  XOR U10116 ( .A(n10638), .B(n10639), .Z(n10634) );
  AND U10117 ( .A(n10640), .B(n10641), .Z(n10639) );
  XNOR U10118 ( .A(p_input[7157]), .B(n10638), .Z(n10641) );
  XOR U10119 ( .A(n10638), .B(p_input[7125]), .Z(n10640) );
  XOR U10120 ( .A(n10642), .B(n10643), .Z(n10638) );
  AND U10121 ( .A(n10644), .B(n10645), .Z(n10643) );
  XNOR U10122 ( .A(p_input[7156]), .B(n10642), .Z(n10645) );
  XOR U10123 ( .A(n10642), .B(p_input[7124]), .Z(n10644) );
  XOR U10124 ( .A(n10646), .B(n10647), .Z(n10642) );
  AND U10125 ( .A(n10648), .B(n10649), .Z(n10647) );
  XNOR U10126 ( .A(p_input[7155]), .B(n10646), .Z(n10649) );
  XOR U10127 ( .A(n10646), .B(p_input[7123]), .Z(n10648) );
  XOR U10128 ( .A(n10650), .B(n10651), .Z(n10646) );
  AND U10129 ( .A(n10652), .B(n10653), .Z(n10651) );
  XNOR U10130 ( .A(p_input[7154]), .B(n10650), .Z(n10653) );
  XOR U10131 ( .A(n10650), .B(p_input[7122]), .Z(n10652) );
  XOR U10132 ( .A(n10654), .B(n10655), .Z(n10650) );
  AND U10133 ( .A(n10656), .B(n10657), .Z(n10655) );
  XNOR U10134 ( .A(p_input[7153]), .B(n10654), .Z(n10657) );
  XOR U10135 ( .A(n10654), .B(p_input[7121]), .Z(n10656) );
  XOR U10136 ( .A(n10658), .B(n10659), .Z(n10654) );
  AND U10137 ( .A(n10660), .B(n10661), .Z(n10659) );
  XNOR U10138 ( .A(p_input[7152]), .B(n10658), .Z(n10661) );
  XOR U10139 ( .A(n10658), .B(p_input[7120]), .Z(n10660) );
  XOR U10140 ( .A(n10662), .B(n10663), .Z(n10658) );
  AND U10141 ( .A(n10664), .B(n10665), .Z(n10663) );
  XNOR U10142 ( .A(p_input[7151]), .B(n10662), .Z(n10665) );
  XOR U10143 ( .A(n10662), .B(p_input[7119]), .Z(n10664) );
  XOR U10144 ( .A(n10666), .B(n10667), .Z(n10662) );
  AND U10145 ( .A(n10668), .B(n10669), .Z(n10667) );
  XNOR U10146 ( .A(p_input[7150]), .B(n10666), .Z(n10669) );
  XOR U10147 ( .A(n10666), .B(p_input[7118]), .Z(n10668) );
  XOR U10148 ( .A(n10670), .B(n10671), .Z(n10666) );
  AND U10149 ( .A(n10672), .B(n10673), .Z(n10671) );
  XNOR U10150 ( .A(p_input[7149]), .B(n10670), .Z(n10673) );
  XOR U10151 ( .A(n10670), .B(p_input[7117]), .Z(n10672) );
  XOR U10152 ( .A(n10674), .B(n10675), .Z(n10670) );
  AND U10153 ( .A(n10676), .B(n10677), .Z(n10675) );
  XNOR U10154 ( .A(p_input[7148]), .B(n10674), .Z(n10677) );
  XOR U10155 ( .A(n10674), .B(p_input[7116]), .Z(n10676) );
  XOR U10156 ( .A(n10678), .B(n10679), .Z(n10674) );
  AND U10157 ( .A(n10680), .B(n10681), .Z(n10679) );
  XNOR U10158 ( .A(p_input[7147]), .B(n10678), .Z(n10681) );
  XOR U10159 ( .A(n10678), .B(p_input[7115]), .Z(n10680) );
  XOR U10160 ( .A(n10682), .B(n10683), .Z(n10678) );
  AND U10161 ( .A(n10684), .B(n10685), .Z(n10683) );
  XNOR U10162 ( .A(p_input[7146]), .B(n10682), .Z(n10685) );
  XOR U10163 ( .A(n10682), .B(p_input[7114]), .Z(n10684) );
  XOR U10164 ( .A(n10686), .B(n10687), .Z(n10682) );
  AND U10165 ( .A(n10688), .B(n10689), .Z(n10687) );
  XNOR U10166 ( .A(p_input[7145]), .B(n10686), .Z(n10689) );
  XOR U10167 ( .A(n10686), .B(p_input[7113]), .Z(n10688) );
  XOR U10168 ( .A(n10690), .B(n10691), .Z(n10686) );
  AND U10169 ( .A(n10692), .B(n10693), .Z(n10691) );
  XNOR U10170 ( .A(p_input[7144]), .B(n10690), .Z(n10693) );
  XOR U10171 ( .A(n10690), .B(p_input[7112]), .Z(n10692) );
  XOR U10172 ( .A(n10694), .B(n10695), .Z(n10690) );
  AND U10173 ( .A(n10696), .B(n10697), .Z(n10695) );
  XNOR U10174 ( .A(p_input[7143]), .B(n10694), .Z(n10697) );
  XOR U10175 ( .A(n10694), .B(p_input[7111]), .Z(n10696) );
  XOR U10176 ( .A(n10698), .B(n10699), .Z(n10694) );
  AND U10177 ( .A(n10700), .B(n10701), .Z(n10699) );
  XNOR U10178 ( .A(p_input[7142]), .B(n10698), .Z(n10701) );
  XOR U10179 ( .A(n10698), .B(p_input[7110]), .Z(n10700) );
  XOR U10180 ( .A(n10702), .B(n10703), .Z(n10698) );
  AND U10181 ( .A(n10704), .B(n10705), .Z(n10703) );
  XNOR U10182 ( .A(p_input[7141]), .B(n10702), .Z(n10705) );
  XOR U10183 ( .A(n10702), .B(p_input[7109]), .Z(n10704) );
  XOR U10184 ( .A(n10706), .B(n10707), .Z(n10702) );
  AND U10185 ( .A(n10708), .B(n10709), .Z(n10707) );
  XNOR U10186 ( .A(p_input[7140]), .B(n10706), .Z(n10709) );
  XOR U10187 ( .A(n10706), .B(p_input[7108]), .Z(n10708) );
  XOR U10188 ( .A(n10710), .B(n10711), .Z(n10706) );
  AND U10189 ( .A(n10712), .B(n10713), .Z(n10711) );
  XNOR U10190 ( .A(p_input[7139]), .B(n10710), .Z(n10713) );
  XOR U10191 ( .A(n10710), .B(p_input[7107]), .Z(n10712) );
  XOR U10192 ( .A(n10714), .B(n10715), .Z(n10710) );
  AND U10193 ( .A(n10716), .B(n10717), .Z(n10715) );
  XNOR U10194 ( .A(p_input[7138]), .B(n10714), .Z(n10717) );
  XOR U10195 ( .A(n10714), .B(p_input[7106]), .Z(n10716) );
  XNOR U10196 ( .A(n10718), .B(n10719), .Z(n10714) );
  AND U10197 ( .A(n10720), .B(n10721), .Z(n10719) );
  XOR U10198 ( .A(p_input[7137]), .B(n10718), .Z(n10721) );
  XNOR U10199 ( .A(p_input[7105]), .B(n10718), .Z(n10720) );
  AND U10200 ( .A(p_input[7136]), .B(n10722), .Z(n10718) );
  IV U10201 ( .A(p_input[7104]), .Z(n10722) );
  XNOR U10202 ( .A(p_input[7040]), .B(n10723), .Z(n10316) );
  AND U10203 ( .A(n245), .B(n10724), .Z(n10723) );
  XOR U10204 ( .A(p_input[7072]), .B(p_input[7040]), .Z(n10724) );
  XOR U10205 ( .A(n10725), .B(n10726), .Z(n245) );
  AND U10206 ( .A(n10727), .B(n10728), .Z(n10726) );
  XNOR U10207 ( .A(p_input[7103]), .B(n10725), .Z(n10728) );
  XOR U10208 ( .A(n10725), .B(p_input[7071]), .Z(n10727) );
  XOR U10209 ( .A(n10729), .B(n10730), .Z(n10725) );
  AND U10210 ( .A(n10731), .B(n10732), .Z(n10730) );
  XNOR U10211 ( .A(p_input[7102]), .B(n10729), .Z(n10732) );
  XNOR U10212 ( .A(n10729), .B(n10331), .Z(n10731) );
  IV U10213 ( .A(p_input[7070]), .Z(n10331) );
  XOR U10214 ( .A(n10733), .B(n10734), .Z(n10729) );
  AND U10215 ( .A(n10735), .B(n10736), .Z(n10734) );
  XNOR U10216 ( .A(p_input[7101]), .B(n10733), .Z(n10736) );
  XNOR U10217 ( .A(n10733), .B(n10340), .Z(n10735) );
  IV U10218 ( .A(p_input[7069]), .Z(n10340) );
  XOR U10219 ( .A(n10737), .B(n10738), .Z(n10733) );
  AND U10220 ( .A(n10739), .B(n10740), .Z(n10738) );
  XNOR U10221 ( .A(p_input[7100]), .B(n10737), .Z(n10740) );
  XNOR U10222 ( .A(n10737), .B(n10349), .Z(n10739) );
  IV U10223 ( .A(p_input[7068]), .Z(n10349) );
  XOR U10224 ( .A(n10741), .B(n10742), .Z(n10737) );
  AND U10225 ( .A(n10743), .B(n10744), .Z(n10742) );
  XNOR U10226 ( .A(p_input[7099]), .B(n10741), .Z(n10744) );
  XNOR U10227 ( .A(n10741), .B(n10358), .Z(n10743) );
  IV U10228 ( .A(p_input[7067]), .Z(n10358) );
  XOR U10229 ( .A(n10745), .B(n10746), .Z(n10741) );
  AND U10230 ( .A(n10747), .B(n10748), .Z(n10746) );
  XNOR U10231 ( .A(p_input[7098]), .B(n10745), .Z(n10748) );
  XNOR U10232 ( .A(n10745), .B(n10367), .Z(n10747) );
  IV U10233 ( .A(p_input[7066]), .Z(n10367) );
  XOR U10234 ( .A(n10749), .B(n10750), .Z(n10745) );
  AND U10235 ( .A(n10751), .B(n10752), .Z(n10750) );
  XNOR U10236 ( .A(p_input[7097]), .B(n10749), .Z(n10752) );
  XNOR U10237 ( .A(n10749), .B(n10376), .Z(n10751) );
  IV U10238 ( .A(p_input[7065]), .Z(n10376) );
  XOR U10239 ( .A(n10753), .B(n10754), .Z(n10749) );
  AND U10240 ( .A(n10755), .B(n10756), .Z(n10754) );
  XNOR U10241 ( .A(p_input[7096]), .B(n10753), .Z(n10756) );
  XNOR U10242 ( .A(n10753), .B(n10385), .Z(n10755) );
  IV U10243 ( .A(p_input[7064]), .Z(n10385) );
  XOR U10244 ( .A(n10757), .B(n10758), .Z(n10753) );
  AND U10245 ( .A(n10759), .B(n10760), .Z(n10758) );
  XNOR U10246 ( .A(p_input[7095]), .B(n10757), .Z(n10760) );
  XNOR U10247 ( .A(n10757), .B(n10394), .Z(n10759) );
  IV U10248 ( .A(p_input[7063]), .Z(n10394) );
  XOR U10249 ( .A(n10761), .B(n10762), .Z(n10757) );
  AND U10250 ( .A(n10763), .B(n10764), .Z(n10762) );
  XNOR U10251 ( .A(p_input[7094]), .B(n10761), .Z(n10764) );
  XNOR U10252 ( .A(n10761), .B(n10403), .Z(n10763) );
  IV U10253 ( .A(p_input[7062]), .Z(n10403) );
  XOR U10254 ( .A(n10765), .B(n10766), .Z(n10761) );
  AND U10255 ( .A(n10767), .B(n10768), .Z(n10766) );
  XNOR U10256 ( .A(p_input[7093]), .B(n10765), .Z(n10768) );
  XNOR U10257 ( .A(n10765), .B(n10412), .Z(n10767) );
  IV U10258 ( .A(p_input[7061]), .Z(n10412) );
  XOR U10259 ( .A(n10769), .B(n10770), .Z(n10765) );
  AND U10260 ( .A(n10771), .B(n10772), .Z(n10770) );
  XNOR U10261 ( .A(p_input[7092]), .B(n10769), .Z(n10772) );
  XNOR U10262 ( .A(n10769), .B(n10421), .Z(n10771) );
  IV U10263 ( .A(p_input[7060]), .Z(n10421) );
  XOR U10264 ( .A(n10773), .B(n10774), .Z(n10769) );
  AND U10265 ( .A(n10775), .B(n10776), .Z(n10774) );
  XNOR U10266 ( .A(p_input[7091]), .B(n10773), .Z(n10776) );
  XNOR U10267 ( .A(n10773), .B(n10430), .Z(n10775) );
  IV U10268 ( .A(p_input[7059]), .Z(n10430) );
  XOR U10269 ( .A(n10777), .B(n10778), .Z(n10773) );
  AND U10270 ( .A(n10779), .B(n10780), .Z(n10778) );
  XNOR U10271 ( .A(p_input[7090]), .B(n10777), .Z(n10780) );
  XNOR U10272 ( .A(n10777), .B(n10439), .Z(n10779) );
  IV U10273 ( .A(p_input[7058]), .Z(n10439) );
  XOR U10274 ( .A(n10781), .B(n10782), .Z(n10777) );
  AND U10275 ( .A(n10783), .B(n10784), .Z(n10782) );
  XNOR U10276 ( .A(p_input[7089]), .B(n10781), .Z(n10784) );
  XNOR U10277 ( .A(n10781), .B(n10448), .Z(n10783) );
  IV U10278 ( .A(p_input[7057]), .Z(n10448) );
  XOR U10279 ( .A(n10785), .B(n10786), .Z(n10781) );
  AND U10280 ( .A(n10787), .B(n10788), .Z(n10786) );
  XNOR U10281 ( .A(p_input[7088]), .B(n10785), .Z(n10788) );
  XNOR U10282 ( .A(n10785), .B(n10457), .Z(n10787) );
  IV U10283 ( .A(p_input[7056]), .Z(n10457) );
  XOR U10284 ( .A(n10789), .B(n10790), .Z(n10785) );
  AND U10285 ( .A(n10791), .B(n10792), .Z(n10790) );
  XNOR U10286 ( .A(p_input[7087]), .B(n10789), .Z(n10792) );
  XNOR U10287 ( .A(n10789), .B(n10466), .Z(n10791) );
  IV U10288 ( .A(p_input[7055]), .Z(n10466) );
  XOR U10289 ( .A(n10793), .B(n10794), .Z(n10789) );
  AND U10290 ( .A(n10795), .B(n10796), .Z(n10794) );
  XNOR U10291 ( .A(p_input[7086]), .B(n10793), .Z(n10796) );
  XNOR U10292 ( .A(n10793), .B(n10475), .Z(n10795) );
  IV U10293 ( .A(p_input[7054]), .Z(n10475) );
  XOR U10294 ( .A(n10797), .B(n10798), .Z(n10793) );
  AND U10295 ( .A(n10799), .B(n10800), .Z(n10798) );
  XNOR U10296 ( .A(p_input[7085]), .B(n10797), .Z(n10800) );
  XNOR U10297 ( .A(n10797), .B(n10484), .Z(n10799) );
  IV U10298 ( .A(p_input[7053]), .Z(n10484) );
  XOR U10299 ( .A(n10801), .B(n10802), .Z(n10797) );
  AND U10300 ( .A(n10803), .B(n10804), .Z(n10802) );
  XNOR U10301 ( .A(p_input[7084]), .B(n10801), .Z(n10804) );
  XNOR U10302 ( .A(n10801), .B(n10493), .Z(n10803) );
  IV U10303 ( .A(p_input[7052]), .Z(n10493) );
  XOR U10304 ( .A(n10805), .B(n10806), .Z(n10801) );
  AND U10305 ( .A(n10807), .B(n10808), .Z(n10806) );
  XNOR U10306 ( .A(p_input[7083]), .B(n10805), .Z(n10808) );
  XNOR U10307 ( .A(n10805), .B(n10502), .Z(n10807) );
  IV U10308 ( .A(p_input[7051]), .Z(n10502) );
  XOR U10309 ( .A(n10809), .B(n10810), .Z(n10805) );
  AND U10310 ( .A(n10811), .B(n10812), .Z(n10810) );
  XNOR U10311 ( .A(p_input[7082]), .B(n10809), .Z(n10812) );
  XNOR U10312 ( .A(n10809), .B(n10511), .Z(n10811) );
  IV U10313 ( .A(p_input[7050]), .Z(n10511) );
  XOR U10314 ( .A(n10813), .B(n10814), .Z(n10809) );
  AND U10315 ( .A(n10815), .B(n10816), .Z(n10814) );
  XNOR U10316 ( .A(p_input[7081]), .B(n10813), .Z(n10816) );
  XNOR U10317 ( .A(n10813), .B(n10520), .Z(n10815) );
  IV U10318 ( .A(p_input[7049]), .Z(n10520) );
  XOR U10319 ( .A(n10817), .B(n10818), .Z(n10813) );
  AND U10320 ( .A(n10819), .B(n10820), .Z(n10818) );
  XNOR U10321 ( .A(p_input[7080]), .B(n10817), .Z(n10820) );
  XNOR U10322 ( .A(n10817), .B(n10529), .Z(n10819) );
  IV U10323 ( .A(p_input[7048]), .Z(n10529) );
  XOR U10324 ( .A(n10821), .B(n10822), .Z(n10817) );
  AND U10325 ( .A(n10823), .B(n10824), .Z(n10822) );
  XNOR U10326 ( .A(p_input[7079]), .B(n10821), .Z(n10824) );
  XNOR U10327 ( .A(n10821), .B(n10538), .Z(n10823) );
  IV U10328 ( .A(p_input[7047]), .Z(n10538) );
  XOR U10329 ( .A(n10825), .B(n10826), .Z(n10821) );
  AND U10330 ( .A(n10827), .B(n10828), .Z(n10826) );
  XNOR U10331 ( .A(p_input[7078]), .B(n10825), .Z(n10828) );
  XNOR U10332 ( .A(n10825), .B(n10547), .Z(n10827) );
  IV U10333 ( .A(p_input[7046]), .Z(n10547) );
  XOR U10334 ( .A(n10829), .B(n10830), .Z(n10825) );
  AND U10335 ( .A(n10831), .B(n10832), .Z(n10830) );
  XNOR U10336 ( .A(p_input[7077]), .B(n10829), .Z(n10832) );
  XNOR U10337 ( .A(n10829), .B(n10556), .Z(n10831) );
  IV U10338 ( .A(p_input[7045]), .Z(n10556) );
  XOR U10339 ( .A(n10833), .B(n10834), .Z(n10829) );
  AND U10340 ( .A(n10835), .B(n10836), .Z(n10834) );
  XNOR U10341 ( .A(p_input[7076]), .B(n10833), .Z(n10836) );
  XNOR U10342 ( .A(n10833), .B(n10565), .Z(n10835) );
  IV U10343 ( .A(p_input[7044]), .Z(n10565) );
  XOR U10344 ( .A(n10837), .B(n10838), .Z(n10833) );
  AND U10345 ( .A(n10839), .B(n10840), .Z(n10838) );
  XNOR U10346 ( .A(p_input[7075]), .B(n10837), .Z(n10840) );
  XNOR U10347 ( .A(n10837), .B(n10574), .Z(n10839) );
  IV U10348 ( .A(p_input[7043]), .Z(n10574) );
  XOR U10349 ( .A(n10841), .B(n10842), .Z(n10837) );
  AND U10350 ( .A(n10843), .B(n10844), .Z(n10842) );
  XNOR U10351 ( .A(p_input[7074]), .B(n10841), .Z(n10844) );
  XNOR U10352 ( .A(n10841), .B(n10583), .Z(n10843) );
  IV U10353 ( .A(p_input[7042]), .Z(n10583) );
  XNOR U10354 ( .A(n10845), .B(n10846), .Z(n10841) );
  AND U10355 ( .A(n10847), .B(n10848), .Z(n10846) );
  XOR U10356 ( .A(p_input[7073]), .B(n10845), .Z(n10848) );
  XNOR U10357 ( .A(p_input[7041]), .B(n10845), .Z(n10847) );
  AND U10358 ( .A(p_input[7072]), .B(n10849), .Z(n10845) );
  IV U10359 ( .A(p_input[7040]), .Z(n10849) );
  XOR U10360 ( .A(n10850), .B(n10851), .Z(n9939) );
  AND U10361 ( .A(n465), .B(n10852), .Z(n10851) );
  XNOR U10362 ( .A(n10853), .B(n10850), .Z(n10852) );
  XOR U10363 ( .A(n10854), .B(n10855), .Z(n465) );
  AND U10364 ( .A(n10856), .B(n10857), .Z(n10855) );
  XNOR U10365 ( .A(n9954), .B(n10854), .Z(n10857) );
  AND U10366 ( .A(p_input[7039]), .B(p_input[7007]), .Z(n9954) );
  XNOR U10367 ( .A(n10854), .B(n9951), .Z(n10856) );
  IV U10368 ( .A(n10858), .Z(n9951) );
  AND U10369 ( .A(p_input[6943]), .B(p_input[6975]), .Z(n10858) );
  XOR U10370 ( .A(n10859), .B(n10860), .Z(n10854) );
  AND U10371 ( .A(n10861), .B(n10862), .Z(n10860) );
  XOR U10372 ( .A(n10859), .B(n9966), .Z(n10862) );
  XNOR U10373 ( .A(p_input[7006]), .B(n10863), .Z(n9966) );
  AND U10374 ( .A(n251), .B(n10864), .Z(n10863) );
  XOR U10375 ( .A(p_input[7038]), .B(p_input[7006]), .Z(n10864) );
  XNOR U10376 ( .A(n9963), .B(n10859), .Z(n10861) );
  XOR U10377 ( .A(n10865), .B(n10866), .Z(n9963) );
  AND U10378 ( .A(n248), .B(n10867), .Z(n10866) );
  XOR U10379 ( .A(p_input[6974]), .B(p_input[6942]), .Z(n10867) );
  XOR U10380 ( .A(n10868), .B(n10869), .Z(n10859) );
  AND U10381 ( .A(n10870), .B(n10871), .Z(n10869) );
  XOR U10382 ( .A(n10868), .B(n9978), .Z(n10871) );
  XNOR U10383 ( .A(p_input[7005]), .B(n10872), .Z(n9978) );
  AND U10384 ( .A(n251), .B(n10873), .Z(n10872) );
  XOR U10385 ( .A(p_input[7037]), .B(p_input[7005]), .Z(n10873) );
  XNOR U10386 ( .A(n9975), .B(n10868), .Z(n10870) );
  XOR U10387 ( .A(n10874), .B(n10875), .Z(n9975) );
  AND U10388 ( .A(n248), .B(n10876), .Z(n10875) );
  XOR U10389 ( .A(p_input[6973]), .B(p_input[6941]), .Z(n10876) );
  XOR U10390 ( .A(n10877), .B(n10878), .Z(n10868) );
  AND U10391 ( .A(n10879), .B(n10880), .Z(n10878) );
  XOR U10392 ( .A(n10877), .B(n9990), .Z(n10880) );
  XNOR U10393 ( .A(p_input[7004]), .B(n10881), .Z(n9990) );
  AND U10394 ( .A(n251), .B(n10882), .Z(n10881) );
  XOR U10395 ( .A(p_input[7036]), .B(p_input[7004]), .Z(n10882) );
  XNOR U10396 ( .A(n9987), .B(n10877), .Z(n10879) );
  XOR U10397 ( .A(n10883), .B(n10884), .Z(n9987) );
  AND U10398 ( .A(n248), .B(n10885), .Z(n10884) );
  XOR U10399 ( .A(p_input[6972]), .B(p_input[6940]), .Z(n10885) );
  XOR U10400 ( .A(n10886), .B(n10887), .Z(n10877) );
  AND U10401 ( .A(n10888), .B(n10889), .Z(n10887) );
  XOR U10402 ( .A(n10886), .B(n10002), .Z(n10889) );
  XNOR U10403 ( .A(p_input[7003]), .B(n10890), .Z(n10002) );
  AND U10404 ( .A(n251), .B(n10891), .Z(n10890) );
  XOR U10405 ( .A(p_input[7035]), .B(p_input[7003]), .Z(n10891) );
  XNOR U10406 ( .A(n9999), .B(n10886), .Z(n10888) );
  XOR U10407 ( .A(n10892), .B(n10893), .Z(n9999) );
  AND U10408 ( .A(n248), .B(n10894), .Z(n10893) );
  XOR U10409 ( .A(p_input[6971]), .B(p_input[6939]), .Z(n10894) );
  XOR U10410 ( .A(n10895), .B(n10896), .Z(n10886) );
  AND U10411 ( .A(n10897), .B(n10898), .Z(n10896) );
  XOR U10412 ( .A(n10895), .B(n10014), .Z(n10898) );
  XNOR U10413 ( .A(p_input[7002]), .B(n10899), .Z(n10014) );
  AND U10414 ( .A(n251), .B(n10900), .Z(n10899) );
  XOR U10415 ( .A(p_input[7034]), .B(p_input[7002]), .Z(n10900) );
  XNOR U10416 ( .A(n10011), .B(n10895), .Z(n10897) );
  XOR U10417 ( .A(n10901), .B(n10902), .Z(n10011) );
  AND U10418 ( .A(n248), .B(n10903), .Z(n10902) );
  XOR U10419 ( .A(p_input[6970]), .B(p_input[6938]), .Z(n10903) );
  XOR U10420 ( .A(n10904), .B(n10905), .Z(n10895) );
  AND U10421 ( .A(n10906), .B(n10907), .Z(n10905) );
  XOR U10422 ( .A(n10904), .B(n10026), .Z(n10907) );
  XNOR U10423 ( .A(p_input[7001]), .B(n10908), .Z(n10026) );
  AND U10424 ( .A(n251), .B(n10909), .Z(n10908) );
  XOR U10425 ( .A(p_input[7033]), .B(p_input[7001]), .Z(n10909) );
  XNOR U10426 ( .A(n10023), .B(n10904), .Z(n10906) );
  XOR U10427 ( .A(n10910), .B(n10911), .Z(n10023) );
  AND U10428 ( .A(n248), .B(n10912), .Z(n10911) );
  XOR U10429 ( .A(p_input[6969]), .B(p_input[6937]), .Z(n10912) );
  XOR U10430 ( .A(n10913), .B(n10914), .Z(n10904) );
  AND U10431 ( .A(n10915), .B(n10916), .Z(n10914) );
  XOR U10432 ( .A(n10913), .B(n10038), .Z(n10916) );
  XNOR U10433 ( .A(p_input[7000]), .B(n10917), .Z(n10038) );
  AND U10434 ( .A(n251), .B(n10918), .Z(n10917) );
  XOR U10435 ( .A(p_input[7032]), .B(p_input[7000]), .Z(n10918) );
  XNOR U10436 ( .A(n10035), .B(n10913), .Z(n10915) );
  XOR U10437 ( .A(n10919), .B(n10920), .Z(n10035) );
  AND U10438 ( .A(n248), .B(n10921), .Z(n10920) );
  XOR U10439 ( .A(p_input[6968]), .B(p_input[6936]), .Z(n10921) );
  XOR U10440 ( .A(n10922), .B(n10923), .Z(n10913) );
  AND U10441 ( .A(n10924), .B(n10925), .Z(n10923) );
  XOR U10442 ( .A(n10922), .B(n10050), .Z(n10925) );
  XNOR U10443 ( .A(p_input[6999]), .B(n10926), .Z(n10050) );
  AND U10444 ( .A(n251), .B(n10927), .Z(n10926) );
  XOR U10445 ( .A(p_input[7031]), .B(p_input[6999]), .Z(n10927) );
  XNOR U10446 ( .A(n10047), .B(n10922), .Z(n10924) );
  XOR U10447 ( .A(n10928), .B(n10929), .Z(n10047) );
  AND U10448 ( .A(n248), .B(n10930), .Z(n10929) );
  XOR U10449 ( .A(p_input[6967]), .B(p_input[6935]), .Z(n10930) );
  XOR U10450 ( .A(n10931), .B(n10932), .Z(n10922) );
  AND U10451 ( .A(n10933), .B(n10934), .Z(n10932) );
  XOR U10452 ( .A(n10931), .B(n10062), .Z(n10934) );
  XNOR U10453 ( .A(p_input[6998]), .B(n10935), .Z(n10062) );
  AND U10454 ( .A(n251), .B(n10936), .Z(n10935) );
  XOR U10455 ( .A(p_input[7030]), .B(p_input[6998]), .Z(n10936) );
  XNOR U10456 ( .A(n10059), .B(n10931), .Z(n10933) );
  XOR U10457 ( .A(n10937), .B(n10938), .Z(n10059) );
  AND U10458 ( .A(n248), .B(n10939), .Z(n10938) );
  XOR U10459 ( .A(p_input[6966]), .B(p_input[6934]), .Z(n10939) );
  XOR U10460 ( .A(n10940), .B(n10941), .Z(n10931) );
  AND U10461 ( .A(n10942), .B(n10943), .Z(n10941) );
  XOR U10462 ( .A(n10940), .B(n10074), .Z(n10943) );
  XNOR U10463 ( .A(p_input[6997]), .B(n10944), .Z(n10074) );
  AND U10464 ( .A(n251), .B(n10945), .Z(n10944) );
  XOR U10465 ( .A(p_input[7029]), .B(p_input[6997]), .Z(n10945) );
  XNOR U10466 ( .A(n10071), .B(n10940), .Z(n10942) );
  XOR U10467 ( .A(n10946), .B(n10947), .Z(n10071) );
  AND U10468 ( .A(n248), .B(n10948), .Z(n10947) );
  XOR U10469 ( .A(p_input[6965]), .B(p_input[6933]), .Z(n10948) );
  XOR U10470 ( .A(n10949), .B(n10950), .Z(n10940) );
  AND U10471 ( .A(n10951), .B(n10952), .Z(n10950) );
  XOR U10472 ( .A(n10949), .B(n10086), .Z(n10952) );
  XNOR U10473 ( .A(p_input[6996]), .B(n10953), .Z(n10086) );
  AND U10474 ( .A(n251), .B(n10954), .Z(n10953) );
  XOR U10475 ( .A(p_input[7028]), .B(p_input[6996]), .Z(n10954) );
  XNOR U10476 ( .A(n10083), .B(n10949), .Z(n10951) );
  XOR U10477 ( .A(n10955), .B(n10956), .Z(n10083) );
  AND U10478 ( .A(n248), .B(n10957), .Z(n10956) );
  XOR U10479 ( .A(p_input[6964]), .B(p_input[6932]), .Z(n10957) );
  XOR U10480 ( .A(n10958), .B(n10959), .Z(n10949) );
  AND U10481 ( .A(n10960), .B(n10961), .Z(n10959) );
  XOR U10482 ( .A(n10958), .B(n10098), .Z(n10961) );
  XNOR U10483 ( .A(p_input[6995]), .B(n10962), .Z(n10098) );
  AND U10484 ( .A(n251), .B(n10963), .Z(n10962) );
  XOR U10485 ( .A(p_input[7027]), .B(p_input[6995]), .Z(n10963) );
  XNOR U10486 ( .A(n10095), .B(n10958), .Z(n10960) );
  XOR U10487 ( .A(n10964), .B(n10965), .Z(n10095) );
  AND U10488 ( .A(n248), .B(n10966), .Z(n10965) );
  XOR U10489 ( .A(p_input[6963]), .B(p_input[6931]), .Z(n10966) );
  XOR U10490 ( .A(n10967), .B(n10968), .Z(n10958) );
  AND U10491 ( .A(n10969), .B(n10970), .Z(n10968) );
  XOR U10492 ( .A(n10967), .B(n10110), .Z(n10970) );
  XNOR U10493 ( .A(p_input[6994]), .B(n10971), .Z(n10110) );
  AND U10494 ( .A(n251), .B(n10972), .Z(n10971) );
  XOR U10495 ( .A(p_input[7026]), .B(p_input[6994]), .Z(n10972) );
  XNOR U10496 ( .A(n10107), .B(n10967), .Z(n10969) );
  XOR U10497 ( .A(n10973), .B(n10974), .Z(n10107) );
  AND U10498 ( .A(n248), .B(n10975), .Z(n10974) );
  XOR U10499 ( .A(p_input[6962]), .B(p_input[6930]), .Z(n10975) );
  XOR U10500 ( .A(n10976), .B(n10977), .Z(n10967) );
  AND U10501 ( .A(n10978), .B(n10979), .Z(n10977) );
  XOR U10502 ( .A(n10976), .B(n10122), .Z(n10979) );
  XNOR U10503 ( .A(p_input[6993]), .B(n10980), .Z(n10122) );
  AND U10504 ( .A(n251), .B(n10981), .Z(n10980) );
  XOR U10505 ( .A(p_input[7025]), .B(p_input[6993]), .Z(n10981) );
  XNOR U10506 ( .A(n10119), .B(n10976), .Z(n10978) );
  XOR U10507 ( .A(n10982), .B(n10983), .Z(n10119) );
  AND U10508 ( .A(n248), .B(n10984), .Z(n10983) );
  XOR U10509 ( .A(p_input[6961]), .B(p_input[6929]), .Z(n10984) );
  XOR U10510 ( .A(n10985), .B(n10986), .Z(n10976) );
  AND U10511 ( .A(n10987), .B(n10988), .Z(n10986) );
  XOR U10512 ( .A(n10985), .B(n10134), .Z(n10988) );
  XNOR U10513 ( .A(p_input[6992]), .B(n10989), .Z(n10134) );
  AND U10514 ( .A(n251), .B(n10990), .Z(n10989) );
  XOR U10515 ( .A(p_input[7024]), .B(p_input[6992]), .Z(n10990) );
  XNOR U10516 ( .A(n10131), .B(n10985), .Z(n10987) );
  XOR U10517 ( .A(n10991), .B(n10992), .Z(n10131) );
  AND U10518 ( .A(n248), .B(n10993), .Z(n10992) );
  XOR U10519 ( .A(p_input[6960]), .B(p_input[6928]), .Z(n10993) );
  XOR U10520 ( .A(n10994), .B(n10995), .Z(n10985) );
  AND U10521 ( .A(n10996), .B(n10997), .Z(n10995) );
  XOR U10522 ( .A(n10994), .B(n10146), .Z(n10997) );
  XNOR U10523 ( .A(p_input[6991]), .B(n10998), .Z(n10146) );
  AND U10524 ( .A(n251), .B(n10999), .Z(n10998) );
  XOR U10525 ( .A(p_input[7023]), .B(p_input[6991]), .Z(n10999) );
  XNOR U10526 ( .A(n10143), .B(n10994), .Z(n10996) );
  XOR U10527 ( .A(n11000), .B(n11001), .Z(n10143) );
  AND U10528 ( .A(n248), .B(n11002), .Z(n11001) );
  XOR U10529 ( .A(p_input[6959]), .B(p_input[6927]), .Z(n11002) );
  XOR U10530 ( .A(n11003), .B(n11004), .Z(n10994) );
  AND U10531 ( .A(n11005), .B(n11006), .Z(n11004) );
  XOR U10532 ( .A(n11003), .B(n10158), .Z(n11006) );
  XNOR U10533 ( .A(p_input[6990]), .B(n11007), .Z(n10158) );
  AND U10534 ( .A(n251), .B(n11008), .Z(n11007) );
  XOR U10535 ( .A(p_input[7022]), .B(p_input[6990]), .Z(n11008) );
  XNOR U10536 ( .A(n10155), .B(n11003), .Z(n11005) );
  XOR U10537 ( .A(n11009), .B(n11010), .Z(n10155) );
  AND U10538 ( .A(n248), .B(n11011), .Z(n11010) );
  XOR U10539 ( .A(p_input[6958]), .B(p_input[6926]), .Z(n11011) );
  XOR U10540 ( .A(n11012), .B(n11013), .Z(n11003) );
  AND U10541 ( .A(n11014), .B(n11015), .Z(n11013) );
  XOR U10542 ( .A(n11012), .B(n10170), .Z(n11015) );
  XNOR U10543 ( .A(p_input[6989]), .B(n11016), .Z(n10170) );
  AND U10544 ( .A(n251), .B(n11017), .Z(n11016) );
  XOR U10545 ( .A(p_input[7021]), .B(p_input[6989]), .Z(n11017) );
  XNOR U10546 ( .A(n10167), .B(n11012), .Z(n11014) );
  XOR U10547 ( .A(n11018), .B(n11019), .Z(n10167) );
  AND U10548 ( .A(n248), .B(n11020), .Z(n11019) );
  XOR U10549 ( .A(p_input[6957]), .B(p_input[6925]), .Z(n11020) );
  XOR U10550 ( .A(n11021), .B(n11022), .Z(n11012) );
  AND U10551 ( .A(n11023), .B(n11024), .Z(n11022) );
  XOR U10552 ( .A(n11021), .B(n10182), .Z(n11024) );
  XNOR U10553 ( .A(p_input[6988]), .B(n11025), .Z(n10182) );
  AND U10554 ( .A(n251), .B(n11026), .Z(n11025) );
  XOR U10555 ( .A(p_input[7020]), .B(p_input[6988]), .Z(n11026) );
  XNOR U10556 ( .A(n10179), .B(n11021), .Z(n11023) );
  XOR U10557 ( .A(n11027), .B(n11028), .Z(n10179) );
  AND U10558 ( .A(n248), .B(n11029), .Z(n11028) );
  XOR U10559 ( .A(p_input[6956]), .B(p_input[6924]), .Z(n11029) );
  XOR U10560 ( .A(n11030), .B(n11031), .Z(n11021) );
  AND U10561 ( .A(n11032), .B(n11033), .Z(n11031) );
  XOR U10562 ( .A(n11030), .B(n10194), .Z(n11033) );
  XNOR U10563 ( .A(p_input[6987]), .B(n11034), .Z(n10194) );
  AND U10564 ( .A(n251), .B(n11035), .Z(n11034) );
  XOR U10565 ( .A(p_input[7019]), .B(p_input[6987]), .Z(n11035) );
  XNOR U10566 ( .A(n10191), .B(n11030), .Z(n11032) );
  XOR U10567 ( .A(n11036), .B(n11037), .Z(n10191) );
  AND U10568 ( .A(n248), .B(n11038), .Z(n11037) );
  XOR U10569 ( .A(p_input[6955]), .B(p_input[6923]), .Z(n11038) );
  XOR U10570 ( .A(n11039), .B(n11040), .Z(n11030) );
  AND U10571 ( .A(n11041), .B(n11042), .Z(n11040) );
  XOR U10572 ( .A(n11039), .B(n10206), .Z(n11042) );
  XNOR U10573 ( .A(p_input[6986]), .B(n11043), .Z(n10206) );
  AND U10574 ( .A(n251), .B(n11044), .Z(n11043) );
  XOR U10575 ( .A(p_input[7018]), .B(p_input[6986]), .Z(n11044) );
  XNOR U10576 ( .A(n10203), .B(n11039), .Z(n11041) );
  XOR U10577 ( .A(n11045), .B(n11046), .Z(n10203) );
  AND U10578 ( .A(n248), .B(n11047), .Z(n11046) );
  XOR U10579 ( .A(p_input[6954]), .B(p_input[6922]), .Z(n11047) );
  XOR U10580 ( .A(n11048), .B(n11049), .Z(n11039) );
  AND U10581 ( .A(n11050), .B(n11051), .Z(n11049) );
  XOR U10582 ( .A(n11048), .B(n10218), .Z(n11051) );
  XNOR U10583 ( .A(p_input[6985]), .B(n11052), .Z(n10218) );
  AND U10584 ( .A(n251), .B(n11053), .Z(n11052) );
  XOR U10585 ( .A(p_input[7017]), .B(p_input[6985]), .Z(n11053) );
  XNOR U10586 ( .A(n10215), .B(n11048), .Z(n11050) );
  XOR U10587 ( .A(n11054), .B(n11055), .Z(n10215) );
  AND U10588 ( .A(n248), .B(n11056), .Z(n11055) );
  XOR U10589 ( .A(p_input[6953]), .B(p_input[6921]), .Z(n11056) );
  XOR U10590 ( .A(n11057), .B(n11058), .Z(n11048) );
  AND U10591 ( .A(n11059), .B(n11060), .Z(n11058) );
  XOR U10592 ( .A(n11057), .B(n10230), .Z(n11060) );
  XNOR U10593 ( .A(p_input[6984]), .B(n11061), .Z(n10230) );
  AND U10594 ( .A(n251), .B(n11062), .Z(n11061) );
  XOR U10595 ( .A(p_input[7016]), .B(p_input[6984]), .Z(n11062) );
  XNOR U10596 ( .A(n10227), .B(n11057), .Z(n11059) );
  XOR U10597 ( .A(n11063), .B(n11064), .Z(n10227) );
  AND U10598 ( .A(n248), .B(n11065), .Z(n11064) );
  XOR U10599 ( .A(p_input[6952]), .B(p_input[6920]), .Z(n11065) );
  XOR U10600 ( .A(n11066), .B(n11067), .Z(n11057) );
  AND U10601 ( .A(n11068), .B(n11069), .Z(n11067) );
  XOR U10602 ( .A(n11066), .B(n10242), .Z(n11069) );
  XNOR U10603 ( .A(p_input[6983]), .B(n11070), .Z(n10242) );
  AND U10604 ( .A(n251), .B(n11071), .Z(n11070) );
  XOR U10605 ( .A(p_input[7015]), .B(p_input[6983]), .Z(n11071) );
  XNOR U10606 ( .A(n10239), .B(n11066), .Z(n11068) );
  XOR U10607 ( .A(n11072), .B(n11073), .Z(n10239) );
  AND U10608 ( .A(n248), .B(n11074), .Z(n11073) );
  XOR U10609 ( .A(p_input[6951]), .B(p_input[6919]), .Z(n11074) );
  XOR U10610 ( .A(n11075), .B(n11076), .Z(n11066) );
  AND U10611 ( .A(n11077), .B(n11078), .Z(n11076) );
  XOR U10612 ( .A(n11075), .B(n10254), .Z(n11078) );
  XNOR U10613 ( .A(p_input[6982]), .B(n11079), .Z(n10254) );
  AND U10614 ( .A(n251), .B(n11080), .Z(n11079) );
  XOR U10615 ( .A(p_input[7014]), .B(p_input[6982]), .Z(n11080) );
  XNOR U10616 ( .A(n10251), .B(n11075), .Z(n11077) );
  XOR U10617 ( .A(n11081), .B(n11082), .Z(n10251) );
  AND U10618 ( .A(n248), .B(n11083), .Z(n11082) );
  XOR U10619 ( .A(p_input[6950]), .B(p_input[6918]), .Z(n11083) );
  XOR U10620 ( .A(n11084), .B(n11085), .Z(n11075) );
  AND U10621 ( .A(n11086), .B(n11087), .Z(n11085) );
  XOR U10622 ( .A(n11084), .B(n10266), .Z(n11087) );
  XNOR U10623 ( .A(p_input[6981]), .B(n11088), .Z(n10266) );
  AND U10624 ( .A(n251), .B(n11089), .Z(n11088) );
  XOR U10625 ( .A(p_input[7013]), .B(p_input[6981]), .Z(n11089) );
  XNOR U10626 ( .A(n10263), .B(n11084), .Z(n11086) );
  XOR U10627 ( .A(n11090), .B(n11091), .Z(n10263) );
  AND U10628 ( .A(n248), .B(n11092), .Z(n11091) );
  XOR U10629 ( .A(p_input[6949]), .B(p_input[6917]), .Z(n11092) );
  XOR U10630 ( .A(n11093), .B(n11094), .Z(n11084) );
  AND U10631 ( .A(n11095), .B(n11096), .Z(n11094) );
  XOR U10632 ( .A(n11093), .B(n10278), .Z(n11096) );
  XNOR U10633 ( .A(p_input[6980]), .B(n11097), .Z(n10278) );
  AND U10634 ( .A(n251), .B(n11098), .Z(n11097) );
  XOR U10635 ( .A(p_input[7012]), .B(p_input[6980]), .Z(n11098) );
  XNOR U10636 ( .A(n10275), .B(n11093), .Z(n11095) );
  XOR U10637 ( .A(n11099), .B(n11100), .Z(n10275) );
  AND U10638 ( .A(n248), .B(n11101), .Z(n11100) );
  XOR U10639 ( .A(p_input[6948]), .B(p_input[6916]), .Z(n11101) );
  XOR U10640 ( .A(n11102), .B(n11103), .Z(n11093) );
  AND U10641 ( .A(n11104), .B(n11105), .Z(n11103) );
  XOR U10642 ( .A(n11102), .B(n10290), .Z(n11105) );
  XNOR U10643 ( .A(p_input[6979]), .B(n11106), .Z(n10290) );
  AND U10644 ( .A(n251), .B(n11107), .Z(n11106) );
  XOR U10645 ( .A(p_input[7011]), .B(p_input[6979]), .Z(n11107) );
  XNOR U10646 ( .A(n10287), .B(n11102), .Z(n11104) );
  XOR U10647 ( .A(n11108), .B(n11109), .Z(n10287) );
  AND U10648 ( .A(n248), .B(n11110), .Z(n11109) );
  XOR U10649 ( .A(p_input[6947]), .B(p_input[6915]), .Z(n11110) );
  XOR U10650 ( .A(n11111), .B(n11112), .Z(n11102) );
  AND U10651 ( .A(n11113), .B(n11114), .Z(n11112) );
  XOR U10652 ( .A(n11111), .B(n10302), .Z(n11114) );
  XNOR U10653 ( .A(p_input[6978]), .B(n11115), .Z(n10302) );
  AND U10654 ( .A(n251), .B(n11116), .Z(n11115) );
  XOR U10655 ( .A(p_input[7010]), .B(p_input[6978]), .Z(n11116) );
  XNOR U10656 ( .A(n10299), .B(n11111), .Z(n11113) );
  XOR U10657 ( .A(n11117), .B(n11118), .Z(n10299) );
  AND U10658 ( .A(n248), .B(n11119), .Z(n11118) );
  XOR U10659 ( .A(p_input[6946]), .B(p_input[6914]), .Z(n11119) );
  XOR U10660 ( .A(n11120), .B(n11121), .Z(n11111) );
  AND U10661 ( .A(n11122), .B(n11123), .Z(n11121) );
  XNOR U10662 ( .A(n11124), .B(n10315), .Z(n11123) );
  XNOR U10663 ( .A(p_input[6977]), .B(n11125), .Z(n10315) );
  AND U10664 ( .A(n251), .B(n11126), .Z(n11125) );
  XNOR U10665 ( .A(p_input[7009]), .B(n11127), .Z(n11126) );
  IV U10666 ( .A(p_input[6977]), .Z(n11127) );
  XNOR U10667 ( .A(n10312), .B(n11120), .Z(n11122) );
  XNOR U10668 ( .A(p_input[6913]), .B(n11128), .Z(n10312) );
  AND U10669 ( .A(n248), .B(n11129), .Z(n11128) );
  XOR U10670 ( .A(p_input[6945]), .B(p_input[6913]), .Z(n11129) );
  IV U10671 ( .A(n11124), .Z(n11120) );
  AND U10672 ( .A(n10850), .B(n10853), .Z(n11124) );
  XOR U10673 ( .A(p_input[6976]), .B(n11130), .Z(n10853) );
  AND U10674 ( .A(n251), .B(n11131), .Z(n11130) );
  XOR U10675 ( .A(p_input[7008]), .B(p_input[6976]), .Z(n11131) );
  XOR U10676 ( .A(n11132), .B(n11133), .Z(n251) );
  AND U10677 ( .A(n11134), .B(n11135), .Z(n11133) );
  XNOR U10678 ( .A(p_input[7039]), .B(n11132), .Z(n11135) );
  XOR U10679 ( .A(n11132), .B(p_input[7007]), .Z(n11134) );
  XOR U10680 ( .A(n11136), .B(n11137), .Z(n11132) );
  AND U10681 ( .A(n11138), .B(n11139), .Z(n11137) );
  XNOR U10682 ( .A(p_input[7038]), .B(n11136), .Z(n11139) );
  XOR U10683 ( .A(n11136), .B(p_input[7006]), .Z(n11138) );
  XOR U10684 ( .A(n11140), .B(n11141), .Z(n11136) );
  AND U10685 ( .A(n11142), .B(n11143), .Z(n11141) );
  XNOR U10686 ( .A(p_input[7037]), .B(n11140), .Z(n11143) );
  XOR U10687 ( .A(n11140), .B(p_input[7005]), .Z(n11142) );
  XOR U10688 ( .A(n11144), .B(n11145), .Z(n11140) );
  AND U10689 ( .A(n11146), .B(n11147), .Z(n11145) );
  XNOR U10690 ( .A(p_input[7036]), .B(n11144), .Z(n11147) );
  XOR U10691 ( .A(n11144), .B(p_input[7004]), .Z(n11146) );
  XOR U10692 ( .A(n11148), .B(n11149), .Z(n11144) );
  AND U10693 ( .A(n11150), .B(n11151), .Z(n11149) );
  XNOR U10694 ( .A(p_input[7035]), .B(n11148), .Z(n11151) );
  XOR U10695 ( .A(n11148), .B(p_input[7003]), .Z(n11150) );
  XOR U10696 ( .A(n11152), .B(n11153), .Z(n11148) );
  AND U10697 ( .A(n11154), .B(n11155), .Z(n11153) );
  XNOR U10698 ( .A(p_input[7034]), .B(n11152), .Z(n11155) );
  XOR U10699 ( .A(n11152), .B(p_input[7002]), .Z(n11154) );
  XOR U10700 ( .A(n11156), .B(n11157), .Z(n11152) );
  AND U10701 ( .A(n11158), .B(n11159), .Z(n11157) );
  XNOR U10702 ( .A(p_input[7033]), .B(n11156), .Z(n11159) );
  XOR U10703 ( .A(n11156), .B(p_input[7001]), .Z(n11158) );
  XOR U10704 ( .A(n11160), .B(n11161), .Z(n11156) );
  AND U10705 ( .A(n11162), .B(n11163), .Z(n11161) );
  XNOR U10706 ( .A(p_input[7032]), .B(n11160), .Z(n11163) );
  XOR U10707 ( .A(n11160), .B(p_input[7000]), .Z(n11162) );
  XOR U10708 ( .A(n11164), .B(n11165), .Z(n11160) );
  AND U10709 ( .A(n11166), .B(n11167), .Z(n11165) );
  XNOR U10710 ( .A(p_input[7031]), .B(n11164), .Z(n11167) );
  XOR U10711 ( .A(n11164), .B(p_input[6999]), .Z(n11166) );
  XOR U10712 ( .A(n11168), .B(n11169), .Z(n11164) );
  AND U10713 ( .A(n11170), .B(n11171), .Z(n11169) );
  XNOR U10714 ( .A(p_input[7030]), .B(n11168), .Z(n11171) );
  XOR U10715 ( .A(n11168), .B(p_input[6998]), .Z(n11170) );
  XOR U10716 ( .A(n11172), .B(n11173), .Z(n11168) );
  AND U10717 ( .A(n11174), .B(n11175), .Z(n11173) );
  XNOR U10718 ( .A(p_input[7029]), .B(n11172), .Z(n11175) );
  XOR U10719 ( .A(n11172), .B(p_input[6997]), .Z(n11174) );
  XOR U10720 ( .A(n11176), .B(n11177), .Z(n11172) );
  AND U10721 ( .A(n11178), .B(n11179), .Z(n11177) );
  XNOR U10722 ( .A(p_input[7028]), .B(n11176), .Z(n11179) );
  XOR U10723 ( .A(n11176), .B(p_input[6996]), .Z(n11178) );
  XOR U10724 ( .A(n11180), .B(n11181), .Z(n11176) );
  AND U10725 ( .A(n11182), .B(n11183), .Z(n11181) );
  XNOR U10726 ( .A(p_input[7027]), .B(n11180), .Z(n11183) );
  XOR U10727 ( .A(n11180), .B(p_input[6995]), .Z(n11182) );
  XOR U10728 ( .A(n11184), .B(n11185), .Z(n11180) );
  AND U10729 ( .A(n11186), .B(n11187), .Z(n11185) );
  XNOR U10730 ( .A(p_input[7026]), .B(n11184), .Z(n11187) );
  XOR U10731 ( .A(n11184), .B(p_input[6994]), .Z(n11186) );
  XOR U10732 ( .A(n11188), .B(n11189), .Z(n11184) );
  AND U10733 ( .A(n11190), .B(n11191), .Z(n11189) );
  XNOR U10734 ( .A(p_input[7025]), .B(n11188), .Z(n11191) );
  XOR U10735 ( .A(n11188), .B(p_input[6993]), .Z(n11190) );
  XOR U10736 ( .A(n11192), .B(n11193), .Z(n11188) );
  AND U10737 ( .A(n11194), .B(n11195), .Z(n11193) );
  XNOR U10738 ( .A(p_input[7024]), .B(n11192), .Z(n11195) );
  XOR U10739 ( .A(n11192), .B(p_input[6992]), .Z(n11194) );
  XOR U10740 ( .A(n11196), .B(n11197), .Z(n11192) );
  AND U10741 ( .A(n11198), .B(n11199), .Z(n11197) );
  XNOR U10742 ( .A(p_input[7023]), .B(n11196), .Z(n11199) );
  XOR U10743 ( .A(n11196), .B(p_input[6991]), .Z(n11198) );
  XOR U10744 ( .A(n11200), .B(n11201), .Z(n11196) );
  AND U10745 ( .A(n11202), .B(n11203), .Z(n11201) );
  XNOR U10746 ( .A(p_input[7022]), .B(n11200), .Z(n11203) );
  XOR U10747 ( .A(n11200), .B(p_input[6990]), .Z(n11202) );
  XOR U10748 ( .A(n11204), .B(n11205), .Z(n11200) );
  AND U10749 ( .A(n11206), .B(n11207), .Z(n11205) );
  XNOR U10750 ( .A(p_input[7021]), .B(n11204), .Z(n11207) );
  XOR U10751 ( .A(n11204), .B(p_input[6989]), .Z(n11206) );
  XOR U10752 ( .A(n11208), .B(n11209), .Z(n11204) );
  AND U10753 ( .A(n11210), .B(n11211), .Z(n11209) );
  XNOR U10754 ( .A(p_input[7020]), .B(n11208), .Z(n11211) );
  XOR U10755 ( .A(n11208), .B(p_input[6988]), .Z(n11210) );
  XOR U10756 ( .A(n11212), .B(n11213), .Z(n11208) );
  AND U10757 ( .A(n11214), .B(n11215), .Z(n11213) );
  XNOR U10758 ( .A(p_input[7019]), .B(n11212), .Z(n11215) );
  XOR U10759 ( .A(n11212), .B(p_input[6987]), .Z(n11214) );
  XOR U10760 ( .A(n11216), .B(n11217), .Z(n11212) );
  AND U10761 ( .A(n11218), .B(n11219), .Z(n11217) );
  XNOR U10762 ( .A(p_input[7018]), .B(n11216), .Z(n11219) );
  XOR U10763 ( .A(n11216), .B(p_input[6986]), .Z(n11218) );
  XOR U10764 ( .A(n11220), .B(n11221), .Z(n11216) );
  AND U10765 ( .A(n11222), .B(n11223), .Z(n11221) );
  XNOR U10766 ( .A(p_input[7017]), .B(n11220), .Z(n11223) );
  XOR U10767 ( .A(n11220), .B(p_input[6985]), .Z(n11222) );
  XOR U10768 ( .A(n11224), .B(n11225), .Z(n11220) );
  AND U10769 ( .A(n11226), .B(n11227), .Z(n11225) );
  XNOR U10770 ( .A(p_input[7016]), .B(n11224), .Z(n11227) );
  XOR U10771 ( .A(n11224), .B(p_input[6984]), .Z(n11226) );
  XOR U10772 ( .A(n11228), .B(n11229), .Z(n11224) );
  AND U10773 ( .A(n11230), .B(n11231), .Z(n11229) );
  XNOR U10774 ( .A(p_input[7015]), .B(n11228), .Z(n11231) );
  XOR U10775 ( .A(n11228), .B(p_input[6983]), .Z(n11230) );
  XOR U10776 ( .A(n11232), .B(n11233), .Z(n11228) );
  AND U10777 ( .A(n11234), .B(n11235), .Z(n11233) );
  XNOR U10778 ( .A(p_input[7014]), .B(n11232), .Z(n11235) );
  XOR U10779 ( .A(n11232), .B(p_input[6982]), .Z(n11234) );
  XOR U10780 ( .A(n11236), .B(n11237), .Z(n11232) );
  AND U10781 ( .A(n11238), .B(n11239), .Z(n11237) );
  XNOR U10782 ( .A(p_input[7013]), .B(n11236), .Z(n11239) );
  XOR U10783 ( .A(n11236), .B(p_input[6981]), .Z(n11238) );
  XOR U10784 ( .A(n11240), .B(n11241), .Z(n11236) );
  AND U10785 ( .A(n11242), .B(n11243), .Z(n11241) );
  XNOR U10786 ( .A(p_input[7012]), .B(n11240), .Z(n11243) );
  XOR U10787 ( .A(n11240), .B(p_input[6980]), .Z(n11242) );
  XOR U10788 ( .A(n11244), .B(n11245), .Z(n11240) );
  AND U10789 ( .A(n11246), .B(n11247), .Z(n11245) );
  XNOR U10790 ( .A(p_input[7011]), .B(n11244), .Z(n11247) );
  XOR U10791 ( .A(n11244), .B(p_input[6979]), .Z(n11246) );
  XOR U10792 ( .A(n11248), .B(n11249), .Z(n11244) );
  AND U10793 ( .A(n11250), .B(n11251), .Z(n11249) );
  XNOR U10794 ( .A(p_input[7010]), .B(n11248), .Z(n11251) );
  XOR U10795 ( .A(n11248), .B(p_input[6978]), .Z(n11250) );
  XNOR U10796 ( .A(n11252), .B(n11253), .Z(n11248) );
  AND U10797 ( .A(n11254), .B(n11255), .Z(n11253) );
  XOR U10798 ( .A(p_input[7009]), .B(n11252), .Z(n11255) );
  XNOR U10799 ( .A(p_input[6977]), .B(n11252), .Z(n11254) );
  AND U10800 ( .A(p_input[7008]), .B(n11256), .Z(n11252) );
  IV U10801 ( .A(p_input[6976]), .Z(n11256) );
  XNOR U10802 ( .A(p_input[6912]), .B(n11257), .Z(n10850) );
  AND U10803 ( .A(n248), .B(n11258), .Z(n11257) );
  XOR U10804 ( .A(p_input[6944]), .B(p_input[6912]), .Z(n11258) );
  XOR U10805 ( .A(n11259), .B(n11260), .Z(n248) );
  AND U10806 ( .A(n11261), .B(n11262), .Z(n11260) );
  XNOR U10807 ( .A(p_input[6975]), .B(n11259), .Z(n11262) );
  XOR U10808 ( .A(n11259), .B(p_input[6943]), .Z(n11261) );
  XOR U10809 ( .A(n11263), .B(n11264), .Z(n11259) );
  AND U10810 ( .A(n11265), .B(n11266), .Z(n11264) );
  XNOR U10811 ( .A(p_input[6974]), .B(n11263), .Z(n11266) );
  XNOR U10812 ( .A(n11263), .B(n10865), .Z(n11265) );
  IV U10813 ( .A(p_input[6942]), .Z(n10865) );
  XOR U10814 ( .A(n11267), .B(n11268), .Z(n11263) );
  AND U10815 ( .A(n11269), .B(n11270), .Z(n11268) );
  XNOR U10816 ( .A(p_input[6973]), .B(n11267), .Z(n11270) );
  XNOR U10817 ( .A(n11267), .B(n10874), .Z(n11269) );
  IV U10818 ( .A(p_input[6941]), .Z(n10874) );
  XOR U10819 ( .A(n11271), .B(n11272), .Z(n11267) );
  AND U10820 ( .A(n11273), .B(n11274), .Z(n11272) );
  XNOR U10821 ( .A(p_input[6972]), .B(n11271), .Z(n11274) );
  XNOR U10822 ( .A(n11271), .B(n10883), .Z(n11273) );
  IV U10823 ( .A(p_input[6940]), .Z(n10883) );
  XOR U10824 ( .A(n11275), .B(n11276), .Z(n11271) );
  AND U10825 ( .A(n11277), .B(n11278), .Z(n11276) );
  XNOR U10826 ( .A(p_input[6971]), .B(n11275), .Z(n11278) );
  XNOR U10827 ( .A(n11275), .B(n10892), .Z(n11277) );
  IV U10828 ( .A(p_input[6939]), .Z(n10892) );
  XOR U10829 ( .A(n11279), .B(n11280), .Z(n11275) );
  AND U10830 ( .A(n11281), .B(n11282), .Z(n11280) );
  XNOR U10831 ( .A(p_input[6970]), .B(n11279), .Z(n11282) );
  XNOR U10832 ( .A(n11279), .B(n10901), .Z(n11281) );
  IV U10833 ( .A(p_input[6938]), .Z(n10901) );
  XOR U10834 ( .A(n11283), .B(n11284), .Z(n11279) );
  AND U10835 ( .A(n11285), .B(n11286), .Z(n11284) );
  XNOR U10836 ( .A(p_input[6969]), .B(n11283), .Z(n11286) );
  XNOR U10837 ( .A(n11283), .B(n10910), .Z(n11285) );
  IV U10838 ( .A(p_input[6937]), .Z(n10910) );
  XOR U10839 ( .A(n11287), .B(n11288), .Z(n11283) );
  AND U10840 ( .A(n11289), .B(n11290), .Z(n11288) );
  XNOR U10841 ( .A(p_input[6968]), .B(n11287), .Z(n11290) );
  XNOR U10842 ( .A(n11287), .B(n10919), .Z(n11289) );
  IV U10843 ( .A(p_input[6936]), .Z(n10919) );
  XOR U10844 ( .A(n11291), .B(n11292), .Z(n11287) );
  AND U10845 ( .A(n11293), .B(n11294), .Z(n11292) );
  XNOR U10846 ( .A(p_input[6967]), .B(n11291), .Z(n11294) );
  XNOR U10847 ( .A(n11291), .B(n10928), .Z(n11293) );
  IV U10848 ( .A(p_input[6935]), .Z(n10928) );
  XOR U10849 ( .A(n11295), .B(n11296), .Z(n11291) );
  AND U10850 ( .A(n11297), .B(n11298), .Z(n11296) );
  XNOR U10851 ( .A(p_input[6966]), .B(n11295), .Z(n11298) );
  XNOR U10852 ( .A(n11295), .B(n10937), .Z(n11297) );
  IV U10853 ( .A(p_input[6934]), .Z(n10937) );
  XOR U10854 ( .A(n11299), .B(n11300), .Z(n11295) );
  AND U10855 ( .A(n11301), .B(n11302), .Z(n11300) );
  XNOR U10856 ( .A(p_input[6965]), .B(n11299), .Z(n11302) );
  XNOR U10857 ( .A(n11299), .B(n10946), .Z(n11301) );
  IV U10858 ( .A(p_input[6933]), .Z(n10946) );
  XOR U10859 ( .A(n11303), .B(n11304), .Z(n11299) );
  AND U10860 ( .A(n11305), .B(n11306), .Z(n11304) );
  XNOR U10861 ( .A(p_input[6964]), .B(n11303), .Z(n11306) );
  XNOR U10862 ( .A(n11303), .B(n10955), .Z(n11305) );
  IV U10863 ( .A(p_input[6932]), .Z(n10955) );
  XOR U10864 ( .A(n11307), .B(n11308), .Z(n11303) );
  AND U10865 ( .A(n11309), .B(n11310), .Z(n11308) );
  XNOR U10866 ( .A(p_input[6963]), .B(n11307), .Z(n11310) );
  XNOR U10867 ( .A(n11307), .B(n10964), .Z(n11309) );
  IV U10868 ( .A(p_input[6931]), .Z(n10964) );
  XOR U10869 ( .A(n11311), .B(n11312), .Z(n11307) );
  AND U10870 ( .A(n11313), .B(n11314), .Z(n11312) );
  XNOR U10871 ( .A(p_input[6962]), .B(n11311), .Z(n11314) );
  XNOR U10872 ( .A(n11311), .B(n10973), .Z(n11313) );
  IV U10873 ( .A(p_input[6930]), .Z(n10973) );
  XOR U10874 ( .A(n11315), .B(n11316), .Z(n11311) );
  AND U10875 ( .A(n11317), .B(n11318), .Z(n11316) );
  XNOR U10876 ( .A(p_input[6961]), .B(n11315), .Z(n11318) );
  XNOR U10877 ( .A(n11315), .B(n10982), .Z(n11317) );
  IV U10878 ( .A(p_input[6929]), .Z(n10982) );
  XOR U10879 ( .A(n11319), .B(n11320), .Z(n11315) );
  AND U10880 ( .A(n11321), .B(n11322), .Z(n11320) );
  XNOR U10881 ( .A(p_input[6960]), .B(n11319), .Z(n11322) );
  XNOR U10882 ( .A(n11319), .B(n10991), .Z(n11321) );
  IV U10883 ( .A(p_input[6928]), .Z(n10991) );
  XOR U10884 ( .A(n11323), .B(n11324), .Z(n11319) );
  AND U10885 ( .A(n11325), .B(n11326), .Z(n11324) );
  XNOR U10886 ( .A(p_input[6959]), .B(n11323), .Z(n11326) );
  XNOR U10887 ( .A(n11323), .B(n11000), .Z(n11325) );
  IV U10888 ( .A(p_input[6927]), .Z(n11000) );
  XOR U10889 ( .A(n11327), .B(n11328), .Z(n11323) );
  AND U10890 ( .A(n11329), .B(n11330), .Z(n11328) );
  XNOR U10891 ( .A(p_input[6958]), .B(n11327), .Z(n11330) );
  XNOR U10892 ( .A(n11327), .B(n11009), .Z(n11329) );
  IV U10893 ( .A(p_input[6926]), .Z(n11009) );
  XOR U10894 ( .A(n11331), .B(n11332), .Z(n11327) );
  AND U10895 ( .A(n11333), .B(n11334), .Z(n11332) );
  XNOR U10896 ( .A(p_input[6957]), .B(n11331), .Z(n11334) );
  XNOR U10897 ( .A(n11331), .B(n11018), .Z(n11333) );
  IV U10898 ( .A(p_input[6925]), .Z(n11018) );
  XOR U10899 ( .A(n11335), .B(n11336), .Z(n11331) );
  AND U10900 ( .A(n11337), .B(n11338), .Z(n11336) );
  XNOR U10901 ( .A(p_input[6956]), .B(n11335), .Z(n11338) );
  XNOR U10902 ( .A(n11335), .B(n11027), .Z(n11337) );
  IV U10903 ( .A(p_input[6924]), .Z(n11027) );
  XOR U10904 ( .A(n11339), .B(n11340), .Z(n11335) );
  AND U10905 ( .A(n11341), .B(n11342), .Z(n11340) );
  XNOR U10906 ( .A(p_input[6955]), .B(n11339), .Z(n11342) );
  XNOR U10907 ( .A(n11339), .B(n11036), .Z(n11341) );
  IV U10908 ( .A(p_input[6923]), .Z(n11036) );
  XOR U10909 ( .A(n11343), .B(n11344), .Z(n11339) );
  AND U10910 ( .A(n11345), .B(n11346), .Z(n11344) );
  XNOR U10911 ( .A(p_input[6954]), .B(n11343), .Z(n11346) );
  XNOR U10912 ( .A(n11343), .B(n11045), .Z(n11345) );
  IV U10913 ( .A(p_input[6922]), .Z(n11045) );
  XOR U10914 ( .A(n11347), .B(n11348), .Z(n11343) );
  AND U10915 ( .A(n11349), .B(n11350), .Z(n11348) );
  XNOR U10916 ( .A(p_input[6953]), .B(n11347), .Z(n11350) );
  XNOR U10917 ( .A(n11347), .B(n11054), .Z(n11349) );
  IV U10918 ( .A(p_input[6921]), .Z(n11054) );
  XOR U10919 ( .A(n11351), .B(n11352), .Z(n11347) );
  AND U10920 ( .A(n11353), .B(n11354), .Z(n11352) );
  XNOR U10921 ( .A(p_input[6952]), .B(n11351), .Z(n11354) );
  XNOR U10922 ( .A(n11351), .B(n11063), .Z(n11353) );
  IV U10923 ( .A(p_input[6920]), .Z(n11063) );
  XOR U10924 ( .A(n11355), .B(n11356), .Z(n11351) );
  AND U10925 ( .A(n11357), .B(n11358), .Z(n11356) );
  XNOR U10926 ( .A(p_input[6951]), .B(n11355), .Z(n11358) );
  XNOR U10927 ( .A(n11355), .B(n11072), .Z(n11357) );
  IV U10928 ( .A(p_input[6919]), .Z(n11072) );
  XOR U10929 ( .A(n11359), .B(n11360), .Z(n11355) );
  AND U10930 ( .A(n11361), .B(n11362), .Z(n11360) );
  XNOR U10931 ( .A(p_input[6950]), .B(n11359), .Z(n11362) );
  XNOR U10932 ( .A(n11359), .B(n11081), .Z(n11361) );
  IV U10933 ( .A(p_input[6918]), .Z(n11081) );
  XOR U10934 ( .A(n11363), .B(n11364), .Z(n11359) );
  AND U10935 ( .A(n11365), .B(n11366), .Z(n11364) );
  XNOR U10936 ( .A(p_input[6949]), .B(n11363), .Z(n11366) );
  XNOR U10937 ( .A(n11363), .B(n11090), .Z(n11365) );
  IV U10938 ( .A(p_input[6917]), .Z(n11090) );
  XOR U10939 ( .A(n11367), .B(n11368), .Z(n11363) );
  AND U10940 ( .A(n11369), .B(n11370), .Z(n11368) );
  XNOR U10941 ( .A(p_input[6948]), .B(n11367), .Z(n11370) );
  XNOR U10942 ( .A(n11367), .B(n11099), .Z(n11369) );
  IV U10943 ( .A(p_input[6916]), .Z(n11099) );
  XOR U10944 ( .A(n11371), .B(n11372), .Z(n11367) );
  AND U10945 ( .A(n11373), .B(n11374), .Z(n11372) );
  XNOR U10946 ( .A(p_input[6947]), .B(n11371), .Z(n11374) );
  XNOR U10947 ( .A(n11371), .B(n11108), .Z(n11373) );
  IV U10948 ( .A(p_input[6915]), .Z(n11108) );
  XOR U10949 ( .A(n11375), .B(n11376), .Z(n11371) );
  AND U10950 ( .A(n11377), .B(n11378), .Z(n11376) );
  XNOR U10951 ( .A(p_input[6946]), .B(n11375), .Z(n11378) );
  XNOR U10952 ( .A(n11375), .B(n11117), .Z(n11377) );
  IV U10953 ( .A(p_input[6914]), .Z(n11117) );
  XNOR U10954 ( .A(n11379), .B(n11380), .Z(n11375) );
  AND U10955 ( .A(n11381), .B(n11382), .Z(n11380) );
  XOR U10956 ( .A(p_input[6945]), .B(n11379), .Z(n11382) );
  XNOR U10957 ( .A(p_input[6913]), .B(n11379), .Z(n11381) );
  AND U10958 ( .A(p_input[6944]), .B(n11383), .Z(n11379) );
  IV U10959 ( .A(p_input[6912]), .Z(n11383) );
  XOR U10960 ( .A(n11384), .B(n11385), .Z(n9562) );
  AND U10961 ( .A(n825), .B(n11386), .Z(n11385) );
  XNOR U10962 ( .A(n11387), .B(n11384), .Z(n11386) );
  XOR U10963 ( .A(n11388), .B(n11389), .Z(n825) );
  AND U10964 ( .A(n11390), .B(n11391), .Z(n11389) );
  XOR U10965 ( .A(n11388), .B(n9577), .Z(n11391) );
  XNOR U10966 ( .A(n11392), .B(n11393), .Z(n9577) );
  AND U10967 ( .A(n11394), .B(n471), .Z(n11393) );
  AND U10968 ( .A(n11392), .B(n11395), .Z(n11394) );
  XNOR U10969 ( .A(n9574), .B(n11388), .Z(n11390) );
  XOR U10970 ( .A(n11396), .B(n11397), .Z(n9574) );
  AND U10971 ( .A(n11398), .B(n468), .Z(n11397) );
  NOR U10972 ( .A(n11396), .B(n11399), .Z(n11398) );
  XOR U10973 ( .A(n11400), .B(n11401), .Z(n11388) );
  AND U10974 ( .A(n11402), .B(n11403), .Z(n11401) );
  XOR U10975 ( .A(n11400), .B(n9589), .Z(n11403) );
  XOR U10976 ( .A(n11404), .B(n11405), .Z(n9589) );
  AND U10977 ( .A(n471), .B(n11406), .Z(n11405) );
  XOR U10978 ( .A(n11407), .B(n11404), .Z(n11406) );
  XNOR U10979 ( .A(n9586), .B(n11400), .Z(n11402) );
  XOR U10980 ( .A(n11408), .B(n11409), .Z(n9586) );
  AND U10981 ( .A(n468), .B(n11410), .Z(n11409) );
  XOR U10982 ( .A(n11411), .B(n11408), .Z(n11410) );
  XOR U10983 ( .A(n11412), .B(n11413), .Z(n11400) );
  AND U10984 ( .A(n11414), .B(n11415), .Z(n11413) );
  XOR U10985 ( .A(n11412), .B(n9601), .Z(n11415) );
  XOR U10986 ( .A(n11416), .B(n11417), .Z(n9601) );
  AND U10987 ( .A(n471), .B(n11418), .Z(n11417) );
  XOR U10988 ( .A(n11419), .B(n11416), .Z(n11418) );
  XNOR U10989 ( .A(n9598), .B(n11412), .Z(n11414) );
  XOR U10990 ( .A(n11420), .B(n11421), .Z(n9598) );
  AND U10991 ( .A(n468), .B(n11422), .Z(n11421) );
  XOR U10992 ( .A(n11423), .B(n11420), .Z(n11422) );
  XOR U10993 ( .A(n11424), .B(n11425), .Z(n11412) );
  AND U10994 ( .A(n11426), .B(n11427), .Z(n11425) );
  XOR U10995 ( .A(n11424), .B(n9613), .Z(n11427) );
  XOR U10996 ( .A(n11428), .B(n11429), .Z(n9613) );
  AND U10997 ( .A(n471), .B(n11430), .Z(n11429) );
  XOR U10998 ( .A(n11431), .B(n11428), .Z(n11430) );
  XNOR U10999 ( .A(n9610), .B(n11424), .Z(n11426) );
  XOR U11000 ( .A(n11432), .B(n11433), .Z(n9610) );
  AND U11001 ( .A(n468), .B(n11434), .Z(n11433) );
  XOR U11002 ( .A(n11435), .B(n11432), .Z(n11434) );
  XOR U11003 ( .A(n11436), .B(n11437), .Z(n11424) );
  AND U11004 ( .A(n11438), .B(n11439), .Z(n11437) );
  XOR U11005 ( .A(n11436), .B(n9625), .Z(n11439) );
  XOR U11006 ( .A(n11440), .B(n11441), .Z(n9625) );
  AND U11007 ( .A(n471), .B(n11442), .Z(n11441) );
  XOR U11008 ( .A(n11443), .B(n11440), .Z(n11442) );
  XNOR U11009 ( .A(n9622), .B(n11436), .Z(n11438) );
  XOR U11010 ( .A(n11444), .B(n11445), .Z(n9622) );
  AND U11011 ( .A(n468), .B(n11446), .Z(n11445) );
  XOR U11012 ( .A(n11447), .B(n11444), .Z(n11446) );
  XOR U11013 ( .A(n11448), .B(n11449), .Z(n11436) );
  AND U11014 ( .A(n11450), .B(n11451), .Z(n11449) );
  XOR U11015 ( .A(n11448), .B(n9637), .Z(n11451) );
  XOR U11016 ( .A(n11452), .B(n11453), .Z(n9637) );
  AND U11017 ( .A(n471), .B(n11454), .Z(n11453) );
  XOR U11018 ( .A(n11455), .B(n11452), .Z(n11454) );
  XNOR U11019 ( .A(n9634), .B(n11448), .Z(n11450) );
  XOR U11020 ( .A(n11456), .B(n11457), .Z(n9634) );
  AND U11021 ( .A(n468), .B(n11458), .Z(n11457) );
  XOR U11022 ( .A(n11459), .B(n11456), .Z(n11458) );
  XOR U11023 ( .A(n11460), .B(n11461), .Z(n11448) );
  AND U11024 ( .A(n11462), .B(n11463), .Z(n11461) );
  XOR U11025 ( .A(n11460), .B(n9649), .Z(n11463) );
  XOR U11026 ( .A(n11464), .B(n11465), .Z(n9649) );
  AND U11027 ( .A(n471), .B(n11466), .Z(n11465) );
  XOR U11028 ( .A(n11467), .B(n11464), .Z(n11466) );
  XNOR U11029 ( .A(n9646), .B(n11460), .Z(n11462) );
  XOR U11030 ( .A(n11468), .B(n11469), .Z(n9646) );
  AND U11031 ( .A(n468), .B(n11470), .Z(n11469) );
  XOR U11032 ( .A(n11471), .B(n11468), .Z(n11470) );
  XOR U11033 ( .A(n11472), .B(n11473), .Z(n11460) );
  AND U11034 ( .A(n11474), .B(n11475), .Z(n11473) );
  XOR U11035 ( .A(n11472), .B(n9661), .Z(n11475) );
  XOR U11036 ( .A(n11476), .B(n11477), .Z(n9661) );
  AND U11037 ( .A(n471), .B(n11478), .Z(n11477) );
  XOR U11038 ( .A(n11479), .B(n11476), .Z(n11478) );
  XNOR U11039 ( .A(n9658), .B(n11472), .Z(n11474) );
  XOR U11040 ( .A(n11480), .B(n11481), .Z(n9658) );
  AND U11041 ( .A(n468), .B(n11482), .Z(n11481) );
  XOR U11042 ( .A(n11483), .B(n11480), .Z(n11482) );
  XOR U11043 ( .A(n11484), .B(n11485), .Z(n11472) );
  AND U11044 ( .A(n11486), .B(n11487), .Z(n11485) );
  XOR U11045 ( .A(n11484), .B(n9673), .Z(n11487) );
  XOR U11046 ( .A(n11488), .B(n11489), .Z(n9673) );
  AND U11047 ( .A(n471), .B(n11490), .Z(n11489) );
  XOR U11048 ( .A(n11491), .B(n11488), .Z(n11490) );
  XNOR U11049 ( .A(n9670), .B(n11484), .Z(n11486) );
  XOR U11050 ( .A(n11492), .B(n11493), .Z(n9670) );
  AND U11051 ( .A(n468), .B(n11494), .Z(n11493) );
  XOR U11052 ( .A(n11495), .B(n11492), .Z(n11494) );
  XOR U11053 ( .A(n11496), .B(n11497), .Z(n11484) );
  AND U11054 ( .A(n11498), .B(n11499), .Z(n11497) );
  XOR U11055 ( .A(n11496), .B(n9685), .Z(n11499) );
  XOR U11056 ( .A(n11500), .B(n11501), .Z(n9685) );
  AND U11057 ( .A(n471), .B(n11502), .Z(n11501) );
  XOR U11058 ( .A(n11503), .B(n11500), .Z(n11502) );
  XNOR U11059 ( .A(n9682), .B(n11496), .Z(n11498) );
  XOR U11060 ( .A(n11504), .B(n11505), .Z(n9682) );
  AND U11061 ( .A(n468), .B(n11506), .Z(n11505) );
  XOR U11062 ( .A(n11507), .B(n11504), .Z(n11506) );
  XOR U11063 ( .A(n11508), .B(n11509), .Z(n11496) );
  AND U11064 ( .A(n11510), .B(n11511), .Z(n11509) );
  XOR U11065 ( .A(n11508), .B(n9697), .Z(n11511) );
  XOR U11066 ( .A(n11512), .B(n11513), .Z(n9697) );
  AND U11067 ( .A(n471), .B(n11514), .Z(n11513) );
  XOR U11068 ( .A(n11515), .B(n11512), .Z(n11514) );
  XNOR U11069 ( .A(n9694), .B(n11508), .Z(n11510) );
  XOR U11070 ( .A(n11516), .B(n11517), .Z(n9694) );
  AND U11071 ( .A(n468), .B(n11518), .Z(n11517) );
  XOR U11072 ( .A(n11519), .B(n11516), .Z(n11518) );
  XOR U11073 ( .A(n11520), .B(n11521), .Z(n11508) );
  AND U11074 ( .A(n11522), .B(n11523), .Z(n11521) );
  XOR U11075 ( .A(n11520), .B(n9709), .Z(n11523) );
  XOR U11076 ( .A(n11524), .B(n11525), .Z(n9709) );
  AND U11077 ( .A(n471), .B(n11526), .Z(n11525) );
  XOR U11078 ( .A(n11527), .B(n11524), .Z(n11526) );
  XNOR U11079 ( .A(n9706), .B(n11520), .Z(n11522) );
  XOR U11080 ( .A(n11528), .B(n11529), .Z(n9706) );
  AND U11081 ( .A(n468), .B(n11530), .Z(n11529) );
  XOR U11082 ( .A(n11531), .B(n11528), .Z(n11530) );
  XOR U11083 ( .A(n11532), .B(n11533), .Z(n11520) );
  AND U11084 ( .A(n11534), .B(n11535), .Z(n11533) );
  XOR U11085 ( .A(n11532), .B(n9721), .Z(n11535) );
  XOR U11086 ( .A(n11536), .B(n11537), .Z(n9721) );
  AND U11087 ( .A(n471), .B(n11538), .Z(n11537) );
  XOR U11088 ( .A(n11539), .B(n11536), .Z(n11538) );
  XNOR U11089 ( .A(n9718), .B(n11532), .Z(n11534) );
  XOR U11090 ( .A(n11540), .B(n11541), .Z(n9718) );
  AND U11091 ( .A(n468), .B(n11542), .Z(n11541) );
  XOR U11092 ( .A(n11543), .B(n11540), .Z(n11542) );
  XOR U11093 ( .A(n11544), .B(n11545), .Z(n11532) );
  AND U11094 ( .A(n11546), .B(n11547), .Z(n11545) );
  XOR U11095 ( .A(n11544), .B(n9733), .Z(n11547) );
  XOR U11096 ( .A(n11548), .B(n11549), .Z(n9733) );
  AND U11097 ( .A(n471), .B(n11550), .Z(n11549) );
  XOR U11098 ( .A(n11551), .B(n11548), .Z(n11550) );
  XNOR U11099 ( .A(n9730), .B(n11544), .Z(n11546) );
  XOR U11100 ( .A(n11552), .B(n11553), .Z(n9730) );
  AND U11101 ( .A(n468), .B(n11554), .Z(n11553) );
  XOR U11102 ( .A(n11555), .B(n11552), .Z(n11554) );
  XOR U11103 ( .A(n11556), .B(n11557), .Z(n11544) );
  AND U11104 ( .A(n11558), .B(n11559), .Z(n11557) );
  XOR U11105 ( .A(n11556), .B(n9745), .Z(n11559) );
  XOR U11106 ( .A(n11560), .B(n11561), .Z(n9745) );
  AND U11107 ( .A(n471), .B(n11562), .Z(n11561) );
  XOR U11108 ( .A(n11563), .B(n11560), .Z(n11562) );
  XNOR U11109 ( .A(n9742), .B(n11556), .Z(n11558) );
  XOR U11110 ( .A(n11564), .B(n11565), .Z(n9742) );
  AND U11111 ( .A(n468), .B(n11566), .Z(n11565) );
  XOR U11112 ( .A(n11567), .B(n11564), .Z(n11566) );
  XOR U11113 ( .A(n11568), .B(n11569), .Z(n11556) );
  AND U11114 ( .A(n11570), .B(n11571), .Z(n11569) );
  XOR U11115 ( .A(n11568), .B(n9757), .Z(n11571) );
  XOR U11116 ( .A(n11572), .B(n11573), .Z(n9757) );
  AND U11117 ( .A(n471), .B(n11574), .Z(n11573) );
  XOR U11118 ( .A(n11575), .B(n11572), .Z(n11574) );
  XNOR U11119 ( .A(n9754), .B(n11568), .Z(n11570) );
  XOR U11120 ( .A(n11576), .B(n11577), .Z(n9754) );
  AND U11121 ( .A(n468), .B(n11578), .Z(n11577) );
  XOR U11122 ( .A(n11579), .B(n11576), .Z(n11578) );
  XOR U11123 ( .A(n11580), .B(n11581), .Z(n11568) );
  AND U11124 ( .A(n11582), .B(n11583), .Z(n11581) );
  XOR U11125 ( .A(n11580), .B(n9769), .Z(n11583) );
  XOR U11126 ( .A(n11584), .B(n11585), .Z(n9769) );
  AND U11127 ( .A(n471), .B(n11586), .Z(n11585) );
  XOR U11128 ( .A(n11587), .B(n11584), .Z(n11586) );
  XNOR U11129 ( .A(n9766), .B(n11580), .Z(n11582) );
  XOR U11130 ( .A(n11588), .B(n11589), .Z(n9766) );
  AND U11131 ( .A(n468), .B(n11590), .Z(n11589) );
  XOR U11132 ( .A(n11591), .B(n11588), .Z(n11590) );
  XOR U11133 ( .A(n11592), .B(n11593), .Z(n11580) );
  AND U11134 ( .A(n11594), .B(n11595), .Z(n11593) );
  XOR U11135 ( .A(n11592), .B(n9781), .Z(n11595) );
  XOR U11136 ( .A(n11596), .B(n11597), .Z(n9781) );
  AND U11137 ( .A(n471), .B(n11598), .Z(n11597) );
  XOR U11138 ( .A(n11599), .B(n11596), .Z(n11598) );
  XNOR U11139 ( .A(n9778), .B(n11592), .Z(n11594) );
  XOR U11140 ( .A(n11600), .B(n11601), .Z(n9778) );
  AND U11141 ( .A(n468), .B(n11602), .Z(n11601) );
  XOR U11142 ( .A(n11603), .B(n11600), .Z(n11602) );
  XOR U11143 ( .A(n11604), .B(n11605), .Z(n11592) );
  AND U11144 ( .A(n11606), .B(n11607), .Z(n11605) );
  XOR U11145 ( .A(n11604), .B(n9793), .Z(n11607) );
  XOR U11146 ( .A(n11608), .B(n11609), .Z(n9793) );
  AND U11147 ( .A(n471), .B(n11610), .Z(n11609) );
  XOR U11148 ( .A(n11611), .B(n11608), .Z(n11610) );
  XNOR U11149 ( .A(n9790), .B(n11604), .Z(n11606) );
  XOR U11150 ( .A(n11612), .B(n11613), .Z(n9790) );
  AND U11151 ( .A(n468), .B(n11614), .Z(n11613) );
  XOR U11152 ( .A(n11615), .B(n11612), .Z(n11614) );
  XOR U11153 ( .A(n11616), .B(n11617), .Z(n11604) );
  AND U11154 ( .A(n11618), .B(n11619), .Z(n11617) );
  XOR U11155 ( .A(n11616), .B(n9805), .Z(n11619) );
  XOR U11156 ( .A(n11620), .B(n11621), .Z(n9805) );
  AND U11157 ( .A(n471), .B(n11622), .Z(n11621) );
  XOR U11158 ( .A(n11623), .B(n11620), .Z(n11622) );
  XNOR U11159 ( .A(n9802), .B(n11616), .Z(n11618) );
  XOR U11160 ( .A(n11624), .B(n11625), .Z(n9802) );
  AND U11161 ( .A(n468), .B(n11626), .Z(n11625) );
  XOR U11162 ( .A(n11627), .B(n11624), .Z(n11626) );
  XOR U11163 ( .A(n11628), .B(n11629), .Z(n11616) );
  AND U11164 ( .A(n11630), .B(n11631), .Z(n11629) );
  XOR U11165 ( .A(n11628), .B(n9817), .Z(n11631) );
  XOR U11166 ( .A(n11632), .B(n11633), .Z(n9817) );
  AND U11167 ( .A(n471), .B(n11634), .Z(n11633) );
  XOR U11168 ( .A(n11635), .B(n11632), .Z(n11634) );
  XNOR U11169 ( .A(n9814), .B(n11628), .Z(n11630) );
  XOR U11170 ( .A(n11636), .B(n11637), .Z(n9814) );
  AND U11171 ( .A(n468), .B(n11638), .Z(n11637) );
  XOR U11172 ( .A(n11639), .B(n11636), .Z(n11638) );
  XOR U11173 ( .A(n11640), .B(n11641), .Z(n11628) );
  AND U11174 ( .A(n11642), .B(n11643), .Z(n11641) );
  XOR U11175 ( .A(n11640), .B(n9829), .Z(n11643) );
  XOR U11176 ( .A(n11644), .B(n11645), .Z(n9829) );
  AND U11177 ( .A(n471), .B(n11646), .Z(n11645) );
  XOR U11178 ( .A(n11647), .B(n11644), .Z(n11646) );
  XNOR U11179 ( .A(n9826), .B(n11640), .Z(n11642) );
  XOR U11180 ( .A(n11648), .B(n11649), .Z(n9826) );
  AND U11181 ( .A(n468), .B(n11650), .Z(n11649) );
  XOR U11182 ( .A(n11651), .B(n11648), .Z(n11650) );
  XOR U11183 ( .A(n11652), .B(n11653), .Z(n11640) );
  AND U11184 ( .A(n11654), .B(n11655), .Z(n11653) );
  XOR U11185 ( .A(n11652), .B(n9841), .Z(n11655) );
  XOR U11186 ( .A(n11656), .B(n11657), .Z(n9841) );
  AND U11187 ( .A(n471), .B(n11658), .Z(n11657) );
  XOR U11188 ( .A(n11659), .B(n11656), .Z(n11658) );
  XNOR U11189 ( .A(n9838), .B(n11652), .Z(n11654) );
  XOR U11190 ( .A(n11660), .B(n11661), .Z(n9838) );
  AND U11191 ( .A(n468), .B(n11662), .Z(n11661) );
  XOR U11192 ( .A(n11663), .B(n11660), .Z(n11662) );
  XOR U11193 ( .A(n11664), .B(n11665), .Z(n11652) );
  AND U11194 ( .A(n11666), .B(n11667), .Z(n11665) );
  XOR U11195 ( .A(n11664), .B(n9853), .Z(n11667) );
  XOR U11196 ( .A(n11668), .B(n11669), .Z(n9853) );
  AND U11197 ( .A(n471), .B(n11670), .Z(n11669) );
  XOR U11198 ( .A(n11671), .B(n11668), .Z(n11670) );
  XNOR U11199 ( .A(n9850), .B(n11664), .Z(n11666) );
  XOR U11200 ( .A(n11672), .B(n11673), .Z(n9850) );
  AND U11201 ( .A(n468), .B(n11674), .Z(n11673) );
  XOR U11202 ( .A(n11675), .B(n11672), .Z(n11674) );
  XOR U11203 ( .A(n11676), .B(n11677), .Z(n11664) );
  AND U11204 ( .A(n11678), .B(n11679), .Z(n11677) );
  XOR U11205 ( .A(n11676), .B(n9865), .Z(n11679) );
  XOR U11206 ( .A(n11680), .B(n11681), .Z(n9865) );
  AND U11207 ( .A(n471), .B(n11682), .Z(n11681) );
  XOR U11208 ( .A(n11683), .B(n11680), .Z(n11682) );
  XNOR U11209 ( .A(n9862), .B(n11676), .Z(n11678) );
  XOR U11210 ( .A(n11684), .B(n11685), .Z(n9862) );
  AND U11211 ( .A(n468), .B(n11686), .Z(n11685) );
  XOR U11212 ( .A(n11687), .B(n11684), .Z(n11686) );
  XOR U11213 ( .A(n11688), .B(n11689), .Z(n11676) );
  AND U11214 ( .A(n11690), .B(n11691), .Z(n11689) );
  XOR U11215 ( .A(n11688), .B(n9877), .Z(n11691) );
  XOR U11216 ( .A(n11692), .B(n11693), .Z(n9877) );
  AND U11217 ( .A(n471), .B(n11694), .Z(n11693) );
  XOR U11218 ( .A(n11695), .B(n11692), .Z(n11694) );
  XNOR U11219 ( .A(n9874), .B(n11688), .Z(n11690) );
  XOR U11220 ( .A(n11696), .B(n11697), .Z(n9874) );
  AND U11221 ( .A(n468), .B(n11698), .Z(n11697) );
  XOR U11222 ( .A(n11699), .B(n11696), .Z(n11698) );
  XOR U11223 ( .A(n11700), .B(n11701), .Z(n11688) );
  AND U11224 ( .A(n11702), .B(n11703), .Z(n11701) );
  XOR U11225 ( .A(n11700), .B(n9889), .Z(n11703) );
  XOR U11226 ( .A(n11704), .B(n11705), .Z(n9889) );
  AND U11227 ( .A(n471), .B(n11706), .Z(n11705) );
  XOR U11228 ( .A(n11707), .B(n11704), .Z(n11706) );
  XNOR U11229 ( .A(n9886), .B(n11700), .Z(n11702) );
  XOR U11230 ( .A(n11708), .B(n11709), .Z(n9886) );
  AND U11231 ( .A(n468), .B(n11710), .Z(n11709) );
  XOR U11232 ( .A(n11711), .B(n11708), .Z(n11710) );
  XOR U11233 ( .A(n11712), .B(n11713), .Z(n11700) );
  AND U11234 ( .A(n11714), .B(n11715), .Z(n11713) );
  XOR U11235 ( .A(n11712), .B(n9901), .Z(n11715) );
  XOR U11236 ( .A(n11716), .B(n11717), .Z(n9901) );
  AND U11237 ( .A(n471), .B(n11718), .Z(n11717) );
  XOR U11238 ( .A(n11719), .B(n11716), .Z(n11718) );
  XNOR U11239 ( .A(n9898), .B(n11712), .Z(n11714) );
  XOR U11240 ( .A(n11720), .B(n11721), .Z(n9898) );
  AND U11241 ( .A(n468), .B(n11722), .Z(n11721) );
  XOR U11242 ( .A(n11723), .B(n11720), .Z(n11722) );
  XOR U11243 ( .A(n11724), .B(n11725), .Z(n11712) );
  AND U11244 ( .A(n11726), .B(n11727), .Z(n11725) );
  XOR U11245 ( .A(n11724), .B(n9913), .Z(n11727) );
  XOR U11246 ( .A(n11728), .B(n11729), .Z(n9913) );
  AND U11247 ( .A(n471), .B(n11730), .Z(n11729) );
  XOR U11248 ( .A(n11731), .B(n11728), .Z(n11730) );
  XNOR U11249 ( .A(n9910), .B(n11724), .Z(n11726) );
  XOR U11250 ( .A(n11732), .B(n11733), .Z(n9910) );
  AND U11251 ( .A(n468), .B(n11734), .Z(n11733) );
  XOR U11252 ( .A(n11735), .B(n11732), .Z(n11734) );
  XOR U11253 ( .A(n11736), .B(n11737), .Z(n11724) );
  AND U11254 ( .A(n11738), .B(n11739), .Z(n11737) );
  XOR U11255 ( .A(n11736), .B(n9925), .Z(n11739) );
  XOR U11256 ( .A(n11740), .B(n11741), .Z(n9925) );
  AND U11257 ( .A(n471), .B(n11742), .Z(n11741) );
  XOR U11258 ( .A(n11743), .B(n11740), .Z(n11742) );
  XNOR U11259 ( .A(n9922), .B(n11736), .Z(n11738) );
  XOR U11260 ( .A(n11744), .B(n11745), .Z(n9922) );
  AND U11261 ( .A(n468), .B(n11746), .Z(n11745) );
  XOR U11262 ( .A(n11747), .B(n11744), .Z(n11746) );
  XOR U11263 ( .A(n11748), .B(n11749), .Z(n11736) );
  AND U11264 ( .A(n11750), .B(n11751), .Z(n11749) );
  XNOR U11265 ( .A(n11752), .B(n9938), .Z(n11751) );
  XOR U11266 ( .A(n11753), .B(n11754), .Z(n9938) );
  AND U11267 ( .A(n471), .B(n11755), .Z(n11754) );
  XOR U11268 ( .A(n11753), .B(n11756), .Z(n11755) );
  XNOR U11269 ( .A(n9935), .B(n11748), .Z(n11750) );
  XOR U11270 ( .A(n11757), .B(n11758), .Z(n9935) );
  AND U11271 ( .A(n468), .B(n11759), .Z(n11758) );
  XOR U11272 ( .A(n11757), .B(n11760), .Z(n11759) );
  IV U11273 ( .A(n11752), .Z(n11748) );
  AND U11274 ( .A(n11384), .B(n11387), .Z(n11752) );
  XNOR U11275 ( .A(n11761), .B(n11762), .Z(n11387) );
  AND U11276 ( .A(n471), .B(n11763), .Z(n11762) );
  XNOR U11277 ( .A(n11764), .B(n11761), .Z(n11763) );
  XOR U11278 ( .A(n11765), .B(n11766), .Z(n471) );
  AND U11279 ( .A(n11767), .B(n11768), .Z(n11766) );
  XOR U11280 ( .A(n11395), .B(n11765), .Z(n11768) );
  IV U11281 ( .A(n11769), .Z(n11395) );
  AND U11282 ( .A(p_input[6911]), .B(p_input[6879]), .Z(n11769) );
  XOR U11283 ( .A(n11765), .B(n11392), .Z(n11767) );
  AND U11284 ( .A(p_input[6815]), .B(p_input[6847]), .Z(n11392) );
  XOR U11285 ( .A(n11770), .B(n11771), .Z(n11765) );
  AND U11286 ( .A(n11772), .B(n11773), .Z(n11771) );
  XOR U11287 ( .A(n11770), .B(n11407), .Z(n11773) );
  XNOR U11288 ( .A(p_input[6878]), .B(n11774), .Z(n11407) );
  AND U11289 ( .A(n259), .B(n11775), .Z(n11774) );
  XOR U11290 ( .A(p_input[6910]), .B(p_input[6878]), .Z(n11775) );
  XNOR U11291 ( .A(n11404), .B(n11770), .Z(n11772) );
  XOR U11292 ( .A(n11776), .B(n11777), .Z(n11404) );
  AND U11293 ( .A(n257), .B(n11778), .Z(n11777) );
  XOR U11294 ( .A(p_input[6846]), .B(p_input[6814]), .Z(n11778) );
  XOR U11295 ( .A(n11779), .B(n11780), .Z(n11770) );
  AND U11296 ( .A(n11781), .B(n11782), .Z(n11780) );
  XOR U11297 ( .A(n11779), .B(n11419), .Z(n11782) );
  XNOR U11298 ( .A(p_input[6877]), .B(n11783), .Z(n11419) );
  AND U11299 ( .A(n259), .B(n11784), .Z(n11783) );
  XOR U11300 ( .A(p_input[6909]), .B(p_input[6877]), .Z(n11784) );
  XNOR U11301 ( .A(n11416), .B(n11779), .Z(n11781) );
  XOR U11302 ( .A(n11785), .B(n11786), .Z(n11416) );
  AND U11303 ( .A(n257), .B(n11787), .Z(n11786) );
  XOR U11304 ( .A(p_input[6845]), .B(p_input[6813]), .Z(n11787) );
  XOR U11305 ( .A(n11788), .B(n11789), .Z(n11779) );
  AND U11306 ( .A(n11790), .B(n11791), .Z(n11789) );
  XOR U11307 ( .A(n11788), .B(n11431), .Z(n11791) );
  XNOR U11308 ( .A(p_input[6876]), .B(n11792), .Z(n11431) );
  AND U11309 ( .A(n259), .B(n11793), .Z(n11792) );
  XOR U11310 ( .A(p_input[6908]), .B(p_input[6876]), .Z(n11793) );
  XNOR U11311 ( .A(n11428), .B(n11788), .Z(n11790) );
  XOR U11312 ( .A(n11794), .B(n11795), .Z(n11428) );
  AND U11313 ( .A(n257), .B(n11796), .Z(n11795) );
  XOR U11314 ( .A(p_input[6844]), .B(p_input[6812]), .Z(n11796) );
  XOR U11315 ( .A(n11797), .B(n11798), .Z(n11788) );
  AND U11316 ( .A(n11799), .B(n11800), .Z(n11798) );
  XOR U11317 ( .A(n11797), .B(n11443), .Z(n11800) );
  XNOR U11318 ( .A(p_input[6875]), .B(n11801), .Z(n11443) );
  AND U11319 ( .A(n259), .B(n11802), .Z(n11801) );
  XOR U11320 ( .A(p_input[6907]), .B(p_input[6875]), .Z(n11802) );
  XNOR U11321 ( .A(n11440), .B(n11797), .Z(n11799) );
  XOR U11322 ( .A(n11803), .B(n11804), .Z(n11440) );
  AND U11323 ( .A(n257), .B(n11805), .Z(n11804) );
  XOR U11324 ( .A(p_input[6843]), .B(p_input[6811]), .Z(n11805) );
  XOR U11325 ( .A(n11806), .B(n11807), .Z(n11797) );
  AND U11326 ( .A(n11808), .B(n11809), .Z(n11807) );
  XOR U11327 ( .A(n11806), .B(n11455), .Z(n11809) );
  XNOR U11328 ( .A(p_input[6874]), .B(n11810), .Z(n11455) );
  AND U11329 ( .A(n259), .B(n11811), .Z(n11810) );
  XOR U11330 ( .A(p_input[6906]), .B(p_input[6874]), .Z(n11811) );
  XNOR U11331 ( .A(n11452), .B(n11806), .Z(n11808) );
  XOR U11332 ( .A(n11812), .B(n11813), .Z(n11452) );
  AND U11333 ( .A(n257), .B(n11814), .Z(n11813) );
  XOR U11334 ( .A(p_input[6842]), .B(p_input[6810]), .Z(n11814) );
  XOR U11335 ( .A(n11815), .B(n11816), .Z(n11806) );
  AND U11336 ( .A(n11817), .B(n11818), .Z(n11816) );
  XOR U11337 ( .A(n11815), .B(n11467), .Z(n11818) );
  XNOR U11338 ( .A(p_input[6873]), .B(n11819), .Z(n11467) );
  AND U11339 ( .A(n259), .B(n11820), .Z(n11819) );
  XOR U11340 ( .A(p_input[6905]), .B(p_input[6873]), .Z(n11820) );
  XNOR U11341 ( .A(n11464), .B(n11815), .Z(n11817) );
  XOR U11342 ( .A(n11821), .B(n11822), .Z(n11464) );
  AND U11343 ( .A(n257), .B(n11823), .Z(n11822) );
  XOR U11344 ( .A(p_input[6841]), .B(p_input[6809]), .Z(n11823) );
  XOR U11345 ( .A(n11824), .B(n11825), .Z(n11815) );
  AND U11346 ( .A(n11826), .B(n11827), .Z(n11825) );
  XOR U11347 ( .A(n11824), .B(n11479), .Z(n11827) );
  XNOR U11348 ( .A(p_input[6872]), .B(n11828), .Z(n11479) );
  AND U11349 ( .A(n259), .B(n11829), .Z(n11828) );
  XOR U11350 ( .A(p_input[6904]), .B(p_input[6872]), .Z(n11829) );
  XNOR U11351 ( .A(n11476), .B(n11824), .Z(n11826) );
  XOR U11352 ( .A(n11830), .B(n11831), .Z(n11476) );
  AND U11353 ( .A(n257), .B(n11832), .Z(n11831) );
  XOR U11354 ( .A(p_input[6840]), .B(p_input[6808]), .Z(n11832) );
  XOR U11355 ( .A(n11833), .B(n11834), .Z(n11824) );
  AND U11356 ( .A(n11835), .B(n11836), .Z(n11834) );
  XOR U11357 ( .A(n11833), .B(n11491), .Z(n11836) );
  XNOR U11358 ( .A(p_input[6871]), .B(n11837), .Z(n11491) );
  AND U11359 ( .A(n259), .B(n11838), .Z(n11837) );
  XOR U11360 ( .A(p_input[6903]), .B(p_input[6871]), .Z(n11838) );
  XNOR U11361 ( .A(n11488), .B(n11833), .Z(n11835) );
  XOR U11362 ( .A(n11839), .B(n11840), .Z(n11488) );
  AND U11363 ( .A(n257), .B(n11841), .Z(n11840) );
  XOR U11364 ( .A(p_input[6839]), .B(p_input[6807]), .Z(n11841) );
  XOR U11365 ( .A(n11842), .B(n11843), .Z(n11833) );
  AND U11366 ( .A(n11844), .B(n11845), .Z(n11843) );
  XOR U11367 ( .A(n11842), .B(n11503), .Z(n11845) );
  XNOR U11368 ( .A(p_input[6870]), .B(n11846), .Z(n11503) );
  AND U11369 ( .A(n259), .B(n11847), .Z(n11846) );
  XOR U11370 ( .A(p_input[6902]), .B(p_input[6870]), .Z(n11847) );
  XNOR U11371 ( .A(n11500), .B(n11842), .Z(n11844) );
  XOR U11372 ( .A(n11848), .B(n11849), .Z(n11500) );
  AND U11373 ( .A(n257), .B(n11850), .Z(n11849) );
  XOR U11374 ( .A(p_input[6838]), .B(p_input[6806]), .Z(n11850) );
  XOR U11375 ( .A(n11851), .B(n11852), .Z(n11842) );
  AND U11376 ( .A(n11853), .B(n11854), .Z(n11852) );
  XOR U11377 ( .A(n11851), .B(n11515), .Z(n11854) );
  XNOR U11378 ( .A(p_input[6869]), .B(n11855), .Z(n11515) );
  AND U11379 ( .A(n259), .B(n11856), .Z(n11855) );
  XOR U11380 ( .A(p_input[6901]), .B(p_input[6869]), .Z(n11856) );
  XNOR U11381 ( .A(n11512), .B(n11851), .Z(n11853) );
  XOR U11382 ( .A(n11857), .B(n11858), .Z(n11512) );
  AND U11383 ( .A(n257), .B(n11859), .Z(n11858) );
  XOR U11384 ( .A(p_input[6837]), .B(p_input[6805]), .Z(n11859) );
  XOR U11385 ( .A(n11860), .B(n11861), .Z(n11851) );
  AND U11386 ( .A(n11862), .B(n11863), .Z(n11861) );
  XOR U11387 ( .A(n11860), .B(n11527), .Z(n11863) );
  XNOR U11388 ( .A(p_input[6868]), .B(n11864), .Z(n11527) );
  AND U11389 ( .A(n259), .B(n11865), .Z(n11864) );
  XOR U11390 ( .A(p_input[6900]), .B(p_input[6868]), .Z(n11865) );
  XNOR U11391 ( .A(n11524), .B(n11860), .Z(n11862) );
  XOR U11392 ( .A(n11866), .B(n11867), .Z(n11524) );
  AND U11393 ( .A(n257), .B(n11868), .Z(n11867) );
  XOR U11394 ( .A(p_input[6836]), .B(p_input[6804]), .Z(n11868) );
  XOR U11395 ( .A(n11869), .B(n11870), .Z(n11860) );
  AND U11396 ( .A(n11871), .B(n11872), .Z(n11870) );
  XOR U11397 ( .A(n11869), .B(n11539), .Z(n11872) );
  XNOR U11398 ( .A(p_input[6867]), .B(n11873), .Z(n11539) );
  AND U11399 ( .A(n259), .B(n11874), .Z(n11873) );
  XOR U11400 ( .A(p_input[6899]), .B(p_input[6867]), .Z(n11874) );
  XNOR U11401 ( .A(n11536), .B(n11869), .Z(n11871) );
  XOR U11402 ( .A(n11875), .B(n11876), .Z(n11536) );
  AND U11403 ( .A(n257), .B(n11877), .Z(n11876) );
  XOR U11404 ( .A(p_input[6835]), .B(p_input[6803]), .Z(n11877) );
  XOR U11405 ( .A(n11878), .B(n11879), .Z(n11869) );
  AND U11406 ( .A(n11880), .B(n11881), .Z(n11879) );
  XOR U11407 ( .A(n11878), .B(n11551), .Z(n11881) );
  XNOR U11408 ( .A(p_input[6866]), .B(n11882), .Z(n11551) );
  AND U11409 ( .A(n259), .B(n11883), .Z(n11882) );
  XOR U11410 ( .A(p_input[6898]), .B(p_input[6866]), .Z(n11883) );
  XNOR U11411 ( .A(n11548), .B(n11878), .Z(n11880) );
  XOR U11412 ( .A(n11884), .B(n11885), .Z(n11548) );
  AND U11413 ( .A(n257), .B(n11886), .Z(n11885) );
  XOR U11414 ( .A(p_input[6834]), .B(p_input[6802]), .Z(n11886) );
  XOR U11415 ( .A(n11887), .B(n11888), .Z(n11878) );
  AND U11416 ( .A(n11889), .B(n11890), .Z(n11888) );
  XOR U11417 ( .A(n11887), .B(n11563), .Z(n11890) );
  XNOR U11418 ( .A(p_input[6865]), .B(n11891), .Z(n11563) );
  AND U11419 ( .A(n259), .B(n11892), .Z(n11891) );
  XOR U11420 ( .A(p_input[6897]), .B(p_input[6865]), .Z(n11892) );
  XNOR U11421 ( .A(n11560), .B(n11887), .Z(n11889) );
  XOR U11422 ( .A(n11893), .B(n11894), .Z(n11560) );
  AND U11423 ( .A(n257), .B(n11895), .Z(n11894) );
  XOR U11424 ( .A(p_input[6833]), .B(p_input[6801]), .Z(n11895) );
  XOR U11425 ( .A(n11896), .B(n11897), .Z(n11887) );
  AND U11426 ( .A(n11898), .B(n11899), .Z(n11897) );
  XOR U11427 ( .A(n11896), .B(n11575), .Z(n11899) );
  XNOR U11428 ( .A(p_input[6864]), .B(n11900), .Z(n11575) );
  AND U11429 ( .A(n259), .B(n11901), .Z(n11900) );
  XOR U11430 ( .A(p_input[6896]), .B(p_input[6864]), .Z(n11901) );
  XNOR U11431 ( .A(n11572), .B(n11896), .Z(n11898) );
  XOR U11432 ( .A(n11902), .B(n11903), .Z(n11572) );
  AND U11433 ( .A(n257), .B(n11904), .Z(n11903) );
  XOR U11434 ( .A(p_input[6832]), .B(p_input[6800]), .Z(n11904) );
  XOR U11435 ( .A(n11905), .B(n11906), .Z(n11896) );
  AND U11436 ( .A(n11907), .B(n11908), .Z(n11906) );
  XOR U11437 ( .A(n11905), .B(n11587), .Z(n11908) );
  XNOR U11438 ( .A(p_input[6863]), .B(n11909), .Z(n11587) );
  AND U11439 ( .A(n259), .B(n11910), .Z(n11909) );
  XOR U11440 ( .A(p_input[6895]), .B(p_input[6863]), .Z(n11910) );
  XNOR U11441 ( .A(n11584), .B(n11905), .Z(n11907) );
  XOR U11442 ( .A(n11911), .B(n11912), .Z(n11584) );
  AND U11443 ( .A(n257), .B(n11913), .Z(n11912) );
  XOR U11444 ( .A(p_input[6831]), .B(p_input[6799]), .Z(n11913) );
  XOR U11445 ( .A(n11914), .B(n11915), .Z(n11905) );
  AND U11446 ( .A(n11916), .B(n11917), .Z(n11915) );
  XOR U11447 ( .A(n11914), .B(n11599), .Z(n11917) );
  XNOR U11448 ( .A(p_input[6862]), .B(n11918), .Z(n11599) );
  AND U11449 ( .A(n259), .B(n11919), .Z(n11918) );
  XOR U11450 ( .A(p_input[6894]), .B(p_input[6862]), .Z(n11919) );
  XNOR U11451 ( .A(n11596), .B(n11914), .Z(n11916) );
  XOR U11452 ( .A(n11920), .B(n11921), .Z(n11596) );
  AND U11453 ( .A(n257), .B(n11922), .Z(n11921) );
  XOR U11454 ( .A(p_input[6830]), .B(p_input[6798]), .Z(n11922) );
  XOR U11455 ( .A(n11923), .B(n11924), .Z(n11914) );
  AND U11456 ( .A(n11925), .B(n11926), .Z(n11924) );
  XOR U11457 ( .A(n11923), .B(n11611), .Z(n11926) );
  XNOR U11458 ( .A(p_input[6861]), .B(n11927), .Z(n11611) );
  AND U11459 ( .A(n259), .B(n11928), .Z(n11927) );
  XOR U11460 ( .A(p_input[6893]), .B(p_input[6861]), .Z(n11928) );
  XNOR U11461 ( .A(n11608), .B(n11923), .Z(n11925) );
  XOR U11462 ( .A(n11929), .B(n11930), .Z(n11608) );
  AND U11463 ( .A(n257), .B(n11931), .Z(n11930) );
  XOR U11464 ( .A(p_input[6829]), .B(p_input[6797]), .Z(n11931) );
  XOR U11465 ( .A(n11932), .B(n11933), .Z(n11923) );
  AND U11466 ( .A(n11934), .B(n11935), .Z(n11933) );
  XOR U11467 ( .A(n11932), .B(n11623), .Z(n11935) );
  XNOR U11468 ( .A(p_input[6860]), .B(n11936), .Z(n11623) );
  AND U11469 ( .A(n259), .B(n11937), .Z(n11936) );
  XOR U11470 ( .A(p_input[6892]), .B(p_input[6860]), .Z(n11937) );
  XNOR U11471 ( .A(n11620), .B(n11932), .Z(n11934) );
  XOR U11472 ( .A(n11938), .B(n11939), .Z(n11620) );
  AND U11473 ( .A(n257), .B(n11940), .Z(n11939) );
  XOR U11474 ( .A(p_input[6828]), .B(p_input[6796]), .Z(n11940) );
  XOR U11475 ( .A(n11941), .B(n11942), .Z(n11932) );
  AND U11476 ( .A(n11943), .B(n11944), .Z(n11942) );
  XOR U11477 ( .A(n11941), .B(n11635), .Z(n11944) );
  XNOR U11478 ( .A(p_input[6859]), .B(n11945), .Z(n11635) );
  AND U11479 ( .A(n259), .B(n11946), .Z(n11945) );
  XOR U11480 ( .A(p_input[6891]), .B(p_input[6859]), .Z(n11946) );
  XNOR U11481 ( .A(n11632), .B(n11941), .Z(n11943) );
  XOR U11482 ( .A(n11947), .B(n11948), .Z(n11632) );
  AND U11483 ( .A(n257), .B(n11949), .Z(n11948) );
  XOR U11484 ( .A(p_input[6827]), .B(p_input[6795]), .Z(n11949) );
  XOR U11485 ( .A(n11950), .B(n11951), .Z(n11941) );
  AND U11486 ( .A(n11952), .B(n11953), .Z(n11951) );
  XOR U11487 ( .A(n11950), .B(n11647), .Z(n11953) );
  XNOR U11488 ( .A(p_input[6858]), .B(n11954), .Z(n11647) );
  AND U11489 ( .A(n259), .B(n11955), .Z(n11954) );
  XOR U11490 ( .A(p_input[6890]), .B(p_input[6858]), .Z(n11955) );
  XNOR U11491 ( .A(n11644), .B(n11950), .Z(n11952) );
  XOR U11492 ( .A(n11956), .B(n11957), .Z(n11644) );
  AND U11493 ( .A(n257), .B(n11958), .Z(n11957) );
  XOR U11494 ( .A(p_input[6826]), .B(p_input[6794]), .Z(n11958) );
  XOR U11495 ( .A(n11959), .B(n11960), .Z(n11950) );
  AND U11496 ( .A(n11961), .B(n11962), .Z(n11960) );
  XOR U11497 ( .A(n11959), .B(n11659), .Z(n11962) );
  XNOR U11498 ( .A(p_input[6857]), .B(n11963), .Z(n11659) );
  AND U11499 ( .A(n259), .B(n11964), .Z(n11963) );
  XOR U11500 ( .A(p_input[6889]), .B(p_input[6857]), .Z(n11964) );
  XNOR U11501 ( .A(n11656), .B(n11959), .Z(n11961) );
  XOR U11502 ( .A(n11965), .B(n11966), .Z(n11656) );
  AND U11503 ( .A(n257), .B(n11967), .Z(n11966) );
  XOR U11504 ( .A(p_input[6825]), .B(p_input[6793]), .Z(n11967) );
  XOR U11505 ( .A(n11968), .B(n11969), .Z(n11959) );
  AND U11506 ( .A(n11970), .B(n11971), .Z(n11969) );
  XOR U11507 ( .A(n11968), .B(n11671), .Z(n11971) );
  XNOR U11508 ( .A(p_input[6856]), .B(n11972), .Z(n11671) );
  AND U11509 ( .A(n259), .B(n11973), .Z(n11972) );
  XOR U11510 ( .A(p_input[6888]), .B(p_input[6856]), .Z(n11973) );
  XNOR U11511 ( .A(n11668), .B(n11968), .Z(n11970) );
  XOR U11512 ( .A(n11974), .B(n11975), .Z(n11668) );
  AND U11513 ( .A(n257), .B(n11976), .Z(n11975) );
  XOR U11514 ( .A(p_input[6824]), .B(p_input[6792]), .Z(n11976) );
  XOR U11515 ( .A(n11977), .B(n11978), .Z(n11968) );
  AND U11516 ( .A(n11979), .B(n11980), .Z(n11978) );
  XOR U11517 ( .A(n11977), .B(n11683), .Z(n11980) );
  XNOR U11518 ( .A(p_input[6855]), .B(n11981), .Z(n11683) );
  AND U11519 ( .A(n259), .B(n11982), .Z(n11981) );
  XOR U11520 ( .A(p_input[6887]), .B(p_input[6855]), .Z(n11982) );
  XNOR U11521 ( .A(n11680), .B(n11977), .Z(n11979) );
  XOR U11522 ( .A(n11983), .B(n11984), .Z(n11680) );
  AND U11523 ( .A(n257), .B(n11985), .Z(n11984) );
  XOR U11524 ( .A(p_input[6823]), .B(p_input[6791]), .Z(n11985) );
  XOR U11525 ( .A(n11986), .B(n11987), .Z(n11977) );
  AND U11526 ( .A(n11988), .B(n11989), .Z(n11987) );
  XOR U11527 ( .A(n11986), .B(n11695), .Z(n11989) );
  XNOR U11528 ( .A(p_input[6854]), .B(n11990), .Z(n11695) );
  AND U11529 ( .A(n259), .B(n11991), .Z(n11990) );
  XOR U11530 ( .A(p_input[6886]), .B(p_input[6854]), .Z(n11991) );
  XNOR U11531 ( .A(n11692), .B(n11986), .Z(n11988) );
  XOR U11532 ( .A(n11992), .B(n11993), .Z(n11692) );
  AND U11533 ( .A(n257), .B(n11994), .Z(n11993) );
  XOR U11534 ( .A(p_input[6822]), .B(p_input[6790]), .Z(n11994) );
  XOR U11535 ( .A(n11995), .B(n11996), .Z(n11986) );
  AND U11536 ( .A(n11997), .B(n11998), .Z(n11996) );
  XOR U11537 ( .A(n11995), .B(n11707), .Z(n11998) );
  XNOR U11538 ( .A(p_input[6853]), .B(n11999), .Z(n11707) );
  AND U11539 ( .A(n259), .B(n12000), .Z(n11999) );
  XOR U11540 ( .A(p_input[6885]), .B(p_input[6853]), .Z(n12000) );
  XNOR U11541 ( .A(n11704), .B(n11995), .Z(n11997) );
  XOR U11542 ( .A(n12001), .B(n12002), .Z(n11704) );
  AND U11543 ( .A(n257), .B(n12003), .Z(n12002) );
  XOR U11544 ( .A(p_input[6821]), .B(p_input[6789]), .Z(n12003) );
  XOR U11545 ( .A(n12004), .B(n12005), .Z(n11995) );
  AND U11546 ( .A(n12006), .B(n12007), .Z(n12005) );
  XOR U11547 ( .A(n12004), .B(n11719), .Z(n12007) );
  XNOR U11548 ( .A(p_input[6852]), .B(n12008), .Z(n11719) );
  AND U11549 ( .A(n259), .B(n12009), .Z(n12008) );
  XOR U11550 ( .A(p_input[6884]), .B(p_input[6852]), .Z(n12009) );
  XNOR U11551 ( .A(n11716), .B(n12004), .Z(n12006) );
  XOR U11552 ( .A(n12010), .B(n12011), .Z(n11716) );
  AND U11553 ( .A(n257), .B(n12012), .Z(n12011) );
  XOR U11554 ( .A(p_input[6820]), .B(p_input[6788]), .Z(n12012) );
  XOR U11555 ( .A(n12013), .B(n12014), .Z(n12004) );
  AND U11556 ( .A(n12015), .B(n12016), .Z(n12014) );
  XOR U11557 ( .A(n12013), .B(n11731), .Z(n12016) );
  XNOR U11558 ( .A(p_input[6851]), .B(n12017), .Z(n11731) );
  AND U11559 ( .A(n259), .B(n12018), .Z(n12017) );
  XOR U11560 ( .A(p_input[6883]), .B(p_input[6851]), .Z(n12018) );
  XNOR U11561 ( .A(n11728), .B(n12013), .Z(n12015) );
  XOR U11562 ( .A(n12019), .B(n12020), .Z(n11728) );
  AND U11563 ( .A(n257), .B(n12021), .Z(n12020) );
  XOR U11564 ( .A(p_input[6819]), .B(p_input[6787]), .Z(n12021) );
  XOR U11565 ( .A(n12022), .B(n12023), .Z(n12013) );
  AND U11566 ( .A(n12024), .B(n12025), .Z(n12023) );
  XOR U11567 ( .A(n12022), .B(n11743), .Z(n12025) );
  XNOR U11568 ( .A(p_input[6850]), .B(n12026), .Z(n11743) );
  AND U11569 ( .A(n259), .B(n12027), .Z(n12026) );
  XOR U11570 ( .A(p_input[6882]), .B(p_input[6850]), .Z(n12027) );
  XNOR U11571 ( .A(n11740), .B(n12022), .Z(n12024) );
  XOR U11572 ( .A(n12028), .B(n12029), .Z(n11740) );
  AND U11573 ( .A(n257), .B(n12030), .Z(n12029) );
  XOR U11574 ( .A(p_input[6818]), .B(p_input[6786]), .Z(n12030) );
  XOR U11575 ( .A(n12031), .B(n12032), .Z(n12022) );
  AND U11576 ( .A(n12033), .B(n12034), .Z(n12032) );
  XNOR U11577 ( .A(n12035), .B(n11756), .Z(n12034) );
  XNOR U11578 ( .A(p_input[6849]), .B(n12036), .Z(n11756) );
  AND U11579 ( .A(n259), .B(n12037), .Z(n12036) );
  XNOR U11580 ( .A(p_input[6881]), .B(n12038), .Z(n12037) );
  IV U11581 ( .A(p_input[6849]), .Z(n12038) );
  XNOR U11582 ( .A(n11753), .B(n12031), .Z(n12033) );
  XNOR U11583 ( .A(p_input[6785]), .B(n12039), .Z(n11753) );
  AND U11584 ( .A(n257), .B(n12040), .Z(n12039) );
  XOR U11585 ( .A(p_input[6817]), .B(p_input[6785]), .Z(n12040) );
  IV U11586 ( .A(n12035), .Z(n12031) );
  AND U11587 ( .A(n11761), .B(n11764), .Z(n12035) );
  XOR U11588 ( .A(p_input[6848]), .B(n12041), .Z(n11764) );
  AND U11589 ( .A(n259), .B(n12042), .Z(n12041) );
  XOR U11590 ( .A(p_input[6880]), .B(p_input[6848]), .Z(n12042) );
  XOR U11591 ( .A(n12043), .B(n12044), .Z(n259) );
  AND U11592 ( .A(n12045), .B(n12046), .Z(n12044) );
  XNOR U11593 ( .A(p_input[6911]), .B(n12043), .Z(n12046) );
  XOR U11594 ( .A(n12043), .B(p_input[6879]), .Z(n12045) );
  XOR U11595 ( .A(n12047), .B(n12048), .Z(n12043) );
  AND U11596 ( .A(n12049), .B(n12050), .Z(n12048) );
  XNOR U11597 ( .A(p_input[6910]), .B(n12047), .Z(n12050) );
  XOR U11598 ( .A(n12047), .B(p_input[6878]), .Z(n12049) );
  XOR U11599 ( .A(n12051), .B(n12052), .Z(n12047) );
  AND U11600 ( .A(n12053), .B(n12054), .Z(n12052) );
  XNOR U11601 ( .A(p_input[6909]), .B(n12051), .Z(n12054) );
  XOR U11602 ( .A(n12051), .B(p_input[6877]), .Z(n12053) );
  XOR U11603 ( .A(n12055), .B(n12056), .Z(n12051) );
  AND U11604 ( .A(n12057), .B(n12058), .Z(n12056) );
  XNOR U11605 ( .A(p_input[6908]), .B(n12055), .Z(n12058) );
  XOR U11606 ( .A(n12055), .B(p_input[6876]), .Z(n12057) );
  XOR U11607 ( .A(n12059), .B(n12060), .Z(n12055) );
  AND U11608 ( .A(n12061), .B(n12062), .Z(n12060) );
  XNOR U11609 ( .A(p_input[6907]), .B(n12059), .Z(n12062) );
  XOR U11610 ( .A(n12059), .B(p_input[6875]), .Z(n12061) );
  XOR U11611 ( .A(n12063), .B(n12064), .Z(n12059) );
  AND U11612 ( .A(n12065), .B(n12066), .Z(n12064) );
  XNOR U11613 ( .A(p_input[6906]), .B(n12063), .Z(n12066) );
  XOR U11614 ( .A(n12063), .B(p_input[6874]), .Z(n12065) );
  XOR U11615 ( .A(n12067), .B(n12068), .Z(n12063) );
  AND U11616 ( .A(n12069), .B(n12070), .Z(n12068) );
  XNOR U11617 ( .A(p_input[6905]), .B(n12067), .Z(n12070) );
  XOR U11618 ( .A(n12067), .B(p_input[6873]), .Z(n12069) );
  XOR U11619 ( .A(n12071), .B(n12072), .Z(n12067) );
  AND U11620 ( .A(n12073), .B(n12074), .Z(n12072) );
  XNOR U11621 ( .A(p_input[6904]), .B(n12071), .Z(n12074) );
  XOR U11622 ( .A(n12071), .B(p_input[6872]), .Z(n12073) );
  XOR U11623 ( .A(n12075), .B(n12076), .Z(n12071) );
  AND U11624 ( .A(n12077), .B(n12078), .Z(n12076) );
  XNOR U11625 ( .A(p_input[6903]), .B(n12075), .Z(n12078) );
  XOR U11626 ( .A(n12075), .B(p_input[6871]), .Z(n12077) );
  XOR U11627 ( .A(n12079), .B(n12080), .Z(n12075) );
  AND U11628 ( .A(n12081), .B(n12082), .Z(n12080) );
  XNOR U11629 ( .A(p_input[6902]), .B(n12079), .Z(n12082) );
  XOR U11630 ( .A(n12079), .B(p_input[6870]), .Z(n12081) );
  XOR U11631 ( .A(n12083), .B(n12084), .Z(n12079) );
  AND U11632 ( .A(n12085), .B(n12086), .Z(n12084) );
  XNOR U11633 ( .A(p_input[6901]), .B(n12083), .Z(n12086) );
  XOR U11634 ( .A(n12083), .B(p_input[6869]), .Z(n12085) );
  XOR U11635 ( .A(n12087), .B(n12088), .Z(n12083) );
  AND U11636 ( .A(n12089), .B(n12090), .Z(n12088) );
  XNOR U11637 ( .A(p_input[6900]), .B(n12087), .Z(n12090) );
  XOR U11638 ( .A(n12087), .B(p_input[6868]), .Z(n12089) );
  XOR U11639 ( .A(n12091), .B(n12092), .Z(n12087) );
  AND U11640 ( .A(n12093), .B(n12094), .Z(n12092) );
  XNOR U11641 ( .A(p_input[6899]), .B(n12091), .Z(n12094) );
  XOR U11642 ( .A(n12091), .B(p_input[6867]), .Z(n12093) );
  XOR U11643 ( .A(n12095), .B(n12096), .Z(n12091) );
  AND U11644 ( .A(n12097), .B(n12098), .Z(n12096) );
  XNOR U11645 ( .A(p_input[6898]), .B(n12095), .Z(n12098) );
  XOR U11646 ( .A(n12095), .B(p_input[6866]), .Z(n12097) );
  XOR U11647 ( .A(n12099), .B(n12100), .Z(n12095) );
  AND U11648 ( .A(n12101), .B(n12102), .Z(n12100) );
  XNOR U11649 ( .A(p_input[6897]), .B(n12099), .Z(n12102) );
  XOR U11650 ( .A(n12099), .B(p_input[6865]), .Z(n12101) );
  XOR U11651 ( .A(n12103), .B(n12104), .Z(n12099) );
  AND U11652 ( .A(n12105), .B(n12106), .Z(n12104) );
  XNOR U11653 ( .A(p_input[6896]), .B(n12103), .Z(n12106) );
  XOR U11654 ( .A(n12103), .B(p_input[6864]), .Z(n12105) );
  XOR U11655 ( .A(n12107), .B(n12108), .Z(n12103) );
  AND U11656 ( .A(n12109), .B(n12110), .Z(n12108) );
  XNOR U11657 ( .A(p_input[6895]), .B(n12107), .Z(n12110) );
  XOR U11658 ( .A(n12107), .B(p_input[6863]), .Z(n12109) );
  XOR U11659 ( .A(n12111), .B(n12112), .Z(n12107) );
  AND U11660 ( .A(n12113), .B(n12114), .Z(n12112) );
  XNOR U11661 ( .A(p_input[6894]), .B(n12111), .Z(n12114) );
  XOR U11662 ( .A(n12111), .B(p_input[6862]), .Z(n12113) );
  XOR U11663 ( .A(n12115), .B(n12116), .Z(n12111) );
  AND U11664 ( .A(n12117), .B(n12118), .Z(n12116) );
  XNOR U11665 ( .A(p_input[6893]), .B(n12115), .Z(n12118) );
  XOR U11666 ( .A(n12115), .B(p_input[6861]), .Z(n12117) );
  XOR U11667 ( .A(n12119), .B(n12120), .Z(n12115) );
  AND U11668 ( .A(n12121), .B(n12122), .Z(n12120) );
  XNOR U11669 ( .A(p_input[6892]), .B(n12119), .Z(n12122) );
  XOR U11670 ( .A(n12119), .B(p_input[6860]), .Z(n12121) );
  XOR U11671 ( .A(n12123), .B(n12124), .Z(n12119) );
  AND U11672 ( .A(n12125), .B(n12126), .Z(n12124) );
  XNOR U11673 ( .A(p_input[6891]), .B(n12123), .Z(n12126) );
  XOR U11674 ( .A(n12123), .B(p_input[6859]), .Z(n12125) );
  XOR U11675 ( .A(n12127), .B(n12128), .Z(n12123) );
  AND U11676 ( .A(n12129), .B(n12130), .Z(n12128) );
  XNOR U11677 ( .A(p_input[6890]), .B(n12127), .Z(n12130) );
  XOR U11678 ( .A(n12127), .B(p_input[6858]), .Z(n12129) );
  XOR U11679 ( .A(n12131), .B(n12132), .Z(n12127) );
  AND U11680 ( .A(n12133), .B(n12134), .Z(n12132) );
  XNOR U11681 ( .A(p_input[6889]), .B(n12131), .Z(n12134) );
  XOR U11682 ( .A(n12131), .B(p_input[6857]), .Z(n12133) );
  XOR U11683 ( .A(n12135), .B(n12136), .Z(n12131) );
  AND U11684 ( .A(n12137), .B(n12138), .Z(n12136) );
  XNOR U11685 ( .A(p_input[6888]), .B(n12135), .Z(n12138) );
  XOR U11686 ( .A(n12135), .B(p_input[6856]), .Z(n12137) );
  XOR U11687 ( .A(n12139), .B(n12140), .Z(n12135) );
  AND U11688 ( .A(n12141), .B(n12142), .Z(n12140) );
  XNOR U11689 ( .A(p_input[6887]), .B(n12139), .Z(n12142) );
  XOR U11690 ( .A(n12139), .B(p_input[6855]), .Z(n12141) );
  XOR U11691 ( .A(n12143), .B(n12144), .Z(n12139) );
  AND U11692 ( .A(n12145), .B(n12146), .Z(n12144) );
  XNOR U11693 ( .A(p_input[6886]), .B(n12143), .Z(n12146) );
  XOR U11694 ( .A(n12143), .B(p_input[6854]), .Z(n12145) );
  XOR U11695 ( .A(n12147), .B(n12148), .Z(n12143) );
  AND U11696 ( .A(n12149), .B(n12150), .Z(n12148) );
  XNOR U11697 ( .A(p_input[6885]), .B(n12147), .Z(n12150) );
  XOR U11698 ( .A(n12147), .B(p_input[6853]), .Z(n12149) );
  XOR U11699 ( .A(n12151), .B(n12152), .Z(n12147) );
  AND U11700 ( .A(n12153), .B(n12154), .Z(n12152) );
  XNOR U11701 ( .A(p_input[6884]), .B(n12151), .Z(n12154) );
  XOR U11702 ( .A(n12151), .B(p_input[6852]), .Z(n12153) );
  XOR U11703 ( .A(n12155), .B(n12156), .Z(n12151) );
  AND U11704 ( .A(n12157), .B(n12158), .Z(n12156) );
  XNOR U11705 ( .A(p_input[6883]), .B(n12155), .Z(n12158) );
  XOR U11706 ( .A(n12155), .B(p_input[6851]), .Z(n12157) );
  XOR U11707 ( .A(n12159), .B(n12160), .Z(n12155) );
  AND U11708 ( .A(n12161), .B(n12162), .Z(n12160) );
  XNOR U11709 ( .A(p_input[6882]), .B(n12159), .Z(n12162) );
  XOR U11710 ( .A(n12159), .B(p_input[6850]), .Z(n12161) );
  XNOR U11711 ( .A(n12163), .B(n12164), .Z(n12159) );
  AND U11712 ( .A(n12165), .B(n12166), .Z(n12164) );
  XOR U11713 ( .A(p_input[6881]), .B(n12163), .Z(n12166) );
  XNOR U11714 ( .A(p_input[6849]), .B(n12163), .Z(n12165) );
  AND U11715 ( .A(p_input[6880]), .B(n12167), .Z(n12163) );
  IV U11716 ( .A(p_input[6848]), .Z(n12167) );
  XNOR U11717 ( .A(p_input[6784]), .B(n12168), .Z(n11761) );
  AND U11718 ( .A(n257), .B(n12169), .Z(n12168) );
  XOR U11719 ( .A(p_input[6816]), .B(p_input[6784]), .Z(n12169) );
  XOR U11720 ( .A(n12170), .B(n12171), .Z(n257) );
  AND U11721 ( .A(n12172), .B(n12173), .Z(n12171) );
  XNOR U11722 ( .A(p_input[6847]), .B(n12170), .Z(n12173) );
  XOR U11723 ( .A(n12170), .B(p_input[6815]), .Z(n12172) );
  XOR U11724 ( .A(n12174), .B(n12175), .Z(n12170) );
  AND U11725 ( .A(n12176), .B(n12177), .Z(n12175) );
  XNOR U11726 ( .A(p_input[6846]), .B(n12174), .Z(n12177) );
  XNOR U11727 ( .A(n12174), .B(n11776), .Z(n12176) );
  IV U11728 ( .A(p_input[6814]), .Z(n11776) );
  XOR U11729 ( .A(n12178), .B(n12179), .Z(n12174) );
  AND U11730 ( .A(n12180), .B(n12181), .Z(n12179) );
  XNOR U11731 ( .A(p_input[6845]), .B(n12178), .Z(n12181) );
  XNOR U11732 ( .A(n12178), .B(n11785), .Z(n12180) );
  IV U11733 ( .A(p_input[6813]), .Z(n11785) );
  XOR U11734 ( .A(n12182), .B(n12183), .Z(n12178) );
  AND U11735 ( .A(n12184), .B(n12185), .Z(n12183) );
  XNOR U11736 ( .A(p_input[6844]), .B(n12182), .Z(n12185) );
  XNOR U11737 ( .A(n12182), .B(n11794), .Z(n12184) );
  IV U11738 ( .A(p_input[6812]), .Z(n11794) );
  XOR U11739 ( .A(n12186), .B(n12187), .Z(n12182) );
  AND U11740 ( .A(n12188), .B(n12189), .Z(n12187) );
  XNOR U11741 ( .A(p_input[6843]), .B(n12186), .Z(n12189) );
  XNOR U11742 ( .A(n12186), .B(n11803), .Z(n12188) );
  IV U11743 ( .A(p_input[6811]), .Z(n11803) );
  XOR U11744 ( .A(n12190), .B(n12191), .Z(n12186) );
  AND U11745 ( .A(n12192), .B(n12193), .Z(n12191) );
  XNOR U11746 ( .A(p_input[6842]), .B(n12190), .Z(n12193) );
  XNOR U11747 ( .A(n12190), .B(n11812), .Z(n12192) );
  IV U11748 ( .A(p_input[6810]), .Z(n11812) );
  XOR U11749 ( .A(n12194), .B(n12195), .Z(n12190) );
  AND U11750 ( .A(n12196), .B(n12197), .Z(n12195) );
  XNOR U11751 ( .A(p_input[6841]), .B(n12194), .Z(n12197) );
  XNOR U11752 ( .A(n12194), .B(n11821), .Z(n12196) );
  IV U11753 ( .A(p_input[6809]), .Z(n11821) );
  XOR U11754 ( .A(n12198), .B(n12199), .Z(n12194) );
  AND U11755 ( .A(n12200), .B(n12201), .Z(n12199) );
  XNOR U11756 ( .A(p_input[6840]), .B(n12198), .Z(n12201) );
  XNOR U11757 ( .A(n12198), .B(n11830), .Z(n12200) );
  IV U11758 ( .A(p_input[6808]), .Z(n11830) );
  XOR U11759 ( .A(n12202), .B(n12203), .Z(n12198) );
  AND U11760 ( .A(n12204), .B(n12205), .Z(n12203) );
  XNOR U11761 ( .A(p_input[6839]), .B(n12202), .Z(n12205) );
  XNOR U11762 ( .A(n12202), .B(n11839), .Z(n12204) );
  IV U11763 ( .A(p_input[6807]), .Z(n11839) );
  XOR U11764 ( .A(n12206), .B(n12207), .Z(n12202) );
  AND U11765 ( .A(n12208), .B(n12209), .Z(n12207) );
  XNOR U11766 ( .A(p_input[6838]), .B(n12206), .Z(n12209) );
  XNOR U11767 ( .A(n12206), .B(n11848), .Z(n12208) );
  IV U11768 ( .A(p_input[6806]), .Z(n11848) );
  XOR U11769 ( .A(n12210), .B(n12211), .Z(n12206) );
  AND U11770 ( .A(n12212), .B(n12213), .Z(n12211) );
  XNOR U11771 ( .A(p_input[6837]), .B(n12210), .Z(n12213) );
  XNOR U11772 ( .A(n12210), .B(n11857), .Z(n12212) );
  IV U11773 ( .A(p_input[6805]), .Z(n11857) );
  XOR U11774 ( .A(n12214), .B(n12215), .Z(n12210) );
  AND U11775 ( .A(n12216), .B(n12217), .Z(n12215) );
  XNOR U11776 ( .A(p_input[6836]), .B(n12214), .Z(n12217) );
  XNOR U11777 ( .A(n12214), .B(n11866), .Z(n12216) );
  IV U11778 ( .A(p_input[6804]), .Z(n11866) );
  XOR U11779 ( .A(n12218), .B(n12219), .Z(n12214) );
  AND U11780 ( .A(n12220), .B(n12221), .Z(n12219) );
  XNOR U11781 ( .A(p_input[6835]), .B(n12218), .Z(n12221) );
  XNOR U11782 ( .A(n12218), .B(n11875), .Z(n12220) );
  IV U11783 ( .A(p_input[6803]), .Z(n11875) );
  XOR U11784 ( .A(n12222), .B(n12223), .Z(n12218) );
  AND U11785 ( .A(n12224), .B(n12225), .Z(n12223) );
  XNOR U11786 ( .A(p_input[6834]), .B(n12222), .Z(n12225) );
  XNOR U11787 ( .A(n12222), .B(n11884), .Z(n12224) );
  IV U11788 ( .A(p_input[6802]), .Z(n11884) );
  XOR U11789 ( .A(n12226), .B(n12227), .Z(n12222) );
  AND U11790 ( .A(n12228), .B(n12229), .Z(n12227) );
  XNOR U11791 ( .A(p_input[6833]), .B(n12226), .Z(n12229) );
  XNOR U11792 ( .A(n12226), .B(n11893), .Z(n12228) );
  IV U11793 ( .A(p_input[6801]), .Z(n11893) );
  XOR U11794 ( .A(n12230), .B(n12231), .Z(n12226) );
  AND U11795 ( .A(n12232), .B(n12233), .Z(n12231) );
  XNOR U11796 ( .A(p_input[6832]), .B(n12230), .Z(n12233) );
  XNOR U11797 ( .A(n12230), .B(n11902), .Z(n12232) );
  IV U11798 ( .A(p_input[6800]), .Z(n11902) );
  XOR U11799 ( .A(n12234), .B(n12235), .Z(n12230) );
  AND U11800 ( .A(n12236), .B(n12237), .Z(n12235) );
  XNOR U11801 ( .A(p_input[6831]), .B(n12234), .Z(n12237) );
  XNOR U11802 ( .A(n12234), .B(n11911), .Z(n12236) );
  IV U11803 ( .A(p_input[6799]), .Z(n11911) );
  XOR U11804 ( .A(n12238), .B(n12239), .Z(n12234) );
  AND U11805 ( .A(n12240), .B(n12241), .Z(n12239) );
  XNOR U11806 ( .A(p_input[6830]), .B(n12238), .Z(n12241) );
  XNOR U11807 ( .A(n12238), .B(n11920), .Z(n12240) );
  IV U11808 ( .A(p_input[6798]), .Z(n11920) );
  XOR U11809 ( .A(n12242), .B(n12243), .Z(n12238) );
  AND U11810 ( .A(n12244), .B(n12245), .Z(n12243) );
  XNOR U11811 ( .A(p_input[6829]), .B(n12242), .Z(n12245) );
  XNOR U11812 ( .A(n12242), .B(n11929), .Z(n12244) );
  IV U11813 ( .A(p_input[6797]), .Z(n11929) );
  XOR U11814 ( .A(n12246), .B(n12247), .Z(n12242) );
  AND U11815 ( .A(n12248), .B(n12249), .Z(n12247) );
  XNOR U11816 ( .A(p_input[6828]), .B(n12246), .Z(n12249) );
  XNOR U11817 ( .A(n12246), .B(n11938), .Z(n12248) );
  IV U11818 ( .A(p_input[6796]), .Z(n11938) );
  XOR U11819 ( .A(n12250), .B(n12251), .Z(n12246) );
  AND U11820 ( .A(n12252), .B(n12253), .Z(n12251) );
  XNOR U11821 ( .A(p_input[6827]), .B(n12250), .Z(n12253) );
  XNOR U11822 ( .A(n12250), .B(n11947), .Z(n12252) );
  IV U11823 ( .A(p_input[6795]), .Z(n11947) );
  XOR U11824 ( .A(n12254), .B(n12255), .Z(n12250) );
  AND U11825 ( .A(n12256), .B(n12257), .Z(n12255) );
  XNOR U11826 ( .A(p_input[6826]), .B(n12254), .Z(n12257) );
  XNOR U11827 ( .A(n12254), .B(n11956), .Z(n12256) );
  IV U11828 ( .A(p_input[6794]), .Z(n11956) );
  XOR U11829 ( .A(n12258), .B(n12259), .Z(n12254) );
  AND U11830 ( .A(n12260), .B(n12261), .Z(n12259) );
  XNOR U11831 ( .A(p_input[6825]), .B(n12258), .Z(n12261) );
  XNOR U11832 ( .A(n12258), .B(n11965), .Z(n12260) );
  IV U11833 ( .A(p_input[6793]), .Z(n11965) );
  XOR U11834 ( .A(n12262), .B(n12263), .Z(n12258) );
  AND U11835 ( .A(n12264), .B(n12265), .Z(n12263) );
  XNOR U11836 ( .A(p_input[6824]), .B(n12262), .Z(n12265) );
  XNOR U11837 ( .A(n12262), .B(n11974), .Z(n12264) );
  IV U11838 ( .A(p_input[6792]), .Z(n11974) );
  XOR U11839 ( .A(n12266), .B(n12267), .Z(n12262) );
  AND U11840 ( .A(n12268), .B(n12269), .Z(n12267) );
  XNOR U11841 ( .A(p_input[6823]), .B(n12266), .Z(n12269) );
  XNOR U11842 ( .A(n12266), .B(n11983), .Z(n12268) );
  IV U11843 ( .A(p_input[6791]), .Z(n11983) );
  XOR U11844 ( .A(n12270), .B(n12271), .Z(n12266) );
  AND U11845 ( .A(n12272), .B(n12273), .Z(n12271) );
  XNOR U11846 ( .A(p_input[6822]), .B(n12270), .Z(n12273) );
  XNOR U11847 ( .A(n12270), .B(n11992), .Z(n12272) );
  IV U11848 ( .A(p_input[6790]), .Z(n11992) );
  XOR U11849 ( .A(n12274), .B(n12275), .Z(n12270) );
  AND U11850 ( .A(n12276), .B(n12277), .Z(n12275) );
  XNOR U11851 ( .A(p_input[6821]), .B(n12274), .Z(n12277) );
  XNOR U11852 ( .A(n12274), .B(n12001), .Z(n12276) );
  IV U11853 ( .A(p_input[6789]), .Z(n12001) );
  XOR U11854 ( .A(n12278), .B(n12279), .Z(n12274) );
  AND U11855 ( .A(n12280), .B(n12281), .Z(n12279) );
  XNOR U11856 ( .A(p_input[6820]), .B(n12278), .Z(n12281) );
  XNOR U11857 ( .A(n12278), .B(n12010), .Z(n12280) );
  IV U11858 ( .A(p_input[6788]), .Z(n12010) );
  XOR U11859 ( .A(n12282), .B(n12283), .Z(n12278) );
  AND U11860 ( .A(n12284), .B(n12285), .Z(n12283) );
  XNOR U11861 ( .A(p_input[6819]), .B(n12282), .Z(n12285) );
  XNOR U11862 ( .A(n12282), .B(n12019), .Z(n12284) );
  IV U11863 ( .A(p_input[6787]), .Z(n12019) );
  XOR U11864 ( .A(n12286), .B(n12287), .Z(n12282) );
  AND U11865 ( .A(n12288), .B(n12289), .Z(n12287) );
  XNOR U11866 ( .A(p_input[6818]), .B(n12286), .Z(n12289) );
  XNOR U11867 ( .A(n12286), .B(n12028), .Z(n12288) );
  IV U11868 ( .A(p_input[6786]), .Z(n12028) );
  XNOR U11869 ( .A(n12290), .B(n12291), .Z(n12286) );
  AND U11870 ( .A(n12292), .B(n12293), .Z(n12291) );
  XOR U11871 ( .A(p_input[6817]), .B(n12290), .Z(n12293) );
  XNOR U11872 ( .A(p_input[6785]), .B(n12290), .Z(n12292) );
  AND U11873 ( .A(p_input[6816]), .B(n12294), .Z(n12290) );
  IV U11874 ( .A(p_input[6784]), .Z(n12294) );
  XOR U11875 ( .A(n12295), .B(n12296), .Z(n11384) );
  AND U11876 ( .A(n468), .B(n12297), .Z(n12296) );
  XNOR U11877 ( .A(n12298), .B(n12295), .Z(n12297) );
  XOR U11878 ( .A(n12299), .B(n12300), .Z(n468) );
  AND U11879 ( .A(n12301), .B(n12302), .Z(n12300) );
  XNOR U11880 ( .A(n11399), .B(n12299), .Z(n12302) );
  AND U11881 ( .A(p_input[6783]), .B(p_input[6751]), .Z(n11399) );
  XNOR U11882 ( .A(n12299), .B(n11396), .Z(n12301) );
  IV U11883 ( .A(n12303), .Z(n11396) );
  AND U11884 ( .A(p_input[6687]), .B(p_input[6719]), .Z(n12303) );
  XOR U11885 ( .A(n12304), .B(n12305), .Z(n12299) );
  AND U11886 ( .A(n12306), .B(n12307), .Z(n12305) );
  XOR U11887 ( .A(n12304), .B(n11411), .Z(n12307) );
  XNOR U11888 ( .A(p_input[6750]), .B(n12308), .Z(n11411) );
  AND U11889 ( .A(n263), .B(n12309), .Z(n12308) );
  XOR U11890 ( .A(p_input[6782]), .B(p_input[6750]), .Z(n12309) );
  XNOR U11891 ( .A(n11408), .B(n12304), .Z(n12306) );
  XOR U11892 ( .A(n12310), .B(n12311), .Z(n11408) );
  AND U11893 ( .A(n260), .B(n12312), .Z(n12311) );
  XOR U11894 ( .A(p_input[6718]), .B(p_input[6686]), .Z(n12312) );
  XOR U11895 ( .A(n12313), .B(n12314), .Z(n12304) );
  AND U11896 ( .A(n12315), .B(n12316), .Z(n12314) );
  XOR U11897 ( .A(n12313), .B(n11423), .Z(n12316) );
  XNOR U11898 ( .A(p_input[6749]), .B(n12317), .Z(n11423) );
  AND U11899 ( .A(n263), .B(n12318), .Z(n12317) );
  XOR U11900 ( .A(p_input[6781]), .B(p_input[6749]), .Z(n12318) );
  XNOR U11901 ( .A(n11420), .B(n12313), .Z(n12315) );
  XOR U11902 ( .A(n12319), .B(n12320), .Z(n11420) );
  AND U11903 ( .A(n260), .B(n12321), .Z(n12320) );
  XOR U11904 ( .A(p_input[6717]), .B(p_input[6685]), .Z(n12321) );
  XOR U11905 ( .A(n12322), .B(n12323), .Z(n12313) );
  AND U11906 ( .A(n12324), .B(n12325), .Z(n12323) );
  XOR U11907 ( .A(n12322), .B(n11435), .Z(n12325) );
  XNOR U11908 ( .A(p_input[6748]), .B(n12326), .Z(n11435) );
  AND U11909 ( .A(n263), .B(n12327), .Z(n12326) );
  XOR U11910 ( .A(p_input[6780]), .B(p_input[6748]), .Z(n12327) );
  XNOR U11911 ( .A(n11432), .B(n12322), .Z(n12324) );
  XOR U11912 ( .A(n12328), .B(n12329), .Z(n11432) );
  AND U11913 ( .A(n260), .B(n12330), .Z(n12329) );
  XOR U11914 ( .A(p_input[6716]), .B(p_input[6684]), .Z(n12330) );
  XOR U11915 ( .A(n12331), .B(n12332), .Z(n12322) );
  AND U11916 ( .A(n12333), .B(n12334), .Z(n12332) );
  XOR U11917 ( .A(n12331), .B(n11447), .Z(n12334) );
  XNOR U11918 ( .A(p_input[6747]), .B(n12335), .Z(n11447) );
  AND U11919 ( .A(n263), .B(n12336), .Z(n12335) );
  XOR U11920 ( .A(p_input[6779]), .B(p_input[6747]), .Z(n12336) );
  XNOR U11921 ( .A(n11444), .B(n12331), .Z(n12333) );
  XOR U11922 ( .A(n12337), .B(n12338), .Z(n11444) );
  AND U11923 ( .A(n260), .B(n12339), .Z(n12338) );
  XOR U11924 ( .A(p_input[6715]), .B(p_input[6683]), .Z(n12339) );
  XOR U11925 ( .A(n12340), .B(n12341), .Z(n12331) );
  AND U11926 ( .A(n12342), .B(n12343), .Z(n12341) );
  XOR U11927 ( .A(n12340), .B(n11459), .Z(n12343) );
  XNOR U11928 ( .A(p_input[6746]), .B(n12344), .Z(n11459) );
  AND U11929 ( .A(n263), .B(n12345), .Z(n12344) );
  XOR U11930 ( .A(p_input[6778]), .B(p_input[6746]), .Z(n12345) );
  XNOR U11931 ( .A(n11456), .B(n12340), .Z(n12342) );
  XOR U11932 ( .A(n12346), .B(n12347), .Z(n11456) );
  AND U11933 ( .A(n260), .B(n12348), .Z(n12347) );
  XOR U11934 ( .A(p_input[6714]), .B(p_input[6682]), .Z(n12348) );
  XOR U11935 ( .A(n12349), .B(n12350), .Z(n12340) );
  AND U11936 ( .A(n12351), .B(n12352), .Z(n12350) );
  XOR U11937 ( .A(n12349), .B(n11471), .Z(n12352) );
  XNOR U11938 ( .A(p_input[6745]), .B(n12353), .Z(n11471) );
  AND U11939 ( .A(n263), .B(n12354), .Z(n12353) );
  XOR U11940 ( .A(p_input[6777]), .B(p_input[6745]), .Z(n12354) );
  XNOR U11941 ( .A(n11468), .B(n12349), .Z(n12351) );
  XOR U11942 ( .A(n12355), .B(n12356), .Z(n11468) );
  AND U11943 ( .A(n260), .B(n12357), .Z(n12356) );
  XOR U11944 ( .A(p_input[6713]), .B(p_input[6681]), .Z(n12357) );
  XOR U11945 ( .A(n12358), .B(n12359), .Z(n12349) );
  AND U11946 ( .A(n12360), .B(n12361), .Z(n12359) );
  XOR U11947 ( .A(n12358), .B(n11483), .Z(n12361) );
  XNOR U11948 ( .A(p_input[6744]), .B(n12362), .Z(n11483) );
  AND U11949 ( .A(n263), .B(n12363), .Z(n12362) );
  XOR U11950 ( .A(p_input[6776]), .B(p_input[6744]), .Z(n12363) );
  XNOR U11951 ( .A(n11480), .B(n12358), .Z(n12360) );
  XOR U11952 ( .A(n12364), .B(n12365), .Z(n11480) );
  AND U11953 ( .A(n260), .B(n12366), .Z(n12365) );
  XOR U11954 ( .A(p_input[6712]), .B(p_input[6680]), .Z(n12366) );
  XOR U11955 ( .A(n12367), .B(n12368), .Z(n12358) );
  AND U11956 ( .A(n12369), .B(n12370), .Z(n12368) );
  XOR U11957 ( .A(n12367), .B(n11495), .Z(n12370) );
  XNOR U11958 ( .A(p_input[6743]), .B(n12371), .Z(n11495) );
  AND U11959 ( .A(n263), .B(n12372), .Z(n12371) );
  XOR U11960 ( .A(p_input[6775]), .B(p_input[6743]), .Z(n12372) );
  XNOR U11961 ( .A(n11492), .B(n12367), .Z(n12369) );
  XOR U11962 ( .A(n12373), .B(n12374), .Z(n11492) );
  AND U11963 ( .A(n260), .B(n12375), .Z(n12374) );
  XOR U11964 ( .A(p_input[6711]), .B(p_input[6679]), .Z(n12375) );
  XOR U11965 ( .A(n12376), .B(n12377), .Z(n12367) );
  AND U11966 ( .A(n12378), .B(n12379), .Z(n12377) );
  XOR U11967 ( .A(n12376), .B(n11507), .Z(n12379) );
  XNOR U11968 ( .A(p_input[6742]), .B(n12380), .Z(n11507) );
  AND U11969 ( .A(n263), .B(n12381), .Z(n12380) );
  XOR U11970 ( .A(p_input[6774]), .B(p_input[6742]), .Z(n12381) );
  XNOR U11971 ( .A(n11504), .B(n12376), .Z(n12378) );
  XOR U11972 ( .A(n12382), .B(n12383), .Z(n11504) );
  AND U11973 ( .A(n260), .B(n12384), .Z(n12383) );
  XOR U11974 ( .A(p_input[6710]), .B(p_input[6678]), .Z(n12384) );
  XOR U11975 ( .A(n12385), .B(n12386), .Z(n12376) );
  AND U11976 ( .A(n12387), .B(n12388), .Z(n12386) );
  XOR U11977 ( .A(n12385), .B(n11519), .Z(n12388) );
  XNOR U11978 ( .A(p_input[6741]), .B(n12389), .Z(n11519) );
  AND U11979 ( .A(n263), .B(n12390), .Z(n12389) );
  XOR U11980 ( .A(p_input[6773]), .B(p_input[6741]), .Z(n12390) );
  XNOR U11981 ( .A(n11516), .B(n12385), .Z(n12387) );
  XOR U11982 ( .A(n12391), .B(n12392), .Z(n11516) );
  AND U11983 ( .A(n260), .B(n12393), .Z(n12392) );
  XOR U11984 ( .A(p_input[6709]), .B(p_input[6677]), .Z(n12393) );
  XOR U11985 ( .A(n12394), .B(n12395), .Z(n12385) );
  AND U11986 ( .A(n12396), .B(n12397), .Z(n12395) );
  XOR U11987 ( .A(n12394), .B(n11531), .Z(n12397) );
  XNOR U11988 ( .A(p_input[6740]), .B(n12398), .Z(n11531) );
  AND U11989 ( .A(n263), .B(n12399), .Z(n12398) );
  XOR U11990 ( .A(p_input[6772]), .B(p_input[6740]), .Z(n12399) );
  XNOR U11991 ( .A(n11528), .B(n12394), .Z(n12396) );
  XOR U11992 ( .A(n12400), .B(n12401), .Z(n11528) );
  AND U11993 ( .A(n260), .B(n12402), .Z(n12401) );
  XOR U11994 ( .A(p_input[6708]), .B(p_input[6676]), .Z(n12402) );
  XOR U11995 ( .A(n12403), .B(n12404), .Z(n12394) );
  AND U11996 ( .A(n12405), .B(n12406), .Z(n12404) );
  XOR U11997 ( .A(n12403), .B(n11543), .Z(n12406) );
  XNOR U11998 ( .A(p_input[6739]), .B(n12407), .Z(n11543) );
  AND U11999 ( .A(n263), .B(n12408), .Z(n12407) );
  XOR U12000 ( .A(p_input[6771]), .B(p_input[6739]), .Z(n12408) );
  XNOR U12001 ( .A(n11540), .B(n12403), .Z(n12405) );
  XOR U12002 ( .A(n12409), .B(n12410), .Z(n11540) );
  AND U12003 ( .A(n260), .B(n12411), .Z(n12410) );
  XOR U12004 ( .A(p_input[6707]), .B(p_input[6675]), .Z(n12411) );
  XOR U12005 ( .A(n12412), .B(n12413), .Z(n12403) );
  AND U12006 ( .A(n12414), .B(n12415), .Z(n12413) );
  XOR U12007 ( .A(n12412), .B(n11555), .Z(n12415) );
  XNOR U12008 ( .A(p_input[6738]), .B(n12416), .Z(n11555) );
  AND U12009 ( .A(n263), .B(n12417), .Z(n12416) );
  XOR U12010 ( .A(p_input[6770]), .B(p_input[6738]), .Z(n12417) );
  XNOR U12011 ( .A(n11552), .B(n12412), .Z(n12414) );
  XOR U12012 ( .A(n12418), .B(n12419), .Z(n11552) );
  AND U12013 ( .A(n260), .B(n12420), .Z(n12419) );
  XOR U12014 ( .A(p_input[6706]), .B(p_input[6674]), .Z(n12420) );
  XOR U12015 ( .A(n12421), .B(n12422), .Z(n12412) );
  AND U12016 ( .A(n12423), .B(n12424), .Z(n12422) );
  XOR U12017 ( .A(n12421), .B(n11567), .Z(n12424) );
  XNOR U12018 ( .A(p_input[6737]), .B(n12425), .Z(n11567) );
  AND U12019 ( .A(n263), .B(n12426), .Z(n12425) );
  XOR U12020 ( .A(p_input[6769]), .B(p_input[6737]), .Z(n12426) );
  XNOR U12021 ( .A(n11564), .B(n12421), .Z(n12423) );
  XOR U12022 ( .A(n12427), .B(n12428), .Z(n11564) );
  AND U12023 ( .A(n260), .B(n12429), .Z(n12428) );
  XOR U12024 ( .A(p_input[6705]), .B(p_input[6673]), .Z(n12429) );
  XOR U12025 ( .A(n12430), .B(n12431), .Z(n12421) );
  AND U12026 ( .A(n12432), .B(n12433), .Z(n12431) );
  XOR U12027 ( .A(n12430), .B(n11579), .Z(n12433) );
  XNOR U12028 ( .A(p_input[6736]), .B(n12434), .Z(n11579) );
  AND U12029 ( .A(n263), .B(n12435), .Z(n12434) );
  XOR U12030 ( .A(p_input[6768]), .B(p_input[6736]), .Z(n12435) );
  XNOR U12031 ( .A(n11576), .B(n12430), .Z(n12432) );
  XOR U12032 ( .A(n12436), .B(n12437), .Z(n11576) );
  AND U12033 ( .A(n260), .B(n12438), .Z(n12437) );
  XOR U12034 ( .A(p_input[6704]), .B(p_input[6672]), .Z(n12438) );
  XOR U12035 ( .A(n12439), .B(n12440), .Z(n12430) );
  AND U12036 ( .A(n12441), .B(n12442), .Z(n12440) );
  XOR U12037 ( .A(n12439), .B(n11591), .Z(n12442) );
  XNOR U12038 ( .A(p_input[6735]), .B(n12443), .Z(n11591) );
  AND U12039 ( .A(n263), .B(n12444), .Z(n12443) );
  XOR U12040 ( .A(p_input[6767]), .B(p_input[6735]), .Z(n12444) );
  XNOR U12041 ( .A(n11588), .B(n12439), .Z(n12441) );
  XOR U12042 ( .A(n12445), .B(n12446), .Z(n11588) );
  AND U12043 ( .A(n260), .B(n12447), .Z(n12446) );
  XOR U12044 ( .A(p_input[6703]), .B(p_input[6671]), .Z(n12447) );
  XOR U12045 ( .A(n12448), .B(n12449), .Z(n12439) );
  AND U12046 ( .A(n12450), .B(n12451), .Z(n12449) );
  XOR U12047 ( .A(n12448), .B(n11603), .Z(n12451) );
  XNOR U12048 ( .A(p_input[6734]), .B(n12452), .Z(n11603) );
  AND U12049 ( .A(n263), .B(n12453), .Z(n12452) );
  XOR U12050 ( .A(p_input[6766]), .B(p_input[6734]), .Z(n12453) );
  XNOR U12051 ( .A(n11600), .B(n12448), .Z(n12450) );
  XOR U12052 ( .A(n12454), .B(n12455), .Z(n11600) );
  AND U12053 ( .A(n260), .B(n12456), .Z(n12455) );
  XOR U12054 ( .A(p_input[6702]), .B(p_input[6670]), .Z(n12456) );
  XOR U12055 ( .A(n12457), .B(n12458), .Z(n12448) );
  AND U12056 ( .A(n12459), .B(n12460), .Z(n12458) );
  XOR U12057 ( .A(n12457), .B(n11615), .Z(n12460) );
  XNOR U12058 ( .A(p_input[6733]), .B(n12461), .Z(n11615) );
  AND U12059 ( .A(n263), .B(n12462), .Z(n12461) );
  XOR U12060 ( .A(p_input[6765]), .B(p_input[6733]), .Z(n12462) );
  XNOR U12061 ( .A(n11612), .B(n12457), .Z(n12459) );
  XOR U12062 ( .A(n12463), .B(n12464), .Z(n11612) );
  AND U12063 ( .A(n260), .B(n12465), .Z(n12464) );
  XOR U12064 ( .A(p_input[6701]), .B(p_input[6669]), .Z(n12465) );
  XOR U12065 ( .A(n12466), .B(n12467), .Z(n12457) );
  AND U12066 ( .A(n12468), .B(n12469), .Z(n12467) );
  XOR U12067 ( .A(n12466), .B(n11627), .Z(n12469) );
  XNOR U12068 ( .A(p_input[6732]), .B(n12470), .Z(n11627) );
  AND U12069 ( .A(n263), .B(n12471), .Z(n12470) );
  XOR U12070 ( .A(p_input[6764]), .B(p_input[6732]), .Z(n12471) );
  XNOR U12071 ( .A(n11624), .B(n12466), .Z(n12468) );
  XOR U12072 ( .A(n12472), .B(n12473), .Z(n11624) );
  AND U12073 ( .A(n260), .B(n12474), .Z(n12473) );
  XOR U12074 ( .A(p_input[6700]), .B(p_input[6668]), .Z(n12474) );
  XOR U12075 ( .A(n12475), .B(n12476), .Z(n12466) );
  AND U12076 ( .A(n12477), .B(n12478), .Z(n12476) );
  XOR U12077 ( .A(n12475), .B(n11639), .Z(n12478) );
  XNOR U12078 ( .A(p_input[6731]), .B(n12479), .Z(n11639) );
  AND U12079 ( .A(n263), .B(n12480), .Z(n12479) );
  XOR U12080 ( .A(p_input[6763]), .B(p_input[6731]), .Z(n12480) );
  XNOR U12081 ( .A(n11636), .B(n12475), .Z(n12477) );
  XOR U12082 ( .A(n12481), .B(n12482), .Z(n11636) );
  AND U12083 ( .A(n260), .B(n12483), .Z(n12482) );
  XOR U12084 ( .A(p_input[6699]), .B(p_input[6667]), .Z(n12483) );
  XOR U12085 ( .A(n12484), .B(n12485), .Z(n12475) );
  AND U12086 ( .A(n12486), .B(n12487), .Z(n12485) );
  XOR U12087 ( .A(n12484), .B(n11651), .Z(n12487) );
  XNOR U12088 ( .A(p_input[6730]), .B(n12488), .Z(n11651) );
  AND U12089 ( .A(n263), .B(n12489), .Z(n12488) );
  XOR U12090 ( .A(p_input[6762]), .B(p_input[6730]), .Z(n12489) );
  XNOR U12091 ( .A(n11648), .B(n12484), .Z(n12486) );
  XOR U12092 ( .A(n12490), .B(n12491), .Z(n11648) );
  AND U12093 ( .A(n260), .B(n12492), .Z(n12491) );
  XOR U12094 ( .A(p_input[6698]), .B(p_input[6666]), .Z(n12492) );
  XOR U12095 ( .A(n12493), .B(n12494), .Z(n12484) );
  AND U12096 ( .A(n12495), .B(n12496), .Z(n12494) );
  XOR U12097 ( .A(n12493), .B(n11663), .Z(n12496) );
  XNOR U12098 ( .A(p_input[6729]), .B(n12497), .Z(n11663) );
  AND U12099 ( .A(n263), .B(n12498), .Z(n12497) );
  XOR U12100 ( .A(p_input[6761]), .B(p_input[6729]), .Z(n12498) );
  XNOR U12101 ( .A(n11660), .B(n12493), .Z(n12495) );
  XOR U12102 ( .A(n12499), .B(n12500), .Z(n11660) );
  AND U12103 ( .A(n260), .B(n12501), .Z(n12500) );
  XOR U12104 ( .A(p_input[6697]), .B(p_input[6665]), .Z(n12501) );
  XOR U12105 ( .A(n12502), .B(n12503), .Z(n12493) );
  AND U12106 ( .A(n12504), .B(n12505), .Z(n12503) );
  XOR U12107 ( .A(n12502), .B(n11675), .Z(n12505) );
  XNOR U12108 ( .A(p_input[6728]), .B(n12506), .Z(n11675) );
  AND U12109 ( .A(n263), .B(n12507), .Z(n12506) );
  XOR U12110 ( .A(p_input[6760]), .B(p_input[6728]), .Z(n12507) );
  XNOR U12111 ( .A(n11672), .B(n12502), .Z(n12504) );
  XOR U12112 ( .A(n12508), .B(n12509), .Z(n11672) );
  AND U12113 ( .A(n260), .B(n12510), .Z(n12509) );
  XOR U12114 ( .A(p_input[6696]), .B(p_input[6664]), .Z(n12510) );
  XOR U12115 ( .A(n12511), .B(n12512), .Z(n12502) );
  AND U12116 ( .A(n12513), .B(n12514), .Z(n12512) );
  XOR U12117 ( .A(n12511), .B(n11687), .Z(n12514) );
  XNOR U12118 ( .A(p_input[6727]), .B(n12515), .Z(n11687) );
  AND U12119 ( .A(n263), .B(n12516), .Z(n12515) );
  XOR U12120 ( .A(p_input[6759]), .B(p_input[6727]), .Z(n12516) );
  XNOR U12121 ( .A(n11684), .B(n12511), .Z(n12513) );
  XOR U12122 ( .A(n12517), .B(n12518), .Z(n11684) );
  AND U12123 ( .A(n260), .B(n12519), .Z(n12518) );
  XOR U12124 ( .A(p_input[6695]), .B(p_input[6663]), .Z(n12519) );
  XOR U12125 ( .A(n12520), .B(n12521), .Z(n12511) );
  AND U12126 ( .A(n12522), .B(n12523), .Z(n12521) );
  XOR U12127 ( .A(n12520), .B(n11699), .Z(n12523) );
  XNOR U12128 ( .A(p_input[6726]), .B(n12524), .Z(n11699) );
  AND U12129 ( .A(n263), .B(n12525), .Z(n12524) );
  XOR U12130 ( .A(p_input[6758]), .B(p_input[6726]), .Z(n12525) );
  XNOR U12131 ( .A(n11696), .B(n12520), .Z(n12522) );
  XOR U12132 ( .A(n12526), .B(n12527), .Z(n11696) );
  AND U12133 ( .A(n260), .B(n12528), .Z(n12527) );
  XOR U12134 ( .A(p_input[6694]), .B(p_input[6662]), .Z(n12528) );
  XOR U12135 ( .A(n12529), .B(n12530), .Z(n12520) );
  AND U12136 ( .A(n12531), .B(n12532), .Z(n12530) );
  XOR U12137 ( .A(n12529), .B(n11711), .Z(n12532) );
  XNOR U12138 ( .A(p_input[6725]), .B(n12533), .Z(n11711) );
  AND U12139 ( .A(n263), .B(n12534), .Z(n12533) );
  XOR U12140 ( .A(p_input[6757]), .B(p_input[6725]), .Z(n12534) );
  XNOR U12141 ( .A(n11708), .B(n12529), .Z(n12531) );
  XOR U12142 ( .A(n12535), .B(n12536), .Z(n11708) );
  AND U12143 ( .A(n260), .B(n12537), .Z(n12536) );
  XOR U12144 ( .A(p_input[6693]), .B(p_input[6661]), .Z(n12537) );
  XOR U12145 ( .A(n12538), .B(n12539), .Z(n12529) );
  AND U12146 ( .A(n12540), .B(n12541), .Z(n12539) );
  XOR U12147 ( .A(n12538), .B(n11723), .Z(n12541) );
  XNOR U12148 ( .A(p_input[6724]), .B(n12542), .Z(n11723) );
  AND U12149 ( .A(n263), .B(n12543), .Z(n12542) );
  XOR U12150 ( .A(p_input[6756]), .B(p_input[6724]), .Z(n12543) );
  XNOR U12151 ( .A(n11720), .B(n12538), .Z(n12540) );
  XOR U12152 ( .A(n12544), .B(n12545), .Z(n11720) );
  AND U12153 ( .A(n260), .B(n12546), .Z(n12545) );
  XOR U12154 ( .A(p_input[6692]), .B(p_input[6660]), .Z(n12546) );
  XOR U12155 ( .A(n12547), .B(n12548), .Z(n12538) );
  AND U12156 ( .A(n12549), .B(n12550), .Z(n12548) );
  XOR U12157 ( .A(n12547), .B(n11735), .Z(n12550) );
  XNOR U12158 ( .A(p_input[6723]), .B(n12551), .Z(n11735) );
  AND U12159 ( .A(n263), .B(n12552), .Z(n12551) );
  XOR U12160 ( .A(p_input[6755]), .B(p_input[6723]), .Z(n12552) );
  XNOR U12161 ( .A(n11732), .B(n12547), .Z(n12549) );
  XOR U12162 ( .A(n12553), .B(n12554), .Z(n11732) );
  AND U12163 ( .A(n260), .B(n12555), .Z(n12554) );
  XOR U12164 ( .A(p_input[6691]), .B(p_input[6659]), .Z(n12555) );
  XOR U12165 ( .A(n12556), .B(n12557), .Z(n12547) );
  AND U12166 ( .A(n12558), .B(n12559), .Z(n12557) );
  XOR U12167 ( .A(n12556), .B(n11747), .Z(n12559) );
  XNOR U12168 ( .A(p_input[6722]), .B(n12560), .Z(n11747) );
  AND U12169 ( .A(n263), .B(n12561), .Z(n12560) );
  XOR U12170 ( .A(p_input[6754]), .B(p_input[6722]), .Z(n12561) );
  XNOR U12171 ( .A(n11744), .B(n12556), .Z(n12558) );
  XOR U12172 ( .A(n12562), .B(n12563), .Z(n11744) );
  AND U12173 ( .A(n260), .B(n12564), .Z(n12563) );
  XOR U12174 ( .A(p_input[6690]), .B(p_input[6658]), .Z(n12564) );
  XOR U12175 ( .A(n12565), .B(n12566), .Z(n12556) );
  AND U12176 ( .A(n12567), .B(n12568), .Z(n12566) );
  XNOR U12177 ( .A(n12569), .B(n11760), .Z(n12568) );
  XNOR U12178 ( .A(p_input[6721]), .B(n12570), .Z(n11760) );
  AND U12179 ( .A(n263), .B(n12571), .Z(n12570) );
  XNOR U12180 ( .A(p_input[6753]), .B(n12572), .Z(n12571) );
  IV U12181 ( .A(p_input[6721]), .Z(n12572) );
  XNOR U12182 ( .A(n11757), .B(n12565), .Z(n12567) );
  XNOR U12183 ( .A(p_input[6657]), .B(n12573), .Z(n11757) );
  AND U12184 ( .A(n260), .B(n12574), .Z(n12573) );
  XOR U12185 ( .A(p_input[6689]), .B(p_input[6657]), .Z(n12574) );
  IV U12186 ( .A(n12569), .Z(n12565) );
  AND U12187 ( .A(n12295), .B(n12298), .Z(n12569) );
  XOR U12188 ( .A(p_input[6720]), .B(n12575), .Z(n12298) );
  AND U12189 ( .A(n263), .B(n12576), .Z(n12575) );
  XOR U12190 ( .A(p_input[6752]), .B(p_input[6720]), .Z(n12576) );
  XOR U12191 ( .A(n12577), .B(n12578), .Z(n263) );
  AND U12192 ( .A(n12579), .B(n12580), .Z(n12578) );
  XNOR U12193 ( .A(p_input[6783]), .B(n12577), .Z(n12580) );
  XOR U12194 ( .A(n12577), .B(p_input[6751]), .Z(n12579) );
  XOR U12195 ( .A(n12581), .B(n12582), .Z(n12577) );
  AND U12196 ( .A(n12583), .B(n12584), .Z(n12582) );
  XNOR U12197 ( .A(p_input[6782]), .B(n12581), .Z(n12584) );
  XOR U12198 ( .A(n12581), .B(p_input[6750]), .Z(n12583) );
  XOR U12199 ( .A(n12585), .B(n12586), .Z(n12581) );
  AND U12200 ( .A(n12587), .B(n12588), .Z(n12586) );
  XNOR U12201 ( .A(p_input[6781]), .B(n12585), .Z(n12588) );
  XOR U12202 ( .A(n12585), .B(p_input[6749]), .Z(n12587) );
  XOR U12203 ( .A(n12589), .B(n12590), .Z(n12585) );
  AND U12204 ( .A(n12591), .B(n12592), .Z(n12590) );
  XNOR U12205 ( .A(p_input[6780]), .B(n12589), .Z(n12592) );
  XOR U12206 ( .A(n12589), .B(p_input[6748]), .Z(n12591) );
  XOR U12207 ( .A(n12593), .B(n12594), .Z(n12589) );
  AND U12208 ( .A(n12595), .B(n12596), .Z(n12594) );
  XNOR U12209 ( .A(p_input[6779]), .B(n12593), .Z(n12596) );
  XOR U12210 ( .A(n12593), .B(p_input[6747]), .Z(n12595) );
  XOR U12211 ( .A(n12597), .B(n12598), .Z(n12593) );
  AND U12212 ( .A(n12599), .B(n12600), .Z(n12598) );
  XNOR U12213 ( .A(p_input[6778]), .B(n12597), .Z(n12600) );
  XOR U12214 ( .A(n12597), .B(p_input[6746]), .Z(n12599) );
  XOR U12215 ( .A(n12601), .B(n12602), .Z(n12597) );
  AND U12216 ( .A(n12603), .B(n12604), .Z(n12602) );
  XNOR U12217 ( .A(p_input[6777]), .B(n12601), .Z(n12604) );
  XOR U12218 ( .A(n12601), .B(p_input[6745]), .Z(n12603) );
  XOR U12219 ( .A(n12605), .B(n12606), .Z(n12601) );
  AND U12220 ( .A(n12607), .B(n12608), .Z(n12606) );
  XNOR U12221 ( .A(p_input[6776]), .B(n12605), .Z(n12608) );
  XOR U12222 ( .A(n12605), .B(p_input[6744]), .Z(n12607) );
  XOR U12223 ( .A(n12609), .B(n12610), .Z(n12605) );
  AND U12224 ( .A(n12611), .B(n12612), .Z(n12610) );
  XNOR U12225 ( .A(p_input[6775]), .B(n12609), .Z(n12612) );
  XOR U12226 ( .A(n12609), .B(p_input[6743]), .Z(n12611) );
  XOR U12227 ( .A(n12613), .B(n12614), .Z(n12609) );
  AND U12228 ( .A(n12615), .B(n12616), .Z(n12614) );
  XNOR U12229 ( .A(p_input[6774]), .B(n12613), .Z(n12616) );
  XOR U12230 ( .A(n12613), .B(p_input[6742]), .Z(n12615) );
  XOR U12231 ( .A(n12617), .B(n12618), .Z(n12613) );
  AND U12232 ( .A(n12619), .B(n12620), .Z(n12618) );
  XNOR U12233 ( .A(p_input[6773]), .B(n12617), .Z(n12620) );
  XOR U12234 ( .A(n12617), .B(p_input[6741]), .Z(n12619) );
  XOR U12235 ( .A(n12621), .B(n12622), .Z(n12617) );
  AND U12236 ( .A(n12623), .B(n12624), .Z(n12622) );
  XNOR U12237 ( .A(p_input[6772]), .B(n12621), .Z(n12624) );
  XOR U12238 ( .A(n12621), .B(p_input[6740]), .Z(n12623) );
  XOR U12239 ( .A(n12625), .B(n12626), .Z(n12621) );
  AND U12240 ( .A(n12627), .B(n12628), .Z(n12626) );
  XNOR U12241 ( .A(p_input[6771]), .B(n12625), .Z(n12628) );
  XOR U12242 ( .A(n12625), .B(p_input[6739]), .Z(n12627) );
  XOR U12243 ( .A(n12629), .B(n12630), .Z(n12625) );
  AND U12244 ( .A(n12631), .B(n12632), .Z(n12630) );
  XNOR U12245 ( .A(p_input[6770]), .B(n12629), .Z(n12632) );
  XOR U12246 ( .A(n12629), .B(p_input[6738]), .Z(n12631) );
  XOR U12247 ( .A(n12633), .B(n12634), .Z(n12629) );
  AND U12248 ( .A(n12635), .B(n12636), .Z(n12634) );
  XNOR U12249 ( .A(p_input[6769]), .B(n12633), .Z(n12636) );
  XOR U12250 ( .A(n12633), .B(p_input[6737]), .Z(n12635) );
  XOR U12251 ( .A(n12637), .B(n12638), .Z(n12633) );
  AND U12252 ( .A(n12639), .B(n12640), .Z(n12638) );
  XNOR U12253 ( .A(p_input[6768]), .B(n12637), .Z(n12640) );
  XOR U12254 ( .A(n12637), .B(p_input[6736]), .Z(n12639) );
  XOR U12255 ( .A(n12641), .B(n12642), .Z(n12637) );
  AND U12256 ( .A(n12643), .B(n12644), .Z(n12642) );
  XNOR U12257 ( .A(p_input[6767]), .B(n12641), .Z(n12644) );
  XOR U12258 ( .A(n12641), .B(p_input[6735]), .Z(n12643) );
  XOR U12259 ( .A(n12645), .B(n12646), .Z(n12641) );
  AND U12260 ( .A(n12647), .B(n12648), .Z(n12646) );
  XNOR U12261 ( .A(p_input[6766]), .B(n12645), .Z(n12648) );
  XOR U12262 ( .A(n12645), .B(p_input[6734]), .Z(n12647) );
  XOR U12263 ( .A(n12649), .B(n12650), .Z(n12645) );
  AND U12264 ( .A(n12651), .B(n12652), .Z(n12650) );
  XNOR U12265 ( .A(p_input[6765]), .B(n12649), .Z(n12652) );
  XOR U12266 ( .A(n12649), .B(p_input[6733]), .Z(n12651) );
  XOR U12267 ( .A(n12653), .B(n12654), .Z(n12649) );
  AND U12268 ( .A(n12655), .B(n12656), .Z(n12654) );
  XNOR U12269 ( .A(p_input[6764]), .B(n12653), .Z(n12656) );
  XOR U12270 ( .A(n12653), .B(p_input[6732]), .Z(n12655) );
  XOR U12271 ( .A(n12657), .B(n12658), .Z(n12653) );
  AND U12272 ( .A(n12659), .B(n12660), .Z(n12658) );
  XNOR U12273 ( .A(p_input[6763]), .B(n12657), .Z(n12660) );
  XOR U12274 ( .A(n12657), .B(p_input[6731]), .Z(n12659) );
  XOR U12275 ( .A(n12661), .B(n12662), .Z(n12657) );
  AND U12276 ( .A(n12663), .B(n12664), .Z(n12662) );
  XNOR U12277 ( .A(p_input[6762]), .B(n12661), .Z(n12664) );
  XOR U12278 ( .A(n12661), .B(p_input[6730]), .Z(n12663) );
  XOR U12279 ( .A(n12665), .B(n12666), .Z(n12661) );
  AND U12280 ( .A(n12667), .B(n12668), .Z(n12666) );
  XNOR U12281 ( .A(p_input[6761]), .B(n12665), .Z(n12668) );
  XOR U12282 ( .A(n12665), .B(p_input[6729]), .Z(n12667) );
  XOR U12283 ( .A(n12669), .B(n12670), .Z(n12665) );
  AND U12284 ( .A(n12671), .B(n12672), .Z(n12670) );
  XNOR U12285 ( .A(p_input[6760]), .B(n12669), .Z(n12672) );
  XOR U12286 ( .A(n12669), .B(p_input[6728]), .Z(n12671) );
  XOR U12287 ( .A(n12673), .B(n12674), .Z(n12669) );
  AND U12288 ( .A(n12675), .B(n12676), .Z(n12674) );
  XNOR U12289 ( .A(p_input[6759]), .B(n12673), .Z(n12676) );
  XOR U12290 ( .A(n12673), .B(p_input[6727]), .Z(n12675) );
  XOR U12291 ( .A(n12677), .B(n12678), .Z(n12673) );
  AND U12292 ( .A(n12679), .B(n12680), .Z(n12678) );
  XNOR U12293 ( .A(p_input[6758]), .B(n12677), .Z(n12680) );
  XOR U12294 ( .A(n12677), .B(p_input[6726]), .Z(n12679) );
  XOR U12295 ( .A(n12681), .B(n12682), .Z(n12677) );
  AND U12296 ( .A(n12683), .B(n12684), .Z(n12682) );
  XNOR U12297 ( .A(p_input[6757]), .B(n12681), .Z(n12684) );
  XOR U12298 ( .A(n12681), .B(p_input[6725]), .Z(n12683) );
  XOR U12299 ( .A(n12685), .B(n12686), .Z(n12681) );
  AND U12300 ( .A(n12687), .B(n12688), .Z(n12686) );
  XNOR U12301 ( .A(p_input[6756]), .B(n12685), .Z(n12688) );
  XOR U12302 ( .A(n12685), .B(p_input[6724]), .Z(n12687) );
  XOR U12303 ( .A(n12689), .B(n12690), .Z(n12685) );
  AND U12304 ( .A(n12691), .B(n12692), .Z(n12690) );
  XNOR U12305 ( .A(p_input[6755]), .B(n12689), .Z(n12692) );
  XOR U12306 ( .A(n12689), .B(p_input[6723]), .Z(n12691) );
  XOR U12307 ( .A(n12693), .B(n12694), .Z(n12689) );
  AND U12308 ( .A(n12695), .B(n12696), .Z(n12694) );
  XNOR U12309 ( .A(p_input[6754]), .B(n12693), .Z(n12696) );
  XOR U12310 ( .A(n12693), .B(p_input[6722]), .Z(n12695) );
  XNOR U12311 ( .A(n12697), .B(n12698), .Z(n12693) );
  AND U12312 ( .A(n12699), .B(n12700), .Z(n12698) );
  XOR U12313 ( .A(p_input[6753]), .B(n12697), .Z(n12700) );
  XNOR U12314 ( .A(p_input[6721]), .B(n12697), .Z(n12699) );
  AND U12315 ( .A(p_input[6752]), .B(n12701), .Z(n12697) );
  IV U12316 ( .A(p_input[6720]), .Z(n12701) );
  XNOR U12317 ( .A(p_input[6656]), .B(n12702), .Z(n12295) );
  AND U12318 ( .A(n260), .B(n12703), .Z(n12702) );
  XOR U12319 ( .A(p_input[6688]), .B(p_input[6656]), .Z(n12703) );
  XOR U12320 ( .A(n12704), .B(n12705), .Z(n260) );
  AND U12321 ( .A(n12706), .B(n12707), .Z(n12705) );
  XNOR U12322 ( .A(p_input[6719]), .B(n12704), .Z(n12707) );
  XOR U12323 ( .A(n12704), .B(p_input[6687]), .Z(n12706) );
  XOR U12324 ( .A(n12708), .B(n12709), .Z(n12704) );
  AND U12325 ( .A(n12710), .B(n12711), .Z(n12709) );
  XNOR U12326 ( .A(p_input[6718]), .B(n12708), .Z(n12711) );
  XNOR U12327 ( .A(n12708), .B(n12310), .Z(n12710) );
  IV U12328 ( .A(p_input[6686]), .Z(n12310) );
  XOR U12329 ( .A(n12712), .B(n12713), .Z(n12708) );
  AND U12330 ( .A(n12714), .B(n12715), .Z(n12713) );
  XNOR U12331 ( .A(p_input[6717]), .B(n12712), .Z(n12715) );
  XNOR U12332 ( .A(n12712), .B(n12319), .Z(n12714) );
  IV U12333 ( .A(p_input[6685]), .Z(n12319) );
  XOR U12334 ( .A(n12716), .B(n12717), .Z(n12712) );
  AND U12335 ( .A(n12718), .B(n12719), .Z(n12717) );
  XNOR U12336 ( .A(p_input[6716]), .B(n12716), .Z(n12719) );
  XNOR U12337 ( .A(n12716), .B(n12328), .Z(n12718) );
  IV U12338 ( .A(p_input[6684]), .Z(n12328) );
  XOR U12339 ( .A(n12720), .B(n12721), .Z(n12716) );
  AND U12340 ( .A(n12722), .B(n12723), .Z(n12721) );
  XNOR U12341 ( .A(p_input[6715]), .B(n12720), .Z(n12723) );
  XNOR U12342 ( .A(n12720), .B(n12337), .Z(n12722) );
  IV U12343 ( .A(p_input[6683]), .Z(n12337) );
  XOR U12344 ( .A(n12724), .B(n12725), .Z(n12720) );
  AND U12345 ( .A(n12726), .B(n12727), .Z(n12725) );
  XNOR U12346 ( .A(p_input[6714]), .B(n12724), .Z(n12727) );
  XNOR U12347 ( .A(n12724), .B(n12346), .Z(n12726) );
  IV U12348 ( .A(p_input[6682]), .Z(n12346) );
  XOR U12349 ( .A(n12728), .B(n12729), .Z(n12724) );
  AND U12350 ( .A(n12730), .B(n12731), .Z(n12729) );
  XNOR U12351 ( .A(p_input[6713]), .B(n12728), .Z(n12731) );
  XNOR U12352 ( .A(n12728), .B(n12355), .Z(n12730) );
  IV U12353 ( .A(p_input[6681]), .Z(n12355) );
  XOR U12354 ( .A(n12732), .B(n12733), .Z(n12728) );
  AND U12355 ( .A(n12734), .B(n12735), .Z(n12733) );
  XNOR U12356 ( .A(p_input[6712]), .B(n12732), .Z(n12735) );
  XNOR U12357 ( .A(n12732), .B(n12364), .Z(n12734) );
  IV U12358 ( .A(p_input[6680]), .Z(n12364) );
  XOR U12359 ( .A(n12736), .B(n12737), .Z(n12732) );
  AND U12360 ( .A(n12738), .B(n12739), .Z(n12737) );
  XNOR U12361 ( .A(p_input[6711]), .B(n12736), .Z(n12739) );
  XNOR U12362 ( .A(n12736), .B(n12373), .Z(n12738) );
  IV U12363 ( .A(p_input[6679]), .Z(n12373) );
  XOR U12364 ( .A(n12740), .B(n12741), .Z(n12736) );
  AND U12365 ( .A(n12742), .B(n12743), .Z(n12741) );
  XNOR U12366 ( .A(p_input[6710]), .B(n12740), .Z(n12743) );
  XNOR U12367 ( .A(n12740), .B(n12382), .Z(n12742) );
  IV U12368 ( .A(p_input[6678]), .Z(n12382) );
  XOR U12369 ( .A(n12744), .B(n12745), .Z(n12740) );
  AND U12370 ( .A(n12746), .B(n12747), .Z(n12745) );
  XNOR U12371 ( .A(p_input[6709]), .B(n12744), .Z(n12747) );
  XNOR U12372 ( .A(n12744), .B(n12391), .Z(n12746) );
  IV U12373 ( .A(p_input[6677]), .Z(n12391) );
  XOR U12374 ( .A(n12748), .B(n12749), .Z(n12744) );
  AND U12375 ( .A(n12750), .B(n12751), .Z(n12749) );
  XNOR U12376 ( .A(p_input[6708]), .B(n12748), .Z(n12751) );
  XNOR U12377 ( .A(n12748), .B(n12400), .Z(n12750) );
  IV U12378 ( .A(p_input[6676]), .Z(n12400) );
  XOR U12379 ( .A(n12752), .B(n12753), .Z(n12748) );
  AND U12380 ( .A(n12754), .B(n12755), .Z(n12753) );
  XNOR U12381 ( .A(p_input[6707]), .B(n12752), .Z(n12755) );
  XNOR U12382 ( .A(n12752), .B(n12409), .Z(n12754) );
  IV U12383 ( .A(p_input[6675]), .Z(n12409) );
  XOR U12384 ( .A(n12756), .B(n12757), .Z(n12752) );
  AND U12385 ( .A(n12758), .B(n12759), .Z(n12757) );
  XNOR U12386 ( .A(p_input[6706]), .B(n12756), .Z(n12759) );
  XNOR U12387 ( .A(n12756), .B(n12418), .Z(n12758) );
  IV U12388 ( .A(p_input[6674]), .Z(n12418) );
  XOR U12389 ( .A(n12760), .B(n12761), .Z(n12756) );
  AND U12390 ( .A(n12762), .B(n12763), .Z(n12761) );
  XNOR U12391 ( .A(p_input[6705]), .B(n12760), .Z(n12763) );
  XNOR U12392 ( .A(n12760), .B(n12427), .Z(n12762) );
  IV U12393 ( .A(p_input[6673]), .Z(n12427) );
  XOR U12394 ( .A(n12764), .B(n12765), .Z(n12760) );
  AND U12395 ( .A(n12766), .B(n12767), .Z(n12765) );
  XNOR U12396 ( .A(p_input[6704]), .B(n12764), .Z(n12767) );
  XNOR U12397 ( .A(n12764), .B(n12436), .Z(n12766) );
  IV U12398 ( .A(p_input[6672]), .Z(n12436) );
  XOR U12399 ( .A(n12768), .B(n12769), .Z(n12764) );
  AND U12400 ( .A(n12770), .B(n12771), .Z(n12769) );
  XNOR U12401 ( .A(p_input[6703]), .B(n12768), .Z(n12771) );
  XNOR U12402 ( .A(n12768), .B(n12445), .Z(n12770) );
  IV U12403 ( .A(p_input[6671]), .Z(n12445) );
  XOR U12404 ( .A(n12772), .B(n12773), .Z(n12768) );
  AND U12405 ( .A(n12774), .B(n12775), .Z(n12773) );
  XNOR U12406 ( .A(p_input[6702]), .B(n12772), .Z(n12775) );
  XNOR U12407 ( .A(n12772), .B(n12454), .Z(n12774) );
  IV U12408 ( .A(p_input[6670]), .Z(n12454) );
  XOR U12409 ( .A(n12776), .B(n12777), .Z(n12772) );
  AND U12410 ( .A(n12778), .B(n12779), .Z(n12777) );
  XNOR U12411 ( .A(p_input[6701]), .B(n12776), .Z(n12779) );
  XNOR U12412 ( .A(n12776), .B(n12463), .Z(n12778) );
  IV U12413 ( .A(p_input[6669]), .Z(n12463) );
  XOR U12414 ( .A(n12780), .B(n12781), .Z(n12776) );
  AND U12415 ( .A(n12782), .B(n12783), .Z(n12781) );
  XNOR U12416 ( .A(p_input[6700]), .B(n12780), .Z(n12783) );
  XNOR U12417 ( .A(n12780), .B(n12472), .Z(n12782) );
  IV U12418 ( .A(p_input[6668]), .Z(n12472) );
  XOR U12419 ( .A(n12784), .B(n12785), .Z(n12780) );
  AND U12420 ( .A(n12786), .B(n12787), .Z(n12785) );
  XNOR U12421 ( .A(p_input[6699]), .B(n12784), .Z(n12787) );
  XNOR U12422 ( .A(n12784), .B(n12481), .Z(n12786) );
  IV U12423 ( .A(p_input[6667]), .Z(n12481) );
  XOR U12424 ( .A(n12788), .B(n12789), .Z(n12784) );
  AND U12425 ( .A(n12790), .B(n12791), .Z(n12789) );
  XNOR U12426 ( .A(p_input[6698]), .B(n12788), .Z(n12791) );
  XNOR U12427 ( .A(n12788), .B(n12490), .Z(n12790) );
  IV U12428 ( .A(p_input[6666]), .Z(n12490) );
  XOR U12429 ( .A(n12792), .B(n12793), .Z(n12788) );
  AND U12430 ( .A(n12794), .B(n12795), .Z(n12793) );
  XNOR U12431 ( .A(p_input[6697]), .B(n12792), .Z(n12795) );
  XNOR U12432 ( .A(n12792), .B(n12499), .Z(n12794) );
  IV U12433 ( .A(p_input[6665]), .Z(n12499) );
  XOR U12434 ( .A(n12796), .B(n12797), .Z(n12792) );
  AND U12435 ( .A(n12798), .B(n12799), .Z(n12797) );
  XNOR U12436 ( .A(p_input[6696]), .B(n12796), .Z(n12799) );
  XNOR U12437 ( .A(n12796), .B(n12508), .Z(n12798) );
  IV U12438 ( .A(p_input[6664]), .Z(n12508) );
  XOR U12439 ( .A(n12800), .B(n12801), .Z(n12796) );
  AND U12440 ( .A(n12802), .B(n12803), .Z(n12801) );
  XNOR U12441 ( .A(p_input[6695]), .B(n12800), .Z(n12803) );
  XNOR U12442 ( .A(n12800), .B(n12517), .Z(n12802) );
  IV U12443 ( .A(p_input[6663]), .Z(n12517) );
  XOR U12444 ( .A(n12804), .B(n12805), .Z(n12800) );
  AND U12445 ( .A(n12806), .B(n12807), .Z(n12805) );
  XNOR U12446 ( .A(p_input[6694]), .B(n12804), .Z(n12807) );
  XNOR U12447 ( .A(n12804), .B(n12526), .Z(n12806) );
  IV U12448 ( .A(p_input[6662]), .Z(n12526) );
  XOR U12449 ( .A(n12808), .B(n12809), .Z(n12804) );
  AND U12450 ( .A(n12810), .B(n12811), .Z(n12809) );
  XNOR U12451 ( .A(p_input[6693]), .B(n12808), .Z(n12811) );
  XNOR U12452 ( .A(n12808), .B(n12535), .Z(n12810) );
  IV U12453 ( .A(p_input[6661]), .Z(n12535) );
  XOR U12454 ( .A(n12812), .B(n12813), .Z(n12808) );
  AND U12455 ( .A(n12814), .B(n12815), .Z(n12813) );
  XNOR U12456 ( .A(p_input[6692]), .B(n12812), .Z(n12815) );
  XNOR U12457 ( .A(n12812), .B(n12544), .Z(n12814) );
  IV U12458 ( .A(p_input[6660]), .Z(n12544) );
  XOR U12459 ( .A(n12816), .B(n12817), .Z(n12812) );
  AND U12460 ( .A(n12818), .B(n12819), .Z(n12817) );
  XNOR U12461 ( .A(p_input[6691]), .B(n12816), .Z(n12819) );
  XNOR U12462 ( .A(n12816), .B(n12553), .Z(n12818) );
  IV U12463 ( .A(p_input[6659]), .Z(n12553) );
  XOR U12464 ( .A(n12820), .B(n12821), .Z(n12816) );
  AND U12465 ( .A(n12822), .B(n12823), .Z(n12821) );
  XNOR U12466 ( .A(p_input[6690]), .B(n12820), .Z(n12823) );
  XNOR U12467 ( .A(n12820), .B(n12562), .Z(n12822) );
  IV U12468 ( .A(p_input[6658]), .Z(n12562) );
  XNOR U12469 ( .A(n12824), .B(n12825), .Z(n12820) );
  AND U12470 ( .A(n12826), .B(n12827), .Z(n12825) );
  XOR U12471 ( .A(p_input[6689]), .B(n12824), .Z(n12827) );
  XNOR U12472 ( .A(p_input[6657]), .B(n12824), .Z(n12826) );
  AND U12473 ( .A(p_input[6688]), .B(n12828), .Z(n12824) );
  IV U12474 ( .A(p_input[6656]), .Z(n12828) );
  XOR U12475 ( .A(n12829), .B(n12830), .Z(n9185) );
  AND U12476 ( .A(n1000), .B(n12831), .Z(n12830) );
  XNOR U12477 ( .A(n12832), .B(n12829), .Z(n12831) );
  XOR U12478 ( .A(n12833), .B(n12834), .Z(n1000) );
  AND U12479 ( .A(n12835), .B(n12836), .Z(n12834) );
  XOR U12480 ( .A(n12833), .B(n9200), .Z(n12836) );
  XOR U12481 ( .A(n12837), .B(n12838), .Z(n9200) );
  AND U12482 ( .A(n831), .B(n12839), .Z(n12838) );
  XOR U12483 ( .A(n12840), .B(n12837), .Z(n12839) );
  XNOR U12484 ( .A(n9197), .B(n12833), .Z(n12835) );
  XOR U12485 ( .A(n12841), .B(n12842), .Z(n9197) );
  AND U12486 ( .A(n828), .B(n12843), .Z(n12842) );
  XOR U12487 ( .A(n12844), .B(n12841), .Z(n12843) );
  XOR U12488 ( .A(n12845), .B(n12846), .Z(n12833) );
  AND U12489 ( .A(n12847), .B(n12848), .Z(n12846) );
  XOR U12490 ( .A(n12845), .B(n9212), .Z(n12848) );
  XOR U12491 ( .A(n12849), .B(n12850), .Z(n9212) );
  AND U12492 ( .A(n831), .B(n12851), .Z(n12850) );
  XOR U12493 ( .A(n12852), .B(n12849), .Z(n12851) );
  XNOR U12494 ( .A(n9209), .B(n12845), .Z(n12847) );
  XOR U12495 ( .A(n12853), .B(n12854), .Z(n9209) );
  AND U12496 ( .A(n828), .B(n12855), .Z(n12854) );
  XOR U12497 ( .A(n12856), .B(n12853), .Z(n12855) );
  XOR U12498 ( .A(n12857), .B(n12858), .Z(n12845) );
  AND U12499 ( .A(n12859), .B(n12860), .Z(n12858) );
  XOR U12500 ( .A(n12857), .B(n9224), .Z(n12860) );
  XOR U12501 ( .A(n12861), .B(n12862), .Z(n9224) );
  AND U12502 ( .A(n831), .B(n12863), .Z(n12862) );
  XOR U12503 ( .A(n12864), .B(n12861), .Z(n12863) );
  XNOR U12504 ( .A(n9221), .B(n12857), .Z(n12859) );
  XOR U12505 ( .A(n12865), .B(n12866), .Z(n9221) );
  AND U12506 ( .A(n828), .B(n12867), .Z(n12866) );
  XOR U12507 ( .A(n12868), .B(n12865), .Z(n12867) );
  XOR U12508 ( .A(n12869), .B(n12870), .Z(n12857) );
  AND U12509 ( .A(n12871), .B(n12872), .Z(n12870) );
  XOR U12510 ( .A(n12869), .B(n9236), .Z(n12872) );
  XOR U12511 ( .A(n12873), .B(n12874), .Z(n9236) );
  AND U12512 ( .A(n831), .B(n12875), .Z(n12874) );
  XOR U12513 ( .A(n12876), .B(n12873), .Z(n12875) );
  XNOR U12514 ( .A(n9233), .B(n12869), .Z(n12871) );
  XOR U12515 ( .A(n12877), .B(n12878), .Z(n9233) );
  AND U12516 ( .A(n828), .B(n12879), .Z(n12878) );
  XOR U12517 ( .A(n12880), .B(n12877), .Z(n12879) );
  XOR U12518 ( .A(n12881), .B(n12882), .Z(n12869) );
  AND U12519 ( .A(n12883), .B(n12884), .Z(n12882) );
  XOR U12520 ( .A(n12881), .B(n9248), .Z(n12884) );
  XOR U12521 ( .A(n12885), .B(n12886), .Z(n9248) );
  AND U12522 ( .A(n831), .B(n12887), .Z(n12886) );
  XOR U12523 ( .A(n12888), .B(n12885), .Z(n12887) );
  XNOR U12524 ( .A(n9245), .B(n12881), .Z(n12883) );
  XOR U12525 ( .A(n12889), .B(n12890), .Z(n9245) );
  AND U12526 ( .A(n828), .B(n12891), .Z(n12890) );
  XOR U12527 ( .A(n12892), .B(n12889), .Z(n12891) );
  XOR U12528 ( .A(n12893), .B(n12894), .Z(n12881) );
  AND U12529 ( .A(n12895), .B(n12896), .Z(n12894) );
  XOR U12530 ( .A(n12893), .B(n9260), .Z(n12896) );
  XOR U12531 ( .A(n12897), .B(n12898), .Z(n9260) );
  AND U12532 ( .A(n831), .B(n12899), .Z(n12898) );
  XOR U12533 ( .A(n12900), .B(n12897), .Z(n12899) );
  XNOR U12534 ( .A(n9257), .B(n12893), .Z(n12895) );
  XOR U12535 ( .A(n12901), .B(n12902), .Z(n9257) );
  AND U12536 ( .A(n828), .B(n12903), .Z(n12902) );
  XOR U12537 ( .A(n12904), .B(n12901), .Z(n12903) );
  XOR U12538 ( .A(n12905), .B(n12906), .Z(n12893) );
  AND U12539 ( .A(n12907), .B(n12908), .Z(n12906) );
  XOR U12540 ( .A(n12905), .B(n9272), .Z(n12908) );
  XOR U12541 ( .A(n12909), .B(n12910), .Z(n9272) );
  AND U12542 ( .A(n831), .B(n12911), .Z(n12910) );
  XOR U12543 ( .A(n12912), .B(n12909), .Z(n12911) );
  XNOR U12544 ( .A(n9269), .B(n12905), .Z(n12907) );
  XOR U12545 ( .A(n12913), .B(n12914), .Z(n9269) );
  AND U12546 ( .A(n828), .B(n12915), .Z(n12914) );
  XOR U12547 ( .A(n12916), .B(n12913), .Z(n12915) );
  XOR U12548 ( .A(n12917), .B(n12918), .Z(n12905) );
  AND U12549 ( .A(n12919), .B(n12920), .Z(n12918) );
  XOR U12550 ( .A(n12917), .B(n9284), .Z(n12920) );
  XOR U12551 ( .A(n12921), .B(n12922), .Z(n9284) );
  AND U12552 ( .A(n831), .B(n12923), .Z(n12922) );
  XOR U12553 ( .A(n12924), .B(n12921), .Z(n12923) );
  XNOR U12554 ( .A(n9281), .B(n12917), .Z(n12919) );
  XOR U12555 ( .A(n12925), .B(n12926), .Z(n9281) );
  AND U12556 ( .A(n828), .B(n12927), .Z(n12926) );
  XOR U12557 ( .A(n12928), .B(n12925), .Z(n12927) );
  XOR U12558 ( .A(n12929), .B(n12930), .Z(n12917) );
  AND U12559 ( .A(n12931), .B(n12932), .Z(n12930) );
  XOR U12560 ( .A(n12929), .B(n9296), .Z(n12932) );
  XOR U12561 ( .A(n12933), .B(n12934), .Z(n9296) );
  AND U12562 ( .A(n831), .B(n12935), .Z(n12934) );
  XOR U12563 ( .A(n12936), .B(n12933), .Z(n12935) );
  XNOR U12564 ( .A(n9293), .B(n12929), .Z(n12931) );
  XOR U12565 ( .A(n12937), .B(n12938), .Z(n9293) );
  AND U12566 ( .A(n828), .B(n12939), .Z(n12938) );
  XOR U12567 ( .A(n12940), .B(n12937), .Z(n12939) );
  XOR U12568 ( .A(n12941), .B(n12942), .Z(n12929) );
  AND U12569 ( .A(n12943), .B(n12944), .Z(n12942) );
  XOR U12570 ( .A(n12941), .B(n9308), .Z(n12944) );
  XOR U12571 ( .A(n12945), .B(n12946), .Z(n9308) );
  AND U12572 ( .A(n831), .B(n12947), .Z(n12946) );
  XOR U12573 ( .A(n12948), .B(n12945), .Z(n12947) );
  XNOR U12574 ( .A(n9305), .B(n12941), .Z(n12943) );
  XOR U12575 ( .A(n12949), .B(n12950), .Z(n9305) );
  AND U12576 ( .A(n828), .B(n12951), .Z(n12950) );
  XOR U12577 ( .A(n12952), .B(n12949), .Z(n12951) );
  XOR U12578 ( .A(n12953), .B(n12954), .Z(n12941) );
  AND U12579 ( .A(n12955), .B(n12956), .Z(n12954) );
  XOR U12580 ( .A(n12953), .B(n9320), .Z(n12956) );
  XOR U12581 ( .A(n12957), .B(n12958), .Z(n9320) );
  AND U12582 ( .A(n831), .B(n12959), .Z(n12958) );
  XOR U12583 ( .A(n12960), .B(n12957), .Z(n12959) );
  XNOR U12584 ( .A(n9317), .B(n12953), .Z(n12955) );
  XOR U12585 ( .A(n12961), .B(n12962), .Z(n9317) );
  AND U12586 ( .A(n828), .B(n12963), .Z(n12962) );
  XOR U12587 ( .A(n12964), .B(n12961), .Z(n12963) );
  XOR U12588 ( .A(n12965), .B(n12966), .Z(n12953) );
  AND U12589 ( .A(n12967), .B(n12968), .Z(n12966) );
  XOR U12590 ( .A(n12965), .B(n9332), .Z(n12968) );
  XOR U12591 ( .A(n12969), .B(n12970), .Z(n9332) );
  AND U12592 ( .A(n831), .B(n12971), .Z(n12970) );
  XOR U12593 ( .A(n12972), .B(n12969), .Z(n12971) );
  XNOR U12594 ( .A(n9329), .B(n12965), .Z(n12967) );
  XOR U12595 ( .A(n12973), .B(n12974), .Z(n9329) );
  AND U12596 ( .A(n828), .B(n12975), .Z(n12974) );
  XOR U12597 ( .A(n12976), .B(n12973), .Z(n12975) );
  XOR U12598 ( .A(n12977), .B(n12978), .Z(n12965) );
  AND U12599 ( .A(n12979), .B(n12980), .Z(n12978) );
  XOR U12600 ( .A(n12977), .B(n9344), .Z(n12980) );
  XOR U12601 ( .A(n12981), .B(n12982), .Z(n9344) );
  AND U12602 ( .A(n831), .B(n12983), .Z(n12982) );
  XOR U12603 ( .A(n12984), .B(n12981), .Z(n12983) );
  XNOR U12604 ( .A(n9341), .B(n12977), .Z(n12979) );
  XOR U12605 ( .A(n12985), .B(n12986), .Z(n9341) );
  AND U12606 ( .A(n828), .B(n12987), .Z(n12986) );
  XOR U12607 ( .A(n12988), .B(n12985), .Z(n12987) );
  XOR U12608 ( .A(n12989), .B(n12990), .Z(n12977) );
  AND U12609 ( .A(n12991), .B(n12992), .Z(n12990) );
  XOR U12610 ( .A(n12989), .B(n9356), .Z(n12992) );
  XOR U12611 ( .A(n12993), .B(n12994), .Z(n9356) );
  AND U12612 ( .A(n831), .B(n12995), .Z(n12994) );
  XOR U12613 ( .A(n12996), .B(n12993), .Z(n12995) );
  XNOR U12614 ( .A(n9353), .B(n12989), .Z(n12991) );
  XOR U12615 ( .A(n12997), .B(n12998), .Z(n9353) );
  AND U12616 ( .A(n828), .B(n12999), .Z(n12998) );
  XOR U12617 ( .A(n13000), .B(n12997), .Z(n12999) );
  XOR U12618 ( .A(n13001), .B(n13002), .Z(n12989) );
  AND U12619 ( .A(n13003), .B(n13004), .Z(n13002) );
  XOR U12620 ( .A(n13001), .B(n9368), .Z(n13004) );
  XOR U12621 ( .A(n13005), .B(n13006), .Z(n9368) );
  AND U12622 ( .A(n831), .B(n13007), .Z(n13006) );
  XOR U12623 ( .A(n13008), .B(n13005), .Z(n13007) );
  XNOR U12624 ( .A(n9365), .B(n13001), .Z(n13003) );
  XOR U12625 ( .A(n13009), .B(n13010), .Z(n9365) );
  AND U12626 ( .A(n828), .B(n13011), .Z(n13010) );
  XOR U12627 ( .A(n13012), .B(n13009), .Z(n13011) );
  XOR U12628 ( .A(n13013), .B(n13014), .Z(n13001) );
  AND U12629 ( .A(n13015), .B(n13016), .Z(n13014) );
  XOR U12630 ( .A(n13013), .B(n9380), .Z(n13016) );
  XOR U12631 ( .A(n13017), .B(n13018), .Z(n9380) );
  AND U12632 ( .A(n831), .B(n13019), .Z(n13018) );
  XOR U12633 ( .A(n13020), .B(n13017), .Z(n13019) );
  XNOR U12634 ( .A(n9377), .B(n13013), .Z(n13015) );
  XOR U12635 ( .A(n13021), .B(n13022), .Z(n9377) );
  AND U12636 ( .A(n828), .B(n13023), .Z(n13022) );
  XOR U12637 ( .A(n13024), .B(n13021), .Z(n13023) );
  XOR U12638 ( .A(n13025), .B(n13026), .Z(n13013) );
  AND U12639 ( .A(n13027), .B(n13028), .Z(n13026) );
  XOR U12640 ( .A(n13025), .B(n9392), .Z(n13028) );
  XOR U12641 ( .A(n13029), .B(n13030), .Z(n9392) );
  AND U12642 ( .A(n831), .B(n13031), .Z(n13030) );
  XOR U12643 ( .A(n13032), .B(n13029), .Z(n13031) );
  XNOR U12644 ( .A(n9389), .B(n13025), .Z(n13027) );
  XOR U12645 ( .A(n13033), .B(n13034), .Z(n9389) );
  AND U12646 ( .A(n828), .B(n13035), .Z(n13034) );
  XOR U12647 ( .A(n13036), .B(n13033), .Z(n13035) );
  XOR U12648 ( .A(n13037), .B(n13038), .Z(n13025) );
  AND U12649 ( .A(n13039), .B(n13040), .Z(n13038) );
  XOR U12650 ( .A(n13037), .B(n9404), .Z(n13040) );
  XOR U12651 ( .A(n13041), .B(n13042), .Z(n9404) );
  AND U12652 ( .A(n831), .B(n13043), .Z(n13042) );
  XOR U12653 ( .A(n13044), .B(n13041), .Z(n13043) );
  XNOR U12654 ( .A(n9401), .B(n13037), .Z(n13039) );
  XOR U12655 ( .A(n13045), .B(n13046), .Z(n9401) );
  AND U12656 ( .A(n828), .B(n13047), .Z(n13046) );
  XOR U12657 ( .A(n13048), .B(n13045), .Z(n13047) );
  XOR U12658 ( .A(n13049), .B(n13050), .Z(n13037) );
  AND U12659 ( .A(n13051), .B(n13052), .Z(n13050) );
  XOR U12660 ( .A(n13049), .B(n9416), .Z(n13052) );
  XOR U12661 ( .A(n13053), .B(n13054), .Z(n9416) );
  AND U12662 ( .A(n831), .B(n13055), .Z(n13054) );
  XOR U12663 ( .A(n13056), .B(n13053), .Z(n13055) );
  XNOR U12664 ( .A(n9413), .B(n13049), .Z(n13051) );
  XOR U12665 ( .A(n13057), .B(n13058), .Z(n9413) );
  AND U12666 ( .A(n828), .B(n13059), .Z(n13058) );
  XOR U12667 ( .A(n13060), .B(n13057), .Z(n13059) );
  XOR U12668 ( .A(n13061), .B(n13062), .Z(n13049) );
  AND U12669 ( .A(n13063), .B(n13064), .Z(n13062) );
  XOR U12670 ( .A(n13061), .B(n9428), .Z(n13064) );
  XOR U12671 ( .A(n13065), .B(n13066), .Z(n9428) );
  AND U12672 ( .A(n831), .B(n13067), .Z(n13066) );
  XOR U12673 ( .A(n13068), .B(n13065), .Z(n13067) );
  XNOR U12674 ( .A(n9425), .B(n13061), .Z(n13063) );
  XOR U12675 ( .A(n13069), .B(n13070), .Z(n9425) );
  AND U12676 ( .A(n828), .B(n13071), .Z(n13070) );
  XOR U12677 ( .A(n13072), .B(n13069), .Z(n13071) );
  XOR U12678 ( .A(n13073), .B(n13074), .Z(n13061) );
  AND U12679 ( .A(n13075), .B(n13076), .Z(n13074) );
  XOR U12680 ( .A(n13073), .B(n9440), .Z(n13076) );
  XOR U12681 ( .A(n13077), .B(n13078), .Z(n9440) );
  AND U12682 ( .A(n831), .B(n13079), .Z(n13078) );
  XOR U12683 ( .A(n13080), .B(n13077), .Z(n13079) );
  XNOR U12684 ( .A(n9437), .B(n13073), .Z(n13075) );
  XOR U12685 ( .A(n13081), .B(n13082), .Z(n9437) );
  AND U12686 ( .A(n828), .B(n13083), .Z(n13082) );
  XOR U12687 ( .A(n13084), .B(n13081), .Z(n13083) );
  XOR U12688 ( .A(n13085), .B(n13086), .Z(n13073) );
  AND U12689 ( .A(n13087), .B(n13088), .Z(n13086) );
  XOR U12690 ( .A(n13085), .B(n9452), .Z(n13088) );
  XOR U12691 ( .A(n13089), .B(n13090), .Z(n9452) );
  AND U12692 ( .A(n831), .B(n13091), .Z(n13090) );
  XOR U12693 ( .A(n13092), .B(n13089), .Z(n13091) );
  XNOR U12694 ( .A(n9449), .B(n13085), .Z(n13087) );
  XOR U12695 ( .A(n13093), .B(n13094), .Z(n9449) );
  AND U12696 ( .A(n828), .B(n13095), .Z(n13094) );
  XOR U12697 ( .A(n13096), .B(n13093), .Z(n13095) );
  XOR U12698 ( .A(n13097), .B(n13098), .Z(n13085) );
  AND U12699 ( .A(n13099), .B(n13100), .Z(n13098) );
  XOR U12700 ( .A(n13097), .B(n9464), .Z(n13100) );
  XOR U12701 ( .A(n13101), .B(n13102), .Z(n9464) );
  AND U12702 ( .A(n831), .B(n13103), .Z(n13102) );
  XOR U12703 ( .A(n13104), .B(n13101), .Z(n13103) );
  XNOR U12704 ( .A(n9461), .B(n13097), .Z(n13099) );
  XOR U12705 ( .A(n13105), .B(n13106), .Z(n9461) );
  AND U12706 ( .A(n828), .B(n13107), .Z(n13106) );
  XOR U12707 ( .A(n13108), .B(n13105), .Z(n13107) );
  XOR U12708 ( .A(n13109), .B(n13110), .Z(n13097) );
  AND U12709 ( .A(n13111), .B(n13112), .Z(n13110) );
  XOR U12710 ( .A(n13109), .B(n9476), .Z(n13112) );
  XOR U12711 ( .A(n13113), .B(n13114), .Z(n9476) );
  AND U12712 ( .A(n831), .B(n13115), .Z(n13114) );
  XOR U12713 ( .A(n13116), .B(n13113), .Z(n13115) );
  XNOR U12714 ( .A(n9473), .B(n13109), .Z(n13111) );
  XOR U12715 ( .A(n13117), .B(n13118), .Z(n9473) );
  AND U12716 ( .A(n828), .B(n13119), .Z(n13118) );
  XOR U12717 ( .A(n13120), .B(n13117), .Z(n13119) );
  XOR U12718 ( .A(n13121), .B(n13122), .Z(n13109) );
  AND U12719 ( .A(n13123), .B(n13124), .Z(n13122) );
  XOR U12720 ( .A(n13121), .B(n9488), .Z(n13124) );
  XOR U12721 ( .A(n13125), .B(n13126), .Z(n9488) );
  AND U12722 ( .A(n831), .B(n13127), .Z(n13126) );
  XOR U12723 ( .A(n13128), .B(n13125), .Z(n13127) );
  XNOR U12724 ( .A(n9485), .B(n13121), .Z(n13123) );
  XOR U12725 ( .A(n13129), .B(n13130), .Z(n9485) );
  AND U12726 ( .A(n828), .B(n13131), .Z(n13130) );
  XOR U12727 ( .A(n13132), .B(n13129), .Z(n13131) );
  XOR U12728 ( .A(n13133), .B(n13134), .Z(n13121) );
  AND U12729 ( .A(n13135), .B(n13136), .Z(n13134) );
  XOR U12730 ( .A(n13133), .B(n9500), .Z(n13136) );
  XOR U12731 ( .A(n13137), .B(n13138), .Z(n9500) );
  AND U12732 ( .A(n831), .B(n13139), .Z(n13138) );
  XOR U12733 ( .A(n13140), .B(n13137), .Z(n13139) );
  XNOR U12734 ( .A(n9497), .B(n13133), .Z(n13135) );
  XOR U12735 ( .A(n13141), .B(n13142), .Z(n9497) );
  AND U12736 ( .A(n828), .B(n13143), .Z(n13142) );
  XOR U12737 ( .A(n13144), .B(n13141), .Z(n13143) );
  XOR U12738 ( .A(n13145), .B(n13146), .Z(n13133) );
  AND U12739 ( .A(n13147), .B(n13148), .Z(n13146) );
  XOR U12740 ( .A(n13145), .B(n9512), .Z(n13148) );
  XOR U12741 ( .A(n13149), .B(n13150), .Z(n9512) );
  AND U12742 ( .A(n831), .B(n13151), .Z(n13150) );
  XOR U12743 ( .A(n13152), .B(n13149), .Z(n13151) );
  XNOR U12744 ( .A(n9509), .B(n13145), .Z(n13147) );
  XOR U12745 ( .A(n13153), .B(n13154), .Z(n9509) );
  AND U12746 ( .A(n828), .B(n13155), .Z(n13154) );
  XOR U12747 ( .A(n13156), .B(n13153), .Z(n13155) );
  XOR U12748 ( .A(n13157), .B(n13158), .Z(n13145) );
  AND U12749 ( .A(n13159), .B(n13160), .Z(n13158) );
  XOR U12750 ( .A(n13157), .B(n9524), .Z(n13160) );
  XOR U12751 ( .A(n13161), .B(n13162), .Z(n9524) );
  AND U12752 ( .A(n831), .B(n13163), .Z(n13162) );
  XOR U12753 ( .A(n13164), .B(n13161), .Z(n13163) );
  XNOR U12754 ( .A(n9521), .B(n13157), .Z(n13159) );
  XOR U12755 ( .A(n13165), .B(n13166), .Z(n9521) );
  AND U12756 ( .A(n828), .B(n13167), .Z(n13166) );
  XOR U12757 ( .A(n13168), .B(n13165), .Z(n13167) );
  XOR U12758 ( .A(n13169), .B(n13170), .Z(n13157) );
  AND U12759 ( .A(n13171), .B(n13172), .Z(n13170) );
  XOR U12760 ( .A(n13169), .B(n9536), .Z(n13172) );
  XOR U12761 ( .A(n13173), .B(n13174), .Z(n9536) );
  AND U12762 ( .A(n831), .B(n13175), .Z(n13174) );
  XOR U12763 ( .A(n13176), .B(n13173), .Z(n13175) );
  XNOR U12764 ( .A(n9533), .B(n13169), .Z(n13171) );
  XOR U12765 ( .A(n13177), .B(n13178), .Z(n9533) );
  AND U12766 ( .A(n828), .B(n13179), .Z(n13178) );
  XOR U12767 ( .A(n13180), .B(n13177), .Z(n13179) );
  XOR U12768 ( .A(n13181), .B(n13182), .Z(n13169) );
  AND U12769 ( .A(n13183), .B(n13184), .Z(n13182) );
  XOR U12770 ( .A(n13181), .B(n9548), .Z(n13184) );
  XOR U12771 ( .A(n13185), .B(n13186), .Z(n9548) );
  AND U12772 ( .A(n831), .B(n13187), .Z(n13186) );
  XOR U12773 ( .A(n13188), .B(n13185), .Z(n13187) );
  XNOR U12774 ( .A(n9545), .B(n13181), .Z(n13183) );
  XOR U12775 ( .A(n13189), .B(n13190), .Z(n9545) );
  AND U12776 ( .A(n828), .B(n13191), .Z(n13190) );
  XOR U12777 ( .A(n13192), .B(n13189), .Z(n13191) );
  XOR U12778 ( .A(n13193), .B(n13194), .Z(n13181) );
  AND U12779 ( .A(n13195), .B(n13196), .Z(n13194) );
  XNOR U12780 ( .A(n13197), .B(n9561), .Z(n13196) );
  XOR U12781 ( .A(n13198), .B(n13199), .Z(n9561) );
  AND U12782 ( .A(n831), .B(n13200), .Z(n13199) );
  XOR U12783 ( .A(n13198), .B(n13201), .Z(n13200) );
  XNOR U12784 ( .A(n9558), .B(n13193), .Z(n13195) );
  XOR U12785 ( .A(n13202), .B(n13203), .Z(n9558) );
  AND U12786 ( .A(n828), .B(n13204), .Z(n13203) );
  XOR U12787 ( .A(n13202), .B(n13205), .Z(n13204) );
  IV U12788 ( .A(n13197), .Z(n13193) );
  AND U12789 ( .A(n12829), .B(n12832), .Z(n13197) );
  XNOR U12790 ( .A(n13206), .B(n13207), .Z(n12832) );
  AND U12791 ( .A(n831), .B(n13208), .Z(n13207) );
  XNOR U12792 ( .A(n13209), .B(n13206), .Z(n13208) );
  XOR U12793 ( .A(n13210), .B(n13211), .Z(n831) );
  AND U12794 ( .A(n13212), .B(n13213), .Z(n13211) );
  XOR U12795 ( .A(n13210), .B(n12840), .Z(n13213) );
  XNOR U12796 ( .A(n13214), .B(n13215), .Z(n12840) );
  AND U12797 ( .A(n13216), .B(n479), .Z(n13215) );
  AND U12798 ( .A(n13214), .B(n13217), .Z(n13216) );
  XNOR U12799 ( .A(n12837), .B(n13210), .Z(n13212) );
  XOR U12800 ( .A(n13218), .B(n13219), .Z(n12837) );
  AND U12801 ( .A(n13220), .B(n477), .Z(n13219) );
  NOR U12802 ( .A(n13218), .B(n13221), .Z(n13220) );
  XOR U12803 ( .A(n13222), .B(n13223), .Z(n13210) );
  AND U12804 ( .A(n13224), .B(n13225), .Z(n13223) );
  XOR U12805 ( .A(n13222), .B(n12852), .Z(n13225) );
  XOR U12806 ( .A(n13226), .B(n13227), .Z(n12852) );
  AND U12807 ( .A(n479), .B(n13228), .Z(n13227) );
  XOR U12808 ( .A(n13229), .B(n13226), .Z(n13228) );
  XNOR U12809 ( .A(n12849), .B(n13222), .Z(n13224) );
  XOR U12810 ( .A(n13230), .B(n13231), .Z(n12849) );
  AND U12811 ( .A(n477), .B(n13232), .Z(n13231) );
  XOR U12812 ( .A(n13233), .B(n13230), .Z(n13232) );
  XOR U12813 ( .A(n13234), .B(n13235), .Z(n13222) );
  AND U12814 ( .A(n13236), .B(n13237), .Z(n13235) );
  XOR U12815 ( .A(n13234), .B(n12864), .Z(n13237) );
  XOR U12816 ( .A(n13238), .B(n13239), .Z(n12864) );
  AND U12817 ( .A(n479), .B(n13240), .Z(n13239) );
  XOR U12818 ( .A(n13241), .B(n13238), .Z(n13240) );
  XNOR U12819 ( .A(n12861), .B(n13234), .Z(n13236) );
  XOR U12820 ( .A(n13242), .B(n13243), .Z(n12861) );
  AND U12821 ( .A(n477), .B(n13244), .Z(n13243) );
  XOR U12822 ( .A(n13245), .B(n13242), .Z(n13244) );
  XOR U12823 ( .A(n13246), .B(n13247), .Z(n13234) );
  AND U12824 ( .A(n13248), .B(n13249), .Z(n13247) );
  XOR U12825 ( .A(n13246), .B(n12876), .Z(n13249) );
  XOR U12826 ( .A(n13250), .B(n13251), .Z(n12876) );
  AND U12827 ( .A(n479), .B(n13252), .Z(n13251) );
  XOR U12828 ( .A(n13253), .B(n13250), .Z(n13252) );
  XNOR U12829 ( .A(n12873), .B(n13246), .Z(n13248) );
  XOR U12830 ( .A(n13254), .B(n13255), .Z(n12873) );
  AND U12831 ( .A(n477), .B(n13256), .Z(n13255) );
  XOR U12832 ( .A(n13257), .B(n13254), .Z(n13256) );
  XOR U12833 ( .A(n13258), .B(n13259), .Z(n13246) );
  AND U12834 ( .A(n13260), .B(n13261), .Z(n13259) );
  XOR U12835 ( .A(n13258), .B(n12888), .Z(n13261) );
  XOR U12836 ( .A(n13262), .B(n13263), .Z(n12888) );
  AND U12837 ( .A(n479), .B(n13264), .Z(n13263) );
  XOR U12838 ( .A(n13265), .B(n13262), .Z(n13264) );
  XNOR U12839 ( .A(n12885), .B(n13258), .Z(n13260) );
  XOR U12840 ( .A(n13266), .B(n13267), .Z(n12885) );
  AND U12841 ( .A(n477), .B(n13268), .Z(n13267) );
  XOR U12842 ( .A(n13269), .B(n13266), .Z(n13268) );
  XOR U12843 ( .A(n13270), .B(n13271), .Z(n13258) );
  AND U12844 ( .A(n13272), .B(n13273), .Z(n13271) );
  XOR U12845 ( .A(n13270), .B(n12900), .Z(n13273) );
  XOR U12846 ( .A(n13274), .B(n13275), .Z(n12900) );
  AND U12847 ( .A(n479), .B(n13276), .Z(n13275) );
  XOR U12848 ( .A(n13277), .B(n13274), .Z(n13276) );
  XNOR U12849 ( .A(n12897), .B(n13270), .Z(n13272) );
  XOR U12850 ( .A(n13278), .B(n13279), .Z(n12897) );
  AND U12851 ( .A(n477), .B(n13280), .Z(n13279) );
  XOR U12852 ( .A(n13281), .B(n13278), .Z(n13280) );
  XOR U12853 ( .A(n13282), .B(n13283), .Z(n13270) );
  AND U12854 ( .A(n13284), .B(n13285), .Z(n13283) );
  XOR U12855 ( .A(n13282), .B(n12912), .Z(n13285) );
  XOR U12856 ( .A(n13286), .B(n13287), .Z(n12912) );
  AND U12857 ( .A(n479), .B(n13288), .Z(n13287) );
  XOR U12858 ( .A(n13289), .B(n13286), .Z(n13288) );
  XNOR U12859 ( .A(n12909), .B(n13282), .Z(n13284) );
  XOR U12860 ( .A(n13290), .B(n13291), .Z(n12909) );
  AND U12861 ( .A(n477), .B(n13292), .Z(n13291) );
  XOR U12862 ( .A(n13293), .B(n13290), .Z(n13292) );
  XOR U12863 ( .A(n13294), .B(n13295), .Z(n13282) );
  AND U12864 ( .A(n13296), .B(n13297), .Z(n13295) );
  XOR U12865 ( .A(n13294), .B(n12924), .Z(n13297) );
  XOR U12866 ( .A(n13298), .B(n13299), .Z(n12924) );
  AND U12867 ( .A(n479), .B(n13300), .Z(n13299) );
  XOR U12868 ( .A(n13301), .B(n13298), .Z(n13300) );
  XNOR U12869 ( .A(n12921), .B(n13294), .Z(n13296) );
  XOR U12870 ( .A(n13302), .B(n13303), .Z(n12921) );
  AND U12871 ( .A(n477), .B(n13304), .Z(n13303) );
  XOR U12872 ( .A(n13305), .B(n13302), .Z(n13304) );
  XOR U12873 ( .A(n13306), .B(n13307), .Z(n13294) );
  AND U12874 ( .A(n13308), .B(n13309), .Z(n13307) );
  XOR U12875 ( .A(n13306), .B(n12936), .Z(n13309) );
  XOR U12876 ( .A(n13310), .B(n13311), .Z(n12936) );
  AND U12877 ( .A(n479), .B(n13312), .Z(n13311) );
  XOR U12878 ( .A(n13313), .B(n13310), .Z(n13312) );
  XNOR U12879 ( .A(n12933), .B(n13306), .Z(n13308) );
  XOR U12880 ( .A(n13314), .B(n13315), .Z(n12933) );
  AND U12881 ( .A(n477), .B(n13316), .Z(n13315) );
  XOR U12882 ( .A(n13317), .B(n13314), .Z(n13316) );
  XOR U12883 ( .A(n13318), .B(n13319), .Z(n13306) );
  AND U12884 ( .A(n13320), .B(n13321), .Z(n13319) );
  XOR U12885 ( .A(n13318), .B(n12948), .Z(n13321) );
  XOR U12886 ( .A(n13322), .B(n13323), .Z(n12948) );
  AND U12887 ( .A(n479), .B(n13324), .Z(n13323) );
  XOR U12888 ( .A(n13325), .B(n13322), .Z(n13324) );
  XNOR U12889 ( .A(n12945), .B(n13318), .Z(n13320) );
  XOR U12890 ( .A(n13326), .B(n13327), .Z(n12945) );
  AND U12891 ( .A(n477), .B(n13328), .Z(n13327) );
  XOR U12892 ( .A(n13329), .B(n13326), .Z(n13328) );
  XOR U12893 ( .A(n13330), .B(n13331), .Z(n13318) );
  AND U12894 ( .A(n13332), .B(n13333), .Z(n13331) );
  XOR U12895 ( .A(n13330), .B(n12960), .Z(n13333) );
  XOR U12896 ( .A(n13334), .B(n13335), .Z(n12960) );
  AND U12897 ( .A(n479), .B(n13336), .Z(n13335) );
  XOR U12898 ( .A(n13337), .B(n13334), .Z(n13336) );
  XNOR U12899 ( .A(n12957), .B(n13330), .Z(n13332) );
  XOR U12900 ( .A(n13338), .B(n13339), .Z(n12957) );
  AND U12901 ( .A(n477), .B(n13340), .Z(n13339) );
  XOR U12902 ( .A(n13341), .B(n13338), .Z(n13340) );
  XOR U12903 ( .A(n13342), .B(n13343), .Z(n13330) );
  AND U12904 ( .A(n13344), .B(n13345), .Z(n13343) );
  XOR U12905 ( .A(n13342), .B(n12972), .Z(n13345) );
  XOR U12906 ( .A(n13346), .B(n13347), .Z(n12972) );
  AND U12907 ( .A(n479), .B(n13348), .Z(n13347) );
  XOR U12908 ( .A(n13349), .B(n13346), .Z(n13348) );
  XNOR U12909 ( .A(n12969), .B(n13342), .Z(n13344) );
  XOR U12910 ( .A(n13350), .B(n13351), .Z(n12969) );
  AND U12911 ( .A(n477), .B(n13352), .Z(n13351) );
  XOR U12912 ( .A(n13353), .B(n13350), .Z(n13352) );
  XOR U12913 ( .A(n13354), .B(n13355), .Z(n13342) );
  AND U12914 ( .A(n13356), .B(n13357), .Z(n13355) );
  XOR U12915 ( .A(n13354), .B(n12984), .Z(n13357) );
  XOR U12916 ( .A(n13358), .B(n13359), .Z(n12984) );
  AND U12917 ( .A(n479), .B(n13360), .Z(n13359) );
  XOR U12918 ( .A(n13361), .B(n13358), .Z(n13360) );
  XNOR U12919 ( .A(n12981), .B(n13354), .Z(n13356) );
  XOR U12920 ( .A(n13362), .B(n13363), .Z(n12981) );
  AND U12921 ( .A(n477), .B(n13364), .Z(n13363) );
  XOR U12922 ( .A(n13365), .B(n13362), .Z(n13364) );
  XOR U12923 ( .A(n13366), .B(n13367), .Z(n13354) );
  AND U12924 ( .A(n13368), .B(n13369), .Z(n13367) );
  XOR U12925 ( .A(n13366), .B(n12996), .Z(n13369) );
  XOR U12926 ( .A(n13370), .B(n13371), .Z(n12996) );
  AND U12927 ( .A(n479), .B(n13372), .Z(n13371) );
  XOR U12928 ( .A(n13373), .B(n13370), .Z(n13372) );
  XNOR U12929 ( .A(n12993), .B(n13366), .Z(n13368) );
  XOR U12930 ( .A(n13374), .B(n13375), .Z(n12993) );
  AND U12931 ( .A(n477), .B(n13376), .Z(n13375) );
  XOR U12932 ( .A(n13377), .B(n13374), .Z(n13376) );
  XOR U12933 ( .A(n13378), .B(n13379), .Z(n13366) );
  AND U12934 ( .A(n13380), .B(n13381), .Z(n13379) );
  XOR U12935 ( .A(n13378), .B(n13008), .Z(n13381) );
  XOR U12936 ( .A(n13382), .B(n13383), .Z(n13008) );
  AND U12937 ( .A(n479), .B(n13384), .Z(n13383) );
  XOR U12938 ( .A(n13385), .B(n13382), .Z(n13384) );
  XNOR U12939 ( .A(n13005), .B(n13378), .Z(n13380) );
  XOR U12940 ( .A(n13386), .B(n13387), .Z(n13005) );
  AND U12941 ( .A(n477), .B(n13388), .Z(n13387) );
  XOR U12942 ( .A(n13389), .B(n13386), .Z(n13388) );
  XOR U12943 ( .A(n13390), .B(n13391), .Z(n13378) );
  AND U12944 ( .A(n13392), .B(n13393), .Z(n13391) );
  XOR U12945 ( .A(n13390), .B(n13020), .Z(n13393) );
  XOR U12946 ( .A(n13394), .B(n13395), .Z(n13020) );
  AND U12947 ( .A(n479), .B(n13396), .Z(n13395) );
  XOR U12948 ( .A(n13397), .B(n13394), .Z(n13396) );
  XNOR U12949 ( .A(n13017), .B(n13390), .Z(n13392) );
  XOR U12950 ( .A(n13398), .B(n13399), .Z(n13017) );
  AND U12951 ( .A(n477), .B(n13400), .Z(n13399) );
  XOR U12952 ( .A(n13401), .B(n13398), .Z(n13400) );
  XOR U12953 ( .A(n13402), .B(n13403), .Z(n13390) );
  AND U12954 ( .A(n13404), .B(n13405), .Z(n13403) );
  XOR U12955 ( .A(n13402), .B(n13032), .Z(n13405) );
  XOR U12956 ( .A(n13406), .B(n13407), .Z(n13032) );
  AND U12957 ( .A(n479), .B(n13408), .Z(n13407) );
  XOR U12958 ( .A(n13409), .B(n13406), .Z(n13408) );
  XNOR U12959 ( .A(n13029), .B(n13402), .Z(n13404) );
  XOR U12960 ( .A(n13410), .B(n13411), .Z(n13029) );
  AND U12961 ( .A(n477), .B(n13412), .Z(n13411) );
  XOR U12962 ( .A(n13413), .B(n13410), .Z(n13412) );
  XOR U12963 ( .A(n13414), .B(n13415), .Z(n13402) );
  AND U12964 ( .A(n13416), .B(n13417), .Z(n13415) );
  XOR U12965 ( .A(n13414), .B(n13044), .Z(n13417) );
  XOR U12966 ( .A(n13418), .B(n13419), .Z(n13044) );
  AND U12967 ( .A(n479), .B(n13420), .Z(n13419) );
  XOR U12968 ( .A(n13421), .B(n13418), .Z(n13420) );
  XNOR U12969 ( .A(n13041), .B(n13414), .Z(n13416) );
  XOR U12970 ( .A(n13422), .B(n13423), .Z(n13041) );
  AND U12971 ( .A(n477), .B(n13424), .Z(n13423) );
  XOR U12972 ( .A(n13425), .B(n13422), .Z(n13424) );
  XOR U12973 ( .A(n13426), .B(n13427), .Z(n13414) );
  AND U12974 ( .A(n13428), .B(n13429), .Z(n13427) );
  XOR U12975 ( .A(n13426), .B(n13056), .Z(n13429) );
  XOR U12976 ( .A(n13430), .B(n13431), .Z(n13056) );
  AND U12977 ( .A(n479), .B(n13432), .Z(n13431) );
  XOR U12978 ( .A(n13433), .B(n13430), .Z(n13432) );
  XNOR U12979 ( .A(n13053), .B(n13426), .Z(n13428) );
  XOR U12980 ( .A(n13434), .B(n13435), .Z(n13053) );
  AND U12981 ( .A(n477), .B(n13436), .Z(n13435) );
  XOR U12982 ( .A(n13437), .B(n13434), .Z(n13436) );
  XOR U12983 ( .A(n13438), .B(n13439), .Z(n13426) );
  AND U12984 ( .A(n13440), .B(n13441), .Z(n13439) );
  XOR U12985 ( .A(n13438), .B(n13068), .Z(n13441) );
  XOR U12986 ( .A(n13442), .B(n13443), .Z(n13068) );
  AND U12987 ( .A(n479), .B(n13444), .Z(n13443) );
  XOR U12988 ( .A(n13445), .B(n13442), .Z(n13444) );
  XNOR U12989 ( .A(n13065), .B(n13438), .Z(n13440) );
  XOR U12990 ( .A(n13446), .B(n13447), .Z(n13065) );
  AND U12991 ( .A(n477), .B(n13448), .Z(n13447) );
  XOR U12992 ( .A(n13449), .B(n13446), .Z(n13448) );
  XOR U12993 ( .A(n13450), .B(n13451), .Z(n13438) );
  AND U12994 ( .A(n13452), .B(n13453), .Z(n13451) );
  XOR U12995 ( .A(n13450), .B(n13080), .Z(n13453) );
  XOR U12996 ( .A(n13454), .B(n13455), .Z(n13080) );
  AND U12997 ( .A(n479), .B(n13456), .Z(n13455) );
  XOR U12998 ( .A(n13457), .B(n13454), .Z(n13456) );
  XNOR U12999 ( .A(n13077), .B(n13450), .Z(n13452) );
  XOR U13000 ( .A(n13458), .B(n13459), .Z(n13077) );
  AND U13001 ( .A(n477), .B(n13460), .Z(n13459) );
  XOR U13002 ( .A(n13461), .B(n13458), .Z(n13460) );
  XOR U13003 ( .A(n13462), .B(n13463), .Z(n13450) );
  AND U13004 ( .A(n13464), .B(n13465), .Z(n13463) );
  XOR U13005 ( .A(n13462), .B(n13092), .Z(n13465) );
  XOR U13006 ( .A(n13466), .B(n13467), .Z(n13092) );
  AND U13007 ( .A(n479), .B(n13468), .Z(n13467) );
  XOR U13008 ( .A(n13469), .B(n13466), .Z(n13468) );
  XNOR U13009 ( .A(n13089), .B(n13462), .Z(n13464) );
  XOR U13010 ( .A(n13470), .B(n13471), .Z(n13089) );
  AND U13011 ( .A(n477), .B(n13472), .Z(n13471) );
  XOR U13012 ( .A(n13473), .B(n13470), .Z(n13472) );
  XOR U13013 ( .A(n13474), .B(n13475), .Z(n13462) );
  AND U13014 ( .A(n13476), .B(n13477), .Z(n13475) );
  XOR U13015 ( .A(n13474), .B(n13104), .Z(n13477) );
  XOR U13016 ( .A(n13478), .B(n13479), .Z(n13104) );
  AND U13017 ( .A(n479), .B(n13480), .Z(n13479) );
  XOR U13018 ( .A(n13481), .B(n13478), .Z(n13480) );
  XNOR U13019 ( .A(n13101), .B(n13474), .Z(n13476) );
  XOR U13020 ( .A(n13482), .B(n13483), .Z(n13101) );
  AND U13021 ( .A(n477), .B(n13484), .Z(n13483) );
  XOR U13022 ( .A(n13485), .B(n13482), .Z(n13484) );
  XOR U13023 ( .A(n13486), .B(n13487), .Z(n13474) );
  AND U13024 ( .A(n13488), .B(n13489), .Z(n13487) );
  XOR U13025 ( .A(n13486), .B(n13116), .Z(n13489) );
  XOR U13026 ( .A(n13490), .B(n13491), .Z(n13116) );
  AND U13027 ( .A(n479), .B(n13492), .Z(n13491) );
  XOR U13028 ( .A(n13493), .B(n13490), .Z(n13492) );
  XNOR U13029 ( .A(n13113), .B(n13486), .Z(n13488) );
  XOR U13030 ( .A(n13494), .B(n13495), .Z(n13113) );
  AND U13031 ( .A(n477), .B(n13496), .Z(n13495) );
  XOR U13032 ( .A(n13497), .B(n13494), .Z(n13496) );
  XOR U13033 ( .A(n13498), .B(n13499), .Z(n13486) );
  AND U13034 ( .A(n13500), .B(n13501), .Z(n13499) );
  XOR U13035 ( .A(n13498), .B(n13128), .Z(n13501) );
  XOR U13036 ( .A(n13502), .B(n13503), .Z(n13128) );
  AND U13037 ( .A(n479), .B(n13504), .Z(n13503) );
  XOR U13038 ( .A(n13505), .B(n13502), .Z(n13504) );
  XNOR U13039 ( .A(n13125), .B(n13498), .Z(n13500) );
  XOR U13040 ( .A(n13506), .B(n13507), .Z(n13125) );
  AND U13041 ( .A(n477), .B(n13508), .Z(n13507) );
  XOR U13042 ( .A(n13509), .B(n13506), .Z(n13508) );
  XOR U13043 ( .A(n13510), .B(n13511), .Z(n13498) );
  AND U13044 ( .A(n13512), .B(n13513), .Z(n13511) );
  XOR U13045 ( .A(n13510), .B(n13140), .Z(n13513) );
  XOR U13046 ( .A(n13514), .B(n13515), .Z(n13140) );
  AND U13047 ( .A(n479), .B(n13516), .Z(n13515) );
  XOR U13048 ( .A(n13517), .B(n13514), .Z(n13516) );
  XNOR U13049 ( .A(n13137), .B(n13510), .Z(n13512) );
  XOR U13050 ( .A(n13518), .B(n13519), .Z(n13137) );
  AND U13051 ( .A(n477), .B(n13520), .Z(n13519) );
  XOR U13052 ( .A(n13521), .B(n13518), .Z(n13520) );
  XOR U13053 ( .A(n13522), .B(n13523), .Z(n13510) );
  AND U13054 ( .A(n13524), .B(n13525), .Z(n13523) );
  XOR U13055 ( .A(n13522), .B(n13152), .Z(n13525) );
  XOR U13056 ( .A(n13526), .B(n13527), .Z(n13152) );
  AND U13057 ( .A(n479), .B(n13528), .Z(n13527) );
  XOR U13058 ( .A(n13529), .B(n13526), .Z(n13528) );
  XNOR U13059 ( .A(n13149), .B(n13522), .Z(n13524) );
  XOR U13060 ( .A(n13530), .B(n13531), .Z(n13149) );
  AND U13061 ( .A(n477), .B(n13532), .Z(n13531) );
  XOR U13062 ( .A(n13533), .B(n13530), .Z(n13532) );
  XOR U13063 ( .A(n13534), .B(n13535), .Z(n13522) );
  AND U13064 ( .A(n13536), .B(n13537), .Z(n13535) );
  XOR U13065 ( .A(n13534), .B(n13164), .Z(n13537) );
  XOR U13066 ( .A(n13538), .B(n13539), .Z(n13164) );
  AND U13067 ( .A(n479), .B(n13540), .Z(n13539) );
  XOR U13068 ( .A(n13541), .B(n13538), .Z(n13540) );
  XNOR U13069 ( .A(n13161), .B(n13534), .Z(n13536) );
  XOR U13070 ( .A(n13542), .B(n13543), .Z(n13161) );
  AND U13071 ( .A(n477), .B(n13544), .Z(n13543) );
  XOR U13072 ( .A(n13545), .B(n13542), .Z(n13544) );
  XOR U13073 ( .A(n13546), .B(n13547), .Z(n13534) );
  AND U13074 ( .A(n13548), .B(n13549), .Z(n13547) );
  XOR U13075 ( .A(n13546), .B(n13176), .Z(n13549) );
  XOR U13076 ( .A(n13550), .B(n13551), .Z(n13176) );
  AND U13077 ( .A(n479), .B(n13552), .Z(n13551) );
  XOR U13078 ( .A(n13553), .B(n13550), .Z(n13552) );
  XNOR U13079 ( .A(n13173), .B(n13546), .Z(n13548) );
  XOR U13080 ( .A(n13554), .B(n13555), .Z(n13173) );
  AND U13081 ( .A(n477), .B(n13556), .Z(n13555) );
  XOR U13082 ( .A(n13557), .B(n13554), .Z(n13556) );
  XOR U13083 ( .A(n13558), .B(n13559), .Z(n13546) );
  AND U13084 ( .A(n13560), .B(n13561), .Z(n13559) );
  XOR U13085 ( .A(n13558), .B(n13188), .Z(n13561) );
  XOR U13086 ( .A(n13562), .B(n13563), .Z(n13188) );
  AND U13087 ( .A(n479), .B(n13564), .Z(n13563) );
  XOR U13088 ( .A(n13565), .B(n13562), .Z(n13564) );
  XNOR U13089 ( .A(n13185), .B(n13558), .Z(n13560) );
  XOR U13090 ( .A(n13566), .B(n13567), .Z(n13185) );
  AND U13091 ( .A(n477), .B(n13568), .Z(n13567) );
  XOR U13092 ( .A(n13569), .B(n13566), .Z(n13568) );
  XOR U13093 ( .A(n13570), .B(n13571), .Z(n13558) );
  AND U13094 ( .A(n13572), .B(n13573), .Z(n13571) );
  XNOR U13095 ( .A(n13574), .B(n13201), .Z(n13573) );
  XOR U13096 ( .A(n13575), .B(n13576), .Z(n13201) );
  AND U13097 ( .A(n479), .B(n13577), .Z(n13576) );
  XOR U13098 ( .A(n13575), .B(n13578), .Z(n13577) );
  XNOR U13099 ( .A(n13198), .B(n13570), .Z(n13572) );
  XOR U13100 ( .A(n13579), .B(n13580), .Z(n13198) );
  AND U13101 ( .A(n477), .B(n13581), .Z(n13580) );
  XOR U13102 ( .A(n13579), .B(n13582), .Z(n13581) );
  IV U13103 ( .A(n13574), .Z(n13570) );
  AND U13104 ( .A(n13206), .B(n13209), .Z(n13574) );
  XNOR U13105 ( .A(n13583), .B(n13584), .Z(n13209) );
  AND U13106 ( .A(n479), .B(n13585), .Z(n13584) );
  XNOR U13107 ( .A(n13586), .B(n13583), .Z(n13585) );
  XOR U13108 ( .A(n13587), .B(n13588), .Z(n479) );
  AND U13109 ( .A(n13589), .B(n13590), .Z(n13588) );
  XOR U13110 ( .A(n13217), .B(n13587), .Z(n13590) );
  IV U13111 ( .A(n13591), .Z(n13217) );
  AND U13112 ( .A(p_input[6655]), .B(p_input[6623]), .Z(n13591) );
  XOR U13113 ( .A(n13587), .B(n13214), .Z(n13589) );
  AND U13114 ( .A(p_input[6559]), .B(p_input[6591]), .Z(n13214) );
  XOR U13115 ( .A(n13592), .B(n13593), .Z(n13587) );
  AND U13116 ( .A(n13594), .B(n13595), .Z(n13593) );
  XOR U13117 ( .A(n13592), .B(n13229), .Z(n13595) );
  XNOR U13118 ( .A(p_input[6622]), .B(n13596), .Z(n13229) );
  AND U13119 ( .A(n275), .B(n13597), .Z(n13596) );
  XOR U13120 ( .A(p_input[6654]), .B(p_input[6622]), .Z(n13597) );
  XNOR U13121 ( .A(n13226), .B(n13592), .Z(n13594) );
  XOR U13122 ( .A(n13598), .B(n13599), .Z(n13226) );
  AND U13123 ( .A(n273), .B(n13600), .Z(n13599) );
  XOR U13124 ( .A(p_input[6590]), .B(p_input[6558]), .Z(n13600) );
  XOR U13125 ( .A(n13601), .B(n13602), .Z(n13592) );
  AND U13126 ( .A(n13603), .B(n13604), .Z(n13602) );
  XOR U13127 ( .A(n13601), .B(n13241), .Z(n13604) );
  XNOR U13128 ( .A(p_input[6621]), .B(n13605), .Z(n13241) );
  AND U13129 ( .A(n275), .B(n13606), .Z(n13605) );
  XOR U13130 ( .A(p_input[6653]), .B(p_input[6621]), .Z(n13606) );
  XNOR U13131 ( .A(n13238), .B(n13601), .Z(n13603) );
  XOR U13132 ( .A(n13607), .B(n13608), .Z(n13238) );
  AND U13133 ( .A(n273), .B(n13609), .Z(n13608) );
  XOR U13134 ( .A(p_input[6589]), .B(p_input[6557]), .Z(n13609) );
  XOR U13135 ( .A(n13610), .B(n13611), .Z(n13601) );
  AND U13136 ( .A(n13612), .B(n13613), .Z(n13611) );
  XOR U13137 ( .A(n13610), .B(n13253), .Z(n13613) );
  XNOR U13138 ( .A(p_input[6620]), .B(n13614), .Z(n13253) );
  AND U13139 ( .A(n275), .B(n13615), .Z(n13614) );
  XOR U13140 ( .A(p_input[6652]), .B(p_input[6620]), .Z(n13615) );
  XNOR U13141 ( .A(n13250), .B(n13610), .Z(n13612) );
  XOR U13142 ( .A(n13616), .B(n13617), .Z(n13250) );
  AND U13143 ( .A(n273), .B(n13618), .Z(n13617) );
  XOR U13144 ( .A(p_input[6588]), .B(p_input[6556]), .Z(n13618) );
  XOR U13145 ( .A(n13619), .B(n13620), .Z(n13610) );
  AND U13146 ( .A(n13621), .B(n13622), .Z(n13620) );
  XOR U13147 ( .A(n13619), .B(n13265), .Z(n13622) );
  XNOR U13148 ( .A(p_input[6619]), .B(n13623), .Z(n13265) );
  AND U13149 ( .A(n275), .B(n13624), .Z(n13623) );
  XOR U13150 ( .A(p_input[6651]), .B(p_input[6619]), .Z(n13624) );
  XNOR U13151 ( .A(n13262), .B(n13619), .Z(n13621) );
  XOR U13152 ( .A(n13625), .B(n13626), .Z(n13262) );
  AND U13153 ( .A(n273), .B(n13627), .Z(n13626) );
  XOR U13154 ( .A(p_input[6587]), .B(p_input[6555]), .Z(n13627) );
  XOR U13155 ( .A(n13628), .B(n13629), .Z(n13619) );
  AND U13156 ( .A(n13630), .B(n13631), .Z(n13629) );
  XOR U13157 ( .A(n13628), .B(n13277), .Z(n13631) );
  XNOR U13158 ( .A(p_input[6618]), .B(n13632), .Z(n13277) );
  AND U13159 ( .A(n275), .B(n13633), .Z(n13632) );
  XOR U13160 ( .A(p_input[6650]), .B(p_input[6618]), .Z(n13633) );
  XNOR U13161 ( .A(n13274), .B(n13628), .Z(n13630) );
  XOR U13162 ( .A(n13634), .B(n13635), .Z(n13274) );
  AND U13163 ( .A(n273), .B(n13636), .Z(n13635) );
  XOR U13164 ( .A(p_input[6586]), .B(p_input[6554]), .Z(n13636) );
  XOR U13165 ( .A(n13637), .B(n13638), .Z(n13628) );
  AND U13166 ( .A(n13639), .B(n13640), .Z(n13638) );
  XOR U13167 ( .A(n13637), .B(n13289), .Z(n13640) );
  XNOR U13168 ( .A(p_input[6617]), .B(n13641), .Z(n13289) );
  AND U13169 ( .A(n275), .B(n13642), .Z(n13641) );
  XOR U13170 ( .A(p_input[6649]), .B(p_input[6617]), .Z(n13642) );
  XNOR U13171 ( .A(n13286), .B(n13637), .Z(n13639) );
  XOR U13172 ( .A(n13643), .B(n13644), .Z(n13286) );
  AND U13173 ( .A(n273), .B(n13645), .Z(n13644) );
  XOR U13174 ( .A(p_input[6585]), .B(p_input[6553]), .Z(n13645) );
  XOR U13175 ( .A(n13646), .B(n13647), .Z(n13637) );
  AND U13176 ( .A(n13648), .B(n13649), .Z(n13647) );
  XOR U13177 ( .A(n13646), .B(n13301), .Z(n13649) );
  XNOR U13178 ( .A(p_input[6616]), .B(n13650), .Z(n13301) );
  AND U13179 ( .A(n275), .B(n13651), .Z(n13650) );
  XOR U13180 ( .A(p_input[6648]), .B(p_input[6616]), .Z(n13651) );
  XNOR U13181 ( .A(n13298), .B(n13646), .Z(n13648) );
  XOR U13182 ( .A(n13652), .B(n13653), .Z(n13298) );
  AND U13183 ( .A(n273), .B(n13654), .Z(n13653) );
  XOR U13184 ( .A(p_input[6584]), .B(p_input[6552]), .Z(n13654) );
  XOR U13185 ( .A(n13655), .B(n13656), .Z(n13646) );
  AND U13186 ( .A(n13657), .B(n13658), .Z(n13656) );
  XOR U13187 ( .A(n13655), .B(n13313), .Z(n13658) );
  XNOR U13188 ( .A(p_input[6615]), .B(n13659), .Z(n13313) );
  AND U13189 ( .A(n275), .B(n13660), .Z(n13659) );
  XOR U13190 ( .A(p_input[6647]), .B(p_input[6615]), .Z(n13660) );
  XNOR U13191 ( .A(n13310), .B(n13655), .Z(n13657) );
  XOR U13192 ( .A(n13661), .B(n13662), .Z(n13310) );
  AND U13193 ( .A(n273), .B(n13663), .Z(n13662) );
  XOR U13194 ( .A(p_input[6583]), .B(p_input[6551]), .Z(n13663) );
  XOR U13195 ( .A(n13664), .B(n13665), .Z(n13655) );
  AND U13196 ( .A(n13666), .B(n13667), .Z(n13665) );
  XOR U13197 ( .A(n13664), .B(n13325), .Z(n13667) );
  XNOR U13198 ( .A(p_input[6614]), .B(n13668), .Z(n13325) );
  AND U13199 ( .A(n275), .B(n13669), .Z(n13668) );
  XOR U13200 ( .A(p_input[6646]), .B(p_input[6614]), .Z(n13669) );
  XNOR U13201 ( .A(n13322), .B(n13664), .Z(n13666) );
  XOR U13202 ( .A(n13670), .B(n13671), .Z(n13322) );
  AND U13203 ( .A(n273), .B(n13672), .Z(n13671) );
  XOR U13204 ( .A(p_input[6582]), .B(p_input[6550]), .Z(n13672) );
  XOR U13205 ( .A(n13673), .B(n13674), .Z(n13664) );
  AND U13206 ( .A(n13675), .B(n13676), .Z(n13674) );
  XOR U13207 ( .A(n13673), .B(n13337), .Z(n13676) );
  XNOR U13208 ( .A(p_input[6613]), .B(n13677), .Z(n13337) );
  AND U13209 ( .A(n275), .B(n13678), .Z(n13677) );
  XOR U13210 ( .A(p_input[6645]), .B(p_input[6613]), .Z(n13678) );
  XNOR U13211 ( .A(n13334), .B(n13673), .Z(n13675) );
  XOR U13212 ( .A(n13679), .B(n13680), .Z(n13334) );
  AND U13213 ( .A(n273), .B(n13681), .Z(n13680) );
  XOR U13214 ( .A(p_input[6581]), .B(p_input[6549]), .Z(n13681) );
  XOR U13215 ( .A(n13682), .B(n13683), .Z(n13673) );
  AND U13216 ( .A(n13684), .B(n13685), .Z(n13683) );
  XOR U13217 ( .A(n13682), .B(n13349), .Z(n13685) );
  XNOR U13218 ( .A(p_input[6612]), .B(n13686), .Z(n13349) );
  AND U13219 ( .A(n275), .B(n13687), .Z(n13686) );
  XOR U13220 ( .A(p_input[6644]), .B(p_input[6612]), .Z(n13687) );
  XNOR U13221 ( .A(n13346), .B(n13682), .Z(n13684) );
  XOR U13222 ( .A(n13688), .B(n13689), .Z(n13346) );
  AND U13223 ( .A(n273), .B(n13690), .Z(n13689) );
  XOR U13224 ( .A(p_input[6580]), .B(p_input[6548]), .Z(n13690) );
  XOR U13225 ( .A(n13691), .B(n13692), .Z(n13682) );
  AND U13226 ( .A(n13693), .B(n13694), .Z(n13692) );
  XOR U13227 ( .A(n13691), .B(n13361), .Z(n13694) );
  XNOR U13228 ( .A(p_input[6611]), .B(n13695), .Z(n13361) );
  AND U13229 ( .A(n275), .B(n13696), .Z(n13695) );
  XOR U13230 ( .A(p_input[6643]), .B(p_input[6611]), .Z(n13696) );
  XNOR U13231 ( .A(n13358), .B(n13691), .Z(n13693) );
  XOR U13232 ( .A(n13697), .B(n13698), .Z(n13358) );
  AND U13233 ( .A(n273), .B(n13699), .Z(n13698) );
  XOR U13234 ( .A(p_input[6579]), .B(p_input[6547]), .Z(n13699) );
  XOR U13235 ( .A(n13700), .B(n13701), .Z(n13691) );
  AND U13236 ( .A(n13702), .B(n13703), .Z(n13701) );
  XOR U13237 ( .A(n13700), .B(n13373), .Z(n13703) );
  XNOR U13238 ( .A(p_input[6610]), .B(n13704), .Z(n13373) );
  AND U13239 ( .A(n275), .B(n13705), .Z(n13704) );
  XOR U13240 ( .A(p_input[6642]), .B(p_input[6610]), .Z(n13705) );
  XNOR U13241 ( .A(n13370), .B(n13700), .Z(n13702) );
  XOR U13242 ( .A(n13706), .B(n13707), .Z(n13370) );
  AND U13243 ( .A(n273), .B(n13708), .Z(n13707) );
  XOR U13244 ( .A(p_input[6578]), .B(p_input[6546]), .Z(n13708) );
  XOR U13245 ( .A(n13709), .B(n13710), .Z(n13700) );
  AND U13246 ( .A(n13711), .B(n13712), .Z(n13710) );
  XOR U13247 ( .A(n13709), .B(n13385), .Z(n13712) );
  XNOR U13248 ( .A(p_input[6609]), .B(n13713), .Z(n13385) );
  AND U13249 ( .A(n275), .B(n13714), .Z(n13713) );
  XOR U13250 ( .A(p_input[6641]), .B(p_input[6609]), .Z(n13714) );
  XNOR U13251 ( .A(n13382), .B(n13709), .Z(n13711) );
  XOR U13252 ( .A(n13715), .B(n13716), .Z(n13382) );
  AND U13253 ( .A(n273), .B(n13717), .Z(n13716) );
  XOR U13254 ( .A(p_input[6577]), .B(p_input[6545]), .Z(n13717) );
  XOR U13255 ( .A(n13718), .B(n13719), .Z(n13709) );
  AND U13256 ( .A(n13720), .B(n13721), .Z(n13719) );
  XOR U13257 ( .A(n13718), .B(n13397), .Z(n13721) );
  XNOR U13258 ( .A(p_input[6608]), .B(n13722), .Z(n13397) );
  AND U13259 ( .A(n275), .B(n13723), .Z(n13722) );
  XOR U13260 ( .A(p_input[6640]), .B(p_input[6608]), .Z(n13723) );
  XNOR U13261 ( .A(n13394), .B(n13718), .Z(n13720) );
  XOR U13262 ( .A(n13724), .B(n13725), .Z(n13394) );
  AND U13263 ( .A(n273), .B(n13726), .Z(n13725) );
  XOR U13264 ( .A(p_input[6576]), .B(p_input[6544]), .Z(n13726) );
  XOR U13265 ( .A(n13727), .B(n13728), .Z(n13718) );
  AND U13266 ( .A(n13729), .B(n13730), .Z(n13728) );
  XOR U13267 ( .A(n13727), .B(n13409), .Z(n13730) );
  XNOR U13268 ( .A(p_input[6607]), .B(n13731), .Z(n13409) );
  AND U13269 ( .A(n275), .B(n13732), .Z(n13731) );
  XOR U13270 ( .A(p_input[6639]), .B(p_input[6607]), .Z(n13732) );
  XNOR U13271 ( .A(n13406), .B(n13727), .Z(n13729) );
  XOR U13272 ( .A(n13733), .B(n13734), .Z(n13406) );
  AND U13273 ( .A(n273), .B(n13735), .Z(n13734) );
  XOR U13274 ( .A(p_input[6575]), .B(p_input[6543]), .Z(n13735) );
  XOR U13275 ( .A(n13736), .B(n13737), .Z(n13727) );
  AND U13276 ( .A(n13738), .B(n13739), .Z(n13737) );
  XOR U13277 ( .A(n13736), .B(n13421), .Z(n13739) );
  XNOR U13278 ( .A(p_input[6606]), .B(n13740), .Z(n13421) );
  AND U13279 ( .A(n275), .B(n13741), .Z(n13740) );
  XOR U13280 ( .A(p_input[6638]), .B(p_input[6606]), .Z(n13741) );
  XNOR U13281 ( .A(n13418), .B(n13736), .Z(n13738) );
  XOR U13282 ( .A(n13742), .B(n13743), .Z(n13418) );
  AND U13283 ( .A(n273), .B(n13744), .Z(n13743) );
  XOR U13284 ( .A(p_input[6574]), .B(p_input[6542]), .Z(n13744) );
  XOR U13285 ( .A(n13745), .B(n13746), .Z(n13736) );
  AND U13286 ( .A(n13747), .B(n13748), .Z(n13746) );
  XOR U13287 ( .A(n13745), .B(n13433), .Z(n13748) );
  XNOR U13288 ( .A(p_input[6605]), .B(n13749), .Z(n13433) );
  AND U13289 ( .A(n275), .B(n13750), .Z(n13749) );
  XOR U13290 ( .A(p_input[6637]), .B(p_input[6605]), .Z(n13750) );
  XNOR U13291 ( .A(n13430), .B(n13745), .Z(n13747) );
  XOR U13292 ( .A(n13751), .B(n13752), .Z(n13430) );
  AND U13293 ( .A(n273), .B(n13753), .Z(n13752) );
  XOR U13294 ( .A(p_input[6573]), .B(p_input[6541]), .Z(n13753) );
  XOR U13295 ( .A(n13754), .B(n13755), .Z(n13745) );
  AND U13296 ( .A(n13756), .B(n13757), .Z(n13755) );
  XOR U13297 ( .A(n13754), .B(n13445), .Z(n13757) );
  XNOR U13298 ( .A(p_input[6604]), .B(n13758), .Z(n13445) );
  AND U13299 ( .A(n275), .B(n13759), .Z(n13758) );
  XOR U13300 ( .A(p_input[6636]), .B(p_input[6604]), .Z(n13759) );
  XNOR U13301 ( .A(n13442), .B(n13754), .Z(n13756) );
  XOR U13302 ( .A(n13760), .B(n13761), .Z(n13442) );
  AND U13303 ( .A(n273), .B(n13762), .Z(n13761) );
  XOR U13304 ( .A(p_input[6572]), .B(p_input[6540]), .Z(n13762) );
  XOR U13305 ( .A(n13763), .B(n13764), .Z(n13754) );
  AND U13306 ( .A(n13765), .B(n13766), .Z(n13764) );
  XOR U13307 ( .A(n13763), .B(n13457), .Z(n13766) );
  XNOR U13308 ( .A(p_input[6603]), .B(n13767), .Z(n13457) );
  AND U13309 ( .A(n275), .B(n13768), .Z(n13767) );
  XOR U13310 ( .A(p_input[6635]), .B(p_input[6603]), .Z(n13768) );
  XNOR U13311 ( .A(n13454), .B(n13763), .Z(n13765) );
  XOR U13312 ( .A(n13769), .B(n13770), .Z(n13454) );
  AND U13313 ( .A(n273), .B(n13771), .Z(n13770) );
  XOR U13314 ( .A(p_input[6571]), .B(p_input[6539]), .Z(n13771) );
  XOR U13315 ( .A(n13772), .B(n13773), .Z(n13763) );
  AND U13316 ( .A(n13774), .B(n13775), .Z(n13773) );
  XOR U13317 ( .A(n13772), .B(n13469), .Z(n13775) );
  XNOR U13318 ( .A(p_input[6602]), .B(n13776), .Z(n13469) );
  AND U13319 ( .A(n275), .B(n13777), .Z(n13776) );
  XOR U13320 ( .A(p_input[6634]), .B(p_input[6602]), .Z(n13777) );
  XNOR U13321 ( .A(n13466), .B(n13772), .Z(n13774) );
  XOR U13322 ( .A(n13778), .B(n13779), .Z(n13466) );
  AND U13323 ( .A(n273), .B(n13780), .Z(n13779) );
  XOR U13324 ( .A(p_input[6570]), .B(p_input[6538]), .Z(n13780) );
  XOR U13325 ( .A(n13781), .B(n13782), .Z(n13772) );
  AND U13326 ( .A(n13783), .B(n13784), .Z(n13782) );
  XOR U13327 ( .A(n13781), .B(n13481), .Z(n13784) );
  XNOR U13328 ( .A(p_input[6601]), .B(n13785), .Z(n13481) );
  AND U13329 ( .A(n275), .B(n13786), .Z(n13785) );
  XOR U13330 ( .A(p_input[6633]), .B(p_input[6601]), .Z(n13786) );
  XNOR U13331 ( .A(n13478), .B(n13781), .Z(n13783) );
  XOR U13332 ( .A(n13787), .B(n13788), .Z(n13478) );
  AND U13333 ( .A(n273), .B(n13789), .Z(n13788) );
  XOR U13334 ( .A(p_input[6569]), .B(p_input[6537]), .Z(n13789) );
  XOR U13335 ( .A(n13790), .B(n13791), .Z(n13781) );
  AND U13336 ( .A(n13792), .B(n13793), .Z(n13791) );
  XOR U13337 ( .A(n13790), .B(n13493), .Z(n13793) );
  XNOR U13338 ( .A(p_input[6600]), .B(n13794), .Z(n13493) );
  AND U13339 ( .A(n275), .B(n13795), .Z(n13794) );
  XOR U13340 ( .A(p_input[6632]), .B(p_input[6600]), .Z(n13795) );
  XNOR U13341 ( .A(n13490), .B(n13790), .Z(n13792) );
  XOR U13342 ( .A(n13796), .B(n13797), .Z(n13490) );
  AND U13343 ( .A(n273), .B(n13798), .Z(n13797) );
  XOR U13344 ( .A(p_input[6568]), .B(p_input[6536]), .Z(n13798) );
  XOR U13345 ( .A(n13799), .B(n13800), .Z(n13790) );
  AND U13346 ( .A(n13801), .B(n13802), .Z(n13800) );
  XOR U13347 ( .A(n13799), .B(n13505), .Z(n13802) );
  XNOR U13348 ( .A(p_input[6599]), .B(n13803), .Z(n13505) );
  AND U13349 ( .A(n275), .B(n13804), .Z(n13803) );
  XOR U13350 ( .A(p_input[6631]), .B(p_input[6599]), .Z(n13804) );
  XNOR U13351 ( .A(n13502), .B(n13799), .Z(n13801) );
  XOR U13352 ( .A(n13805), .B(n13806), .Z(n13502) );
  AND U13353 ( .A(n273), .B(n13807), .Z(n13806) );
  XOR U13354 ( .A(p_input[6567]), .B(p_input[6535]), .Z(n13807) );
  XOR U13355 ( .A(n13808), .B(n13809), .Z(n13799) );
  AND U13356 ( .A(n13810), .B(n13811), .Z(n13809) );
  XOR U13357 ( .A(n13808), .B(n13517), .Z(n13811) );
  XNOR U13358 ( .A(p_input[6598]), .B(n13812), .Z(n13517) );
  AND U13359 ( .A(n275), .B(n13813), .Z(n13812) );
  XOR U13360 ( .A(p_input[6630]), .B(p_input[6598]), .Z(n13813) );
  XNOR U13361 ( .A(n13514), .B(n13808), .Z(n13810) );
  XOR U13362 ( .A(n13814), .B(n13815), .Z(n13514) );
  AND U13363 ( .A(n273), .B(n13816), .Z(n13815) );
  XOR U13364 ( .A(p_input[6566]), .B(p_input[6534]), .Z(n13816) );
  XOR U13365 ( .A(n13817), .B(n13818), .Z(n13808) );
  AND U13366 ( .A(n13819), .B(n13820), .Z(n13818) );
  XOR U13367 ( .A(n13817), .B(n13529), .Z(n13820) );
  XNOR U13368 ( .A(p_input[6597]), .B(n13821), .Z(n13529) );
  AND U13369 ( .A(n275), .B(n13822), .Z(n13821) );
  XOR U13370 ( .A(p_input[6629]), .B(p_input[6597]), .Z(n13822) );
  XNOR U13371 ( .A(n13526), .B(n13817), .Z(n13819) );
  XOR U13372 ( .A(n13823), .B(n13824), .Z(n13526) );
  AND U13373 ( .A(n273), .B(n13825), .Z(n13824) );
  XOR U13374 ( .A(p_input[6565]), .B(p_input[6533]), .Z(n13825) );
  XOR U13375 ( .A(n13826), .B(n13827), .Z(n13817) );
  AND U13376 ( .A(n13828), .B(n13829), .Z(n13827) );
  XOR U13377 ( .A(n13826), .B(n13541), .Z(n13829) );
  XNOR U13378 ( .A(p_input[6596]), .B(n13830), .Z(n13541) );
  AND U13379 ( .A(n275), .B(n13831), .Z(n13830) );
  XOR U13380 ( .A(p_input[6628]), .B(p_input[6596]), .Z(n13831) );
  XNOR U13381 ( .A(n13538), .B(n13826), .Z(n13828) );
  XOR U13382 ( .A(n13832), .B(n13833), .Z(n13538) );
  AND U13383 ( .A(n273), .B(n13834), .Z(n13833) );
  XOR U13384 ( .A(p_input[6564]), .B(p_input[6532]), .Z(n13834) );
  XOR U13385 ( .A(n13835), .B(n13836), .Z(n13826) );
  AND U13386 ( .A(n13837), .B(n13838), .Z(n13836) );
  XOR U13387 ( .A(n13835), .B(n13553), .Z(n13838) );
  XNOR U13388 ( .A(p_input[6595]), .B(n13839), .Z(n13553) );
  AND U13389 ( .A(n275), .B(n13840), .Z(n13839) );
  XOR U13390 ( .A(p_input[6627]), .B(p_input[6595]), .Z(n13840) );
  XNOR U13391 ( .A(n13550), .B(n13835), .Z(n13837) );
  XOR U13392 ( .A(n13841), .B(n13842), .Z(n13550) );
  AND U13393 ( .A(n273), .B(n13843), .Z(n13842) );
  XOR U13394 ( .A(p_input[6563]), .B(p_input[6531]), .Z(n13843) );
  XOR U13395 ( .A(n13844), .B(n13845), .Z(n13835) );
  AND U13396 ( .A(n13846), .B(n13847), .Z(n13845) );
  XOR U13397 ( .A(n13844), .B(n13565), .Z(n13847) );
  XNOR U13398 ( .A(p_input[6594]), .B(n13848), .Z(n13565) );
  AND U13399 ( .A(n275), .B(n13849), .Z(n13848) );
  XOR U13400 ( .A(p_input[6626]), .B(p_input[6594]), .Z(n13849) );
  XNOR U13401 ( .A(n13562), .B(n13844), .Z(n13846) );
  XOR U13402 ( .A(n13850), .B(n13851), .Z(n13562) );
  AND U13403 ( .A(n273), .B(n13852), .Z(n13851) );
  XOR U13404 ( .A(p_input[6562]), .B(p_input[6530]), .Z(n13852) );
  XOR U13405 ( .A(n13853), .B(n13854), .Z(n13844) );
  AND U13406 ( .A(n13855), .B(n13856), .Z(n13854) );
  XNOR U13407 ( .A(n13857), .B(n13578), .Z(n13856) );
  XNOR U13408 ( .A(p_input[6593]), .B(n13858), .Z(n13578) );
  AND U13409 ( .A(n275), .B(n13859), .Z(n13858) );
  XNOR U13410 ( .A(p_input[6625]), .B(n13860), .Z(n13859) );
  IV U13411 ( .A(p_input[6593]), .Z(n13860) );
  XNOR U13412 ( .A(n13575), .B(n13853), .Z(n13855) );
  XNOR U13413 ( .A(p_input[6529]), .B(n13861), .Z(n13575) );
  AND U13414 ( .A(n273), .B(n13862), .Z(n13861) );
  XOR U13415 ( .A(p_input[6561]), .B(p_input[6529]), .Z(n13862) );
  IV U13416 ( .A(n13857), .Z(n13853) );
  AND U13417 ( .A(n13583), .B(n13586), .Z(n13857) );
  XOR U13418 ( .A(p_input[6592]), .B(n13863), .Z(n13586) );
  AND U13419 ( .A(n275), .B(n13864), .Z(n13863) );
  XOR U13420 ( .A(p_input[6624]), .B(p_input[6592]), .Z(n13864) );
  XOR U13421 ( .A(n13865), .B(n13866), .Z(n275) );
  AND U13422 ( .A(n13867), .B(n13868), .Z(n13866) );
  XNOR U13423 ( .A(p_input[6655]), .B(n13865), .Z(n13868) );
  XOR U13424 ( .A(n13865), .B(p_input[6623]), .Z(n13867) );
  XOR U13425 ( .A(n13869), .B(n13870), .Z(n13865) );
  AND U13426 ( .A(n13871), .B(n13872), .Z(n13870) );
  XNOR U13427 ( .A(p_input[6654]), .B(n13869), .Z(n13872) );
  XOR U13428 ( .A(n13869), .B(p_input[6622]), .Z(n13871) );
  XOR U13429 ( .A(n13873), .B(n13874), .Z(n13869) );
  AND U13430 ( .A(n13875), .B(n13876), .Z(n13874) );
  XNOR U13431 ( .A(p_input[6653]), .B(n13873), .Z(n13876) );
  XOR U13432 ( .A(n13873), .B(p_input[6621]), .Z(n13875) );
  XOR U13433 ( .A(n13877), .B(n13878), .Z(n13873) );
  AND U13434 ( .A(n13879), .B(n13880), .Z(n13878) );
  XNOR U13435 ( .A(p_input[6652]), .B(n13877), .Z(n13880) );
  XOR U13436 ( .A(n13877), .B(p_input[6620]), .Z(n13879) );
  XOR U13437 ( .A(n13881), .B(n13882), .Z(n13877) );
  AND U13438 ( .A(n13883), .B(n13884), .Z(n13882) );
  XNOR U13439 ( .A(p_input[6651]), .B(n13881), .Z(n13884) );
  XOR U13440 ( .A(n13881), .B(p_input[6619]), .Z(n13883) );
  XOR U13441 ( .A(n13885), .B(n13886), .Z(n13881) );
  AND U13442 ( .A(n13887), .B(n13888), .Z(n13886) );
  XNOR U13443 ( .A(p_input[6650]), .B(n13885), .Z(n13888) );
  XOR U13444 ( .A(n13885), .B(p_input[6618]), .Z(n13887) );
  XOR U13445 ( .A(n13889), .B(n13890), .Z(n13885) );
  AND U13446 ( .A(n13891), .B(n13892), .Z(n13890) );
  XNOR U13447 ( .A(p_input[6649]), .B(n13889), .Z(n13892) );
  XOR U13448 ( .A(n13889), .B(p_input[6617]), .Z(n13891) );
  XOR U13449 ( .A(n13893), .B(n13894), .Z(n13889) );
  AND U13450 ( .A(n13895), .B(n13896), .Z(n13894) );
  XNOR U13451 ( .A(p_input[6648]), .B(n13893), .Z(n13896) );
  XOR U13452 ( .A(n13893), .B(p_input[6616]), .Z(n13895) );
  XOR U13453 ( .A(n13897), .B(n13898), .Z(n13893) );
  AND U13454 ( .A(n13899), .B(n13900), .Z(n13898) );
  XNOR U13455 ( .A(p_input[6647]), .B(n13897), .Z(n13900) );
  XOR U13456 ( .A(n13897), .B(p_input[6615]), .Z(n13899) );
  XOR U13457 ( .A(n13901), .B(n13902), .Z(n13897) );
  AND U13458 ( .A(n13903), .B(n13904), .Z(n13902) );
  XNOR U13459 ( .A(p_input[6646]), .B(n13901), .Z(n13904) );
  XOR U13460 ( .A(n13901), .B(p_input[6614]), .Z(n13903) );
  XOR U13461 ( .A(n13905), .B(n13906), .Z(n13901) );
  AND U13462 ( .A(n13907), .B(n13908), .Z(n13906) );
  XNOR U13463 ( .A(p_input[6645]), .B(n13905), .Z(n13908) );
  XOR U13464 ( .A(n13905), .B(p_input[6613]), .Z(n13907) );
  XOR U13465 ( .A(n13909), .B(n13910), .Z(n13905) );
  AND U13466 ( .A(n13911), .B(n13912), .Z(n13910) );
  XNOR U13467 ( .A(p_input[6644]), .B(n13909), .Z(n13912) );
  XOR U13468 ( .A(n13909), .B(p_input[6612]), .Z(n13911) );
  XOR U13469 ( .A(n13913), .B(n13914), .Z(n13909) );
  AND U13470 ( .A(n13915), .B(n13916), .Z(n13914) );
  XNOR U13471 ( .A(p_input[6643]), .B(n13913), .Z(n13916) );
  XOR U13472 ( .A(n13913), .B(p_input[6611]), .Z(n13915) );
  XOR U13473 ( .A(n13917), .B(n13918), .Z(n13913) );
  AND U13474 ( .A(n13919), .B(n13920), .Z(n13918) );
  XNOR U13475 ( .A(p_input[6642]), .B(n13917), .Z(n13920) );
  XOR U13476 ( .A(n13917), .B(p_input[6610]), .Z(n13919) );
  XOR U13477 ( .A(n13921), .B(n13922), .Z(n13917) );
  AND U13478 ( .A(n13923), .B(n13924), .Z(n13922) );
  XNOR U13479 ( .A(p_input[6641]), .B(n13921), .Z(n13924) );
  XOR U13480 ( .A(n13921), .B(p_input[6609]), .Z(n13923) );
  XOR U13481 ( .A(n13925), .B(n13926), .Z(n13921) );
  AND U13482 ( .A(n13927), .B(n13928), .Z(n13926) );
  XNOR U13483 ( .A(p_input[6640]), .B(n13925), .Z(n13928) );
  XOR U13484 ( .A(n13925), .B(p_input[6608]), .Z(n13927) );
  XOR U13485 ( .A(n13929), .B(n13930), .Z(n13925) );
  AND U13486 ( .A(n13931), .B(n13932), .Z(n13930) );
  XNOR U13487 ( .A(p_input[6639]), .B(n13929), .Z(n13932) );
  XOR U13488 ( .A(n13929), .B(p_input[6607]), .Z(n13931) );
  XOR U13489 ( .A(n13933), .B(n13934), .Z(n13929) );
  AND U13490 ( .A(n13935), .B(n13936), .Z(n13934) );
  XNOR U13491 ( .A(p_input[6638]), .B(n13933), .Z(n13936) );
  XOR U13492 ( .A(n13933), .B(p_input[6606]), .Z(n13935) );
  XOR U13493 ( .A(n13937), .B(n13938), .Z(n13933) );
  AND U13494 ( .A(n13939), .B(n13940), .Z(n13938) );
  XNOR U13495 ( .A(p_input[6637]), .B(n13937), .Z(n13940) );
  XOR U13496 ( .A(n13937), .B(p_input[6605]), .Z(n13939) );
  XOR U13497 ( .A(n13941), .B(n13942), .Z(n13937) );
  AND U13498 ( .A(n13943), .B(n13944), .Z(n13942) );
  XNOR U13499 ( .A(p_input[6636]), .B(n13941), .Z(n13944) );
  XOR U13500 ( .A(n13941), .B(p_input[6604]), .Z(n13943) );
  XOR U13501 ( .A(n13945), .B(n13946), .Z(n13941) );
  AND U13502 ( .A(n13947), .B(n13948), .Z(n13946) );
  XNOR U13503 ( .A(p_input[6635]), .B(n13945), .Z(n13948) );
  XOR U13504 ( .A(n13945), .B(p_input[6603]), .Z(n13947) );
  XOR U13505 ( .A(n13949), .B(n13950), .Z(n13945) );
  AND U13506 ( .A(n13951), .B(n13952), .Z(n13950) );
  XNOR U13507 ( .A(p_input[6634]), .B(n13949), .Z(n13952) );
  XOR U13508 ( .A(n13949), .B(p_input[6602]), .Z(n13951) );
  XOR U13509 ( .A(n13953), .B(n13954), .Z(n13949) );
  AND U13510 ( .A(n13955), .B(n13956), .Z(n13954) );
  XNOR U13511 ( .A(p_input[6633]), .B(n13953), .Z(n13956) );
  XOR U13512 ( .A(n13953), .B(p_input[6601]), .Z(n13955) );
  XOR U13513 ( .A(n13957), .B(n13958), .Z(n13953) );
  AND U13514 ( .A(n13959), .B(n13960), .Z(n13958) );
  XNOR U13515 ( .A(p_input[6632]), .B(n13957), .Z(n13960) );
  XOR U13516 ( .A(n13957), .B(p_input[6600]), .Z(n13959) );
  XOR U13517 ( .A(n13961), .B(n13962), .Z(n13957) );
  AND U13518 ( .A(n13963), .B(n13964), .Z(n13962) );
  XNOR U13519 ( .A(p_input[6631]), .B(n13961), .Z(n13964) );
  XOR U13520 ( .A(n13961), .B(p_input[6599]), .Z(n13963) );
  XOR U13521 ( .A(n13965), .B(n13966), .Z(n13961) );
  AND U13522 ( .A(n13967), .B(n13968), .Z(n13966) );
  XNOR U13523 ( .A(p_input[6630]), .B(n13965), .Z(n13968) );
  XOR U13524 ( .A(n13965), .B(p_input[6598]), .Z(n13967) );
  XOR U13525 ( .A(n13969), .B(n13970), .Z(n13965) );
  AND U13526 ( .A(n13971), .B(n13972), .Z(n13970) );
  XNOR U13527 ( .A(p_input[6629]), .B(n13969), .Z(n13972) );
  XOR U13528 ( .A(n13969), .B(p_input[6597]), .Z(n13971) );
  XOR U13529 ( .A(n13973), .B(n13974), .Z(n13969) );
  AND U13530 ( .A(n13975), .B(n13976), .Z(n13974) );
  XNOR U13531 ( .A(p_input[6628]), .B(n13973), .Z(n13976) );
  XOR U13532 ( .A(n13973), .B(p_input[6596]), .Z(n13975) );
  XOR U13533 ( .A(n13977), .B(n13978), .Z(n13973) );
  AND U13534 ( .A(n13979), .B(n13980), .Z(n13978) );
  XNOR U13535 ( .A(p_input[6627]), .B(n13977), .Z(n13980) );
  XOR U13536 ( .A(n13977), .B(p_input[6595]), .Z(n13979) );
  XOR U13537 ( .A(n13981), .B(n13982), .Z(n13977) );
  AND U13538 ( .A(n13983), .B(n13984), .Z(n13982) );
  XNOR U13539 ( .A(p_input[6626]), .B(n13981), .Z(n13984) );
  XOR U13540 ( .A(n13981), .B(p_input[6594]), .Z(n13983) );
  XNOR U13541 ( .A(n13985), .B(n13986), .Z(n13981) );
  AND U13542 ( .A(n13987), .B(n13988), .Z(n13986) );
  XOR U13543 ( .A(p_input[6625]), .B(n13985), .Z(n13988) );
  XNOR U13544 ( .A(p_input[6593]), .B(n13985), .Z(n13987) );
  AND U13545 ( .A(p_input[6624]), .B(n13989), .Z(n13985) );
  IV U13546 ( .A(p_input[6592]), .Z(n13989) );
  XNOR U13547 ( .A(p_input[6528]), .B(n13990), .Z(n13583) );
  AND U13548 ( .A(n273), .B(n13991), .Z(n13990) );
  XOR U13549 ( .A(p_input[6560]), .B(p_input[6528]), .Z(n13991) );
  XOR U13550 ( .A(n13992), .B(n13993), .Z(n273) );
  AND U13551 ( .A(n13994), .B(n13995), .Z(n13993) );
  XNOR U13552 ( .A(p_input[6591]), .B(n13992), .Z(n13995) );
  XOR U13553 ( .A(n13992), .B(p_input[6559]), .Z(n13994) );
  XOR U13554 ( .A(n13996), .B(n13997), .Z(n13992) );
  AND U13555 ( .A(n13998), .B(n13999), .Z(n13997) );
  XNOR U13556 ( .A(p_input[6590]), .B(n13996), .Z(n13999) );
  XNOR U13557 ( .A(n13996), .B(n13598), .Z(n13998) );
  IV U13558 ( .A(p_input[6558]), .Z(n13598) );
  XOR U13559 ( .A(n14000), .B(n14001), .Z(n13996) );
  AND U13560 ( .A(n14002), .B(n14003), .Z(n14001) );
  XNOR U13561 ( .A(p_input[6589]), .B(n14000), .Z(n14003) );
  XNOR U13562 ( .A(n14000), .B(n13607), .Z(n14002) );
  IV U13563 ( .A(p_input[6557]), .Z(n13607) );
  XOR U13564 ( .A(n14004), .B(n14005), .Z(n14000) );
  AND U13565 ( .A(n14006), .B(n14007), .Z(n14005) );
  XNOR U13566 ( .A(p_input[6588]), .B(n14004), .Z(n14007) );
  XNOR U13567 ( .A(n14004), .B(n13616), .Z(n14006) );
  IV U13568 ( .A(p_input[6556]), .Z(n13616) );
  XOR U13569 ( .A(n14008), .B(n14009), .Z(n14004) );
  AND U13570 ( .A(n14010), .B(n14011), .Z(n14009) );
  XNOR U13571 ( .A(p_input[6587]), .B(n14008), .Z(n14011) );
  XNOR U13572 ( .A(n14008), .B(n13625), .Z(n14010) );
  IV U13573 ( .A(p_input[6555]), .Z(n13625) );
  XOR U13574 ( .A(n14012), .B(n14013), .Z(n14008) );
  AND U13575 ( .A(n14014), .B(n14015), .Z(n14013) );
  XNOR U13576 ( .A(p_input[6586]), .B(n14012), .Z(n14015) );
  XNOR U13577 ( .A(n14012), .B(n13634), .Z(n14014) );
  IV U13578 ( .A(p_input[6554]), .Z(n13634) );
  XOR U13579 ( .A(n14016), .B(n14017), .Z(n14012) );
  AND U13580 ( .A(n14018), .B(n14019), .Z(n14017) );
  XNOR U13581 ( .A(p_input[6585]), .B(n14016), .Z(n14019) );
  XNOR U13582 ( .A(n14016), .B(n13643), .Z(n14018) );
  IV U13583 ( .A(p_input[6553]), .Z(n13643) );
  XOR U13584 ( .A(n14020), .B(n14021), .Z(n14016) );
  AND U13585 ( .A(n14022), .B(n14023), .Z(n14021) );
  XNOR U13586 ( .A(p_input[6584]), .B(n14020), .Z(n14023) );
  XNOR U13587 ( .A(n14020), .B(n13652), .Z(n14022) );
  IV U13588 ( .A(p_input[6552]), .Z(n13652) );
  XOR U13589 ( .A(n14024), .B(n14025), .Z(n14020) );
  AND U13590 ( .A(n14026), .B(n14027), .Z(n14025) );
  XNOR U13591 ( .A(p_input[6583]), .B(n14024), .Z(n14027) );
  XNOR U13592 ( .A(n14024), .B(n13661), .Z(n14026) );
  IV U13593 ( .A(p_input[6551]), .Z(n13661) );
  XOR U13594 ( .A(n14028), .B(n14029), .Z(n14024) );
  AND U13595 ( .A(n14030), .B(n14031), .Z(n14029) );
  XNOR U13596 ( .A(p_input[6582]), .B(n14028), .Z(n14031) );
  XNOR U13597 ( .A(n14028), .B(n13670), .Z(n14030) );
  IV U13598 ( .A(p_input[6550]), .Z(n13670) );
  XOR U13599 ( .A(n14032), .B(n14033), .Z(n14028) );
  AND U13600 ( .A(n14034), .B(n14035), .Z(n14033) );
  XNOR U13601 ( .A(p_input[6581]), .B(n14032), .Z(n14035) );
  XNOR U13602 ( .A(n14032), .B(n13679), .Z(n14034) );
  IV U13603 ( .A(p_input[6549]), .Z(n13679) );
  XOR U13604 ( .A(n14036), .B(n14037), .Z(n14032) );
  AND U13605 ( .A(n14038), .B(n14039), .Z(n14037) );
  XNOR U13606 ( .A(p_input[6580]), .B(n14036), .Z(n14039) );
  XNOR U13607 ( .A(n14036), .B(n13688), .Z(n14038) );
  IV U13608 ( .A(p_input[6548]), .Z(n13688) );
  XOR U13609 ( .A(n14040), .B(n14041), .Z(n14036) );
  AND U13610 ( .A(n14042), .B(n14043), .Z(n14041) );
  XNOR U13611 ( .A(p_input[6579]), .B(n14040), .Z(n14043) );
  XNOR U13612 ( .A(n14040), .B(n13697), .Z(n14042) );
  IV U13613 ( .A(p_input[6547]), .Z(n13697) );
  XOR U13614 ( .A(n14044), .B(n14045), .Z(n14040) );
  AND U13615 ( .A(n14046), .B(n14047), .Z(n14045) );
  XNOR U13616 ( .A(p_input[6578]), .B(n14044), .Z(n14047) );
  XNOR U13617 ( .A(n14044), .B(n13706), .Z(n14046) );
  IV U13618 ( .A(p_input[6546]), .Z(n13706) );
  XOR U13619 ( .A(n14048), .B(n14049), .Z(n14044) );
  AND U13620 ( .A(n14050), .B(n14051), .Z(n14049) );
  XNOR U13621 ( .A(p_input[6577]), .B(n14048), .Z(n14051) );
  XNOR U13622 ( .A(n14048), .B(n13715), .Z(n14050) );
  IV U13623 ( .A(p_input[6545]), .Z(n13715) );
  XOR U13624 ( .A(n14052), .B(n14053), .Z(n14048) );
  AND U13625 ( .A(n14054), .B(n14055), .Z(n14053) );
  XNOR U13626 ( .A(p_input[6576]), .B(n14052), .Z(n14055) );
  XNOR U13627 ( .A(n14052), .B(n13724), .Z(n14054) );
  IV U13628 ( .A(p_input[6544]), .Z(n13724) );
  XOR U13629 ( .A(n14056), .B(n14057), .Z(n14052) );
  AND U13630 ( .A(n14058), .B(n14059), .Z(n14057) );
  XNOR U13631 ( .A(p_input[6575]), .B(n14056), .Z(n14059) );
  XNOR U13632 ( .A(n14056), .B(n13733), .Z(n14058) );
  IV U13633 ( .A(p_input[6543]), .Z(n13733) );
  XOR U13634 ( .A(n14060), .B(n14061), .Z(n14056) );
  AND U13635 ( .A(n14062), .B(n14063), .Z(n14061) );
  XNOR U13636 ( .A(p_input[6574]), .B(n14060), .Z(n14063) );
  XNOR U13637 ( .A(n14060), .B(n13742), .Z(n14062) );
  IV U13638 ( .A(p_input[6542]), .Z(n13742) );
  XOR U13639 ( .A(n14064), .B(n14065), .Z(n14060) );
  AND U13640 ( .A(n14066), .B(n14067), .Z(n14065) );
  XNOR U13641 ( .A(p_input[6573]), .B(n14064), .Z(n14067) );
  XNOR U13642 ( .A(n14064), .B(n13751), .Z(n14066) );
  IV U13643 ( .A(p_input[6541]), .Z(n13751) );
  XOR U13644 ( .A(n14068), .B(n14069), .Z(n14064) );
  AND U13645 ( .A(n14070), .B(n14071), .Z(n14069) );
  XNOR U13646 ( .A(p_input[6572]), .B(n14068), .Z(n14071) );
  XNOR U13647 ( .A(n14068), .B(n13760), .Z(n14070) );
  IV U13648 ( .A(p_input[6540]), .Z(n13760) );
  XOR U13649 ( .A(n14072), .B(n14073), .Z(n14068) );
  AND U13650 ( .A(n14074), .B(n14075), .Z(n14073) );
  XNOR U13651 ( .A(p_input[6571]), .B(n14072), .Z(n14075) );
  XNOR U13652 ( .A(n14072), .B(n13769), .Z(n14074) );
  IV U13653 ( .A(p_input[6539]), .Z(n13769) );
  XOR U13654 ( .A(n14076), .B(n14077), .Z(n14072) );
  AND U13655 ( .A(n14078), .B(n14079), .Z(n14077) );
  XNOR U13656 ( .A(p_input[6570]), .B(n14076), .Z(n14079) );
  XNOR U13657 ( .A(n14076), .B(n13778), .Z(n14078) );
  IV U13658 ( .A(p_input[6538]), .Z(n13778) );
  XOR U13659 ( .A(n14080), .B(n14081), .Z(n14076) );
  AND U13660 ( .A(n14082), .B(n14083), .Z(n14081) );
  XNOR U13661 ( .A(p_input[6569]), .B(n14080), .Z(n14083) );
  XNOR U13662 ( .A(n14080), .B(n13787), .Z(n14082) );
  IV U13663 ( .A(p_input[6537]), .Z(n13787) );
  XOR U13664 ( .A(n14084), .B(n14085), .Z(n14080) );
  AND U13665 ( .A(n14086), .B(n14087), .Z(n14085) );
  XNOR U13666 ( .A(p_input[6568]), .B(n14084), .Z(n14087) );
  XNOR U13667 ( .A(n14084), .B(n13796), .Z(n14086) );
  IV U13668 ( .A(p_input[6536]), .Z(n13796) );
  XOR U13669 ( .A(n14088), .B(n14089), .Z(n14084) );
  AND U13670 ( .A(n14090), .B(n14091), .Z(n14089) );
  XNOR U13671 ( .A(p_input[6567]), .B(n14088), .Z(n14091) );
  XNOR U13672 ( .A(n14088), .B(n13805), .Z(n14090) );
  IV U13673 ( .A(p_input[6535]), .Z(n13805) );
  XOR U13674 ( .A(n14092), .B(n14093), .Z(n14088) );
  AND U13675 ( .A(n14094), .B(n14095), .Z(n14093) );
  XNOR U13676 ( .A(p_input[6566]), .B(n14092), .Z(n14095) );
  XNOR U13677 ( .A(n14092), .B(n13814), .Z(n14094) );
  IV U13678 ( .A(p_input[6534]), .Z(n13814) );
  XOR U13679 ( .A(n14096), .B(n14097), .Z(n14092) );
  AND U13680 ( .A(n14098), .B(n14099), .Z(n14097) );
  XNOR U13681 ( .A(p_input[6565]), .B(n14096), .Z(n14099) );
  XNOR U13682 ( .A(n14096), .B(n13823), .Z(n14098) );
  IV U13683 ( .A(p_input[6533]), .Z(n13823) );
  XOR U13684 ( .A(n14100), .B(n14101), .Z(n14096) );
  AND U13685 ( .A(n14102), .B(n14103), .Z(n14101) );
  XNOR U13686 ( .A(p_input[6564]), .B(n14100), .Z(n14103) );
  XNOR U13687 ( .A(n14100), .B(n13832), .Z(n14102) );
  IV U13688 ( .A(p_input[6532]), .Z(n13832) );
  XOR U13689 ( .A(n14104), .B(n14105), .Z(n14100) );
  AND U13690 ( .A(n14106), .B(n14107), .Z(n14105) );
  XNOR U13691 ( .A(p_input[6563]), .B(n14104), .Z(n14107) );
  XNOR U13692 ( .A(n14104), .B(n13841), .Z(n14106) );
  IV U13693 ( .A(p_input[6531]), .Z(n13841) );
  XOR U13694 ( .A(n14108), .B(n14109), .Z(n14104) );
  AND U13695 ( .A(n14110), .B(n14111), .Z(n14109) );
  XNOR U13696 ( .A(p_input[6562]), .B(n14108), .Z(n14111) );
  XNOR U13697 ( .A(n14108), .B(n13850), .Z(n14110) );
  IV U13698 ( .A(p_input[6530]), .Z(n13850) );
  XNOR U13699 ( .A(n14112), .B(n14113), .Z(n14108) );
  AND U13700 ( .A(n14114), .B(n14115), .Z(n14113) );
  XOR U13701 ( .A(p_input[6561]), .B(n14112), .Z(n14115) );
  XNOR U13702 ( .A(p_input[6529]), .B(n14112), .Z(n14114) );
  AND U13703 ( .A(p_input[6560]), .B(n14116), .Z(n14112) );
  IV U13704 ( .A(p_input[6528]), .Z(n14116) );
  XOR U13705 ( .A(n14117), .B(n14118), .Z(n13206) );
  AND U13706 ( .A(n477), .B(n14119), .Z(n14118) );
  XNOR U13707 ( .A(n14120), .B(n14117), .Z(n14119) );
  XOR U13708 ( .A(n14121), .B(n14122), .Z(n477) );
  AND U13709 ( .A(n14123), .B(n14124), .Z(n14122) );
  XNOR U13710 ( .A(n13221), .B(n14121), .Z(n14124) );
  AND U13711 ( .A(p_input[6527]), .B(p_input[6495]), .Z(n13221) );
  XNOR U13712 ( .A(n14121), .B(n13218), .Z(n14123) );
  IV U13713 ( .A(n14125), .Z(n13218) );
  AND U13714 ( .A(p_input[6431]), .B(p_input[6463]), .Z(n14125) );
  XOR U13715 ( .A(n14126), .B(n14127), .Z(n14121) );
  AND U13716 ( .A(n14128), .B(n14129), .Z(n14127) );
  XOR U13717 ( .A(n14126), .B(n13233), .Z(n14129) );
  XNOR U13718 ( .A(p_input[6494]), .B(n14130), .Z(n13233) );
  AND U13719 ( .A(n279), .B(n14131), .Z(n14130) );
  XOR U13720 ( .A(p_input[6526]), .B(p_input[6494]), .Z(n14131) );
  XNOR U13721 ( .A(n13230), .B(n14126), .Z(n14128) );
  XOR U13722 ( .A(n14132), .B(n14133), .Z(n13230) );
  AND U13723 ( .A(n276), .B(n14134), .Z(n14133) );
  XOR U13724 ( .A(p_input[6462]), .B(p_input[6430]), .Z(n14134) );
  XOR U13725 ( .A(n14135), .B(n14136), .Z(n14126) );
  AND U13726 ( .A(n14137), .B(n14138), .Z(n14136) );
  XOR U13727 ( .A(n14135), .B(n13245), .Z(n14138) );
  XNOR U13728 ( .A(p_input[6493]), .B(n14139), .Z(n13245) );
  AND U13729 ( .A(n279), .B(n14140), .Z(n14139) );
  XOR U13730 ( .A(p_input[6525]), .B(p_input[6493]), .Z(n14140) );
  XNOR U13731 ( .A(n13242), .B(n14135), .Z(n14137) );
  XOR U13732 ( .A(n14141), .B(n14142), .Z(n13242) );
  AND U13733 ( .A(n276), .B(n14143), .Z(n14142) );
  XOR U13734 ( .A(p_input[6461]), .B(p_input[6429]), .Z(n14143) );
  XOR U13735 ( .A(n14144), .B(n14145), .Z(n14135) );
  AND U13736 ( .A(n14146), .B(n14147), .Z(n14145) );
  XOR U13737 ( .A(n14144), .B(n13257), .Z(n14147) );
  XNOR U13738 ( .A(p_input[6492]), .B(n14148), .Z(n13257) );
  AND U13739 ( .A(n279), .B(n14149), .Z(n14148) );
  XOR U13740 ( .A(p_input[6524]), .B(p_input[6492]), .Z(n14149) );
  XNOR U13741 ( .A(n13254), .B(n14144), .Z(n14146) );
  XOR U13742 ( .A(n14150), .B(n14151), .Z(n13254) );
  AND U13743 ( .A(n276), .B(n14152), .Z(n14151) );
  XOR U13744 ( .A(p_input[6460]), .B(p_input[6428]), .Z(n14152) );
  XOR U13745 ( .A(n14153), .B(n14154), .Z(n14144) );
  AND U13746 ( .A(n14155), .B(n14156), .Z(n14154) );
  XOR U13747 ( .A(n14153), .B(n13269), .Z(n14156) );
  XNOR U13748 ( .A(p_input[6491]), .B(n14157), .Z(n13269) );
  AND U13749 ( .A(n279), .B(n14158), .Z(n14157) );
  XOR U13750 ( .A(p_input[6523]), .B(p_input[6491]), .Z(n14158) );
  XNOR U13751 ( .A(n13266), .B(n14153), .Z(n14155) );
  XOR U13752 ( .A(n14159), .B(n14160), .Z(n13266) );
  AND U13753 ( .A(n276), .B(n14161), .Z(n14160) );
  XOR U13754 ( .A(p_input[6459]), .B(p_input[6427]), .Z(n14161) );
  XOR U13755 ( .A(n14162), .B(n14163), .Z(n14153) );
  AND U13756 ( .A(n14164), .B(n14165), .Z(n14163) );
  XOR U13757 ( .A(n14162), .B(n13281), .Z(n14165) );
  XNOR U13758 ( .A(p_input[6490]), .B(n14166), .Z(n13281) );
  AND U13759 ( .A(n279), .B(n14167), .Z(n14166) );
  XOR U13760 ( .A(p_input[6522]), .B(p_input[6490]), .Z(n14167) );
  XNOR U13761 ( .A(n13278), .B(n14162), .Z(n14164) );
  XOR U13762 ( .A(n14168), .B(n14169), .Z(n13278) );
  AND U13763 ( .A(n276), .B(n14170), .Z(n14169) );
  XOR U13764 ( .A(p_input[6458]), .B(p_input[6426]), .Z(n14170) );
  XOR U13765 ( .A(n14171), .B(n14172), .Z(n14162) );
  AND U13766 ( .A(n14173), .B(n14174), .Z(n14172) );
  XOR U13767 ( .A(n14171), .B(n13293), .Z(n14174) );
  XNOR U13768 ( .A(p_input[6489]), .B(n14175), .Z(n13293) );
  AND U13769 ( .A(n279), .B(n14176), .Z(n14175) );
  XOR U13770 ( .A(p_input[6521]), .B(p_input[6489]), .Z(n14176) );
  XNOR U13771 ( .A(n13290), .B(n14171), .Z(n14173) );
  XOR U13772 ( .A(n14177), .B(n14178), .Z(n13290) );
  AND U13773 ( .A(n276), .B(n14179), .Z(n14178) );
  XOR U13774 ( .A(p_input[6457]), .B(p_input[6425]), .Z(n14179) );
  XOR U13775 ( .A(n14180), .B(n14181), .Z(n14171) );
  AND U13776 ( .A(n14182), .B(n14183), .Z(n14181) );
  XOR U13777 ( .A(n14180), .B(n13305), .Z(n14183) );
  XNOR U13778 ( .A(p_input[6488]), .B(n14184), .Z(n13305) );
  AND U13779 ( .A(n279), .B(n14185), .Z(n14184) );
  XOR U13780 ( .A(p_input[6520]), .B(p_input[6488]), .Z(n14185) );
  XNOR U13781 ( .A(n13302), .B(n14180), .Z(n14182) );
  XOR U13782 ( .A(n14186), .B(n14187), .Z(n13302) );
  AND U13783 ( .A(n276), .B(n14188), .Z(n14187) );
  XOR U13784 ( .A(p_input[6456]), .B(p_input[6424]), .Z(n14188) );
  XOR U13785 ( .A(n14189), .B(n14190), .Z(n14180) );
  AND U13786 ( .A(n14191), .B(n14192), .Z(n14190) );
  XOR U13787 ( .A(n14189), .B(n13317), .Z(n14192) );
  XNOR U13788 ( .A(p_input[6487]), .B(n14193), .Z(n13317) );
  AND U13789 ( .A(n279), .B(n14194), .Z(n14193) );
  XOR U13790 ( .A(p_input[6519]), .B(p_input[6487]), .Z(n14194) );
  XNOR U13791 ( .A(n13314), .B(n14189), .Z(n14191) );
  XOR U13792 ( .A(n14195), .B(n14196), .Z(n13314) );
  AND U13793 ( .A(n276), .B(n14197), .Z(n14196) );
  XOR U13794 ( .A(p_input[6455]), .B(p_input[6423]), .Z(n14197) );
  XOR U13795 ( .A(n14198), .B(n14199), .Z(n14189) );
  AND U13796 ( .A(n14200), .B(n14201), .Z(n14199) );
  XOR U13797 ( .A(n14198), .B(n13329), .Z(n14201) );
  XNOR U13798 ( .A(p_input[6486]), .B(n14202), .Z(n13329) );
  AND U13799 ( .A(n279), .B(n14203), .Z(n14202) );
  XOR U13800 ( .A(p_input[6518]), .B(p_input[6486]), .Z(n14203) );
  XNOR U13801 ( .A(n13326), .B(n14198), .Z(n14200) );
  XOR U13802 ( .A(n14204), .B(n14205), .Z(n13326) );
  AND U13803 ( .A(n276), .B(n14206), .Z(n14205) );
  XOR U13804 ( .A(p_input[6454]), .B(p_input[6422]), .Z(n14206) );
  XOR U13805 ( .A(n14207), .B(n14208), .Z(n14198) );
  AND U13806 ( .A(n14209), .B(n14210), .Z(n14208) );
  XOR U13807 ( .A(n14207), .B(n13341), .Z(n14210) );
  XNOR U13808 ( .A(p_input[6485]), .B(n14211), .Z(n13341) );
  AND U13809 ( .A(n279), .B(n14212), .Z(n14211) );
  XOR U13810 ( .A(p_input[6517]), .B(p_input[6485]), .Z(n14212) );
  XNOR U13811 ( .A(n13338), .B(n14207), .Z(n14209) );
  XOR U13812 ( .A(n14213), .B(n14214), .Z(n13338) );
  AND U13813 ( .A(n276), .B(n14215), .Z(n14214) );
  XOR U13814 ( .A(p_input[6453]), .B(p_input[6421]), .Z(n14215) );
  XOR U13815 ( .A(n14216), .B(n14217), .Z(n14207) );
  AND U13816 ( .A(n14218), .B(n14219), .Z(n14217) );
  XOR U13817 ( .A(n14216), .B(n13353), .Z(n14219) );
  XNOR U13818 ( .A(p_input[6484]), .B(n14220), .Z(n13353) );
  AND U13819 ( .A(n279), .B(n14221), .Z(n14220) );
  XOR U13820 ( .A(p_input[6516]), .B(p_input[6484]), .Z(n14221) );
  XNOR U13821 ( .A(n13350), .B(n14216), .Z(n14218) );
  XOR U13822 ( .A(n14222), .B(n14223), .Z(n13350) );
  AND U13823 ( .A(n276), .B(n14224), .Z(n14223) );
  XOR U13824 ( .A(p_input[6452]), .B(p_input[6420]), .Z(n14224) );
  XOR U13825 ( .A(n14225), .B(n14226), .Z(n14216) );
  AND U13826 ( .A(n14227), .B(n14228), .Z(n14226) );
  XOR U13827 ( .A(n14225), .B(n13365), .Z(n14228) );
  XNOR U13828 ( .A(p_input[6483]), .B(n14229), .Z(n13365) );
  AND U13829 ( .A(n279), .B(n14230), .Z(n14229) );
  XOR U13830 ( .A(p_input[6515]), .B(p_input[6483]), .Z(n14230) );
  XNOR U13831 ( .A(n13362), .B(n14225), .Z(n14227) );
  XOR U13832 ( .A(n14231), .B(n14232), .Z(n13362) );
  AND U13833 ( .A(n276), .B(n14233), .Z(n14232) );
  XOR U13834 ( .A(p_input[6451]), .B(p_input[6419]), .Z(n14233) );
  XOR U13835 ( .A(n14234), .B(n14235), .Z(n14225) );
  AND U13836 ( .A(n14236), .B(n14237), .Z(n14235) );
  XOR U13837 ( .A(n14234), .B(n13377), .Z(n14237) );
  XNOR U13838 ( .A(p_input[6482]), .B(n14238), .Z(n13377) );
  AND U13839 ( .A(n279), .B(n14239), .Z(n14238) );
  XOR U13840 ( .A(p_input[6514]), .B(p_input[6482]), .Z(n14239) );
  XNOR U13841 ( .A(n13374), .B(n14234), .Z(n14236) );
  XOR U13842 ( .A(n14240), .B(n14241), .Z(n13374) );
  AND U13843 ( .A(n276), .B(n14242), .Z(n14241) );
  XOR U13844 ( .A(p_input[6450]), .B(p_input[6418]), .Z(n14242) );
  XOR U13845 ( .A(n14243), .B(n14244), .Z(n14234) );
  AND U13846 ( .A(n14245), .B(n14246), .Z(n14244) );
  XOR U13847 ( .A(n14243), .B(n13389), .Z(n14246) );
  XNOR U13848 ( .A(p_input[6481]), .B(n14247), .Z(n13389) );
  AND U13849 ( .A(n279), .B(n14248), .Z(n14247) );
  XOR U13850 ( .A(p_input[6513]), .B(p_input[6481]), .Z(n14248) );
  XNOR U13851 ( .A(n13386), .B(n14243), .Z(n14245) );
  XOR U13852 ( .A(n14249), .B(n14250), .Z(n13386) );
  AND U13853 ( .A(n276), .B(n14251), .Z(n14250) );
  XOR U13854 ( .A(p_input[6449]), .B(p_input[6417]), .Z(n14251) );
  XOR U13855 ( .A(n14252), .B(n14253), .Z(n14243) );
  AND U13856 ( .A(n14254), .B(n14255), .Z(n14253) );
  XOR U13857 ( .A(n14252), .B(n13401), .Z(n14255) );
  XNOR U13858 ( .A(p_input[6480]), .B(n14256), .Z(n13401) );
  AND U13859 ( .A(n279), .B(n14257), .Z(n14256) );
  XOR U13860 ( .A(p_input[6512]), .B(p_input[6480]), .Z(n14257) );
  XNOR U13861 ( .A(n13398), .B(n14252), .Z(n14254) );
  XOR U13862 ( .A(n14258), .B(n14259), .Z(n13398) );
  AND U13863 ( .A(n276), .B(n14260), .Z(n14259) );
  XOR U13864 ( .A(p_input[6448]), .B(p_input[6416]), .Z(n14260) );
  XOR U13865 ( .A(n14261), .B(n14262), .Z(n14252) );
  AND U13866 ( .A(n14263), .B(n14264), .Z(n14262) );
  XOR U13867 ( .A(n14261), .B(n13413), .Z(n14264) );
  XNOR U13868 ( .A(p_input[6479]), .B(n14265), .Z(n13413) );
  AND U13869 ( .A(n279), .B(n14266), .Z(n14265) );
  XOR U13870 ( .A(p_input[6511]), .B(p_input[6479]), .Z(n14266) );
  XNOR U13871 ( .A(n13410), .B(n14261), .Z(n14263) );
  XOR U13872 ( .A(n14267), .B(n14268), .Z(n13410) );
  AND U13873 ( .A(n276), .B(n14269), .Z(n14268) );
  XOR U13874 ( .A(p_input[6447]), .B(p_input[6415]), .Z(n14269) );
  XOR U13875 ( .A(n14270), .B(n14271), .Z(n14261) );
  AND U13876 ( .A(n14272), .B(n14273), .Z(n14271) );
  XOR U13877 ( .A(n14270), .B(n13425), .Z(n14273) );
  XNOR U13878 ( .A(p_input[6478]), .B(n14274), .Z(n13425) );
  AND U13879 ( .A(n279), .B(n14275), .Z(n14274) );
  XOR U13880 ( .A(p_input[6510]), .B(p_input[6478]), .Z(n14275) );
  XNOR U13881 ( .A(n13422), .B(n14270), .Z(n14272) );
  XOR U13882 ( .A(n14276), .B(n14277), .Z(n13422) );
  AND U13883 ( .A(n276), .B(n14278), .Z(n14277) );
  XOR U13884 ( .A(p_input[6446]), .B(p_input[6414]), .Z(n14278) );
  XOR U13885 ( .A(n14279), .B(n14280), .Z(n14270) );
  AND U13886 ( .A(n14281), .B(n14282), .Z(n14280) );
  XOR U13887 ( .A(n14279), .B(n13437), .Z(n14282) );
  XNOR U13888 ( .A(p_input[6477]), .B(n14283), .Z(n13437) );
  AND U13889 ( .A(n279), .B(n14284), .Z(n14283) );
  XOR U13890 ( .A(p_input[6509]), .B(p_input[6477]), .Z(n14284) );
  XNOR U13891 ( .A(n13434), .B(n14279), .Z(n14281) );
  XOR U13892 ( .A(n14285), .B(n14286), .Z(n13434) );
  AND U13893 ( .A(n276), .B(n14287), .Z(n14286) );
  XOR U13894 ( .A(p_input[6445]), .B(p_input[6413]), .Z(n14287) );
  XOR U13895 ( .A(n14288), .B(n14289), .Z(n14279) );
  AND U13896 ( .A(n14290), .B(n14291), .Z(n14289) );
  XOR U13897 ( .A(n14288), .B(n13449), .Z(n14291) );
  XNOR U13898 ( .A(p_input[6476]), .B(n14292), .Z(n13449) );
  AND U13899 ( .A(n279), .B(n14293), .Z(n14292) );
  XOR U13900 ( .A(p_input[6508]), .B(p_input[6476]), .Z(n14293) );
  XNOR U13901 ( .A(n13446), .B(n14288), .Z(n14290) );
  XOR U13902 ( .A(n14294), .B(n14295), .Z(n13446) );
  AND U13903 ( .A(n276), .B(n14296), .Z(n14295) );
  XOR U13904 ( .A(p_input[6444]), .B(p_input[6412]), .Z(n14296) );
  XOR U13905 ( .A(n14297), .B(n14298), .Z(n14288) );
  AND U13906 ( .A(n14299), .B(n14300), .Z(n14298) );
  XOR U13907 ( .A(n14297), .B(n13461), .Z(n14300) );
  XNOR U13908 ( .A(p_input[6475]), .B(n14301), .Z(n13461) );
  AND U13909 ( .A(n279), .B(n14302), .Z(n14301) );
  XOR U13910 ( .A(p_input[6507]), .B(p_input[6475]), .Z(n14302) );
  XNOR U13911 ( .A(n13458), .B(n14297), .Z(n14299) );
  XOR U13912 ( .A(n14303), .B(n14304), .Z(n13458) );
  AND U13913 ( .A(n276), .B(n14305), .Z(n14304) );
  XOR U13914 ( .A(p_input[6443]), .B(p_input[6411]), .Z(n14305) );
  XOR U13915 ( .A(n14306), .B(n14307), .Z(n14297) );
  AND U13916 ( .A(n14308), .B(n14309), .Z(n14307) );
  XOR U13917 ( .A(n14306), .B(n13473), .Z(n14309) );
  XNOR U13918 ( .A(p_input[6474]), .B(n14310), .Z(n13473) );
  AND U13919 ( .A(n279), .B(n14311), .Z(n14310) );
  XOR U13920 ( .A(p_input[6506]), .B(p_input[6474]), .Z(n14311) );
  XNOR U13921 ( .A(n13470), .B(n14306), .Z(n14308) );
  XOR U13922 ( .A(n14312), .B(n14313), .Z(n13470) );
  AND U13923 ( .A(n276), .B(n14314), .Z(n14313) );
  XOR U13924 ( .A(p_input[6442]), .B(p_input[6410]), .Z(n14314) );
  XOR U13925 ( .A(n14315), .B(n14316), .Z(n14306) );
  AND U13926 ( .A(n14317), .B(n14318), .Z(n14316) );
  XOR U13927 ( .A(n14315), .B(n13485), .Z(n14318) );
  XNOR U13928 ( .A(p_input[6473]), .B(n14319), .Z(n13485) );
  AND U13929 ( .A(n279), .B(n14320), .Z(n14319) );
  XOR U13930 ( .A(p_input[6505]), .B(p_input[6473]), .Z(n14320) );
  XNOR U13931 ( .A(n13482), .B(n14315), .Z(n14317) );
  XOR U13932 ( .A(n14321), .B(n14322), .Z(n13482) );
  AND U13933 ( .A(n276), .B(n14323), .Z(n14322) );
  XOR U13934 ( .A(p_input[6441]), .B(p_input[6409]), .Z(n14323) );
  XOR U13935 ( .A(n14324), .B(n14325), .Z(n14315) );
  AND U13936 ( .A(n14326), .B(n14327), .Z(n14325) );
  XOR U13937 ( .A(n14324), .B(n13497), .Z(n14327) );
  XNOR U13938 ( .A(p_input[6472]), .B(n14328), .Z(n13497) );
  AND U13939 ( .A(n279), .B(n14329), .Z(n14328) );
  XOR U13940 ( .A(p_input[6504]), .B(p_input[6472]), .Z(n14329) );
  XNOR U13941 ( .A(n13494), .B(n14324), .Z(n14326) );
  XOR U13942 ( .A(n14330), .B(n14331), .Z(n13494) );
  AND U13943 ( .A(n276), .B(n14332), .Z(n14331) );
  XOR U13944 ( .A(p_input[6440]), .B(p_input[6408]), .Z(n14332) );
  XOR U13945 ( .A(n14333), .B(n14334), .Z(n14324) );
  AND U13946 ( .A(n14335), .B(n14336), .Z(n14334) );
  XOR U13947 ( .A(n14333), .B(n13509), .Z(n14336) );
  XNOR U13948 ( .A(p_input[6471]), .B(n14337), .Z(n13509) );
  AND U13949 ( .A(n279), .B(n14338), .Z(n14337) );
  XOR U13950 ( .A(p_input[6503]), .B(p_input[6471]), .Z(n14338) );
  XNOR U13951 ( .A(n13506), .B(n14333), .Z(n14335) );
  XOR U13952 ( .A(n14339), .B(n14340), .Z(n13506) );
  AND U13953 ( .A(n276), .B(n14341), .Z(n14340) );
  XOR U13954 ( .A(p_input[6439]), .B(p_input[6407]), .Z(n14341) );
  XOR U13955 ( .A(n14342), .B(n14343), .Z(n14333) );
  AND U13956 ( .A(n14344), .B(n14345), .Z(n14343) );
  XOR U13957 ( .A(n14342), .B(n13521), .Z(n14345) );
  XNOR U13958 ( .A(p_input[6470]), .B(n14346), .Z(n13521) );
  AND U13959 ( .A(n279), .B(n14347), .Z(n14346) );
  XOR U13960 ( .A(p_input[6502]), .B(p_input[6470]), .Z(n14347) );
  XNOR U13961 ( .A(n13518), .B(n14342), .Z(n14344) );
  XOR U13962 ( .A(n14348), .B(n14349), .Z(n13518) );
  AND U13963 ( .A(n276), .B(n14350), .Z(n14349) );
  XOR U13964 ( .A(p_input[6438]), .B(p_input[6406]), .Z(n14350) );
  XOR U13965 ( .A(n14351), .B(n14352), .Z(n14342) );
  AND U13966 ( .A(n14353), .B(n14354), .Z(n14352) );
  XOR U13967 ( .A(n14351), .B(n13533), .Z(n14354) );
  XNOR U13968 ( .A(p_input[6469]), .B(n14355), .Z(n13533) );
  AND U13969 ( .A(n279), .B(n14356), .Z(n14355) );
  XOR U13970 ( .A(p_input[6501]), .B(p_input[6469]), .Z(n14356) );
  XNOR U13971 ( .A(n13530), .B(n14351), .Z(n14353) );
  XOR U13972 ( .A(n14357), .B(n14358), .Z(n13530) );
  AND U13973 ( .A(n276), .B(n14359), .Z(n14358) );
  XOR U13974 ( .A(p_input[6437]), .B(p_input[6405]), .Z(n14359) );
  XOR U13975 ( .A(n14360), .B(n14361), .Z(n14351) );
  AND U13976 ( .A(n14362), .B(n14363), .Z(n14361) );
  XOR U13977 ( .A(n14360), .B(n13545), .Z(n14363) );
  XNOR U13978 ( .A(p_input[6468]), .B(n14364), .Z(n13545) );
  AND U13979 ( .A(n279), .B(n14365), .Z(n14364) );
  XOR U13980 ( .A(p_input[6500]), .B(p_input[6468]), .Z(n14365) );
  XNOR U13981 ( .A(n13542), .B(n14360), .Z(n14362) );
  XOR U13982 ( .A(n14366), .B(n14367), .Z(n13542) );
  AND U13983 ( .A(n276), .B(n14368), .Z(n14367) );
  XOR U13984 ( .A(p_input[6436]), .B(p_input[6404]), .Z(n14368) );
  XOR U13985 ( .A(n14369), .B(n14370), .Z(n14360) );
  AND U13986 ( .A(n14371), .B(n14372), .Z(n14370) );
  XOR U13987 ( .A(n14369), .B(n13557), .Z(n14372) );
  XNOR U13988 ( .A(p_input[6467]), .B(n14373), .Z(n13557) );
  AND U13989 ( .A(n279), .B(n14374), .Z(n14373) );
  XOR U13990 ( .A(p_input[6499]), .B(p_input[6467]), .Z(n14374) );
  XNOR U13991 ( .A(n13554), .B(n14369), .Z(n14371) );
  XOR U13992 ( .A(n14375), .B(n14376), .Z(n13554) );
  AND U13993 ( .A(n276), .B(n14377), .Z(n14376) );
  XOR U13994 ( .A(p_input[6435]), .B(p_input[6403]), .Z(n14377) );
  XOR U13995 ( .A(n14378), .B(n14379), .Z(n14369) );
  AND U13996 ( .A(n14380), .B(n14381), .Z(n14379) );
  XOR U13997 ( .A(n14378), .B(n13569), .Z(n14381) );
  XNOR U13998 ( .A(p_input[6466]), .B(n14382), .Z(n13569) );
  AND U13999 ( .A(n279), .B(n14383), .Z(n14382) );
  XOR U14000 ( .A(p_input[6498]), .B(p_input[6466]), .Z(n14383) );
  XNOR U14001 ( .A(n13566), .B(n14378), .Z(n14380) );
  XOR U14002 ( .A(n14384), .B(n14385), .Z(n13566) );
  AND U14003 ( .A(n276), .B(n14386), .Z(n14385) );
  XOR U14004 ( .A(p_input[6434]), .B(p_input[6402]), .Z(n14386) );
  XOR U14005 ( .A(n14387), .B(n14388), .Z(n14378) );
  AND U14006 ( .A(n14389), .B(n14390), .Z(n14388) );
  XNOR U14007 ( .A(n14391), .B(n13582), .Z(n14390) );
  XNOR U14008 ( .A(p_input[6465]), .B(n14392), .Z(n13582) );
  AND U14009 ( .A(n279), .B(n14393), .Z(n14392) );
  XNOR U14010 ( .A(p_input[6497]), .B(n14394), .Z(n14393) );
  IV U14011 ( .A(p_input[6465]), .Z(n14394) );
  XNOR U14012 ( .A(n13579), .B(n14387), .Z(n14389) );
  XNOR U14013 ( .A(p_input[6401]), .B(n14395), .Z(n13579) );
  AND U14014 ( .A(n276), .B(n14396), .Z(n14395) );
  XOR U14015 ( .A(p_input[6433]), .B(p_input[6401]), .Z(n14396) );
  IV U14016 ( .A(n14391), .Z(n14387) );
  AND U14017 ( .A(n14117), .B(n14120), .Z(n14391) );
  XOR U14018 ( .A(p_input[6464]), .B(n14397), .Z(n14120) );
  AND U14019 ( .A(n279), .B(n14398), .Z(n14397) );
  XOR U14020 ( .A(p_input[6496]), .B(p_input[6464]), .Z(n14398) );
  XOR U14021 ( .A(n14399), .B(n14400), .Z(n279) );
  AND U14022 ( .A(n14401), .B(n14402), .Z(n14400) );
  XNOR U14023 ( .A(p_input[6527]), .B(n14399), .Z(n14402) );
  XOR U14024 ( .A(n14399), .B(p_input[6495]), .Z(n14401) );
  XOR U14025 ( .A(n14403), .B(n14404), .Z(n14399) );
  AND U14026 ( .A(n14405), .B(n14406), .Z(n14404) );
  XNOR U14027 ( .A(p_input[6526]), .B(n14403), .Z(n14406) );
  XOR U14028 ( .A(n14403), .B(p_input[6494]), .Z(n14405) );
  XOR U14029 ( .A(n14407), .B(n14408), .Z(n14403) );
  AND U14030 ( .A(n14409), .B(n14410), .Z(n14408) );
  XNOR U14031 ( .A(p_input[6525]), .B(n14407), .Z(n14410) );
  XOR U14032 ( .A(n14407), .B(p_input[6493]), .Z(n14409) );
  XOR U14033 ( .A(n14411), .B(n14412), .Z(n14407) );
  AND U14034 ( .A(n14413), .B(n14414), .Z(n14412) );
  XNOR U14035 ( .A(p_input[6524]), .B(n14411), .Z(n14414) );
  XOR U14036 ( .A(n14411), .B(p_input[6492]), .Z(n14413) );
  XOR U14037 ( .A(n14415), .B(n14416), .Z(n14411) );
  AND U14038 ( .A(n14417), .B(n14418), .Z(n14416) );
  XNOR U14039 ( .A(p_input[6523]), .B(n14415), .Z(n14418) );
  XOR U14040 ( .A(n14415), .B(p_input[6491]), .Z(n14417) );
  XOR U14041 ( .A(n14419), .B(n14420), .Z(n14415) );
  AND U14042 ( .A(n14421), .B(n14422), .Z(n14420) );
  XNOR U14043 ( .A(p_input[6522]), .B(n14419), .Z(n14422) );
  XOR U14044 ( .A(n14419), .B(p_input[6490]), .Z(n14421) );
  XOR U14045 ( .A(n14423), .B(n14424), .Z(n14419) );
  AND U14046 ( .A(n14425), .B(n14426), .Z(n14424) );
  XNOR U14047 ( .A(p_input[6521]), .B(n14423), .Z(n14426) );
  XOR U14048 ( .A(n14423), .B(p_input[6489]), .Z(n14425) );
  XOR U14049 ( .A(n14427), .B(n14428), .Z(n14423) );
  AND U14050 ( .A(n14429), .B(n14430), .Z(n14428) );
  XNOR U14051 ( .A(p_input[6520]), .B(n14427), .Z(n14430) );
  XOR U14052 ( .A(n14427), .B(p_input[6488]), .Z(n14429) );
  XOR U14053 ( .A(n14431), .B(n14432), .Z(n14427) );
  AND U14054 ( .A(n14433), .B(n14434), .Z(n14432) );
  XNOR U14055 ( .A(p_input[6519]), .B(n14431), .Z(n14434) );
  XOR U14056 ( .A(n14431), .B(p_input[6487]), .Z(n14433) );
  XOR U14057 ( .A(n14435), .B(n14436), .Z(n14431) );
  AND U14058 ( .A(n14437), .B(n14438), .Z(n14436) );
  XNOR U14059 ( .A(p_input[6518]), .B(n14435), .Z(n14438) );
  XOR U14060 ( .A(n14435), .B(p_input[6486]), .Z(n14437) );
  XOR U14061 ( .A(n14439), .B(n14440), .Z(n14435) );
  AND U14062 ( .A(n14441), .B(n14442), .Z(n14440) );
  XNOR U14063 ( .A(p_input[6517]), .B(n14439), .Z(n14442) );
  XOR U14064 ( .A(n14439), .B(p_input[6485]), .Z(n14441) );
  XOR U14065 ( .A(n14443), .B(n14444), .Z(n14439) );
  AND U14066 ( .A(n14445), .B(n14446), .Z(n14444) );
  XNOR U14067 ( .A(p_input[6516]), .B(n14443), .Z(n14446) );
  XOR U14068 ( .A(n14443), .B(p_input[6484]), .Z(n14445) );
  XOR U14069 ( .A(n14447), .B(n14448), .Z(n14443) );
  AND U14070 ( .A(n14449), .B(n14450), .Z(n14448) );
  XNOR U14071 ( .A(p_input[6515]), .B(n14447), .Z(n14450) );
  XOR U14072 ( .A(n14447), .B(p_input[6483]), .Z(n14449) );
  XOR U14073 ( .A(n14451), .B(n14452), .Z(n14447) );
  AND U14074 ( .A(n14453), .B(n14454), .Z(n14452) );
  XNOR U14075 ( .A(p_input[6514]), .B(n14451), .Z(n14454) );
  XOR U14076 ( .A(n14451), .B(p_input[6482]), .Z(n14453) );
  XOR U14077 ( .A(n14455), .B(n14456), .Z(n14451) );
  AND U14078 ( .A(n14457), .B(n14458), .Z(n14456) );
  XNOR U14079 ( .A(p_input[6513]), .B(n14455), .Z(n14458) );
  XOR U14080 ( .A(n14455), .B(p_input[6481]), .Z(n14457) );
  XOR U14081 ( .A(n14459), .B(n14460), .Z(n14455) );
  AND U14082 ( .A(n14461), .B(n14462), .Z(n14460) );
  XNOR U14083 ( .A(p_input[6512]), .B(n14459), .Z(n14462) );
  XOR U14084 ( .A(n14459), .B(p_input[6480]), .Z(n14461) );
  XOR U14085 ( .A(n14463), .B(n14464), .Z(n14459) );
  AND U14086 ( .A(n14465), .B(n14466), .Z(n14464) );
  XNOR U14087 ( .A(p_input[6511]), .B(n14463), .Z(n14466) );
  XOR U14088 ( .A(n14463), .B(p_input[6479]), .Z(n14465) );
  XOR U14089 ( .A(n14467), .B(n14468), .Z(n14463) );
  AND U14090 ( .A(n14469), .B(n14470), .Z(n14468) );
  XNOR U14091 ( .A(p_input[6510]), .B(n14467), .Z(n14470) );
  XOR U14092 ( .A(n14467), .B(p_input[6478]), .Z(n14469) );
  XOR U14093 ( .A(n14471), .B(n14472), .Z(n14467) );
  AND U14094 ( .A(n14473), .B(n14474), .Z(n14472) );
  XNOR U14095 ( .A(p_input[6509]), .B(n14471), .Z(n14474) );
  XOR U14096 ( .A(n14471), .B(p_input[6477]), .Z(n14473) );
  XOR U14097 ( .A(n14475), .B(n14476), .Z(n14471) );
  AND U14098 ( .A(n14477), .B(n14478), .Z(n14476) );
  XNOR U14099 ( .A(p_input[6508]), .B(n14475), .Z(n14478) );
  XOR U14100 ( .A(n14475), .B(p_input[6476]), .Z(n14477) );
  XOR U14101 ( .A(n14479), .B(n14480), .Z(n14475) );
  AND U14102 ( .A(n14481), .B(n14482), .Z(n14480) );
  XNOR U14103 ( .A(p_input[6507]), .B(n14479), .Z(n14482) );
  XOR U14104 ( .A(n14479), .B(p_input[6475]), .Z(n14481) );
  XOR U14105 ( .A(n14483), .B(n14484), .Z(n14479) );
  AND U14106 ( .A(n14485), .B(n14486), .Z(n14484) );
  XNOR U14107 ( .A(p_input[6506]), .B(n14483), .Z(n14486) );
  XOR U14108 ( .A(n14483), .B(p_input[6474]), .Z(n14485) );
  XOR U14109 ( .A(n14487), .B(n14488), .Z(n14483) );
  AND U14110 ( .A(n14489), .B(n14490), .Z(n14488) );
  XNOR U14111 ( .A(p_input[6505]), .B(n14487), .Z(n14490) );
  XOR U14112 ( .A(n14487), .B(p_input[6473]), .Z(n14489) );
  XOR U14113 ( .A(n14491), .B(n14492), .Z(n14487) );
  AND U14114 ( .A(n14493), .B(n14494), .Z(n14492) );
  XNOR U14115 ( .A(p_input[6504]), .B(n14491), .Z(n14494) );
  XOR U14116 ( .A(n14491), .B(p_input[6472]), .Z(n14493) );
  XOR U14117 ( .A(n14495), .B(n14496), .Z(n14491) );
  AND U14118 ( .A(n14497), .B(n14498), .Z(n14496) );
  XNOR U14119 ( .A(p_input[6503]), .B(n14495), .Z(n14498) );
  XOR U14120 ( .A(n14495), .B(p_input[6471]), .Z(n14497) );
  XOR U14121 ( .A(n14499), .B(n14500), .Z(n14495) );
  AND U14122 ( .A(n14501), .B(n14502), .Z(n14500) );
  XNOR U14123 ( .A(p_input[6502]), .B(n14499), .Z(n14502) );
  XOR U14124 ( .A(n14499), .B(p_input[6470]), .Z(n14501) );
  XOR U14125 ( .A(n14503), .B(n14504), .Z(n14499) );
  AND U14126 ( .A(n14505), .B(n14506), .Z(n14504) );
  XNOR U14127 ( .A(p_input[6501]), .B(n14503), .Z(n14506) );
  XOR U14128 ( .A(n14503), .B(p_input[6469]), .Z(n14505) );
  XOR U14129 ( .A(n14507), .B(n14508), .Z(n14503) );
  AND U14130 ( .A(n14509), .B(n14510), .Z(n14508) );
  XNOR U14131 ( .A(p_input[6500]), .B(n14507), .Z(n14510) );
  XOR U14132 ( .A(n14507), .B(p_input[6468]), .Z(n14509) );
  XOR U14133 ( .A(n14511), .B(n14512), .Z(n14507) );
  AND U14134 ( .A(n14513), .B(n14514), .Z(n14512) );
  XNOR U14135 ( .A(p_input[6499]), .B(n14511), .Z(n14514) );
  XOR U14136 ( .A(n14511), .B(p_input[6467]), .Z(n14513) );
  XOR U14137 ( .A(n14515), .B(n14516), .Z(n14511) );
  AND U14138 ( .A(n14517), .B(n14518), .Z(n14516) );
  XNOR U14139 ( .A(p_input[6498]), .B(n14515), .Z(n14518) );
  XOR U14140 ( .A(n14515), .B(p_input[6466]), .Z(n14517) );
  XNOR U14141 ( .A(n14519), .B(n14520), .Z(n14515) );
  AND U14142 ( .A(n14521), .B(n14522), .Z(n14520) );
  XOR U14143 ( .A(p_input[6497]), .B(n14519), .Z(n14522) );
  XNOR U14144 ( .A(p_input[6465]), .B(n14519), .Z(n14521) );
  AND U14145 ( .A(p_input[6496]), .B(n14523), .Z(n14519) );
  IV U14146 ( .A(p_input[6464]), .Z(n14523) );
  XNOR U14147 ( .A(p_input[6400]), .B(n14524), .Z(n14117) );
  AND U14148 ( .A(n276), .B(n14525), .Z(n14524) );
  XOR U14149 ( .A(p_input[6432]), .B(p_input[6400]), .Z(n14525) );
  XOR U14150 ( .A(n14526), .B(n14527), .Z(n276) );
  AND U14151 ( .A(n14528), .B(n14529), .Z(n14527) );
  XNOR U14152 ( .A(p_input[6463]), .B(n14526), .Z(n14529) );
  XOR U14153 ( .A(n14526), .B(p_input[6431]), .Z(n14528) );
  XOR U14154 ( .A(n14530), .B(n14531), .Z(n14526) );
  AND U14155 ( .A(n14532), .B(n14533), .Z(n14531) );
  XNOR U14156 ( .A(p_input[6462]), .B(n14530), .Z(n14533) );
  XNOR U14157 ( .A(n14530), .B(n14132), .Z(n14532) );
  IV U14158 ( .A(p_input[6430]), .Z(n14132) );
  XOR U14159 ( .A(n14534), .B(n14535), .Z(n14530) );
  AND U14160 ( .A(n14536), .B(n14537), .Z(n14535) );
  XNOR U14161 ( .A(p_input[6461]), .B(n14534), .Z(n14537) );
  XNOR U14162 ( .A(n14534), .B(n14141), .Z(n14536) );
  IV U14163 ( .A(p_input[6429]), .Z(n14141) );
  XOR U14164 ( .A(n14538), .B(n14539), .Z(n14534) );
  AND U14165 ( .A(n14540), .B(n14541), .Z(n14539) );
  XNOR U14166 ( .A(p_input[6460]), .B(n14538), .Z(n14541) );
  XNOR U14167 ( .A(n14538), .B(n14150), .Z(n14540) );
  IV U14168 ( .A(p_input[6428]), .Z(n14150) );
  XOR U14169 ( .A(n14542), .B(n14543), .Z(n14538) );
  AND U14170 ( .A(n14544), .B(n14545), .Z(n14543) );
  XNOR U14171 ( .A(p_input[6459]), .B(n14542), .Z(n14545) );
  XNOR U14172 ( .A(n14542), .B(n14159), .Z(n14544) );
  IV U14173 ( .A(p_input[6427]), .Z(n14159) );
  XOR U14174 ( .A(n14546), .B(n14547), .Z(n14542) );
  AND U14175 ( .A(n14548), .B(n14549), .Z(n14547) );
  XNOR U14176 ( .A(p_input[6458]), .B(n14546), .Z(n14549) );
  XNOR U14177 ( .A(n14546), .B(n14168), .Z(n14548) );
  IV U14178 ( .A(p_input[6426]), .Z(n14168) );
  XOR U14179 ( .A(n14550), .B(n14551), .Z(n14546) );
  AND U14180 ( .A(n14552), .B(n14553), .Z(n14551) );
  XNOR U14181 ( .A(p_input[6457]), .B(n14550), .Z(n14553) );
  XNOR U14182 ( .A(n14550), .B(n14177), .Z(n14552) );
  IV U14183 ( .A(p_input[6425]), .Z(n14177) );
  XOR U14184 ( .A(n14554), .B(n14555), .Z(n14550) );
  AND U14185 ( .A(n14556), .B(n14557), .Z(n14555) );
  XNOR U14186 ( .A(p_input[6456]), .B(n14554), .Z(n14557) );
  XNOR U14187 ( .A(n14554), .B(n14186), .Z(n14556) );
  IV U14188 ( .A(p_input[6424]), .Z(n14186) );
  XOR U14189 ( .A(n14558), .B(n14559), .Z(n14554) );
  AND U14190 ( .A(n14560), .B(n14561), .Z(n14559) );
  XNOR U14191 ( .A(p_input[6455]), .B(n14558), .Z(n14561) );
  XNOR U14192 ( .A(n14558), .B(n14195), .Z(n14560) );
  IV U14193 ( .A(p_input[6423]), .Z(n14195) );
  XOR U14194 ( .A(n14562), .B(n14563), .Z(n14558) );
  AND U14195 ( .A(n14564), .B(n14565), .Z(n14563) );
  XNOR U14196 ( .A(p_input[6454]), .B(n14562), .Z(n14565) );
  XNOR U14197 ( .A(n14562), .B(n14204), .Z(n14564) );
  IV U14198 ( .A(p_input[6422]), .Z(n14204) );
  XOR U14199 ( .A(n14566), .B(n14567), .Z(n14562) );
  AND U14200 ( .A(n14568), .B(n14569), .Z(n14567) );
  XNOR U14201 ( .A(p_input[6453]), .B(n14566), .Z(n14569) );
  XNOR U14202 ( .A(n14566), .B(n14213), .Z(n14568) );
  IV U14203 ( .A(p_input[6421]), .Z(n14213) );
  XOR U14204 ( .A(n14570), .B(n14571), .Z(n14566) );
  AND U14205 ( .A(n14572), .B(n14573), .Z(n14571) );
  XNOR U14206 ( .A(p_input[6452]), .B(n14570), .Z(n14573) );
  XNOR U14207 ( .A(n14570), .B(n14222), .Z(n14572) );
  IV U14208 ( .A(p_input[6420]), .Z(n14222) );
  XOR U14209 ( .A(n14574), .B(n14575), .Z(n14570) );
  AND U14210 ( .A(n14576), .B(n14577), .Z(n14575) );
  XNOR U14211 ( .A(p_input[6451]), .B(n14574), .Z(n14577) );
  XNOR U14212 ( .A(n14574), .B(n14231), .Z(n14576) );
  IV U14213 ( .A(p_input[6419]), .Z(n14231) );
  XOR U14214 ( .A(n14578), .B(n14579), .Z(n14574) );
  AND U14215 ( .A(n14580), .B(n14581), .Z(n14579) );
  XNOR U14216 ( .A(p_input[6450]), .B(n14578), .Z(n14581) );
  XNOR U14217 ( .A(n14578), .B(n14240), .Z(n14580) );
  IV U14218 ( .A(p_input[6418]), .Z(n14240) );
  XOR U14219 ( .A(n14582), .B(n14583), .Z(n14578) );
  AND U14220 ( .A(n14584), .B(n14585), .Z(n14583) );
  XNOR U14221 ( .A(p_input[6449]), .B(n14582), .Z(n14585) );
  XNOR U14222 ( .A(n14582), .B(n14249), .Z(n14584) );
  IV U14223 ( .A(p_input[6417]), .Z(n14249) );
  XOR U14224 ( .A(n14586), .B(n14587), .Z(n14582) );
  AND U14225 ( .A(n14588), .B(n14589), .Z(n14587) );
  XNOR U14226 ( .A(p_input[6448]), .B(n14586), .Z(n14589) );
  XNOR U14227 ( .A(n14586), .B(n14258), .Z(n14588) );
  IV U14228 ( .A(p_input[6416]), .Z(n14258) );
  XOR U14229 ( .A(n14590), .B(n14591), .Z(n14586) );
  AND U14230 ( .A(n14592), .B(n14593), .Z(n14591) );
  XNOR U14231 ( .A(p_input[6447]), .B(n14590), .Z(n14593) );
  XNOR U14232 ( .A(n14590), .B(n14267), .Z(n14592) );
  IV U14233 ( .A(p_input[6415]), .Z(n14267) );
  XOR U14234 ( .A(n14594), .B(n14595), .Z(n14590) );
  AND U14235 ( .A(n14596), .B(n14597), .Z(n14595) );
  XNOR U14236 ( .A(p_input[6446]), .B(n14594), .Z(n14597) );
  XNOR U14237 ( .A(n14594), .B(n14276), .Z(n14596) );
  IV U14238 ( .A(p_input[6414]), .Z(n14276) );
  XOR U14239 ( .A(n14598), .B(n14599), .Z(n14594) );
  AND U14240 ( .A(n14600), .B(n14601), .Z(n14599) );
  XNOR U14241 ( .A(p_input[6445]), .B(n14598), .Z(n14601) );
  XNOR U14242 ( .A(n14598), .B(n14285), .Z(n14600) );
  IV U14243 ( .A(p_input[6413]), .Z(n14285) );
  XOR U14244 ( .A(n14602), .B(n14603), .Z(n14598) );
  AND U14245 ( .A(n14604), .B(n14605), .Z(n14603) );
  XNOR U14246 ( .A(p_input[6444]), .B(n14602), .Z(n14605) );
  XNOR U14247 ( .A(n14602), .B(n14294), .Z(n14604) );
  IV U14248 ( .A(p_input[6412]), .Z(n14294) );
  XOR U14249 ( .A(n14606), .B(n14607), .Z(n14602) );
  AND U14250 ( .A(n14608), .B(n14609), .Z(n14607) );
  XNOR U14251 ( .A(p_input[6443]), .B(n14606), .Z(n14609) );
  XNOR U14252 ( .A(n14606), .B(n14303), .Z(n14608) );
  IV U14253 ( .A(p_input[6411]), .Z(n14303) );
  XOR U14254 ( .A(n14610), .B(n14611), .Z(n14606) );
  AND U14255 ( .A(n14612), .B(n14613), .Z(n14611) );
  XNOR U14256 ( .A(p_input[6442]), .B(n14610), .Z(n14613) );
  XNOR U14257 ( .A(n14610), .B(n14312), .Z(n14612) );
  IV U14258 ( .A(p_input[6410]), .Z(n14312) );
  XOR U14259 ( .A(n14614), .B(n14615), .Z(n14610) );
  AND U14260 ( .A(n14616), .B(n14617), .Z(n14615) );
  XNOR U14261 ( .A(p_input[6441]), .B(n14614), .Z(n14617) );
  XNOR U14262 ( .A(n14614), .B(n14321), .Z(n14616) );
  IV U14263 ( .A(p_input[6409]), .Z(n14321) );
  XOR U14264 ( .A(n14618), .B(n14619), .Z(n14614) );
  AND U14265 ( .A(n14620), .B(n14621), .Z(n14619) );
  XNOR U14266 ( .A(p_input[6440]), .B(n14618), .Z(n14621) );
  XNOR U14267 ( .A(n14618), .B(n14330), .Z(n14620) );
  IV U14268 ( .A(p_input[6408]), .Z(n14330) );
  XOR U14269 ( .A(n14622), .B(n14623), .Z(n14618) );
  AND U14270 ( .A(n14624), .B(n14625), .Z(n14623) );
  XNOR U14271 ( .A(p_input[6439]), .B(n14622), .Z(n14625) );
  XNOR U14272 ( .A(n14622), .B(n14339), .Z(n14624) );
  IV U14273 ( .A(p_input[6407]), .Z(n14339) );
  XOR U14274 ( .A(n14626), .B(n14627), .Z(n14622) );
  AND U14275 ( .A(n14628), .B(n14629), .Z(n14627) );
  XNOR U14276 ( .A(p_input[6438]), .B(n14626), .Z(n14629) );
  XNOR U14277 ( .A(n14626), .B(n14348), .Z(n14628) );
  IV U14278 ( .A(p_input[6406]), .Z(n14348) );
  XOR U14279 ( .A(n14630), .B(n14631), .Z(n14626) );
  AND U14280 ( .A(n14632), .B(n14633), .Z(n14631) );
  XNOR U14281 ( .A(p_input[6437]), .B(n14630), .Z(n14633) );
  XNOR U14282 ( .A(n14630), .B(n14357), .Z(n14632) );
  IV U14283 ( .A(p_input[6405]), .Z(n14357) );
  XOR U14284 ( .A(n14634), .B(n14635), .Z(n14630) );
  AND U14285 ( .A(n14636), .B(n14637), .Z(n14635) );
  XNOR U14286 ( .A(p_input[6436]), .B(n14634), .Z(n14637) );
  XNOR U14287 ( .A(n14634), .B(n14366), .Z(n14636) );
  IV U14288 ( .A(p_input[6404]), .Z(n14366) );
  XOR U14289 ( .A(n14638), .B(n14639), .Z(n14634) );
  AND U14290 ( .A(n14640), .B(n14641), .Z(n14639) );
  XNOR U14291 ( .A(p_input[6435]), .B(n14638), .Z(n14641) );
  XNOR U14292 ( .A(n14638), .B(n14375), .Z(n14640) );
  IV U14293 ( .A(p_input[6403]), .Z(n14375) );
  XOR U14294 ( .A(n14642), .B(n14643), .Z(n14638) );
  AND U14295 ( .A(n14644), .B(n14645), .Z(n14643) );
  XNOR U14296 ( .A(p_input[6434]), .B(n14642), .Z(n14645) );
  XNOR U14297 ( .A(n14642), .B(n14384), .Z(n14644) );
  IV U14298 ( .A(p_input[6402]), .Z(n14384) );
  XNOR U14299 ( .A(n14646), .B(n14647), .Z(n14642) );
  AND U14300 ( .A(n14648), .B(n14649), .Z(n14647) );
  XOR U14301 ( .A(p_input[6433]), .B(n14646), .Z(n14649) );
  XNOR U14302 ( .A(p_input[6401]), .B(n14646), .Z(n14648) );
  AND U14303 ( .A(p_input[6432]), .B(n14650), .Z(n14646) );
  IV U14304 ( .A(p_input[6400]), .Z(n14650) );
  XOR U14305 ( .A(n14651), .B(n14652), .Z(n12829) );
  AND U14306 ( .A(n828), .B(n14653), .Z(n14652) );
  XNOR U14307 ( .A(n14654), .B(n14651), .Z(n14653) );
  XOR U14308 ( .A(n14655), .B(n14656), .Z(n828) );
  AND U14309 ( .A(n14657), .B(n14658), .Z(n14656) );
  XOR U14310 ( .A(n14655), .B(n12844), .Z(n14658) );
  XNOR U14311 ( .A(n14659), .B(n14660), .Z(n12844) );
  AND U14312 ( .A(n14661), .B(n483), .Z(n14660) );
  AND U14313 ( .A(n14659), .B(n14662), .Z(n14661) );
  XNOR U14314 ( .A(n12841), .B(n14655), .Z(n14657) );
  XOR U14315 ( .A(n14663), .B(n14664), .Z(n12841) );
  AND U14316 ( .A(n14665), .B(n480), .Z(n14664) );
  NOR U14317 ( .A(n14663), .B(n14666), .Z(n14665) );
  XOR U14318 ( .A(n14667), .B(n14668), .Z(n14655) );
  AND U14319 ( .A(n14669), .B(n14670), .Z(n14668) );
  XOR U14320 ( .A(n14667), .B(n12856), .Z(n14670) );
  XOR U14321 ( .A(n14671), .B(n14672), .Z(n12856) );
  AND U14322 ( .A(n483), .B(n14673), .Z(n14672) );
  XOR U14323 ( .A(n14674), .B(n14671), .Z(n14673) );
  XNOR U14324 ( .A(n12853), .B(n14667), .Z(n14669) );
  XOR U14325 ( .A(n14675), .B(n14676), .Z(n12853) );
  AND U14326 ( .A(n480), .B(n14677), .Z(n14676) );
  XOR U14327 ( .A(n14678), .B(n14675), .Z(n14677) );
  XOR U14328 ( .A(n14679), .B(n14680), .Z(n14667) );
  AND U14329 ( .A(n14681), .B(n14682), .Z(n14680) );
  XOR U14330 ( .A(n14679), .B(n12868), .Z(n14682) );
  XOR U14331 ( .A(n14683), .B(n14684), .Z(n12868) );
  AND U14332 ( .A(n483), .B(n14685), .Z(n14684) );
  XOR U14333 ( .A(n14686), .B(n14683), .Z(n14685) );
  XNOR U14334 ( .A(n12865), .B(n14679), .Z(n14681) );
  XOR U14335 ( .A(n14687), .B(n14688), .Z(n12865) );
  AND U14336 ( .A(n480), .B(n14689), .Z(n14688) );
  XOR U14337 ( .A(n14690), .B(n14687), .Z(n14689) );
  XOR U14338 ( .A(n14691), .B(n14692), .Z(n14679) );
  AND U14339 ( .A(n14693), .B(n14694), .Z(n14692) );
  XOR U14340 ( .A(n14691), .B(n12880), .Z(n14694) );
  XOR U14341 ( .A(n14695), .B(n14696), .Z(n12880) );
  AND U14342 ( .A(n483), .B(n14697), .Z(n14696) );
  XOR U14343 ( .A(n14698), .B(n14695), .Z(n14697) );
  XNOR U14344 ( .A(n12877), .B(n14691), .Z(n14693) );
  XOR U14345 ( .A(n14699), .B(n14700), .Z(n12877) );
  AND U14346 ( .A(n480), .B(n14701), .Z(n14700) );
  XOR U14347 ( .A(n14702), .B(n14699), .Z(n14701) );
  XOR U14348 ( .A(n14703), .B(n14704), .Z(n14691) );
  AND U14349 ( .A(n14705), .B(n14706), .Z(n14704) );
  XOR U14350 ( .A(n14703), .B(n12892), .Z(n14706) );
  XOR U14351 ( .A(n14707), .B(n14708), .Z(n12892) );
  AND U14352 ( .A(n483), .B(n14709), .Z(n14708) );
  XOR U14353 ( .A(n14710), .B(n14707), .Z(n14709) );
  XNOR U14354 ( .A(n12889), .B(n14703), .Z(n14705) );
  XOR U14355 ( .A(n14711), .B(n14712), .Z(n12889) );
  AND U14356 ( .A(n480), .B(n14713), .Z(n14712) );
  XOR U14357 ( .A(n14714), .B(n14711), .Z(n14713) );
  XOR U14358 ( .A(n14715), .B(n14716), .Z(n14703) );
  AND U14359 ( .A(n14717), .B(n14718), .Z(n14716) );
  XOR U14360 ( .A(n14715), .B(n12904), .Z(n14718) );
  XOR U14361 ( .A(n14719), .B(n14720), .Z(n12904) );
  AND U14362 ( .A(n483), .B(n14721), .Z(n14720) );
  XOR U14363 ( .A(n14722), .B(n14719), .Z(n14721) );
  XNOR U14364 ( .A(n12901), .B(n14715), .Z(n14717) );
  XOR U14365 ( .A(n14723), .B(n14724), .Z(n12901) );
  AND U14366 ( .A(n480), .B(n14725), .Z(n14724) );
  XOR U14367 ( .A(n14726), .B(n14723), .Z(n14725) );
  XOR U14368 ( .A(n14727), .B(n14728), .Z(n14715) );
  AND U14369 ( .A(n14729), .B(n14730), .Z(n14728) );
  XOR U14370 ( .A(n14727), .B(n12916), .Z(n14730) );
  XOR U14371 ( .A(n14731), .B(n14732), .Z(n12916) );
  AND U14372 ( .A(n483), .B(n14733), .Z(n14732) );
  XOR U14373 ( .A(n14734), .B(n14731), .Z(n14733) );
  XNOR U14374 ( .A(n12913), .B(n14727), .Z(n14729) );
  XOR U14375 ( .A(n14735), .B(n14736), .Z(n12913) );
  AND U14376 ( .A(n480), .B(n14737), .Z(n14736) );
  XOR U14377 ( .A(n14738), .B(n14735), .Z(n14737) );
  XOR U14378 ( .A(n14739), .B(n14740), .Z(n14727) );
  AND U14379 ( .A(n14741), .B(n14742), .Z(n14740) );
  XOR U14380 ( .A(n14739), .B(n12928), .Z(n14742) );
  XOR U14381 ( .A(n14743), .B(n14744), .Z(n12928) );
  AND U14382 ( .A(n483), .B(n14745), .Z(n14744) );
  XOR U14383 ( .A(n14746), .B(n14743), .Z(n14745) );
  XNOR U14384 ( .A(n12925), .B(n14739), .Z(n14741) );
  XOR U14385 ( .A(n14747), .B(n14748), .Z(n12925) );
  AND U14386 ( .A(n480), .B(n14749), .Z(n14748) );
  XOR U14387 ( .A(n14750), .B(n14747), .Z(n14749) );
  XOR U14388 ( .A(n14751), .B(n14752), .Z(n14739) );
  AND U14389 ( .A(n14753), .B(n14754), .Z(n14752) );
  XOR U14390 ( .A(n14751), .B(n12940), .Z(n14754) );
  XOR U14391 ( .A(n14755), .B(n14756), .Z(n12940) );
  AND U14392 ( .A(n483), .B(n14757), .Z(n14756) );
  XOR U14393 ( .A(n14758), .B(n14755), .Z(n14757) );
  XNOR U14394 ( .A(n12937), .B(n14751), .Z(n14753) );
  XOR U14395 ( .A(n14759), .B(n14760), .Z(n12937) );
  AND U14396 ( .A(n480), .B(n14761), .Z(n14760) );
  XOR U14397 ( .A(n14762), .B(n14759), .Z(n14761) );
  XOR U14398 ( .A(n14763), .B(n14764), .Z(n14751) );
  AND U14399 ( .A(n14765), .B(n14766), .Z(n14764) );
  XOR U14400 ( .A(n14763), .B(n12952), .Z(n14766) );
  XOR U14401 ( .A(n14767), .B(n14768), .Z(n12952) );
  AND U14402 ( .A(n483), .B(n14769), .Z(n14768) );
  XOR U14403 ( .A(n14770), .B(n14767), .Z(n14769) );
  XNOR U14404 ( .A(n12949), .B(n14763), .Z(n14765) );
  XOR U14405 ( .A(n14771), .B(n14772), .Z(n12949) );
  AND U14406 ( .A(n480), .B(n14773), .Z(n14772) );
  XOR U14407 ( .A(n14774), .B(n14771), .Z(n14773) );
  XOR U14408 ( .A(n14775), .B(n14776), .Z(n14763) );
  AND U14409 ( .A(n14777), .B(n14778), .Z(n14776) );
  XOR U14410 ( .A(n14775), .B(n12964), .Z(n14778) );
  XOR U14411 ( .A(n14779), .B(n14780), .Z(n12964) );
  AND U14412 ( .A(n483), .B(n14781), .Z(n14780) );
  XOR U14413 ( .A(n14782), .B(n14779), .Z(n14781) );
  XNOR U14414 ( .A(n12961), .B(n14775), .Z(n14777) );
  XOR U14415 ( .A(n14783), .B(n14784), .Z(n12961) );
  AND U14416 ( .A(n480), .B(n14785), .Z(n14784) );
  XOR U14417 ( .A(n14786), .B(n14783), .Z(n14785) );
  XOR U14418 ( .A(n14787), .B(n14788), .Z(n14775) );
  AND U14419 ( .A(n14789), .B(n14790), .Z(n14788) );
  XOR U14420 ( .A(n14787), .B(n12976), .Z(n14790) );
  XOR U14421 ( .A(n14791), .B(n14792), .Z(n12976) );
  AND U14422 ( .A(n483), .B(n14793), .Z(n14792) );
  XOR U14423 ( .A(n14794), .B(n14791), .Z(n14793) );
  XNOR U14424 ( .A(n12973), .B(n14787), .Z(n14789) );
  XOR U14425 ( .A(n14795), .B(n14796), .Z(n12973) );
  AND U14426 ( .A(n480), .B(n14797), .Z(n14796) );
  XOR U14427 ( .A(n14798), .B(n14795), .Z(n14797) );
  XOR U14428 ( .A(n14799), .B(n14800), .Z(n14787) );
  AND U14429 ( .A(n14801), .B(n14802), .Z(n14800) );
  XOR U14430 ( .A(n14799), .B(n12988), .Z(n14802) );
  XOR U14431 ( .A(n14803), .B(n14804), .Z(n12988) );
  AND U14432 ( .A(n483), .B(n14805), .Z(n14804) );
  XOR U14433 ( .A(n14806), .B(n14803), .Z(n14805) );
  XNOR U14434 ( .A(n12985), .B(n14799), .Z(n14801) );
  XOR U14435 ( .A(n14807), .B(n14808), .Z(n12985) );
  AND U14436 ( .A(n480), .B(n14809), .Z(n14808) );
  XOR U14437 ( .A(n14810), .B(n14807), .Z(n14809) );
  XOR U14438 ( .A(n14811), .B(n14812), .Z(n14799) );
  AND U14439 ( .A(n14813), .B(n14814), .Z(n14812) );
  XOR U14440 ( .A(n14811), .B(n13000), .Z(n14814) );
  XOR U14441 ( .A(n14815), .B(n14816), .Z(n13000) );
  AND U14442 ( .A(n483), .B(n14817), .Z(n14816) );
  XOR U14443 ( .A(n14818), .B(n14815), .Z(n14817) );
  XNOR U14444 ( .A(n12997), .B(n14811), .Z(n14813) );
  XOR U14445 ( .A(n14819), .B(n14820), .Z(n12997) );
  AND U14446 ( .A(n480), .B(n14821), .Z(n14820) );
  XOR U14447 ( .A(n14822), .B(n14819), .Z(n14821) );
  XOR U14448 ( .A(n14823), .B(n14824), .Z(n14811) );
  AND U14449 ( .A(n14825), .B(n14826), .Z(n14824) );
  XOR U14450 ( .A(n14823), .B(n13012), .Z(n14826) );
  XOR U14451 ( .A(n14827), .B(n14828), .Z(n13012) );
  AND U14452 ( .A(n483), .B(n14829), .Z(n14828) );
  XOR U14453 ( .A(n14830), .B(n14827), .Z(n14829) );
  XNOR U14454 ( .A(n13009), .B(n14823), .Z(n14825) );
  XOR U14455 ( .A(n14831), .B(n14832), .Z(n13009) );
  AND U14456 ( .A(n480), .B(n14833), .Z(n14832) );
  XOR U14457 ( .A(n14834), .B(n14831), .Z(n14833) );
  XOR U14458 ( .A(n14835), .B(n14836), .Z(n14823) );
  AND U14459 ( .A(n14837), .B(n14838), .Z(n14836) );
  XOR U14460 ( .A(n14835), .B(n13024), .Z(n14838) );
  XOR U14461 ( .A(n14839), .B(n14840), .Z(n13024) );
  AND U14462 ( .A(n483), .B(n14841), .Z(n14840) );
  XOR U14463 ( .A(n14842), .B(n14839), .Z(n14841) );
  XNOR U14464 ( .A(n13021), .B(n14835), .Z(n14837) );
  XOR U14465 ( .A(n14843), .B(n14844), .Z(n13021) );
  AND U14466 ( .A(n480), .B(n14845), .Z(n14844) );
  XOR U14467 ( .A(n14846), .B(n14843), .Z(n14845) );
  XOR U14468 ( .A(n14847), .B(n14848), .Z(n14835) );
  AND U14469 ( .A(n14849), .B(n14850), .Z(n14848) );
  XOR U14470 ( .A(n14847), .B(n13036), .Z(n14850) );
  XOR U14471 ( .A(n14851), .B(n14852), .Z(n13036) );
  AND U14472 ( .A(n483), .B(n14853), .Z(n14852) );
  XOR U14473 ( .A(n14854), .B(n14851), .Z(n14853) );
  XNOR U14474 ( .A(n13033), .B(n14847), .Z(n14849) );
  XOR U14475 ( .A(n14855), .B(n14856), .Z(n13033) );
  AND U14476 ( .A(n480), .B(n14857), .Z(n14856) );
  XOR U14477 ( .A(n14858), .B(n14855), .Z(n14857) );
  XOR U14478 ( .A(n14859), .B(n14860), .Z(n14847) );
  AND U14479 ( .A(n14861), .B(n14862), .Z(n14860) );
  XOR U14480 ( .A(n14859), .B(n13048), .Z(n14862) );
  XOR U14481 ( .A(n14863), .B(n14864), .Z(n13048) );
  AND U14482 ( .A(n483), .B(n14865), .Z(n14864) );
  XOR U14483 ( .A(n14866), .B(n14863), .Z(n14865) );
  XNOR U14484 ( .A(n13045), .B(n14859), .Z(n14861) );
  XOR U14485 ( .A(n14867), .B(n14868), .Z(n13045) );
  AND U14486 ( .A(n480), .B(n14869), .Z(n14868) );
  XOR U14487 ( .A(n14870), .B(n14867), .Z(n14869) );
  XOR U14488 ( .A(n14871), .B(n14872), .Z(n14859) );
  AND U14489 ( .A(n14873), .B(n14874), .Z(n14872) );
  XOR U14490 ( .A(n14871), .B(n13060), .Z(n14874) );
  XOR U14491 ( .A(n14875), .B(n14876), .Z(n13060) );
  AND U14492 ( .A(n483), .B(n14877), .Z(n14876) );
  XOR U14493 ( .A(n14878), .B(n14875), .Z(n14877) );
  XNOR U14494 ( .A(n13057), .B(n14871), .Z(n14873) );
  XOR U14495 ( .A(n14879), .B(n14880), .Z(n13057) );
  AND U14496 ( .A(n480), .B(n14881), .Z(n14880) );
  XOR U14497 ( .A(n14882), .B(n14879), .Z(n14881) );
  XOR U14498 ( .A(n14883), .B(n14884), .Z(n14871) );
  AND U14499 ( .A(n14885), .B(n14886), .Z(n14884) );
  XOR U14500 ( .A(n14883), .B(n13072), .Z(n14886) );
  XOR U14501 ( .A(n14887), .B(n14888), .Z(n13072) );
  AND U14502 ( .A(n483), .B(n14889), .Z(n14888) );
  XOR U14503 ( .A(n14890), .B(n14887), .Z(n14889) );
  XNOR U14504 ( .A(n13069), .B(n14883), .Z(n14885) );
  XOR U14505 ( .A(n14891), .B(n14892), .Z(n13069) );
  AND U14506 ( .A(n480), .B(n14893), .Z(n14892) );
  XOR U14507 ( .A(n14894), .B(n14891), .Z(n14893) );
  XOR U14508 ( .A(n14895), .B(n14896), .Z(n14883) );
  AND U14509 ( .A(n14897), .B(n14898), .Z(n14896) );
  XOR U14510 ( .A(n14895), .B(n13084), .Z(n14898) );
  XOR U14511 ( .A(n14899), .B(n14900), .Z(n13084) );
  AND U14512 ( .A(n483), .B(n14901), .Z(n14900) );
  XOR U14513 ( .A(n14902), .B(n14899), .Z(n14901) );
  XNOR U14514 ( .A(n13081), .B(n14895), .Z(n14897) );
  XOR U14515 ( .A(n14903), .B(n14904), .Z(n13081) );
  AND U14516 ( .A(n480), .B(n14905), .Z(n14904) );
  XOR U14517 ( .A(n14906), .B(n14903), .Z(n14905) );
  XOR U14518 ( .A(n14907), .B(n14908), .Z(n14895) );
  AND U14519 ( .A(n14909), .B(n14910), .Z(n14908) );
  XOR U14520 ( .A(n14907), .B(n13096), .Z(n14910) );
  XOR U14521 ( .A(n14911), .B(n14912), .Z(n13096) );
  AND U14522 ( .A(n483), .B(n14913), .Z(n14912) );
  XOR U14523 ( .A(n14914), .B(n14911), .Z(n14913) );
  XNOR U14524 ( .A(n13093), .B(n14907), .Z(n14909) );
  XOR U14525 ( .A(n14915), .B(n14916), .Z(n13093) );
  AND U14526 ( .A(n480), .B(n14917), .Z(n14916) );
  XOR U14527 ( .A(n14918), .B(n14915), .Z(n14917) );
  XOR U14528 ( .A(n14919), .B(n14920), .Z(n14907) );
  AND U14529 ( .A(n14921), .B(n14922), .Z(n14920) );
  XOR U14530 ( .A(n14919), .B(n13108), .Z(n14922) );
  XOR U14531 ( .A(n14923), .B(n14924), .Z(n13108) );
  AND U14532 ( .A(n483), .B(n14925), .Z(n14924) );
  XOR U14533 ( .A(n14926), .B(n14923), .Z(n14925) );
  XNOR U14534 ( .A(n13105), .B(n14919), .Z(n14921) );
  XOR U14535 ( .A(n14927), .B(n14928), .Z(n13105) );
  AND U14536 ( .A(n480), .B(n14929), .Z(n14928) );
  XOR U14537 ( .A(n14930), .B(n14927), .Z(n14929) );
  XOR U14538 ( .A(n14931), .B(n14932), .Z(n14919) );
  AND U14539 ( .A(n14933), .B(n14934), .Z(n14932) );
  XOR U14540 ( .A(n14931), .B(n13120), .Z(n14934) );
  XOR U14541 ( .A(n14935), .B(n14936), .Z(n13120) );
  AND U14542 ( .A(n483), .B(n14937), .Z(n14936) );
  XOR U14543 ( .A(n14938), .B(n14935), .Z(n14937) );
  XNOR U14544 ( .A(n13117), .B(n14931), .Z(n14933) );
  XOR U14545 ( .A(n14939), .B(n14940), .Z(n13117) );
  AND U14546 ( .A(n480), .B(n14941), .Z(n14940) );
  XOR U14547 ( .A(n14942), .B(n14939), .Z(n14941) );
  XOR U14548 ( .A(n14943), .B(n14944), .Z(n14931) );
  AND U14549 ( .A(n14945), .B(n14946), .Z(n14944) );
  XOR U14550 ( .A(n14943), .B(n13132), .Z(n14946) );
  XOR U14551 ( .A(n14947), .B(n14948), .Z(n13132) );
  AND U14552 ( .A(n483), .B(n14949), .Z(n14948) );
  XOR U14553 ( .A(n14950), .B(n14947), .Z(n14949) );
  XNOR U14554 ( .A(n13129), .B(n14943), .Z(n14945) );
  XOR U14555 ( .A(n14951), .B(n14952), .Z(n13129) );
  AND U14556 ( .A(n480), .B(n14953), .Z(n14952) );
  XOR U14557 ( .A(n14954), .B(n14951), .Z(n14953) );
  XOR U14558 ( .A(n14955), .B(n14956), .Z(n14943) );
  AND U14559 ( .A(n14957), .B(n14958), .Z(n14956) );
  XOR U14560 ( .A(n14955), .B(n13144), .Z(n14958) );
  XOR U14561 ( .A(n14959), .B(n14960), .Z(n13144) );
  AND U14562 ( .A(n483), .B(n14961), .Z(n14960) );
  XOR U14563 ( .A(n14962), .B(n14959), .Z(n14961) );
  XNOR U14564 ( .A(n13141), .B(n14955), .Z(n14957) );
  XOR U14565 ( .A(n14963), .B(n14964), .Z(n13141) );
  AND U14566 ( .A(n480), .B(n14965), .Z(n14964) );
  XOR U14567 ( .A(n14966), .B(n14963), .Z(n14965) );
  XOR U14568 ( .A(n14967), .B(n14968), .Z(n14955) );
  AND U14569 ( .A(n14969), .B(n14970), .Z(n14968) );
  XOR U14570 ( .A(n14967), .B(n13156), .Z(n14970) );
  XOR U14571 ( .A(n14971), .B(n14972), .Z(n13156) );
  AND U14572 ( .A(n483), .B(n14973), .Z(n14972) );
  XOR U14573 ( .A(n14974), .B(n14971), .Z(n14973) );
  XNOR U14574 ( .A(n13153), .B(n14967), .Z(n14969) );
  XOR U14575 ( .A(n14975), .B(n14976), .Z(n13153) );
  AND U14576 ( .A(n480), .B(n14977), .Z(n14976) );
  XOR U14577 ( .A(n14978), .B(n14975), .Z(n14977) );
  XOR U14578 ( .A(n14979), .B(n14980), .Z(n14967) );
  AND U14579 ( .A(n14981), .B(n14982), .Z(n14980) );
  XOR U14580 ( .A(n14979), .B(n13168), .Z(n14982) );
  XOR U14581 ( .A(n14983), .B(n14984), .Z(n13168) );
  AND U14582 ( .A(n483), .B(n14985), .Z(n14984) );
  XOR U14583 ( .A(n14986), .B(n14983), .Z(n14985) );
  XNOR U14584 ( .A(n13165), .B(n14979), .Z(n14981) );
  XOR U14585 ( .A(n14987), .B(n14988), .Z(n13165) );
  AND U14586 ( .A(n480), .B(n14989), .Z(n14988) );
  XOR U14587 ( .A(n14990), .B(n14987), .Z(n14989) );
  XOR U14588 ( .A(n14991), .B(n14992), .Z(n14979) );
  AND U14589 ( .A(n14993), .B(n14994), .Z(n14992) );
  XOR U14590 ( .A(n14991), .B(n13180), .Z(n14994) );
  XOR U14591 ( .A(n14995), .B(n14996), .Z(n13180) );
  AND U14592 ( .A(n483), .B(n14997), .Z(n14996) );
  XOR U14593 ( .A(n14998), .B(n14995), .Z(n14997) );
  XNOR U14594 ( .A(n13177), .B(n14991), .Z(n14993) );
  XOR U14595 ( .A(n14999), .B(n15000), .Z(n13177) );
  AND U14596 ( .A(n480), .B(n15001), .Z(n15000) );
  XOR U14597 ( .A(n15002), .B(n14999), .Z(n15001) );
  XOR U14598 ( .A(n15003), .B(n15004), .Z(n14991) );
  AND U14599 ( .A(n15005), .B(n15006), .Z(n15004) );
  XOR U14600 ( .A(n15003), .B(n13192), .Z(n15006) );
  XOR U14601 ( .A(n15007), .B(n15008), .Z(n13192) );
  AND U14602 ( .A(n483), .B(n15009), .Z(n15008) );
  XOR U14603 ( .A(n15010), .B(n15007), .Z(n15009) );
  XNOR U14604 ( .A(n13189), .B(n15003), .Z(n15005) );
  XOR U14605 ( .A(n15011), .B(n15012), .Z(n13189) );
  AND U14606 ( .A(n480), .B(n15013), .Z(n15012) );
  XOR U14607 ( .A(n15014), .B(n15011), .Z(n15013) );
  XOR U14608 ( .A(n15015), .B(n15016), .Z(n15003) );
  AND U14609 ( .A(n15017), .B(n15018), .Z(n15016) );
  XNOR U14610 ( .A(n15019), .B(n13205), .Z(n15018) );
  XOR U14611 ( .A(n15020), .B(n15021), .Z(n13205) );
  AND U14612 ( .A(n483), .B(n15022), .Z(n15021) );
  XOR U14613 ( .A(n15020), .B(n15023), .Z(n15022) );
  XNOR U14614 ( .A(n13202), .B(n15015), .Z(n15017) );
  XOR U14615 ( .A(n15024), .B(n15025), .Z(n13202) );
  AND U14616 ( .A(n480), .B(n15026), .Z(n15025) );
  XOR U14617 ( .A(n15024), .B(n15027), .Z(n15026) );
  IV U14618 ( .A(n15019), .Z(n15015) );
  AND U14619 ( .A(n14651), .B(n14654), .Z(n15019) );
  XNOR U14620 ( .A(n15028), .B(n15029), .Z(n14654) );
  AND U14621 ( .A(n483), .B(n15030), .Z(n15029) );
  XNOR U14622 ( .A(n15031), .B(n15028), .Z(n15030) );
  XOR U14623 ( .A(n15032), .B(n15033), .Z(n483) );
  AND U14624 ( .A(n15034), .B(n15035), .Z(n15033) );
  XOR U14625 ( .A(n14662), .B(n15032), .Z(n15035) );
  IV U14626 ( .A(n15036), .Z(n14662) );
  AND U14627 ( .A(p_input[6399]), .B(p_input[6367]), .Z(n15036) );
  XOR U14628 ( .A(n15032), .B(n14659), .Z(n15034) );
  AND U14629 ( .A(p_input[6303]), .B(p_input[6335]), .Z(n14659) );
  XOR U14630 ( .A(n15037), .B(n15038), .Z(n15032) );
  AND U14631 ( .A(n15039), .B(n15040), .Z(n15038) );
  XOR U14632 ( .A(n15037), .B(n14674), .Z(n15040) );
  XNOR U14633 ( .A(p_input[6366]), .B(n15041), .Z(n14674) );
  AND U14634 ( .A(n287), .B(n15042), .Z(n15041) );
  XOR U14635 ( .A(p_input[6398]), .B(p_input[6366]), .Z(n15042) );
  XNOR U14636 ( .A(n14671), .B(n15037), .Z(n15039) );
  XOR U14637 ( .A(n15043), .B(n15044), .Z(n14671) );
  AND U14638 ( .A(n285), .B(n15045), .Z(n15044) );
  XOR U14639 ( .A(p_input[6334]), .B(p_input[6302]), .Z(n15045) );
  XOR U14640 ( .A(n15046), .B(n15047), .Z(n15037) );
  AND U14641 ( .A(n15048), .B(n15049), .Z(n15047) );
  XOR U14642 ( .A(n15046), .B(n14686), .Z(n15049) );
  XNOR U14643 ( .A(p_input[6365]), .B(n15050), .Z(n14686) );
  AND U14644 ( .A(n287), .B(n15051), .Z(n15050) );
  XOR U14645 ( .A(p_input[6397]), .B(p_input[6365]), .Z(n15051) );
  XNOR U14646 ( .A(n14683), .B(n15046), .Z(n15048) );
  XOR U14647 ( .A(n15052), .B(n15053), .Z(n14683) );
  AND U14648 ( .A(n285), .B(n15054), .Z(n15053) );
  XOR U14649 ( .A(p_input[6333]), .B(p_input[6301]), .Z(n15054) );
  XOR U14650 ( .A(n15055), .B(n15056), .Z(n15046) );
  AND U14651 ( .A(n15057), .B(n15058), .Z(n15056) );
  XOR U14652 ( .A(n15055), .B(n14698), .Z(n15058) );
  XNOR U14653 ( .A(p_input[6364]), .B(n15059), .Z(n14698) );
  AND U14654 ( .A(n287), .B(n15060), .Z(n15059) );
  XOR U14655 ( .A(p_input[6396]), .B(p_input[6364]), .Z(n15060) );
  XNOR U14656 ( .A(n14695), .B(n15055), .Z(n15057) );
  XOR U14657 ( .A(n15061), .B(n15062), .Z(n14695) );
  AND U14658 ( .A(n285), .B(n15063), .Z(n15062) );
  XOR U14659 ( .A(p_input[6332]), .B(p_input[6300]), .Z(n15063) );
  XOR U14660 ( .A(n15064), .B(n15065), .Z(n15055) );
  AND U14661 ( .A(n15066), .B(n15067), .Z(n15065) );
  XOR U14662 ( .A(n15064), .B(n14710), .Z(n15067) );
  XNOR U14663 ( .A(p_input[6363]), .B(n15068), .Z(n14710) );
  AND U14664 ( .A(n287), .B(n15069), .Z(n15068) );
  XOR U14665 ( .A(p_input[6395]), .B(p_input[6363]), .Z(n15069) );
  XNOR U14666 ( .A(n14707), .B(n15064), .Z(n15066) );
  XOR U14667 ( .A(n15070), .B(n15071), .Z(n14707) );
  AND U14668 ( .A(n285), .B(n15072), .Z(n15071) );
  XOR U14669 ( .A(p_input[6331]), .B(p_input[6299]), .Z(n15072) );
  XOR U14670 ( .A(n15073), .B(n15074), .Z(n15064) );
  AND U14671 ( .A(n15075), .B(n15076), .Z(n15074) );
  XOR U14672 ( .A(n15073), .B(n14722), .Z(n15076) );
  XNOR U14673 ( .A(p_input[6362]), .B(n15077), .Z(n14722) );
  AND U14674 ( .A(n287), .B(n15078), .Z(n15077) );
  XOR U14675 ( .A(p_input[6394]), .B(p_input[6362]), .Z(n15078) );
  XNOR U14676 ( .A(n14719), .B(n15073), .Z(n15075) );
  XOR U14677 ( .A(n15079), .B(n15080), .Z(n14719) );
  AND U14678 ( .A(n285), .B(n15081), .Z(n15080) );
  XOR U14679 ( .A(p_input[6330]), .B(p_input[6298]), .Z(n15081) );
  XOR U14680 ( .A(n15082), .B(n15083), .Z(n15073) );
  AND U14681 ( .A(n15084), .B(n15085), .Z(n15083) );
  XOR U14682 ( .A(n15082), .B(n14734), .Z(n15085) );
  XNOR U14683 ( .A(p_input[6361]), .B(n15086), .Z(n14734) );
  AND U14684 ( .A(n287), .B(n15087), .Z(n15086) );
  XOR U14685 ( .A(p_input[6393]), .B(p_input[6361]), .Z(n15087) );
  XNOR U14686 ( .A(n14731), .B(n15082), .Z(n15084) );
  XOR U14687 ( .A(n15088), .B(n15089), .Z(n14731) );
  AND U14688 ( .A(n285), .B(n15090), .Z(n15089) );
  XOR U14689 ( .A(p_input[6329]), .B(p_input[6297]), .Z(n15090) );
  XOR U14690 ( .A(n15091), .B(n15092), .Z(n15082) );
  AND U14691 ( .A(n15093), .B(n15094), .Z(n15092) );
  XOR U14692 ( .A(n15091), .B(n14746), .Z(n15094) );
  XNOR U14693 ( .A(p_input[6360]), .B(n15095), .Z(n14746) );
  AND U14694 ( .A(n287), .B(n15096), .Z(n15095) );
  XOR U14695 ( .A(p_input[6392]), .B(p_input[6360]), .Z(n15096) );
  XNOR U14696 ( .A(n14743), .B(n15091), .Z(n15093) );
  XOR U14697 ( .A(n15097), .B(n15098), .Z(n14743) );
  AND U14698 ( .A(n285), .B(n15099), .Z(n15098) );
  XOR U14699 ( .A(p_input[6328]), .B(p_input[6296]), .Z(n15099) );
  XOR U14700 ( .A(n15100), .B(n15101), .Z(n15091) );
  AND U14701 ( .A(n15102), .B(n15103), .Z(n15101) );
  XOR U14702 ( .A(n15100), .B(n14758), .Z(n15103) );
  XNOR U14703 ( .A(p_input[6359]), .B(n15104), .Z(n14758) );
  AND U14704 ( .A(n287), .B(n15105), .Z(n15104) );
  XOR U14705 ( .A(p_input[6391]), .B(p_input[6359]), .Z(n15105) );
  XNOR U14706 ( .A(n14755), .B(n15100), .Z(n15102) );
  XOR U14707 ( .A(n15106), .B(n15107), .Z(n14755) );
  AND U14708 ( .A(n285), .B(n15108), .Z(n15107) );
  XOR U14709 ( .A(p_input[6327]), .B(p_input[6295]), .Z(n15108) );
  XOR U14710 ( .A(n15109), .B(n15110), .Z(n15100) );
  AND U14711 ( .A(n15111), .B(n15112), .Z(n15110) );
  XOR U14712 ( .A(n15109), .B(n14770), .Z(n15112) );
  XNOR U14713 ( .A(p_input[6358]), .B(n15113), .Z(n14770) );
  AND U14714 ( .A(n287), .B(n15114), .Z(n15113) );
  XOR U14715 ( .A(p_input[6390]), .B(p_input[6358]), .Z(n15114) );
  XNOR U14716 ( .A(n14767), .B(n15109), .Z(n15111) );
  XOR U14717 ( .A(n15115), .B(n15116), .Z(n14767) );
  AND U14718 ( .A(n285), .B(n15117), .Z(n15116) );
  XOR U14719 ( .A(p_input[6326]), .B(p_input[6294]), .Z(n15117) );
  XOR U14720 ( .A(n15118), .B(n15119), .Z(n15109) );
  AND U14721 ( .A(n15120), .B(n15121), .Z(n15119) );
  XOR U14722 ( .A(n15118), .B(n14782), .Z(n15121) );
  XNOR U14723 ( .A(p_input[6357]), .B(n15122), .Z(n14782) );
  AND U14724 ( .A(n287), .B(n15123), .Z(n15122) );
  XOR U14725 ( .A(p_input[6389]), .B(p_input[6357]), .Z(n15123) );
  XNOR U14726 ( .A(n14779), .B(n15118), .Z(n15120) );
  XOR U14727 ( .A(n15124), .B(n15125), .Z(n14779) );
  AND U14728 ( .A(n285), .B(n15126), .Z(n15125) );
  XOR U14729 ( .A(p_input[6325]), .B(p_input[6293]), .Z(n15126) );
  XOR U14730 ( .A(n15127), .B(n15128), .Z(n15118) );
  AND U14731 ( .A(n15129), .B(n15130), .Z(n15128) );
  XOR U14732 ( .A(n15127), .B(n14794), .Z(n15130) );
  XNOR U14733 ( .A(p_input[6356]), .B(n15131), .Z(n14794) );
  AND U14734 ( .A(n287), .B(n15132), .Z(n15131) );
  XOR U14735 ( .A(p_input[6388]), .B(p_input[6356]), .Z(n15132) );
  XNOR U14736 ( .A(n14791), .B(n15127), .Z(n15129) );
  XOR U14737 ( .A(n15133), .B(n15134), .Z(n14791) );
  AND U14738 ( .A(n285), .B(n15135), .Z(n15134) );
  XOR U14739 ( .A(p_input[6324]), .B(p_input[6292]), .Z(n15135) );
  XOR U14740 ( .A(n15136), .B(n15137), .Z(n15127) );
  AND U14741 ( .A(n15138), .B(n15139), .Z(n15137) );
  XOR U14742 ( .A(n15136), .B(n14806), .Z(n15139) );
  XNOR U14743 ( .A(p_input[6355]), .B(n15140), .Z(n14806) );
  AND U14744 ( .A(n287), .B(n15141), .Z(n15140) );
  XOR U14745 ( .A(p_input[6387]), .B(p_input[6355]), .Z(n15141) );
  XNOR U14746 ( .A(n14803), .B(n15136), .Z(n15138) );
  XOR U14747 ( .A(n15142), .B(n15143), .Z(n14803) );
  AND U14748 ( .A(n285), .B(n15144), .Z(n15143) );
  XOR U14749 ( .A(p_input[6323]), .B(p_input[6291]), .Z(n15144) );
  XOR U14750 ( .A(n15145), .B(n15146), .Z(n15136) );
  AND U14751 ( .A(n15147), .B(n15148), .Z(n15146) );
  XOR U14752 ( .A(n15145), .B(n14818), .Z(n15148) );
  XNOR U14753 ( .A(p_input[6354]), .B(n15149), .Z(n14818) );
  AND U14754 ( .A(n287), .B(n15150), .Z(n15149) );
  XOR U14755 ( .A(p_input[6386]), .B(p_input[6354]), .Z(n15150) );
  XNOR U14756 ( .A(n14815), .B(n15145), .Z(n15147) );
  XOR U14757 ( .A(n15151), .B(n15152), .Z(n14815) );
  AND U14758 ( .A(n285), .B(n15153), .Z(n15152) );
  XOR U14759 ( .A(p_input[6322]), .B(p_input[6290]), .Z(n15153) );
  XOR U14760 ( .A(n15154), .B(n15155), .Z(n15145) );
  AND U14761 ( .A(n15156), .B(n15157), .Z(n15155) );
  XOR U14762 ( .A(n15154), .B(n14830), .Z(n15157) );
  XNOR U14763 ( .A(p_input[6353]), .B(n15158), .Z(n14830) );
  AND U14764 ( .A(n287), .B(n15159), .Z(n15158) );
  XOR U14765 ( .A(p_input[6385]), .B(p_input[6353]), .Z(n15159) );
  XNOR U14766 ( .A(n14827), .B(n15154), .Z(n15156) );
  XOR U14767 ( .A(n15160), .B(n15161), .Z(n14827) );
  AND U14768 ( .A(n285), .B(n15162), .Z(n15161) );
  XOR U14769 ( .A(p_input[6321]), .B(p_input[6289]), .Z(n15162) );
  XOR U14770 ( .A(n15163), .B(n15164), .Z(n15154) );
  AND U14771 ( .A(n15165), .B(n15166), .Z(n15164) );
  XOR U14772 ( .A(n15163), .B(n14842), .Z(n15166) );
  XNOR U14773 ( .A(p_input[6352]), .B(n15167), .Z(n14842) );
  AND U14774 ( .A(n287), .B(n15168), .Z(n15167) );
  XOR U14775 ( .A(p_input[6384]), .B(p_input[6352]), .Z(n15168) );
  XNOR U14776 ( .A(n14839), .B(n15163), .Z(n15165) );
  XOR U14777 ( .A(n15169), .B(n15170), .Z(n14839) );
  AND U14778 ( .A(n285), .B(n15171), .Z(n15170) );
  XOR U14779 ( .A(p_input[6320]), .B(p_input[6288]), .Z(n15171) );
  XOR U14780 ( .A(n15172), .B(n15173), .Z(n15163) );
  AND U14781 ( .A(n15174), .B(n15175), .Z(n15173) );
  XOR U14782 ( .A(n15172), .B(n14854), .Z(n15175) );
  XNOR U14783 ( .A(p_input[6351]), .B(n15176), .Z(n14854) );
  AND U14784 ( .A(n287), .B(n15177), .Z(n15176) );
  XOR U14785 ( .A(p_input[6383]), .B(p_input[6351]), .Z(n15177) );
  XNOR U14786 ( .A(n14851), .B(n15172), .Z(n15174) );
  XOR U14787 ( .A(n15178), .B(n15179), .Z(n14851) );
  AND U14788 ( .A(n285), .B(n15180), .Z(n15179) );
  XOR U14789 ( .A(p_input[6319]), .B(p_input[6287]), .Z(n15180) );
  XOR U14790 ( .A(n15181), .B(n15182), .Z(n15172) );
  AND U14791 ( .A(n15183), .B(n15184), .Z(n15182) );
  XOR U14792 ( .A(n15181), .B(n14866), .Z(n15184) );
  XNOR U14793 ( .A(p_input[6350]), .B(n15185), .Z(n14866) );
  AND U14794 ( .A(n287), .B(n15186), .Z(n15185) );
  XOR U14795 ( .A(p_input[6382]), .B(p_input[6350]), .Z(n15186) );
  XNOR U14796 ( .A(n14863), .B(n15181), .Z(n15183) );
  XOR U14797 ( .A(n15187), .B(n15188), .Z(n14863) );
  AND U14798 ( .A(n285), .B(n15189), .Z(n15188) );
  XOR U14799 ( .A(p_input[6318]), .B(p_input[6286]), .Z(n15189) );
  XOR U14800 ( .A(n15190), .B(n15191), .Z(n15181) );
  AND U14801 ( .A(n15192), .B(n15193), .Z(n15191) );
  XOR U14802 ( .A(n15190), .B(n14878), .Z(n15193) );
  XNOR U14803 ( .A(p_input[6349]), .B(n15194), .Z(n14878) );
  AND U14804 ( .A(n287), .B(n15195), .Z(n15194) );
  XOR U14805 ( .A(p_input[6381]), .B(p_input[6349]), .Z(n15195) );
  XNOR U14806 ( .A(n14875), .B(n15190), .Z(n15192) );
  XOR U14807 ( .A(n15196), .B(n15197), .Z(n14875) );
  AND U14808 ( .A(n285), .B(n15198), .Z(n15197) );
  XOR U14809 ( .A(p_input[6317]), .B(p_input[6285]), .Z(n15198) );
  XOR U14810 ( .A(n15199), .B(n15200), .Z(n15190) );
  AND U14811 ( .A(n15201), .B(n15202), .Z(n15200) );
  XOR U14812 ( .A(n15199), .B(n14890), .Z(n15202) );
  XNOR U14813 ( .A(p_input[6348]), .B(n15203), .Z(n14890) );
  AND U14814 ( .A(n287), .B(n15204), .Z(n15203) );
  XOR U14815 ( .A(p_input[6380]), .B(p_input[6348]), .Z(n15204) );
  XNOR U14816 ( .A(n14887), .B(n15199), .Z(n15201) );
  XOR U14817 ( .A(n15205), .B(n15206), .Z(n14887) );
  AND U14818 ( .A(n285), .B(n15207), .Z(n15206) );
  XOR U14819 ( .A(p_input[6316]), .B(p_input[6284]), .Z(n15207) );
  XOR U14820 ( .A(n15208), .B(n15209), .Z(n15199) );
  AND U14821 ( .A(n15210), .B(n15211), .Z(n15209) );
  XOR U14822 ( .A(n15208), .B(n14902), .Z(n15211) );
  XNOR U14823 ( .A(p_input[6347]), .B(n15212), .Z(n14902) );
  AND U14824 ( .A(n287), .B(n15213), .Z(n15212) );
  XOR U14825 ( .A(p_input[6379]), .B(p_input[6347]), .Z(n15213) );
  XNOR U14826 ( .A(n14899), .B(n15208), .Z(n15210) );
  XOR U14827 ( .A(n15214), .B(n15215), .Z(n14899) );
  AND U14828 ( .A(n285), .B(n15216), .Z(n15215) );
  XOR U14829 ( .A(p_input[6315]), .B(p_input[6283]), .Z(n15216) );
  XOR U14830 ( .A(n15217), .B(n15218), .Z(n15208) );
  AND U14831 ( .A(n15219), .B(n15220), .Z(n15218) );
  XOR U14832 ( .A(n15217), .B(n14914), .Z(n15220) );
  XNOR U14833 ( .A(p_input[6346]), .B(n15221), .Z(n14914) );
  AND U14834 ( .A(n287), .B(n15222), .Z(n15221) );
  XOR U14835 ( .A(p_input[6378]), .B(p_input[6346]), .Z(n15222) );
  XNOR U14836 ( .A(n14911), .B(n15217), .Z(n15219) );
  XOR U14837 ( .A(n15223), .B(n15224), .Z(n14911) );
  AND U14838 ( .A(n285), .B(n15225), .Z(n15224) );
  XOR U14839 ( .A(p_input[6314]), .B(p_input[6282]), .Z(n15225) );
  XOR U14840 ( .A(n15226), .B(n15227), .Z(n15217) );
  AND U14841 ( .A(n15228), .B(n15229), .Z(n15227) );
  XOR U14842 ( .A(n15226), .B(n14926), .Z(n15229) );
  XNOR U14843 ( .A(p_input[6345]), .B(n15230), .Z(n14926) );
  AND U14844 ( .A(n287), .B(n15231), .Z(n15230) );
  XOR U14845 ( .A(p_input[6377]), .B(p_input[6345]), .Z(n15231) );
  XNOR U14846 ( .A(n14923), .B(n15226), .Z(n15228) );
  XOR U14847 ( .A(n15232), .B(n15233), .Z(n14923) );
  AND U14848 ( .A(n285), .B(n15234), .Z(n15233) );
  XOR U14849 ( .A(p_input[6313]), .B(p_input[6281]), .Z(n15234) );
  XOR U14850 ( .A(n15235), .B(n15236), .Z(n15226) );
  AND U14851 ( .A(n15237), .B(n15238), .Z(n15236) );
  XOR U14852 ( .A(n15235), .B(n14938), .Z(n15238) );
  XNOR U14853 ( .A(p_input[6344]), .B(n15239), .Z(n14938) );
  AND U14854 ( .A(n287), .B(n15240), .Z(n15239) );
  XOR U14855 ( .A(p_input[6376]), .B(p_input[6344]), .Z(n15240) );
  XNOR U14856 ( .A(n14935), .B(n15235), .Z(n15237) );
  XOR U14857 ( .A(n15241), .B(n15242), .Z(n14935) );
  AND U14858 ( .A(n285), .B(n15243), .Z(n15242) );
  XOR U14859 ( .A(p_input[6312]), .B(p_input[6280]), .Z(n15243) );
  XOR U14860 ( .A(n15244), .B(n15245), .Z(n15235) );
  AND U14861 ( .A(n15246), .B(n15247), .Z(n15245) );
  XOR U14862 ( .A(n15244), .B(n14950), .Z(n15247) );
  XNOR U14863 ( .A(p_input[6343]), .B(n15248), .Z(n14950) );
  AND U14864 ( .A(n287), .B(n15249), .Z(n15248) );
  XOR U14865 ( .A(p_input[6375]), .B(p_input[6343]), .Z(n15249) );
  XNOR U14866 ( .A(n14947), .B(n15244), .Z(n15246) );
  XOR U14867 ( .A(n15250), .B(n15251), .Z(n14947) );
  AND U14868 ( .A(n285), .B(n15252), .Z(n15251) );
  XOR U14869 ( .A(p_input[6311]), .B(p_input[6279]), .Z(n15252) );
  XOR U14870 ( .A(n15253), .B(n15254), .Z(n15244) );
  AND U14871 ( .A(n15255), .B(n15256), .Z(n15254) );
  XOR U14872 ( .A(n15253), .B(n14962), .Z(n15256) );
  XNOR U14873 ( .A(p_input[6342]), .B(n15257), .Z(n14962) );
  AND U14874 ( .A(n287), .B(n15258), .Z(n15257) );
  XOR U14875 ( .A(p_input[6374]), .B(p_input[6342]), .Z(n15258) );
  XNOR U14876 ( .A(n14959), .B(n15253), .Z(n15255) );
  XOR U14877 ( .A(n15259), .B(n15260), .Z(n14959) );
  AND U14878 ( .A(n285), .B(n15261), .Z(n15260) );
  XOR U14879 ( .A(p_input[6310]), .B(p_input[6278]), .Z(n15261) );
  XOR U14880 ( .A(n15262), .B(n15263), .Z(n15253) );
  AND U14881 ( .A(n15264), .B(n15265), .Z(n15263) );
  XOR U14882 ( .A(n15262), .B(n14974), .Z(n15265) );
  XNOR U14883 ( .A(p_input[6341]), .B(n15266), .Z(n14974) );
  AND U14884 ( .A(n287), .B(n15267), .Z(n15266) );
  XOR U14885 ( .A(p_input[6373]), .B(p_input[6341]), .Z(n15267) );
  XNOR U14886 ( .A(n14971), .B(n15262), .Z(n15264) );
  XOR U14887 ( .A(n15268), .B(n15269), .Z(n14971) );
  AND U14888 ( .A(n285), .B(n15270), .Z(n15269) );
  XOR U14889 ( .A(p_input[6309]), .B(p_input[6277]), .Z(n15270) );
  XOR U14890 ( .A(n15271), .B(n15272), .Z(n15262) );
  AND U14891 ( .A(n15273), .B(n15274), .Z(n15272) );
  XOR U14892 ( .A(n15271), .B(n14986), .Z(n15274) );
  XNOR U14893 ( .A(p_input[6340]), .B(n15275), .Z(n14986) );
  AND U14894 ( .A(n287), .B(n15276), .Z(n15275) );
  XOR U14895 ( .A(p_input[6372]), .B(p_input[6340]), .Z(n15276) );
  XNOR U14896 ( .A(n14983), .B(n15271), .Z(n15273) );
  XOR U14897 ( .A(n15277), .B(n15278), .Z(n14983) );
  AND U14898 ( .A(n285), .B(n15279), .Z(n15278) );
  XOR U14899 ( .A(p_input[6308]), .B(p_input[6276]), .Z(n15279) );
  XOR U14900 ( .A(n15280), .B(n15281), .Z(n15271) );
  AND U14901 ( .A(n15282), .B(n15283), .Z(n15281) );
  XOR U14902 ( .A(n15280), .B(n14998), .Z(n15283) );
  XNOR U14903 ( .A(p_input[6339]), .B(n15284), .Z(n14998) );
  AND U14904 ( .A(n287), .B(n15285), .Z(n15284) );
  XOR U14905 ( .A(p_input[6371]), .B(p_input[6339]), .Z(n15285) );
  XNOR U14906 ( .A(n14995), .B(n15280), .Z(n15282) );
  XOR U14907 ( .A(n15286), .B(n15287), .Z(n14995) );
  AND U14908 ( .A(n285), .B(n15288), .Z(n15287) );
  XOR U14909 ( .A(p_input[6307]), .B(p_input[6275]), .Z(n15288) );
  XOR U14910 ( .A(n15289), .B(n15290), .Z(n15280) );
  AND U14911 ( .A(n15291), .B(n15292), .Z(n15290) );
  XOR U14912 ( .A(n15289), .B(n15010), .Z(n15292) );
  XNOR U14913 ( .A(p_input[6338]), .B(n15293), .Z(n15010) );
  AND U14914 ( .A(n287), .B(n15294), .Z(n15293) );
  XOR U14915 ( .A(p_input[6370]), .B(p_input[6338]), .Z(n15294) );
  XNOR U14916 ( .A(n15007), .B(n15289), .Z(n15291) );
  XOR U14917 ( .A(n15295), .B(n15296), .Z(n15007) );
  AND U14918 ( .A(n285), .B(n15297), .Z(n15296) );
  XOR U14919 ( .A(p_input[6306]), .B(p_input[6274]), .Z(n15297) );
  XOR U14920 ( .A(n15298), .B(n15299), .Z(n15289) );
  AND U14921 ( .A(n15300), .B(n15301), .Z(n15299) );
  XNOR U14922 ( .A(n15302), .B(n15023), .Z(n15301) );
  XNOR U14923 ( .A(p_input[6337]), .B(n15303), .Z(n15023) );
  AND U14924 ( .A(n287), .B(n15304), .Z(n15303) );
  XNOR U14925 ( .A(p_input[6369]), .B(n15305), .Z(n15304) );
  IV U14926 ( .A(p_input[6337]), .Z(n15305) );
  XNOR U14927 ( .A(n15020), .B(n15298), .Z(n15300) );
  XNOR U14928 ( .A(p_input[6273]), .B(n15306), .Z(n15020) );
  AND U14929 ( .A(n285), .B(n15307), .Z(n15306) );
  XOR U14930 ( .A(p_input[6305]), .B(p_input[6273]), .Z(n15307) );
  IV U14931 ( .A(n15302), .Z(n15298) );
  AND U14932 ( .A(n15028), .B(n15031), .Z(n15302) );
  XOR U14933 ( .A(p_input[6336]), .B(n15308), .Z(n15031) );
  AND U14934 ( .A(n287), .B(n15309), .Z(n15308) );
  XOR U14935 ( .A(p_input[6368]), .B(p_input[6336]), .Z(n15309) );
  XOR U14936 ( .A(n15310), .B(n15311), .Z(n287) );
  AND U14937 ( .A(n15312), .B(n15313), .Z(n15311) );
  XNOR U14938 ( .A(p_input[6399]), .B(n15310), .Z(n15313) );
  XOR U14939 ( .A(n15310), .B(p_input[6367]), .Z(n15312) );
  XOR U14940 ( .A(n15314), .B(n15315), .Z(n15310) );
  AND U14941 ( .A(n15316), .B(n15317), .Z(n15315) );
  XNOR U14942 ( .A(p_input[6398]), .B(n15314), .Z(n15317) );
  XOR U14943 ( .A(n15314), .B(p_input[6366]), .Z(n15316) );
  XOR U14944 ( .A(n15318), .B(n15319), .Z(n15314) );
  AND U14945 ( .A(n15320), .B(n15321), .Z(n15319) );
  XNOR U14946 ( .A(p_input[6397]), .B(n15318), .Z(n15321) );
  XOR U14947 ( .A(n15318), .B(p_input[6365]), .Z(n15320) );
  XOR U14948 ( .A(n15322), .B(n15323), .Z(n15318) );
  AND U14949 ( .A(n15324), .B(n15325), .Z(n15323) );
  XNOR U14950 ( .A(p_input[6396]), .B(n15322), .Z(n15325) );
  XOR U14951 ( .A(n15322), .B(p_input[6364]), .Z(n15324) );
  XOR U14952 ( .A(n15326), .B(n15327), .Z(n15322) );
  AND U14953 ( .A(n15328), .B(n15329), .Z(n15327) );
  XNOR U14954 ( .A(p_input[6395]), .B(n15326), .Z(n15329) );
  XOR U14955 ( .A(n15326), .B(p_input[6363]), .Z(n15328) );
  XOR U14956 ( .A(n15330), .B(n15331), .Z(n15326) );
  AND U14957 ( .A(n15332), .B(n15333), .Z(n15331) );
  XNOR U14958 ( .A(p_input[6394]), .B(n15330), .Z(n15333) );
  XOR U14959 ( .A(n15330), .B(p_input[6362]), .Z(n15332) );
  XOR U14960 ( .A(n15334), .B(n15335), .Z(n15330) );
  AND U14961 ( .A(n15336), .B(n15337), .Z(n15335) );
  XNOR U14962 ( .A(p_input[6393]), .B(n15334), .Z(n15337) );
  XOR U14963 ( .A(n15334), .B(p_input[6361]), .Z(n15336) );
  XOR U14964 ( .A(n15338), .B(n15339), .Z(n15334) );
  AND U14965 ( .A(n15340), .B(n15341), .Z(n15339) );
  XNOR U14966 ( .A(p_input[6392]), .B(n15338), .Z(n15341) );
  XOR U14967 ( .A(n15338), .B(p_input[6360]), .Z(n15340) );
  XOR U14968 ( .A(n15342), .B(n15343), .Z(n15338) );
  AND U14969 ( .A(n15344), .B(n15345), .Z(n15343) );
  XNOR U14970 ( .A(p_input[6391]), .B(n15342), .Z(n15345) );
  XOR U14971 ( .A(n15342), .B(p_input[6359]), .Z(n15344) );
  XOR U14972 ( .A(n15346), .B(n15347), .Z(n15342) );
  AND U14973 ( .A(n15348), .B(n15349), .Z(n15347) );
  XNOR U14974 ( .A(p_input[6390]), .B(n15346), .Z(n15349) );
  XOR U14975 ( .A(n15346), .B(p_input[6358]), .Z(n15348) );
  XOR U14976 ( .A(n15350), .B(n15351), .Z(n15346) );
  AND U14977 ( .A(n15352), .B(n15353), .Z(n15351) );
  XNOR U14978 ( .A(p_input[6389]), .B(n15350), .Z(n15353) );
  XOR U14979 ( .A(n15350), .B(p_input[6357]), .Z(n15352) );
  XOR U14980 ( .A(n15354), .B(n15355), .Z(n15350) );
  AND U14981 ( .A(n15356), .B(n15357), .Z(n15355) );
  XNOR U14982 ( .A(p_input[6388]), .B(n15354), .Z(n15357) );
  XOR U14983 ( .A(n15354), .B(p_input[6356]), .Z(n15356) );
  XOR U14984 ( .A(n15358), .B(n15359), .Z(n15354) );
  AND U14985 ( .A(n15360), .B(n15361), .Z(n15359) );
  XNOR U14986 ( .A(p_input[6387]), .B(n15358), .Z(n15361) );
  XOR U14987 ( .A(n15358), .B(p_input[6355]), .Z(n15360) );
  XOR U14988 ( .A(n15362), .B(n15363), .Z(n15358) );
  AND U14989 ( .A(n15364), .B(n15365), .Z(n15363) );
  XNOR U14990 ( .A(p_input[6386]), .B(n15362), .Z(n15365) );
  XOR U14991 ( .A(n15362), .B(p_input[6354]), .Z(n15364) );
  XOR U14992 ( .A(n15366), .B(n15367), .Z(n15362) );
  AND U14993 ( .A(n15368), .B(n15369), .Z(n15367) );
  XNOR U14994 ( .A(p_input[6385]), .B(n15366), .Z(n15369) );
  XOR U14995 ( .A(n15366), .B(p_input[6353]), .Z(n15368) );
  XOR U14996 ( .A(n15370), .B(n15371), .Z(n15366) );
  AND U14997 ( .A(n15372), .B(n15373), .Z(n15371) );
  XNOR U14998 ( .A(p_input[6384]), .B(n15370), .Z(n15373) );
  XOR U14999 ( .A(n15370), .B(p_input[6352]), .Z(n15372) );
  XOR U15000 ( .A(n15374), .B(n15375), .Z(n15370) );
  AND U15001 ( .A(n15376), .B(n15377), .Z(n15375) );
  XNOR U15002 ( .A(p_input[6383]), .B(n15374), .Z(n15377) );
  XOR U15003 ( .A(n15374), .B(p_input[6351]), .Z(n15376) );
  XOR U15004 ( .A(n15378), .B(n15379), .Z(n15374) );
  AND U15005 ( .A(n15380), .B(n15381), .Z(n15379) );
  XNOR U15006 ( .A(p_input[6382]), .B(n15378), .Z(n15381) );
  XOR U15007 ( .A(n15378), .B(p_input[6350]), .Z(n15380) );
  XOR U15008 ( .A(n15382), .B(n15383), .Z(n15378) );
  AND U15009 ( .A(n15384), .B(n15385), .Z(n15383) );
  XNOR U15010 ( .A(p_input[6381]), .B(n15382), .Z(n15385) );
  XOR U15011 ( .A(n15382), .B(p_input[6349]), .Z(n15384) );
  XOR U15012 ( .A(n15386), .B(n15387), .Z(n15382) );
  AND U15013 ( .A(n15388), .B(n15389), .Z(n15387) );
  XNOR U15014 ( .A(p_input[6380]), .B(n15386), .Z(n15389) );
  XOR U15015 ( .A(n15386), .B(p_input[6348]), .Z(n15388) );
  XOR U15016 ( .A(n15390), .B(n15391), .Z(n15386) );
  AND U15017 ( .A(n15392), .B(n15393), .Z(n15391) );
  XNOR U15018 ( .A(p_input[6379]), .B(n15390), .Z(n15393) );
  XOR U15019 ( .A(n15390), .B(p_input[6347]), .Z(n15392) );
  XOR U15020 ( .A(n15394), .B(n15395), .Z(n15390) );
  AND U15021 ( .A(n15396), .B(n15397), .Z(n15395) );
  XNOR U15022 ( .A(p_input[6378]), .B(n15394), .Z(n15397) );
  XOR U15023 ( .A(n15394), .B(p_input[6346]), .Z(n15396) );
  XOR U15024 ( .A(n15398), .B(n15399), .Z(n15394) );
  AND U15025 ( .A(n15400), .B(n15401), .Z(n15399) );
  XNOR U15026 ( .A(p_input[6377]), .B(n15398), .Z(n15401) );
  XOR U15027 ( .A(n15398), .B(p_input[6345]), .Z(n15400) );
  XOR U15028 ( .A(n15402), .B(n15403), .Z(n15398) );
  AND U15029 ( .A(n15404), .B(n15405), .Z(n15403) );
  XNOR U15030 ( .A(p_input[6376]), .B(n15402), .Z(n15405) );
  XOR U15031 ( .A(n15402), .B(p_input[6344]), .Z(n15404) );
  XOR U15032 ( .A(n15406), .B(n15407), .Z(n15402) );
  AND U15033 ( .A(n15408), .B(n15409), .Z(n15407) );
  XNOR U15034 ( .A(p_input[6375]), .B(n15406), .Z(n15409) );
  XOR U15035 ( .A(n15406), .B(p_input[6343]), .Z(n15408) );
  XOR U15036 ( .A(n15410), .B(n15411), .Z(n15406) );
  AND U15037 ( .A(n15412), .B(n15413), .Z(n15411) );
  XNOR U15038 ( .A(p_input[6374]), .B(n15410), .Z(n15413) );
  XOR U15039 ( .A(n15410), .B(p_input[6342]), .Z(n15412) );
  XOR U15040 ( .A(n15414), .B(n15415), .Z(n15410) );
  AND U15041 ( .A(n15416), .B(n15417), .Z(n15415) );
  XNOR U15042 ( .A(p_input[6373]), .B(n15414), .Z(n15417) );
  XOR U15043 ( .A(n15414), .B(p_input[6341]), .Z(n15416) );
  XOR U15044 ( .A(n15418), .B(n15419), .Z(n15414) );
  AND U15045 ( .A(n15420), .B(n15421), .Z(n15419) );
  XNOR U15046 ( .A(p_input[6372]), .B(n15418), .Z(n15421) );
  XOR U15047 ( .A(n15418), .B(p_input[6340]), .Z(n15420) );
  XOR U15048 ( .A(n15422), .B(n15423), .Z(n15418) );
  AND U15049 ( .A(n15424), .B(n15425), .Z(n15423) );
  XNOR U15050 ( .A(p_input[6371]), .B(n15422), .Z(n15425) );
  XOR U15051 ( .A(n15422), .B(p_input[6339]), .Z(n15424) );
  XOR U15052 ( .A(n15426), .B(n15427), .Z(n15422) );
  AND U15053 ( .A(n15428), .B(n15429), .Z(n15427) );
  XNOR U15054 ( .A(p_input[6370]), .B(n15426), .Z(n15429) );
  XOR U15055 ( .A(n15426), .B(p_input[6338]), .Z(n15428) );
  XNOR U15056 ( .A(n15430), .B(n15431), .Z(n15426) );
  AND U15057 ( .A(n15432), .B(n15433), .Z(n15431) );
  XOR U15058 ( .A(p_input[6369]), .B(n15430), .Z(n15433) );
  XNOR U15059 ( .A(p_input[6337]), .B(n15430), .Z(n15432) );
  AND U15060 ( .A(p_input[6368]), .B(n15434), .Z(n15430) );
  IV U15061 ( .A(p_input[6336]), .Z(n15434) );
  XNOR U15062 ( .A(p_input[6272]), .B(n15435), .Z(n15028) );
  AND U15063 ( .A(n285), .B(n15436), .Z(n15435) );
  XOR U15064 ( .A(p_input[6304]), .B(p_input[6272]), .Z(n15436) );
  XOR U15065 ( .A(n15437), .B(n15438), .Z(n285) );
  AND U15066 ( .A(n15439), .B(n15440), .Z(n15438) );
  XNOR U15067 ( .A(p_input[6335]), .B(n15437), .Z(n15440) );
  XOR U15068 ( .A(n15437), .B(p_input[6303]), .Z(n15439) );
  XOR U15069 ( .A(n15441), .B(n15442), .Z(n15437) );
  AND U15070 ( .A(n15443), .B(n15444), .Z(n15442) );
  XNOR U15071 ( .A(p_input[6334]), .B(n15441), .Z(n15444) );
  XNOR U15072 ( .A(n15441), .B(n15043), .Z(n15443) );
  IV U15073 ( .A(p_input[6302]), .Z(n15043) );
  XOR U15074 ( .A(n15445), .B(n15446), .Z(n15441) );
  AND U15075 ( .A(n15447), .B(n15448), .Z(n15446) );
  XNOR U15076 ( .A(p_input[6333]), .B(n15445), .Z(n15448) );
  XNOR U15077 ( .A(n15445), .B(n15052), .Z(n15447) );
  IV U15078 ( .A(p_input[6301]), .Z(n15052) );
  XOR U15079 ( .A(n15449), .B(n15450), .Z(n15445) );
  AND U15080 ( .A(n15451), .B(n15452), .Z(n15450) );
  XNOR U15081 ( .A(p_input[6332]), .B(n15449), .Z(n15452) );
  XNOR U15082 ( .A(n15449), .B(n15061), .Z(n15451) );
  IV U15083 ( .A(p_input[6300]), .Z(n15061) );
  XOR U15084 ( .A(n15453), .B(n15454), .Z(n15449) );
  AND U15085 ( .A(n15455), .B(n15456), .Z(n15454) );
  XNOR U15086 ( .A(p_input[6331]), .B(n15453), .Z(n15456) );
  XNOR U15087 ( .A(n15453), .B(n15070), .Z(n15455) );
  IV U15088 ( .A(p_input[6299]), .Z(n15070) );
  XOR U15089 ( .A(n15457), .B(n15458), .Z(n15453) );
  AND U15090 ( .A(n15459), .B(n15460), .Z(n15458) );
  XNOR U15091 ( .A(p_input[6330]), .B(n15457), .Z(n15460) );
  XNOR U15092 ( .A(n15457), .B(n15079), .Z(n15459) );
  IV U15093 ( .A(p_input[6298]), .Z(n15079) );
  XOR U15094 ( .A(n15461), .B(n15462), .Z(n15457) );
  AND U15095 ( .A(n15463), .B(n15464), .Z(n15462) );
  XNOR U15096 ( .A(p_input[6329]), .B(n15461), .Z(n15464) );
  XNOR U15097 ( .A(n15461), .B(n15088), .Z(n15463) );
  IV U15098 ( .A(p_input[6297]), .Z(n15088) );
  XOR U15099 ( .A(n15465), .B(n15466), .Z(n15461) );
  AND U15100 ( .A(n15467), .B(n15468), .Z(n15466) );
  XNOR U15101 ( .A(p_input[6328]), .B(n15465), .Z(n15468) );
  XNOR U15102 ( .A(n15465), .B(n15097), .Z(n15467) );
  IV U15103 ( .A(p_input[6296]), .Z(n15097) );
  XOR U15104 ( .A(n15469), .B(n15470), .Z(n15465) );
  AND U15105 ( .A(n15471), .B(n15472), .Z(n15470) );
  XNOR U15106 ( .A(p_input[6327]), .B(n15469), .Z(n15472) );
  XNOR U15107 ( .A(n15469), .B(n15106), .Z(n15471) );
  IV U15108 ( .A(p_input[6295]), .Z(n15106) );
  XOR U15109 ( .A(n15473), .B(n15474), .Z(n15469) );
  AND U15110 ( .A(n15475), .B(n15476), .Z(n15474) );
  XNOR U15111 ( .A(p_input[6326]), .B(n15473), .Z(n15476) );
  XNOR U15112 ( .A(n15473), .B(n15115), .Z(n15475) );
  IV U15113 ( .A(p_input[6294]), .Z(n15115) );
  XOR U15114 ( .A(n15477), .B(n15478), .Z(n15473) );
  AND U15115 ( .A(n15479), .B(n15480), .Z(n15478) );
  XNOR U15116 ( .A(p_input[6325]), .B(n15477), .Z(n15480) );
  XNOR U15117 ( .A(n15477), .B(n15124), .Z(n15479) );
  IV U15118 ( .A(p_input[6293]), .Z(n15124) );
  XOR U15119 ( .A(n15481), .B(n15482), .Z(n15477) );
  AND U15120 ( .A(n15483), .B(n15484), .Z(n15482) );
  XNOR U15121 ( .A(p_input[6324]), .B(n15481), .Z(n15484) );
  XNOR U15122 ( .A(n15481), .B(n15133), .Z(n15483) );
  IV U15123 ( .A(p_input[6292]), .Z(n15133) );
  XOR U15124 ( .A(n15485), .B(n15486), .Z(n15481) );
  AND U15125 ( .A(n15487), .B(n15488), .Z(n15486) );
  XNOR U15126 ( .A(p_input[6323]), .B(n15485), .Z(n15488) );
  XNOR U15127 ( .A(n15485), .B(n15142), .Z(n15487) );
  IV U15128 ( .A(p_input[6291]), .Z(n15142) );
  XOR U15129 ( .A(n15489), .B(n15490), .Z(n15485) );
  AND U15130 ( .A(n15491), .B(n15492), .Z(n15490) );
  XNOR U15131 ( .A(p_input[6322]), .B(n15489), .Z(n15492) );
  XNOR U15132 ( .A(n15489), .B(n15151), .Z(n15491) );
  IV U15133 ( .A(p_input[6290]), .Z(n15151) );
  XOR U15134 ( .A(n15493), .B(n15494), .Z(n15489) );
  AND U15135 ( .A(n15495), .B(n15496), .Z(n15494) );
  XNOR U15136 ( .A(p_input[6321]), .B(n15493), .Z(n15496) );
  XNOR U15137 ( .A(n15493), .B(n15160), .Z(n15495) );
  IV U15138 ( .A(p_input[6289]), .Z(n15160) );
  XOR U15139 ( .A(n15497), .B(n15498), .Z(n15493) );
  AND U15140 ( .A(n15499), .B(n15500), .Z(n15498) );
  XNOR U15141 ( .A(p_input[6320]), .B(n15497), .Z(n15500) );
  XNOR U15142 ( .A(n15497), .B(n15169), .Z(n15499) );
  IV U15143 ( .A(p_input[6288]), .Z(n15169) );
  XOR U15144 ( .A(n15501), .B(n15502), .Z(n15497) );
  AND U15145 ( .A(n15503), .B(n15504), .Z(n15502) );
  XNOR U15146 ( .A(p_input[6319]), .B(n15501), .Z(n15504) );
  XNOR U15147 ( .A(n15501), .B(n15178), .Z(n15503) );
  IV U15148 ( .A(p_input[6287]), .Z(n15178) );
  XOR U15149 ( .A(n15505), .B(n15506), .Z(n15501) );
  AND U15150 ( .A(n15507), .B(n15508), .Z(n15506) );
  XNOR U15151 ( .A(p_input[6318]), .B(n15505), .Z(n15508) );
  XNOR U15152 ( .A(n15505), .B(n15187), .Z(n15507) );
  IV U15153 ( .A(p_input[6286]), .Z(n15187) );
  XOR U15154 ( .A(n15509), .B(n15510), .Z(n15505) );
  AND U15155 ( .A(n15511), .B(n15512), .Z(n15510) );
  XNOR U15156 ( .A(p_input[6317]), .B(n15509), .Z(n15512) );
  XNOR U15157 ( .A(n15509), .B(n15196), .Z(n15511) );
  IV U15158 ( .A(p_input[6285]), .Z(n15196) );
  XOR U15159 ( .A(n15513), .B(n15514), .Z(n15509) );
  AND U15160 ( .A(n15515), .B(n15516), .Z(n15514) );
  XNOR U15161 ( .A(p_input[6316]), .B(n15513), .Z(n15516) );
  XNOR U15162 ( .A(n15513), .B(n15205), .Z(n15515) );
  IV U15163 ( .A(p_input[6284]), .Z(n15205) );
  XOR U15164 ( .A(n15517), .B(n15518), .Z(n15513) );
  AND U15165 ( .A(n15519), .B(n15520), .Z(n15518) );
  XNOR U15166 ( .A(p_input[6315]), .B(n15517), .Z(n15520) );
  XNOR U15167 ( .A(n15517), .B(n15214), .Z(n15519) );
  IV U15168 ( .A(p_input[6283]), .Z(n15214) );
  XOR U15169 ( .A(n15521), .B(n15522), .Z(n15517) );
  AND U15170 ( .A(n15523), .B(n15524), .Z(n15522) );
  XNOR U15171 ( .A(p_input[6314]), .B(n15521), .Z(n15524) );
  XNOR U15172 ( .A(n15521), .B(n15223), .Z(n15523) );
  IV U15173 ( .A(p_input[6282]), .Z(n15223) );
  XOR U15174 ( .A(n15525), .B(n15526), .Z(n15521) );
  AND U15175 ( .A(n15527), .B(n15528), .Z(n15526) );
  XNOR U15176 ( .A(p_input[6313]), .B(n15525), .Z(n15528) );
  XNOR U15177 ( .A(n15525), .B(n15232), .Z(n15527) );
  IV U15178 ( .A(p_input[6281]), .Z(n15232) );
  XOR U15179 ( .A(n15529), .B(n15530), .Z(n15525) );
  AND U15180 ( .A(n15531), .B(n15532), .Z(n15530) );
  XNOR U15181 ( .A(p_input[6312]), .B(n15529), .Z(n15532) );
  XNOR U15182 ( .A(n15529), .B(n15241), .Z(n15531) );
  IV U15183 ( .A(p_input[6280]), .Z(n15241) );
  XOR U15184 ( .A(n15533), .B(n15534), .Z(n15529) );
  AND U15185 ( .A(n15535), .B(n15536), .Z(n15534) );
  XNOR U15186 ( .A(p_input[6311]), .B(n15533), .Z(n15536) );
  XNOR U15187 ( .A(n15533), .B(n15250), .Z(n15535) );
  IV U15188 ( .A(p_input[6279]), .Z(n15250) );
  XOR U15189 ( .A(n15537), .B(n15538), .Z(n15533) );
  AND U15190 ( .A(n15539), .B(n15540), .Z(n15538) );
  XNOR U15191 ( .A(p_input[6310]), .B(n15537), .Z(n15540) );
  XNOR U15192 ( .A(n15537), .B(n15259), .Z(n15539) );
  IV U15193 ( .A(p_input[6278]), .Z(n15259) );
  XOR U15194 ( .A(n15541), .B(n15542), .Z(n15537) );
  AND U15195 ( .A(n15543), .B(n15544), .Z(n15542) );
  XNOR U15196 ( .A(p_input[6309]), .B(n15541), .Z(n15544) );
  XNOR U15197 ( .A(n15541), .B(n15268), .Z(n15543) );
  IV U15198 ( .A(p_input[6277]), .Z(n15268) );
  XOR U15199 ( .A(n15545), .B(n15546), .Z(n15541) );
  AND U15200 ( .A(n15547), .B(n15548), .Z(n15546) );
  XNOR U15201 ( .A(p_input[6308]), .B(n15545), .Z(n15548) );
  XNOR U15202 ( .A(n15545), .B(n15277), .Z(n15547) );
  IV U15203 ( .A(p_input[6276]), .Z(n15277) );
  XOR U15204 ( .A(n15549), .B(n15550), .Z(n15545) );
  AND U15205 ( .A(n15551), .B(n15552), .Z(n15550) );
  XNOR U15206 ( .A(p_input[6307]), .B(n15549), .Z(n15552) );
  XNOR U15207 ( .A(n15549), .B(n15286), .Z(n15551) );
  IV U15208 ( .A(p_input[6275]), .Z(n15286) );
  XOR U15209 ( .A(n15553), .B(n15554), .Z(n15549) );
  AND U15210 ( .A(n15555), .B(n15556), .Z(n15554) );
  XNOR U15211 ( .A(p_input[6306]), .B(n15553), .Z(n15556) );
  XNOR U15212 ( .A(n15553), .B(n15295), .Z(n15555) );
  IV U15213 ( .A(p_input[6274]), .Z(n15295) );
  XNOR U15214 ( .A(n15557), .B(n15558), .Z(n15553) );
  AND U15215 ( .A(n15559), .B(n15560), .Z(n15558) );
  XOR U15216 ( .A(p_input[6305]), .B(n15557), .Z(n15560) );
  XNOR U15217 ( .A(p_input[6273]), .B(n15557), .Z(n15559) );
  AND U15218 ( .A(p_input[6304]), .B(n15561), .Z(n15557) );
  IV U15219 ( .A(p_input[6272]), .Z(n15561) );
  XOR U15220 ( .A(n15562), .B(n15563), .Z(n14651) );
  AND U15221 ( .A(n480), .B(n15564), .Z(n15563) );
  XNOR U15222 ( .A(n15565), .B(n15562), .Z(n15564) );
  XOR U15223 ( .A(n15566), .B(n15567), .Z(n480) );
  AND U15224 ( .A(n15568), .B(n15569), .Z(n15567) );
  XNOR U15225 ( .A(n14666), .B(n15566), .Z(n15569) );
  AND U15226 ( .A(p_input[6271]), .B(p_input[6239]), .Z(n14666) );
  XNOR U15227 ( .A(n15566), .B(n14663), .Z(n15568) );
  IV U15228 ( .A(n15570), .Z(n14663) );
  AND U15229 ( .A(p_input[6175]), .B(p_input[6207]), .Z(n15570) );
  XOR U15230 ( .A(n15571), .B(n15572), .Z(n15566) );
  AND U15231 ( .A(n15573), .B(n15574), .Z(n15572) );
  XOR U15232 ( .A(n15571), .B(n14678), .Z(n15574) );
  XNOR U15233 ( .A(p_input[6238]), .B(n15575), .Z(n14678) );
  AND U15234 ( .A(n291), .B(n15576), .Z(n15575) );
  XOR U15235 ( .A(p_input[6270]), .B(p_input[6238]), .Z(n15576) );
  XNOR U15236 ( .A(n14675), .B(n15571), .Z(n15573) );
  XOR U15237 ( .A(n15577), .B(n15578), .Z(n14675) );
  AND U15238 ( .A(n288), .B(n15579), .Z(n15578) );
  XOR U15239 ( .A(p_input[6206]), .B(p_input[6174]), .Z(n15579) );
  XOR U15240 ( .A(n15580), .B(n15581), .Z(n15571) );
  AND U15241 ( .A(n15582), .B(n15583), .Z(n15581) );
  XOR U15242 ( .A(n15580), .B(n14690), .Z(n15583) );
  XNOR U15243 ( .A(p_input[6237]), .B(n15584), .Z(n14690) );
  AND U15244 ( .A(n291), .B(n15585), .Z(n15584) );
  XOR U15245 ( .A(p_input[6269]), .B(p_input[6237]), .Z(n15585) );
  XNOR U15246 ( .A(n14687), .B(n15580), .Z(n15582) );
  XOR U15247 ( .A(n15586), .B(n15587), .Z(n14687) );
  AND U15248 ( .A(n288), .B(n15588), .Z(n15587) );
  XOR U15249 ( .A(p_input[6205]), .B(p_input[6173]), .Z(n15588) );
  XOR U15250 ( .A(n15589), .B(n15590), .Z(n15580) );
  AND U15251 ( .A(n15591), .B(n15592), .Z(n15590) );
  XOR U15252 ( .A(n15589), .B(n14702), .Z(n15592) );
  XNOR U15253 ( .A(p_input[6236]), .B(n15593), .Z(n14702) );
  AND U15254 ( .A(n291), .B(n15594), .Z(n15593) );
  XOR U15255 ( .A(p_input[6268]), .B(p_input[6236]), .Z(n15594) );
  XNOR U15256 ( .A(n14699), .B(n15589), .Z(n15591) );
  XOR U15257 ( .A(n15595), .B(n15596), .Z(n14699) );
  AND U15258 ( .A(n288), .B(n15597), .Z(n15596) );
  XOR U15259 ( .A(p_input[6204]), .B(p_input[6172]), .Z(n15597) );
  XOR U15260 ( .A(n15598), .B(n15599), .Z(n15589) );
  AND U15261 ( .A(n15600), .B(n15601), .Z(n15599) );
  XOR U15262 ( .A(n15598), .B(n14714), .Z(n15601) );
  XNOR U15263 ( .A(p_input[6235]), .B(n15602), .Z(n14714) );
  AND U15264 ( .A(n291), .B(n15603), .Z(n15602) );
  XOR U15265 ( .A(p_input[6267]), .B(p_input[6235]), .Z(n15603) );
  XNOR U15266 ( .A(n14711), .B(n15598), .Z(n15600) );
  XOR U15267 ( .A(n15604), .B(n15605), .Z(n14711) );
  AND U15268 ( .A(n288), .B(n15606), .Z(n15605) );
  XOR U15269 ( .A(p_input[6203]), .B(p_input[6171]), .Z(n15606) );
  XOR U15270 ( .A(n15607), .B(n15608), .Z(n15598) );
  AND U15271 ( .A(n15609), .B(n15610), .Z(n15608) );
  XOR U15272 ( .A(n15607), .B(n14726), .Z(n15610) );
  XNOR U15273 ( .A(p_input[6234]), .B(n15611), .Z(n14726) );
  AND U15274 ( .A(n291), .B(n15612), .Z(n15611) );
  XOR U15275 ( .A(p_input[6266]), .B(p_input[6234]), .Z(n15612) );
  XNOR U15276 ( .A(n14723), .B(n15607), .Z(n15609) );
  XOR U15277 ( .A(n15613), .B(n15614), .Z(n14723) );
  AND U15278 ( .A(n288), .B(n15615), .Z(n15614) );
  XOR U15279 ( .A(p_input[6202]), .B(p_input[6170]), .Z(n15615) );
  XOR U15280 ( .A(n15616), .B(n15617), .Z(n15607) );
  AND U15281 ( .A(n15618), .B(n15619), .Z(n15617) );
  XOR U15282 ( .A(n15616), .B(n14738), .Z(n15619) );
  XNOR U15283 ( .A(p_input[6233]), .B(n15620), .Z(n14738) );
  AND U15284 ( .A(n291), .B(n15621), .Z(n15620) );
  XOR U15285 ( .A(p_input[6265]), .B(p_input[6233]), .Z(n15621) );
  XNOR U15286 ( .A(n14735), .B(n15616), .Z(n15618) );
  XOR U15287 ( .A(n15622), .B(n15623), .Z(n14735) );
  AND U15288 ( .A(n288), .B(n15624), .Z(n15623) );
  XOR U15289 ( .A(p_input[6201]), .B(p_input[6169]), .Z(n15624) );
  XOR U15290 ( .A(n15625), .B(n15626), .Z(n15616) );
  AND U15291 ( .A(n15627), .B(n15628), .Z(n15626) );
  XOR U15292 ( .A(n15625), .B(n14750), .Z(n15628) );
  XNOR U15293 ( .A(p_input[6232]), .B(n15629), .Z(n14750) );
  AND U15294 ( .A(n291), .B(n15630), .Z(n15629) );
  XOR U15295 ( .A(p_input[6264]), .B(p_input[6232]), .Z(n15630) );
  XNOR U15296 ( .A(n14747), .B(n15625), .Z(n15627) );
  XOR U15297 ( .A(n15631), .B(n15632), .Z(n14747) );
  AND U15298 ( .A(n288), .B(n15633), .Z(n15632) );
  XOR U15299 ( .A(p_input[6200]), .B(p_input[6168]), .Z(n15633) );
  XOR U15300 ( .A(n15634), .B(n15635), .Z(n15625) );
  AND U15301 ( .A(n15636), .B(n15637), .Z(n15635) );
  XOR U15302 ( .A(n15634), .B(n14762), .Z(n15637) );
  XNOR U15303 ( .A(p_input[6231]), .B(n15638), .Z(n14762) );
  AND U15304 ( .A(n291), .B(n15639), .Z(n15638) );
  XOR U15305 ( .A(p_input[6263]), .B(p_input[6231]), .Z(n15639) );
  XNOR U15306 ( .A(n14759), .B(n15634), .Z(n15636) );
  XOR U15307 ( .A(n15640), .B(n15641), .Z(n14759) );
  AND U15308 ( .A(n288), .B(n15642), .Z(n15641) );
  XOR U15309 ( .A(p_input[6199]), .B(p_input[6167]), .Z(n15642) );
  XOR U15310 ( .A(n15643), .B(n15644), .Z(n15634) );
  AND U15311 ( .A(n15645), .B(n15646), .Z(n15644) );
  XOR U15312 ( .A(n15643), .B(n14774), .Z(n15646) );
  XNOR U15313 ( .A(p_input[6230]), .B(n15647), .Z(n14774) );
  AND U15314 ( .A(n291), .B(n15648), .Z(n15647) );
  XOR U15315 ( .A(p_input[6262]), .B(p_input[6230]), .Z(n15648) );
  XNOR U15316 ( .A(n14771), .B(n15643), .Z(n15645) );
  XOR U15317 ( .A(n15649), .B(n15650), .Z(n14771) );
  AND U15318 ( .A(n288), .B(n15651), .Z(n15650) );
  XOR U15319 ( .A(p_input[6198]), .B(p_input[6166]), .Z(n15651) );
  XOR U15320 ( .A(n15652), .B(n15653), .Z(n15643) );
  AND U15321 ( .A(n15654), .B(n15655), .Z(n15653) );
  XOR U15322 ( .A(n15652), .B(n14786), .Z(n15655) );
  XNOR U15323 ( .A(p_input[6229]), .B(n15656), .Z(n14786) );
  AND U15324 ( .A(n291), .B(n15657), .Z(n15656) );
  XOR U15325 ( .A(p_input[6261]), .B(p_input[6229]), .Z(n15657) );
  XNOR U15326 ( .A(n14783), .B(n15652), .Z(n15654) );
  XOR U15327 ( .A(n15658), .B(n15659), .Z(n14783) );
  AND U15328 ( .A(n288), .B(n15660), .Z(n15659) );
  XOR U15329 ( .A(p_input[6197]), .B(p_input[6165]), .Z(n15660) );
  XOR U15330 ( .A(n15661), .B(n15662), .Z(n15652) );
  AND U15331 ( .A(n15663), .B(n15664), .Z(n15662) );
  XOR U15332 ( .A(n15661), .B(n14798), .Z(n15664) );
  XNOR U15333 ( .A(p_input[6228]), .B(n15665), .Z(n14798) );
  AND U15334 ( .A(n291), .B(n15666), .Z(n15665) );
  XOR U15335 ( .A(p_input[6260]), .B(p_input[6228]), .Z(n15666) );
  XNOR U15336 ( .A(n14795), .B(n15661), .Z(n15663) );
  XOR U15337 ( .A(n15667), .B(n15668), .Z(n14795) );
  AND U15338 ( .A(n288), .B(n15669), .Z(n15668) );
  XOR U15339 ( .A(p_input[6196]), .B(p_input[6164]), .Z(n15669) );
  XOR U15340 ( .A(n15670), .B(n15671), .Z(n15661) );
  AND U15341 ( .A(n15672), .B(n15673), .Z(n15671) );
  XOR U15342 ( .A(n15670), .B(n14810), .Z(n15673) );
  XNOR U15343 ( .A(p_input[6227]), .B(n15674), .Z(n14810) );
  AND U15344 ( .A(n291), .B(n15675), .Z(n15674) );
  XOR U15345 ( .A(p_input[6259]), .B(p_input[6227]), .Z(n15675) );
  XNOR U15346 ( .A(n14807), .B(n15670), .Z(n15672) );
  XOR U15347 ( .A(n15676), .B(n15677), .Z(n14807) );
  AND U15348 ( .A(n288), .B(n15678), .Z(n15677) );
  XOR U15349 ( .A(p_input[6195]), .B(p_input[6163]), .Z(n15678) );
  XOR U15350 ( .A(n15679), .B(n15680), .Z(n15670) );
  AND U15351 ( .A(n15681), .B(n15682), .Z(n15680) );
  XOR U15352 ( .A(n15679), .B(n14822), .Z(n15682) );
  XNOR U15353 ( .A(p_input[6226]), .B(n15683), .Z(n14822) );
  AND U15354 ( .A(n291), .B(n15684), .Z(n15683) );
  XOR U15355 ( .A(p_input[6258]), .B(p_input[6226]), .Z(n15684) );
  XNOR U15356 ( .A(n14819), .B(n15679), .Z(n15681) );
  XOR U15357 ( .A(n15685), .B(n15686), .Z(n14819) );
  AND U15358 ( .A(n288), .B(n15687), .Z(n15686) );
  XOR U15359 ( .A(p_input[6194]), .B(p_input[6162]), .Z(n15687) );
  XOR U15360 ( .A(n15688), .B(n15689), .Z(n15679) );
  AND U15361 ( .A(n15690), .B(n15691), .Z(n15689) );
  XOR U15362 ( .A(n15688), .B(n14834), .Z(n15691) );
  XNOR U15363 ( .A(p_input[6225]), .B(n15692), .Z(n14834) );
  AND U15364 ( .A(n291), .B(n15693), .Z(n15692) );
  XOR U15365 ( .A(p_input[6257]), .B(p_input[6225]), .Z(n15693) );
  XNOR U15366 ( .A(n14831), .B(n15688), .Z(n15690) );
  XOR U15367 ( .A(n15694), .B(n15695), .Z(n14831) );
  AND U15368 ( .A(n288), .B(n15696), .Z(n15695) );
  XOR U15369 ( .A(p_input[6193]), .B(p_input[6161]), .Z(n15696) );
  XOR U15370 ( .A(n15697), .B(n15698), .Z(n15688) );
  AND U15371 ( .A(n15699), .B(n15700), .Z(n15698) );
  XOR U15372 ( .A(n15697), .B(n14846), .Z(n15700) );
  XNOR U15373 ( .A(p_input[6224]), .B(n15701), .Z(n14846) );
  AND U15374 ( .A(n291), .B(n15702), .Z(n15701) );
  XOR U15375 ( .A(p_input[6256]), .B(p_input[6224]), .Z(n15702) );
  XNOR U15376 ( .A(n14843), .B(n15697), .Z(n15699) );
  XOR U15377 ( .A(n15703), .B(n15704), .Z(n14843) );
  AND U15378 ( .A(n288), .B(n15705), .Z(n15704) );
  XOR U15379 ( .A(p_input[6192]), .B(p_input[6160]), .Z(n15705) );
  XOR U15380 ( .A(n15706), .B(n15707), .Z(n15697) );
  AND U15381 ( .A(n15708), .B(n15709), .Z(n15707) );
  XOR U15382 ( .A(n15706), .B(n14858), .Z(n15709) );
  XNOR U15383 ( .A(p_input[6223]), .B(n15710), .Z(n14858) );
  AND U15384 ( .A(n291), .B(n15711), .Z(n15710) );
  XOR U15385 ( .A(p_input[6255]), .B(p_input[6223]), .Z(n15711) );
  XNOR U15386 ( .A(n14855), .B(n15706), .Z(n15708) );
  XOR U15387 ( .A(n15712), .B(n15713), .Z(n14855) );
  AND U15388 ( .A(n288), .B(n15714), .Z(n15713) );
  XOR U15389 ( .A(p_input[6191]), .B(p_input[6159]), .Z(n15714) );
  XOR U15390 ( .A(n15715), .B(n15716), .Z(n15706) );
  AND U15391 ( .A(n15717), .B(n15718), .Z(n15716) );
  XOR U15392 ( .A(n15715), .B(n14870), .Z(n15718) );
  XNOR U15393 ( .A(p_input[6222]), .B(n15719), .Z(n14870) );
  AND U15394 ( .A(n291), .B(n15720), .Z(n15719) );
  XOR U15395 ( .A(p_input[6254]), .B(p_input[6222]), .Z(n15720) );
  XNOR U15396 ( .A(n14867), .B(n15715), .Z(n15717) );
  XOR U15397 ( .A(n15721), .B(n15722), .Z(n14867) );
  AND U15398 ( .A(n288), .B(n15723), .Z(n15722) );
  XOR U15399 ( .A(p_input[6190]), .B(p_input[6158]), .Z(n15723) );
  XOR U15400 ( .A(n15724), .B(n15725), .Z(n15715) );
  AND U15401 ( .A(n15726), .B(n15727), .Z(n15725) );
  XOR U15402 ( .A(n15724), .B(n14882), .Z(n15727) );
  XNOR U15403 ( .A(p_input[6221]), .B(n15728), .Z(n14882) );
  AND U15404 ( .A(n291), .B(n15729), .Z(n15728) );
  XOR U15405 ( .A(p_input[6253]), .B(p_input[6221]), .Z(n15729) );
  XNOR U15406 ( .A(n14879), .B(n15724), .Z(n15726) );
  XOR U15407 ( .A(n15730), .B(n15731), .Z(n14879) );
  AND U15408 ( .A(n288), .B(n15732), .Z(n15731) );
  XOR U15409 ( .A(p_input[6189]), .B(p_input[6157]), .Z(n15732) );
  XOR U15410 ( .A(n15733), .B(n15734), .Z(n15724) );
  AND U15411 ( .A(n15735), .B(n15736), .Z(n15734) );
  XOR U15412 ( .A(n15733), .B(n14894), .Z(n15736) );
  XNOR U15413 ( .A(p_input[6220]), .B(n15737), .Z(n14894) );
  AND U15414 ( .A(n291), .B(n15738), .Z(n15737) );
  XOR U15415 ( .A(p_input[6252]), .B(p_input[6220]), .Z(n15738) );
  XNOR U15416 ( .A(n14891), .B(n15733), .Z(n15735) );
  XOR U15417 ( .A(n15739), .B(n15740), .Z(n14891) );
  AND U15418 ( .A(n288), .B(n15741), .Z(n15740) );
  XOR U15419 ( .A(p_input[6188]), .B(p_input[6156]), .Z(n15741) );
  XOR U15420 ( .A(n15742), .B(n15743), .Z(n15733) );
  AND U15421 ( .A(n15744), .B(n15745), .Z(n15743) );
  XOR U15422 ( .A(n15742), .B(n14906), .Z(n15745) );
  XNOR U15423 ( .A(p_input[6219]), .B(n15746), .Z(n14906) );
  AND U15424 ( .A(n291), .B(n15747), .Z(n15746) );
  XOR U15425 ( .A(p_input[6251]), .B(p_input[6219]), .Z(n15747) );
  XNOR U15426 ( .A(n14903), .B(n15742), .Z(n15744) );
  XOR U15427 ( .A(n15748), .B(n15749), .Z(n14903) );
  AND U15428 ( .A(n288), .B(n15750), .Z(n15749) );
  XOR U15429 ( .A(p_input[6187]), .B(p_input[6155]), .Z(n15750) );
  XOR U15430 ( .A(n15751), .B(n15752), .Z(n15742) );
  AND U15431 ( .A(n15753), .B(n15754), .Z(n15752) );
  XOR U15432 ( .A(n15751), .B(n14918), .Z(n15754) );
  XNOR U15433 ( .A(p_input[6218]), .B(n15755), .Z(n14918) );
  AND U15434 ( .A(n291), .B(n15756), .Z(n15755) );
  XOR U15435 ( .A(p_input[6250]), .B(p_input[6218]), .Z(n15756) );
  XNOR U15436 ( .A(n14915), .B(n15751), .Z(n15753) );
  XOR U15437 ( .A(n15757), .B(n15758), .Z(n14915) );
  AND U15438 ( .A(n288), .B(n15759), .Z(n15758) );
  XOR U15439 ( .A(p_input[6186]), .B(p_input[6154]), .Z(n15759) );
  XOR U15440 ( .A(n15760), .B(n15761), .Z(n15751) );
  AND U15441 ( .A(n15762), .B(n15763), .Z(n15761) );
  XOR U15442 ( .A(n15760), .B(n14930), .Z(n15763) );
  XNOR U15443 ( .A(p_input[6217]), .B(n15764), .Z(n14930) );
  AND U15444 ( .A(n291), .B(n15765), .Z(n15764) );
  XOR U15445 ( .A(p_input[6249]), .B(p_input[6217]), .Z(n15765) );
  XNOR U15446 ( .A(n14927), .B(n15760), .Z(n15762) );
  XOR U15447 ( .A(n15766), .B(n15767), .Z(n14927) );
  AND U15448 ( .A(n288), .B(n15768), .Z(n15767) );
  XOR U15449 ( .A(p_input[6185]), .B(p_input[6153]), .Z(n15768) );
  XOR U15450 ( .A(n15769), .B(n15770), .Z(n15760) );
  AND U15451 ( .A(n15771), .B(n15772), .Z(n15770) );
  XOR U15452 ( .A(n15769), .B(n14942), .Z(n15772) );
  XNOR U15453 ( .A(p_input[6216]), .B(n15773), .Z(n14942) );
  AND U15454 ( .A(n291), .B(n15774), .Z(n15773) );
  XOR U15455 ( .A(p_input[6248]), .B(p_input[6216]), .Z(n15774) );
  XNOR U15456 ( .A(n14939), .B(n15769), .Z(n15771) );
  XOR U15457 ( .A(n15775), .B(n15776), .Z(n14939) );
  AND U15458 ( .A(n288), .B(n15777), .Z(n15776) );
  XOR U15459 ( .A(p_input[6184]), .B(p_input[6152]), .Z(n15777) );
  XOR U15460 ( .A(n15778), .B(n15779), .Z(n15769) );
  AND U15461 ( .A(n15780), .B(n15781), .Z(n15779) );
  XOR U15462 ( .A(n15778), .B(n14954), .Z(n15781) );
  XNOR U15463 ( .A(p_input[6215]), .B(n15782), .Z(n14954) );
  AND U15464 ( .A(n291), .B(n15783), .Z(n15782) );
  XOR U15465 ( .A(p_input[6247]), .B(p_input[6215]), .Z(n15783) );
  XNOR U15466 ( .A(n14951), .B(n15778), .Z(n15780) );
  XOR U15467 ( .A(n15784), .B(n15785), .Z(n14951) );
  AND U15468 ( .A(n288), .B(n15786), .Z(n15785) );
  XOR U15469 ( .A(p_input[6183]), .B(p_input[6151]), .Z(n15786) );
  XOR U15470 ( .A(n15787), .B(n15788), .Z(n15778) );
  AND U15471 ( .A(n15789), .B(n15790), .Z(n15788) );
  XOR U15472 ( .A(n15787), .B(n14966), .Z(n15790) );
  XNOR U15473 ( .A(p_input[6214]), .B(n15791), .Z(n14966) );
  AND U15474 ( .A(n291), .B(n15792), .Z(n15791) );
  XOR U15475 ( .A(p_input[6246]), .B(p_input[6214]), .Z(n15792) );
  XNOR U15476 ( .A(n14963), .B(n15787), .Z(n15789) );
  XOR U15477 ( .A(n15793), .B(n15794), .Z(n14963) );
  AND U15478 ( .A(n288), .B(n15795), .Z(n15794) );
  XOR U15479 ( .A(p_input[6182]), .B(p_input[6150]), .Z(n15795) );
  XOR U15480 ( .A(n15796), .B(n15797), .Z(n15787) );
  AND U15481 ( .A(n15798), .B(n15799), .Z(n15797) );
  XOR U15482 ( .A(n15796), .B(n14978), .Z(n15799) );
  XNOR U15483 ( .A(p_input[6213]), .B(n15800), .Z(n14978) );
  AND U15484 ( .A(n291), .B(n15801), .Z(n15800) );
  XOR U15485 ( .A(p_input[6245]), .B(p_input[6213]), .Z(n15801) );
  XNOR U15486 ( .A(n14975), .B(n15796), .Z(n15798) );
  XOR U15487 ( .A(n15802), .B(n15803), .Z(n14975) );
  AND U15488 ( .A(n288), .B(n15804), .Z(n15803) );
  XOR U15489 ( .A(p_input[6181]), .B(p_input[6149]), .Z(n15804) );
  XOR U15490 ( .A(n15805), .B(n15806), .Z(n15796) );
  AND U15491 ( .A(n15807), .B(n15808), .Z(n15806) );
  XOR U15492 ( .A(n15805), .B(n14990), .Z(n15808) );
  XNOR U15493 ( .A(p_input[6212]), .B(n15809), .Z(n14990) );
  AND U15494 ( .A(n291), .B(n15810), .Z(n15809) );
  XOR U15495 ( .A(p_input[6244]), .B(p_input[6212]), .Z(n15810) );
  XNOR U15496 ( .A(n14987), .B(n15805), .Z(n15807) );
  XOR U15497 ( .A(n15811), .B(n15812), .Z(n14987) );
  AND U15498 ( .A(n288), .B(n15813), .Z(n15812) );
  XOR U15499 ( .A(p_input[6180]), .B(p_input[6148]), .Z(n15813) );
  XOR U15500 ( .A(n15814), .B(n15815), .Z(n15805) );
  AND U15501 ( .A(n15816), .B(n15817), .Z(n15815) );
  XOR U15502 ( .A(n15814), .B(n15002), .Z(n15817) );
  XNOR U15503 ( .A(p_input[6211]), .B(n15818), .Z(n15002) );
  AND U15504 ( .A(n291), .B(n15819), .Z(n15818) );
  XOR U15505 ( .A(p_input[6243]), .B(p_input[6211]), .Z(n15819) );
  XNOR U15506 ( .A(n14999), .B(n15814), .Z(n15816) );
  XOR U15507 ( .A(n15820), .B(n15821), .Z(n14999) );
  AND U15508 ( .A(n288), .B(n15822), .Z(n15821) );
  XOR U15509 ( .A(p_input[6179]), .B(p_input[6147]), .Z(n15822) );
  XOR U15510 ( .A(n15823), .B(n15824), .Z(n15814) );
  AND U15511 ( .A(n15825), .B(n15826), .Z(n15824) );
  XOR U15512 ( .A(n15823), .B(n15014), .Z(n15826) );
  XNOR U15513 ( .A(p_input[6210]), .B(n15827), .Z(n15014) );
  AND U15514 ( .A(n291), .B(n15828), .Z(n15827) );
  XOR U15515 ( .A(p_input[6242]), .B(p_input[6210]), .Z(n15828) );
  XNOR U15516 ( .A(n15011), .B(n15823), .Z(n15825) );
  XOR U15517 ( .A(n15829), .B(n15830), .Z(n15011) );
  AND U15518 ( .A(n288), .B(n15831), .Z(n15830) );
  XOR U15519 ( .A(p_input[6178]), .B(p_input[6146]), .Z(n15831) );
  XOR U15520 ( .A(n15832), .B(n15833), .Z(n15823) );
  AND U15521 ( .A(n15834), .B(n15835), .Z(n15833) );
  XNOR U15522 ( .A(n15836), .B(n15027), .Z(n15835) );
  XNOR U15523 ( .A(p_input[6209]), .B(n15837), .Z(n15027) );
  AND U15524 ( .A(n291), .B(n15838), .Z(n15837) );
  XNOR U15525 ( .A(p_input[6241]), .B(n15839), .Z(n15838) );
  IV U15526 ( .A(p_input[6209]), .Z(n15839) );
  XNOR U15527 ( .A(n15024), .B(n15832), .Z(n15834) );
  XNOR U15528 ( .A(p_input[6145]), .B(n15840), .Z(n15024) );
  AND U15529 ( .A(n288), .B(n15841), .Z(n15840) );
  XOR U15530 ( .A(p_input[6177]), .B(p_input[6145]), .Z(n15841) );
  IV U15531 ( .A(n15836), .Z(n15832) );
  AND U15532 ( .A(n15562), .B(n15565), .Z(n15836) );
  XOR U15533 ( .A(p_input[6208]), .B(n15842), .Z(n15565) );
  AND U15534 ( .A(n291), .B(n15843), .Z(n15842) );
  XOR U15535 ( .A(p_input[6240]), .B(p_input[6208]), .Z(n15843) );
  XOR U15536 ( .A(n15844), .B(n15845), .Z(n291) );
  AND U15537 ( .A(n15846), .B(n15847), .Z(n15845) );
  XNOR U15538 ( .A(p_input[6271]), .B(n15844), .Z(n15847) );
  XOR U15539 ( .A(n15844), .B(p_input[6239]), .Z(n15846) );
  XOR U15540 ( .A(n15848), .B(n15849), .Z(n15844) );
  AND U15541 ( .A(n15850), .B(n15851), .Z(n15849) );
  XNOR U15542 ( .A(p_input[6270]), .B(n15848), .Z(n15851) );
  XOR U15543 ( .A(n15848), .B(p_input[6238]), .Z(n15850) );
  XOR U15544 ( .A(n15852), .B(n15853), .Z(n15848) );
  AND U15545 ( .A(n15854), .B(n15855), .Z(n15853) );
  XNOR U15546 ( .A(p_input[6269]), .B(n15852), .Z(n15855) );
  XOR U15547 ( .A(n15852), .B(p_input[6237]), .Z(n15854) );
  XOR U15548 ( .A(n15856), .B(n15857), .Z(n15852) );
  AND U15549 ( .A(n15858), .B(n15859), .Z(n15857) );
  XNOR U15550 ( .A(p_input[6268]), .B(n15856), .Z(n15859) );
  XOR U15551 ( .A(n15856), .B(p_input[6236]), .Z(n15858) );
  XOR U15552 ( .A(n15860), .B(n15861), .Z(n15856) );
  AND U15553 ( .A(n15862), .B(n15863), .Z(n15861) );
  XNOR U15554 ( .A(p_input[6267]), .B(n15860), .Z(n15863) );
  XOR U15555 ( .A(n15860), .B(p_input[6235]), .Z(n15862) );
  XOR U15556 ( .A(n15864), .B(n15865), .Z(n15860) );
  AND U15557 ( .A(n15866), .B(n15867), .Z(n15865) );
  XNOR U15558 ( .A(p_input[6266]), .B(n15864), .Z(n15867) );
  XOR U15559 ( .A(n15864), .B(p_input[6234]), .Z(n15866) );
  XOR U15560 ( .A(n15868), .B(n15869), .Z(n15864) );
  AND U15561 ( .A(n15870), .B(n15871), .Z(n15869) );
  XNOR U15562 ( .A(p_input[6265]), .B(n15868), .Z(n15871) );
  XOR U15563 ( .A(n15868), .B(p_input[6233]), .Z(n15870) );
  XOR U15564 ( .A(n15872), .B(n15873), .Z(n15868) );
  AND U15565 ( .A(n15874), .B(n15875), .Z(n15873) );
  XNOR U15566 ( .A(p_input[6264]), .B(n15872), .Z(n15875) );
  XOR U15567 ( .A(n15872), .B(p_input[6232]), .Z(n15874) );
  XOR U15568 ( .A(n15876), .B(n15877), .Z(n15872) );
  AND U15569 ( .A(n15878), .B(n15879), .Z(n15877) );
  XNOR U15570 ( .A(p_input[6263]), .B(n15876), .Z(n15879) );
  XOR U15571 ( .A(n15876), .B(p_input[6231]), .Z(n15878) );
  XOR U15572 ( .A(n15880), .B(n15881), .Z(n15876) );
  AND U15573 ( .A(n15882), .B(n15883), .Z(n15881) );
  XNOR U15574 ( .A(p_input[6262]), .B(n15880), .Z(n15883) );
  XOR U15575 ( .A(n15880), .B(p_input[6230]), .Z(n15882) );
  XOR U15576 ( .A(n15884), .B(n15885), .Z(n15880) );
  AND U15577 ( .A(n15886), .B(n15887), .Z(n15885) );
  XNOR U15578 ( .A(p_input[6261]), .B(n15884), .Z(n15887) );
  XOR U15579 ( .A(n15884), .B(p_input[6229]), .Z(n15886) );
  XOR U15580 ( .A(n15888), .B(n15889), .Z(n15884) );
  AND U15581 ( .A(n15890), .B(n15891), .Z(n15889) );
  XNOR U15582 ( .A(p_input[6260]), .B(n15888), .Z(n15891) );
  XOR U15583 ( .A(n15888), .B(p_input[6228]), .Z(n15890) );
  XOR U15584 ( .A(n15892), .B(n15893), .Z(n15888) );
  AND U15585 ( .A(n15894), .B(n15895), .Z(n15893) );
  XNOR U15586 ( .A(p_input[6259]), .B(n15892), .Z(n15895) );
  XOR U15587 ( .A(n15892), .B(p_input[6227]), .Z(n15894) );
  XOR U15588 ( .A(n15896), .B(n15897), .Z(n15892) );
  AND U15589 ( .A(n15898), .B(n15899), .Z(n15897) );
  XNOR U15590 ( .A(p_input[6258]), .B(n15896), .Z(n15899) );
  XOR U15591 ( .A(n15896), .B(p_input[6226]), .Z(n15898) );
  XOR U15592 ( .A(n15900), .B(n15901), .Z(n15896) );
  AND U15593 ( .A(n15902), .B(n15903), .Z(n15901) );
  XNOR U15594 ( .A(p_input[6257]), .B(n15900), .Z(n15903) );
  XOR U15595 ( .A(n15900), .B(p_input[6225]), .Z(n15902) );
  XOR U15596 ( .A(n15904), .B(n15905), .Z(n15900) );
  AND U15597 ( .A(n15906), .B(n15907), .Z(n15905) );
  XNOR U15598 ( .A(p_input[6256]), .B(n15904), .Z(n15907) );
  XOR U15599 ( .A(n15904), .B(p_input[6224]), .Z(n15906) );
  XOR U15600 ( .A(n15908), .B(n15909), .Z(n15904) );
  AND U15601 ( .A(n15910), .B(n15911), .Z(n15909) );
  XNOR U15602 ( .A(p_input[6255]), .B(n15908), .Z(n15911) );
  XOR U15603 ( .A(n15908), .B(p_input[6223]), .Z(n15910) );
  XOR U15604 ( .A(n15912), .B(n15913), .Z(n15908) );
  AND U15605 ( .A(n15914), .B(n15915), .Z(n15913) );
  XNOR U15606 ( .A(p_input[6254]), .B(n15912), .Z(n15915) );
  XOR U15607 ( .A(n15912), .B(p_input[6222]), .Z(n15914) );
  XOR U15608 ( .A(n15916), .B(n15917), .Z(n15912) );
  AND U15609 ( .A(n15918), .B(n15919), .Z(n15917) );
  XNOR U15610 ( .A(p_input[6253]), .B(n15916), .Z(n15919) );
  XOR U15611 ( .A(n15916), .B(p_input[6221]), .Z(n15918) );
  XOR U15612 ( .A(n15920), .B(n15921), .Z(n15916) );
  AND U15613 ( .A(n15922), .B(n15923), .Z(n15921) );
  XNOR U15614 ( .A(p_input[6252]), .B(n15920), .Z(n15923) );
  XOR U15615 ( .A(n15920), .B(p_input[6220]), .Z(n15922) );
  XOR U15616 ( .A(n15924), .B(n15925), .Z(n15920) );
  AND U15617 ( .A(n15926), .B(n15927), .Z(n15925) );
  XNOR U15618 ( .A(p_input[6251]), .B(n15924), .Z(n15927) );
  XOR U15619 ( .A(n15924), .B(p_input[6219]), .Z(n15926) );
  XOR U15620 ( .A(n15928), .B(n15929), .Z(n15924) );
  AND U15621 ( .A(n15930), .B(n15931), .Z(n15929) );
  XNOR U15622 ( .A(p_input[6250]), .B(n15928), .Z(n15931) );
  XOR U15623 ( .A(n15928), .B(p_input[6218]), .Z(n15930) );
  XOR U15624 ( .A(n15932), .B(n15933), .Z(n15928) );
  AND U15625 ( .A(n15934), .B(n15935), .Z(n15933) );
  XNOR U15626 ( .A(p_input[6249]), .B(n15932), .Z(n15935) );
  XOR U15627 ( .A(n15932), .B(p_input[6217]), .Z(n15934) );
  XOR U15628 ( .A(n15936), .B(n15937), .Z(n15932) );
  AND U15629 ( .A(n15938), .B(n15939), .Z(n15937) );
  XNOR U15630 ( .A(p_input[6248]), .B(n15936), .Z(n15939) );
  XOR U15631 ( .A(n15936), .B(p_input[6216]), .Z(n15938) );
  XOR U15632 ( .A(n15940), .B(n15941), .Z(n15936) );
  AND U15633 ( .A(n15942), .B(n15943), .Z(n15941) );
  XNOR U15634 ( .A(p_input[6247]), .B(n15940), .Z(n15943) );
  XOR U15635 ( .A(n15940), .B(p_input[6215]), .Z(n15942) );
  XOR U15636 ( .A(n15944), .B(n15945), .Z(n15940) );
  AND U15637 ( .A(n15946), .B(n15947), .Z(n15945) );
  XNOR U15638 ( .A(p_input[6246]), .B(n15944), .Z(n15947) );
  XOR U15639 ( .A(n15944), .B(p_input[6214]), .Z(n15946) );
  XOR U15640 ( .A(n15948), .B(n15949), .Z(n15944) );
  AND U15641 ( .A(n15950), .B(n15951), .Z(n15949) );
  XNOR U15642 ( .A(p_input[6245]), .B(n15948), .Z(n15951) );
  XOR U15643 ( .A(n15948), .B(p_input[6213]), .Z(n15950) );
  XOR U15644 ( .A(n15952), .B(n15953), .Z(n15948) );
  AND U15645 ( .A(n15954), .B(n15955), .Z(n15953) );
  XNOR U15646 ( .A(p_input[6244]), .B(n15952), .Z(n15955) );
  XOR U15647 ( .A(n15952), .B(p_input[6212]), .Z(n15954) );
  XOR U15648 ( .A(n15956), .B(n15957), .Z(n15952) );
  AND U15649 ( .A(n15958), .B(n15959), .Z(n15957) );
  XNOR U15650 ( .A(p_input[6243]), .B(n15956), .Z(n15959) );
  XOR U15651 ( .A(n15956), .B(p_input[6211]), .Z(n15958) );
  XOR U15652 ( .A(n15960), .B(n15961), .Z(n15956) );
  AND U15653 ( .A(n15962), .B(n15963), .Z(n15961) );
  XNOR U15654 ( .A(p_input[6242]), .B(n15960), .Z(n15963) );
  XOR U15655 ( .A(n15960), .B(p_input[6210]), .Z(n15962) );
  XNOR U15656 ( .A(n15964), .B(n15965), .Z(n15960) );
  AND U15657 ( .A(n15966), .B(n15967), .Z(n15965) );
  XOR U15658 ( .A(p_input[6241]), .B(n15964), .Z(n15967) );
  XNOR U15659 ( .A(p_input[6209]), .B(n15964), .Z(n15966) );
  AND U15660 ( .A(p_input[6240]), .B(n15968), .Z(n15964) );
  IV U15661 ( .A(p_input[6208]), .Z(n15968) );
  XNOR U15662 ( .A(p_input[6144]), .B(n15969), .Z(n15562) );
  AND U15663 ( .A(n288), .B(n15970), .Z(n15969) );
  XOR U15664 ( .A(p_input[6176]), .B(p_input[6144]), .Z(n15970) );
  XOR U15665 ( .A(n15971), .B(n15972), .Z(n288) );
  AND U15666 ( .A(n15973), .B(n15974), .Z(n15972) );
  XNOR U15667 ( .A(p_input[6207]), .B(n15971), .Z(n15974) );
  XOR U15668 ( .A(n15971), .B(p_input[6175]), .Z(n15973) );
  XOR U15669 ( .A(n15975), .B(n15976), .Z(n15971) );
  AND U15670 ( .A(n15977), .B(n15978), .Z(n15976) );
  XNOR U15671 ( .A(p_input[6206]), .B(n15975), .Z(n15978) );
  XNOR U15672 ( .A(n15975), .B(n15577), .Z(n15977) );
  IV U15673 ( .A(p_input[6174]), .Z(n15577) );
  XOR U15674 ( .A(n15979), .B(n15980), .Z(n15975) );
  AND U15675 ( .A(n15981), .B(n15982), .Z(n15980) );
  XNOR U15676 ( .A(p_input[6205]), .B(n15979), .Z(n15982) );
  XNOR U15677 ( .A(n15979), .B(n15586), .Z(n15981) );
  IV U15678 ( .A(p_input[6173]), .Z(n15586) );
  XOR U15679 ( .A(n15983), .B(n15984), .Z(n15979) );
  AND U15680 ( .A(n15985), .B(n15986), .Z(n15984) );
  XNOR U15681 ( .A(p_input[6204]), .B(n15983), .Z(n15986) );
  XNOR U15682 ( .A(n15983), .B(n15595), .Z(n15985) );
  IV U15683 ( .A(p_input[6172]), .Z(n15595) );
  XOR U15684 ( .A(n15987), .B(n15988), .Z(n15983) );
  AND U15685 ( .A(n15989), .B(n15990), .Z(n15988) );
  XNOR U15686 ( .A(p_input[6203]), .B(n15987), .Z(n15990) );
  XNOR U15687 ( .A(n15987), .B(n15604), .Z(n15989) );
  IV U15688 ( .A(p_input[6171]), .Z(n15604) );
  XOR U15689 ( .A(n15991), .B(n15992), .Z(n15987) );
  AND U15690 ( .A(n15993), .B(n15994), .Z(n15992) );
  XNOR U15691 ( .A(p_input[6202]), .B(n15991), .Z(n15994) );
  XNOR U15692 ( .A(n15991), .B(n15613), .Z(n15993) );
  IV U15693 ( .A(p_input[6170]), .Z(n15613) );
  XOR U15694 ( .A(n15995), .B(n15996), .Z(n15991) );
  AND U15695 ( .A(n15997), .B(n15998), .Z(n15996) );
  XNOR U15696 ( .A(p_input[6201]), .B(n15995), .Z(n15998) );
  XNOR U15697 ( .A(n15995), .B(n15622), .Z(n15997) );
  IV U15698 ( .A(p_input[6169]), .Z(n15622) );
  XOR U15699 ( .A(n15999), .B(n16000), .Z(n15995) );
  AND U15700 ( .A(n16001), .B(n16002), .Z(n16000) );
  XNOR U15701 ( .A(p_input[6200]), .B(n15999), .Z(n16002) );
  XNOR U15702 ( .A(n15999), .B(n15631), .Z(n16001) );
  IV U15703 ( .A(p_input[6168]), .Z(n15631) );
  XOR U15704 ( .A(n16003), .B(n16004), .Z(n15999) );
  AND U15705 ( .A(n16005), .B(n16006), .Z(n16004) );
  XNOR U15706 ( .A(p_input[6199]), .B(n16003), .Z(n16006) );
  XNOR U15707 ( .A(n16003), .B(n15640), .Z(n16005) );
  IV U15708 ( .A(p_input[6167]), .Z(n15640) );
  XOR U15709 ( .A(n16007), .B(n16008), .Z(n16003) );
  AND U15710 ( .A(n16009), .B(n16010), .Z(n16008) );
  XNOR U15711 ( .A(p_input[6198]), .B(n16007), .Z(n16010) );
  XNOR U15712 ( .A(n16007), .B(n15649), .Z(n16009) );
  IV U15713 ( .A(p_input[6166]), .Z(n15649) );
  XOR U15714 ( .A(n16011), .B(n16012), .Z(n16007) );
  AND U15715 ( .A(n16013), .B(n16014), .Z(n16012) );
  XNOR U15716 ( .A(p_input[6197]), .B(n16011), .Z(n16014) );
  XNOR U15717 ( .A(n16011), .B(n15658), .Z(n16013) );
  IV U15718 ( .A(p_input[6165]), .Z(n15658) );
  XOR U15719 ( .A(n16015), .B(n16016), .Z(n16011) );
  AND U15720 ( .A(n16017), .B(n16018), .Z(n16016) );
  XNOR U15721 ( .A(p_input[6196]), .B(n16015), .Z(n16018) );
  XNOR U15722 ( .A(n16015), .B(n15667), .Z(n16017) );
  IV U15723 ( .A(p_input[6164]), .Z(n15667) );
  XOR U15724 ( .A(n16019), .B(n16020), .Z(n16015) );
  AND U15725 ( .A(n16021), .B(n16022), .Z(n16020) );
  XNOR U15726 ( .A(p_input[6195]), .B(n16019), .Z(n16022) );
  XNOR U15727 ( .A(n16019), .B(n15676), .Z(n16021) );
  IV U15728 ( .A(p_input[6163]), .Z(n15676) );
  XOR U15729 ( .A(n16023), .B(n16024), .Z(n16019) );
  AND U15730 ( .A(n16025), .B(n16026), .Z(n16024) );
  XNOR U15731 ( .A(p_input[6194]), .B(n16023), .Z(n16026) );
  XNOR U15732 ( .A(n16023), .B(n15685), .Z(n16025) );
  IV U15733 ( .A(p_input[6162]), .Z(n15685) );
  XOR U15734 ( .A(n16027), .B(n16028), .Z(n16023) );
  AND U15735 ( .A(n16029), .B(n16030), .Z(n16028) );
  XNOR U15736 ( .A(p_input[6193]), .B(n16027), .Z(n16030) );
  XNOR U15737 ( .A(n16027), .B(n15694), .Z(n16029) );
  IV U15738 ( .A(p_input[6161]), .Z(n15694) );
  XOR U15739 ( .A(n16031), .B(n16032), .Z(n16027) );
  AND U15740 ( .A(n16033), .B(n16034), .Z(n16032) );
  XNOR U15741 ( .A(p_input[6192]), .B(n16031), .Z(n16034) );
  XNOR U15742 ( .A(n16031), .B(n15703), .Z(n16033) );
  IV U15743 ( .A(p_input[6160]), .Z(n15703) );
  XOR U15744 ( .A(n16035), .B(n16036), .Z(n16031) );
  AND U15745 ( .A(n16037), .B(n16038), .Z(n16036) );
  XNOR U15746 ( .A(p_input[6191]), .B(n16035), .Z(n16038) );
  XNOR U15747 ( .A(n16035), .B(n15712), .Z(n16037) );
  IV U15748 ( .A(p_input[6159]), .Z(n15712) );
  XOR U15749 ( .A(n16039), .B(n16040), .Z(n16035) );
  AND U15750 ( .A(n16041), .B(n16042), .Z(n16040) );
  XNOR U15751 ( .A(p_input[6190]), .B(n16039), .Z(n16042) );
  XNOR U15752 ( .A(n16039), .B(n15721), .Z(n16041) );
  IV U15753 ( .A(p_input[6158]), .Z(n15721) );
  XOR U15754 ( .A(n16043), .B(n16044), .Z(n16039) );
  AND U15755 ( .A(n16045), .B(n16046), .Z(n16044) );
  XNOR U15756 ( .A(p_input[6189]), .B(n16043), .Z(n16046) );
  XNOR U15757 ( .A(n16043), .B(n15730), .Z(n16045) );
  IV U15758 ( .A(p_input[6157]), .Z(n15730) );
  XOR U15759 ( .A(n16047), .B(n16048), .Z(n16043) );
  AND U15760 ( .A(n16049), .B(n16050), .Z(n16048) );
  XNOR U15761 ( .A(p_input[6188]), .B(n16047), .Z(n16050) );
  XNOR U15762 ( .A(n16047), .B(n15739), .Z(n16049) );
  IV U15763 ( .A(p_input[6156]), .Z(n15739) );
  XOR U15764 ( .A(n16051), .B(n16052), .Z(n16047) );
  AND U15765 ( .A(n16053), .B(n16054), .Z(n16052) );
  XNOR U15766 ( .A(p_input[6187]), .B(n16051), .Z(n16054) );
  XNOR U15767 ( .A(n16051), .B(n15748), .Z(n16053) );
  IV U15768 ( .A(p_input[6155]), .Z(n15748) );
  XOR U15769 ( .A(n16055), .B(n16056), .Z(n16051) );
  AND U15770 ( .A(n16057), .B(n16058), .Z(n16056) );
  XNOR U15771 ( .A(p_input[6186]), .B(n16055), .Z(n16058) );
  XNOR U15772 ( .A(n16055), .B(n15757), .Z(n16057) );
  IV U15773 ( .A(p_input[6154]), .Z(n15757) );
  XOR U15774 ( .A(n16059), .B(n16060), .Z(n16055) );
  AND U15775 ( .A(n16061), .B(n16062), .Z(n16060) );
  XNOR U15776 ( .A(p_input[6185]), .B(n16059), .Z(n16062) );
  XNOR U15777 ( .A(n16059), .B(n15766), .Z(n16061) );
  IV U15778 ( .A(p_input[6153]), .Z(n15766) );
  XOR U15779 ( .A(n16063), .B(n16064), .Z(n16059) );
  AND U15780 ( .A(n16065), .B(n16066), .Z(n16064) );
  XNOR U15781 ( .A(p_input[6184]), .B(n16063), .Z(n16066) );
  XNOR U15782 ( .A(n16063), .B(n15775), .Z(n16065) );
  IV U15783 ( .A(p_input[6152]), .Z(n15775) );
  XOR U15784 ( .A(n16067), .B(n16068), .Z(n16063) );
  AND U15785 ( .A(n16069), .B(n16070), .Z(n16068) );
  XNOR U15786 ( .A(p_input[6183]), .B(n16067), .Z(n16070) );
  XNOR U15787 ( .A(n16067), .B(n15784), .Z(n16069) );
  IV U15788 ( .A(p_input[6151]), .Z(n15784) );
  XOR U15789 ( .A(n16071), .B(n16072), .Z(n16067) );
  AND U15790 ( .A(n16073), .B(n16074), .Z(n16072) );
  XNOR U15791 ( .A(p_input[6182]), .B(n16071), .Z(n16074) );
  XNOR U15792 ( .A(n16071), .B(n15793), .Z(n16073) );
  IV U15793 ( .A(p_input[6150]), .Z(n15793) );
  XOR U15794 ( .A(n16075), .B(n16076), .Z(n16071) );
  AND U15795 ( .A(n16077), .B(n16078), .Z(n16076) );
  XNOR U15796 ( .A(p_input[6181]), .B(n16075), .Z(n16078) );
  XNOR U15797 ( .A(n16075), .B(n15802), .Z(n16077) );
  IV U15798 ( .A(p_input[6149]), .Z(n15802) );
  XOR U15799 ( .A(n16079), .B(n16080), .Z(n16075) );
  AND U15800 ( .A(n16081), .B(n16082), .Z(n16080) );
  XNOR U15801 ( .A(p_input[6180]), .B(n16079), .Z(n16082) );
  XNOR U15802 ( .A(n16079), .B(n15811), .Z(n16081) );
  IV U15803 ( .A(p_input[6148]), .Z(n15811) );
  XOR U15804 ( .A(n16083), .B(n16084), .Z(n16079) );
  AND U15805 ( .A(n16085), .B(n16086), .Z(n16084) );
  XNOR U15806 ( .A(p_input[6179]), .B(n16083), .Z(n16086) );
  XNOR U15807 ( .A(n16083), .B(n15820), .Z(n16085) );
  IV U15808 ( .A(p_input[6147]), .Z(n15820) );
  XOR U15809 ( .A(n16087), .B(n16088), .Z(n16083) );
  AND U15810 ( .A(n16089), .B(n16090), .Z(n16088) );
  XNOR U15811 ( .A(p_input[6178]), .B(n16087), .Z(n16090) );
  XNOR U15812 ( .A(n16087), .B(n15829), .Z(n16089) );
  IV U15813 ( .A(p_input[6146]), .Z(n15829) );
  XNOR U15814 ( .A(n16091), .B(n16092), .Z(n16087) );
  AND U15815 ( .A(n16093), .B(n16094), .Z(n16092) );
  XOR U15816 ( .A(p_input[6177]), .B(n16091), .Z(n16094) );
  XNOR U15817 ( .A(p_input[6145]), .B(n16091), .Z(n16093) );
  AND U15818 ( .A(p_input[6176]), .B(n16095), .Z(n16091) );
  IV U15819 ( .A(p_input[6144]), .Z(n16095) );
  XOR U15820 ( .A(n16096), .B(n16097), .Z(n1520) );
  AND U15821 ( .A(n1125), .B(n16098), .Z(n16097) );
  XNOR U15822 ( .A(n16099), .B(n16096), .Z(n16098) );
  XOR U15823 ( .A(n16100), .B(n16101), .Z(n1125) );
  AND U15824 ( .A(n16102), .B(n16103), .Z(n16101) );
  XOR U15825 ( .A(n16100), .B(n1535), .Z(n16103) );
  XOR U15826 ( .A(n16104), .B(n16105), .Z(n1535) );
  AND U15827 ( .A(n1091), .B(n16106), .Z(n16105) );
  XOR U15828 ( .A(n16107), .B(n16104), .Z(n16106) );
  XNOR U15829 ( .A(n1532), .B(n16100), .Z(n16102) );
  XOR U15830 ( .A(n16108), .B(n16109), .Z(n1532) );
  AND U15831 ( .A(n1088), .B(n16110), .Z(n16109) );
  XOR U15832 ( .A(n16111), .B(n16108), .Z(n16110) );
  XOR U15833 ( .A(n16112), .B(n16113), .Z(n16100) );
  AND U15834 ( .A(n16114), .B(n16115), .Z(n16113) );
  XOR U15835 ( .A(n16112), .B(n1547), .Z(n16115) );
  XOR U15836 ( .A(n16116), .B(n16117), .Z(n1547) );
  AND U15837 ( .A(n1091), .B(n16118), .Z(n16117) );
  XOR U15838 ( .A(n16119), .B(n16116), .Z(n16118) );
  XNOR U15839 ( .A(n1544), .B(n16112), .Z(n16114) );
  XOR U15840 ( .A(n16120), .B(n16121), .Z(n1544) );
  AND U15841 ( .A(n1088), .B(n16122), .Z(n16121) );
  XOR U15842 ( .A(n16123), .B(n16120), .Z(n16122) );
  XOR U15843 ( .A(n16124), .B(n16125), .Z(n16112) );
  AND U15844 ( .A(n16126), .B(n16127), .Z(n16125) );
  XOR U15845 ( .A(n16124), .B(n1559), .Z(n16127) );
  XOR U15846 ( .A(n16128), .B(n16129), .Z(n1559) );
  AND U15847 ( .A(n1091), .B(n16130), .Z(n16129) );
  XOR U15848 ( .A(n16131), .B(n16128), .Z(n16130) );
  XNOR U15849 ( .A(n1556), .B(n16124), .Z(n16126) );
  XOR U15850 ( .A(n16132), .B(n16133), .Z(n1556) );
  AND U15851 ( .A(n1088), .B(n16134), .Z(n16133) );
  XOR U15852 ( .A(n16135), .B(n16132), .Z(n16134) );
  XOR U15853 ( .A(n16136), .B(n16137), .Z(n16124) );
  AND U15854 ( .A(n16138), .B(n16139), .Z(n16137) );
  XOR U15855 ( .A(n16136), .B(n1571), .Z(n16139) );
  XOR U15856 ( .A(n16140), .B(n16141), .Z(n1571) );
  AND U15857 ( .A(n1091), .B(n16142), .Z(n16141) );
  XOR U15858 ( .A(n16143), .B(n16140), .Z(n16142) );
  XNOR U15859 ( .A(n1568), .B(n16136), .Z(n16138) );
  XOR U15860 ( .A(n16144), .B(n16145), .Z(n1568) );
  AND U15861 ( .A(n1088), .B(n16146), .Z(n16145) );
  XOR U15862 ( .A(n16147), .B(n16144), .Z(n16146) );
  XOR U15863 ( .A(n16148), .B(n16149), .Z(n16136) );
  AND U15864 ( .A(n16150), .B(n16151), .Z(n16149) );
  XOR U15865 ( .A(n16148), .B(n1583), .Z(n16151) );
  XOR U15866 ( .A(n16152), .B(n16153), .Z(n1583) );
  AND U15867 ( .A(n1091), .B(n16154), .Z(n16153) );
  XOR U15868 ( .A(n16155), .B(n16152), .Z(n16154) );
  XNOR U15869 ( .A(n1580), .B(n16148), .Z(n16150) );
  XOR U15870 ( .A(n16156), .B(n16157), .Z(n1580) );
  AND U15871 ( .A(n1088), .B(n16158), .Z(n16157) );
  XOR U15872 ( .A(n16159), .B(n16156), .Z(n16158) );
  XOR U15873 ( .A(n16160), .B(n16161), .Z(n16148) );
  AND U15874 ( .A(n16162), .B(n16163), .Z(n16161) );
  XOR U15875 ( .A(n16160), .B(n1595), .Z(n16163) );
  XOR U15876 ( .A(n16164), .B(n16165), .Z(n1595) );
  AND U15877 ( .A(n1091), .B(n16166), .Z(n16165) );
  XOR U15878 ( .A(n16167), .B(n16164), .Z(n16166) );
  XNOR U15879 ( .A(n1592), .B(n16160), .Z(n16162) );
  XOR U15880 ( .A(n16168), .B(n16169), .Z(n1592) );
  AND U15881 ( .A(n1088), .B(n16170), .Z(n16169) );
  XOR U15882 ( .A(n16171), .B(n16168), .Z(n16170) );
  XOR U15883 ( .A(n16172), .B(n16173), .Z(n16160) );
  AND U15884 ( .A(n16174), .B(n16175), .Z(n16173) );
  XOR U15885 ( .A(n16172), .B(n1607), .Z(n16175) );
  XOR U15886 ( .A(n16176), .B(n16177), .Z(n1607) );
  AND U15887 ( .A(n1091), .B(n16178), .Z(n16177) );
  XOR U15888 ( .A(n16179), .B(n16176), .Z(n16178) );
  XNOR U15889 ( .A(n1604), .B(n16172), .Z(n16174) );
  XOR U15890 ( .A(n16180), .B(n16181), .Z(n1604) );
  AND U15891 ( .A(n1088), .B(n16182), .Z(n16181) );
  XOR U15892 ( .A(n16183), .B(n16180), .Z(n16182) );
  XOR U15893 ( .A(n16184), .B(n16185), .Z(n16172) );
  AND U15894 ( .A(n16186), .B(n16187), .Z(n16185) );
  XOR U15895 ( .A(n16184), .B(n1619), .Z(n16187) );
  XOR U15896 ( .A(n16188), .B(n16189), .Z(n1619) );
  AND U15897 ( .A(n1091), .B(n16190), .Z(n16189) );
  XOR U15898 ( .A(n16191), .B(n16188), .Z(n16190) );
  XNOR U15899 ( .A(n1616), .B(n16184), .Z(n16186) );
  XOR U15900 ( .A(n16192), .B(n16193), .Z(n1616) );
  AND U15901 ( .A(n1088), .B(n16194), .Z(n16193) );
  XOR U15902 ( .A(n16195), .B(n16192), .Z(n16194) );
  XOR U15903 ( .A(n16196), .B(n16197), .Z(n16184) );
  AND U15904 ( .A(n16198), .B(n16199), .Z(n16197) );
  XOR U15905 ( .A(n16196), .B(n1631), .Z(n16199) );
  XOR U15906 ( .A(n16200), .B(n16201), .Z(n1631) );
  AND U15907 ( .A(n1091), .B(n16202), .Z(n16201) );
  XOR U15908 ( .A(n16203), .B(n16200), .Z(n16202) );
  XNOR U15909 ( .A(n1628), .B(n16196), .Z(n16198) );
  XOR U15910 ( .A(n16204), .B(n16205), .Z(n1628) );
  AND U15911 ( .A(n1088), .B(n16206), .Z(n16205) );
  XOR U15912 ( .A(n16207), .B(n16204), .Z(n16206) );
  XOR U15913 ( .A(n16208), .B(n16209), .Z(n16196) );
  AND U15914 ( .A(n16210), .B(n16211), .Z(n16209) );
  XOR U15915 ( .A(n16208), .B(n1643), .Z(n16211) );
  XOR U15916 ( .A(n16212), .B(n16213), .Z(n1643) );
  AND U15917 ( .A(n1091), .B(n16214), .Z(n16213) );
  XOR U15918 ( .A(n16215), .B(n16212), .Z(n16214) );
  XNOR U15919 ( .A(n1640), .B(n16208), .Z(n16210) );
  XOR U15920 ( .A(n16216), .B(n16217), .Z(n1640) );
  AND U15921 ( .A(n1088), .B(n16218), .Z(n16217) );
  XOR U15922 ( .A(n16219), .B(n16216), .Z(n16218) );
  XOR U15923 ( .A(n16220), .B(n16221), .Z(n16208) );
  AND U15924 ( .A(n16222), .B(n16223), .Z(n16221) );
  XOR U15925 ( .A(n16220), .B(n1655), .Z(n16223) );
  XOR U15926 ( .A(n16224), .B(n16225), .Z(n1655) );
  AND U15927 ( .A(n1091), .B(n16226), .Z(n16225) );
  XOR U15928 ( .A(n16227), .B(n16224), .Z(n16226) );
  XNOR U15929 ( .A(n1652), .B(n16220), .Z(n16222) );
  XOR U15930 ( .A(n16228), .B(n16229), .Z(n1652) );
  AND U15931 ( .A(n1088), .B(n16230), .Z(n16229) );
  XOR U15932 ( .A(n16231), .B(n16228), .Z(n16230) );
  XOR U15933 ( .A(n16232), .B(n16233), .Z(n16220) );
  AND U15934 ( .A(n16234), .B(n16235), .Z(n16233) );
  XOR U15935 ( .A(n16232), .B(n1667), .Z(n16235) );
  XOR U15936 ( .A(n16236), .B(n16237), .Z(n1667) );
  AND U15937 ( .A(n1091), .B(n16238), .Z(n16237) );
  XOR U15938 ( .A(n16239), .B(n16236), .Z(n16238) );
  XNOR U15939 ( .A(n1664), .B(n16232), .Z(n16234) );
  XOR U15940 ( .A(n16240), .B(n16241), .Z(n1664) );
  AND U15941 ( .A(n1088), .B(n16242), .Z(n16241) );
  XOR U15942 ( .A(n16243), .B(n16240), .Z(n16242) );
  XOR U15943 ( .A(n16244), .B(n16245), .Z(n16232) );
  AND U15944 ( .A(n16246), .B(n16247), .Z(n16245) );
  XOR U15945 ( .A(n16244), .B(n1679), .Z(n16247) );
  XOR U15946 ( .A(n16248), .B(n16249), .Z(n1679) );
  AND U15947 ( .A(n1091), .B(n16250), .Z(n16249) );
  XOR U15948 ( .A(n16251), .B(n16248), .Z(n16250) );
  XNOR U15949 ( .A(n1676), .B(n16244), .Z(n16246) );
  XOR U15950 ( .A(n16252), .B(n16253), .Z(n1676) );
  AND U15951 ( .A(n1088), .B(n16254), .Z(n16253) );
  XOR U15952 ( .A(n16255), .B(n16252), .Z(n16254) );
  XOR U15953 ( .A(n16256), .B(n16257), .Z(n16244) );
  AND U15954 ( .A(n16258), .B(n16259), .Z(n16257) );
  XOR U15955 ( .A(n16256), .B(n1691), .Z(n16259) );
  XOR U15956 ( .A(n16260), .B(n16261), .Z(n1691) );
  AND U15957 ( .A(n1091), .B(n16262), .Z(n16261) );
  XOR U15958 ( .A(n16263), .B(n16260), .Z(n16262) );
  XNOR U15959 ( .A(n1688), .B(n16256), .Z(n16258) );
  XOR U15960 ( .A(n16264), .B(n16265), .Z(n1688) );
  AND U15961 ( .A(n1088), .B(n16266), .Z(n16265) );
  XOR U15962 ( .A(n16267), .B(n16264), .Z(n16266) );
  XOR U15963 ( .A(n16268), .B(n16269), .Z(n16256) );
  AND U15964 ( .A(n16270), .B(n16271), .Z(n16269) );
  XOR U15965 ( .A(n16268), .B(n1703), .Z(n16271) );
  XOR U15966 ( .A(n16272), .B(n16273), .Z(n1703) );
  AND U15967 ( .A(n1091), .B(n16274), .Z(n16273) );
  XOR U15968 ( .A(n16275), .B(n16272), .Z(n16274) );
  XNOR U15969 ( .A(n1700), .B(n16268), .Z(n16270) );
  XOR U15970 ( .A(n16276), .B(n16277), .Z(n1700) );
  AND U15971 ( .A(n1088), .B(n16278), .Z(n16277) );
  XOR U15972 ( .A(n16279), .B(n16276), .Z(n16278) );
  XOR U15973 ( .A(n16280), .B(n16281), .Z(n16268) );
  AND U15974 ( .A(n16282), .B(n16283), .Z(n16281) );
  XOR U15975 ( .A(n16280), .B(n1715), .Z(n16283) );
  XOR U15976 ( .A(n16284), .B(n16285), .Z(n1715) );
  AND U15977 ( .A(n1091), .B(n16286), .Z(n16285) );
  XOR U15978 ( .A(n16287), .B(n16284), .Z(n16286) );
  XNOR U15979 ( .A(n1712), .B(n16280), .Z(n16282) );
  XOR U15980 ( .A(n16288), .B(n16289), .Z(n1712) );
  AND U15981 ( .A(n1088), .B(n16290), .Z(n16289) );
  XOR U15982 ( .A(n16291), .B(n16288), .Z(n16290) );
  XOR U15983 ( .A(n16292), .B(n16293), .Z(n16280) );
  AND U15984 ( .A(n16294), .B(n16295), .Z(n16293) );
  XOR U15985 ( .A(n16292), .B(n1727), .Z(n16295) );
  XOR U15986 ( .A(n16296), .B(n16297), .Z(n1727) );
  AND U15987 ( .A(n1091), .B(n16298), .Z(n16297) );
  XOR U15988 ( .A(n16299), .B(n16296), .Z(n16298) );
  XNOR U15989 ( .A(n1724), .B(n16292), .Z(n16294) );
  XOR U15990 ( .A(n16300), .B(n16301), .Z(n1724) );
  AND U15991 ( .A(n1088), .B(n16302), .Z(n16301) );
  XOR U15992 ( .A(n16303), .B(n16300), .Z(n16302) );
  XOR U15993 ( .A(n16304), .B(n16305), .Z(n16292) );
  AND U15994 ( .A(n16306), .B(n16307), .Z(n16305) );
  XOR U15995 ( .A(n16304), .B(n1739), .Z(n16307) );
  XOR U15996 ( .A(n16308), .B(n16309), .Z(n1739) );
  AND U15997 ( .A(n1091), .B(n16310), .Z(n16309) );
  XOR U15998 ( .A(n16311), .B(n16308), .Z(n16310) );
  XNOR U15999 ( .A(n1736), .B(n16304), .Z(n16306) );
  XOR U16000 ( .A(n16312), .B(n16313), .Z(n1736) );
  AND U16001 ( .A(n1088), .B(n16314), .Z(n16313) );
  XOR U16002 ( .A(n16315), .B(n16312), .Z(n16314) );
  XOR U16003 ( .A(n16316), .B(n16317), .Z(n16304) );
  AND U16004 ( .A(n16318), .B(n16319), .Z(n16317) );
  XOR U16005 ( .A(n16316), .B(n1751), .Z(n16319) );
  XOR U16006 ( .A(n16320), .B(n16321), .Z(n1751) );
  AND U16007 ( .A(n1091), .B(n16322), .Z(n16321) );
  XOR U16008 ( .A(n16323), .B(n16320), .Z(n16322) );
  XNOR U16009 ( .A(n1748), .B(n16316), .Z(n16318) );
  XOR U16010 ( .A(n16324), .B(n16325), .Z(n1748) );
  AND U16011 ( .A(n1088), .B(n16326), .Z(n16325) );
  XOR U16012 ( .A(n16327), .B(n16324), .Z(n16326) );
  XOR U16013 ( .A(n16328), .B(n16329), .Z(n16316) );
  AND U16014 ( .A(n16330), .B(n16331), .Z(n16329) );
  XOR U16015 ( .A(n16328), .B(n1763), .Z(n16331) );
  XOR U16016 ( .A(n16332), .B(n16333), .Z(n1763) );
  AND U16017 ( .A(n1091), .B(n16334), .Z(n16333) );
  XOR U16018 ( .A(n16335), .B(n16332), .Z(n16334) );
  XNOR U16019 ( .A(n1760), .B(n16328), .Z(n16330) );
  XOR U16020 ( .A(n16336), .B(n16337), .Z(n1760) );
  AND U16021 ( .A(n1088), .B(n16338), .Z(n16337) );
  XOR U16022 ( .A(n16339), .B(n16336), .Z(n16338) );
  XOR U16023 ( .A(n16340), .B(n16341), .Z(n16328) );
  AND U16024 ( .A(n16342), .B(n16343), .Z(n16341) );
  XOR U16025 ( .A(n16340), .B(n1775), .Z(n16343) );
  XOR U16026 ( .A(n16344), .B(n16345), .Z(n1775) );
  AND U16027 ( .A(n1091), .B(n16346), .Z(n16345) );
  XOR U16028 ( .A(n16347), .B(n16344), .Z(n16346) );
  XNOR U16029 ( .A(n1772), .B(n16340), .Z(n16342) );
  XOR U16030 ( .A(n16348), .B(n16349), .Z(n1772) );
  AND U16031 ( .A(n1088), .B(n16350), .Z(n16349) );
  XOR U16032 ( .A(n16351), .B(n16348), .Z(n16350) );
  XOR U16033 ( .A(n16352), .B(n16353), .Z(n16340) );
  AND U16034 ( .A(n16354), .B(n16355), .Z(n16353) );
  XOR U16035 ( .A(n16352), .B(n1787), .Z(n16355) );
  XOR U16036 ( .A(n16356), .B(n16357), .Z(n1787) );
  AND U16037 ( .A(n1091), .B(n16358), .Z(n16357) );
  XOR U16038 ( .A(n16359), .B(n16356), .Z(n16358) );
  XNOR U16039 ( .A(n1784), .B(n16352), .Z(n16354) );
  XOR U16040 ( .A(n16360), .B(n16361), .Z(n1784) );
  AND U16041 ( .A(n1088), .B(n16362), .Z(n16361) );
  XOR U16042 ( .A(n16363), .B(n16360), .Z(n16362) );
  XOR U16043 ( .A(n16364), .B(n16365), .Z(n16352) );
  AND U16044 ( .A(n16366), .B(n16367), .Z(n16365) );
  XOR U16045 ( .A(n16364), .B(n1799), .Z(n16367) );
  XOR U16046 ( .A(n16368), .B(n16369), .Z(n1799) );
  AND U16047 ( .A(n1091), .B(n16370), .Z(n16369) );
  XOR U16048 ( .A(n16371), .B(n16368), .Z(n16370) );
  XNOR U16049 ( .A(n1796), .B(n16364), .Z(n16366) );
  XOR U16050 ( .A(n16372), .B(n16373), .Z(n1796) );
  AND U16051 ( .A(n1088), .B(n16374), .Z(n16373) );
  XOR U16052 ( .A(n16375), .B(n16372), .Z(n16374) );
  XOR U16053 ( .A(n16376), .B(n16377), .Z(n16364) );
  AND U16054 ( .A(n16378), .B(n16379), .Z(n16377) );
  XOR U16055 ( .A(n16376), .B(n1811), .Z(n16379) );
  XOR U16056 ( .A(n16380), .B(n16381), .Z(n1811) );
  AND U16057 ( .A(n1091), .B(n16382), .Z(n16381) );
  XOR U16058 ( .A(n16383), .B(n16380), .Z(n16382) );
  XNOR U16059 ( .A(n1808), .B(n16376), .Z(n16378) );
  XOR U16060 ( .A(n16384), .B(n16385), .Z(n1808) );
  AND U16061 ( .A(n1088), .B(n16386), .Z(n16385) );
  XOR U16062 ( .A(n16387), .B(n16384), .Z(n16386) );
  XOR U16063 ( .A(n16388), .B(n16389), .Z(n16376) );
  AND U16064 ( .A(n16390), .B(n16391), .Z(n16389) );
  XOR U16065 ( .A(n16388), .B(n1823), .Z(n16391) );
  XOR U16066 ( .A(n16392), .B(n16393), .Z(n1823) );
  AND U16067 ( .A(n1091), .B(n16394), .Z(n16393) );
  XOR U16068 ( .A(n16395), .B(n16392), .Z(n16394) );
  XNOR U16069 ( .A(n1820), .B(n16388), .Z(n16390) );
  XOR U16070 ( .A(n16396), .B(n16397), .Z(n1820) );
  AND U16071 ( .A(n1088), .B(n16398), .Z(n16397) );
  XOR U16072 ( .A(n16399), .B(n16396), .Z(n16398) );
  XOR U16073 ( .A(n16400), .B(n16401), .Z(n16388) );
  AND U16074 ( .A(n16402), .B(n16403), .Z(n16401) );
  XOR U16075 ( .A(n16400), .B(n1835), .Z(n16403) );
  XOR U16076 ( .A(n16404), .B(n16405), .Z(n1835) );
  AND U16077 ( .A(n1091), .B(n16406), .Z(n16405) );
  XOR U16078 ( .A(n16407), .B(n16404), .Z(n16406) );
  XNOR U16079 ( .A(n1832), .B(n16400), .Z(n16402) );
  XOR U16080 ( .A(n16408), .B(n16409), .Z(n1832) );
  AND U16081 ( .A(n1088), .B(n16410), .Z(n16409) );
  XOR U16082 ( .A(n16411), .B(n16408), .Z(n16410) );
  XOR U16083 ( .A(n16412), .B(n16413), .Z(n16400) );
  AND U16084 ( .A(n16414), .B(n16415), .Z(n16413) );
  XOR U16085 ( .A(n16412), .B(n1847), .Z(n16415) );
  XOR U16086 ( .A(n16416), .B(n16417), .Z(n1847) );
  AND U16087 ( .A(n1091), .B(n16418), .Z(n16417) );
  XOR U16088 ( .A(n16419), .B(n16416), .Z(n16418) );
  XNOR U16089 ( .A(n1844), .B(n16412), .Z(n16414) );
  XOR U16090 ( .A(n16420), .B(n16421), .Z(n1844) );
  AND U16091 ( .A(n1088), .B(n16422), .Z(n16421) );
  XOR U16092 ( .A(n16423), .B(n16420), .Z(n16422) );
  XOR U16093 ( .A(n16424), .B(n16425), .Z(n16412) );
  AND U16094 ( .A(n16426), .B(n16427), .Z(n16425) );
  XOR U16095 ( .A(n16424), .B(n1859), .Z(n16427) );
  XOR U16096 ( .A(n16428), .B(n16429), .Z(n1859) );
  AND U16097 ( .A(n1091), .B(n16430), .Z(n16429) );
  XOR U16098 ( .A(n16431), .B(n16428), .Z(n16430) );
  XNOR U16099 ( .A(n1856), .B(n16424), .Z(n16426) );
  XOR U16100 ( .A(n16432), .B(n16433), .Z(n1856) );
  AND U16101 ( .A(n1088), .B(n16434), .Z(n16433) );
  XOR U16102 ( .A(n16435), .B(n16432), .Z(n16434) );
  XOR U16103 ( .A(n16436), .B(n16437), .Z(n16424) );
  AND U16104 ( .A(n16438), .B(n16439), .Z(n16437) );
  XOR U16105 ( .A(n16436), .B(n1871), .Z(n16439) );
  XOR U16106 ( .A(n16440), .B(n16441), .Z(n1871) );
  AND U16107 ( .A(n1091), .B(n16442), .Z(n16441) );
  XOR U16108 ( .A(n16443), .B(n16440), .Z(n16442) );
  XNOR U16109 ( .A(n1868), .B(n16436), .Z(n16438) );
  XOR U16110 ( .A(n16444), .B(n16445), .Z(n1868) );
  AND U16111 ( .A(n1088), .B(n16446), .Z(n16445) );
  XOR U16112 ( .A(n16447), .B(n16444), .Z(n16446) );
  XOR U16113 ( .A(n16448), .B(n16449), .Z(n16436) );
  AND U16114 ( .A(n16450), .B(n16451), .Z(n16449) );
  XOR U16115 ( .A(n16448), .B(n1883), .Z(n16451) );
  XOR U16116 ( .A(n16452), .B(n16453), .Z(n1883) );
  AND U16117 ( .A(n1091), .B(n16454), .Z(n16453) );
  XOR U16118 ( .A(n16455), .B(n16452), .Z(n16454) );
  XNOR U16119 ( .A(n1880), .B(n16448), .Z(n16450) );
  XOR U16120 ( .A(n16456), .B(n16457), .Z(n1880) );
  AND U16121 ( .A(n1088), .B(n16458), .Z(n16457) );
  XOR U16122 ( .A(n16459), .B(n16456), .Z(n16458) );
  XOR U16123 ( .A(n16460), .B(n16461), .Z(n16448) );
  AND U16124 ( .A(n16462), .B(n16463), .Z(n16461) );
  XNOR U16125 ( .A(n16464), .B(n1896), .Z(n16463) );
  XOR U16126 ( .A(n16465), .B(n16466), .Z(n1896) );
  AND U16127 ( .A(n1091), .B(n16467), .Z(n16466) );
  XOR U16128 ( .A(n16465), .B(n16468), .Z(n16467) );
  XNOR U16129 ( .A(n1893), .B(n16460), .Z(n16462) );
  XOR U16130 ( .A(n16469), .B(n16470), .Z(n1893) );
  AND U16131 ( .A(n1088), .B(n16471), .Z(n16470) );
  XOR U16132 ( .A(n16469), .B(n16472), .Z(n16471) );
  IV U16133 ( .A(n16464), .Z(n16460) );
  AND U16134 ( .A(n16096), .B(n16099), .Z(n16464) );
  XNOR U16135 ( .A(n16473), .B(n16474), .Z(n16099) );
  AND U16136 ( .A(n1091), .B(n16475), .Z(n16474) );
  XNOR U16137 ( .A(n16476), .B(n16473), .Z(n16475) );
  XOR U16138 ( .A(n16477), .B(n16478), .Z(n1091) );
  AND U16139 ( .A(n16479), .B(n16480), .Z(n16478) );
  XOR U16140 ( .A(n16477), .B(n16107), .Z(n16480) );
  XOR U16141 ( .A(n16481), .B(n16482), .Z(n16107) );
  AND U16142 ( .A(n1011), .B(n16483), .Z(n16482) );
  XOR U16143 ( .A(n16484), .B(n16481), .Z(n16483) );
  XNOR U16144 ( .A(n16104), .B(n16477), .Z(n16479) );
  XOR U16145 ( .A(n16485), .B(n16486), .Z(n16104) );
  AND U16146 ( .A(n1009), .B(n16487), .Z(n16486) );
  XOR U16147 ( .A(n16488), .B(n16485), .Z(n16487) );
  XOR U16148 ( .A(n16489), .B(n16490), .Z(n16477) );
  AND U16149 ( .A(n16491), .B(n16492), .Z(n16490) );
  XOR U16150 ( .A(n16489), .B(n16119), .Z(n16492) );
  XOR U16151 ( .A(n16493), .B(n16494), .Z(n16119) );
  AND U16152 ( .A(n1011), .B(n16495), .Z(n16494) );
  XOR U16153 ( .A(n16496), .B(n16493), .Z(n16495) );
  XNOR U16154 ( .A(n16116), .B(n16489), .Z(n16491) );
  XOR U16155 ( .A(n16497), .B(n16498), .Z(n16116) );
  AND U16156 ( .A(n1009), .B(n16499), .Z(n16498) );
  XOR U16157 ( .A(n16500), .B(n16497), .Z(n16499) );
  XOR U16158 ( .A(n16501), .B(n16502), .Z(n16489) );
  AND U16159 ( .A(n16503), .B(n16504), .Z(n16502) );
  XOR U16160 ( .A(n16501), .B(n16131), .Z(n16504) );
  XOR U16161 ( .A(n16505), .B(n16506), .Z(n16131) );
  AND U16162 ( .A(n1011), .B(n16507), .Z(n16506) );
  XOR U16163 ( .A(n16508), .B(n16505), .Z(n16507) );
  XNOR U16164 ( .A(n16128), .B(n16501), .Z(n16503) );
  XOR U16165 ( .A(n16509), .B(n16510), .Z(n16128) );
  AND U16166 ( .A(n1009), .B(n16511), .Z(n16510) );
  XOR U16167 ( .A(n16512), .B(n16509), .Z(n16511) );
  XOR U16168 ( .A(n16513), .B(n16514), .Z(n16501) );
  AND U16169 ( .A(n16515), .B(n16516), .Z(n16514) );
  XOR U16170 ( .A(n16513), .B(n16143), .Z(n16516) );
  XOR U16171 ( .A(n16517), .B(n16518), .Z(n16143) );
  AND U16172 ( .A(n1011), .B(n16519), .Z(n16518) );
  XOR U16173 ( .A(n16520), .B(n16517), .Z(n16519) );
  XNOR U16174 ( .A(n16140), .B(n16513), .Z(n16515) );
  XOR U16175 ( .A(n16521), .B(n16522), .Z(n16140) );
  AND U16176 ( .A(n1009), .B(n16523), .Z(n16522) );
  XOR U16177 ( .A(n16524), .B(n16521), .Z(n16523) );
  XOR U16178 ( .A(n16525), .B(n16526), .Z(n16513) );
  AND U16179 ( .A(n16527), .B(n16528), .Z(n16526) );
  XOR U16180 ( .A(n16525), .B(n16155), .Z(n16528) );
  XOR U16181 ( .A(n16529), .B(n16530), .Z(n16155) );
  AND U16182 ( .A(n1011), .B(n16531), .Z(n16530) );
  XOR U16183 ( .A(n16532), .B(n16529), .Z(n16531) );
  XNOR U16184 ( .A(n16152), .B(n16525), .Z(n16527) );
  XOR U16185 ( .A(n16533), .B(n16534), .Z(n16152) );
  AND U16186 ( .A(n1009), .B(n16535), .Z(n16534) );
  XOR U16187 ( .A(n16536), .B(n16533), .Z(n16535) );
  XOR U16188 ( .A(n16537), .B(n16538), .Z(n16525) );
  AND U16189 ( .A(n16539), .B(n16540), .Z(n16538) );
  XOR U16190 ( .A(n16537), .B(n16167), .Z(n16540) );
  XOR U16191 ( .A(n16541), .B(n16542), .Z(n16167) );
  AND U16192 ( .A(n1011), .B(n16543), .Z(n16542) );
  XOR U16193 ( .A(n16544), .B(n16541), .Z(n16543) );
  XNOR U16194 ( .A(n16164), .B(n16537), .Z(n16539) );
  XOR U16195 ( .A(n16545), .B(n16546), .Z(n16164) );
  AND U16196 ( .A(n1009), .B(n16547), .Z(n16546) );
  XOR U16197 ( .A(n16548), .B(n16545), .Z(n16547) );
  XOR U16198 ( .A(n16549), .B(n16550), .Z(n16537) );
  AND U16199 ( .A(n16551), .B(n16552), .Z(n16550) );
  XOR U16200 ( .A(n16549), .B(n16179), .Z(n16552) );
  XOR U16201 ( .A(n16553), .B(n16554), .Z(n16179) );
  AND U16202 ( .A(n1011), .B(n16555), .Z(n16554) );
  XOR U16203 ( .A(n16556), .B(n16553), .Z(n16555) );
  XNOR U16204 ( .A(n16176), .B(n16549), .Z(n16551) );
  XOR U16205 ( .A(n16557), .B(n16558), .Z(n16176) );
  AND U16206 ( .A(n1009), .B(n16559), .Z(n16558) );
  XOR U16207 ( .A(n16560), .B(n16557), .Z(n16559) );
  XOR U16208 ( .A(n16561), .B(n16562), .Z(n16549) );
  AND U16209 ( .A(n16563), .B(n16564), .Z(n16562) );
  XOR U16210 ( .A(n16561), .B(n16191), .Z(n16564) );
  XOR U16211 ( .A(n16565), .B(n16566), .Z(n16191) );
  AND U16212 ( .A(n1011), .B(n16567), .Z(n16566) );
  XOR U16213 ( .A(n16568), .B(n16565), .Z(n16567) );
  XNOR U16214 ( .A(n16188), .B(n16561), .Z(n16563) );
  XOR U16215 ( .A(n16569), .B(n16570), .Z(n16188) );
  AND U16216 ( .A(n1009), .B(n16571), .Z(n16570) );
  XOR U16217 ( .A(n16572), .B(n16569), .Z(n16571) );
  XOR U16218 ( .A(n16573), .B(n16574), .Z(n16561) );
  AND U16219 ( .A(n16575), .B(n16576), .Z(n16574) );
  XOR U16220 ( .A(n16573), .B(n16203), .Z(n16576) );
  XOR U16221 ( .A(n16577), .B(n16578), .Z(n16203) );
  AND U16222 ( .A(n1011), .B(n16579), .Z(n16578) );
  XOR U16223 ( .A(n16580), .B(n16577), .Z(n16579) );
  XNOR U16224 ( .A(n16200), .B(n16573), .Z(n16575) );
  XOR U16225 ( .A(n16581), .B(n16582), .Z(n16200) );
  AND U16226 ( .A(n1009), .B(n16583), .Z(n16582) );
  XOR U16227 ( .A(n16584), .B(n16581), .Z(n16583) );
  XOR U16228 ( .A(n16585), .B(n16586), .Z(n16573) );
  AND U16229 ( .A(n16587), .B(n16588), .Z(n16586) );
  XOR U16230 ( .A(n16585), .B(n16215), .Z(n16588) );
  XOR U16231 ( .A(n16589), .B(n16590), .Z(n16215) );
  AND U16232 ( .A(n1011), .B(n16591), .Z(n16590) );
  XOR U16233 ( .A(n16592), .B(n16589), .Z(n16591) );
  XNOR U16234 ( .A(n16212), .B(n16585), .Z(n16587) );
  XOR U16235 ( .A(n16593), .B(n16594), .Z(n16212) );
  AND U16236 ( .A(n1009), .B(n16595), .Z(n16594) );
  XOR U16237 ( .A(n16596), .B(n16593), .Z(n16595) );
  XOR U16238 ( .A(n16597), .B(n16598), .Z(n16585) );
  AND U16239 ( .A(n16599), .B(n16600), .Z(n16598) );
  XOR U16240 ( .A(n16597), .B(n16227), .Z(n16600) );
  XOR U16241 ( .A(n16601), .B(n16602), .Z(n16227) );
  AND U16242 ( .A(n1011), .B(n16603), .Z(n16602) );
  XOR U16243 ( .A(n16604), .B(n16601), .Z(n16603) );
  XNOR U16244 ( .A(n16224), .B(n16597), .Z(n16599) );
  XOR U16245 ( .A(n16605), .B(n16606), .Z(n16224) );
  AND U16246 ( .A(n1009), .B(n16607), .Z(n16606) );
  XOR U16247 ( .A(n16608), .B(n16605), .Z(n16607) );
  XOR U16248 ( .A(n16609), .B(n16610), .Z(n16597) );
  AND U16249 ( .A(n16611), .B(n16612), .Z(n16610) );
  XOR U16250 ( .A(n16609), .B(n16239), .Z(n16612) );
  XOR U16251 ( .A(n16613), .B(n16614), .Z(n16239) );
  AND U16252 ( .A(n1011), .B(n16615), .Z(n16614) );
  XOR U16253 ( .A(n16616), .B(n16613), .Z(n16615) );
  XNOR U16254 ( .A(n16236), .B(n16609), .Z(n16611) );
  XOR U16255 ( .A(n16617), .B(n16618), .Z(n16236) );
  AND U16256 ( .A(n1009), .B(n16619), .Z(n16618) );
  XOR U16257 ( .A(n16620), .B(n16617), .Z(n16619) );
  XOR U16258 ( .A(n16621), .B(n16622), .Z(n16609) );
  AND U16259 ( .A(n16623), .B(n16624), .Z(n16622) );
  XOR U16260 ( .A(n16621), .B(n16251), .Z(n16624) );
  XOR U16261 ( .A(n16625), .B(n16626), .Z(n16251) );
  AND U16262 ( .A(n1011), .B(n16627), .Z(n16626) );
  XOR U16263 ( .A(n16628), .B(n16625), .Z(n16627) );
  XNOR U16264 ( .A(n16248), .B(n16621), .Z(n16623) );
  XOR U16265 ( .A(n16629), .B(n16630), .Z(n16248) );
  AND U16266 ( .A(n1009), .B(n16631), .Z(n16630) );
  XOR U16267 ( .A(n16632), .B(n16629), .Z(n16631) );
  XOR U16268 ( .A(n16633), .B(n16634), .Z(n16621) );
  AND U16269 ( .A(n16635), .B(n16636), .Z(n16634) );
  XOR U16270 ( .A(n16633), .B(n16263), .Z(n16636) );
  XOR U16271 ( .A(n16637), .B(n16638), .Z(n16263) );
  AND U16272 ( .A(n1011), .B(n16639), .Z(n16638) );
  XOR U16273 ( .A(n16640), .B(n16637), .Z(n16639) );
  XNOR U16274 ( .A(n16260), .B(n16633), .Z(n16635) );
  XOR U16275 ( .A(n16641), .B(n16642), .Z(n16260) );
  AND U16276 ( .A(n1009), .B(n16643), .Z(n16642) );
  XOR U16277 ( .A(n16644), .B(n16641), .Z(n16643) );
  XOR U16278 ( .A(n16645), .B(n16646), .Z(n16633) );
  AND U16279 ( .A(n16647), .B(n16648), .Z(n16646) );
  XOR U16280 ( .A(n16645), .B(n16275), .Z(n16648) );
  XOR U16281 ( .A(n16649), .B(n16650), .Z(n16275) );
  AND U16282 ( .A(n1011), .B(n16651), .Z(n16650) );
  XOR U16283 ( .A(n16652), .B(n16649), .Z(n16651) );
  XNOR U16284 ( .A(n16272), .B(n16645), .Z(n16647) );
  XOR U16285 ( .A(n16653), .B(n16654), .Z(n16272) );
  AND U16286 ( .A(n1009), .B(n16655), .Z(n16654) );
  XOR U16287 ( .A(n16656), .B(n16653), .Z(n16655) );
  XOR U16288 ( .A(n16657), .B(n16658), .Z(n16645) );
  AND U16289 ( .A(n16659), .B(n16660), .Z(n16658) );
  XOR U16290 ( .A(n16657), .B(n16287), .Z(n16660) );
  XOR U16291 ( .A(n16661), .B(n16662), .Z(n16287) );
  AND U16292 ( .A(n1011), .B(n16663), .Z(n16662) );
  XOR U16293 ( .A(n16664), .B(n16661), .Z(n16663) );
  XNOR U16294 ( .A(n16284), .B(n16657), .Z(n16659) );
  XOR U16295 ( .A(n16665), .B(n16666), .Z(n16284) );
  AND U16296 ( .A(n1009), .B(n16667), .Z(n16666) );
  XOR U16297 ( .A(n16668), .B(n16665), .Z(n16667) );
  XOR U16298 ( .A(n16669), .B(n16670), .Z(n16657) );
  AND U16299 ( .A(n16671), .B(n16672), .Z(n16670) );
  XOR U16300 ( .A(n16669), .B(n16299), .Z(n16672) );
  XOR U16301 ( .A(n16673), .B(n16674), .Z(n16299) );
  AND U16302 ( .A(n1011), .B(n16675), .Z(n16674) );
  XOR U16303 ( .A(n16676), .B(n16673), .Z(n16675) );
  XNOR U16304 ( .A(n16296), .B(n16669), .Z(n16671) );
  XOR U16305 ( .A(n16677), .B(n16678), .Z(n16296) );
  AND U16306 ( .A(n1009), .B(n16679), .Z(n16678) );
  XOR U16307 ( .A(n16680), .B(n16677), .Z(n16679) );
  XOR U16308 ( .A(n16681), .B(n16682), .Z(n16669) );
  AND U16309 ( .A(n16683), .B(n16684), .Z(n16682) );
  XOR U16310 ( .A(n16681), .B(n16311), .Z(n16684) );
  XOR U16311 ( .A(n16685), .B(n16686), .Z(n16311) );
  AND U16312 ( .A(n1011), .B(n16687), .Z(n16686) );
  XOR U16313 ( .A(n16688), .B(n16685), .Z(n16687) );
  XNOR U16314 ( .A(n16308), .B(n16681), .Z(n16683) );
  XOR U16315 ( .A(n16689), .B(n16690), .Z(n16308) );
  AND U16316 ( .A(n1009), .B(n16691), .Z(n16690) );
  XOR U16317 ( .A(n16692), .B(n16689), .Z(n16691) );
  XOR U16318 ( .A(n16693), .B(n16694), .Z(n16681) );
  AND U16319 ( .A(n16695), .B(n16696), .Z(n16694) );
  XOR U16320 ( .A(n16693), .B(n16323), .Z(n16696) );
  XOR U16321 ( .A(n16697), .B(n16698), .Z(n16323) );
  AND U16322 ( .A(n1011), .B(n16699), .Z(n16698) );
  XOR U16323 ( .A(n16700), .B(n16697), .Z(n16699) );
  XNOR U16324 ( .A(n16320), .B(n16693), .Z(n16695) );
  XOR U16325 ( .A(n16701), .B(n16702), .Z(n16320) );
  AND U16326 ( .A(n1009), .B(n16703), .Z(n16702) );
  XOR U16327 ( .A(n16704), .B(n16701), .Z(n16703) );
  XOR U16328 ( .A(n16705), .B(n16706), .Z(n16693) );
  AND U16329 ( .A(n16707), .B(n16708), .Z(n16706) );
  XOR U16330 ( .A(n16705), .B(n16335), .Z(n16708) );
  XOR U16331 ( .A(n16709), .B(n16710), .Z(n16335) );
  AND U16332 ( .A(n1011), .B(n16711), .Z(n16710) );
  XOR U16333 ( .A(n16712), .B(n16709), .Z(n16711) );
  XNOR U16334 ( .A(n16332), .B(n16705), .Z(n16707) );
  XOR U16335 ( .A(n16713), .B(n16714), .Z(n16332) );
  AND U16336 ( .A(n1009), .B(n16715), .Z(n16714) );
  XOR U16337 ( .A(n16716), .B(n16713), .Z(n16715) );
  XOR U16338 ( .A(n16717), .B(n16718), .Z(n16705) );
  AND U16339 ( .A(n16719), .B(n16720), .Z(n16718) );
  XOR U16340 ( .A(n16717), .B(n16347), .Z(n16720) );
  XOR U16341 ( .A(n16721), .B(n16722), .Z(n16347) );
  AND U16342 ( .A(n1011), .B(n16723), .Z(n16722) );
  XOR U16343 ( .A(n16724), .B(n16721), .Z(n16723) );
  XNOR U16344 ( .A(n16344), .B(n16717), .Z(n16719) );
  XOR U16345 ( .A(n16725), .B(n16726), .Z(n16344) );
  AND U16346 ( .A(n1009), .B(n16727), .Z(n16726) );
  XOR U16347 ( .A(n16728), .B(n16725), .Z(n16727) );
  XOR U16348 ( .A(n16729), .B(n16730), .Z(n16717) );
  AND U16349 ( .A(n16731), .B(n16732), .Z(n16730) );
  XOR U16350 ( .A(n16729), .B(n16359), .Z(n16732) );
  XOR U16351 ( .A(n16733), .B(n16734), .Z(n16359) );
  AND U16352 ( .A(n1011), .B(n16735), .Z(n16734) );
  XOR U16353 ( .A(n16736), .B(n16733), .Z(n16735) );
  XNOR U16354 ( .A(n16356), .B(n16729), .Z(n16731) );
  XOR U16355 ( .A(n16737), .B(n16738), .Z(n16356) );
  AND U16356 ( .A(n1009), .B(n16739), .Z(n16738) );
  XOR U16357 ( .A(n16740), .B(n16737), .Z(n16739) );
  XOR U16358 ( .A(n16741), .B(n16742), .Z(n16729) );
  AND U16359 ( .A(n16743), .B(n16744), .Z(n16742) );
  XOR U16360 ( .A(n16741), .B(n16371), .Z(n16744) );
  XOR U16361 ( .A(n16745), .B(n16746), .Z(n16371) );
  AND U16362 ( .A(n1011), .B(n16747), .Z(n16746) );
  XOR U16363 ( .A(n16748), .B(n16745), .Z(n16747) );
  XNOR U16364 ( .A(n16368), .B(n16741), .Z(n16743) );
  XOR U16365 ( .A(n16749), .B(n16750), .Z(n16368) );
  AND U16366 ( .A(n1009), .B(n16751), .Z(n16750) );
  XOR U16367 ( .A(n16752), .B(n16749), .Z(n16751) );
  XOR U16368 ( .A(n16753), .B(n16754), .Z(n16741) );
  AND U16369 ( .A(n16755), .B(n16756), .Z(n16754) );
  XOR U16370 ( .A(n16753), .B(n16383), .Z(n16756) );
  XOR U16371 ( .A(n16757), .B(n16758), .Z(n16383) );
  AND U16372 ( .A(n1011), .B(n16759), .Z(n16758) );
  XOR U16373 ( .A(n16760), .B(n16757), .Z(n16759) );
  XNOR U16374 ( .A(n16380), .B(n16753), .Z(n16755) );
  XOR U16375 ( .A(n16761), .B(n16762), .Z(n16380) );
  AND U16376 ( .A(n1009), .B(n16763), .Z(n16762) );
  XOR U16377 ( .A(n16764), .B(n16761), .Z(n16763) );
  XOR U16378 ( .A(n16765), .B(n16766), .Z(n16753) );
  AND U16379 ( .A(n16767), .B(n16768), .Z(n16766) );
  XOR U16380 ( .A(n16765), .B(n16395), .Z(n16768) );
  XOR U16381 ( .A(n16769), .B(n16770), .Z(n16395) );
  AND U16382 ( .A(n1011), .B(n16771), .Z(n16770) );
  XOR U16383 ( .A(n16772), .B(n16769), .Z(n16771) );
  XNOR U16384 ( .A(n16392), .B(n16765), .Z(n16767) );
  XOR U16385 ( .A(n16773), .B(n16774), .Z(n16392) );
  AND U16386 ( .A(n1009), .B(n16775), .Z(n16774) );
  XOR U16387 ( .A(n16776), .B(n16773), .Z(n16775) );
  XOR U16388 ( .A(n16777), .B(n16778), .Z(n16765) );
  AND U16389 ( .A(n16779), .B(n16780), .Z(n16778) );
  XOR U16390 ( .A(n16777), .B(n16407), .Z(n16780) );
  XOR U16391 ( .A(n16781), .B(n16782), .Z(n16407) );
  AND U16392 ( .A(n1011), .B(n16783), .Z(n16782) );
  XOR U16393 ( .A(n16784), .B(n16781), .Z(n16783) );
  XNOR U16394 ( .A(n16404), .B(n16777), .Z(n16779) );
  XOR U16395 ( .A(n16785), .B(n16786), .Z(n16404) );
  AND U16396 ( .A(n1009), .B(n16787), .Z(n16786) );
  XOR U16397 ( .A(n16788), .B(n16785), .Z(n16787) );
  XOR U16398 ( .A(n16789), .B(n16790), .Z(n16777) );
  AND U16399 ( .A(n16791), .B(n16792), .Z(n16790) );
  XOR U16400 ( .A(n16789), .B(n16419), .Z(n16792) );
  XOR U16401 ( .A(n16793), .B(n16794), .Z(n16419) );
  AND U16402 ( .A(n1011), .B(n16795), .Z(n16794) );
  XOR U16403 ( .A(n16796), .B(n16793), .Z(n16795) );
  XNOR U16404 ( .A(n16416), .B(n16789), .Z(n16791) );
  XOR U16405 ( .A(n16797), .B(n16798), .Z(n16416) );
  AND U16406 ( .A(n1009), .B(n16799), .Z(n16798) );
  XOR U16407 ( .A(n16800), .B(n16797), .Z(n16799) );
  XOR U16408 ( .A(n16801), .B(n16802), .Z(n16789) );
  AND U16409 ( .A(n16803), .B(n16804), .Z(n16802) );
  XOR U16410 ( .A(n16801), .B(n16431), .Z(n16804) );
  XOR U16411 ( .A(n16805), .B(n16806), .Z(n16431) );
  AND U16412 ( .A(n1011), .B(n16807), .Z(n16806) );
  XOR U16413 ( .A(n16808), .B(n16805), .Z(n16807) );
  XNOR U16414 ( .A(n16428), .B(n16801), .Z(n16803) );
  XOR U16415 ( .A(n16809), .B(n16810), .Z(n16428) );
  AND U16416 ( .A(n1009), .B(n16811), .Z(n16810) );
  XOR U16417 ( .A(n16812), .B(n16809), .Z(n16811) );
  XOR U16418 ( .A(n16813), .B(n16814), .Z(n16801) );
  AND U16419 ( .A(n16815), .B(n16816), .Z(n16814) );
  XOR U16420 ( .A(n16813), .B(n16443), .Z(n16816) );
  XOR U16421 ( .A(n16817), .B(n16818), .Z(n16443) );
  AND U16422 ( .A(n1011), .B(n16819), .Z(n16818) );
  XOR U16423 ( .A(n16820), .B(n16817), .Z(n16819) );
  XNOR U16424 ( .A(n16440), .B(n16813), .Z(n16815) );
  XOR U16425 ( .A(n16821), .B(n16822), .Z(n16440) );
  AND U16426 ( .A(n1009), .B(n16823), .Z(n16822) );
  XOR U16427 ( .A(n16824), .B(n16821), .Z(n16823) );
  XOR U16428 ( .A(n16825), .B(n16826), .Z(n16813) );
  AND U16429 ( .A(n16827), .B(n16828), .Z(n16826) );
  XOR U16430 ( .A(n16825), .B(n16455), .Z(n16828) );
  XOR U16431 ( .A(n16829), .B(n16830), .Z(n16455) );
  AND U16432 ( .A(n1011), .B(n16831), .Z(n16830) );
  XOR U16433 ( .A(n16832), .B(n16829), .Z(n16831) );
  XNOR U16434 ( .A(n16452), .B(n16825), .Z(n16827) );
  XOR U16435 ( .A(n16833), .B(n16834), .Z(n16452) );
  AND U16436 ( .A(n1009), .B(n16835), .Z(n16834) );
  XOR U16437 ( .A(n16836), .B(n16833), .Z(n16835) );
  XOR U16438 ( .A(n16837), .B(n16838), .Z(n16825) );
  AND U16439 ( .A(n16839), .B(n16840), .Z(n16838) );
  XNOR U16440 ( .A(n16841), .B(n16468), .Z(n16840) );
  XOR U16441 ( .A(n16842), .B(n16843), .Z(n16468) );
  AND U16442 ( .A(n1011), .B(n16844), .Z(n16843) );
  XOR U16443 ( .A(n16842), .B(n16845), .Z(n16844) );
  XNOR U16444 ( .A(n16465), .B(n16837), .Z(n16839) );
  XOR U16445 ( .A(n16846), .B(n16847), .Z(n16465) );
  AND U16446 ( .A(n1009), .B(n16848), .Z(n16847) );
  XOR U16447 ( .A(n16846), .B(n16849), .Z(n16848) );
  IV U16448 ( .A(n16841), .Z(n16837) );
  AND U16449 ( .A(n16473), .B(n16476), .Z(n16841) );
  XNOR U16450 ( .A(n16850), .B(n16851), .Z(n16476) );
  AND U16451 ( .A(n1011), .B(n16852), .Z(n16851) );
  XNOR U16452 ( .A(n16853), .B(n16850), .Z(n16852) );
  XOR U16453 ( .A(n16854), .B(n16855), .Z(n1011) );
  AND U16454 ( .A(n16856), .B(n16857), .Z(n16855) );
  XOR U16455 ( .A(n16854), .B(n16484), .Z(n16857) );
  XOR U16456 ( .A(n16858), .B(n16859), .Z(n16484) );
  AND U16457 ( .A(n843), .B(n16860), .Z(n16859) );
  XOR U16458 ( .A(n16861), .B(n16858), .Z(n16860) );
  XNOR U16459 ( .A(n16481), .B(n16854), .Z(n16856) );
  XOR U16460 ( .A(n16862), .B(n16863), .Z(n16481) );
  AND U16461 ( .A(n841), .B(n16864), .Z(n16863) );
  XOR U16462 ( .A(n16865), .B(n16862), .Z(n16864) );
  XOR U16463 ( .A(n16866), .B(n16867), .Z(n16854) );
  AND U16464 ( .A(n16868), .B(n16869), .Z(n16867) );
  XOR U16465 ( .A(n16866), .B(n16496), .Z(n16869) );
  XOR U16466 ( .A(n16870), .B(n16871), .Z(n16496) );
  AND U16467 ( .A(n843), .B(n16872), .Z(n16871) );
  XOR U16468 ( .A(n16873), .B(n16870), .Z(n16872) );
  XNOR U16469 ( .A(n16493), .B(n16866), .Z(n16868) );
  XOR U16470 ( .A(n16874), .B(n16875), .Z(n16493) );
  AND U16471 ( .A(n841), .B(n16876), .Z(n16875) );
  XOR U16472 ( .A(n16877), .B(n16874), .Z(n16876) );
  XOR U16473 ( .A(n16878), .B(n16879), .Z(n16866) );
  AND U16474 ( .A(n16880), .B(n16881), .Z(n16879) );
  XOR U16475 ( .A(n16878), .B(n16508), .Z(n16881) );
  XOR U16476 ( .A(n16882), .B(n16883), .Z(n16508) );
  AND U16477 ( .A(n843), .B(n16884), .Z(n16883) );
  XOR U16478 ( .A(n16885), .B(n16882), .Z(n16884) );
  XNOR U16479 ( .A(n16505), .B(n16878), .Z(n16880) );
  XOR U16480 ( .A(n16886), .B(n16887), .Z(n16505) );
  AND U16481 ( .A(n841), .B(n16888), .Z(n16887) );
  XOR U16482 ( .A(n16889), .B(n16886), .Z(n16888) );
  XOR U16483 ( .A(n16890), .B(n16891), .Z(n16878) );
  AND U16484 ( .A(n16892), .B(n16893), .Z(n16891) );
  XOR U16485 ( .A(n16890), .B(n16520), .Z(n16893) );
  XOR U16486 ( .A(n16894), .B(n16895), .Z(n16520) );
  AND U16487 ( .A(n843), .B(n16896), .Z(n16895) );
  XOR U16488 ( .A(n16897), .B(n16894), .Z(n16896) );
  XNOR U16489 ( .A(n16517), .B(n16890), .Z(n16892) );
  XOR U16490 ( .A(n16898), .B(n16899), .Z(n16517) );
  AND U16491 ( .A(n841), .B(n16900), .Z(n16899) );
  XOR U16492 ( .A(n16901), .B(n16898), .Z(n16900) );
  XOR U16493 ( .A(n16902), .B(n16903), .Z(n16890) );
  AND U16494 ( .A(n16904), .B(n16905), .Z(n16903) );
  XOR U16495 ( .A(n16902), .B(n16532), .Z(n16905) );
  XOR U16496 ( .A(n16906), .B(n16907), .Z(n16532) );
  AND U16497 ( .A(n843), .B(n16908), .Z(n16907) );
  XOR U16498 ( .A(n16909), .B(n16906), .Z(n16908) );
  XNOR U16499 ( .A(n16529), .B(n16902), .Z(n16904) );
  XOR U16500 ( .A(n16910), .B(n16911), .Z(n16529) );
  AND U16501 ( .A(n841), .B(n16912), .Z(n16911) );
  XOR U16502 ( .A(n16913), .B(n16910), .Z(n16912) );
  XOR U16503 ( .A(n16914), .B(n16915), .Z(n16902) );
  AND U16504 ( .A(n16916), .B(n16917), .Z(n16915) );
  XOR U16505 ( .A(n16914), .B(n16544), .Z(n16917) );
  XOR U16506 ( .A(n16918), .B(n16919), .Z(n16544) );
  AND U16507 ( .A(n843), .B(n16920), .Z(n16919) );
  XOR U16508 ( .A(n16921), .B(n16918), .Z(n16920) );
  XNOR U16509 ( .A(n16541), .B(n16914), .Z(n16916) );
  XOR U16510 ( .A(n16922), .B(n16923), .Z(n16541) );
  AND U16511 ( .A(n841), .B(n16924), .Z(n16923) );
  XOR U16512 ( .A(n16925), .B(n16922), .Z(n16924) );
  XOR U16513 ( .A(n16926), .B(n16927), .Z(n16914) );
  AND U16514 ( .A(n16928), .B(n16929), .Z(n16927) );
  XOR U16515 ( .A(n16926), .B(n16556), .Z(n16929) );
  XOR U16516 ( .A(n16930), .B(n16931), .Z(n16556) );
  AND U16517 ( .A(n843), .B(n16932), .Z(n16931) );
  XOR U16518 ( .A(n16933), .B(n16930), .Z(n16932) );
  XNOR U16519 ( .A(n16553), .B(n16926), .Z(n16928) );
  XOR U16520 ( .A(n16934), .B(n16935), .Z(n16553) );
  AND U16521 ( .A(n841), .B(n16936), .Z(n16935) );
  XOR U16522 ( .A(n16937), .B(n16934), .Z(n16936) );
  XOR U16523 ( .A(n16938), .B(n16939), .Z(n16926) );
  AND U16524 ( .A(n16940), .B(n16941), .Z(n16939) );
  XOR U16525 ( .A(n16938), .B(n16568), .Z(n16941) );
  XOR U16526 ( .A(n16942), .B(n16943), .Z(n16568) );
  AND U16527 ( .A(n843), .B(n16944), .Z(n16943) );
  XOR U16528 ( .A(n16945), .B(n16942), .Z(n16944) );
  XNOR U16529 ( .A(n16565), .B(n16938), .Z(n16940) );
  XOR U16530 ( .A(n16946), .B(n16947), .Z(n16565) );
  AND U16531 ( .A(n841), .B(n16948), .Z(n16947) );
  XOR U16532 ( .A(n16949), .B(n16946), .Z(n16948) );
  XOR U16533 ( .A(n16950), .B(n16951), .Z(n16938) );
  AND U16534 ( .A(n16952), .B(n16953), .Z(n16951) );
  XOR U16535 ( .A(n16950), .B(n16580), .Z(n16953) );
  XOR U16536 ( .A(n16954), .B(n16955), .Z(n16580) );
  AND U16537 ( .A(n843), .B(n16956), .Z(n16955) );
  XOR U16538 ( .A(n16957), .B(n16954), .Z(n16956) );
  XNOR U16539 ( .A(n16577), .B(n16950), .Z(n16952) );
  XOR U16540 ( .A(n16958), .B(n16959), .Z(n16577) );
  AND U16541 ( .A(n841), .B(n16960), .Z(n16959) );
  XOR U16542 ( .A(n16961), .B(n16958), .Z(n16960) );
  XOR U16543 ( .A(n16962), .B(n16963), .Z(n16950) );
  AND U16544 ( .A(n16964), .B(n16965), .Z(n16963) );
  XOR U16545 ( .A(n16962), .B(n16592), .Z(n16965) );
  XOR U16546 ( .A(n16966), .B(n16967), .Z(n16592) );
  AND U16547 ( .A(n843), .B(n16968), .Z(n16967) );
  XOR U16548 ( .A(n16969), .B(n16966), .Z(n16968) );
  XNOR U16549 ( .A(n16589), .B(n16962), .Z(n16964) );
  XOR U16550 ( .A(n16970), .B(n16971), .Z(n16589) );
  AND U16551 ( .A(n841), .B(n16972), .Z(n16971) );
  XOR U16552 ( .A(n16973), .B(n16970), .Z(n16972) );
  XOR U16553 ( .A(n16974), .B(n16975), .Z(n16962) );
  AND U16554 ( .A(n16976), .B(n16977), .Z(n16975) );
  XOR U16555 ( .A(n16974), .B(n16604), .Z(n16977) );
  XOR U16556 ( .A(n16978), .B(n16979), .Z(n16604) );
  AND U16557 ( .A(n843), .B(n16980), .Z(n16979) );
  XOR U16558 ( .A(n16981), .B(n16978), .Z(n16980) );
  XNOR U16559 ( .A(n16601), .B(n16974), .Z(n16976) );
  XOR U16560 ( .A(n16982), .B(n16983), .Z(n16601) );
  AND U16561 ( .A(n841), .B(n16984), .Z(n16983) );
  XOR U16562 ( .A(n16985), .B(n16982), .Z(n16984) );
  XOR U16563 ( .A(n16986), .B(n16987), .Z(n16974) );
  AND U16564 ( .A(n16988), .B(n16989), .Z(n16987) );
  XOR U16565 ( .A(n16986), .B(n16616), .Z(n16989) );
  XOR U16566 ( .A(n16990), .B(n16991), .Z(n16616) );
  AND U16567 ( .A(n843), .B(n16992), .Z(n16991) );
  XOR U16568 ( .A(n16993), .B(n16990), .Z(n16992) );
  XNOR U16569 ( .A(n16613), .B(n16986), .Z(n16988) );
  XOR U16570 ( .A(n16994), .B(n16995), .Z(n16613) );
  AND U16571 ( .A(n841), .B(n16996), .Z(n16995) );
  XOR U16572 ( .A(n16997), .B(n16994), .Z(n16996) );
  XOR U16573 ( .A(n16998), .B(n16999), .Z(n16986) );
  AND U16574 ( .A(n17000), .B(n17001), .Z(n16999) );
  XOR U16575 ( .A(n16998), .B(n16628), .Z(n17001) );
  XOR U16576 ( .A(n17002), .B(n17003), .Z(n16628) );
  AND U16577 ( .A(n843), .B(n17004), .Z(n17003) );
  XOR U16578 ( .A(n17005), .B(n17002), .Z(n17004) );
  XNOR U16579 ( .A(n16625), .B(n16998), .Z(n17000) );
  XOR U16580 ( .A(n17006), .B(n17007), .Z(n16625) );
  AND U16581 ( .A(n841), .B(n17008), .Z(n17007) );
  XOR U16582 ( .A(n17009), .B(n17006), .Z(n17008) );
  XOR U16583 ( .A(n17010), .B(n17011), .Z(n16998) );
  AND U16584 ( .A(n17012), .B(n17013), .Z(n17011) );
  XOR U16585 ( .A(n17010), .B(n16640), .Z(n17013) );
  XOR U16586 ( .A(n17014), .B(n17015), .Z(n16640) );
  AND U16587 ( .A(n843), .B(n17016), .Z(n17015) );
  XOR U16588 ( .A(n17017), .B(n17014), .Z(n17016) );
  XNOR U16589 ( .A(n16637), .B(n17010), .Z(n17012) );
  XOR U16590 ( .A(n17018), .B(n17019), .Z(n16637) );
  AND U16591 ( .A(n841), .B(n17020), .Z(n17019) );
  XOR U16592 ( .A(n17021), .B(n17018), .Z(n17020) );
  XOR U16593 ( .A(n17022), .B(n17023), .Z(n17010) );
  AND U16594 ( .A(n17024), .B(n17025), .Z(n17023) );
  XOR U16595 ( .A(n17022), .B(n16652), .Z(n17025) );
  XOR U16596 ( .A(n17026), .B(n17027), .Z(n16652) );
  AND U16597 ( .A(n843), .B(n17028), .Z(n17027) );
  XOR U16598 ( .A(n17029), .B(n17026), .Z(n17028) );
  XNOR U16599 ( .A(n16649), .B(n17022), .Z(n17024) );
  XOR U16600 ( .A(n17030), .B(n17031), .Z(n16649) );
  AND U16601 ( .A(n841), .B(n17032), .Z(n17031) );
  XOR U16602 ( .A(n17033), .B(n17030), .Z(n17032) );
  XOR U16603 ( .A(n17034), .B(n17035), .Z(n17022) );
  AND U16604 ( .A(n17036), .B(n17037), .Z(n17035) );
  XOR U16605 ( .A(n17034), .B(n16664), .Z(n17037) );
  XOR U16606 ( .A(n17038), .B(n17039), .Z(n16664) );
  AND U16607 ( .A(n843), .B(n17040), .Z(n17039) );
  XOR U16608 ( .A(n17041), .B(n17038), .Z(n17040) );
  XNOR U16609 ( .A(n16661), .B(n17034), .Z(n17036) );
  XOR U16610 ( .A(n17042), .B(n17043), .Z(n16661) );
  AND U16611 ( .A(n841), .B(n17044), .Z(n17043) );
  XOR U16612 ( .A(n17045), .B(n17042), .Z(n17044) );
  XOR U16613 ( .A(n17046), .B(n17047), .Z(n17034) );
  AND U16614 ( .A(n17048), .B(n17049), .Z(n17047) );
  XOR U16615 ( .A(n17046), .B(n16676), .Z(n17049) );
  XOR U16616 ( .A(n17050), .B(n17051), .Z(n16676) );
  AND U16617 ( .A(n843), .B(n17052), .Z(n17051) );
  XOR U16618 ( .A(n17053), .B(n17050), .Z(n17052) );
  XNOR U16619 ( .A(n16673), .B(n17046), .Z(n17048) );
  XOR U16620 ( .A(n17054), .B(n17055), .Z(n16673) );
  AND U16621 ( .A(n841), .B(n17056), .Z(n17055) );
  XOR U16622 ( .A(n17057), .B(n17054), .Z(n17056) );
  XOR U16623 ( .A(n17058), .B(n17059), .Z(n17046) );
  AND U16624 ( .A(n17060), .B(n17061), .Z(n17059) );
  XOR U16625 ( .A(n17058), .B(n16688), .Z(n17061) );
  XOR U16626 ( .A(n17062), .B(n17063), .Z(n16688) );
  AND U16627 ( .A(n843), .B(n17064), .Z(n17063) );
  XOR U16628 ( .A(n17065), .B(n17062), .Z(n17064) );
  XNOR U16629 ( .A(n16685), .B(n17058), .Z(n17060) );
  XOR U16630 ( .A(n17066), .B(n17067), .Z(n16685) );
  AND U16631 ( .A(n841), .B(n17068), .Z(n17067) );
  XOR U16632 ( .A(n17069), .B(n17066), .Z(n17068) );
  XOR U16633 ( .A(n17070), .B(n17071), .Z(n17058) );
  AND U16634 ( .A(n17072), .B(n17073), .Z(n17071) );
  XOR U16635 ( .A(n17070), .B(n16700), .Z(n17073) );
  XOR U16636 ( .A(n17074), .B(n17075), .Z(n16700) );
  AND U16637 ( .A(n843), .B(n17076), .Z(n17075) );
  XOR U16638 ( .A(n17077), .B(n17074), .Z(n17076) );
  XNOR U16639 ( .A(n16697), .B(n17070), .Z(n17072) );
  XOR U16640 ( .A(n17078), .B(n17079), .Z(n16697) );
  AND U16641 ( .A(n841), .B(n17080), .Z(n17079) );
  XOR U16642 ( .A(n17081), .B(n17078), .Z(n17080) );
  XOR U16643 ( .A(n17082), .B(n17083), .Z(n17070) );
  AND U16644 ( .A(n17084), .B(n17085), .Z(n17083) );
  XOR U16645 ( .A(n17082), .B(n16712), .Z(n17085) );
  XOR U16646 ( .A(n17086), .B(n17087), .Z(n16712) );
  AND U16647 ( .A(n843), .B(n17088), .Z(n17087) );
  XOR U16648 ( .A(n17089), .B(n17086), .Z(n17088) );
  XNOR U16649 ( .A(n16709), .B(n17082), .Z(n17084) );
  XOR U16650 ( .A(n17090), .B(n17091), .Z(n16709) );
  AND U16651 ( .A(n841), .B(n17092), .Z(n17091) );
  XOR U16652 ( .A(n17093), .B(n17090), .Z(n17092) );
  XOR U16653 ( .A(n17094), .B(n17095), .Z(n17082) );
  AND U16654 ( .A(n17096), .B(n17097), .Z(n17095) );
  XOR U16655 ( .A(n17094), .B(n16724), .Z(n17097) );
  XOR U16656 ( .A(n17098), .B(n17099), .Z(n16724) );
  AND U16657 ( .A(n843), .B(n17100), .Z(n17099) );
  XOR U16658 ( .A(n17101), .B(n17098), .Z(n17100) );
  XNOR U16659 ( .A(n16721), .B(n17094), .Z(n17096) );
  XOR U16660 ( .A(n17102), .B(n17103), .Z(n16721) );
  AND U16661 ( .A(n841), .B(n17104), .Z(n17103) );
  XOR U16662 ( .A(n17105), .B(n17102), .Z(n17104) );
  XOR U16663 ( .A(n17106), .B(n17107), .Z(n17094) );
  AND U16664 ( .A(n17108), .B(n17109), .Z(n17107) );
  XOR U16665 ( .A(n17106), .B(n16736), .Z(n17109) );
  XOR U16666 ( .A(n17110), .B(n17111), .Z(n16736) );
  AND U16667 ( .A(n843), .B(n17112), .Z(n17111) );
  XOR U16668 ( .A(n17113), .B(n17110), .Z(n17112) );
  XNOR U16669 ( .A(n16733), .B(n17106), .Z(n17108) );
  XOR U16670 ( .A(n17114), .B(n17115), .Z(n16733) );
  AND U16671 ( .A(n841), .B(n17116), .Z(n17115) );
  XOR U16672 ( .A(n17117), .B(n17114), .Z(n17116) );
  XOR U16673 ( .A(n17118), .B(n17119), .Z(n17106) );
  AND U16674 ( .A(n17120), .B(n17121), .Z(n17119) );
  XOR U16675 ( .A(n17118), .B(n16748), .Z(n17121) );
  XOR U16676 ( .A(n17122), .B(n17123), .Z(n16748) );
  AND U16677 ( .A(n843), .B(n17124), .Z(n17123) );
  XOR U16678 ( .A(n17125), .B(n17122), .Z(n17124) );
  XNOR U16679 ( .A(n16745), .B(n17118), .Z(n17120) );
  XOR U16680 ( .A(n17126), .B(n17127), .Z(n16745) );
  AND U16681 ( .A(n841), .B(n17128), .Z(n17127) );
  XOR U16682 ( .A(n17129), .B(n17126), .Z(n17128) );
  XOR U16683 ( .A(n17130), .B(n17131), .Z(n17118) );
  AND U16684 ( .A(n17132), .B(n17133), .Z(n17131) );
  XOR U16685 ( .A(n17130), .B(n16760), .Z(n17133) );
  XOR U16686 ( .A(n17134), .B(n17135), .Z(n16760) );
  AND U16687 ( .A(n843), .B(n17136), .Z(n17135) );
  XOR U16688 ( .A(n17137), .B(n17134), .Z(n17136) );
  XNOR U16689 ( .A(n16757), .B(n17130), .Z(n17132) );
  XOR U16690 ( .A(n17138), .B(n17139), .Z(n16757) );
  AND U16691 ( .A(n841), .B(n17140), .Z(n17139) );
  XOR U16692 ( .A(n17141), .B(n17138), .Z(n17140) );
  XOR U16693 ( .A(n17142), .B(n17143), .Z(n17130) );
  AND U16694 ( .A(n17144), .B(n17145), .Z(n17143) );
  XOR U16695 ( .A(n17142), .B(n16772), .Z(n17145) );
  XOR U16696 ( .A(n17146), .B(n17147), .Z(n16772) );
  AND U16697 ( .A(n843), .B(n17148), .Z(n17147) );
  XOR U16698 ( .A(n17149), .B(n17146), .Z(n17148) );
  XNOR U16699 ( .A(n16769), .B(n17142), .Z(n17144) );
  XOR U16700 ( .A(n17150), .B(n17151), .Z(n16769) );
  AND U16701 ( .A(n841), .B(n17152), .Z(n17151) );
  XOR U16702 ( .A(n17153), .B(n17150), .Z(n17152) );
  XOR U16703 ( .A(n17154), .B(n17155), .Z(n17142) );
  AND U16704 ( .A(n17156), .B(n17157), .Z(n17155) );
  XOR U16705 ( .A(n17154), .B(n16784), .Z(n17157) );
  XOR U16706 ( .A(n17158), .B(n17159), .Z(n16784) );
  AND U16707 ( .A(n843), .B(n17160), .Z(n17159) );
  XOR U16708 ( .A(n17161), .B(n17158), .Z(n17160) );
  XNOR U16709 ( .A(n16781), .B(n17154), .Z(n17156) );
  XOR U16710 ( .A(n17162), .B(n17163), .Z(n16781) );
  AND U16711 ( .A(n841), .B(n17164), .Z(n17163) );
  XOR U16712 ( .A(n17165), .B(n17162), .Z(n17164) );
  XOR U16713 ( .A(n17166), .B(n17167), .Z(n17154) );
  AND U16714 ( .A(n17168), .B(n17169), .Z(n17167) );
  XOR U16715 ( .A(n17166), .B(n16796), .Z(n17169) );
  XOR U16716 ( .A(n17170), .B(n17171), .Z(n16796) );
  AND U16717 ( .A(n843), .B(n17172), .Z(n17171) );
  XOR U16718 ( .A(n17173), .B(n17170), .Z(n17172) );
  XNOR U16719 ( .A(n16793), .B(n17166), .Z(n17168) );
  XOR U16720 ( .A(n17174), .B(n17175), .Z(n16793) );
  AND U16721 ( .A(n841), .B(n17176), .Z(n17175) );
  XOR U16722 ( .A(n17177), .B(n17174), .Z(n17176) );
  XOR U16723 ( .A(n17178), .B(n17179), .Z(n17166) );
  AND U16724 ( .A(n17180), .B(n17181), .Z(n17179) );
  XOR U16725 ( .A(n17178), .B(n16808), .Z(n17181) );
  XOR U16726 ( .A(n17182), .B(n17183), .Z(n16808) );
  AND U16727 ( .A(n843), .B(n17184), .Z(n17183) );
  XOR U16728 ( .A(n17185), .B(n17182), .Z(n17184) );
  XNOR U16729 ( .A(n16805), .B(n17178), .Z(n17180) );
  XOR U16730 ( .A(n17186), .B(n17187), .Z(n16805) );
  AND U16731 ( .A(n841), .B(n17188), .Z(n17187) );
  XOR U16732 ( .A(n17189), .B(n17186), .Z(n17188) );
  XOR U16733 ( .A(n17190), .B(n17191), .Z(n17178) );
  AND U16734 ( .A(n17192), .B(n17193), .Z(n17191) );
  XOR U16735 ( .A(n17190), .B(n16820), .Z(n17193) );
  XOR U16736 ( .A(n17194), .B(n17195), .Z(n16820) );
  AND U16737 ( .A(n843), .B(n17196), .Z(n17195) );
  XOR U16738 ( .A(n17197), .B(n17194), .Z(n17196) );
  XNOR U16739 ( .A(n16817), .B(n17190), .Z(n17192) );
  XOR U16740 ( .A(n17198), .B(n17199), .Z(n16817) );
  AND U16741 ( .A(n841), .B(n17200), .Z(n17199) );
  XOR U16742 ( .A(n17201), .B(n17198), .Z(n17200) );
  XOR U16743 ( .A(n17202), .B(n17203), .Z(n17190) );
  AND U16744 ( .A(n17204), .B(n17205), .Z(n17203) );
  XOR U16745 ( .A(n17202), .B(n16832), .Z(n17205) );
  XOR U16746 ( .A(n17206), .B(n17207), .Z(n16832) );
  AND U16747 ( .A(n843), .B(n17208), .Z(n17207) );
  XOR U16748 ( .A(n17209), .B(n17206), .Z(n17208) );
  XNOR U16749 ( .A(n16829), .B(n17202), .Z(n17204) );
  XOR U16750 ( .A(n17210), .B(n17211), .Z(n16829) );
  AND U16751 ( .A(n841), .B(n17212), .Z(n17211) );
  XOR U16752 ( .A(n17213), .B(n17210), .Z(n17212) );
  XOR U16753 ( .A(n17214), .B(n17215), .Z(n17202) );
  AND U16754 ( .A(n17216), .B(n17217), .Z(n17215) );
  XNOR U16755 ( .A(n17218), .B(n16845), .Z(n17217) );
  XOR U16756 ( .A(n17219), .B(n17220), .Z(n16845) );
  AND U16757 ( .A(n843), .B(n17221), .Z(n17220) );
  XOR U16758 ( .A(n17219), .B(n17222), .Z(n17221) );
  XNOR U16759 ( .A(n16842), .B(n17214), .Z(n17216) );
  XOR U16760 ( .A(n17223), .B(n17224), .Z(n16842) );
  AND U16761 ( .A(n841), .B(n17225), .Z(n17224) );
  XOR U16762 ( .A(n17223), .B(n17226), .Z(n17225) );
  IV U16763 ( .A(n17218), .Z(n17214) );
  AND U16764 ( .A(n16850), .B(n16853), .Z(n17218) );
  XNOR U16765 ( .A(n17227), .B(n17228), .Z(n16853) );
  AND U16766 ( .A(n843), .B(n17229), .Z(n17228) );
  XNOR U16767 ( .A(n17230), .B(n17227), .Z(n17229) );
  XOR U16768 ( .A(n17231), .B(n17232), .Z(n843) );
  AND U16769 ( .A(n17233), .B(n17234), .Z(n17232) );
  XOR U16770 ( .A(n17231), .B(n16861), .Z(n17234) );
  XNOR U16771 ( .A(n17235), .B(n17236), .Z(n16861) );
  AND U16772 ( .A(n17237), .B(n499), .Z(n17236) );
  AND U16773 ( .A(n17235), .B(n17238), .Z(n17237) );
  XNOR U16774 ( .A(n16858), .B(n17231), .Z(n17233) );
  XOR U16775 ( .A(n17239), .B(n17240), .Z(n16858) );
  AND U16776 ( .A(n17241), .B(n497), .Z(n17240) );
  NOR U16777 ( .A(n17239), .B(n17242), .Z(n17241) );
  XOR U16778 ( .A(n17243), .B(n17244), .Z(n17231) );
  AND U16779 ( .A(n17245), .B(n17246), .Z(n17244) );
  XOR U16780 ( .A(n17243), .B(n16873), .Z(n17246) );
  XOR U16781 ( .A(n17247), .B(n17248), .Z(n16873) );
  AND U16782 ( .A(n499), .B(n17249), .Z(n17248) );
  XOR U16783 ( .A(n17250), .B(n17247), .Z(n17249) );
  XNOR U16784 ( .A(n16870), .B(n17243), .Z(n17245) );
  XOR U16785 ( .A(n17251), .B(n17252), .Z(n16870) );
  AND U16786 ( .A(n497), .B(n17253), .Z(n17252) );
  XOR U16787 ( .A(n17254), .B(n17251), .Z(n17253) );
  XOR U16788 ( .A(n17255), .B(n17256), .Z(n17243) );
  AND U16789 ( .A(n17257), .B(n17258), .Z(n17256) );
  XOR U16790 ( .A(n17255), .B(n16885), .Z(n17258) );
  XOR U16791 ( .A(n17259), .B(n17260), .Z(n16885) );
  AND U16792 ( .A(n499), .B(n17261), .Z(n17260) );
  XOR U16793 ( .A(n17262), .B(n17259), .Z(n17261) );
  XNOR U16794 ( .A(n16882), .B(n17255), .Z(n17257) );
  XOR U16795 ( .A(n17263), .B(n17264), .Z(n16882) );
  AND U16796 ( .A(n497), .B(n17265), .Z(n17264) );
  XOR U16797 ( .A(n17266), .B(n17263), .Z(n17265) );
  XOR U16798 ( .A(n17267), .B(n17268), .Z(n17255) );
  AND U16799 ( .A(n17269), .B(n17270), .Z(n17268) );
  XOR U16800 ( .A(n17267), .B(n16897), .Z(n17270) );
  XOR U16801 ( .A(n17271), .B(n17272), .Z(n16897) );
  AND U16802 ( .A(n499), .B(n17273), .Z(n17272) );
  XOR U16803 ( .A(n17274), .B(n17271), .Z(n17273) );
  XNOR U16804 ( .A(n16894), .B(n17267), .Z(n17269) );
  XOR U16805 ( .A(n17275), .B(n17276), .Z(n16894) );
  AND U16806 ( .A(n497), .B(n17277), .Z(n17276) );
  XOR U16807 ( .A(n17278), .B(n17275), .Z(n17277) );
  XOR U16808 ( .A(n17279), .B(n17280), .Z(n17267) );
  AND U16809 ( .A(n17281), .B(n17282), .Z(n17280) );
  XOR U16810 ( .A(n17279), .B(n16909), .Z(n17282) );
  XOR U16811 ( .A(n17283), .B(n17284), .Z(n16909) );
  AND U16812 ( .A(n499), .B(n17285), .Z(n17284) );
  XOR U16813 ( .A(n17286), .B(n17283), .Z(n17285) );
  XNOR U16814 ( .A(n16906), .B(n17279), .Z(n17281) );
  XOR U16815 ( .A(n17287), .B(n17288), .Z(n16906) );
  AND U16816 ( .A(n497), .B(n17289), .Z(n17288) );
  XOR U16817 ( .A(n17290), .B(n17287), .Z(n17289) );
  XOR U16818 ( .A(n17291), .B(n17292), .Z(n17279) );
  AND U16819 ( .A(n17293), .B(n17294), .Z(n17292) );
  XOR U16820 ( .A(n17291), .B(n16921), .Z(n17294) );
  XOR U16821 ( .A(n17295), .B(n17296), .Z(n16921) );
  AND U16822 ( .A(n499), .B(n17297), .Z(n17296) );
  XOR U16823 ( .A(n17298), .B(n17295), .Z(n17297) );
  XNOR U16824 ( .A(n16918), .B(n17291), .Z(n17293) );
  XOR U16825 ( .A(n17299), .B(n17300), .Z(n16918) );
  AND U16826 ( .A(n497), .B(n17301), .Z(n17300) );
  XOR U16827 ( .A(n17302), .B(n17299), .Z(n17301) );
  XOR U16828 ( .A(n17303), .B(n17304), .Z(n17291) );
  AND U16829 ( .A(n17305), .B(n17306), .Z(n17304) );
  XOR U16830 ( .A(n17303), .B(n16933), .Z(n17306) );
  XOR U16831 ( .A(n17307), .B(n17308), .Z(n16933) );
  AND U16832 ( .A(n499), .B(n17309), .Z(n17308) );
  XOR U16833 ( .A(n17310), .B(n17307), .Z(n17309) );
  XNOR U16834 ( .A(n16930), .B(n17303), .Z(n17305) );
  XOR U16835 ( .A(n17311), .B(n17312), .Z(n16930) );
  AND U16836 ( .A(n497), .B(n17313), .Z(n17312) );
  XOR U16837 ( .A(n17314), .B(n17311), .Z(n17313) );
  XOR U16838 ( .A(n17315), .B(n17316), .Z(n17303) );
  AND U16839 ( .A(n17317), .B(n17318), .Z(n17316) );
  XOR U16840 ( .A(n17315), .B(n16945), .Z(n17318) );
  XOR U16841 ( .A(n17319), .B(n17320), .Z(n16945) );
  AND U16842 ( .A(n499), .B(n17321), .Z(n17320) );
  XOR U16843 ( .A(n17322), .B(n17319), .Z(n17321) );
  XNOR U16844 ( .A(n16942), .B(n17315), .Z(n17317) );
  XOR U16845 ( .A(n17323), .B(n17324), .Z(n16942) );
  AND U16846 ( .A(n497), .B(n17325), .Z(n17324) );
  XOR U16847 ( .A(n17326), .B(n17323), .Z(n17325) );
  XOR U16848 ( .A(n17327), .B(n17328), .Z(n17315) );
  AND U16849 ( .A(n17329), .B(n17330), .Z(n17328) );
  XOR U16850 ( .A(n17327), .B(n16957), .Z(n17330) );
  XOR U16851 ( .A(n17331), .B(n17332), .Z(n16957) );
  AND U16852 ( .A(n499), .B(n17333), .Z(n17332) );
  XOR U16853 ( .A(n17334), .B(n17331), .Z(n17333) );
  XNOR U16854 ( .A(n16954), .B(n17327), .Z(n17329) );
  XOR U16855 ( .A(n17335), .B(n17336), .Z(n16954) );
  AND U16856 ( .A(n497), .B(n17337), .Z(n17336) );
  XOR U16857 ( .A(n17338), .B(n17335), .Z(n17337) );
  XOR U16858 ( .A(n17339), .B(n17340), .Z(n17327) );
  AND U16859 ( .A(n17341), .B(n17342), .Z(n17340) );
  XOR U16860 ( .A(n17339), .B(n16969), .Z(n17342) );
  XOR U16861 ( .A(n17343), .B(n17344), .Z(n16969) );
  AND U16862 ( .A(n499), .B(n17345), .Z(n17344) );
  XOR U16863 ( .A(n17346), .B(n17343), .Z(n17345) );
  XNOR U16864 ( .A(n16966), .B(n17339), .Z(n17341) );
  XOR U16865 ( .A(n17347), .B(n17348), .Z(n16966) );
  AND U16866 ( .A(n497), .B(n17349), .Z(n17348) );
  XOR U16867 ( .A(n17350), .B(n17347), .Z(n17349) );
  XOR U16868 ( .A(n17351), .B(n17352), .Z(n17339) );
  AND U16869 ( .A(n17353), .B(n17354), .Z(n17352) );
  XOR U16870 ( .A(n17351), .B(n16981), .Z(n17354) );
  XOR U16871 ( .A(n17355), .B(n17356), .Z(n16981) );
  AND U16872 ( .A(n499), .B(n17357), .Z(n17356) );
  XOR U16873 ( .A(n17358), .B(n17355), .Z(n17357) );
  XNOR U16874 ( .A(n16978), .B(n17351), .Z(n17353) );
  XOR U16875 ( .A(n17359), .B(n17360), .Z(n16978) );
  AND U16876 ( .A(n497), .B(n17361), .Z(n17360) );
  XOR U16877 ( .A(n17362), .B(n17359), .Z(n17361) );
  XOR U16878 ( .A(n17363), .B(n17364), .Z(n17351) );
  AND U16879 ( .A(n17365), .B(n17366), .Z(n17364) );
  XOR U16880 ( .A(n17363), .B(n16993), .Z(n17366) );
  XOR U16881 ( .A(n17367), .B(n17368), .Z(n16993) );
  AND U16882 ( .A(n499), .B(n17369), .Z(n17368) );
  XOR U16883 ( .A(n17370), .B(n17367), .Z(n17369) );
  XNOR U16884 ( .A(n16990), .B(n17363), .Z(n17365) );
  XOR U16885 ( .A(n17371), .B(n17372), .Z(n16990) );
  AND U16886 ( .A(n497), .B(n17373), .Z(n17372) );
  XOR U16887 ( .A(n17374), .B(n17371), .Z(n17373) );
  XOR U16888 ( .A(n17375), .B(n17376), .Z(n17363) );
  AND U16889 ( .A(n17377), .B(n17378), .Z(n17376) );
  XOR U16890 ( .A(n17375), .B(n17005), .Z(n17378) );
  XOR U16891 ( .A(n17379), .B(n17380), .Z(n17005) );
  AND U16892 ( .A(n499), .B(n17381), .Z(n17380) );
  XOR U16893 ( .A(n17382), .B(n17379), .Z(n17381) );
  XNOR U16894 ( .A(n17002), .B(n17375), .Z(n17377) );
  XOR U16895 ( .A(n17383), .B(n17384), .Z(n17002) );
  AND U16896 ( .A(n497), .B(n17385), .Z(n17384) );
  XOR U16897 ( .A(n17386), .B(n17383), .Z(n17385) );
  XOR U16898 ( .A(n17387), .B(n17388), .Z(n17375) );
  AND U16899 ( .A(n17389), .B(n17390), .Z(n17388) );
  XOR U16900 ( .A(n17387), .B(n17017), .Z(n17390) );
  XOR U16901 ( .A(n17391), .B(n17392), .Z(n17017) );
  AND U16902 ( .A(n499), .B(n17393), .Z(n17392) );
  XOR U16903 ( .A(n17394), .B(n17391), .Z(n17393) );
  XNOR U16904 ( .A(n17014), .B(n17387), .Z(n17389) );
  XOR U16905 ( .A(n17395), .B(n17396), .Z(n17014) );
  AND U16906 ( .A(n497), .B(n17397), .Z(n17396) );
  XOR U16907 ( .A(n17398), .B(n17395), .Z(n17397) );
  XOR U16908 ( .A(n17399), .B(n17400), .Z(n17387) );
  AND U16909 ( .A(n17401), .B(n17402), .Z(n17400) );
  XOR U16910 ( .A(n17399), .B(n17029), .Z(n17402) );
  XOR U16911 ( .A(n17403), .B(n17404), .Z(n17029) );
  AND U16912 ( .A(n499), .B(n17405), .Z(n17404) );
  XOR U16913 ( .A(n17406), .B(n17403), .Z(n17405) );
  XNOR U16914 ( .A(n17026), .B(n17399), .Z(n17401) );
  XOR U16915 ( .A(n17407), .B(n17408), .Z(n17026) );
  AND U16916 ( .A(n497), .B(n17409), .Z(n17408) );
  XOR U16917 ( .A(n17410), .B(n17407), .Z(n17409) );
  XOR U16918 ( .A(n17411), .B(n17412), .Z(n17399) );
  AND U16919 ( .A(n17413), .B(n17414), .Z(n17412) );
  XOR U16920 ( .A(n17411), .B(n17041), .Z(n17414) );
  XOR U16921 ( .A(n17415), .B(n17416), .Z(n17041) );
  AND U16922 ( .A(n499), .B(n17417), .Z(n17416) );
  XOR U16923 ( .A(n17418), .B(n17415), .Z(n17417) );
  XNOR U16924 ( .A(n17038), .B(n17411), .Z(n17413) );
  XOR U16925 ( .A(n17419), .B(n17420), .Z(n17038) );
  AND U16926 ( .A(n497), .B(n17421), .Z(n17420) );
  XOR U16927 ( .A(n17422), .B(n17419), .Z(n17421) );
  XOR U16928 ( .A(n17423), .B(n17424), .Z(n17411) );
  AND U16929 ( .A(n17425), .B(n17426), .Z(n17424) );
  XOR U16930 ( .A(n17423), .B(n17053), .Z(n17426) );
  XOR U16931 ( .A(n17427), .B(n17428), .Z(n17053) );
  AND U16932 ( .A(n499), .B(n17429), .Z(n17428) );
  XOR U16933 ( .A(n17430), .B(n17427), .Z(n17429) );
  XNOR U16934 ( .A(n17050), .B(n17423), .Z(n17425) );
  XOR U16935 ( .A(n17431), .B(n17432), .Z(n17050) );
  AND U16936 ( .A(n497), .B(n17433), .Z(n17432) );
  XOR U16937 ( .A(n17434), .B(n17431), .Z(n17433) );
  XOR U16938 ( .A(n17435), .B(n17436), .Z(n17423) );
  AND U16939 ( .A(n17437), .B(n17438), .Z(n17436) );
  XOR U16940 ( .A(n17435), .B(n17065), .Z(n17438) );
  XOR U16941 ( .A(n17439), .B(n17440), .Z(n17065) );
  AND U16942 ( .A(n499), .B(n17441), .Z(n17440) );
  XOR U16943 ( .A(n17442), .B(n17439), .Z(n17441) );
  XNOR U16944 ( .A(n17062), .B(n17435), .Z(n17437) );
  XOR U16945 ( .A(n17443), .B(n17444), .Z(n17062) );
  AND U16946 ( .A(n497), .B(n17445), .Z(n17444) );
  XOR U16947 ( .A(n17446), .B(n17443), .Z(n17445) );
  XOR U16948 ( .A(n17447), .B(n17448), .Z(n17435) );
  AND U16949 ( .A(n17449), .B(n17450), .Z(n17448) );
  XOR U16950 ( .A(n17447), .B(n17077), .Z(n17450) );
  XOR U16951 ( .A(n17451), .B(n17452), .Z(n17077) );
  AND U16952 ( .A(n499), .B(n17453), .Z(n17452) );
  XOR U16953 ( .A(n17454), .B(n17451), .Z(n17453) );
  XNOR U16954 ( .A(n17074), .B(n17447), .Z(n17449) );
  XOR U16955 ( .A(n17455), .B(n17456), .Z(n17074) );
  AND U16956 ( .A(n497), .B(n17457), .Z(n17456) );
  XOR U16957 ( .A(n17458), .B(n17455), .Z(n17457) );
  XOR U16958 ( .A(n17459), .B(n17460), .Z(n17447) );
  AND U16959 ( .A(n17461), .B(n17462), .Z(n17460) );
  XOR U16960 ( .A(n17459), .B(n17089), .Z(n17462) );
  XOR U16961 ( .A(n17463), .B(n17464), .Z(n17089) );
  AND U16962 ( .A(n499), .B(n17465), .Z(n17464) );
  XOR U16963 ( .A(n17466), .B(n17463), .Z(n17465) );
  XNOR U16964 ( .A(n17086), .B(n17459), .Z(n17461) );
  XOR U16965 ( .A(n17467), .B(n17468), .Z(n17086) );
  AND U16966 ( .A(n497), .B(n17469), .Z(n17468) );
  XOR U16967 ( .A(n17470), .B(n17467), .Z(n17469) );
  XOR U16968 ( .A(n17471), .B(n17472), .Z(n17459) );
  AND U16969 ( .A(n17473), .B(n17474), .Z(n17472) );
  XOR U16970 ( .A(n17471), .B(n17101), .Z(n17474) );
  XOR U16971 ( .A(n17475), .B(n17476), .Z(n17101) );
  AND U16972 ( .A(n499), .B(n17477), .Z(n17476) );
  XOR U16973 ( .A(n17478), .B(n17475), .Z(n17477) );
  XNOR U16974 ( .A(n17098), .B(n17471), .Z(n17473) );
  XOR U16975 ( .A(n17479), .B(n17480), .Z(n17098) );
  AND U16976 ( .A(n497), .B(n17481), .Z(n17480) );
  XOR U16977 ( .A(n17482), .B(n17479), .Z(n17481) );
  XOR U16978 ( .A(n17483), .B(n17484), .Z(n17471) );
  AND U16979 ( .A(n17485), .B(n17486), .Z(n17484) );
  XOR U16980 ( .A(n17483), .B(n17113), .Z(n17486) );
  XOR U16981 ( .A(n17487), .B(n17488), .Z(n17113) );
  AND U16982 ( .A(n499), .B(n17489), .Z(n17488) );
  XOR U16983 ( .A(n17490), .B(n17487), .Z(n17489) );
  XNOR U16984 ( .A(n17110), .B(n17483), .Z(n17485) );
  XOR U16985 ( .A(n17491), .B(n17492), .Z(n17110) );
  AND U16986 ( .A(n497), .B(n17493), .Z(n17492) );
  XOR U16987 ( .A(n17494), .B(n17491), .Z(n17493) );
  XOR U16988 ( .A(n17495), .B(n17496), .Z(n17483) );
  AND U16989 ( .A(n17497), .B(n17498), .Z(n17496) );
  XOR U16990 ( .A(n17495), .B(n17125), .Z(n17498) );
  XOR U16991 ( .A(n17499), .B(n17500), .Z(n17125) );
  AND U16992 ( .A(n499), .B(n17501), .Z(n17500) );
  XOR U16993 ( .A(n17502), .B(n17499), .Z(n17501) );
  XNOR U16994 ( .A(n17122), .B(n17495), .Z(n17497) );
  XOR U16995 ( .A(n17503), .B(n17504), .Z(n17122) );
  AND U16996 ( .A(n497), .B(n17505), .Z(n17504) );
  XOR U16997 ( .A(n17506), .B(n17503), .Z(n17505) );
  XOR U16998 ( .A(n17507), .B(n17508), .Z(n17495) );
  AND U16999 ( .A(n17509), .B(n17510), .Z(n17508) );
  XOR U17000 ( .A(n17507), .B(n17137), .Z(n17510) );
  XOR U17001 ( .A(n17511), .B(n17512), .Z(n17137) );
  AND U17002 ( .A(n499), .B(n17513), .Z(n17512) );
  XOR U17003 ( .A(n17514), .B(n17511), .Z(n17513) );
  XNOR U17004 ( .A(n17134), .B(n17507), .Z(n17509) );
  XOR U17005 ( .A(n17515), .B(n17516), .Z(n17134) );
  AND U17006 ( .A(n497), .B(n17517), .Z(n17516) );
  XOR U17007 ( .A(n17518), .B(n17515), .Z(n17517) );
  XOR U17008 ( .A(n17519), .B(n17520), .Z(n17507) );
  AND U17009 ( .A(n17521), .B(n17522), .Z(n17520) );
  XOR U17010 ( .A(n17519), .B(n17149), .Z(n17522) );
  XOR U17011 ( .A(n17523), .B(n17524), .Z(n17149) );
  AND U17012 ( .A(n499), .B(n17525), .Z(n17524) );
  XOR U17013 ( .A(n17526), .B(n17523), .Z(n17525) );
  XNOR U17014 ( .A(n17146), .B(n17519), .Z(n17521) );
  XOR U17015 ( .A(n17527), .B(n17528), .Z(n17146) );
  AND U17016 ( .A(n497), .B(n17529), .Z(n17528) );
  XOR U17017 ( .A(n17530), .B(n17527), .Z(n17529) );
  XOR U17018 ( .A(n17531), .B(n17532), .Z(n17519) );
  AND U17019 ( .A(n17533), .B(n17534), .Z(n17532) );
  XOR U17020 ( .A(n17531), .B(n17161), .Z(n17534) );
  XOR U17021 ( .A(n17535), .B(n17536), .Z(n17161) );
  AND U17022 ( .A(n499), .B(n17537), .Z(n17536) );
  XOR U17023 ( .A(n17538), .B(n17535), .Z(n17537) );
  XNOR U17024 ( .A(n17158), .B(n17531), .Z(n17533) );
  XOR U17025 ( .A(n17539), .B(n17540), .Z(n17158) );
  AND U17026 ( .A(n497), .B(n17541), .Z(n17540) );
  XOR U17027 ( .A(n17542), .B(n17539), .Z(n17541) );
  XOR U17028 ( .A(n17543), .B(n17544), .Z(n17531) );
  AND U17029 ( .A(n17545), .B(n17546), .Z(n17544) );
  XOR U17030 ( .A(n17543), .B(n17173), .Z(n17546) );
  XOR U17031 ( .A(n17547), .B(n17548), .Z(n17173) );
  AND U17032 ( .A(n499), .B(n17549), .Z(n17548) );
  XOR U17033 ( .A(n17550), .B(n17547), .Z(n17549) );
  XNOR U17034 ( .A(n17170), .B(n17543), .Z(n17545) );
  XOR U17035 ( .A(n17551), .B(n17552), .Z(n17170) );
  AND U17036 ( .A(n497), .B(n17553), .Z(n17552) );
  XOR U17037 ( .A(n17554), .B(n17551), .Z(n17553) );
  XOR U17038 ( .A(n17555), .B(n17556), .Z(n17543) );
  AND U17039 ( .A(n17557), .B(n17558), .Z(n17556) );
  XOR U17040 ( .A(n17555), .B(n17185), .Z(n17558) );
  XOR U17041 ( .A(n17559), .B(n17560), .Z(n17185) );
  AND U17042 ( .A(n499), .B(n17561), .Z(n17560) );
  XOR U17043 ( .A(n17562), .B(n17559), .Z(n17561) );
  XNOR U17044 ( .A(n17182), .B(n17555), .Z(n17557) );
  XOR U17045 ( .A(n17563), .B(n17564), .Z(n17182) );
  AND U17046 ( .A(n497), .B(n17565), .Z(n17564) );
  XOR U17047 ( .A(n17566), .B(n17563), .Z(n17565) );
  XOR U17048 ( .A(n17567), .B(n17568), .Z(n17555) );
  AND U17049 ( .A(n17569), .B(n17570), .Z(n17568) );
  XOR U17050 ( .A(n17567), .B(n17197), .Z(n17570) );
  XOR U17051 ( .A(n17571), .B(n17572), .Z(n17197) );
  AND U17052 ( .A(n499), .B(n17573), .Z(n17572) );
  XOR U17053 ( .A(n17574), .B(n17571), .Z(n17573) );
  XNOR U17054 ( .A(n17194), .B(n17567), .Z(n17569) );
  XOR U17055 ( .A(n17575), .B(n17576), .Z(n17194) );
  AND U17056 ( .A(n497), .B(n17577), .Z(n17576) );
  XOR U17057 ( .A(n17578), .B(n17575), .Z(n17577) );
  XOR U17058 ( .A(n17579), .B(n17580), .Z(n17567) );
  AND U17059 ( .A(n17581), .B(n17582), .Z(n17580) );
  XOR U17060 ( .A(n17579), .B(n17209), .Z(n17582) );
  XOR U17061 ( .A(n17583), .B(n17584), .Z(n17209) );
  AND U17062 ( .A(n499), .B(n17585), .Z(n17584) );
  XOR U17063 ( .A(n17586), .B(n17583), .Z(n17585) );
  XNOR U17064 ( .A(n17206), .B(n17579), .Z(n17581) );
  XOR U17065 ( .A(n17587), .B(n17588), .Z(n17206) );
  AND U17066 ( .A(n497), .B(n17589), .Z(n17588) );
  XOR U17067 ( .A(n17590), .B(n17587), .Z(n17589) );
  XOR U17068 ( .A(n17591), .B(n17592), .Z(n17579) );
  AND U17069 ( .A(n17593), .B(n17594), .Z(n17592) );
  XNOR U17070 ( .A(n17595), .B(n17222), .Z(n17594) );
  XOR U17071 ( .A(n17596), .B(n17597), .Z(n17222) );
  AND U17072 ( .A(n499), .B(n17598), .Z(n17597) );
  XOR U17073 ( .A(n17596), .B(n17599), .Z(n17598) );
  XNOR U17074 ( .A(n17219), .B(n17591), .Z(n17593) );
  XOR U17075 ( .A(n17600), .B(n17601), .Z(n17219) );
  AND U17076 ( .A(n497), .B(n17602), .Z(n17601) );
  XOR U17077 ( .A(n17600), .B(n17603), .Z(n17602) );
  IV U17078 ( .A(n17595), .Z(n17591) );
  AND U17079 ( .A(n17227), .B(n17230), .Z(n17595) );
  XNOR U17080 ( .A(n17604), .B(n17605), .Z(n17230) );
  AND U17081 ( .A(n499), .B(n17606), .Z(n17605) );
  XNOR U17082 ( .A(n17607), .B(n17604), .Z(n17606) );
  XOR U17083 ( .A(n17608), .B(n17609), .Z(n499) );
  AND U17084 ( .A(n17610), .B(n17611), .Z(n17609) );
  XOR U17085 ( .A(n17238), .B(n17608), .Z(n17611) );
  IV U17086 ( .A(n17612), .Z(n17238) );
  AND U17087 ( .A(p_input[6143]), .B(p_input[6111]), .Z(n17612) );
  XOR U17088 ( .A(n17608), .B(n17235), .Z(n17610) );
  AND U17089 ( .A(p_input[6047]), .B(p_input[6079]), .Z(n17235) );
  XOR U17090 ( .A(n17613), .B(n17614), .Z(n17608) );
  AND U17091 ( .A(n17615), .B(n17616), .Z(n17614) );
  XOR U17092 ( .A(n17613), .B(n17250), .Z(n17616) );
  XNOR U17093 ( .A(p_input[6110]), .B(n17617), .Z(n17250) );
  AND U17094 ( .A(n311), .B(n17618), .Z(n17617) );
  XOR U17095 ( .A(p_input[6142]), .B(p_input[6110]), .Z(n17618) );
  XNOR U17096 ( .A(n17247), .B(n17613), .Z(n17615) );
  XOR U17097 ( .A(n17619), .B(n17620), .Z(n17247) );
  AND U17098 ( .A(n309), .B(n17621), .Z(n17620) );
  XOR U17099 ( .A(p_input[6078]), .B(p_input[6046]), .Z(n17621) );
  XOR U17100 ( .A(n17622), .B(n17623), .Z(n17613) );
  AND U17101 ( .A(n17624), .B(n17625), .Z(n17623) );
  XOR U17102 ( .A(n17622), .B(n17262), .Z(n17625) );
  XNOR U17103 ( .A(p_input[6109]), .B(n17626), .Z(n17262) );
  AND U17104 ( .A(n311), .B(n17627), .Z(n17626) );
  XOR U17105 ( .A(p_input[6141]), .B(p_input[6109]), .Z(n17627) );
  XNOR U17106 ( .A(n17259), .B(n17622), .Z(n17624) );
  XOR U17107 ( .A(n17628), .B(n17629), .Z(n17259) );
  AND U17108 ( .A(n309), .B(n17630), .Z(n17629) );
  XOR U17109 ( .A(p_input[6077]), .B(p_input[6045]), .Z(n17630) );
  XOR U17110 ( .A(n17631), .B(n17632), .Z(n17622) );
  AND U17111 ( .A(n17633), .B(n17634), .Z(n17632) );
  XOR U17112 ( .A(n17631), .B(n17274), .Z(n17634) );
  XNOR U17113 ( .A(p_input[6108]), .B(n17635), .Z(n17274) );
  AND U17114 ( .A(n311), .B(n17636), .Z(n17635) );
  XOR U17115 ( .A(p_input[6140]), .B(p_input[6108]), .Z(n17636) );
  XNOR U17116 ( .A(n17271), .B(n17631), .Z(n17633) );
  XOR U17117 ( .A(n17637), .B(n17638), .Z(n17271) );
  AND U17118 ( .A(n309), .B(n17639), .Z(n17638) );
  XOR U17119 ( .A(p_input[6076]), .B(p_input[6044]), .Z(n17639) );
  XOR U17120 ( .A(n17640), .B(n17641), .Z(n17631) );
  AND U17121 ( .A(n17642), .B(n17643), .Z(n17641) );
  XOR U17122 ( .A(n17640), .B(n17286), .Z(n17643) );
  XNOR U17123 ( .A(p_input[6107]), .B(n17644), .Z(n17286) );
  AND U17124 ( .A(n311), .B(n17645), .Z(n17644) );
  XOR U17125 ( .A(p_input[6139]), .B(p_input[6107]), .Z(n17645) );
  XNOR U17126 ( .A(n17283), .B(n17640), .Z(n17642) );
  XOR U17127 ( .A(n17646), .B(n17647), .Z(n17283) );
  AND U17128 ( .A(n309), .B(n17648), .Z(n17647) );
  XOR U17129 ( .A(p_input[6075]), .B(p_input[6043]), .Z(n17648) );
  XOR U17130 ( .A(n17649), .B(n17650), .Z(n17640) );
  AND U17131 ( .A(n17651), .B(n17652), .Z(n17650) );
  XOR U17132 ( .A(n17649), .B(n17298), .Z(n17652) );
  XNOR U17133 ( .A(p_input[6106]), .B(n17653), .Z(n17298) );
  AND U17134 ( .A(n311), .B(n17654), .Z(n17653) );
  XOR U17135 ( .A(p_input[6138]), .B(p_input[6106]), .Z(n17654) );
  XNOR U17136 ( .A(n17295), .B(n17649), .Z(n17651) );
  XOR U17137 ( .A(n17655), .B(n17656), .Z(n17295) );
  AND U17138 ( .A(n309), .B(n17657), .Z(n17656) );
  XOR U17139 ( .A(p_input[6074]), .B(p_input[6042]), .Z(n17657) );
  XOR U17140 ( .A(n17658), .B(n17659), .Z(n17649) );
  AND U17141 ( .A(n17660), .B(n17661), .Z(n17659) );
  XOR U17142 ( .A(n17658), .B(n17310), .Z(n17661) );
  XNOR U17143 ( .A(p_input[6105]), .B(n17662), .Z(n17310) );
  AND U17144 ( .A(n311), .B(n17663), .Z(n17662) );
  XOR U17145 ( .A(p_input[6137]), .B(p_input[6105]), .Z(n17663) );
  XNOR U17146 ( .A(n17307), .B(n17658), .Z(n17660) );
  XOR U17147 ( .A(n17664), .B(n17665), .Z(n17307) );
  AND U17148 ( .A(n309), .B(n17666), .Z(n17665) );
  XOR U17149 ( .A(p_input[6073]), .B(p_input[6041]), .Z(n17666) );
  XOR U17150 ( .A(n17667), .B(n17668), .Z(n17658) );
  AND U17151 ( .A(n17669), .B(n17670), .Z(n17668) );
  XOR U17152 ( .A(n17667), .B(n17322), .Z(n17670) );
  XNOR U17153 ( .A(p_input[6104]), .B(n17671), .Z(n17322) );
  AND U17154 ( .A(n311), .B(n17672), .Z(n17671) );
  XOR U17155 ( .A(p_input[6136]), .B(p_input[6104]), .Z(n17672) );
  XNOR U17156 ( .A(n17319), .B(n17667), .Z(n17669) );
  XOR U17157 ( .A(n17673), .B(n17674), .Z(n17319) );
  AND U17158 ( .A(n309), .B(n17675), .Z(n17674) );
  XOR U17159 ( .A(p_input[6072]), .B(p_input[6040]), .Z(n17675) );
  XOR U17160 ( .A(n17676), .B(n17677), .Z(n17667) );
  AND U17161 ( .A(n17678), .B(n17679), .Z(n17677) );
  XOR U17162 ( .A(n17676), .B(n17334), .Z(n17679) );
  XNOR U17163 ( .A(p_input[6103]), .B(n17680), .Z(n17334) );
  AND U17164 ( .A(n311), .B(n17681), .Z(n17680) );
  XOR U17165 ( .A(p_input[6135]), .B(p_input[6103]), .Z(n17681) );
  XNOR U17166 ( .A(n17331), .B(n17676), .Z(n17678) );
  XOR U17167 ( .A(n17682), .B(n17683), .Z(n17331) );
  AND U17168 ( .A(n309), .B(n17684), .Z(n17683) );
  XOR U17169 ( .A(p_input[6071]), .B(p_input[6039]), .Z(n17684) );
  XOR U17170 ( .A(n17685), .B(n17686), .Z(n17676) );
  AND U17171 ( .A(n17687), .B(n17688), .Z(n17686) );
  XOR U17172 ( .A(n17685), .B(n17346), .Z(n17688) );
  XNOR U17173 ( .A(p_input[6102]), .B(n17689), .Z(n17346) );
  AND U17174 ( .A(n311), .B(n17690), .Z(n17689) );
  XOR U17175 ( .A(p_input[6134]), .B(p_input[6102]), .Z(n17690) );
  XNOR U17176 ( .A(n17343), .B(n17685), .Z(n17687) );
  XOR U17177 ( .A(n17691), .B(n17692), .Z(n17343) );
  AND U17178 ( .A(n309), .B(n17693), .Z(n17692) );
  XOR U17179 ( .A(p_input[6070]), .B(p_input[6038]), .Z(n17693) );
  XOR U17180 ( .A(n17694), .B(n17695), .Z(n17685) );
  AND U17181 ( .A(n17696), .B(n17697), .Z(n17695) );
  XOR U17182 ( .A(n17694), .B(n17358), .Z(n17697) );
  XNOR U17183 ( .A(p_input[6101]), .B(n17698), .Z(n17358) );
  AND U17184 ( .A(n311), .B(n17699), .Z(n17698) );
  XOR U17185 ( .A(p_input[6133]), .B(p_input[6101]), .Z(n17699) );
  XNOR U17186 ( .A(n17355), .B(n17694), .Z(n17696) );
  XOR U17187 ( .A(n17700), .B(n17701), .Z(n17355) );
  AND U17188 ( .A(n309), .B(n17702), .Z(n17701) );
  XOR U17189 ( .A(p_input[6069]), .B(p_input[6037]), .Z(n17702) );
  XOR U17190 ( .A(n17703), .B(n17704), .Z(n17694) );
  AND U17191 ( .A(n17705), .B(n17706), .Z(n17704) );
  XOR U17192 ( .A(n17703), .B(n17370), .Z(n17706) );
  XNOR U17193 ( .A(p_input[6100]), .B(n17707), .Z(n17370) );
  AND U17194 ( .A(n311), .B(n17708), .Z(n17707) );
  XOR U17195 ( .A(p_input[6132]), .B(p_input[6100]), .Z(n17708) );
  XNOR U17196 ( .A(n17367), .B(n17703), .Z(n17705) );
  XOR U17197 ( .A(n17709), .B(n17710), .Z(n17367) );
  AND U17198 ( .A(n309), .B(n17711), .Z(n17710) );
  XOR U17199 ( .A(p_input[6068]), .B(p_input[6036]), .Z(n17711) );
  XOR U17200 ( .A(n17712), .B(n17713), .Z(n17703) );
  AND U17201 ( .A(n17714), .B(n17715), .Z(n17713) );
  XOR U17202 ( .A(n17712), .B(n17382), .Z(n17715) );
  XNOR U17203 ( .A(p_input[6099]), .B(n17716), .Z(n17382) );
  AND U17204 ( .A(n311), .B(n17717), .Z(n17716) );
  XOR U17205 ( .A(p_input[6131]), .B(p_input[6099]), .Z(n17717) );
  XNOR U17206 ( .A(n17379), .B(n17712), .Z(n17714) );
  XOR U17207 ( .A(n17718), .B(n17719), .Z(n17379) );
  AND U17208 ( .A(n309), .B(n17720), .Z(n17719) );
  XOR U17209 ( .A(p_input[6067]), .B(p_input[6035]), .Z(n17720) );
  XOR U17210 ( .A(n17721), .B(n17722), .Z(n17712) );
  AND U17211 ( .A(n17723), .B(n17724), .Z(n17722) );
  XOR U17212 ( .A(n17721), .B(n17394), .Z(n17724) );
  XNOR U17213 ( .A(p_input[6098]), .B(n17725), .Z(n17394) );
  AND U17214 ( .A(n311), .B(n17726), .Z(n17725) );
  XOR U17215 ( .A(p_input[6130]), .B(p_input[6098]), .Z(n17726) );
  XNOR U17216 ( .A(n17391), .B(n17721), .Z(n17723) );
  XOR U17217 ( .A(n17727), .B(n17728), .Z(n17391) );
  AND U17218 ( .A(n309), .B(n17729), .Z(n17728) );
  XOR U17219 ( .A(p_input[6066]), .B(p_input[6034]), .Z(n17729) );
  XOR U17220 ( .A(n17730), .B(n17731), .Z(n17721) );
  AND U17221 ( .A(n17732), .B(n17733), .Z(n17731) );
  XOR U17222 ( .A(n17730), .B(n17406), .Z(n17733) );
  XNOR U17223 ( .A(p_input[6097]), .B(n17734), .Z(n17406) );
  AND U17224 ( .A(n311), .B(n17735), .Z(n17734) );
  XOR U17225 ( .A(p_input[6129]), .B(p_input[6097]), .Z(n17735) );
  XNOR U17226 ( .A(n17403), .B(n17730), .Z(n17732) );
  XOR U17227 ( .A(n17736), .B(n17737), .Z(n17403) );
  AND U17228 ( .A(n309), .B(n17738), .Z(n17737) );
  XOR U17229 ( .A(p_input[6065]), .B(p_input[6033]), .Z(n17738) );
  XOR U17230 ( .A(n17739), .B(n17740), .Z(n17730) );
  AND U17231 ( .A(n17741), .B(n17742), .Z(n17740) );
  XOR U17232 ( .A(n17739), .B(n17418), .Z(n17742) );
  XNOR U17233 ( .A(p_input[6096]), .B(n17743), .Z(n17418) );
  AND U17234 ( .A(n311), .B(n17744), .Z(n17743) );
  XOR U17235 ( .A(p_input[6128]), .B(p_input[6096]), .Z(n17744) );
  XNOR U17236 ( .A(n17415), .B(n17739), .Z(n17741) );
  XOR U17237 ( .A(n17745), .B(n17746), .Z(n17415) );
  AND U17238 ( .A(n309), .B(n17747), .Z(n17746) );
  XOR U17239 ( .A(p_input[6064]), .B(p_input[6032]), .Z(n17747) );
  XOR U17240 ( .A(n17748), .B(n17749), .Z(n17739) );
  AND U17241 ( .A(n17750), .B(n17751), .Z(n17749) );
  XOR U17242 ( .A(n17748), .B(n17430), .Z(n17751) );
  XNOR U17243 ( .A(p_input[6095]), .B(n17752), .Z(n17430) );
  AND U17244 ( .A(n311), .B(n17753), .Z(n17752) );
  XOR U17245 ( .A(p_input[6127]), .B(p_input[6095]), .Z(n17753) );
  XNOR U17246 ( .A(n17427), .B(n17748), .Z(n17750) );
  XOR U17247 ( .A(n17754), .B(n17755), .Z(n17427) );
  AND U17248 ( .A(n309), .B(n17756), .Z(n17755) );
  XOR U17249 ( .A(p_input[6063]), .B(p_input[6031]), .Z(n17756) );
  XOR U17250 ( .A(n17757), .B(n17758), .Z(n17748) );
  AND U17251 ( .A(n17759), .B(n17760), .Z(n17758) );
  XOR U17252 ( .A(n17757), .B(n17442), .Z(n17760) );
  XNOR U17253 ( .A(p_input[6094]), .B(n17761), .Z(n17442) );
  AND U17254 ( .A(n311), .B(n17762), .Z(n17761) );
  XOR U17255 ( .A(p_input[6126]), .B(p_input[6094]), .Z(n17762) );
  XNOR U17256 ( .A(n17439), .B(n17757), .Z(n17759) );
  XOR U17257 ( .A(n17763), .B(n17764), .Z(n17439) );
  AND U17258 ( .A(n309), .B(n17765), .Z(n17764) );
  XOR U17259 ( .A(p_input[6062]), .B(p_input[6030]), .Z(n17765) );
  XOR U17260 ( .A(n17766), .B(n17767), .Z(n17757) );
  AND U17261 ( .A(n17768), .B(n17769), .Z(n17767) );
  XOR U17262 ( .A(n17766), .B(n17454), .Z(n17769) );
  XNOR U17263 ( .A(p_input[6093]), .B(n17770), .Z(n17454) );
  AND U17264 ( .A(n311), .B(n17771), .Z(n17770) );
  XOR U17265 ( .A(p_input[6125]), .B(p_input[6093]), .Z(n17771) );
  XNOR U17266 ( .A(n17451), .B(n17766), .Z(n17768) );
  XOR U17267 ( .A(n17772), .B(n17773), .Z(n17451) );
  AND U17268 ( .A(n309), .B(n17774), .Z(n17773) );
  XOR U17269 ( .A(p_input[6061]), .B(p_input[6029]), .Z(n17774) );
  XOR U17270 ( .A(n17775), .B(n17776), .Z(n17766) );
  AND U17271 ( .A(n17777), .B(n17778), .Z(n17776) );
  XOR U17272 ( .A(n17775), .B(n17466), .Z(n17778) );
  XNOR U17273 ( .A(p_input[6092]), .B(n17779), .Z(n17466) );
  AND U17274 ( .A(n311), .B(n17780), .Z(n17779) );
  XOR U17275 ( .A(p_input[6124]), .B(p_input[6092]), .Z(n17780) );
  XNOR U17276 ( .A(n17463), .B(n17775), .Z(n17777) );
  XOR U17277 ( .A(n17781), .B(n17782), .Z(n17463) );
  AND U17278 ( .A(n309), .B(n17783), .Z(n17782) );
  XOR U17279 ( .A(p_input[6060]), .B(p_input[6028]), .Z(n17783) );
  XOR U17280 ( .A(n17784), .B(n17785), .Z(n17775) );
  AND U17281 ( .A(n17786), .B(n17787), .Z(n17785) );
  XOR U17282 ( .A(n17784), .B(n17478), .Z(n17787) );
  XNOR U17283 ( .A(p_input[6091]), .B(n17788), .Z(n17478) );
  AND U17284 ( .A(n311), .B(n17789), .Z(n17788) );
  XOR U17285 ( .A(p_input[6123]), .B(p_input[6091]), .Z(n17789) );
  XNOR U17286 ( .A(n17475), .B(n17784), .Z(n17786) );
  XOR U17287 ( .A(n17790), .B(n17791), .Z(n17475) );
  AND U17288 ( .A(n309), .B(n17792), .Z(n17791) );
  XOR U17289 ( .A(p_input[6059]), .B(p_input[6027]), .Z(n17792) );
  XOR U17290 ( .A(n17793), .B(n17794), .Z(n17784) );
  AND U17291 ( .A(n17795), .B(n17796), .Z(n17794) );
  XOR U17292 ( .A(n17793), .B(n17490), .Z(n17796) );
  XNOR U17293 ( .A(p_input[6090]), .B(n17797), .Z(n17490) );
  AND U17294 ( .A(n311), .B(n17798), .Z(n17797) );
  XOR U17295 ( .A(p_input[6122]), .B(p_input[6090]), .Z(n17798) );
  XNOR U17296 ( .A(n17487), .B(n17793), .Z(n17795) );
  XOR U17297 ( .A(n17799), .B(n17800), .Z(n17487) );
  AND U17298 ( .A(n309), .B(n17801), .Z(n17800) );
  XOR U17299 ( .A(p_input[6058]), .B(p_input[6026]), .Z(n17801) );
  XOR U17300 ( .A(n17802), .B(n17803), .Z(n17793) );
  AND U17301 ( .A(n17804), .B(n17805), .Z(n17803) );
  XOR U17302 ( .A(n17802), .B(n17502), .Z(n17805) );
  XNOR U17303 ( .A(p_input[6089]), .B(n17806), .Z(n17502) );
  AND U17304 ( .A(n311), .B(n17807), .Z(n17806) );
  XOR U17305 ( .A(p_input[6121]), .B(p_input[6089]), .Z(n17807) );
  XNOR U17306 ( .A(n17499), .B(n17802), .Z(n17804) );
  XOR U17307 ( .A(n17808), .B(n17809), .Z(n17499) );
  AND U17308 ( .A(n309), .B(n17810), .Z(n17809) );
  XOR U17309 ( .A(p_input[6057]), .B(p_input[6025]), .Z(n17810) );
  XOR U17310 ( .A(n17811), .B(n17812), .Z(n17802) );
  AND U17311 ( .A(n17813), .B(n17814), .Z(n17812) );
  XOR U17312 ( .A(n17811), .B(n17514), .Z(n17814) );
  XNOR U17313 ( .A(p_input[6088]), .B(n17815), .Z(n17514) );
  AND U17314 ( .A(n311), .B(n17816), .Z(n17815) );
  XOR U17315 ( .A(p_input[6120]), .B(p_input[6088]), .Z(n17816) );
  XNOR U17316 ( .A(n17511), .B(n17811), .Z(n17813) );
  XOR U17317 ( .A(n17817), .B(n17818), .Z(n17511) );
  AND U17318 ( .A(n309), .B(n17819), .Z(n17818) );
  XOR U17319 ( .A(p_input[6056]), .B(p_input[6024]), .Z(n17819) );
  XOR U17320 ( .A(n17820), .B(n17821), .Z(n17811) );
  AND U17321 ( .A(n17822), .B(n17823), .Z(n17821) );
  XOR U17322 ( .A(n17820), .B(n17526), .Z(n17823) );
  XNOR U17323 ( .A(p_input[6087]), .B(n17824), .Z(n17526) );
  AND U17324 ( .A(n311), .B(n17825), .Z(n17824) );
  XOR U17325 ( .A(p_input[6119]), .B(p_input[6087]), .Z(n17825) );
  XNOR U17326 ( .A(n17523), .B(n17820), .Z(n17822) );
  XOR U17327 ( .A(n17826), .B(n17827), .Z(n17523) );
  AND U17328 ( .A(n309), .B(n17828), .Z(n17827) );
  XOR U17329 ( .A(p_input[6055]), .B(p_input[6023]), .Z(n17828) );
  XOR U17330 ( .A(n17829), .B(n17830), .Z(n17820) );
  AND U17331 ( .A(n17831), .B(n17832), .Z(n17830) );
  XOR U17332 ( .A(n17829), .B(n17538), .Z(n17832) );
  XNOR U17333 ( .A(p_input[6086]), .B(n17833), .Z(n17538) );
  AND U17334 ( .A(n311), .B(n17834), .Z(n17833) );
  XOR U17335 ( .A(p_input[6118]), .B(p_input[6086]), .Z(n17834) );
  XNOR U17336 ( .A(n17535), .B(n17829), .Z(n17831) );
  XOR U17337 ( .A(n17835), .B(n17836), .Z(n17535) );
  AND U17338 ( .A(n309), .B(n17837), .Z(n17836) );
  XOR U17339 ( .A(p_input[6054]), .B(p_input[6022]), .Z(n17837) );
  XOR U17340 ( .A(n17838), .B(n17839), .Z(n17829) );
  AND U17341 ( .A(n17840), .B(n17841), .Z(n17839) );
  XOR U17342 ( .A(n17838), .B(n17550), .Z(n17841) );
  XNOR U17343 ( .A(p_input[6085]), .B(n17842), .Z(n17550) );
  AND U17344 ( .A(n311), .B(n17843), .Z(n17842) );
  XOR U17345 ( .A(p_input[6117]), .B(p_input[6085]), .Z(n17843) );
  XNOR U17346 ( .A(n17547), .B(n17838), .Z(n17840) );
  XOR U17347 ( .A(n17844), .B(n17845), .Z(n17547) );
  AND U17348 ( .A(n309), .B(n17846), .Z(n17845) );
  XOR U17349 ( .A(p_input[6053]), .B(p_input[6021]), .Z(n17846) );
  XOR U17350 ( .A(n17847), .B(n17848), .Z(n17838) );
  AND U17351 ( .A(n17849), .B(n17850), .Z(n17848) );
  XOR U17352 ( .A(n17847), .B(n17562), .Z(n17850) );
  XNOR U17353 ( .A(p_input[6084]), .B(n17851), .Z(n17562) );
  AND U17354 ( .A(n311), .B(n17852), .Z(n17851) );
  XOR U17355 ( .A(p_input[6116]), .B(p_input[6084]), .Z(n17852) );
  XNOR U17356 ( .A(n17559), .B(n17847), .Z(n17849) );
  XOR U17357 ( .A(n17853), .B(n17854), .Z(n17559) );
  AND U17358 ( .A(n309), .B(n17855), .Z(n17854) );
  XOR U17359 ( .A(p_input[6052]), .B(p_input[6020]), .Z(n17855) );
  XOR U17360 ( .A(n17856), .B(n17857), .Z(n17847) );
  AND U17361 ( .A(n17858), .B(n17859), .Z(n17857) );
  XOR U17362 ( .A(n17856), .B(n17574), .Z(n17859) );
  XNOR U17363 ( .A(p_input[6083]), .B(n17860), .Z(n17574) );
  AND U17364 ( .A(n311), .B(n17861), .Z(n17860) );
  XOR U17365 ( .A(p_input[6115]), .B(p_input[6083]), .Z(n17861) );
  XNOR U17366 ( .A(n17571), .B(n17856), .Z(n17858) );
  XOR U17367 ( .A(n17862), .B(n17863), .Z(n17571) );
  AND U17368 ( .A(n309), .B(n17864), .Z(n17863) );
  XOR U17369 ( .A(p_input[6051]), .B(p_input[6019]), .Z(n17864) );
  XOR U17370 ( .A(n17865), .B(n17866), .Z(n17856) );
  AND U17371 ( .A(n17867), .B(n17868), .Z(n17866) );
  XOR U17372 ( .A(n17865), .B(n17586), .Z(n17868) );
  XNOR U17373 ( .A(p_input[6082]), .B(n17869), .Z(n17586) );
  AND U17374 ( .A(n311), .B(n17870), .Z(n17869) );
  XOR U17375 ( .A(p_input[6114]), .B(p_input[6082]), .Z(n17870) );
  XNOR U17376 ( .A(n17583), .B(n17865), .Z(n17867) );
  XOR U17377 ( .A(n17871), .B(n17872), .Z(n17583) );
  AND U17378 ( .A(n309), .B(n17873), .Z(n17872) );
  XOR U17379 ( .A(p_input[6050]), .B(p_input[6018]), .Z(n17873) );
  XOR U17380 ( .A(n17874), .B(n17875), .Z(n17865) );
  AND U17381 ( .A(n17876), .B(n17877), .Z(n17875) );
  XNOR U17382 ( .A(n17878), .B(n17599), .Z(n17877) );
  XNOR U17383 ( .A(p_input[6081]), .B(n17879), .Z(n17599) );
  AND U17384 ( .A(n311), .B(n17880), .Z(n17879) );
  XNOR U17385 ( .A(p_input[6113]), .B(n17881), .Z(n17880) );
  IV U17386 ( .A(p_input[6081]), .Z(n17881) );
  XNOR U17387 ( .A(n17596), .B(n17874), .Z(n17876) );
  XNOR U17388 ( .A(p_input[6017]), .B(n17882), .Z(n17596) );
  AND U17389 ( .A(n309), .B(n17883), .Z(n17882) );
  XOR U17390 ( .A(p_input[6049]), .B(p_input[6017]), .Z(n17883) );
  IV U17391 ( .A(n17878), .Z(n17874) );
  AND U17392 ( .A(n17604), .B(n17607), .Z(n17878) );
  XOR U17393 ( .A(p_input[6080]), .B(n17884), .Z(n17607) );
  AND U17394 ( .A(n311), .B(n17885), .Z(n17884) );
  XOR U17395 ( .A(p_input[6112]), .B(p_input[6080]), .Z(n17885) );
  XOR U17396 ( .A(n17886), .B(n17887), .Z(n311) );
  AND U17397 ( .A(n17888), .B(n17889), .Z(n17887) );
  XNOR U17398 ( .A(p_input[6143]), .B(n17886), .Z(n17889) );
  XOR U17399 ( .A(n17886), .B(p_input[6111]), .Z(n17888) );
  XOR U17400 ( .A(n17890), .B(n17891), .Z(n17886) );
  AND U17401 ( .A(n17892), .B(n17893), .Z(n17891) );
  XNOR U17402 ( .A(p_input[6142]), .B(n17890), .Z(n17893) );
  XOR U17403 ( .A(n17890), .B(p_input[6110]), .Z(n17892) );
  XOR U17404 ( .A(n17894), .B(n17895), .Z(n17890) );
  AND U17405 ( .A(n17896), .B(n17897), .Z(n17895) );
  XNOR U17406 ( .A(p_input[6141]), .B(n17894), .Z(n17897) );
  XOR U17407 ( .A(n17894), .B(p_input[6109]), .Z(n17896) );
  XOR U17408 ( .A(n17898), .B(n17899), .Z(n17894) );
  AND U17409 ( .A(n17900), .B(n17901), .Z(n17899) );
  XNOR U17410 ( .A(p_input[6140]), .B(n17898), .Z(n17901) );
  XOR U17411 ( .A(n17898), .B(p_input[6108]), .Z(n17900) );
  XOR U17412 ( .A(n17902), .B(n17903), .Z(n17898) );
  AND U17413 ( .A(n17904), .B(n17905), .Z(n17903) );
  XNOR U17414 ( .A(p_input[6139]), .B(n17902), .Z(n17905) );
  XOR U17415 ( .A(n17902), .B(p_input[6107]), .Z(n17904) );
  XOR U17416 ( .A(n17906), .B(n17907), .Z(n17902) );
  AND U17417 ( .A(n17908), .B(n17909), .Z(n17907) );
  XNOR U17418 ( .A(p_input[6138]), .B(n17906), .Z(n17909) );
  XOR U17419 ( .A(n17906), .B(p_input[6106]), .Z(n17908) );
  XOR U17420 ( .A(n17910), .B(n17911), .Z(n17906) );
  AND U17421 ( .A(n17912), .B(n17913), .Z(n17911) );
  XNOR U17422 ( .A(p_input[6137]), .B(n17910), .Z(n17913) );
  XOR U17423 ( .A(n17910), .B(p_input[6105]), .Z(n17912) );
  XOR U17424 ( .A(n17914), .B(n17915), .Z(n17910) );
  AND U17425 ( .A(n17916), .B(n17917), .Z(n17915) );
  XNOR U17426 ( .A(p_input[6136]), .B(n17914), .Z(n17917) );
  XOR U17427 ( .A(n17914), .B(p_input[6104]), .Z(n17916) );
  XOR U17428 ( .A(n17918), .B(n17919), .Z(n17914) );
  AND U17429 ( .A(n17920), .B(n17921), .Z(n17919) );
  XNOR U17430 ( .A(p_input[6135]), .B(n17918), .Z(n17921) );
  XOR U17431 ( .A(n17918), .B(p_input[6103]), .Z(n17920) );
  XOR U17432 ( .A(n17922), .B(n17923), .Z(n17918) );
  AND U17433 ( .A(n17924), .B(n17925), .Z(n17923) );
  XNOR U17434 ( .A(p_input[6134]), .B(n17922), .Z(n17925) );
  XOR U17435 ( .A(n17922), .B(p_input[6102]), .Z(n17924) );
  XOR U17436 ( .A(n17926), .B(n17927), .Z(n17922) );
  AND U17437 ( .A(n17928), .B(n17929), .Z(n17927) );
  XNOR U17438 ( .A(p_input[6133]), .B(n17926), .Z(n17929) );
  XOR U17439 ( .A(n17926), .B(p_input[6101]), .Z(n17928) );
  XOR U17440 ( .A(n17930), .B(n17931), .Z(n17926) );
  AND U17441 ( .A(n17932), .B(n17933), .Z(n17931) );
  XNOR U17442 ( .A(p_input[6132]), .B(n17930), .Z(n17933) );
  XOR U17443 ( .A(n17930), .B(p_input[6100]), .Z(n17932) );
  XOR U17444 ( .A(n17934), .B(n17935), .Z(n17930) );
  AND U17445 ( .A(n17936), .B(n17937), .Z(n17935) );
  XNOR U17446 ( .A(p_input[6131]), .B(n17934), .Z(n17937) );
  XOR U17447 ( .A(n17934), .B(p_input[6099]), .Z(n17936) );
  XOR U17448 ( .A(n17938), .B(n17939), .Z(n17934) );
  AND U17449 ( .A(n17940), .B(n17941), .Z(n17939) );
  XNOR U17450 ( .A(p_input[6130]), .B(n17938), .Z(n17941) );
  XOR U17451 ( .A(n17938), .B(p_input[6098]), .Z(n17940) );
  XOR U17452 ( .A(n17942), .B(n17943), .Z(n17938) );
  AND U17453 ( .A(n17944), .B(n17945), .Z(n17943) );
  XNOR U17454 ( .A(p_input[6129]), .B(n17942), .Z(n17945) );
  XOR U17455 ( .A(n17942), .B(p_input[6097]), .Z(n17944) );
  XOR U17456 ( .A(n17946), .B(n17947), .Z(n17942) );
  AND U17457 ( .A(n17948), .B(n17949), .Z(n17947) );
  XNOR U17458 ( .A(p_input[6128]), .B(n17946), .Z(n17949) );
  XOR U17459 ( .A(n17946), .B(p_input[6096]), .Z(n17948) );
  XOR U17460 ( .A(n17950), .B(n17951), .Z(n17946) );
  AND U17461 ( .A(n17952), .B(n17953), .Z(n17951) );
  XNOR U17462 ( .A(p_input[6127]), .B(n17950), .Z(n17953) );
  XOR U17463 ( .A(n17950), .B(p_input[6095]), .Z(n17952) );
  XOR U17464 ( .A(n17954), .B(n17955), .Z(n17950) );
  AND U17465 ( .A(n17956), .B(n17957), .Z(n17955) );
  XNOR U17466 ( .A(p_input[6126]), .B(n17954), .Z(n17957) );
  XOR U17467 ( .A(n17954), .B(p_input[6094]), .Z(n17956) );
  XOR U17468 ( .A(n17958), .B(n17959), .Z(n17954) );
  AND U17469 ( .A(n17960), .B(n17961), .Z(n17959) );
  XNOR U17470 ( .A(p_input[6125]), .B(n17958), .Z(n17961) );
  XOR U17471 ( .A(n17958), .B(p_input[6093]), .Z(n17960) );
  XOR U17472 ( .A(n17962), .B(n17963), .Z(n17958) );
  AND U17473 ( .A(n17964), .B(n17965), .Z(n17963) );
  XNOR U17474 ( .A(p_input[6124]), .B(n17962), .Z(n17965) );
  XOR U17475 ( .A(n17962), .B(p_input[6092]), .Z(n17964) );
  XOR U17476 ( .A(n17966), .B(n17967), .Z(n17962) );
  AND U17477 ( .A(n17968), .B(n17969), .Z(n17967) );
  XNOR U17478 ( .A(p_input[6123]), .B(n17966), .Z(n17969) );
  XOR U17479 ( .A(n17966), .B(p_input[6091]), .Z(n17968) );
  XOR U17480 ( .A(n17970), .B(n17971), .Z(n17966) );
  AND U17481 ( .A(n17972), .B(n17973), .Z(n17971) );
  XNOR U17482 ( .A(p_input[6122]), .B(n17970), .Z(n17973) );
  XOR U17483 ( .A(n17970), .B(p_input[6090]), .Z(n17972) );
  XOR U17484 ( .A(n17974), .B(n17975), .Z(n17970) );
  AND U17485 ( .A(n17976), .B(n17977), .Z(n17975) );
  XNOR U17486 ( .A(p_input[6121]), .B(n17974), .Z(n17977) );
  XOR U17487 ( .A(n17974), .B(p_input[6089]), .Z(n17976) );
  XOR U17488 ( .A(n17978), .B(n17979), .Z(n17974) );
  AND U17489 ( .A(n17980), .B(n17981), .Z(n17979) );
  XNOR U17490 ( .A(p_input[6120]), .B(n17978), .Z(n17981) );
  XOR U17491 ( .A(n17978), .B(p_input[6088]), .Z(n17980) );
  XOR U17492 ( .A(n17982), .B(n17983), .Z(n17978) );
  AND U17493 ( .A(n17984), .B(n17985), .Z(n17983) );
  XNOR U17494 ( .A(p_input[6119]), .B(n17982), .Z(n17985) );
  XOR U17495 ( .A(n17982), .B(p_input[6087]), .Z(n17984) );
  XOR U17496 ( .A(n17986), .B(n17987), .Z(n17982) );
  AND U17497 ( .A(n17988), .B(n17989), .Z(n17987) );
  XNOR U17498 ( .A(p_input[6118]), .B(n17986), .Z(n17989) );
  XOR U17499 ( .A(n17986), .B(p_input[6086]), .Z(n17988) );
  XOR U17500 ( .A(n17990), .B(n17991), .Z(n17986) );
  AND U17501 ( .A(n17992), .B(n17993), .Z(n17991) );
  XNOR U17502 ( .A(p_input[6117]), .B(n17990), .Z(n17993) );
  XOR U17503 ( .A(n17990), .B(p_input[6085]), .Z(n17992) );
  XOR U17504 ( .A(n17994), .B(n17995), .Z(n17990) );
  AND U17505 ( .A(n17996), .B(n17997), .Z(n17995) );
  XNOR U17506 ( .A(p_input[6116]), .B(n17994), .Z(n17997) );
  XOR U17507 ( .A(n17994), .B(p_input[6084]), .Z(n17996) );
  XOR U17508 ( .A(n17998), .B(n17999), .Z(n17994) );
  AND U17509 ( .A(n18000), .B(n18001), .Z(n17999) );
  XNOR U17510 ( .A(p_input[6115]), .B(n17998), .Z(n18001) );
  XOR U17511 ( .A(n17998), .B(p_input[6083]), .Z(n18000) );
  XOR U17512 ( .A(n18002), .B(n18003), .Z(n17998) );
  AND U17513 ( .A(n18004), .B(n18005), .Z(n18003) );
  XNOR U17514 ( .A(p_input[6114]), .B(n18002), .Z(n18005) );
  XOR U17515 ( .A(n18002), .B(p_input[6082]), .Z(n18004) );
  XNOR U17516 ( .A(n18006), .B(n18007), .Z(n18002) );
  AND U17517 ( .A(n18008), .B(n18009), .Z(n18007) );
  XOR U17518 ( .A(p_input[6113]), .B(n18006), .Z(n18009) );
  XNOR U17519 ( .A(p_input[6081]), .B(n18006), .Z(n18008) );
  AND U17520 ( .A(p_input[6112]), .B(n18010), .Z(n18006) );
  IV U17521 ( .A(p_input[6080]), .Z(n18010) );
  XNOR U17522 ( .A(p_input[6016]), .B(n18011), .Z(n17604) );
  AND U17523 ( .A(n309), .B(n18012), .Z(n18011) );
  XOR U17524 ( .A(p_input[6048]), .B(p_input[6016]), .Z(n18012) );
  XOR U17525 ( .A(n18013), .B(n18014), .Z(n309) );
  AND U17526 ( .A(n18015), .B(n18016), .Z(n18014) );
  XNOR U17527 ( .A(p_input[6079]), .B(n18013), .Z(n18016) );
  XOR U17528 ( .A(n18013), .B(p_input[6047]), .Z(n18015) );
  XOR U17529 ( .A(n18017), .B(n18018), .Z(n18013) );
  AND U17530 ( .A(n18019), .B(n18020), .Z(n18018) );
  XNOR U17531 ( .A(p_input[6078]), .B(n18017), .Z(n18020) );
  XNOR U17532 ( .A(n18017), .B(n17619), .Z(n18019) );
  IV U17533 ( .A(p_input[6046]), .Z(n17619) );
  XOR U17534 ( .A(n18021), .B(n18022), .Z(n18017) );
  AND U17535 ( .A(n18023), .B(n18024), .Z(n18022) );
  XNOR U17536 ( .A(p_input[6077]), .B(n18021), .Z(n18024) );
  XNOR U17537 ( .A(n18021), .B(n17628), .Z(n18023) );
  IV U17538 ( .A(p_input[6045]), .Z(n17628) );
  XOR U17539 ( .A(n18025), .B(n18026), .Z(n18021) );
  AND U17540 ( .A(n18027), .B(n18028), .Z(n18026) );
  XNOR U17541 ( .A(p_input[6076]), .B(n18025), .Z(n18028) );
  XNOR U17542 ( .A(n18025), .B(n17637), .Z(n18027) );
  IV U17543 ( .A(p_input[6044]), .Z(n17637) );
  XOR U17544 ( .A(n18029), .B(n18030), .Z(n18025) );
  AND U17545 ( .A(n18031), .B(n18032), .Z(n18030) );
  XNOR U17546 ( .A(p_input[6075]), .B(n18029), .Z(n18032) );
  XNOR U17547 ( .A(n18029), .B(n17646), .Z(n18031) );
  IV U17548 ( .A(p_input[6043]), .Z(n17646) );
  XOR U17549 ( .A(n18033), .B(n18034), .Z(n18029) );
  AND U17550 ( .A(n18035), .B(n18036), .Z(n18034) );
  XNOR U17551 ( .A(p_input[6074]), .B(n18033), .Z(n18036) );
  XNOR U17552 ( .A(n18033), .B(n17655), .Z(n18035) );
  IV U17553 ( .A(p_input[6042]), .Z(n17655) );
  XOR U17554 ( .A(n18037), .B(n18038), .Z(n18033) );
  AND U17555 ( .A(n18039), .B(n18040), .Z(n18038) );
  XNOR U17556 ( .A(p_input[6073]), .B(n18037), .Z(n18040) );
  XNOR U17557 ( .A(n18037), .B(n17664), .Z(n18039) );
  IV U17558 ( .A(p_input[6041]), .Z(n17664) );
  XOR U17559 ( .A(n18041), .B(n18042), .Z(n18037) );
  AND U17560 ( .A(n18043), .B(n18044), .Z(n18042) );
  XNOR U17561 ( .A(p_input[6072]), .B(n18041), .Z(n18044) );
  XNOR U17562 ( .A(n18041), .B(n17673), .Z(n18043) );
  IV U17563 ( .A(p_input[6040]), .Z(n17673) );
  XOR U17564 ( .A(n18045), .B(n18046), .Z(n18041) );
  AND U17565 ( .A(n18047), .B(n18048), .Z(n18046) );
  XNOR U17566 ( .A(p_input[6071]), .B(n18045), .Z(n18048) );
  XNOR U17567 ( .A(n18045), .B(n17682), .Z(n18047) );
  IV U17568 ( .A(p_input[6039]), .Z(n17682) );
  XOR U17569 ( .A(n18049), .B(n18050), .Z(n18045) );
  AND U17570 ( .A(n18051), .B(n18052), .Z(n18050) );
  XNOR U17571 ( .A(p_input[6070]), .B(n18049), .Z(n18052) );
  XNOR U17572 ( .A(n18049), .B(n17691), .Z(n18051) );
  IV U17573 ( .A(p_input[6038]), .Z(n17691) );
  XOR U17574 ( .A(n18053), .B(n18054), .Z(n18049) );
  AND U17575 ( .A(n18055), .B(n18056), .Z(n18054) );
  XNOR U17576 ( .A(p_input[6069]), .B(n18053), .Z(n18056) );
  XNOR U17577 ( .A(n18053), .B(n17700), .Z(n18055) );
  IV U17578 ( .A(p_input[6037]), .Z(n17700) );
  XOR U17579 ( .A(n18057), .B(n18058), .Z(n18053) );
  AND U17580 ( .A(n18059), .B(n18060), .Z(n18058) );
  XNOR U17581 ( .A(p_input[6068]), .B(n18057), .Z(n18060) );
  XNOR U17582 ( .A(n18057), .B(n17709), .Z(n18059) );
  IV U17583 ( .A(p_input[6036]), .Z(n17709) );
  XOR U17584 ( .A(n18061), .B(n18062), .Z(n18057) );
  AND U17585 ( .A(n18063), .B(n18064), .Z(n18062) );
  XNOR U17586 ( .A(p_input[6067]), .B(n18061), .Z(n18064) );
  XNOR U17587 ( .A(n18061), .B(n17718), .Z(n18063) );
  IV U17588 ( .A(p_input[6035]), .Z(n17718) );
  XOR U17589 ( .A(n18065), .B(n18066), .Z(n18061) );
  AND U17590 ( .A(n18067), .B(n18068), .Z(n18066) );
  XNOR U17591 ( .A(p_input[6066]), .B(n18065), .Z(n18068) );
  XNOR U17592 ( .A(n18065), .B(n17727), .Z(n18067) );
  IV U17593 ( .A(p_input[6034]), .Z(n17727) );
  XOR U17594 ( .A(n18069), .B(n18070), .Z(n18065) );
  AND U17595 ( .A(n18071), .B(n18072), .Z(n18070) );
  XNOR U17596 ( .A(p_input[6065]), .B(n18069), .Z(n18072) );
  XNOR U17597 ( .A(n18069), .B(n17736), .Z(n18071) );
  IV U17598 ( .A(p_input[6033]), .Z(n17736) );
  XOR U17599 ( .A(n18073), .B(n18074), .Z(n18069) );
  AND U17600 ( .A(n18075), .B(n18076), .Z(n18074) );
  XNOR U17601 ( .A(p_input[6064]), .B(n18073), .Z(n18076) );
  XNOR U17602 ( .A(n18073), .B(n17745), .Z(n18075) );
  IV U17603 ( .A(p_input[6032]), .Z(n17745) );
  XOR U17604 ( .A(n18077), .B(n18078), .Z(n18073) );
  AND U17605 ( .A(n18079), .B(n18080), .Z(n18078) );
  XNOR U17606 ( .A(p_input[6063]), .B(n18077), .Z(n18080) );
  XNOR U17607 ( .A(n18077), .B(n17754), .Z(n18079) );
  IV U17608 ( .A(p_input[6031]), .Z(n17754) );
  XOR U17609 ( .A(n18081), .B(n18082), .Z(n18077) );
  AND U17610 ( .A(n18083), .B(n18084), .Z(n18082) );
  XNOR U17611 ( .A(p_input[6062]), .B(n18081), .Z(n18084) );
  XNOR U17612 ( .A(n18081), .B(n17763), .Z(n18083) );
  IV U17613 ( .A(p_input[6030]), .Z(n17763) );
  XOR U17614 ( .A(n18085), .B(n18086), .Z(n18081) );
  AND U17615 ( .A(n18087), .B(n18088), .Z(n18086) );
  XNOR U17616 ( .A(p_input[6061]), .B(n18085), .Z(n18088) );
  XNOR U17617 ( .A(n18085), .B(n17772), .Z(n18087) );
  IV U17618 ( .A(p_input[6029]), .Z(n17772) );
  XOR U17619 ( .A(n18089), .B(n18090), .Z(n18085) );
  AND U17620 ( .A(n18091), .B(n18092), .Z(n18090) );
  XNOR U17621 ( .A(p_input[6060]), .B(n18089), .Z(n18092) );
  XNOR U17622 ( .A(n18089), .B(n17781), .Z(n18091) );
  IV U17623 ( .A(p_input[6028]), .Z(n17781) );
  XOR U17624 ( .A(n18093), .B(n18094), .Z(n18089) );
  AND U17625 ( .A(n18095), .B(n18096), .Z(n18094) );
  XNOR U17626 ( .A(p_input[6059]), .B(n18093), .Z(n18096) );
  XNOR U17627 ( .A(n18093), .B(n17790), .Z(n18095) );
  IV U17628 ( .A(p_input[6027]), .Z(n17790) );
  XOR U17629 ( .A(n18097), .B(n18098), .Z(n18093) );
  AND U17630 ( .A(n18099), .B(n18100), .Z(n18098) );
  XNOR U17631 ( .A(p_input[6058]), .B(n18097), .Z(n18100) );
  XNOR U17632 ( .A(n18097), .B(n17799), .Z(n18099) );
  IV U17633 ( .A(p_input[6026]), .Z(n17799) );
  XOR U17634 ( .A(n18101), .B(n18102), .Z(n18097) );
  AND U17635 ( .A(n18103), .B(n18104), .Z(n18102) );
  XNOR U17636 ( .A(p_input[6057]), .B(n18101), .Z(n18104) );
  XNOR U17637 ( .A(n18101), .B(n17808), .Z(n18103) );
  IV U17638 ( .A(p_input[6025]), .Z(n17808) );
  XOR U17639 ( .A(n18105), .B(n18106), .Z(n18101) );
  AND U17640 ( .A(n18107), .B(n18108), .Z(n18106) );
  XNOR U17641 ( .A(p_input[6056]), .B(n18105), .Z(n18108) );
  XNOR U17642 ( .A(n18105), .B(n17817), .Z(n18107) );
  IV U17643 ( .A(p_input[6024]), .Z(n17817) );
  XOR U17644 ( .A(n18109), .B(n18110), .Z(n18105) );
  AND U17645 ( .A(n18111), .B(n18112), .Z(n18110) );
  XNOR U17646 ( .A(p_input[6055]), .B(n18109), .Z(n18112) );
  XNOR U17647 ( .A(n18109), .B(n17826), .Z(n18111) );
  IV U17648 ( .A(p_input[6023]), .Z(n17826) );
  XOR U17649 ( .A(n18113), .B(n18114), .Z(n18109) );
  AND U17650 ( .A(n18115), .B(n18116), .Z(n18114) );
  XNOR U17651 ( .A(p_input[6054]), .B(n18113), .Z(n18116) );
  XNOR U17652 ( .A(n18113), .B(n17835), .Z(n18115) );
  IV U17653 ( .A(p_input[6022]), .Z(n17835) );
  XOR U17654 ( .A(n18117), .B(n18118), .Z(n18113) );
  AND U17655 ( .A(n18119), .B(n18120), .Z(n18118) );
  XNOR U17656 ( .A(p_input[6053]), .B(n18117), .Z(n18120) );
  XNOR U17657 ( .A(n18117), .B(n17844), .Z(n18119) );
  IV U17658 ( .A(p_input[6021]), .Z(n17844) );
  XOR U17659 ( .A(n18121), .B(n18122), .Z(n18117) );
  AND U17660 ( .A(n18123), .B(n18124), .Z(n18122) );
  XNOR U17661 ( .A(p_input[6052]), .B(n18121), .Z(n18124) );
  XNOR U17662 ( .A(n18121), .B(n17853), .Z(n18123) );
  IV U17663 ( .A(p_input[6020]), .Z(n17853) );
  XOR U17664 ( .A(n18125), .B(n18126), .Z(n18121) );
  AND U17665 ( .A(n18127), .B(n18128), .Z(n18126) );
  XNOR U17666 ( .A(p_input[6051]), .B(n18125), .Z(n18128) );
  XNOR U17667 ( .A(n18125), .B(n17862), .Z(n18127) );
  IV U17668 ( .A(p_input[6019]), .Z(n17862) );
  XOR U17669 ( .A(n18129), .B(n18130), .Z(n18125) );
  AND U17670 ( .A(n18131), .B(n18132), .Z(n18130) );
  XNOR U17671 ( .A(p_input[6050]), .B(n18129), .Z(n18132) );
  XNOR U17672 ( .A(n18129), .B(n17871), .Z(n18131) );
  IV U17673 ( .A(p_input[6018]), .Z(n17871) );
  XNOR U17674 ( .A(n18133), .B(n18134), .Z(n18129) );
  AND U17675 ( .A(n18135), .B(n18136), .Z(n18134) );
  XOR U17676 ( .A(p_input[6049]), .B(n18133), .Z(n18136) );
  XNOR U17677 ( .A(p_input[6017]), .B(n18133), .Z(n18135) );
  AND U17678 ( .A(p_input[6048]), .B(n18137), .Z(n18133) );
  IV U17679 ( .A(p_input[6016]), .Z(n18137) );
  XOR U17680 ( .A(n18138), .B(n18139), .Z(n17227) );
  AND U17681 ( .A(n497), .B(n18140), .Z(n18139) );
  XNOR U17682 ( .A(n18141), .B(n18138), .Z(n18140) );
  XOR U17683 ( .A(n18142), .B(n18143), .Z(n497) );
  AND U17684 ( .A(n18144), .B(n18145), .Z(n18143) );
  XNOR U17685 ( .A(n17242), .B(n18142), .Z(n18145) );
  AND U17686 ( .A(p_input[6015]), .B(p_input[5983]), .Z(n17242) );
  XNOR U17687 ( .A(n18142), .B(n17239), .Z(n18144) );
  IV U17688 ( .A(n18146), .Z(n17239) );
  AND U17689 ( .A(p_input[5919]), .B(p_input[5951]), .Z(n18146) );
  XOR U17690 ( .A(n18147), .B(n18148), .Z(n18142) );
  AND U17691 ( .A(n18149), .B(n18150), .Z(n18148) );
  XOR U17692 ( .A(n18147), .B(n17254), .Z(n18150) );
  XNOR U17693 ( .A(p_input[5982]), .B(n18151), .Z(n17254) );
  AND U17694 ( .A(n315), .B(n18152), .Z(n18151) );
  XOR U17695 ( .A(p_input[6014]), .B(p_input[5982]), .Z(n18152) );
  XNOR U17696 ( .A(n17251), .B(n18147), .Z(n18149) );
  XOR U17697 ( .A(n18153), .B(n18154), .Z(n17251) );
  AND U17698 ( .A(n312), .B(n18155), .Z(n18154) );
  XOR U17699 ( .A(p_input[5950]), .B(p_input[5918]), .Z(n18155) );
  XOR U17700 ( .A(n18156), .B(n18157), .Z(n18147) );
  AND U17701 ( .A(n18158), .B(n18159), .Z(n18157) );
  XOR U17702 ( .A(n18156), .B(n17266), .Z(n18159) );
  XNOR U17703 ( .A(p_input[5981]), .B(n18160), .Z(n17266) );
  AND U17704 ( .A(n315), .B(n18161), .Z(n18160) );
  XOR U17705 ( .A(p_input[6013]), .B(p_input[5981]), .Z(n18161) );
  XNOR U17706 ( .A(n17263), .B(n18156), .Z(n18158) );
  XOR U17707 ( .A(n18162), .B(n18163), .Z(n17263) );
  AND U17708 ( .A(n312), .B(n18164), .Z(n18163) );
  XOR U17709 ( .A(p_input[5949]), .B(p_input[5917]), .Z(n18164) );
  XOR U17710 ( .A(n18165), .B(n18166), .Z(n18156) );
  AND U17711 ( .A(n18167), .B(n18168), .Z(n18166) );
  XOR U17712 ( .A(n18165), .B(n17278), .Z(n18168) );
  XNOR U17713 ( .A(p_input[5980]), .B(n18169), .Z(n17278) );
  AND U17714 ( .A(n315), .B(n18170), .Z(n18169) );
  XOR U17715 ( .A(p_input[6012]), .B(p_input[5980]), .Z(n18170) );
  XNOR U17716 ( .A(n17275), .B(n18165), .Z(n18167) );
  XOR U17717 ( .A(n18171), .B(n18172), .Z(n17275) );
  AND U17718 ( .A(n312), .B(n18173), .Z(n18172) );
  XOR U17719 ( .A(p_input[5948]), .B(p_input[5916]), .Z(n18173) );
  XOR U17720 ( .A(n18174), .B(n18175), .Z(n18165) );
  AND U17721 ( .A(n18176), .B(n18177), .Z(n18175) );
  XOR U17722 ( .A(n18174), .B(n17290), .Z(n18177) );
  XNOR U17723 ( .A(p_input[5979]), .B(n18178), .Z(n17290) );
  AND U17724 ( .A(n315), .B(n18179), .Z(n18178) );
  XOR U17725 ( .A(p_input[6011]), .B(p_input[5979]), .Z(n18179) );
  XNOR U17726 ( .A(n17287), .B(n18174), .Z(n18176) );
  XOR U17727 ( .A(n18180), .B(n18181), .Z(n17287) );
  AND U17728 ( .A(n312), .B(n18182), .Z(n18181) );
  XOR U17729 ( .A(p_input[5947]), .B(p_input[5915]), .Z(n18182) );
  XOR U17730 ( .A(n18183), .B(n18184), .Z(n18174) );
  AND U17731 ( .A(n18185), .B(n18186), .Z(n18184) );
  XOR U17732 ( .A(n18183), .B(n17302), .Z(n18186) );
  XNOR U17733 ( .A(p_input[5978]), .B(n18187), .Z(n17302) );
  AND U17734 ( .A(n315), .B(n18188), .Z(n18187) );
  XOR U17735 ( .A(p_input[6010]), .B(p_input[5978]), .Z(n18188) );
  XNOR U17736 ( .A(n17299), .B(n18183), .Z(n18185) );
  XOR U17737 ( .A(n18189), .B(n18190), .Z(n17299) );
  AND U17738 ( .A(n312), .B(n18191), .Z(n18190) );
  XOR U17739 ( .A(p_input[5946]), .B(p_input[5914]), .Z(n18191) );
  XOR U17740 ( .A(n18192), .B(n18193), .Z(n18183) );
  AND U17741 ( .A(n18194), .B(n18195), .Z(n18193) );
  XOR U17742 ( .A(n18192), .B(n17314), .Z(n18195) );
  XNOR U17743 ( .A(p_input[5977]), .B(n18196), .Z(n17314) );
  AND U17744 ( .A(n315), .B(n18197), .Z(n18196) );
  XOR U17745 ( .A(p_input[6009]), .B(p_input[5977]), .Z(n18197) );
  XNOR U17746 ( .A(n17311), .B(n18192), .Z(n18194) );
  XOR U17747 ( .A(n18198), .B(n18199), .Z(n17311) );
  AND U17748 ( .A(n312), .B(n18200), .Z(n18199) );
  XOR U17749 ( .A(p_input[5945]), .B(p_input[5913]), .Z(n18200) );
  XOR U17750 ( .A(n18201), .B(n18202), .Z(n18192) );
  AND U17751 ( .A(n18203), .B(n18204), .Z(n18202) );
  XOR U17752 ( .A(n18201), .B(n17326), .Z(n18204) );
  XNOR U17753 ( .A(p_input[5976]), .B(n18205), .Z(n17326) );
  AND U17754 ( .A(n315), .B(n18206), .Z(n18205) );
  XOR U17755 ( .A(p_input[6008]), .B(p_input[5976]), .Z(n18206) );
  XNOR U17756 ( .A(n17323), .B(n18201), .Z(n18203) );
  XOR U17757 ( .A(n18207), .B(n18208), .Z(n17323) );
  AND U17758 ( .A(n312), .B(n18209), .Z(n18208) );
  XOR U17759 ( .A(p_input[5944]), .B(p_input[5912]), .Z(n18209) );
  XOR U17760 ( .A(n18210), .B(n18211), .Z(n18201) );
  AND U17761 ( .A(n18212), .B(n18213), .Z(n18211) );
  XOR U17762 ( .A(n18210), .B(n17338), .Z(n18213) );
  XNOR U17763 ( .A(p_input[5975]), .B(n18214), .Z(n17338) );
  AND U17764 ( .A(n315), .B(n18215), .Z(n18214) );
  XOR U17765 ( .A(p_input[6007]), .B(p_input[5975]), .Z(n18215) );
  XNOR U17766 ( .A(n17335), .B(n18210), .Z(n18212) );
  XOR U17767 ( .A(n18216), .B(n18217), .Z(n17335) );
  AND U17768 ( .A(n312), .B(n18218), .Z(n18217) );
  XOR U17769 ( .A(p_input[5943]), .B(p_input[5911]), .Z(n18218) );
  XOR U17770 ( .A(n18219), .B(n18220), .Z(n18210) );
  AND U17771 ( .A(n18221), .B(n18222), .Z(n18220) );
  XOR U17772 ( .A(n18219), .B(n17350), .Z(n18222) );
  XNOR U17773 ( .A(p_input[5974]), .B(n18223), .Z(n17350) );
  AND U17774 ( .A(n315), .B(n18224), .Z(n18223) );
  XOR U17775 ( .A(p_input[6006]), .B(p_input[5974]), .Z(n18224) );
  XNOR U17776 ( .A(n17347), .B(n18219), .Z(n18221) );
  XOR U17777 ( .A(n18225), .B(n18226), .Z(n17347) );
  AND U17778 ( .A(n312), .B(n18227), .Z(n18226) );
  XOR U17779 ( .A(p_input[5942]), .B(p_input[5910]), .Z(n18227) );
  XOR U17780 ( .A(n18228), .B(n18229), .Z(n18219) );
  AND U17781 ( .A(n18230), .B(n18231), .Z(n18229) );
  XOR U17782 ( .A(n18228), .B(n17362), .Z(n18231) );
  XNOR U17783 ( .A(p_input[5973]), .B(n18232), .Z(n17362) );
  AND U17784 ( .A(n315), .B(n18233), .Z(n18232) );
  XOR U17785 ( .A(p_input[6005]), .B(p_input[5973]), .Z(n18233) );
  XNOR U17786 ( .A(n17359), .B(n18228), .Z(n18230) );
  XOR U17787 ( .A(n18234), .B(n18235), .Z(n17359) );
  AND U17788 ( .A(n312), .B(n18236), .Z(n18235) );
  XOR U17789 ( .A(p_input[5941]), .B(p_input[5909]), .Z(n18236) );
  XOR U17790 ( .A(n18237), .B(n18238), .Z(n18228) );
  AND U17791 ( .A(n18239), .B(n18240), .Z(n18238) );
  XOR U17792 ( .A(n18237), .B(n17374), .Z(n18240) );
  XNOR U17793 ( .A(p_input[5972]), .B(n18241), .Z(n17374) );
  AND U17794 ( .A(n315), .B(n18242), .Z(n18241) );
  XOR U17795 ( .A(p_input[6004]), .B(p_input[5972]), .Z(n18242) );
  XNOR U17796 ( .A(n17371), .B(n18237), .Z(n18239) );
  XOR U17797 ( .A(n18243), .B(n18244), .Z(n17371) );
  AND U17798 ( .A(n312), .B(n18245), .Z(n18244) );
  XOR U17799 ( .A(p_input[5940]), .B(p_input[5908]), .Z(n18245) );
  XOR U17800 ( .A(n18246), .B(n18247), .Z(n18237) );
  AND U17801 ( .A(n18248), .B(n18249), .Z(n18247) );
  XOR U17802 ( .A(n18246), .B(n17386), .Z(n18249) );
  XNOR U17803 ( .A(p_input[5971]), .B(n18250), .Z(n17386) );
  AND U17804 ( .A(n315), .B(n18251), .Z(n18250) );
  XOR U17805 ( .A(p_input[6003]), .B(p_input[5971]), .Z(n18251) );
  XNOR U17806 ( .A(n17383), .B(n18246), .Z(n18248) );
  XOR U17807 ( .A(n18252), .B(n18253), .Z(n17383) );
  AND U17808 ( .A(n312), .B(n18254), .Z(n18253) );
  XOR U17809 ( .A(p_input[5939]), .B(p_input[5907]), .Z(n18254) );
  XOR U17810 ( .A(n18255), .B(n18256), .Z(n18246) );
  AND U17811 ( .A(n18257), .B(n18258), .Z(n18256) );
  XOR U17812 ( .A(n18255), .B(n17398), .Z(n18258) );
  XNOR U17813 ( .A(p_input[5970]), .B(n18259), .Z(n17398) );
  AND U17814 ( .A(n315), .B(n18260), .Z(n18259) );
  XOR U17815 ( .A(p_input[6002]), .B(p_input[5970]), .Z(n18260) );
  XNOR U17816 ( .A(n17395), .B(n18255), .Z(n18257) );
  XOR U17817 ( .A(n18261), .B(n18262), .Z(n17395) );
  AND U17818 ( .A(n312), .B(n18263), .Z(n18262) );
  XOR U17819 ( .A(p_input[5938]), .B(p_input[5906]), .Z(n18263) );
  XOR U17820 ( .A(n18264), .B(n18265), .Z(n18255) );
  AND U17821 ( .A(n18266), .B(n18267), .Z(n18265) );
  XOR U17822 ( .A(n18264), .B(n17410), .Z(n18267) );
  XNOR U17823 ( .A(p_input[5969]), .B(n18268), .Z(n17410) );
  AND U17824 ( .A(n315), .B(n18269), .Z(n18268) );
  XOR U17825 ( .A(p_input[6001]), .B(p_input[5969]), .Z(n18269) );
  XNOR U17826 ( .A(n17407), .B(n18264), .Z(n18266) );
  XOR U17827 ( .A(n18270), .B(n18271), .Z(n17407) );
  AND U17828 ( .A(n312), .B(n18272), .Z(n18271) );
  XOR U17829 ( .A(p_input[5937]), .B(p_input[5905]), .Z(n18272) );
  XOR U17830 ( .A(n18273), .B(n18274), .Z(n18264) );
  AND U17831 ( .A(n18275), .B(n18276), .Z(n18274) );
  XOR U17832 ( .A(n18273), .B(n17422), .Z(n18276) );
  XNOR U17833 ( .A(p_input[5968]), .B(n18277), .Z(n17422) );
  AND U17834 ( .A(n315), .B(n18278), .Z(n18277) );
  XOR U17835 ( .A(p_input[6000]), .B(p_input[5968]), .Z(n18278) );
  XNOR U17836 ( .A(n17419), .B(n18273), .Z(n18275) );
  XOR U17837 ( .A(n18279), .B(n18280), .Z(n17419) );
  AND U17838 ( .A(n312), .B(n18281), .Z(n18280) );
  XOR U17839 ( .A(p_input[5936]), .B(p_input[5904]), .Z(n18281) );
  XOR U17840 ( .A(n18282), .B(n18283), .Z(n18273) );
  AND U17841 ( .A(n18284), .B(n18285), .Z(n18283) );
  XOR U17842 ( .A(n18282), .B(n17434), .Z(n18285) );
  XNOR U17843 ( .A(p_input[5967]), .B(n18286), .Z(n17434) );
  AND U17844 ( .A(n315), .B(n18287), .Z(n18286) );
  XOR U17845 ( .A(p_input[5999]), .B(p_input[5967]), .Z(n18287) );
  XNOR U17846 ( .A(n17431), .B(n18282), .Z(n18284) );
  XOR U17847 ( .A(n18288), .B(n18289), .Z(n17431) );
  AND U17848 ( .A(n312), .B(n18290), .Z(n18289) );
  XOR U17849 ( .A(p_input[5935]), .B(p_input[5903]), .Z(n18290) );
  XOR U17850 ( .A(n18291), .B(n18292), .Z(n18282) );
  AND U17851 ( .A(n18293), .B(n18294), .Z(n18292) );
  XOR U17852 ( .A(n18291), .B(n17446), .Z(n18294) );
  XNOR U17853 ( .A(p_input[5966]), .B(n18295), .Z(n17446) );
  AND U17854 ( .A(n315), .B(n18296), .Z(n18295) );
  XOR U17855 ( .A(p_input[5998]), .B(p_input[5966]), .Z(n18296) );
  XNOR U17856 ( .A(n17443), .B(n18291), .Z(n18293) );
  XOR U17857 ( .A(n18297), .B(n18298), .Z(n17443) );
  AND U17858 ( .A(n312), .B(n18299), .Z(n18298) );
  XOR U17859 ( .A(p_input[5934]), .B(p_input[5902]), .Z(n18299) );
  XOR U17860 ( .A(n18300), .B(n18301), .Z(n18291) );
  AND U17861 ( .A(n18302), .B(n18303), .Z(n18301) );
  XOR U17862 ( .A(n18300), .B(n17458), .Z(n18303) );
  XNOR U17863 ( .A(p_input[5965]), .B(n18304), .Z(n17458) );
  AND U17864 ( .A(n315), .B(n18305), .Z(n18304) );
  XOR U17865 ( .A(p_input[5997]), .B(p_input[5965]), .Z(n18305) );
  XNOR U17866 ( .A(n17455), .B(n18300), .Z(n18302) );
  XOR U17867 ( .A(n18306), .B(n18307), .Z(n17455) );
  AND U17868 ( .A(n312), .B(n18308), .Z(n18307) );
  XOR U17869 ( .A(p_input[5933]), .B(p_input[5901]), .Z(n18308) );
  XOR U17870 ( .A(n18309), .B(n18310), .Z(n18300) );
  AND U17871 ( .A(n18311), .B(n18312), .Z(n18310) );
  XOR U17872 ( .A(n18309), .B(n17470), .Z(n18312) );
  XNOR U17873 ( .A(p_input[5964]), .B(n18313), .Z(n17470) );
  AND U17874 ( .A(n315), .B(n18314), .Z(n18313) );
  XOR U17875 ( .A(p_input[5996]), .B(p_input[5964]), .Z(n18314) );
  XNOR U17876 ( .A(n17467), .B(n18309), .Z(n18311) );
  XOR U17877 ( .A(n18315), .B(n18316), .Z(n17467) );
  AND U17878 ( .A(n312), .B(n18317), .Z(n18316) );
  XOR U17879 ( .A(p_input[5932]), .B(p_input[5900]), .Z(n18317) );
  XOR U17880 ( .A(n18318), .B(n18319), .Z(n18309) );
  AND U17881 ( .A(n18320), .B(n18321), .Z(n18319) );
  XOR U17882 ( .A(n18318), .B(n17482), .Z(n18321) );
  XNOR U17883 ( .A(p_input[5963]), .B(n18322), .Z(n17482) );
  AND U17884 ( .A(n315), .B(n18323), .Z(n18322) );
  XOR U17885 ( .A(p_input[5995]), .B(p_input[5963]), .Z(n18323) );
  XNOR U17886 ( .A(n17479), .B(n18318), .Z(n18320) );
  XOR U17887 ( .A(n18324), .B(n18325), .Z(n17479) );
  AND U17888 ( .A(n312), .B(n18326), .Z(n18325) );
  XOR U17889 ( .A(p_input[5931]), .B(p_input[5899]), .Z(n18326) );
  XOR U17890 ( .A(n18327), .B(n18328), .Z(n18318) );
  AND U17891 ( .A(n18329), .B(n18330), .Z(n18328) );
  XOR U17892 ( .A(n18327), .B(n17494), .Z(n18330) );
  XNOR U17893 ( .A(p_input[5962]), .B(n18331), .Z(n17494) );
  AND U17894 ( .A(n315), .B(n18332), .Z(n18331) );
  XOR U17895 ( .A(p_input[5994]), .B(p_input[5962]), .Z(n18332) );
  XNOR U17896 ( .A(n17491), .B(n18327), .Z(n18329) );
  XOR U17897 ( .A(n18333), .B(n18334), .Z(n17491) );
  AND U17898 ( .A(n312), .B(n18335), .Z(n18334) );
  XOR U17899 ( .A(p_input[5930]), .B(p_input[5898]), .Z(n18335) );
  XOR U17900 ( .A(n18336), .B(n18337), .Z(n18327) );
  AND U17901 ( .A(n18338), .B(n18339), .Z(n18337) );
  XOR U17902 ( .A(n18336), .B(n17506), .Z(n18339) );
  XNOR U17903 ( .A(p_input[5961]), .B(n18340), .Z(n17506) );
  AND U17904 ( .A(n315), .B(n18341), .Z(n18340) );
  XOR U17905 ( .A(p_input[5993]), .B(p_input[5961]), .Z(n18341) );
  XNOR U17906 ( .A(n17503), .B(n18336), .Z(n18338) );
  XOR U17907 ( .A(n18342), .B(n18343), .Z(n17503) );
  AND U17908 ( .A(n312), .B(n18344), .Z(n18343) );
  XOR U17909 ( .A(p_input[5929]), .B(p_input[5897]), .Z(n18344) );
  XOR U17910 ( .A(n18345), .B(n18346), .Z(n18336) );
  AND U17911 ( .A(n18347), .B(n18348), .Z(n18346) );
  XOR U17912 ( .A(n18345), .B(n17518), .Z(n18348) );
  XNOR U17913 ( .A(p_input[5960]), .B(n18349), .Z(n17518) );
  AND U17914 ( .A(n315), .B(n18350), .Z(n18349) );
  XOR U17915 ( .A(p_input[5992]), .B(p_input[5960]), .Z(n18350) );
  XNOR U17916 ( .A(n17515), .B(n18345), .Z(n18347) );
  XOR U17917 ( .A(n18351), .B(n18352), .Z(n17515) );
  AND U17918 ( .A(n312), .B(n18353), .Z(n18352) );
  XOR U17919 ( .A(p_input[5928]), .B(p_input[5896]), .Z(n18353) );
  XOR U17920 ( .A(n18354), .B(n18355), .Z(n18345) );
  AND U17921 ( .A(n18356), .B(n18357), .Z(n18355) );
  XOR U17922 ( .A(n18354), .B(n17530), .Z(n18357) );
  XNOR U17923 ( .A(p_input[5959]), .B(n18358), .Z(n17530) );
  AND U17924 ( .A(n315), .B(n18359), .Z(n18358) );
  XOR U17925 ( .A(p_input[5991]), .B(p_input[5959]), .Z(n18359) );
  XNOR U17926 ( .A(n17527), .B(n18354), .Z(n18356) );
  XOR U17927 ( .A(n18360), .B(n18361), .Z(n17527) );
  AND U17928 ( .A(n312), .B(n18362), .Z(n18361) );
  XOR U17929 ( .A(p_input[5927]), .B(p_input[5895]), .Z(n18362) );
  XOR U17930 ( .A(n18363), .B(n18364), .Z(n18354) );
  AND U17931 ( .A(n18365), .B(n18366), .Z(n18364) );
  XOR U17932 ( .A(n18363), .B(n17542), .Z(n18366) );
  XNOR U17933 ( .A(p_input[5958]), .B(n18367), .Z(n17542) );
  AND U17934 ( .A(n315), .B(n18368), .Z(n18367) );
  XOR U17935 ( .A(p_input[5990]), .B(p_input[5958]), .Z(n18368) );
  XNOR U17936 ( .A(n17539), .B(n18363), .Z(n18365) );
  XOR U17937 ( .A(n18369), .B(n18370), .Z(n17539) );
  AND U17938 ( .A(n312), .B(n18371), .Z(n18370) );
  XOR U17939 ( .A(p_input[5926]), .B(p_input[5894]), .Z(n18371) );
  XOR U17940 ( .A(n18372), .B(n18373), .Z(n18363) );
  AND U17941 ( .A(n18374), .B(n18375), .Z(n18373) );
  XOR U17942 ( .A(n18372), .B(n17554), .Z(n18375) );
  XNOR U17943 ( .A(p_input[5957]), .B(n18376), .Z(n17554) );
  AND U17944 ( .A(n315), .B(n18377), .Z(n18376) );
  XOR U17945 ( .A(p_input[5989]), .B(p_input[5957]), .Z(n18377) );
  XNOR U17946 ( .A(n17551), .B(n18372), .Z(n18374) );
  XOR U17947 ( .A(n18378), .B(n18379), .Z(n17551) );
  AND U17948 ( .A(n312), .B(n18380), .Z(n18379) );
  XOR U17949 ( .A(p_input[5925]), .B(p_input[5893]), .Z(n18380) );
  XOR U17950 ( .A(n18381), .B(n18382), .Z(n18372) );
  AND U17951 ( .A(n18383), .B(n18384), .Z(n18382) );
  XOR U17952 ( .A(n18381), .B(n17566), .Z(n18384) );
  XNOR U17953 ( .A(p_input[5956]), .B(n18385), .Z(n17566) );
  AND U17954 ( .A(n315), .B(n18386), .Z(n18385) );
  XOR U17955 ( .A(p_input[5988]), .B(p_input[5956]), .Z(n18386) );
  XNOR U17956 ( .A(n17563), .B(n18381), .Z(n18383) );
  XOR U17957 ( .A(n18387), .B(n18388), .Z(n17563) );
  AND U17958 ( .A(n312), .B(n18389), .Z(n18388) );
  XOR U17959 ( .A(p_input[5924]), .B(p_input[5892]), .Z(n18389) );
  XOR U17960 ( .A(n18390), .B(n18391), .Z(n18381) );
  AND U17961 ( .A(n18392), .B(n18393), .Z(n18391) );
  XOR U17962 ( .A(n18390), .B(n17578), .Z(n18393) );
  XNOR U17963 ( .A(p_input[5955]), .B(n18394), .Z(n17578) );
  AND U17964 ( .A(n315), .B(n18395), .Z(n18394) );
  XOR U17965 ( .A(p_input[5987]), .B(p_input[5955]), .Z(n18395) );
  XNOR U17966 ( .A(n17575), .B(n18390), .Z(n18392) );
  XOR U17967 ( .A(n18396), .B(n18397), .Z(n17575) );
  AND U17968 ( .A(n312), .B(n18398), .Z(n18397) );
  XOR U17969 ( .A(p_input[5923]), .B(p_input[5891]), .Z(n18398) );
  XOR U17970 ( .A(n18399), .B(n18400), .Z(n18390) );
  AND U17971 ( .A(n18401), .B(n18402), .Z(n18400) );
  XOR U17972 ( .A(n18399), .B(n17590), .Z(n18402) );
  XNOR U17973 ( .A(p_input[5954]), .B(n18403), .Z(n17590) );
  AND U17974 ( .A(n315), .B(n18404), .Z(n18403) );
  XOR U17975 ( .A(p_input[5986]), .B(p_input[5954]), .Z(n18404) );
  XNOR U17976 ( .A(n17587), .B(n18399), .Z(n18401) );
  XOR U17977 ( .A(n18405), .B(n18406), .Z(n17587) );
  AND U17978 ( .A(n312), .B(n18407), .Z(n18406) );
  XOR U17979 ( .A(p_input[5922]), .B(p_input[5890]), .Z(n18407) );
  XOR U17980 ( .A(n18408), .B(n18409), .Z(n18399) );
  AND U17981 ( .A(n18410), .B(n18411), .Z(n18409) );
  XNOR U17982 ( .A(n18412), .B(n17603), .Z(n18411) );
  XNOR U17983 ( .A(p_input[5953]), .B(n18413), .Z(n17603) );
  AND U17984 ( .A(n315), .B(n18414), .Z(n18413) );
  XNOR U17985 ( .A(p_input[5985]), .B(n18415), .Z(n18414) );
  IV U17986 ( .A(p_input[5953]), .Z(n18415) );
  XNOR U17987 ( .A(n17600), .B(n18408), .Z(n18410) );
  XNOR U17988 ( .A(p_input[5889]), .B(n18416), .Z(n17600) );
  AND U17989 ( .A(n312), .B(n18417), .Z(n18416) );
  XOR U17990 ( .A(p_input[5921]), .B(p_input[5889]), .Z(n18417) );
  IV U17991 ( .A(n18412), .Z(n18408) );
  AND U17992 ( .A(n18138), .B(n18141), .Z(n18412) );
  XOR U17993 ( .A(p_input[5952]), .B(n18418), .Z(n18141) );
  AND U17994 ( .A(n315), .B(n18419), .Z(n18418) );
  XOR U17995 ( .A(p_input[5984]), .B(p_input[5952]), .Z(n18419) );
  XOR U17996 ( .A(n18420), .B(n18421), .Z(n315) );
  AND U17997 ( .A(n18422), .B(n18423), .Z(n18421) );
  XNOR U17998 ( .A(p_input[6015]), .B(n18420), .Z(n18423) );
  XOR U17999 ( .A(n18420), .B(p_input[5983]), .Z(n18422) );
  XOR U18000 ( .A(n18424), .B(n18425), .Z(n18420) );
  AND U18001 ( .A(n18426), .B(n18427), .Z(n18425) );
  XNOR U18002 ( .A(p_input[6014]), .B(n18424), .Z(n18427) );
  XOR U18003 ( .A(n18424), .B(p_input[5982]), .Z(n18426) );
  XOR U18004 ( .A(n18428), .B(n18429), .Z(n18424) );
  AND U18005 ( .A(n18430), .B(n18431), .Z(n18429) );
  XNOR U18006 ( .A(p_input[6013]), .B(n18428), .Z(n18431) );
  XOR U18007 ( .A(n18428), .B(p_input[5981]), .Z(n18430) );
  XOR U18008 ( .A(n18432), .B(n18433), .Z(n18428) );
  AND U18009 ( .A(n18434), .B(n18435), .Z(n18433) );
  XNOR U18010 ( .A(p_input[6012]), .B(n18432), .Z(n18435) );
  XOR U18011 ( .A(n18432), .B(p_input[5980]), .Z(n18434) );
  XOR U18012 ( .A(n18436), .B(n18437), .Z(n18432) );
  AND U18013 ( .A(n18438), .B(n18439), .Z(n18437) );
  XNOR U18014 ( .A(p_input[6011]), .B(n18436), .Z(n18439) );
  XOR U18015 ( .A(n18436), .B(p_input[5979]), .Z(n18438) );
  XOR U18016 ( .A(n18440), .B(n18441), .Z(n18436) );
  AND U18017 ( .A(n18442), .B(n18443), .Z(n18441) );
  XNOR U18018 ( .A(p_input[6010]), .B(n18440), .Z(n18443) );
  XOR U18019 ( .A(n18440), .B(p_input[5978]), .Z(n18442) );
  XOR U18020 ( .A(n18444), .B(n18445), .Z(n18440) );
  AND U18021 ( .A(n18446), .B(n18447), .Z(n18445) );
  XNOR U18022 ( .A(p_input[6009]), .B(n18444), .Z(n18447) );
  XOR U18023 ( .A(n18444), .B(p_input[5977]), .Z(n18446) );
  XOR U18024 ( .A(n18448), .B(n18449), .Z(n18444) );
  AND U18025 ( .A(n18450), .B(n18451), .Z(n18449) );
  XNOR U18026 ( .A(p_input[6008]), .B(n18448), .Z(n18451) );
  XOR U18027 ( .A(n18448), .B(p_input[5976]), .Z(n18450) );
  XOR U18028 ( .A(n18452), .B(n18453), .Z(n18448) );
  AND U18029 ( .A(n18454), .B(n18455), .Z(n18453) );
  XNOR U18030 ( .A(p_input[6007]), .B(n18452), .Z(n18455) );
  XOR U18031 ( .A(n18452), .B(p_input[5975]), .Z(n18454) );
  XOR U18032 ( .A(n18456), .B(n18457), .Z(n18452) );
  AND U18033 ( .A(n18458), .B(n18459), .Z(n18457) );
  XNOR U18034 ( .A(p_input[6006]), .B(n18456), .Z(n18459) );
  XOR U18035 ( .A(n18456), .B(p_input[5974]), .Z(n18458) );
  XOR U18036 ( .A(n18460), .B(n18461), .Z(n18456) );
  AND U18037 ( .A(n18462), .B(n18463), .Z(n18461) );
  XNOR U18038 ( .A(p_input[6005]), .B(n18460), .Z(n18463) );
  XOR U18039 ( .A(n18460), .B(p_input[5973]), .Z(n18462) );
  XOR U18040 ( .A(n18464), .B(n18465), .Z(n18460) );
  AND U18041 ( .A(n18466), .B(n18467), .Z(n18465) );
  XNOR U18042 ( .A(p_input[6004]), .B(n18464), .Z(n18467) );
  XOR U18043 ( .A(n18464), .B(p_input[5972]), .Z(n18466) );
  XOR U18044 ( .A(n18468), .B(n18469), .Z(n18464) );
  AND U18045 ( .A(n18470), .B(n18471), .Z(n18469) );
  XNOR U18046 ( .A(p_input[6003]), .B(n18468), .Z(n18471) );
  XOR U18047 ( .A(n18468), .B(p_input[5971]), .Z(n18470) );
  XOR U18048 ( .A(n18472), .B(n18473), .Z(n18468) );
  AND U18049 ( .A(n18474), .B(n18475), .Z(n18473) );
  XNOR U18050 ( .A(p_input[6002]), .B(n18472), .Z(n18475) );
  XOR U18051 ( .A(n18472), .B(p_input[5970]), .Z(n18474) );
  XOR U18052 ( .A(n18476), .B(n18477), .Z(n18472) );
  AND U18053 ( .A(n18478), .B(n18479), .Z(n18477) );
  XNOR U18054 ( .A(p_input[6001]), .B(n18476), .Z(n18479) );
  XOR U18055 ( .A(n18476), .B(p_input[5969]), .Z(n18478) );
  XOR U18056 ( .A(n18480), .B(n18481), .Z(n18476) );
  AND U18057 ( .A(n18482), .B(n18483), .Z(n18481) );
  XNOR U18058 ( .A(p_input[6000]), .B(n18480), .Z(n18483) );
  XOR U18059 ( .A(n18480), .B(p_input[5968]), .Z(n18482) );
  XOR U18060 ( .A(n18484), .B(n18485), .Z(n18480) );
  AND U18061 ( .A(n18486), .B(n18487), .Z(n18485) );
  XNOR U18062 ( .A(p_input[5999]), .B(n18484), .Z(n18487) );
  XOR U18063 ( .A(n18484), .B(p_input[5967]), .Z(n18486) );
  XOR U18064 ( .A(n18488), .B(n18489), .Z(n18484) );
  AND U18065 ( .A(n18490), .B(n18491), .Z(n18489) );
  XNOR U18066 ( .A(p_input[5998]), .B(n18488), .Z(n18491) );
  XOR U18067 ( .A(n18488), .B(p_input[5966]), .Z(n18490) );
  XOR U18068 ( .A(n18492), .B(n18493), .Z(n18488) );
  AND U18069 ( .A(n18494), .B(n18495), .Z(n18493) );
  XNOR U18070 ( .A(p_input[5997]), .B(n18492), .Z(n18495) );
  XOR U18071 ( .A(n18492), .B(p_input[5965]), .Z(n18494) );
  XOR U18072 ( .A(n18496), .B(n18497), .Z(n18492) );
  AND U18073 ( .A(n18498), .B(n18499), .Z(n18497) );
  XNOR U18074 ( .A(p_input[5996]), .B(n18496), .Z(n18499) );
  XOR U18075 ( .A(n18496), .B(p_input[5964]), .Z(n18498) );
  XOR U18076 ( .A(n18500), .B(n18501), .Z(n18496) );
  AND U18077 ( .A(n18502), .B(n18503), .Z(n18501) );
  XNOR U18078 ( .A(p_input[5995]), .B(n18500), .Z(n18503) );
  XOR U18079 ( .A(n18500), .B(p_input[5963]), .Z(n18502) );
  XOR U18080 ( .A(n18504), .B(n18505), .Z(n18500) );
  AND U18081 ( .A(n18506), .B(n18507), .Z(n18505) );
  XNOR U18082 ( .A(p_input[5994]), .B(n18504), .Z(n18507) );
  XOR U18083 ( .A(n18504), .B(p_input[5962]), .Z(n18506) );
  XOR U18084 ( .A(n18508), .B(n18509), .Z(n18504) );
  AND U18085 ( .A(n18510), .B(n18511), .Z(n18509) );
  XNOR U18086 ( .A(p_input[5993]), .B(n18508), .Z(n18511) );
  XOR U18087 ( .A(n18508), .B(p_input[5961]), .Z(n18510) );
  XOR U18088 ( .A(n18512), .B(n18513), .Z(n18508) );
  AND U18089 ( .A(n18514), .B(n18515), .Z(n18513) );
  XNOR U18090 ( .A(p_input[5992]), .B(n18512), .Z(n18515) );
  XOR U18091 ( .A(n18512), .B(p_input[5960]), .Z(n18514) );
  XOR U18092 ( .A(n18516), .B(n18517), .Z(n18512) );
  AND U18093 ( .A(n18518), .B(n18519), .Z(n18517) );
  XNOR U18094 ( .A(p_input[5991]), .B(n18516), .Z(n18519) );
  XOR U18095 ( .A(n18516), .B(p_input[5959]), .Z(n18518) );
  XOR U18096 ( .A(n18520), .B(n18521), .Z(n18516) );
  AND U18097 ( .A(n18522), .B(n18523), .Z(n18521) );
  XNOR U18098 ( .A(p_input[5990]), .B(n18520), .Z(n18523) );
  XOR U18099 ( .A(n18520), .B(p_input[5958]), .Z(n18522) );
  XOR U18100 ( .A(n18524), .B(n18525), .Z(n18520) );
  AND U18101 ( .A(n18526), .B(n18527), .Z(n18525) );
  XNOR U18102 ( .A(p_input[5989]), .B(n18524), .Z(n18527) );
  XOR U18103 ( .A(n18524), .B(p_input[5957]), .Z(n18526) );
  XOR U18104 ( .A(n18528), .B(n18529), .Z(n18524) );
  AND U18105 ( .A(n18530), .B(n18531), .Z(n18529) );
  XNOR U18106 ( .A(p_input[5988]), .B(n18528), .Z(n18531) );
  XOR U18107 ( .A(n18528), .B(p_input[5956]), .Z(n18530) );
  XOR U18108 ( .A(n18532), .B(n18533), .Z(n18528) );
  AND U18109 ( .A(n18534), .B(n18535), .Z(n18533) );
  XNOR U18110 ( .A(p_input[5987]), .B(n18532), .Z(n18535) );
  XOR U18111 ( .A(n18532), .B(p_input[5955]), .Z(n18534) );
  XOR U18112 ( .A(n18536), .B(n18537), .Z(n18532) );
  AND U18113 ( .A(n18538), .B(n18539), .Z(n18537) );
  XNOR U18114 ( .A(p_input[5986]), .B(n18536), .Z(n18539) );
  XOR U18115 ( .A(n18536), .B(p_input[5954]), .Z(n18538) );
  XNOR U18116 ( .A(n18540), .B(n18541), .Z(n18536) );
  AND U18117 ( .A(n18542), .B(n18543), .Z(n18541) );
  XOR U18118 ( .A(p_input[5985]), .B(n18540), .Z(n18543) );
  XNOR U18119 ( .A(p_input[5953]), .B(n18540), .Z(n18542) );
  AND U18120 ( .A(p_input[5984]), .B(n18544), .Z(n18540) );
  IV U18121 ( .A(p_input[5952]), .Z(n18544) );
  XNOR U18122 ( .A(p_input[5888]), .B(n18545), .Z(n18138) );
  AND U18123 ( .A(n312), .B(n18546), .Z(n18545) );
  XOR U18124 ( .A(p_input[5920]), .B(p_input[5888]), .Z(n18546) );
  XOR U18125 ( .A(n18547), .B(n18548), .Z(n312) );
  AND U18126 ( .A(n18549), .B(n18550), .Z(n18548) );
  XNOR U18127 ( .A(p_input[5951]), .B(n18547), .Z(n18550) );
  XOR U18128 ( .A(n18547), .B(p_input[5919]), .Z(n18549) );
  XOR U18129 ( .A(n18551), .B(n18552), .Z(n18547) );
  AND U18130 ( .A(n18553), .B(n18554), .Z(n18552) );
  XNOR U18131 ( .A(p_input[5950]), .B(n18551), .Z(n18554) );
  XNOR U18132 ( .A(n18551), .B(n18153), .Z(n18553) );
  IV U18133 ( .A(p_input[5918]), .Z(n18153) );
  XOR U18134 ( .A(n18555), .B(n18556), .Z(n18551) );
  AND U18135 ( .A(n18557), .B(n18558), .Z(n18556) );
  XNOR U18136 ( .A(p_input[5949]), .B(n18555), .Z(n18558) );
  XNOR U18137 ( .A(n18555), .B(n18162), .Z(n18557) );
  IV U18138 ( .A(p_input[5917]), .Z(n18162) );
  XOR U18139 ( .A(n18559), .B(n18560), .Z(n18555) );
  AND U18140 ( .A(n18561), .B(n18562), .Z(n18560) );
  XNOR U18141 ( .A(p_input[5948]), .B(n18559), .Z(n18562) );
  XNOR U18142 ( .A(n18559), .B(n18171), .Z(n18561) );
  IV U18143 ( .A(p_input[5916]), .Z(n18171) );
  XOR U18144 ( .A(n18563), .B(n18564), .Z(n18559) );
  AND U18145 ( .A(n18565), .B(n18566), .Z(n18564) );
  XNOR U18146 ( .A(p_input[5947]), .B(n18563), .Z(n18566) );
  XNOR U18147 ( .A(n18563), .B(n18180), .Z(n18565) );
  IV U18148 ( .A(p_input[5915]), .Z(n18180) );
  XOR U18149 ( .A(n18567), .B(n18568), .Z(n18563) );
  AND U18150 ( .A(n18569), .B(n18570), .Z(n18568) );
  XNOR U18151 ( .A(p_input[5946]), .B(n18567), .Z(n18570) );
  XNOR U18152 ( .A(n18567), .B(n18189), .Z(n18569) );
  IV U18153 ( .A(p_input[5914]), .Z(n18189) );
  XOR U18154 ( .A(n18571), .B(n18572), .Z(n18567) );
  AND U18155 ( .A(n18573), .B(n18574), .Z(n18572) );
  XNOR U18156 ( .A(p_input[5945]), .B(n18571), .Z(n18574) );
  XNOR U18157 ( .A(n18571), .B(n18198), .Z(n18573) );
  IV U18158 ( .A(p_input[5913]), .Z(n18198) );
  XOR U18159 ( .A(n18575), .B(n18576), .Z(n18571) );
  AND U18160 ( .A(n18577), .B(n18578), .Z(n18576) );
  XNOR U18161 ( .A(p_input[5944]), .B(n18575), .Z(n18578) );
  XNOR U18162 ( .A(n18575), .B(n18207), .Z(n18577) );
  IV U18163 ( .A(p_input[5912]), .Z(n18207) );
  XOR U18164 ( .A(n18579), .B(n18580), .Z(n18575) );
  AND U18165 ( .A(n18581), .B(n18582), .Z(n18580) );
  XNOR U18166 ( .A(p_input[5943]), .B(n18579), .Z(n18582) );
  XNOR U18167 ( .A(n18579), .B(n18216), .Z(n18581) );
  IV U18168 ( .A(p_input[5911]), .Z(n18216) );
  XOR U18169 ( .A(n18583), .B(n18584), .Z(n18579) );
  AND U18170 ( .A(n18585), .B(n18586), .Z(n18584) );
  XNOR U18171 ( .A(p_input[5942]), .B(n18583), .Z(n18586) );
  XNOR U18172 ( .A(n18583), .B(n18225), .Z(n18585) );
  IV U18173 ( .A(p_input[5910]), .Z(n18225) );
  XOR U18174 ( .A(n18587), .B(n18588), .Z(n18583) );
  AND U18175 ( .A(n18589), .B(n18590), .Z(n18588) );
  XNOR U18176 ( .A(p_input[5941]), .B(n18587), .Z(n18590) );
  XNOR U18177 ( .A(n18587), .B(n18234), .Z(n18589) );
  IV U18178 ( .A(p_input[5909]), .Z(n18234) );
  XOR U18179 ( .A(n18591), .B(n18592), .Z(n18587) );
  AND U18180 ( .A(n18593), .B(n18594), .Z(n18592) );
  XNOR U18181 ( .A(p_input[5940]), .B(n18591), .Z(n18594) );
  XNOR U18182 ( .A(n18591), .B(n18243), .Z(n18593) );
  IV U18183 ( .A(p_input[5908]), .Z(n18243) );
  XOR U18184 ( .A(n18595), .B(n18596), .Z(n18591) );
  AND U18185 ( .A(n18597), .B(n18598), .Z(n18596) );
  XNOR U18186 ( .A(p_input[5939]), .B(n18595), .Z(n18598) );
  XNOR U18187 ( .A(n18595), .B(n18252), .Z(n18597) );
  IV U18188 ( .A(p_input[5907]), .Z(n18252) );
  XOR U18189 ( .A(n18599), .B(n18600), .Z(n18595) );
  AND U18190 ( .A(n18601), .B(n18602), .Z(n18600) );
  XNOR U18191 ( .A(p_input[5938]), .B(n18599), .Z(n18602) );
  XNOR U18192 ( .A(n18599), .B(n18261), .Z(n18601) );
  IV U18193 ( .A(p_input[5906]), .Z(n18261) );
  XOR U18194 ( .A(n18603), .B(n18604), .Z(n18599) );
  AND U18195 ( .A(n18605), .B(n18606), .Z(n18604) );
  XNOR U18196 ( .A(p_input[5937]), .B(n18603), .Z(n18606) );
  XNOR U18197 ( .A(n18603), .B(n18270), .Z(n18605) );
  IV U18198 ( .A(p_input[5905]), .Z(n18270) );
  XOR U18199 ( .A(n18607), .B(n18608), .Z(n18603) );
  AND U18200 ( .A(n18609), .B(n18610), .Z(n18608) );
  XNOR U18201 ( .A(p_input[5936]), .B(n18607), .Z(n18610) );
  XNOR U18202 ( .A(n18607), .B(n18279), .Z(n18609) );
  IV U18203 ( .A(p_input[5904]), .Z(n18279) );
  XOR U18204 ( .A(n18611), .B(n18612), .Z(n18607) );
  AND U18205 ( .A(n18613), .B(n18614), .Z(n18612) );
  XNOR U18206 ( .A(p_input[5935]), .B(n18611), .Z(n18614) );
  XNOR U18207 ( .A(n18611), .B(n18288), .Z(n18613) );
  IV U18208 ( .A(p_input[5903]), .Z(n18288) );
  XOR U18209 ( .A(n18615), .B(n18616), .Z(n18611) );
  AND U18210 ( .A(n18617), .B(n18618), .Z(n18616) );
  XNOR U18211 ( .A(p_input[5934]), .B(n18615), .Z(n18618) );
  XNOR U18212 ( .A(n18615), .B(n18297), .Z(n18617) );
  IV U18213 ( .A(p_input[5902]), .Z(n18297) );
  XOR U18214 ( .A(n18619), .B(n18620), .Z(n18615) );
  AND U18215 ( .A(n18621), .B(n18622), .Z(n18620) );
  XNOR U18216 ( .A(p_input[5933]), .B(n18619), .Z(n18622) );
  XNOR U18217 ( .A(n18619), .B(n18306), .Z(n18621) );
  IV U18218 ( .A(p_input[5901]), .Z(n18306) );
  XOR U18219 ( .A(n18623), .B(n18624), .Z(n18619) );
  AND U18220 ( .A(n18625), .B(n18626), .Z(n18624) );
  XNOR U18221 ( .A(p_input[5932]), .B(n18623), .Z(n18626) );
  XNOR U18222 ( .A(n18623), .B(n18315), .Z(n18625) );
  IV U18223 ( .A(p_input[5900]), .Z(n18315) );
  XOR U18224 ( .A(n18627), .B(n18628), .Z(n18623) );
  AND U18225 ( .A(n18629), .B(n18630), .Z(n18628) );
  XNOR U18226 ( .A(p_input[5931]), .B(n18627), .Z(n18630) );
  XNOR U18227 ( .A(n18627), .B(n18324), .Z(n18629) );
  IV U18228 ( .A(p_input[5899]), .Z(n18324) );
  XOR U18229 ( .A(n18631), .B(n18632), .Z(n18627) );
  AND U18230 ( .A(n18633), .B(n18634), .Z(n18632) );
  XNOR U18231 ( .A(p_input[5930]), .B(n18631), .Z(n18634) );
  XNOR U18232 ( .A(n18631), .B(n18333), .Z(n18633) );
  IV U18233 ( .A(p_input[5898]), .Z(n18333) );
  XOR U18234 ( .A(n18635), .B(n18636), .Z(n18631) );
  AND U18235 ( .A(n18637), .B(n18638), .Z(n18636) );
  XNOR U18236 ( .A(p_input[5929]), .B(n18635), .Z(n18638) );
  XNOR U18237 ( .A(n18635), .B(n18342), .Z(n18637) );
  IV U18238 ( .A(p_input[5897]), .Z(n18342) );
  XOR U18239 ( .A(n18639), .B(n18640), .Z(n18635) );
  AND U18240 ( .A(n18641), .B(n18642), .Z(n18640) );
  XNOR U18241 ( .A(p_input[5928]), .B(n18639), .Z(n18642) );
  XNOR U18242 ( .A(n18639), .B(n18351), .Z(n18641) );
  IV U18243 ( .A(p_input[5896]), .Z(n18351) );
  XOR U18244 ( .A(n18643), .B(n18644), .Z(n18639) );
  AND U18245 ( .A(n18645), .B(n18646), .Z(n18644) );
  XNOR U18246 ( .A(p_input[5927]), .B(n18643), .Z(n18646) );
  XNOR U18247 ( .A(n18643), .B(n18360), .Z(n18645) );
  IV U18248 ( .A(p_input[5895]), .Z(n18360) );
  XOR U18249 ( .A(n18647), .B(n18648), .Z(n18643) );
  AND U18250 ( .A(n18649), .B(n18650), .Z(n18648) );
  XNOR U18251 ( .A(p_input[5926]), .B(n18647), .Z(n18650) );
  XNOR U18252 ( .A(n18647), .B(n18369), .Z(n18649) );
  IV U18253 ( .A(p_input[5894]), .Z(n18369) );
  XOR U18254 ( .A(n18651), .B(n18652), .Z(n18647) );
  AND U18255 ( .A(n18653), .B(n18654), .Z(n18652) );
  XNOR U18256 ( .A(p_input[5925]), .B(n18651), .Z(n18654) );
  XNOR U18257 ( .A(n18651), .B(n18378), .Z(n18653) );
  IV U18258 ( .A(p_input[5893]), .Z(n18378) );
  XOR U18259 ( .A(n18655), .B(n18656), .Z(n18651) );
  AND U18260 ( .A(n18657), .B(n18658), .Z(n18656) );
  XNOR U18261 ( .A(p_input[5924]), .B(n18655), .Z(n18658) );
  XNOR U18262 ( .A(n18655), .B(n18387), .Z(n18657) );
  IV U18263 ( .A(p_input[5892]), .Z(n18387) );
  XOR U18264 ( .A(n18659), .B(n18660), .Z(n18655) );
  AND U18265 ( .A(n18661), .B(n18662), .Z(n18660) );
  XNOR U18266 ( .A(p_input[5923]), .B(n18659), .Z(n18662) );
  XNOR U18267 ( .A(n18659), .B(n18396), .Z(n18661) );
  IV U18268 ( .A(p_input[5891]), .Z(n18396) );
  XOR U18269 ( .A(n18663), .B(n18664), .Z(n18659) );
  AND U18270 ( .A(n18665), .B(n18666), .Z(n18664) );
  XNOR U18271 ( .A(p_input[5922]), .B(n18663), .Z(n18666) );
  XNOR U18272 ( .A(n18663), .B(n18405), .Z(n18665) );
  IV U18273 ( .A(p_input[5890]), .Z(n18405) );
  XNOR U18274 ( .A(n18667), .B(n18668), .Z(n18663) );
  AND U18275 ( .A(n18669), .B(n18670), .Z(n18668) );
  XOR U18276 ( .A(p_input[5921]), .B(n18667), .Z(n18670) );
  XNOR U18277 ( .A(p_input[5889]), .B(n18667), .Z(n18669) );
  AND U18278 ( .A(p_input[5920]), .B(n18671), .Z(n18667) );
  IV U18279 ( .A(p_input[5888]), .Z(n18671) );
  XOR U18280 ( .A(n18672), .B(n18673), .Z(n16850) );
  AND U18281 ( .A(n841), .B(n18674), .Z(n18673) );
  XNOR U18282 ( .A(n18675), .B(n18672), .Z(n18674) );
  XOR U18283 ( .A(n18676), .B(n18677), .Z(n841) );
  AND U18284 ( .A(n18678), .B(n18679), .Z(n18677) );
  XOR U18285 ( .A(n18676), .B(n16865), .Z(n18679) );
  XNOR U18286 ( .A(n18680), .B(n18681), .Z(n16865) );
  AND U18287 ( .A(n18682), .B(n503), .Z(n18681) );
  AND U18288 ( .A(n18680), .B(n18683), .Z(n18682) );
  XNOR U18289 ( .A(n16862), .B(n18676), .Z(n18678) );
  XOR U18290 ( .A(n18684), .B(n18685), .Z(n16862) );
  AND U18291 ( .A(n18686), .B(n500), .Z(n18685) );
  NOR U18292 ( .A(n18684), .B(n18687), .Z(n18686) );
  XOR U18293 ( .A(n18688), .B(n18689), .Z(n18676) );
  AND U18294 ( .A(n18690), .B(n18691), .Z(n18689) );
  XOR U18295 ( .A(n18688), .B(n16877), .Z(n18691) );
  XOR U18296 ( .A(n18692), .B(n18693), .Z(n16877) );
  AND U18297 ( .A(n503), .B(n18694), .Z(n18693) );
  XOR U18298 ( .A(n18695), .B(n18692), .Z(n18694) );
  XNOR U18299 ( .A(n16874), .B(n18688), .Z(n18690) );
  XOR U18300 ( .A(n18696), .B(n18697), .Z(n16874) );
  AND U18301 ( .A(n500), .B(n18698), .Z(n18697) );
  XOR U18302 ( .A(n18699), .B(n18696), .Z(n18698) );
  XOR U18303 ( .A(n18700), .B(n18701), .Z(n18688) );
  AND U18304 ( .A(n18702), .B(n18703), .Z(n18701) );
  XOR U18305 ( .A(n18700), .B(n16889), .Z(n18703) );
  XOR U18306 ( .A(n18704), .B(n18705), .Z(n16889) );
  AND U18307 ( .A(n503), .B(n18706), .Z(n18705) );
  XOR U18308 ( .A(n18707), .B(n18704), .Z(n18706) );
  XNOR U18309 ( .A(n16886), .B(n18700), .Z(n18702) );
  XOR U18310 ( .A(n18708), .B(n18709), .Z(n16886) );
  AND U18311 ( .A(n500), .B(n18710), .Z(n18709) );
  XOR U18312 ( .A(n18711), .B(n18708), .Z(n18710) );
  XOR U18313 ( .A(n18712), .B(n18713), .Z(n18700) );
  AND U18314 ( .A(n18714), .B(n18715), .Z(n18713) );
  XOR U18315 ( .A(n18712), .B(n16901), .Z(n18715) );
  XOR U18316 ( .A(n18716), .B(n18717), .Z(n16901) );
  AND U18317 ( .A(n503), .B(n18718), .Z(n18717) );
  XOR U18318 ( .A(n18719), .B(n18716), .Z(n18718) );
  XNOR U18319 ( .A(n16898), .B(n18712), .Z(n18714) );
  XOR U18320 ( .A(n18720), .B(n18721), .Z(n16898) );
  AND U18321 ( .A(n500), .B(n18722), .Z(n18721) );
  XOR U18322 ( .A(n18723), .B(n18720), .Z(n18722) );
  XOR U18323 ( .A(n18724), .B(n18725), .Z(n18712) );
  AND U18324 ( .A(n18726), .B(n18727), .Z(n18725) );
  XOR U18325 ( .A(n18724), .B(n16913), .Z(n18727) );
  XOR U18326 ( .A(n18728), .B(n18729), .Z(n16913) );
  AND U18327 ( .A(n503), .B(n18730), .Z(n18729) );
  XOR U18328 ( .A(n18731), .B(n18728), .Z(n18730) );
  XNOR U18329 ( .A(n16910), .B(n18724), .Z(n18726) );
  XOR U18330 ( .A(n18732), .B(n18733), .Z(n16910) );
  AND U18331 ( .A(n500), .B(n18734), .Z(n18733) );
  XOR U18332 ( .A(n18735), .B(n18732), .Z(n18734) );
  XOR U18333 ( .A(n18736), .B(n18737), .Z(n18724) );
  AND U18334 ( .A(n18738), .B(n18739), .Z(n18737) );
  XOR U18335 ( .A(n18736), .B(n16925), .Z(n18739) );
  XOR U18336 ( .A(n18740), .B(n18741), .Z(n16925) );
  AND U18337 ( .A(n503), .B(n18742), .Z(n18741) );
  XOR U18338 ( .A(n18743), .B(n18740), .Z(n18742) );
  XNOR U18339 ( .A(n16922), .B(n18736), .Z(n18738) );
  XOR U18340 ( .A(n18744), .B(n18745), .Z(n16922) );
  AND U18341 ( .A(n500), .B(n18746), .Z(n18745) );
  XOR U18342 ( .A(n18747), .B(n18744), .Z(n18746) );
  XOR U18343 ( .A(n18748), .B(n18749), .Z(n18736) );
  AND U18344 ( .A(n18750), .B(n18751), .Z(n18749) );
  XOR U18345 ( .A(n18748), .B(n16937), .Z(n18751) );
  XOR U18346 ( .A(n18752), .B(n18753), .Z(n16937) );
  AND U18347 ( .A(n503), .B(n18754), .Z(n18753) );
  XOR U18348 ( .A(n18755), .B(n18752), .Z(n18754) );
  XNOR U18349 ( .A(n16934), .B(n18748), .Z(n18750) );
  XOR U18350 ( .A(n18756), .B(n18757), .Z(n16934) );
  AND U18351 ( .A(n500), .B(n18758), .Z(n18757) );
  XOR U18352 ( .A(n18759), .B(n18756), .Z(n18758) );
  XOR U18353 ( .A(n18760), .B(n18761), .Z(n18748) );
  AND U18354 ( .A(n18762), .B(n18763), .Z(n18761) );
  XOR U18355 ( .A(n18760), .B(n16949), .Z(n18763) );
  XOR U18356 ( .A(n18764), .B(n18765), .Z(n16949) );
  AND U18357 ( .A(n503), .B(n18766), .Z(n18765) );
  XOR U18358 ( .A(n18767), .B(n18764), .Z(n18766) );
  XNOR U18359 ( .A(n16946), .B(n18760), .Z(n18762) );
  XOR U18360 ( .A(n18768), .B(n18769), .Z(n16946) );
  AND U18361 ( .A(n500), .B(n18770), .Z(n18769) );
  XOR U18362 ( .A(n18771), .B(n18768), .Z(n18770) );
  XOR U18363 ( .A(n18772), .B(n18773), .Z(n18760) );
  AND U18364 ( .A(n18774), .B(n18775), .Z(n18773) );
  XOR U18365 ( .A(n18772), .B(n16961), .Z(n18775) );
  XOR U18366 ( .A(n18776), .B(n18777), .Z(n16961) );
  AND U18367 ( .A(n503), .B(n18778), .Z(n18777) );
  XOR U18368 ( .A(n18779), .B(n18776), .Z(n18778) );
  XNOR U18369 ( .A(n16958), .B(n18772), .Z(n18774) );
  XOR U18370 ( .A(n18780), .B(n18781), .Z(n16958) );
  AND U18371 ( .A(n500), .B(n18782), .Z(n18781) );
  XOR U18372 ( .A(n18783), .B(n18780), .Z(n18782) );
  XOR U18373 ( .A(n18784), .B(n18785), .Z(n18772) );
  AND U18374 ( .A(n18786), .B(n18787), .Z(n18785) );
  XOR U18375 ( .A(n18784), .B(n16973), .Z(n18787) );
  XOR U18376 ( .A(n18788), .B(n18789), .Z(n16973) );
  AND U18377 ( .A(n503), .B(n18790), .Z(n18789) );
  XOR U18378 ( .A(n18791), .B(n18788), .Z(n18790) );
  XNOR U18379 ( .A(n16970), .B(n18784), .Z(n18786) );
  XOR U18380 ( .A(n18792), .B(n18793), .Z(n16970) );
  AND U18381 ( .A(n500), .B(n18794), .Z(n18793) );
  XOR U18382 ( .A(n18795), .B(n18792), .Z(n18794) );
  XOR U18383 ( .A(n18796), .B(n18797), .Z(n18784) );
  AND U18384 ( .A(n18798), .B(n18799), .Z(n18797) );
  XOR U18385 ( .A(n18796), .B(n16985), .Z(n18799) );
  XOR U18386 ( .A(n18800), .B(n18801), .Z(n16985) );
  AND U18387 ( .A(n503), .B(n18802), .Z(n18801) );
  XOR U18388 ( .A(n18803), .B(n18800), .Z(n18802) );
  XNOR U18389 ( .A(n16982), .B(n18796), .Z(n18798) );
  XOR U18390 ( .A(n18804), .B(n18805), .Z(n16982) );
  AND U18391 ( .A(n500), .B(n18806), .Z(n18805) );
  XOR U18392 ( .A(n18807), .B(n18804), .Z(n18806) );
  XOR U18393 ( .A(n18808), .B(n18809), .Z(n18796) );
  AND U18394 ( .A(n18810), .B(n18811), .Z(n18809) );
  XOR U18395 ( .A(n18808), .B(n16997), .Z(n18811) );
  XOR U18396 ( .A(n18812), .B(n18813), .Z(n16997) );
  AND U18397 ( .A(n503), .B(n18814), .Z(n18813) );
  XOR U18398 ( .A(n18815), .B(n18812), .Z(n18814) );
  XNOR U18399 ( .A(n16994), .B(n18808), .Z(n18810) );
  XOR U18400 ( .A(n18816), .B(n18817), .Z(n16994) );
  AND U18401 ( .A(n500), .B(n18818), .Z(n18817) );
  XOR U18402 ( .A(n18819), .B(n18816), .Z(n18818) );
  XOR U18403 ( .A(n18820), .B(n18821), .Z(n18808) );
  AND U18404 ( .A(n18822), .B(n18823), .Z(n18821) );
  XOR U18405 ( .A(n18820), .B(n17009), .Z(n18823) );
  XOR U18406 ( .A(n18824), .B(n18825), .Z(n17009) );
  AND U18407 ( .A(n503), .B(n18826), .Z(n18825) );
  XOR U18408 ( .A(n18827), .B(n18824), .Z(n18826) );
  XNOR U18409 ( .A(n17006), .B(n18820), .Z(n18822) );
  XOR U18410 ( .A(n18828), .B(n18829), .Z(n17006) );
  AND U18411 ( .A(n500), .B(n18830), .Z(n18829) );
  XOR U18412 ( .A(n18831), .B(n18828), .Z(n18830) );
  XOR U18413 ( .A(n18832), .B(n18833), .Z(n18820) );
  AND U18414 ( .A(n18834), .B(n18835), .Z(n18833) );
  XOR U18415 ( .A(n18832), .B(n17021), .Z(n18835) );
  XOR U18416 ( .A(n18836), .B(n18837), .Z(n17021) );
  AND U18417 ( .A(n503), .B(n18838), .Z(n18837) );
  XOR U18418 ( .A(n18839), .B(n18836), .Z(n18838) );
  XNOR U18419 ( .A(n17018), .B(n18832), .Z(n18834) );
  XOR U18420 ( .A(n18840), .B(n18841), .Z(n17018) );
  AND U18421 ( .A(n500), .B(n18842), .Z(n18841) );
  XOR U18422 ( .A(n18843), .B(n18840), .Z(n18842) );
  XOR U18423 ( .A(n18844), .B(n18845), .Z(n18832) );
  AND U18424 ( .A(n18846), .B(n18847), .Z(n18845) );
  XOR U18425 ( .A(n18844), .B(n17033), .Z(n18847) );
  XOR U18426 ( .A(n18848), .B(n18849), .Z(n17033) );
  AND U18427 ( .A(n503), .B(n18850), .Z(n18849) );
  XOR U18428 ( .A(n18851), .B(n18848), .Z(n18850) );
  XNOR U18429 ( .A(n17030), .B(n18844), .Z(n18846) );
  XOR U18430 ( .A(n18852), .B(n18853), .Z(n17030) );
  AND U18431 ( .A(n500), .B(n18854), .Z(n18853) );
  XOR U18432 ( .A(n18855), .B(n18852), .Z(n18854) );
  XOR U18433 ( .A(n18856), .B(n18857), .Z(n18844) );
  AND U18434 ( .A(n18858), .B(n18859), .Z(n18857) );
  XOR U18435 ( .A(n18856), .B(n17045), .Z(n18859) );
  XOR U18436 ( .A(n18860), .B(n18861), .Z(n17045) );
  AND U18437 ( .A(n503), .B(n18862), .Z(n18861) );
  XOR U18438 ( .A(n18863), .B(n18860), .Z(n18862) );
  XNOR U18439 ( .A(n17042), .B(n18856), .Z(n18858) );
  XOR U18440 ( .A(n18864), .B(n18865), .Z(n17042) );
  AND U18441 ( .A(n500), .B(n18866), .Z(n18865) );
  XOR U18442 ( .A(n18867), .B(n18864), .Z(n18866) );
  XOR U18443 ( .A(n18868), .B(n18869), .Z(n18856) );
  AND U18444 ( .A(n18870), .B(n18871), .Z(n18869) );
  XOR U18445 ( .A(n18868), .B(n17057), .Z(n18871) );
  XOR U18446 ( .A(n18872), .B(n18873), .Z(n17057) );
  AND U18447 ( .A(n503), .B(n18874), .Z(n18873) );
  XOR U18448 ( .A(n18875), .B(n18872), .Z(n18874) );
  XNOR U18449 ( .A(n17054), .B(n18868), .Z(n18870) );
  XOR U18450 ( .A(n18876), .B(n18877), .Z(n17054) );
  AND U18451 ( .A(n500), .B(n18878), .Z(n18877) );
  XOR U18452 ( .A(n18879), .B(n18876), .Z(n18878) );
  XOR U18453 ( .A(n18880), .B(n18881), .Z(n18868) );
  AND U18454 ( .A(n18882), .B(n18883), .Z(n18881) );
  XOR U18455 ( .A(n18880), .B(n17069), .Z(n18883) );
  XOR U18456 ( .A(n18884), .B(n18885), .Z(n17069) );
  AND U18457 ( .A(n503), .B(n18886), .Z(n18885) );
  XOR U18458 ( .A(n18887), .B(n18884), .Z(n18886) );
  XNOR U18459 ( .A(n17066), .B(n18880), .Z(n18882) );
  XOR U18460 ( .A(n18888), .B(n18889), .Z(n17066) );
  AND U18461 ( .A(n500), .B(n18890), .Z(n18889) );
  XOR U18462 ( .A(n18891), .B(n18888), .Z(n18890) );
  XOR U18463 ( .A(n18892), .B(n18893), .Z(n18880) );
  AND U18464 ( .A(n18894), .B(n18895), .Z(n18893) );
  XOR U18465 ( .A(n18892), .B(n17081), .Z(n18895) );
  XOR U18466 ( .A(n18896), .B(n18897), .Z(n17081) );
  AND U18467 ( .A(n503), .B(n18898), .Z(n18897) );
  XOR U18468 ( .A(n18899), .B(n18896), .Z(n18898) );
  XNOR U18469 ( .A(n17078), .B(n18892), .Z(n18894) );
  XOR U18470 ( .A(n18900), .B(n18901), .Z(n17078) );
  AND U18471 ( .A(n500), .B(n18902), .Z(n18901) );
  XOR U18472 ( .A(n18903), .B(n18900), .Z(n18902) );
  XOR U18473 ( .A(n18904), .B(n18905), .Z(n18892) );
  AND U18474 ( .A(n18906), .B(n18907), .Z(n18905) );
  XOR U18475 ( .A(n18904), .B(n17093), .Z(n18907) );
  XOR U18476 ( .A(n18908), .B(n18909), .Z(n17093) );
  AND U18477 ( .A(n503), .B(n18910), .Z(n18909) );
  XOR U18478 ( .A(n18911), .B(n18908), .Z(n18910) );
  XNOR U18479 ( .A(n17090), .B(n18904), .Z(n18906) );
  XOR U18480 ( .A(n18912), .B(n18913), .Z(n17090) );
  AND U18481 ( .A(n500), .B(n18914), .Z(n18913) );
  XOR U18482 ( .A(n18915), .B(n18912), .Z(n18914) );
  XOR U18483 ( .A(n18916), .B(n18917), .Z(n18904) );
  AND U18484 ( .A(n18918), .B(n18919), .Z(n18917) );
  XOR U18485 ( .A(n18916), .B(n17105), .Z(n18919) );
  XOR U18486 ( .A(n18920), .B(n18921), .Z(n17105) );
  AND U18487 ( .A(n503), .B(n18922), .Z(n18921) );
  XOR U18488 ( .A(n18923), .B(n18920), .Z(n18922) );
  XNOR U18489 ( .A(n17102), .B(n18916), .Z(n18918) );
  XOR U18490 ( .A(n18924), .B(n18925), .Z(n17102) );
  AND U18491 ( .A(n500), .B(n18926), .Z(n18925) );
  XOR U18492 ( .A(n18927), .B(n18924), .Z(n18926) );
  XOR U18493 ( .A(n18928), .B(n18929), .Z(n18916) );
  AND U18494 ( .A(n18930), .B(n18931), .Z(n18929) );
  XOR U18495 ( .A(n18928), .B(n17117), .Z(n18931) );
  XOR U18496 ( .A(n18932), .B(n18933), .Z(n17117) );
  AND U18497 ( .A(n503), .B(n18934), .Z(n18933) );
  XOR U18498 ( .A(n18935), .B(n18932), .Z(n18934) );
  XNOR U18499 ( .A(n17114), .B(n18928), .Z(n18930) );
  XOR U18500 ( .A(n18936), .B(n18937), .Z(n17114) );
  AND U18501 ( .A(n500), .B(n18938), .Z(n18937) );
  XOR U18502 ( .A(n18939), .B(n18936), .Z(n18938) );
  XOR U18503 ( .A(n18940), .B(n18941), .Z(n18928) );
  AND U18504 ( .A(n18942), .B(n18943), .Z(n18941) );
  XOR U18505 ( .A(n18940), .B(n17129), .Z(n18943) );
  XOR U18506 ( .A(n18944), .B(n18945), .Z(n17129) );
  AND U18507 ( .A(n503), .B(n18946), .Z(n18945) );
  XOR U18508 ( .A(n18947), .B(n18944), .Z(n18946) );
  XNOR U18509 ( .A(n17126), .B(n18940), .Z(n18942) );
  XOR U18510 ( .A(n18948), .B(n18949), .Z(n17126) );
  AND U18511 ( .A(n500), .B(n18950), .Z(n18949) );
  XOR U18512 ( .A(n18951), .B(n18948), .Z(n18950) );
  XOR U18513 ( .A(n18952), .B(n18953), .Z(n18940) );
  AND U18514 ( .A(n18954), .B(n18955), .Z(n18953) );
  XOR U18515 ( .A(n18952), .B(n17141), .Z(n18955) );
  XOR U18516 ( .A(n18956), .B(n18957), .Z(n17141) );
  AND U18517 ( .A(n503), .B(n18958), .Z(n18957) );
  XOR U18518 ( .A(n18959), .B(n18956), .Z(n18958) );
  XNOR U18519 ( .A(n17138), .B(n18952), .Z(n18954) );
  XOR U18520 ( .A(n18960), .B(n18961), .Z(n17138) );
  AND U18521 ( .A(n500), .B(n18962), .Z(n18961) );
  XOR U18522 ( .A(n18963), .B(n18960), .Z(n18962) );
  XOR U18523 ( .A(n18964), .B(n18965), .Z(n18952) );
  AND U18524 ( .A(n18966), .B(n18967), .Z(n18965) );
  XOR U18525 ( .A(n18964), .B(n17153), .Z(n18967) );
  XOR U18526 ( .A(n18968), .B(n18969), .Z(n17153) );
  AND U18527 ( .A(n503), .B(n18970), .Z(n18969) );
  XOR U18528 ( .A(n18971), .B(n18968), .Z(n18970) );
  XNOR U18529 ( .A(n17150), .B(n18964), .Z(n18966) );
  XOR U18530 ( .A(n18972), .B(n18973), .Z(n17150) );
  AND U18531 ( .A(n500), .B(n18974), .Z(n18973) );
  XOR U18532 ( .A(n18975), .B(n18972), .Z(n18974) );
  XOR U18533 ( .A(n18976), .B(n18977), .Z(n18964) );
  AND U18534 ( .A(n18978), .B(n18979), .Z(n18977) );
  XOR U18535 ( .A(n18976), .B(n17165), .Z(n18979) );
  XOR U18536 ( .A(n18980), .B(n18981), .Z(n17165) );
  AND U18537 ( .A(n503), .B(n18982), .Z(n18981) );
  XOR U18538 ( .A(n18983), .B(n18980), .Z(n18982) );
  XNOR U18539 ( .A(n17162), .B(n18976), .Z(n18978) );
  XOR U18540 ( .A(n18984), .B(n18985), .Z(n17162) );
  AND U18541 ( .A(n500), .B(n18986), .Z(n18985) );
  XOR U18542 ( .A(n18987), .B(n18984), .Z(n18986) );
  XOR U18543 ( .A(n18988), .B(n18989), .Z(n18976) );
  AND U18544 ( .A(n18990), .B(n18991), .Z(n18989) );
  XOR U18545 ( .A(n18988), .B(n17177), .Z(n18991) );
  XOR U18546 ( .A(n18992), .B(n18993), .Z(n17177) );
  AND U18547 ( .A(n503), .B(n18994), .Z(n18993) );
  XOR U18548 ( .A(n18995), .B(n18992), .Z(n18994) );
  XNOR U18549 ( .A(n17174), .B(n18988), .Z(n18990) );
  XOR U18550 ( .A(n18996), .B(n18997), .Z(n17174) );
  AND U18551 ( .A(n500), .B(n18998), .Z(n18997) );
  XOR U18552 ( .A(n18999), .B(n18996), .Z(n18998) );
  XOR U18553 ( .A(n19000), .B(n19001), .Z(n18988) );
  AND U18554 ( .A(n19002), .B(n19003), .Z(n19001) );
  XOR U18555 ( .A(n19000), .B(n17189), .Z(n19003) );
  XOR U18556 ( .A(n19004), .B(n19005), .Z(n17189) );
  AND U18557 ( .A(n503), .B(n19006), .Z(n19005) );
  XOR U18558 ( .A(n19007), .B(n19004), .Z(n19006) );
  XNOR U18559 ( .A(n17186), .B(n19000), .Z(n19002) );
  XOR U18560 ( .A(n19008), .B(n19009), .Z(n17186) );
  AND U18561 ( .A(n500), .B(n19010), .Z(n19009) );
  XOR U18562 ( .A(n19011), .B(n19008), .Z(n19010) );
  XOR U18563 ( .A(n19012), .B(n19013), .Z(n19000) );
  AND U18564 ( .A(n19014), .B(n19015), .Z(n19013) );
  XOR U18565 ( .A(n19012), .B(n17201), .Z(n19015) );
  XOR U18566 ( .A(n19016), .B(n19017), .Z(n17201) );
  AND U18567 ( .A(n503), .B(n19018), .Z(n19017) );
  XOR U18568 ( .A(n19019), .B(n19016), .Z(n19018) );
  XNOR U18569 ( .A(n17198), .B(n19012), .Z(n19014) );
  XOR U18570 ( .A(n19020), .B(n19021), .Z(n17198) );
  AND U18571 ( .A(n500), .B(n19022), .Z(n19021) );
  XOR U18572 ( .A(n19023), .B(n19020), .Z(n19022) );
  XOR U18573 ( .A(n19024), .B(n19025), .Z(n19012) );
  AND U18574 ( .A(n19026), .B(n19027), .Z(n19025) );
  XOR U18575 ( .A(n19024), .B(n17213), .Z(n19027) );
  XOR U18576 ( .A(n19028), .B(n19029), .Z(n17213) );
  AND U18577 ( .A(n503), .B(n19030), .Z(n19029) );
  XOR U18578 ( .A(n19031), .B(n19028), .Z(n19030) );
  XNOR U18579 ( .A(n17210), .B(n19024), .Z(n19026) );
  XOR U18580 ( .A(n19032), .B(n19033), .Z(n17210) );
  AND U18581 ( .A(n500), .B(n19034), .Z(n19033) );
  XOR U18582 ( .A(n19035), .B(n19032), .Z(n19034) );
  XOR U18583 ( .A(n19036), .B(n19037), .Z(n19024) );
  AND U18584 ( .A(n19038), .B(n19039), .Z(n19037) );
  XNOR U18585 ( .A(n19040), .B(n17226), .Z(n19039) );
  XOR U18586 ( .A(n19041), .B(n19042), .Z(n17226) );
  AND U18587 ( .A(n503), .B(n19043), .Z(n19042) );
  XOR U18588 ( .A(n19041), .B(n19044), .Z(n19043) );
  XNOR U18589 ( .A(n17223), .B(n19036), .Z(n19038) );
  XOR U18590 ( .A(n19045), .B(n19046), .Z(n17223) );
  AND U18591 ( .A(n500), .B(n19047), .Z(n19046) );
  XOR U18592 ( .A(n19045), .B(n19048), .Z(n19047) );
  IV U18593 ( .A(n19040), .Z(n19036) );
  AND U18594 ( .A(n18672), .B(n18675), .Z(n19040) );
  XNOR U18595 ( .A(n19049), .B(n19050), .Z(n18675) );
  AND U18596 ( .A(n503), .B(n19051), .Z(n19050) );
  XNOR U18597 ( .A(n19052), .B(n19049), .Z(n19051) );
  XOR U18598 ( .A(n19053), .B(n19054), .Z(n503) );
  AND U18599 ( .A(n19055), .B(n19056), .Z(n19054) );
  XOR U18600 ( .A(n18683), .B(n19053), .Z(n19056) );
  IV U18601 ( .A(n19057), .Z(n18683) );
  AND U18602 ( .A(p_input[5887]), .B(p_input[5855]), .Z(n19057) );
  XOR U18603 ( .A(n19053), .B(n18680), .Z(n19055) );
  AND U18604 ( .A(p_input[5791]), .B(p_input[5823]), .Z(n18680) );
  XOR U18605 ( .A(n19058), .B(n19059), .Z(n19053) );
  AND U18606 ( .A(n19060), .B(n19061), .Z(n19059) );
  XOR U18607 ( .A(n19058), .B(n18695), .Z(n19061) );
  XNOR U18608 ( .A(p_input[5854]), .B(n19062), .Z(n18695) );
  AND U18609 ( .A(n323), .B(n19063), .Z(n19062) );
  XOR U18610 ( .A(p_input[5886]), .B(p_input[5854]), .Z(n19063) );
  XNOR U18611 ( .A(n18692), .B(n19058), .Z(n19060) );
  XOR U18612 ( .A(n19064), .B(n19065), .Z(n18692) );
  AND U18613 ( .A(n321), .B(n19066), .Z(n19065) );
  XOR U18614 ( .A(p_input[5822]), .B(p_input[5790]), .Z(n19066) );
  XOR U18615 ( .A(n19067), .B(n19068), .Z(n19058) );
  AND U18616 ( .A(n19069), .B(n19070), .Z(n19068) );
  XOR U18617 ( .A(n19067), .B(n18707), .Z(n19070) );
  XNOR U18618 ( .A(p_input[5853]), .B(n19071), .Z(n18707) );
  AND U18619 ( .A(n323), .B(n19072), .Z(n19071) );
  XOR U18620 ( .A(p_input[5885]), .B(p_input[5853]), .Z(n19072) );
  XNOR U18621 ( .A(n18704), .B(n19067), .Z(n19069) );
  XOR U18622 ( .A(n19073), .B(n19074), .Z(n18704) );
  AND U18623 ( .A(n321), .B(n19075), .Z(n19074) );
  XOR U18624 ( .A(p_input[5821]), .B(p_input[5789]), .Z(n19075) );
  XOR U18625 ( .A(n19076), .B(n19077), .Z(n19067) );
  AND U18626 ( .A(n19078), .B(n19079), .Z(n19077) );
  XOR U18627 ( .A(n19076), .B(n18719), .Z(n19079) );
  XNOR U18628 ( .A(p_input[5852]), .B(n19080), .Z(n18719) );
  AND U18629 ( .A(n323), .B(n19081), .Z(n19080) );
  XOR U18630 ( .A(p_input[5884]), .B(p_input[5852]), .Z(n19081) );
  XNOR U18631 ( .A(n18716), .B(n19076), .Z(n19078) );
  XOR U18632 ( .A(n19082), .B(n19083), .Z(n18716) );
  AND U18633 ( .A(n321), .B(n19084), .Z(n19083) );
  XOR U18634 ( .A(p_input[5820]), .B(p_input[5788]), .Z(n19084) );
  XOR U18635 ( .A(n19085), .B(n19086), .Z(n19076) );
  AND U18636 ( .A(n19087), .B(n19088), .Z(n19086) );
  XOR U18637 ( .A(n19085), .B(n18731), .Z(n19088) );
  XNOR U18638 ( .A(p_input[5851]), .B(n19089), .Z(n18731) );
  AND U18639 ( .A(n323), .B(n19090), .Z(n19089) );
  XOR U18640 ( .A(p_input[5883]), .B(p_input[5851]), .Z(n19090) );
  XNOR U18641 ( .A(n18728), .B(n19085), .Z(n19087) );
  XOR U18642 ( .A(n19091), .B(n19092), .Z(n18728) );
  AND U18643 ( .A(n321), .B(n19093), .Z(n19092) );
  XOR U18644 ( .A(p_input[5819]), .B(p_input[5787]), .Z(n19093) );
  XOR U18645 ( .A(n19094), .B(n19095), .Z(n19085) );
  AND U18646 ( .A(n19096), .B(n19097), .Z(n19095) );
  XOR U18647 ( .A(n19094), .B(n18743), .Z(n19097) );
  XNOR U18648 ( .A(p_input[5850]), .B(n19098), .Z(n18743) );
  AND U18649 ( .A(n323), .B(n19099), .Z(n19098) );
  XOR U18650 ( .A(p_input[5882]), .B(p_input[5850]), .Z(n19099) );
  XNOR U18651 ( .A(n18740), .B(n19094), .Z(n19096) );
  XOR U18652 ( .A(n19100), .B(n19101), .Z(n18740) );
  AND U18653 ( .A(n321), .B(n19102), .Z(n19101) );
  XOR U18654 ( .A(p_input[5818]), .B(p_input[5786]), .Z(n19102) );
  XOR U18655 ( .A(n19103), .B(n19104), .Z(n19094) );
  AND U18656 ( .A(n19105), .B(n19106), .Z(n19104) );
  XOR U18657 ( .A(n19103), .B(n18755), .Z(n19106) );
  XNOR U18658 ( .A(p_input[5849]), .B(n19107), .Z(n18755) );
  AND U18659 ( .A(n323), .B(n19108), .Z(n19107) );
  XOR U18660 ( .A(p_input[5881]), .B(p_input[5849]), .Z(n19108) );
  XNOR U18661 ( .A(n18752), .B(n19103), .Z(n19105) );
  XOR U18662 ( .A(n19109), .B(n19110), .Z(n18752) );
  AND U18663 ( .A(n321), .B(n19111), .Z(n19110) );
  XOR U18664 ( .A(p_input[5817]), .B(p_input[5785]), .Z(n19111) );
  XOR U18665 ( .A(n19112), .B(n19113), .Z(n19103) );
  AND U18666 ( .A(n19114), .B(n19115), .Z(n19113) );
  XOR U18667 ( .A(n19112), .B(n18767), .Z(n19115) );
  XNOR U18668 ( .A(p_input[5848]), .B(n19116), .Z(n18767) );
  AND U18669 ( .A(n323), .B(n19117), .Z(n19116) );
  XOR U18670 ( .A(p_input[5880]), .B(p_input[5848]), .Z(n19117) );
  XNOR U18671 ( .A(n18764), .B(n19112), .Z(n19114) );
  XOR U18672 ( .A(n19118), .B(n19119), .Z(n18764) );
  AND U18673 ( .A(n321), .B(n19120), .Z(n19119) );
  XOR U18674 ( .A(p_input[5816]), .B(p_input[5784]), .Z(n19120) );
  XOR U18675 ( .A(n19121), .B(n19122), .Z(n19112) );
  AND U18676 ( .A(n19123), .B(n19124), .Z(n19122) );
  XOR U18677 ( .A(n19121), .B(n18779), .Z(n19124) );
  XNOR U18678 ( .A(p_input[5847]), .B(n19125), .Z(n18779) );
  AND U18679 ( .A(n323), .B(n19126), .Z(n19125) );
  XOR U18680 ( .A(p_input[5879]), .B(p_input[5847]), .Z(n19126) );
  XNOR U18681 ( .A(n18776), .B(n19121), .Z(n19123) );
  XOR U18682 ( .A(n19127), .B(n19128), .Z(n18776) );
  AND U18683 ( .A(n321), .B(n19129), .Z(n19128) );
  XOR U18684 ( .A(p_input[5815]), .B(p_input[5783]), .Z(n19129) );
  XOR U18685 ( .A(n19130), .B(n19131), .Z(n19121) );
  AND U18686 ( .A(n19132), .B(n19133), .Z(n19131) );
  XOR U18687 ( .A(n19130), .B(n18791), .Z(n19133) );
  XNOR U18688 ( .A(p_input[5846]), .B(n19134), .Z(n18791) );
  AND U18689 ( .A(n323), .B(n19135), .Z(n19134) );
  XOR U18690 ( .A(p_input[5878]), .B(p_input[5846]), .Z(n19135) );
  XNOR U18691 ( .A(n18788), .B(n19130), .Z(n19132) );
  XOR U18692 ( .A(n19136), .B(n19137), .Z(n18788) );
  AND U18693 ( .A(n321), .B(n19138), .Z(n19137) );
  XOR U18694 ( .A(p_input[5814]), .B(p_input[5782]), .Z(n19138) );
  XOR U18695 ( .A(n19139), .B(n19140), .Z(n19130) );
  AND U18696 ( .A(n19141), .B(n19142), .Z(n19140) );
  XOR U18697 ( .A(n19139), .B(n18803), .Z(n19142) );
  XNOR U18698 ( .A(p_input[5845]), .B(n19143), .Z(n18803) );
  AND U18699 ( .A(n323), .B(n19144), .Z(n19143) );
  XOR U18700 ( .A(p_input[5877]), .B(p_input[5845]), .Z(n19144) );
  XNOR U18701 ( .A(n18800), .B(n19139), .Z(n19141) );
  XOR U18702 ( .A(n19145), .B(n19146), .Z(n18800) );
  AND U18703 ( .A(n321), .B(n19147), .Z(n19146) );
  XOR U18704 ( .A(p_input[5813]), .B(p_input[5781]), .Z(n19147) );
  XOR U18705 ( .A(n19148), .B(n19149), .Z(n19139) );
  AND U18706 ( .A(n19150), .B(n19151), .Z(n19149) );
  XOR U18707 ( .A(n19148), .B(n18815), .Z(n19151) );
  XNOR U18708 ( .A(p_input[5844]), .B(n19152), .Z(n18815) );
  AND U18709 ( .A(n323), .B(n19153), .Z(n19152) );
  XOR U18710 ( .A(p_input[5876]), .B(p_input[5844]), .Z(n19153) );
  XNOR U18711 ( .A(n18812), .B(n19148), .Z(n19150) );
  XOR U18712 ( .A(n19154), .B(n19155), .Z(n18812) );
  AND U18713 ( .A(n321), .B(n19156), .Z(n19155) );
  XOR U18714 ( .A(p_input[5812]), .B(p_input[5780]), .Z(n19156) );
  XOR U18715 ( .A(n19157), .B(n19158), .Z(n19148) );
  AND U18716 ( .A(n19159), .B(n19160), .Z(n19158) );
  XOR U18717 ( .A(n19157), .B(n18827), .Z(n19160) );
  XNOR U18718 ( .A(p_input[5843]), .B(n19161), .Z(n18827) );
  AND U18719 ( .A(n323), .B(n19162), .Z(n19161) );
  XOR U18720 ( .A(p_input[5875]), .B(p_input[5843]), .Z(n19162) );
  XNOR U18721 ( .A(n18824), .B(n19157), .Z(n19159) );
  XOR U18722 ( .A(n19163), .B(n19164), .Z(n18824) );
  AND U18723 ( .A(n321), .B(n19165), .Z(n19164) );
  XOR U18724 ( .A(p_input[5811]), .B(p_input[5779]), .Z(n19165) );
  XOR U18725 ( .A(n19166), .B(n19167), .Z(n19157) );
  AND U18726 ( .A(n19168), .B(n19169), .Z(n19167) );
  XOR U18727 ( .A(n19166), .B(n18839), .Z(n19169) );
  XNOR U18728 ( .A(p_input[5842]), .B(n19170), .Z(n18839) );
  AND U18729 ( .A(n323), .B(n19171), .Z(n19170) );
  XOR U18730 ( .A(p_input[5874]), .B(p_input[5842]), .Z(n19171) );
  XNOR U18731 ( .A(n18836), .B(n19166), .Z(n19168) );
  XOR U18732 ( .A(n19172), .B(n19173), .Z(n18836) );
  AND U18733 ( .A(n321), .B(n19174), .Z(n19173) );
  XOR U18734 ( .A(p_input[5810]), .B(p_input[5778]), .Z(n19174) );
  XOR U18735 ( .A(n19175), .B(n19176), .Z(n19166) );
  AND U18736 ( .A(n19177), .B(n19178), .Z(n19176) );
  XOR U18737 ( .A(n19175), .B(n18851), .Z(n19178) );
  XNOR U18738 ( .A(p_input[5841]), .B(n19179), .Z(n18851) );
  AND U18739 ( .A(n323), .B(n19180), .Z(n19179) );
  XOR U18740 ( .A(p_input[5873]), .B(p_input[5841]), .Z(n19180) );
  XNOR U18741 ( .A(n18848), .B(n19175), .Z(n19177) );
  XOR U18742 ( .A(n19181), .B(n19182), .Z(n18848) );
  AND U18743 ( .A(n321), .B(n19183), .Z(n19182) );
  XOR U18744 ( .A(p_input[5809]), .B(p_input[5777]), .Z(n19183) );
  XOR U18745 ( .A(n19184), .B(n19185), .Z(n19175) );
  AND U18746 ( .A(n19186), .B(n19187), .Z(n19185) );
  XOR U18747 ( .A(n19184), .B(n18863), .Z(n19187) );
  XNOR U18748 ( .A(p_input[5840]), .B(n19188), .Z(n18863) );
  AND U18749 ( .A(n323), .B(n19189), .Z(n19188) );
  XOR U18750 ( .A(p_input[5872]), .B(p_input[5840]), .Z(n19189) );
  XNOR U18751 ( .A(n18860), .B(n19184), .Z(n19186) );
  XOR U18752 ( .A(n19190), .B(n19191), .Z(n18860) );
  AND U18753 ( .A(n321), .B(n19192), .Z(n19191) );
  XOR U18754 ( .A(p_input[5808]), .B(p_input[5776]), .Z(n19192) );
  XOR U18755 ( .A(n19193), .B(n19194), .Z(n19184) );
  AND U18756 ( .A(n19195), .B(n19196), .Z(n19194) );
  XOR U18757 ( .A(n19193), .B(n18875), .Z(n19196) );
  XNOR U18758 ( .A(p_input[5839]), .B(n19197), .Z(n18875) );
  AND U18759 ( .A(n323), .B(n19198), .Z(n19197) );
  XOR U18760 ( .A(p_input[5871]), .B(p_input[5839]), .Z(n19198) );
  XNOR U18761 ( .A(n18872), .B(n19193), .Z(n19195) );
  XOR U18762 ( .A(n19199), .B(n19200), .Z(n18872) );
  AND U18763 ( .A(n321), .B(n19201), .Z(n19200) );
  XOR U18764 ( .A(p_input[5807]), .B(p_input[5775]), .Z(n19201) );
  XOR U18765 ( .A(n19202), .B(n19203), .Z(n19193) );
  AND U18766 ( .A(n19204), .B(n19205), .Z(n19203) );
  XOR U18767 ( .A(n19202), .B(n18887), .Z(n19205) );
  XNOR U18768 ( .A(p_input[5838]), .B(n19206), .Z(n18887) );
  AND U18769 ( .A(n323), .B(n19207), .Z(n19206) );
  XOR U18770 ( .A(p_input[5870]), .B(p_input[5838]), .Z(n19207) );
  XNOR U18771 ( .A(n18884), .B(n19202), .Z(n19204) );
  XOR U18772 ( .A(n19208), .B(n19209), .Z(n18884) );
  AND U18773 ( .A(n321), .B(n19210), .Z(n19209) );
  XOR U18774 ( .A(p_input[5806]), .B(p_input[5774]), .Z(n19210) );
  XOR U18775 ( .A(n19211), .B(n19212), .Z(n19202) );
  AND U18776 ( .A(n19213), .B(n19214), .Z(n19212) );
  XOR U18777 ( .A(n19211), .B(n18899), .Z(n19214) );
  XNOR U18778 ( .A(p_input[5837]), .B(n19215), .Z(n18899) );
  AND U18779 ( .A(n323), .B(n19216), .Z(n19215) );
  XOR U18780 ( .A(p_input[5869]), .B(p_input[5837]), .Z(n19216) );
  XNOR U18781 ( .A(n18896), .B(n19211), .Z(n19213) );
  XOR U18782 ( .A(n19217), .B(n19218), .Z(n18896) );
  AND U18783 ( .A(n321), .B(n19219), .Z(n19218) );
  XOR U18784 ( .A(p_input[5805]), .B(p_input[5773]), .Z(n19219) );
  XOR U18785 ( .A(n19220), .B(n19221), .Z(n19211) );
  AND U18786 ( .A(n19222), .B(n19223), .Z(n19221) );
  XOR U18787 ( .A(n19220), .B(n18911), .Z(n19223) );
  XNOR U18788 ( .A(p_input[5836]), .B(n19224), .Z(n18911) );
  AND U18789 ( .A(n323), .B(n19225), .Z(n19224) );
  XOR U18790 ( .A(p_input[5868]), .B(p_input[5836]), .Z(n19225) );
  XNOR U18791 ( .A(n18908), .B(n19220), .Z(n19222) );
  XOR U18792 ( .A(n19226), .B(n19227), .Z(n18908) );
  AND U18793 ( .A(n321), .B(n19228), .Z(n19227) );
  XOR U18794 ( .A(p_input[5804]), .B(p_input[5772]), .Z(n19228) );
  XOR U18795 ( .A(n19229), .B(n19230), .Z(n19220) );
  AND U18796 ( .A(n19231), .B(n19232), .Z(n19230) );
  XOR U18797 ( .A(n19229), .B(n18923), .Z(n19232) );
  XNOR U18798 ( .A(p_input[5835]), .B(n19233), .Z(n18923) );
  AND U18799 ( .A(n323), .B(n19234), .Z(n19233) );
  XOR U18800 ( .A(p_input[5867]), .B(p_input[5835]), .Z(n19234) );
  XNOR U18801 ( .A(n18920), .B(n19229), .Z(n19231) );
  XOR U18802 ( .A(n19235), .B(n19236), .Z(n18920) );
  AND U18803 ( .A(n321), .B(n19237), .Z(n19236) );
  XOR U18804 ( .A(p_input[5803]), .B(p_input[5771]), .Z(n19237) );
  XOR U18805 ( .A(n19238), .B(n19239), .Z(n19229) );
  AND U18806 ( .A(n19240), .B(n19241), .Z(n19239) );
  XOR U18807 ( .A(n19238), .B(n18935), .Z(n19241) );
  XNOR U18808 ( .A(p_input[5834]), .B(n19242), .Z(n18935) );
  AND U18809 ( .A(n323), .B(n19243), .Z(n19242) );
  XOR U18810 ( .A(p_input[5866]), .B(p_input[5834]), .Z(n19243) );
  XNOR U18811 ( .A(n18932), .B(n19238), .Z(n19240) );
  XOR U18812 ( .A(n19244), .B(n19245), .Z(n18932) );
  AND U18813 ( .A(n321), .B(n19246), .Z(n19245) );
  XOR U18814 ( .A(p_input[5802]), .B(p_input[5770]), .Z(n19246) );
  XOR U18815 ( .A(n19247), .B(n19248), .Z(n19238) );
  AND U18816 ( .A(n19249), .B(n19250), .Z(n19248) );
  XOR U18817 ( .A(n19247), .B(n18947), .Z(n19250) );
  XNOR U18818 ( .A(p_input[5833]), .B(n19251), .Z(n18947) );
  AND U18819 ( .A(n323), .B(n19252), .Z(n19251) );
  XOR U18820 ( .A(p_input[5865]), .B(p_input[5833]), .Z(n19252) );
  XNOR U18821 ( .A(n18944), .B(n19247), .Z(n19249) );
  XOR U18822 ( .A(n19253), .B(n19254), .Z(n18944) );
  AND U18823 ( .A(n321), .B(n19255), .Z(n19254) );
  XOR U18824 ( .A(p_input[5801]), .B(p_input[5769]), .Z(n19255) );
  XOR U18825 ( .A(n19256), .B(n19257), .Z(n19247) );
  AND U18826 ( .A(n19258), .B(n19259), .Z(n19257) );
  XOR U18827 ( .A(n19256), .B(n18959), .Z(n19259) );
  XNOR U18828 ( .A(p_input[5832]), .B(n19260), .Z(n18959) );
  AND U18829 ( .A(n323), .B(n19261), .Z(n19260) );
  XOR U18830 ( .A(p_input[5864]), .B(p_input[5832]), .Z(n19261) );
  XNOR U18831 ( .A(n18956), .B(n19256), .Z(n19258) );
  XOR U18832 ( .A(n19262), .B(n19263), .Z(n18956) );
  AND U18833 ( .A(n321), .B(n19264), .Z(n19263) );
  XOR U18834 ( .A(p_input[5800]), .B(p_input[5768]), .Z(n19264) );
  XOR U18835 ( .A(n19265), .B(n19266), .Z(n19256) );
  AND U18836 ( .A(n19267), .B(n19268), .Z(n19266) );
  XOR U18837 ( .A(n19265), .B(n18971), .Z(n19268) );
  XNOR U18838 ( .A(p_input[5831]), .B(n19269), .Z(n18971) );
  AND U18839 ( .A(n323), .B(n19270), .Z(n19269) );
  XOR U18840 ( .A(p_input[5863]), .B(p_input[5831]), .Z(n19270) );
  XNOR U18841 ( .A(n18968), .B(n19265), .Z(n19267) );
  XOR U18842 ( .A(n19271), .B(n19272), .Z(n18968) );
  AND U18843 ( .A(n321), .B(n19273), .Z(n19272) );
  XOR U18844 ( .A(p_input[5799]), .B(p_input[5767]), .Z(n19273) );
  XOR U18845 ( .A(n19274), .B(n19275), .Z(n19265) );
  AND U18846 ( .A(n19276), .B(n19277), .Z(n19275) );
  XOR U18847 ( .A(n19274), .B(n18983), .Z(n19277) );
  XNOR U18848 ( .A(p_input[5830]), .B(n19278), .Z(n18983) );
  AND U18849 ( .A(n323), .B(n19279), .Z(n19278) );
  XOR U18850 ( .A(p_input[5862]), .B(p_input[5830]), .Z(n19279) );
  XNOR U18851 ( .A(n18980), .B(n19274), .Z(n19276) );
  XOR U18852 ( .A(n19280), .B(n19281), .Z(n18980) );
  AND U18853 ( .A(n321), .B(n19282), .Z(n19281) );
  XOR U18854 ( .A(p_input[5798]), .B(p_input[5766]), .Z(n19282) );
  XOR U18855 ( .A(n19283), .B(n19284), .Z(n19274) );
  AND U18856 ( .A(n19285), .B(n19286), .Z(n19284) );
  XOR U18857 ( .A(n19283), .B(n18995), .Z(n19286) );
  XNOR U18858 ( .A(p_input[5829]), .B(n19287), .Z(n18995) );
  AND U18859 ( .A(n323), .B(n19288), .Z(n19287) );
  XOR U18860 ( .A(p_input[5861]), .B(p_input[5829]), .Z(n19288) );
  XNOR U18861 ( .A(n18992), .B(n19283), .Z(n19285) );
  XOR U18862 ( .A(n19289), .B(n19290), .Z(n18992) );
  AND U18863 ( .A(n321), .B(n19291), .Z(n19290) );
  XOR U18864 ( .A(p_input[5797]), .B(p_input[5765]), .Z(n19291) );
  XOR U18865 ( .A(n19292), .B(n19293), .Z(n19283) );
  AND U18866 ( .A(n19294), .B(n19295), .Z(n19293) );
  XOR U18867 ( .A(n19292), .B(n19007), .Z(n19295) );
  XNOR U18868 ( .A(p_input[5828]), .B(n19296), .Z(n19007) );
  AND U18869 ( .A(n323), .B(n19297), .Z(n19296) );
  XOR U18870 ( .A(p_input[5860]), .B(p_input[5828]), .Z(n19297) );
  XNOR U18871 ( .A(n19004), .B(n19292), .Z(n19294) );
  XOR U18872 ( .A(n19298), .B(n19299), .Z(n19004) );
  AND U18873 ( .A(n321), .B(n19300), .Z(n19299) );
  XOR U18874 ( .A(p_input[5796]), .B(p_input[5764]), .Z(n19300) );
  XOR U18875 ( .A(n19301), .B(n19302), .Z(n19292) );
  AND U18876 ( .A(n19303), .B(n19304), .Z(n19302) );
  XOR U18877 ( .A(n19301), .B(n19019), .Z(n19304) );
  XNOR U18878 ( .A(p_input[5827]), .B(n19305), .Z(n19019) );
  AND U18879 ( .A(n323), .B(n19306), .Z(n19305) );
  XOR U18880 ( .A(p_input[5859]), .B(p_input[5827]), .Z(n19306) );
  XNOR U18881 ( .A(n19016), .B(n19301), .Z(n19303) );
  XOR U18882 ( .A(n19307), .B(n19308), .Z(n19016) );
  AND U18883 ( .A(n321), .B(n19309), .Z(n19308) );
  XOR U18884 ( .A(p_input[5795]), .B(p_input[5763]), .Z(n19309) );
  XOR U18885 ( .A(n19310), .B(n19311), .Z(n19301) );
  AND U18886 ( .A(n19312), .B(n19313), .Z(n19311) );
  XOR U18887 ( .A(n19310), .B(n19031), .Z(n19313) );
  XNOR U18888 ( .A(p_input[5826]), .B(n19314), .Z(n19031) );
  AND U18889 ( .A(n323), .B(n19315), .Z(n19314) );
  XOR U18890 ( .A(p_input[5858]), .B(p_input[5826]), .Z(n19315) );
  XNOR U18891 ( .A(n19028), .B(n19310), .Z(n19312) );
  XOR U18892 ( .A(n19316), .B(n19317), .Z(n19028) );
  AND U18893 ( .A(n321), .B(n19318), .Z(n19317) );
  XOR U18894 ( .A(p_input[5794]), .B(p_input[5762]), .Z(n19318) );
  XOR U18895 ( .A(n19319), .B(n19320), .Z(n19310) );
  AND U18896 ( .A(n19321), .B(n19322), .Z(n19320) );
  XNOR U18897 ( .A(n19323), .B(n19044), .Z(n19322) );
  XNOR U18898 ( .A(p_input[5825]), .B(n19324), .Z(n19044) );
  AND U18899 ( .A(n323), .B(n19325), .Z(n19324) );
  XNOR U18900 ( .A(p_input[5857]), .B(n19326), .Z(n19325) );
  IV U18901 ( .A(p_input[5825]), .Z(n19326) );
  XNOR U18902 ( .A(n19041), .B(n19319), .Z(n19321) );
  XNOR U18903 ( .A(p_input[5761]), .B(n19327), .Z(n19041) );
  AND U18904 ( .A(n321), .B(n19328), .Z(n19327) );
  XOR U18905 ( .A(p_input[5793]), .B(p_input[5761]), .Z(n19328) );
  IV U18906 ( .A(n19323), .Z(n19319) );
  AND U18907 ( .A(n19049), .B(n19052), .Z(n19323) );
  XOR U18908 ( .A(p_input[5824]), .B(n19329), .Z(n19052) );
  AND U18909 ( .A(n323), .B(n19330), .Z(n19329) );
  XOR U18910 ( .A(p_input[5856]), .B(p_input[5824]), .Z(n19330) );
  XOR U18911 ( .A(n19331), .B(n19332), .Z(n323) );
  AND U18912 ( .A(n19333), .B(n19334), .Z(n19332) );
  XNOR U18913 ( .A(p_input[5887]), .B(n19331), .Z(n19334) );
  XOR U18914 ( .A(n19331), .B(p_input[5855]), .Z(n19333) );
  XOR U18915 ( .A(n19335), .B(n19336), .Z(n19331) );
  AND U18916 ( .A(n19337), .B(n19338), .Z(n19336) );
  XNOR U18917 ( .A(p_input[5886]), .B(n19335), .Z(n19338) );
  XOR U18918 ( .A(n19335), .B(p_input[5854]), .Z(n19337) );
  XOR U18919 ( .A(n19339), .B(n19340), .Z(n19335) );
  AND U18920 ( .A(n19341), .B(n19342), .Z(n19340) );
  XNOR U18921 ( .A(p_input[5885]), .B(n19339), .Z(n19342) );
  XOR U18922 ( .A(n19339), .B(p_input[5853]), .Z(n19341) );
  XOR U18923 ( .A(n19343), .B(n19344), .Z(n19339) );
  AND U18924 ( .A(n19345), .B(n19346), .Z(n19344) );
  XNOR U18925 ( .A(p_input[5884]), .B(n19343), .Z(n19346) );
  XOR U18926 ( .A(n19343), .B(p_input[5852]), .Z(n19345) );
  XOR U18927 ( .A(n19347), .B(n19348), .Z(n19343) );
  AND U18928 ( .A(n19349), .B(n19350), .Z(n19348) );
  XNOR U18929 ( .A(p_input[5883]), .B(n19347), .Z(n19350) );
  XOR U18930 ( .A(n19347), .B(p_input[5851]), .Z(n19349) );
  XOR U18931 ( .A(n19351), .B(n19352), .Z(n19347) );
  AND U18932 ( .A(n19353), .B(n19354), .Z(n19352) );
  XNOR U18933 ( .A(p_input[5882]), .B(n19351), .Z(n19354) );
  XOR U18934 ( .A(n19351), .B(p_input[5850]), .Z(n19353) );
  XOR U18935 ( .A(n19355), .B(n19356), .Z(n19351) );
  AND U18936 ( .A(n19357), .B(n19358), .Z(n19356) );
  XNOR U18937 ( .A(p_input[5881]), .B(n19355), .Z(n19358) );
  XOR U18938 ( .A(n19355), .B(p_input[5849]), .Z(n19357) );
  XOR U18939 ( .A(n19359), .B(n19360), .Z(n19355) );
  AND U18940 ( .A(n19361), .B(n19362), .Z(n19360) );
  XNOR U18941 ( .A(p_input[5880]), .B(n19359), .Z(n19362) );
  XOR U18942 ( .A(n19359), .B(p_input[5848]), .Z(n19361) );
  XOR U18943 ( .A(n19363), .B(n19364), .Z(n19359) );
  AND U18944 ( .A(n19365), .B(n19366), .Z(n19364) );
  XNOR U18945 ( .A(p_input[5879]), .B(n19363), .Z(n19366) );
  XOR U18946 ( .A(n19363), .B(p_input[5847]), .Z(n19365) );
  XOR U18947 ( .A(n19367), .B(n19368), .Z(n19363) );
  AND U18948 ( .A(n19369), .B(n19370), .Z(n19368) );
  XNOR U18949 ( .A(p_input[5878]), .B(n19367), .Z(n19370) );
  XOR U18950 ( .A(n19367), .B(p_input[5846]), .Z(n19369) );
  XOR U18951 ( .A(n19371), .B(n19372), .Z(n19367) );
  AND U18952 ( .A(n19373), .B(n19374), .Z(n19372) );
  XNOR U18953 ( .A(p_input[5877]), .B(n19371), .Z(n19374) );
  XOR U18954 ( .A(n19371), .B(p_input[5845]), .Z(n19373) );
  XOR U18955 ( .A(n19375), .B(n19376), .Z(n19371) );
  AND U18956 ( .A(n19377), .B(n19378), .Z(n19376) );
  XNOR U18957 ( .A(p_input[5876]), .B(n19375), .Z(n19378) );
  XOR U18958 ( .A(n19375), .B(p_input[5844]), .Z(n19377) );
  XOR U18959 ( .A(n19379), .B(n19380), .Z(n19375) );
  AND U18960 ( .A(n19381), .B(n19382), .Z(n19380) );
  XNOR U18961 ( .A(p_input[5875]), .B(n19379), .Z(n19382) );
  XOR U18962 ( .A(n19379), .B(p_input[5843]), .Z(n19381) );
  XOR U18963 ( .A(n19383), .B(n19384), .Z(n19379) );
  AND U18964 ( .A(n19385), .B(n19386), .Z(n19384) );
  XNOR U18965 ( .A(p_input[5874]), .B(n19383), .Z(n19386) );
  XOR U18966 ( .A(n19383), .B(p_input[5842]), .Z(n19385) );
  XOR U18967 ( .A(n19387), .B(n19388), .Z(n19383) );
  AND U18968 ( .A(n19389), .B(n19390), .Z(n19388) );
  XNOR U18969 ( .A(p_input[5873]), .B(n19387), .Z(n19390) );
  XOR U18970 ( .A(n19387), .B(p_input[5841]), .Z(n19389) );
  XOR U18971 ( .A(n19391), .B(n19392), .Z(n19387) );
  AND U18972 ( .A(n19393), .B(n19394), .Z(n19392) );
  XNOR U18973 ( .A(p_input[5872]), .B(n19391), .Z(n19394) );
  XOR U18974 ( .A(n19391), .B(p_input[5840]), .Z(n19393) );
  XOR U18975 ( .A(n19395), .B(n19396), .Z(n19391) );
  AND U18976 ( .A(n19397), .B(n19398), .Z(n19396) );
  XNOR U18977 ( .A(p_input[5871]), .B(n19395), .Z(n19398) );
  XOR U18978 ( .A(n19395), .B(p_input[5839]), .Z(n19397) );
  XOR U18979 ( .A(n19399), .B(n19400), .Z(n19395) );
  AND U18980 ( .A(n19401), .B(n19402), .Z(n19400) );
  XNOR U18981 ( .A(p_input[5870]), .B(n19399), .Z(n19402) );
  XOR U18982 ( .A(n19399), .B(p_input[5838]), .Z(n19401) );
  XOR U18983 ( .A(n19403), .B(n19404), .Z(n19399) );
  AND U18984 ( .A(n19405), .B(n19406), .Z(n19404) );
  XNOR U18985 ( .A(p_input[5869]), .B(n19403), .Z(n19406) );
  XOR U18986 ( .A(n19403), .B(p_input[5837]), .Z(n19405) );
  XOR U18987 ( .A(n19407), .B(n19408), .Z(n19403) );
  AND U18988 ( .A(n19409), .B(n19410), .Z(n19408) );
  XNOR U18989 ( .A(p_input[5868]), .B(n19407), .Z(n19410) );
  XOR U18990 ( .A(n19407), .B(p_input[5836]), .Z(n19409) );
  XOR U18991 ( .A(n19411), .B(n19412), .Z(n19407) );
  AND U18992 ( .A(n19413), .B(n19414), .Z(n19412) );
  XNOR U18993 ( .A(p_input[5867]), .B(n19411), .Z(n19414) );
  XOR U18994 ( .A(n19411), .B(p_input[5835]), .Z(n19413) );
  XOR U18995 ( .A(n19415), .B(n19416), .Z(n19411) );
  AND U18996 ( .A(n19417), .B(n19418), .Z(n19416) );
  XNOR U18997 ( .A(p_input[5866]), .B(n19415), .Z(n19418) );
  XOR U18998 ( .A(n19415), .B(p_input[5834]), .Z(n19417) );
  XOR U18999 ( .A(n19419), .B(n19420), .Z(n19415) );
  AND U19000 ( .A(n19421), .B(n19422), .Z(n19420) );
  XNOR U19001 ( .A(p_input[5865]), .B(n19419), .Z(n19422) );
  XOR U19002 ( .A(n19419), .B(p_input[5833]), .Z(n19421) );
  XOR U19003 ( .A(n19423), .B(n19424), .Z(n19419) );
  AND U19004 ( .A(n19425), .B(n19426), .Z(n19424) );
  XNOR U19005 ( .A(p_input[5864]), .B(n19423), .Z(n19426) );
  XOR U19006 ( .A(n19423), .B(p_input[5832]), .Z(n19425) );
  XOR U19007 ( .A(n19427), .B(n19428), .Z(n19423) );
  AND U19008 ( .A(n19429), .B(n19430), .Z(n19428) );
  XNOR U19009 ( .A(p_input[5863]), .B(n19427), .Z(n19430) );
  XOR U19010 ( .A(n19427), .B(p_input[5831]), .Z(n19429) );
  XOR U19011 ( .A(n19431), .B(n19432), .Z(n19427) );
  AND U19012 ( .A(n19433), .B(n19434), .Z(n19432) );
  XNOR U19013 ( .A(p_input[5862]), .B(n19431), .Z(n19434) );
  XOR U19014 ( .A(n19431), .B(p_input[5830]), .Z(n19433) );
  XOR U19015 ( .A(n19435), .B(n19436), .Z(n19431) );
  AND U19016 ( .A(n19437), .B(n19438), .Z(n19436) );
  XNOR U19017 ( .A(p_input[5861]), .B(n19435), .Z(n19438) );
  XOR U19018 ( .A(n19435), .B(p_input[5829]), .Z(n19437) );
  XOR U19019 ( .A(n19439), .B(n19440), .Z(n19435) );
  AND U19020 ( .A(n19441), .B(n19442), .Z(n19440) );
  XNOR U19021 ( .A(p_input[5860]), .B(n19439), .Z(n19442) );
  XOR U19022 ( .A(n19439), .B(p_input[5828]), .Z(n19441) );
  XOR U19023 ( .A(n19443), .B(n19444), .Z(n19439) );
  AND U19024 ( .A(n19445), .B(n19446), .Z(n19444) );
  XNOR U19025 ( .A(p_input[5859]), .B(n19443), .Z(n19446) );
  XOR U19026 ( .A(n19443), .B(p_input[5827]), .Z(n19445) );
  XOR U19027 ( .A(n19447), .B(n19448), .Z(n19443) );
  AND U19028 ( .A(n19449), .B(n19450), .Z(n19448) );
  XNOR U19029 ( .A(p_input[5858]), .B(n19447), .Z(n19450) );
  XOR U19030 ( .A(n19447), .B(p_input[5826]), .Z(n19449) );
  XNOR U19031 ( .A(n19451), .B(n19452), .Z(n19447) );
  AND U19032 ( .A(n19453), .B(n19454), .Z(n19452) );
  XOR U19033 ( .A(p_input[5857]), .B(n19451), .Z(n19454) );
  XNOR U19034 ( .A(p_input[5825]), .B(n19451), .Z(n19453) );
  AND U19035 ( .A(p_input[5856]), .B(n19455), .Z(n19451) );
  IV U19036 ( .A(p_input[5824]), .Z(n19455) );
  XNOR U19037 ( .A(p_input[5760]), .B(n19456), .Z(n19049) );
  AND U19038 ( .A(n321), .B(n19457), .Z(n19456) );
  XOR U19039 ( .A(p_input[5792]), .B(p_input[5760]), .Z(n19457) );
  XOR U19040 ( .A(n19458), .B(n19459), .Z(n321) );
  AND U19041 ( .A(n19460), .B(n19461), .Z(n19459) );
  XNOR U19042 ( .A(p_input[5823]), .B(n19458), .Z(n19461) );
  XOR U19043 ( .A(n19458), .B(p_input[5791]), .Z(n19460) );
  XOR U19044 ( .A(n19462), .B(n19463), .Z(n19458) );
  AND U19045 ( .A(n19464), .B(n19465), .Z(n19463) );
  XNOR U19046 ( .A(p_input[5822]), .B(n19462), .Z(n19465) );
  XNOR U19047 ( .A(n19462), .B(n19064), .Z(n19464) );
  IV U19048 ( .A(p_input[5790]), .Z(n19064) );
  XOR U19049 ( .A(n19466), .B(n19467), .Z(n19462) );
  AND U19050 ( .A(n19468), .B(n19469), .Z(n19467) );
  XNOR U19051 ( .A(p_input[5821]), .B(n19466), .Z(n19469) );
  XNOR U19052 ( .A(n19466), .B(n19073), .Z(n19468) );
  IV U19053 ( .A(p_input[5789]), .Z(n19073) );
  XOR U19054 ( .A(n19470), .B(n19471), .Z(n19466) );
  AND U19055 ( .A(n19472), .B(n19473), .Z(n19471) );
  XNOR U19056 ( .A(p_input[5820]), .B(n19470), .Z(n19473) );
  XNOR U19057 ( .A(n19470), .B(n19082), .Z(n19472) );
  IV U19058 ( .A(p_input[5788]), .Z(n19082) );
  XOR U19059 ( .A(n19474), .B(n19475), .Z(n19470) );
  AND U19060 ( .A(n19476), .B(n19477), .Z(n19475) );
  XNOR U19061 ( .A(p_input[5819]), .B(n19474), .Z(n19477) );
  XNOR U19062 ( .A(n19474), .B(n19091), .Z(n19476) );
  IV U19063 ( .A(p_input[5787]), .Z(n19091) );
  XOR U19064 ( .A(n19478), .B(n19479), .Z(n19474) );
  AND U19065 ( .A(n19480), .B(n19481), .Z(n19479) );
  XNOR U19066 ( .A(p_input[5818]), .B(n19478), .Z(n19481) );
  XNOR U19067 ( .A(n19478), .B(n19100), .Z(n19480) );
  IV U19068 ( .A(p_input[5786]), .Z(n19100) );
  XOR U19069 ( .A(n19482), .B(n19483), .Z(n19478) );
  AND U19070 ( .A(n19484), .B(n19485), .Z(n19483) );
  XNOR U19071 ( .A(p_input[5817]), .B(n19482), .Z(n19485) );
  XNOR U19072 ( .A(n19482), .B(n19109), .Z(n19484) );
  IV U19073 ( .A(p_input[5785]), .Z(n19109) );
  XOR U19074 ( .A(n19486), .B(n19487), .Z(n19482) );
  AND U19075 ( .A(n19488), .B(n19489), .Z(n19487) );
  XNOR U19076 ( .A(p_input[5816]), .B(n19486), .Z(n19489) );
  XNOR U19077 ( .A(n19486), .B(n19118), .Z(n19488) );
  IV U19078 ( .A(p_input[5784]), .Z(n19118) );
  XOR U19079 ( .A(n19490), .B(n19491), .Z(n19486) );
  AND U19080 ( .A(n19492), .B(n19493), .Z(n19491) );
  XNOR U19081 ( .A(p_input[5815]), .B(n19490), .Z(n19493) );
  XNOR U19082 ( .A(n19490), .B(n19127), .Z(n19492) );
  IV U19083 ( .A(p_input[5783]), .Z(n19127) );
  XOR U19084 ( .A(n19494), .B(n19495), .Z(n19490) );
  AND U19085 ( .A(n19496), .B(n19497), .Z(n19495) );
  XNOR U19086 ( .A(p_input[5814]), .B(n19494), .Z(n19497) );
  XNOR U19087 ( .A(n19494), .B(n19136), .Z(n19496) );
  IV U19088 ( .A(p_input[5782]), .Z(n19136) );
  XOR U19089 ( .A(n19498), .B(n19499), .Z(n19494) );
  AND U19090 ( .A(n19500), .B(n19501), .Z(n19499) );
  XNOR U19091 ( .A(p_input[5813]), .B(n19498), .Z(n19501) );
  XNOR U19092 ( .A(n19498), .B(n19145), .Z(n19500) );
  IV U19093 ( .A(p_input[5781]), .Z(n19145) );
  XOR U19094 ( .A(n19502), .B(n19503), .Z(n19498) );
  AND U19095 ( .A(n19504), .B(n19505), .Z(n19503) );
  XNOR U19096 ( .A(p_input[5812]), .B(n19502), .Z(n19505) );
  XNOR U19097 ( .A(n19502), .B(n19154), .Z(n19504) );
  IV U19098 ( .A(p_input[5780]), .Z(n19154) );
  XOR U19099 ( .A(n19506), .B(n19507), .Z(n19502) );
  AND U19100 ( .A(n19508), .B(n19509), .Z(n19507) );
  XNOR U19101 ( .A(p_input[5811]), .B(n19506), .Z(n19509) );
  XNOR U19102 ( .A(n19506), .B(n19163), .Z(n19508) );
  IV U19103 ( .A(p_input[5779]), .Z(n19163) );
  XOR U19104 ( .A(n19510), .B(n19511), .Z(n19506) );
  AND U19105 ( .A(n19512), .B(n19513), .Z(n19511) );
  XNOR U19106 ( .A(p_input[5810]), .B(n19510), .Z(n19513) );
  XNOR U19107 ( .A(n19510), .B(n19172), .Z(n19512) );
  IV U19108 ( .A(p_input[5778]), .Z(n19172) );
  XOR U19109 ( .A(n19514), .B(n19515), .Z(n19510) );
  AND U19110 ( .A(n19516), .B(n19517), .Z(n19515) );
  XNOR U19111 ( .A(p_input[5809]), .B(n19514), .Z(n19517) );
  XNOR U19112 ( .A(n19514), .B(n19181), .Z(n19516) );
  IV U19113 ( .A(p_input[5777]), .Z(n19181) );
  XOR U19114 ( .A(n19518), .B(n19519), .Z(n19514) );
  AND U19115 ( .A(n19520), .B(n19521), .Z(n19519) );
  XNOR U19116 ( .A(p_input[5808]), .B(n19518), .Z(n19521) );
  XNOR U19117 ( .A(n19518), .B(n19190), .Z(n19520) );
  IV U19118 ( .A(p_input[5776]), .Z(n19190) );
  XOR U19119 ( .A(n19522), .B(n19523), .Z(n19518) );
  AND U19120 ( .A(n19524), .B(n19525), .Z(n19523) );
  XNOR U19121 ( .A(p_input[5807]), .B(n19522), .Z(n19525) );
  XNOR U19122 ( .A(n19522), .B(n19199), .Z(n19524) );
  IV U19123 ( .A(p_input[5775]), .Z(n19199) );
  XOR U19124 ( .A(n19526), .B(n19527), .Z(n19522) );
  AND U19125 ( .A(n19528), .B(n19529), .Z(n19527) );
  XNOR U19126 ( .A(p_input[5806]), .B(n19526), .Z(n19529) );
  XNOR U19127 ( .A(n19526), .B(n19208), .Z(n19528) );
  IV U19128 ( .A(p_input[5774]), .Z(n19208) );
  XOR U19129 ( .A(n19530), .B(n19531), .Z(n19526) );
  AND U19130 ( .A(n19532), .B(n19533), .Z(n19531) );
  XNOR U19131 ( .A(p_input[5805]), .B(n19530), .Z(n19533) );
  XNOR U19132 ( .A(n19530), .B(n19217), .Z(n19532) );
  IV U19133 ( .A(p_input[5773]), .Z(n19217) );
  XOR U19134 ( .A(n19534), .B(n19535), .Z(n19530) );
  AND U19135 ( .A(n19536), .B(n19537), .Z(n19535) );
  XNOR U19136 ( .A(p_input[5804]), .B(n19534), .Z(n19537) );
  XNOR U19137 ( .A(n19534), .B(n19226), .Z(n19536) );
  IV U19138 ( .A(p_input[5772]), .Z(n19226) );
  XOR U19139 ( .A(n19538), .B(n19539), .Z(n19534) );
  AND U19140 ( .A(n19540), .B(n19541), .Z(n19539) );
  XNOR U19141 ( .A(p_input[5803]), .B(n19538), .Z(n19541) );
  XNOR U19142 ( .A(n19538), .B(n19235), .Z(n19540) );
  IV U19143 ( .A(p_input[5771]), .Z(n19235) );
  XOR U19144 ( .A(n19542), .B(n19543), .Z(n19538) );
  AND U19145 ( .A(n19544), .B(n19545), .Z(n19543) );
  XNOR U19146 ( .A(p_input[5802]), .B(n19542), .Z(n19545) );
  XNOR U19147 ( .A(n19542), .B(n19244), .Z(n19544) );
  IV U19148 ( .A(p_input[5770]), .Z(n19244) );
  XOR U19149 ( .A(n19546), .B(n19547), .Z(n19542) );
  AND U19150 ( .A(n19548), .B(n19549), .Z(n19547) );
  XNOR U19151 ( .A(p_input[5801]), .B(n19546), .Z(n19549) );
  XNOR U19152 ( .A(n19546), .B(n19253), .Z(n19548) );
  IV U19153 ( .A(p_input[5769]), .Z(n19253) );
  XOR U19154 ( .A(n19550), .B(n19551), .Z(n19546) );
  AND U19155 ( .A(n19552), .B(n19553), .Z(n19551) );
  XNOR U19156 ( .A(p_input[5800]), .B(n19550), .Z(n19553) );
  XNOR U19157 ( .A(n19550), .B(n19262), .Z(n19552) );
  IV U19158 ( .A(p_input[5768]), .Z(n19262) );
  XOR U19159 ( .A(n19554), .B(n19555), .Z(n19550) );
  AND U19160 ( .A(n19556), .B(n19557), .Z(n19555) );
  XNOR U19161 ( .A(p_input[5799]), .B(n19554), .Z(n19557) );
  XNOR U19162 ( .A(n19554), .B(n19271), .Z(n19556) );
  IV U19163 ( .A(p_input[5767]), .Z(n19271) );
  XOR U19164 ( .A(n19558), .B(n19559), .Z(n19554) );
  AND U19165 ( .A(n19560), .B(n19561), .Z(n19559) );
  XNOR U19166 ( .A(p_input[5798]), .B(n19558), .Z(n19561) );
  XNOR U19167 ( .A(n19558), .B(n19280), .Z(n19560) );
  IV U19168 ( .A(p_input[5766]), .Z(n19280) );
  XOR U19169 ( .A(n19562), .B(n19563), .Z(n19558) );
  AND U19170 ( .A(n19564), .B(n19565), .Z(n19563) );
  XNOR U19171 ( .A(p_input[5797]), .B(n19562), .Z(n19565) );
  XNOR U19172 ( .A(n19562), .B(n19289), .Z(n19564) );
  IV U19173 ( .A(p_input[5765]), .Z(n19289) );
  XOR U19174 ( .A(n19566), .B(n19567), .Z(n19562) );
  AND U19175 ( .A(n19568), .B(n19569), .Z(n19567) );
  XNOR U19176 ( .A(p_input[5796]), .B(n19566), .Z(n19569) );
  XNOR U19177 ( .A(n19566), .B(n19298), .Z(n19568) );
  IV U19178 ( .A(p_input[5764]), .Z(n19298) );
  XOR U19179 ( .A(n19570), .B(n19571), .Z(n19566) );
  AND U19180 ( .A(n19572), .B(n19573), .Z(n19571) );
  XNOR U19181 ( .A(p_input[5795]), .B(n19570), .Z(n19573) );
  XNOR U19182 ( .A(n19570), .B(n19307), .Z(n19572) );
  IV U19183 ( .A(p_input[5763]), .Z(n19307) );
  XOR U19184 ( .A(n19574), .B(n19575), .Z(n19570) );
  AND U19185 ( .A(n19576), .B(n19577), .Z(n19575) );
  XNOR U19186 ( .A(p_input[5794]), .B(n19574), .Z(n19577) );
  XNOR U19187 ( .A(n19574), .B(n19316), .Z(n19576) );
  IV U19188 ( .A(p_input[5762]), .Z(n19316) );
  XNOR U19189 ( .A(n19578), .B(n19579), .Z(n19574) );
  AND U19190 ( .A(n19580), .B(n19581), .Z(n19579) );
  XOR U19191 ( .A(p_input[5793]), .B(n19578), .Z(n19581) );
  XNOR U19192 ( .A(p_input[5761]), .B(n19578), .Z(n19580) );
  AND U19193 ( .A(p_input[5792]), .B(n19582), .Z(n19578) );
  IV U19194 ( .A(p_input[5760]), .Z(n19582) );
  XOR U19195 ( .A(n19583), .B(n19584), .Z(n18672) );
  AND U19196 ( .A(n500), .B(n19585), .Z(n19584) );
  XNOR U19197 ( .A(n19586), .B(n19583), .Z(n19585) );
  XOR U19198 ( .A(n19587), .B(n19588), .Z(n500) );
  AND U19199 ( .A(n19589), .B(n19590), .Z(n19588) );
  XNOR U19200 ( .A(n18687), .B(n19587), .Z(n19590) );
  AND U19201 ( .A(p_input[5759]), .B(p_input[5727]), .Z(n18687) );
  XNOR U19202 ( .A(n19587), .B(n18684), .Z(n19589) );
  IV U19203 ( .A(n19591), .Z(n18684) );
  AND U19204 ( .A(p_input[5663]), .B(p_input[5695]), .Z(n19591) );
  XOR U19205 ( .A(n19592), .B(n19593), .Z(n19587) );
  AND U19206 ( .A(n19594), .B(n19595), .Z(n19593) );
  XOR U19207 ( .A(n19592), .B(n18699), .Z(n19595) );
  XNOR U19208 ( .A(p_input[5726]), .B(n19596), .Z(n18699) );
  AND U19209 ( .A(n327), .B(n19597), .Z(n19596) );
  XOR U19210 ( .A(p_input[5758]), .B(p_input[5726]), .Z(n19597) );
  XNOR U19211 ( .A(n18696), .B(n19592), .Z(n19594) );
  XOR U19212 ( .A(n19598), .B(n19599), .Z(n18696) );
  AND U19213 ( .A(n324), .B(n19600), .Z(n19599) );
  XOR U19214 ( .A(p_input[5694]), .B(p_input[5662]), .Z(n19600) );
  XOR U19215 ( .A(n19601), .B(n19602), .Z(n19592) );
  AND U19216 ( .A(n19603), .B(n19604), .Z(n19602) );
  XOR U19217 ( .A(n19601), .B(n18711), .Z(n19604) );
  XNOR U19218 ( .A(p_input[5725]), .B(n19605), .Z(n18711) );
  AND U19219 ( .A(n327), .B(n19606), .Z(n19605) );
  XOR U19220 ( .A(p_input[5757]), .B(p_input[5725]), .Z(n19606) );
  XNOR U19221 ( .A(n18708), .B(n19601), .Z(n19603) );
  XOR U19222 ( .A(n19607), .B(n19608), .Z(n18708) );
  AND U19223 ( .A(n324), .B(n19609), .Z(n19608) );
  XOR U19224 ( .A(p_input[5693]), .B(p_input[5661]), .Z(n19609) );
  XOR U19225 ( .A(n19610), .B(n19611), .Z(n19601) );
  AND U19226 ( .A(n19612), .B(n19613), .Z(n19611) );
  XOR U19227 ( .A(n19610), .B(n18723), .Z(n19613) );
  XNOR U19228 ( .A(p_input[5724]), .B(n19614), .Z(n18723) );
  AND U19229 ( .A(n327), .B(n19615), .Z(n19614) );
  XOR U19230 ( .A(p_input[5756]), .B(p_input[5724]), .Z(n19615) );
  XNOR U19231 ( .A(n18720), .B(n19610), .Z(n19612) );
  XOR U19232 ( .A(n19616), .B(n19617), .Z(n18720) );
  AND U19233 ( .A(n324), .B(n19618), .Z(n19617) );
  XOR U19234 ( .A(p_input[5692]), .B(p_input[5660]), .Z(n19618) );
  XOR U19235 ( .A(n19619), .B(n19620), .Z(n19610) );
  AND U19236 ( .A(n19621), .B(n19622), .Z(n19620) );
  XOR U19237 ( .A(n19619), .B(n18735), .Z(n19622) );
  XNOR U19238 ( .A(p_input[5723]), .B(n19623), .Z(n18735) );
  AND U19239 ( .A(n327), .B(n19624), .Z(n19623) );
  XOR U19240 ( .A(p_input[5755]), .B(p_input[5723]), .Z(n19624) );
  XNOR U19241 ( .A(n18732), .B(n19619), .Z(n19621) );
  XOR U19242 ( .A(n19625), .B(n19626), .Z(n18732) );
  AND U19243 ( .A(n324), .B(n19627), .Z(n19626) );
  XOR U19244 ( .A(p_input[5691]), .B(p_input[5659]), .Z(n19627) );
  XOR U19245 ( .A(n19628), .B(n19629), .Z(n19619) );
  AND U19246 ( .A(n19630), .B(n19631), .Z(n19629) );
  XOR U19247 ( .A(n19628), .B(n18747), .Z(n19631) );
  XNOR U19248 ( .A(p_input[5722]), .B(n19632), .Z(n18747) );
  AND U19249 ( .A(n327), .B(n19633), .Z(n19632) );
  XOR U19250 ( .A(p_input[5754]), .B(p_input[5722]), .Z(n19633) );
  XNOR U19251 ( .A(n18744), .B(n19628), .Z(n19630) );
  XOR U19252 ( .A(n19634), .B(n19635), .Z(n18744) );
  AND U19253 ( .A(n324), .B(n19636), .Z(n19635) );
  XOR U19254 ( .A(p_input[5690]), .B(p_input[5658]), .Z(n19636) );
  XOR U19255 ( .A(n19637), .B(n19638), .Z(n19628) );
  AND U19256 ( .A(n19639), .B(n19640), .Z(n19638) );
  XOR U19257 ( .A(n19637), .B(n18759), .Z(n19640) );
  XNOR U19258 ( .A(p_input[5721]), .B(n19641), .Z(n18759) );
  AND U19259 ( .A(n327), .B(n19642), .Z(n19641) );
  XOR U19260 ( .A(p_input[5753]), .B(p_input[5721]), .Z(n19642) );
  XNOR U19261 ( .A(n18756), .B(n19637), .Z(n19639) );
  XOR U19262 ( .A(n19643), .B(n19644), .Z(n18756) );
  AND U19263 ( .A(n324), .B(n19645), .Z(n19644) );
  XOR U19264 ( .A(p_input[5689]), .B(p_input[5657]), .Z(n19645) );
  XOR U19265 ( .A(n19646), .B(n19647), .Z(n19637) );
  AND U19266 ( .A(n19648), .B(n19649), .Z(n19647) );
  XOR U19267 ( .A(n19646), .B(n18771), .Z(n19649) );
  XNOR U19268 ( .A(p_input[5720]), .B(n19650), .Z(n18771) );
  AND U19269 ( .A(n327), .B(n19651), .Z(n19650) );
  XOR U19270 ( .A(p_input[5752]), .B(p_input[5720]), .Z(n19651) );
  XNOR U19271 ( .A(n18768), .B(n19646), .Z(n19648) );
  XOR U19272 ( .A(n19652), .B(n19653), .Z(n18768) );
  AND U19273 ( .A(n324), .B(n19654), .Z(n19653) );
  XOR U19274 ( .A(p_input[5688]), .B(p_input[5656]), .Z(n19654) );
  XOR U19275 ( .A(n19655), .B(n19656), .Z(n19646) );
  AND U19276 ( .A(n19657), .B(n19658), .Z(n19656) );
  XOR U19277 ( .A(n19655), .B(n18783), .Z(n19658) );
  XNOR U19278 ( .A(p_input[5719]), .B(n19659), .Z(n18783) );
  AND U19279 ( .A(n327), .B(n19660), .Z(n19659) );
  XOR U19280 ( .A(p_input[5751]), .B(p_input[5719]), .Z(n19660) );
  XNOR U19281 ( .A(n18780), .B(n19655), .Z(n19657) );
  XOR U19282 ( .A(n19661), .B(n19662), .Z(n18780) );
  AND U19283 ( .A(n324), .B(n19663), .Z(n19662) );
  XOR U19284 ( .A(p_input[5687]), .B(p_input[5655]), .Z(n19663) );
  XOR U19285 ( .A(n19664), .B(n19665), .Z(n19655) );
  AND U19286 ( .A(n19666), .B(n19667), .Z(n19665) );
  XOR U19287 ( .A(n19664), .B(n18795), .Z(n19667) );
  XNOR U19288 ( .A(p_input[5718]), .B(n19668), .Z(n18795) );
  AND U19289 ( .A(n327), .B(n19669), .Z(n19668) );
  XOR U19290 ( .A(p_input[5750]), .B(p_input[5718]), .Z(n19669) );
  XNOR U19291 ( .A(n18792), .B(n19664), .Z(n19666) );
  XOR U19292 ( .A(n19670), .B(n19671), .Z(n18792) );
  AND U19293 ( .A(n324), .B(n19672), .Z(n19671) );
  XOR U19294 ( .A(p_input[5686]), .B(p_input[5654]), .Z(n19672) );
  XOR U19295 ( .A(n19673), .B(n19674), .Z(n19664) );
  AND U19296 ( .A(n19675), .B(n19676), .Z(n19674) );
  XOR U19297 ( .A(n19673), .B(n18807), .Z(n19676) );
  XNOR U19298 ( .A(p_input[5717]), .B(n19677), .Z(n18807) );
  AND U19299 ( .A(n327), .B(n19678), .Z(n19677) );
  XOR U19300 ( .A(p_input[5749]), .B(p_input[5717]), .Z(n19678) );
  XNOR U19301 ( .A(n18804), .B(n19673), .Z(n19675) );
  XOR U19302 ( .A(n19679), .B(n19680), .Z(n18804) );
  AND U19303 ( .A(n324), .B(n19681), .Z(n19680) );
  XOR U19304 ( .A(p_input[5685]), .B(p_input[5653]), .Z(n19681) );
  XOR U19305 ( .A(n19682), .B(n19683), .Z(n19673) );
  AND U19306 ( .A(n19684), .B(n19685), .Z(n19683) );
  XOR U19307 ( .A(n19682), .B(n18819), .Z(n19685) );
  XNOR U19308 ( .A(p_input[5716]), .B(n19686), .Z(n18819) );
  AND U19309 ( .A(n327), .B(n19687), .Z(n19686) );
  XOR U19310 ( .A(p_input[5748]), .B(p_input[5716]), .Z(n19687) );
  XNOR U19311 ( .A(n18816), .B(n19682), .Z(n19684) );
  XOR U19312 ( .A(n19688), .B(n19689), .Z(n18816) );
  AND U19313 ( .A(n324), .B(n19690), .Z(n19689) );
  XOR U19314 ( .A(p_input[5684]), .B(p_input[5652]), .Z(n19690) );
  XOR U19315 ( .A(n19691), .B(n19692), .Z(n19682) );
  AND U19316 ( .A(n19693), .B(n19694), .Z(n19692) );
  XOR U19317 ( .A(n19691), .B(n18831), .Z(n19694) );
  XNOR U19318 ( .A(p_input[5715]), .B(n19695), .Z(n18831) );
  AND U19319 ( .A(n327), .B(n19696), .Z(n19695) );
  XOR U19320 ( .A(p_input[5747]), .B(p_input[5715]), .Z(n19696) );
  XNOR U19321 ( .A(n18828), .B(n19691), .Z(n19693) );
  XOR U19322 ( .A(n19697), .B(n19698), .Z(n18828) );
  AND U19323 ( .A(n324), .B(n19699), .Z(n19698) );
  XOR U19324 ( .A(p_input[5683]), .B(p_input[5651]), .Z(n19699) );
  XOR U19325 ( .A(n19700), .B(n19701), .Z(n19691) );
  AND U19326 ( .A(n19702), .B(n19703), .Z(n19701) );
  XOR U19327 ( .A(n19700), .B(n18843), .Z(n19703) );
  XNOR U19328 ( .A(p_input[5714]), .B(n19704), .Z(n18843) );
  AND U19329 ( .A(n327), .B(n19705), .Z(n19704) );
  XOR U19330 ( .A(p_input[5746]), .B(p_input[5714]), .Z(n19705) );
  XNOR U19331 ( .A(n18840), .B(n19700), .Z(n19702) );
  XOR U19332 ( .A(n19706), .B(n19707), .Z(n18840) );
  AND U19333 ( .A(n324), .B(n19708), .Z(n19707) );
  XOR U19334 ( .A(p_input[5682]), .B(p_input[5650]), .Z(n19708) );
  XOR U19335 ( .A(n19709), .B(n19710), .Z(n19700) );
  AND U19336 ( .A(n19711), .B(n19712), .Z(n19710) );
  XOR U19337 ( .A(n19709), .B(n18855), .Z(n19712) );
  XNOR U19338 ( .A(p_input[5713]), .B(n19713), .Z(n18855) );
  AND U19339 ( .A(n327), .B(n19714), .Z(n19713) );
  XOR U19340 ( .A(p_input[5745]), .B(p_input[5713]), .Z(n19714) );
  XNOR U19341 ( .A(n18852), .B(n19709), .Z(n19711) );
  XOR U19342 ( .A(n19715), .B(n19716), .Z(n18852) );
  AND U19343 ( .A(n324), .B(n19717), .Z(n19716) );
  XOR U19344 ( .A(p_input[5681]), .B(p_input[5649]), .Z(n19717) );
  XOR U19345 ( .A(n19718), .B(n19719), .Z(n19709) );
  AND U19346 ( .A(n19720), .B(n19721), .Z(n19719) );
  XOR U19347 ( .A(n19718), .B(n18867), .Z(n19721) );
  XNOR U19348 ( .A(p_input[5712]), .B(n19722), .Z(n18867) );
  AND U19349 ( .A(n327), .B(n19723), .Z(n19722) );
  XOR U19350 ( .A(p_input[5744]), .B(p_input[5712]), .Z(n19723) );
  XNOR U19351 ( .A(n18864), .B(n19718), .Z(n19720) );
  XOR U19352 ( .A(n19724), .B(n19725), .Z(n18864) );
  AND U19353 ( .A(n324), .B(n19726), .Z(n19725) );
  XOR U19354 ( .A(p_input[5680]), .B(p_input[5648]), .Z(n19726) );
  XOR U19355 ( .A(n19727), .B(n19728), .Z(n19718) );
  AND U19356 ( .A(n19729), .B(n19730), .Z(n19728) );
  XOR U19357 ( .A(n19727), .B(n18879), .Z(n19730) );
  XNOR U19358 ( .A(p_input[5711]), .B(n19731), .Z(n18879) );
  AND U19359 ( .A(n327), .B(n19732), .Z(n19731) );
  XOR U19360 ( .A(p_input[5743]), .B(p_input[5711]), .Z(n19732) );
  XNOR U19361 ( .A(n18876), .B(n19727), .Z(n19729) );
  XOR U19362 ( .A(n19733), .B(n19734), .Z(n18876) );
  AND U19363 ( .A(n324), .B(n19735), .Z(n19734) );
  XOR U19364 ( .A(p_input[5679]), .B(p_input[5647]), .Z(n19735) );
  XOR U19365 ( .A(n19736), .B(n19737), .Z(n19727) );
  AND U19366 ( .A(n19738), .B(n19739), .Z(n19737) );
  XOR U19367 ( .A(n19736), .B(n18891), .Z(n19739) );
  XNOR U19368 ( .A(p_input[5710]), .B(n19740), .Z(n18891) );
  AND U19369 ( .A(n327), .B(n19741), .Z(n19740) );
  XOR U19370 ( .A(p_input[5742]), .B(p_input[5710]), .Z(n19741) );
  XNOR U19371 ( .A(n18888), .B(n19736), .Z(n19738) );
  XOR U19372 ( .A(n19742), .B(n19743), .Z(n18888) );
  AND U19373 ( .A(n324), .B(n19744), .Z(n19743) );
  XOR U19374 ( .A(p_input[5678]), .B(p_input[5646]), .Z(n19744) );
  XOR U19375 ( .A(n19745), .B(n19746), .Z(n19736) );
  AND U19376 ( .A(n19747), .B(n19748), .Z(n19746) );
  XOR U19377 ( .A(n19745), .B(n18903), .Z(n19748) );
  XNOR U19378 ( .A(p_input[5709]), .B(n19749), .Z(n18903) );
  AND U19379 ( .A(n327), .B(n19750), .Z(n19749) );
  XOR U19380 ( .A(p_input[5741]), .B(p_input[5709]), .Z(n19750) );
  XNOR U19381 ( .A(n18900), .B(n19745), .Z(n19747) );
  XOR U19382 ( .A(n19751), .B(n19752), .Z(n18900) );
  AND U19383 ( .A(n324), .B(n19753), .Z(n19752) );
  XOR U19384 ( .A(p_input[5677]), .B(p_input[5645]), .Z(n19753) );
  XOR U19385 ( .A(n19754), .B(n19755), .Z(n19745) );
  AND U19386 ( .A(n19756), .B(n19757), .Z(n19755) );
  XOR U19387 ( .A(n19754), .B(n18915), .Z(n19757) );
  XNOR U19388 ( .A(p_input[5708]), .B(n19758), .Z(n18915) );
  AND U19389 ( .A(n327), .B(n19759), .Z(n19758) );
  XOR U19390 ( .A(p_input[5740]), .B(p_input[5708]), .Z(n19759) );
  XNOR U19391 ( .A(n18912), .B(n19754), .Z(n19756) );
  XOR U19392 ( .A(n19760), .B(n19761), .Z(n18912) );
  AND U19393 ( .A(n324), .B(n19762), .Z(n19761) );
  XOR U19394 ( .A(p_input[5676]), .B(p_input[5644]), .Z(n19762) );
  XOR U19395 ( .A(n19763), .B(n19764), .Z(n19754) );
  AND U19396 ( .A(n19765), .B(n19766), .Z(n19764) );
  XOR U19397 ( .A(n19763), .B(n18927), .Z(n19766) );
  XNOR U19398 ( .A(p_input[5707]), .B(n19767), .Z(n18927) );
  AND U19399 ( .A(n327), .B(n19768), .Z(n19767) );
  XOR U19400 ( .A(p_input[5739]), .B(p_input[5707]), .Z(n19768) );
  XNOR U19401 ( .A(n18924), .B(n19763), .Z(n19765) );
  XOR U19402 ( .A(n19769), .B(n19770), .Z(n18924) );
  AND U19403 ( .A(n324), .B(n19771), .Z(n19770) );
  XOR U19404 ( .A(p_input[5675]), .B(p_input[5643]), .Z(n19771) );
  XOR U19405 ( .A(n19772), .B(n19773), .Z(n19763) );
  AND U19406 ( .A(n19774), .B(n19775), .Z(n19773) );
  XOR U19407 ( .A(n19772), .B(n18939), .Z(n19775) );
  XNOR U19408 ( .A(p_input[5706]), .B(n19776), .Z(n18939) );
  AND U19409 ( .A(n327), .B(n19777), .Z(n19776) );
  XOR U19410 ( .A(p_input[5738]), .B(p_input[5706]), .Z(n19777) );
  XNOR U19411 ( .A(n18936), .B(n19772), .Z(n19774) );
  XOR U19412 ( .A(n19778), .B(n19779), .Z(n18936) );
  AND U19413 ( .A(n324), .B(n19780), .Z(n19779) );
  XOR U19414 ( .A(p_input[5674]), .B(p_input[5642]), .Z(n19780) );
  XOR U19415 ( .A(n19781), .B(n19782), .Z(n19772) );
  AND U19416 ( .A(n19783), .B(n19784), .Z(n19782) );
  XOR U19417 ( .A(n19781), .B(n18951), .Z(n19784) );
  XNOR U19418 ( .A(p_input[5705]), .B(n19785), .Z(n18951) );
  AND U19419 ( .A(n327), .B(n19786), .Z(n19785) );
  XOR U19420 ( .A(p_input[5737]), .B(p_input[5705]), .Z(n19786) );
  XNOR U19421 ( .A(n18948), .B(n19781), .Z(n19783) );
  XOR U19422 ( .A(n19787), .B(n19788), .Z(n18948) );
  AND U19423 ( .A(n324), .B(n19789), .Z(n19788) );
  XOR U19424 ( .A(p_input[5673]), .B(p_input[5641]), .Z(n19789) );
  XOR U19425 ( .A(n19790), .B(n19791), .Z(n19781) );
  AND U19426 ( .A(n19792), .B(n19793), .Z(n19791) );
  XOR U19427 ( .A(n19790), .B(n18963), .Z(n19793) );
  XNOR U19428 ( .A(p_input[5704]), .B(n19794), .Z(n18963) );
  AND U19429 ( .A(n327), .B(n19795), .Z(n19794) );
  XOR U19430 ( .A(p_input[5736]), .B(p_input[5704]), .Z(n19795) );
  XNOR U19431 ( .A(n18960), .B(n19790), .Z(n19792) );
  XOR U19432 ( .A(n19796), .B(n19797), .Z(n18960) );
  AND U19433 ( .A(n324), .B(n19798), .Z(n19797) );
  XOR U19434 ( .A(p_input[5672]), .B(p_input[5640]), .Z(n19798) );
  XOR U19435 ( .A(n19799), .B(n19800), .Z(n19790) );
  AND U19436 ( .A(n19801), .B(n19802), .Z(n19800) );
  XOR U19437 ( .A(n19799), .B(n18975), .Z(n19802) );
  XNOR U19438 ( .A(p_input[5703]), .B(n19803), .Z(n18975) );
  AND U19439 ( .A(n327), .B(n19804), .Z(n19803) );
  XOR U19440 ( .A(p_input[5735]), .B(p_input[5703]), .Z(n19804) );
  XNOR U19441 ( .A(n18972), .B(n19799), .Z(n19801) );
  XOR U19442 ( .A(n19805), .B(n19806), .Z(n18972) );
  AND U19443 ( .A(n324), .B(n19807), .Z(n19806) );
  XOR U19444 ( .A(p_input[5671]), .B(p_input[5639]), .Z(n19807) );
  XOR U19445 ( .A(n19808), .B(n19809), .Z(n19799) );
  AND U19446 ( .A(n19810), .B(n19811), .Z(n19809) );
  XOR U19447 ( .A(n19808), .B(n18987), .Z(n19811) );
  XNOR U19448 ( .A(p_input[5702]), .B(n19812), .Z(n18987) );
  AND U19449 ( .A(n327), .B(n19813), .Z(n19812) );
  XOR U19450 ( .A(p_input[5734]), .B(p_input[5702]), .Z(n19813) );
  XNOR U19451 ( .A(n18984), .B(n19808), .Z(n19810) );
  XOR U19452 ( .A(n19814), .B(n19815), .Z(n18984) );
  AND U19453 ( .A(n324), .B(n19816), .Z(n19815) );
  XOR U19454 ( .A(p_input[5670]), .B(p_input[5638]), .Z(n19816) );
  XOR U19455 ( .A(n19817), .B(n19818), .Z(n19808) );
  AND U19456 ( .A(n19819), .B(n19820), .Z(n19818) );
  XOR U19457 ( .A(n19817), .B(n18999), .Z(n19820) );
  XNOR U19458 ( .A(p_input[5701]), .B(n19821), .Z(n18999) );
  AND U19459 ( .A(n327), .B(n19822), .Z(n19821) );
  XOR U19460 ( .A(p_input[5733]), .B(p_input[5701]), .Z(n19822) );
  XNOR U19461 ( .A(n18996), .B(n19817), .Z(n19819) );
  XOR U19462 ( .A(n19823), .B(n19824), .Z(n18996) );
  AND U19463 ( .A(n324), .B(n19825), .Z(n19824) );
  XOR U19464 ( .A(p_input[5669]), .B(p_input[5637]), .Z(n19825) );
  XOR U19465 ( .A(n19826), .B(n19827), .Z(n19817) );
  AND U19466 ( .A(n19828), .B(n19829), .Z(n19827) );
  XOR U19467 ( .A(n19826), .B(n19011), .Z(n19829) );
  XNOR U19468 ( .A(p_input[5700]), .B(n19830), .Z(n19011) );
  AND U19469 ( .A(n327), .B(n19831), .Z(n19830) );
  XOR U19470 ( .A(p_input[5732]), .B(p_input[5700]), .Z(n19831) );
  XNOR U19471 ( .A(n19008), .B(n19826), .Z(n19828) );
  XOR U19472 ( .A(n19832), .B(n19833), .Z(n19008) );
  AND U19473 ( .A(n324), .B(n19834), .Z(n19833) );
  XOR U19474 ( .A(p_input[5668]), .B(p_input[5636]), .Z(n19834) );
  XOR U19475 ( .A(n19835), .B(n19836), .Z(n19826) );
  AND U19476 ( .A(n19837), .B(n19838), .Z(n19836) );
  XOR U19477 ( .A(n19835), .B(n19023), .Z(n19838) );
  XNOR U19478 ( .A(p_input[5699]), .B(n19839), .Z(n19023) );
  AND U19479 ( .A(n327), .B(n19840), .Z(n19839) );
  XOR U19480 ( .A(p_input[5731]), .B(p_input[5699]), .Z(n19840) );
  XNOR U19481 ( .A(n19020), .B(n19835), .Z(n19837) );
  XOR U19482 ( .A(n19841), .B(n19842), .Z(n19020) );
  AND U19483 ( .A(n324), .B(n19843), .Z(n19842) );
  XOR U19484 ( .A(p_input[5667]), .B(p_input[5635]), .Z(n19843) );
  XOR U19485 ( .A(n19844), .B(n19845), .Z(n19835) );
  AND U19486 ( .A(n19846), .B(n19847), .Z(n19845) );
  XOR U19487 ( .A(n19844), .B(n19035), .Z(n19847) );
  XNOR U19488 ( .A(p_input[5698]), .B(n19848), .Z(n19035) );
  AND U19489 ( .A(n327), .B(n19849), .Z(n19848) );
  XOR U19490 ( .A(p_input[5730]), .B(p_input[5698]), .Z(n19849) );
  XNOR U19491 ( .A(n19032), .B(n19844), .Z(n19846) );
  XOR U19492 ( .A(n19850), .B(n19851), .Z(n19032) );
  AND U19493 ( .A(n324), .B(n19852), .Z(n19851) );
  XOR U19494 ( .A(p_input[5666]), .B(p_input[5634]), .Z(n19852) );
  XOR U19495 ( .A(n19853), .B(n19854), .Z(n19844) );
  AND U19496 ( .A(n19855), .B(n19856), .Z(n19854) );
  XNOR U19497 ( .A(n19857), .B(n19048), .Z(n19856) );
  XNOR U19498 ( .A(p_input[5697]), .B(n19858), .Z(n19048) );
  AND U19499 ( .A(n327), .B(n19859), .Z(n19858) );
  XNOR U19500 ( .A(p_input[5729]), .B(n19860), .Z(n19859) );
  IV U19501 ( .A(p_input[5697]), .Z(n19860) );
  XNOR U19502 ( .A(n19045), .B(n19853), .Z(n19855) );
  XNOR U19503 ( .A(p_input[5633]), .B(n19861), .Z(n19045) );
  AND U19504 ( .A(n324), .B(n19862), .Z(n19861) );
  XOR U19505 ( .A(p_input[5665]), .B(p_input[5633]), .Z(n19862) );
  IV U19506 ( .A(n19857), .Z(n19853) );
  AND U19507 ( .A(n19583), .B(n19586), .Z(n19857) );
  XOR U19508 ( .A(p_input[5696]), .B(n19863), .Z(n19586) );
  AND U19509 ( .A(n327), .B(n19864), .Z(n19863) );
  XOR U19510 ( .A(p_input[5728]), .B(p_input[5696]), .Z(n19864) );
  XOR U19511 ( .A(n19865), .B(n19866), .Z(n327) );
  AND U19512 ( .A(n19867), .B(n19868), .Z(n19866) );
  XNOR U19513 ( .A(p_input[5759]), .B(n19865), .Z(n19868) );
  XOR U19514 ( .A(n19865), .B(p_input[5727]), .Z(n19867) );
  XOR U19515 ( .A(n19869), .B(n19870), .Z(n19865) );
  AND U19516 ( .A(n19871), .B(n19872), .Z(n19870) );
  XNOR U19517 ( .A(p_input[5758]), .B(n19869), .Z(n19872) );
  XOR U19518 ( .A(n19869), .B(p_input[5726]), .Z(n19871) );
  XOR U19519 ( .A(n19873), .B(n19874), .Z(n19869) );
  AND U19520 ( .A(n19875), .B(n19876), .Z(n19874) );
  XNOR U19521 ( .A(p_input[5757]), .B(n19873), .Z(n19876) );
  XOR U19522 ( .A(n19873), .B(p_input[5725]), .Z(n19875) );
  XOR U19523 ( .A(n19877), .B(n19878), .Z(n19873) );
  AND U19524 ( .A(n19879), .B(n19880), .Z(n19878) );
  XNOR U19525 ( .A(p_input[5756]), .B(n19877), .Z(n19880) );
  XOR U19526 ( .A(n19877), .B(p_input[5724]), .Z(n19879) );
  XOR U19527 ( .A(n19881), .B(n19882), .Z(n19877) );
  AND U19528 ( .A(n19883), .B(n19884), .Z(n19882) );
  XNOR U19529 ( .A(p_input[5755]), .B(n19881), .Z(n19884) );
  XOR U19530 ( .A(n19881), .B(p_input[5723]), .Z(n19883) );
  XOR U19531 ( .A(n19885), .B(n19886), .Z(n19881) );
  AND U19532 ( .A(n19887), .B(n19888), .Z(n19886) );
  XNOR U19533 ( .A(p_input[5754]), .B(n19885), .Z(n19888) );
  XOR U19534 ( .A(n19885), .B(p_input[5722]), .Z(n19887) );
  XOR U19535 ( .A(n19889), .B(n19890), .Z(n19885) );
  AND U19536 ( .A(n19891), .B(n19892), .Z(n19890) );
  XNOR U19537 ( .A(p_input[5753]), .B(n19889), .Z(n19892) );
  XOR U19538 ( .A(n19889), .B(p_input[5721]), .Z(n19891) );
  XOR U19539 ( .A(n19893), .B(n19894), .Z(n19889) );
  AND U19540 ( .A(n19895), .B(n19896), .Z(n19894) );
  XNOR U19541 ( .A(p_input[5752]), .B(n19893), .Z(n19896) );
  XOR U19542 ( .A(n19893), .B(p_input[5720]), .Z(n19895) );
  XOR U19543 ( .A(n19897), .B(n19898), .Z(n19893) );
  AND U19544 ( .A(n19899), .B(n19900), .Z(n19898) );
  XNOR U19545 ( .A(p_input[5751]), .B(n19897), .Z(n19900) );
  XOR U19546 ( .A(n19897), .B(p_input[5719]), .Z(n19899) );
  XOR U19547 ( .A(n19901), .B(n19902), .Z(n19897) );
  AND U19548 ( .A(n19903), .B(n19904), .Z(n19902) );
  XNOR U19549 ( .A(p_input[5750]), .B(n19901), .Z(n19904) );
  XOR U19550 ( .A(n19901), .B(p_input[5718]), .Z(n19903) );
  XOR U19551 ( .A(n19905), .B(n19906), .Z(n19901) );
  AND U19552 ( .A(n19907), .B(n19908), .Z(n19906) );
  XNOR U19553 ( .A(p_input[5749]), .B(n19905), .Z(n19908) );
  XOR U19554 ( .A(n19905), .B(p_input[5717]), .Z(n19907) );
  XOR U19555 ( .A(n19909), .B(n19910), .Z(n19905) );
  AND U19556 ( .A(n19911), .B(n19912), .Z(n19910) );
  XNOR U19557 ( .A(p_input[5748]), .B(n19909), .Z(n19912) );
  XOR U19558 ( .A(n19909), .B(p_input[5716]), .Z(n19911) );
  XOR U19559 ( .A(n19913), .B(n19914), .Z(n19909) );
  AND U19560 ( .A(n19915), .B(n19916), .Z(n19914) );
  XNOR U19561 ( .A(p_input[5747]), .B(n19913), .Z(n19916) );
  XOR U19562 ( .A(n19913), .B(p_input[5715]), .Z(n19915) );
  XOR U19563 ( .A(n19917), .B(n19918), .Z(n19913) );
  AND U19564 ( .A(n19919), .B(n19920), .Z(n19918) );
  XNOR U19565 ( .A(p_input[5746]), .B(n19917), .Z(n19920) );
  XOR U19566 ( .A(n19917), .B(p_input[5714]), .Z(n19919) );
  XOR U19567 ( .A(n19921), .B(n19922), .Z(n19917) );
  AND U19568 ( .A(n19923), .B(n19924), .Z(n19922) );
  XNOR U19569 ( .A(p_input[5745]), .B(n19921), .Z(n19924) );
  XOR U19570 ( .A(n19921), .B(p_input[5713]), .Z(n19923) );
  XOR U19571 ( .A(n19925), .B(n19926), .Z(n19921) );
  AND U19572 ( .A(n19927), .B(n19928), .Z(n19926) );
  XNOR U19573 ( .A(p_input[5744]), .B(n19925), .Z(n19928) );
  XOR U19574 ( .A(n19925), .B(p_input[5712]), .Z(n19927) );
  XOR U19575 ( .A(n19929), .B(n19930), .Z(n19925) );
  AND U19576 ( .A(n19931), .B(n19932), .Z(n19930) );
  XNOR U19577 ( .A(p_input[5743]), .B(n19929), .Z(n19932) );
  XOR U19578 ( .A(n19929), .B(p_input[5711]), .Z(n19931) );
  XOR U19579 ( .A(n19933), .B(n19934), .Z(n19929) );
  AND U19580 ( .A(n19935), .B(n19936), .Z(n19934) );
  XNOR U19581 ( .A(p_input[5742]), .B(n19933), .Z(n19936) );
  XOR U19582 ( .A(n19933), .B(p_input[5710]), .Z(n19935) );
  XOR U19583 ( .A(n19937), .B(n19938), .Z(n19933) );
  AND U19584 ( .A(n19939), .B(n19940), .Z(n19938) );
  XNOR U19585 ( .A(p_input[5741]), .B(n19937), .Z(n19940) );
  XOR U19586 ( .A(n19937), .B(p_input[5709]), .Z(n19939) );
  XOR U19587 ( .A(n19941), .B(n19942), .Z(n19937) );
  AND U19588 ( .A(n19943), .B(n19944), .Z(n19942) );
  XNOR U19589 ( .A(p_input[5740]), .B(n19941), .Z(n19944) );
  XOR U19590 ( .A(n19941), .B(p_input[5708]), .Z(n19943) );
  XOR U19591 ( .A(n19945), .B(n19946), .Z(n19941) );
  AND U19592 ( .A(n19947), .B(n19948), .Z(n19946) );
  XNOR U19593 ( .A(p_input[5739]), .B(n19945), .Z(n19948) );
  XOR U19594 ( .A(n19945), .B(p_input[5707]), .Z(n19947) );
  XOR U19595 ( .A(n19949), .B(n19950), .Z(n19945) );
  AND U19596 ( .A(n19951), .B(n19952), .Z(n19950) );
  XNOR U19597 ( .A(p_input[5738]), .B(n19949), .Z(n19952) );
  XOR U19598 ( .A(n19949), .B(p_input[5706]), .Z(n19951) );
  XOR U19599 ( .A(n19953), .B(n19954), .Z(n19949) );
  AND U19600 ( .A(n19955), .B(n19956), .Z(n19954) );
  XNOR U19601 ( .A(p_input[5737]), .B(n19953), .Z(n19956) );
  XOR U19602 ( .A(n19953), .B(p_input[5705]), .Z(n19955) );
  XOR U19603 ( .A(n19957), .B(n19958), .Z(n19953) );
  AND U19604 ( .A(n19959), .B(n19960), .Z(n19958) );
  XNOR U19605 ( .A(p_input[5736]), .B(n19957), .Z(n19960) );
  XOR U19606 ( .A(n19957), .B(p_input[5704]), .Z(n19959) );
  XOR U19607 ( .A(n19961), .B(n19962), .Z(n19957) );
  AND U19608 ( .A(n19963), .B(n19964), .Z(n19962) );
  XNOR U19609 ( .A(p_input[5735]), .B(n19961), .Z(n19964) );
  XOR U19610 ( .A(n19961), .B(p_input[5703]), .Z(n19963) );
  XOR U19611 ( .A(n19965), .B(n19966), .Z(n19961) );
  AND U19612 ( .A(n19967), .B(n19968), .Z(n19966) );
  XNOR U19613 ( .A(p_input[5734]), .B(n19965), .Z(n19968) );
  XOR U19614 ( .A(n19965), .B(p_input[5702]), .Z(n19967) );
  XOR U19615 ( .A(n19969), .B(n19970), .Z(n19965) );
  AND U19616 ( .A(n19971), .B(n19972), .Z(n19970) );
  XNOR U19617 ( .A(p_input[5733]), .B(n19969), .Z(n19972) );
  XOR U19618 ( .A(n19969), .B(p_input[5701]), .Z(n19971) );
  XOR U19619 ( .A(n19973), .B(n19974), .Z(n19969) );
  AND U19620 ( .A(n19975), .B(n19976), .Z(n19974) );
  XNOR U19621 ( .A(p_input[5732]), .B(n19973), .Z(n19976) );
  XOR U19622 ( .A(n19973), .B(p_input[5700]), .Z(n19975) );
  XOR U19623 ( .A(n19977), .B(n19978), .Z(n19973) );
  AND U19624 ( .A(n19979), .B(n19980), .Z(n19978) );
  XNOR U19625 ( .A(p_input[5731]), .B(n19977), .Z(n19980) );
  XOR U19626 ( .A(n19977), .B(p_input[5699]), .Z(n19979) );
  XOR U19627 ( .A(n19981), .B(n19982), .Z(n19977) );
  AND U19628 ( .A(n19983), .B(n19984), .Z(n19982) );
  XNOR U19629 ( .A(p_input[5730]), .B(n19981), .Z(n19984) );
  XOR U19630 ( .A(n19981), .B(p_input[5698]), .Z(n19983) );
  XNOR U19631 ( .A(n19985), .B(n19986), .Z(n19981) );
  AND U19632 ( .A(n19987), .B(n19988), .Z(n19986) );
  XOR U19633 ( .A(p_input[5729]), .B(n19985), .Z(n19988) );
  XNOR U19634 ( .A(p_input[5697]), .B(n19985), .Z(n19987) );
  AND U19635 ( .A(p_input[5728]), .B(n19989), .Z(n19985) );
  IV U19636 ( .A(p_input[5696]), .Z(n19989) );
  XNOR U19637 ( .A(p_input[5632]), .B(n19990), .Z(n19583) );
  AND U19638 ( .A(n324), .B(n19991), .Z(n19990) );
  XOR U19639 ( .A(p_input[5664]), .B(p_input[5632]), .Z(n19991) );
  XOR U19640 ( .A(n19992), .B(n19993), .Z(n324) );
  AND U19641 ( .A(n19994), .B(n19995), .Z(n19993) );
  XNOR U19642 ( .A(p_input[5695]), .B(n19992), .Z(n19995) );
  XOR U19643 ( .A(n19992), .B(p_input[5663]), .Z(n19994) );
  XOR U19644 ( .A(n19996), .B(n19997), .Z(n19992) );
  AND U19645 ( .A(n19998), .B(n19999), .Z(n19997) );
  XNOR U19646 ( .A(p_input[5694]), .B(n19996), .Z(n19999) );
  XNOR U19647 ( .A(n19996), .B(n19598), .Z(n19998) );
  IV U19648 ( .A(p_input[5662]), .Z(n19598) );
  XOR U19649 ( .A(n20000), .B(n20001), .Z(n19996) );
  AND U19650 ( .A(n20002), .B(n20003), .Z(n20001) );
  XNOR U19651 ( .A(p_input[5693]), .B(n20000), .Z(n20003) );
  XNOR U19652 ( .A(n20000), .B(n19607), .Z(n20002) );
  IV U19653 ( .A(p_input[5661]), .Z(n19607) );
  XOR U19654 ( .A(n20004), .B(n20005), .Z(n20000) );
  AND U19655 ( .A(n20006), .B(n20007), .Z(n20005) );
  XNOR U19656 ( .A(p_input[5692]), .B(n20004), .Z(n20007) );
  XNOR U19657 ( .A(n20004), .B(n19616), .Z(n20006) );
  IV U19658 ( .A(p_input[5660]), .Z(n19616) );
  XOR U19659 ( .A(n20008), .B(n20009), .Z(n20004) );
  AND U19660 ( .A(n20010), .B(n20011), .Z(n20009) );
  XNOR U19661 ( .A(p_input[5691]), .B(n20008), .Z(n20011) );
  XNOR U19662 ( .A(n20008), .B(n19625), .Z(n20010) );
  IV U19663 ( .A(p_input[5659]), .Z(n19625) );
  XOR U19664 ( .A(n20012), .B(n20013), .Z(n20008) );
  AND U19665 ( .A(n20014), .B(n20015), .Z(n20013) );
  XNOR U19666 ( .A(p_input[5690]), .B(n20012), .Z(n20015) );
  XNOR U19667 ( .A(n20012), .B(n19634), .Z(n20014) );
  IV U19668 ( .A(p_input[5658]), .Z(n19634) );
  XOR U19669 ( .A(n20016), .B(n20017), .Z(n20012) );
  AND U19670 ( .A(n20018), .B(n20019), .Z(n20017) );
  XNOR U19671 ( .A(p_input[5689]), .B(n20016), .Z(n20019) );
  XNOR U19672 ( .A(n20016), .B(n19643), .Z(n20018) );
  IV U19673 ( .A(p_input[5657]), .Z(n19643) );
  XOR U19674 ( .A(n20020), .B(n20021), .Z(n20016) );
  AND U19675 ( .A(n20022), .B(n20023), .Z(n20021) );
  XNOR U19676 ( .A(p_input[5688]), .B(n20020), .Z(n20023) );
  XNOR U19677 ( .A(n20020), .B(n19652), .Z(n20022) );
  IV U19678 ( .A(p_input[5656]), .Z(n19652) );
  XOR U19679 ( .A(n20024), .B(n20025), .Z(n20020) );
  AND U19680 ( .A(n20026), .B(n20027), .Z(n20025) );
  XNOR U19681 ( .A(p_input[5687]), .B(n20024), .Z(n20027) );
  XNOR U19682 ( .A(n20024), .B(n19661), .Z(n20026) );
  IV U19683 ( .A(p_input[5655]), .Z(n19661) );
  XOR U19684 ( .A(n20028), .B(n20029), .Z(n20024) );
  AND U19685 ( .A(n20030), .B(n20031), .Z(n20029) );
  XNOR U19686 ( .A(p_input[5686]), .B(n20028), .Z(n20031) );
  XNOR U19687 ( .A(n20028), .B(n19670), .Z(n20030) );
  IV U19688 ( .A(p_input[5654]), .Z(n19670) );
  XOR U19689 ( .A(n20032), .B(n20033), .Z(n20028) );
  AND U19690 ( .A(n20034), .B(n20035), .Z(n20033) );
  XNOR U19691 ( .A(p_input[5685]), .B(n20032), .Z(n20035) );
  XNOR U19692 ( .A(n20032), .B(n19679), .Z(n20034) );
  IV U19693 ( .A(p_input[5653]), .Z(n19679) );
  XOR U19694 ( .A(n20036), .B(n20037), .Z(n20032) );
  AND U19695 ( .A(n20038), .B(n20039), .Z(n20037) );
  XNOR U19696 ( .A(p_input[5684]), .B(n20036), .Z(n20039) );
  XNOR U19697 ( .A(n20036), .B(n19688), .Z(n20038) );
  IV U19698 ( .A(p_input[5652]), .Z(n19688) );
  XOR U19699 ( .A(n20040), .B(n20041), .Z(n20036) );
  AND U19700 ( .A(n20042), .B(n20043), .Z(n20041) );
  XNOR U19701 ( .A(p_input[5683]), .B(n20040), .Z(n20043) );
  XNOR U19702 ( .A(n20040), .B(n19697), .Z(n20042) );
  IV U19703 ( .A(p_input[5651]), .Z(n19697) );
  XOR U19704 ( .A(n20044), .B(n20045), .Z(n20040) );
  AND U19705 ( .A(n20046), .B(n20047), .Z(n20045) );
  XNOR U19706 ( .A(p_input[5682]), .B(n20044), .Z(n20047) );
  XNOR U19707 ( .A(n20044), .B(n19706), .Z(n20046) );
  IV U19708 ( .A(p_input[5650]), .Z(n19706) );
  XOR U19709 ( .A(n20048), .B(n20049), .Z(n20044) );
  AND U19710 ( .A(n20050), .B(n20051), .Z(n20049) );
  XNOR U19711 ( .A(p_input[5681]), .B(n20048), .Z(n20051) );
  XNOR U19712 ( .A(n20048), .B(n19715), .Z(n20050) );
  IV U19713 ( .A(p_input[5649]), .Z(n19715) );
  XOR U19714 ( .A(n20052), .B(n20053), .Z(n20048) );
  AND U19715 ( .A(n20054), .B(n20055), .Z(n20053) );
  XNOR U19716 ( .A(p_input[5680]), .B(n20052), .Z(n20055) );
  XNOR U19717 ( .A(n20052), .B(n19724), .Z(n20054) );
  IV U19718 ( .A(p_input[5648]), .Z(n19724) );
  XOR U19719 ( .A(n20056), .B(n20057), .Z(n20052) );
  AND U19720 ( .A(n20058), .B(n20059), .Z(n20057) );
  XNOR U19721 ( .A(p_input[5679]), .B(n20056), .Z(n20059) );
  XNOR U19722 ( .A(n20056), .B(n19733), .Z(n20058) );
  IV U19723 ( .A(p_input[5647]), .Z(n19733) );
  XOR U19724 ( .A(n20060), .B(n20061), .Z(n20056) );
  AND U19725 ( .A(n20062), .B(n20063), .Z(n20061) );
  XNOR U19726 ( .A(p_input[5678]), .B(n20060), .Z(n20063) );
  XNOR U19727 ( .A(n20060), .B(n19742), .Z(n20062) );
  IV U19728 ( .A(p_input[5646]), .Z(n19742) );
  XOR U19729 ( .A(n20064), .B(n20065), .Z(n20060) );
  AND U19730 ( .A(n20066), .B(n20067), .Z(n20065) );
  XNOR U19731 ( .A(p_input[5677]), .B(n20064), .Z(n20067) );
  XNOR U19732 ( .A(n20064), .B(n19751), .Z(n20066) );
  IV U19733 ( .A(p_input[5645]), .Z(n19751) );
  XOR U19734 ( .A(n20068), .B(n20069), .Z(n20064) );
  AND U19735 ( .A(n20070), .B(n20071), .Z(n20069) );
  XNOR U19736 ( .A(p_input[5676]), .B(n20068), .Z(n20071) );
  XNOR U19737 ( .A(n20068), .B(n19760), .Z(n20070) );
  IV U19738 ( .A(p_input[5644]), .Z(n19760) );
  XOR U19739 ( .A(n20072), .B(n20073), .Z(n20068) );
  AND U19740 ( .A(n20074), .B(n20075), .Z(n20073) );
  XNOR U19741 ( .A(p_input[5675]), .B(n20072), .Z(n20075) );
  XNOR U19742 ( .A(n20072), .B(n19769), .Z(n20074) );
  IV U19743 ( .A(p_input[5643]), .Z(n19769) );
  XOR U19744 ( .A(n20076), .B(n20077), .Z(n20072) );
  AND U19745 ( .A(n20078), .B(n20079), .Z(n20077) );
  XNOR U19746 ( .A(p_input[5674]), .B(n20076), .Z(n20079) );
  XNOR U19747 ( .A(n20076), .B(n19778), .Z(n20078) );
  IV U19748 ( .A(p_input[5642]), .Z(n19778) );
  XOR U19749 ( .A(n20080), .B(n20081), .Z(n20076) );
  AND U19750 ( .A(n20082), .B(n20083), .Z(n20081) );
  XNOR U19751 ( .A(p_input[5673]), .B(n20080), .Z(n20083) );
  XNOR U19752 ( .A(n20080), .B(n19787), .Z(n20082) );
  IV U19753 ( .A(p_input[5641]), .Z(n19787) );
  XOR U19754 ( .A(n20084), .B(n20085), .Z(n20080) );
  AND U19755 ( .A(n20086), .B(n20087), .Z(n20085) );
  XNOR U19756 ( .A(p_input[5672]), .B(n20084), .Z(n20087) );
  XNOR U19757 ( .A(n20084), .B(n19796), .Z(n20086) );
  IV U19758 ( .A(p_input[5640]), .Z(n19796) );
  XOR U19759 ( .A(n20088), .B(n20089), .Z(n20084) );
  AND U19760 ( .A(n20090), .B(n20091), .Z(n20089) );
  XNOR U19761 ( .A(p_input[5671]), .B(n20088), .Z(n20091) );
  XNOR U19762 ( .A(n20088), .B(n19805), .Z(n20090) );
  IV U19763 ( .A(p_input[5639]), .Z(n19805) );
  XOR U19764 ( .A(n20092), .B(n20093), .Z(n20088) );
  AND U19765 ( .A(n20094), .B(n20095), .Z(n20093) );
  XNOR U19766 ( .A(p_input[5670]), .B(n20092), .Z(n20095) );
  XNOR U19767 ( .A(n20092), .B(n19814), .Z(n20094) );
  IV U19768 ( .A(p_input[5638]), .Z(n19814) );
  XOR U19769 ( .A(n20096), .B(n20097), .Z(n20092) );
  AND U19770 ( .A(n20098), .B(n20099), .Z(n20097) );
  XNOR U19771 ( .A(p_input[5669]), .B(n20096), .Z(n20099) );
  XNOR U19772 ( .A(n20096), .B(n19823), .Z(n20098) );
  IV U19773 ( .A(p_input[5637]), .Z(n19823) );
  XOR U19774 ( .A(n20100), .B(n20101), .Z(n20096) );
  AND U19775 ( .A(n20102), .B(n20103), .Z(n20101) );
  XNOR U19776 ( .A(p_input[5668]), .B(n20100), .Z(n20103) );
  XNOR U19777 ( .A(n20100), .B(n19832), .Z(n20102) );
  IV U19778 ( .A(p_input[5636]), .Z(n19832) );
  XOR U19779 ( .A(n20104), .B(n20105), .Z(n20100) );
  AND U19780 ( .A(n20106), .B(n20107), .Z(n20105) );
  XNOR U19781 ( .A(p_input[5667]), .B(n20104), .Z(n20107) );
  XNOR U19782 ( .A(n20104), .B(n19841), .Z(n20106) );
  IV U19783 ( .A(p_input[5635]), .Z(n19841) );
  XOR U19784 ( .A(n20108), .B(n20109), .Z(n20104) );
  AND U19785 ( .A(n20110), .B(n20111), .Z(n20109) );
  XNOR U19786 ( .A(p_input[5666]), .B(n20108), .Z(n20111) );
  XNOR U19787 ( .A(n20108), .B(n19850), .Z(n20110) );
  IV U19788 ( .A(p_input[5634]), .Z(n19850) );
  XNOR U19789 ( .A(n20112), .B(n20113), .Z(n20108) );
  AND U19790 ( .A(n20114), .B(n20115), .Z(n20113) );
  XOR U19791 ( .A(p_input[5665]), .B(n20112), .Z(n20115) );
  XNOR U19792 ( .A(p_input[5633]), .B(n20112), .Z(n20114) );
  AND U19793 ( .A(p_input[5664]), .B(n20116), .Z(n20112) );
  IV U19794 ( .A(p_input[5632]), .Z(n20116) );
  XOR U19795 ( .A(n20117), .B(n20118), .Z(n16473) );
  AND U19796 ( .A(n1009), .B(n20119), .Z(n20118) );
  XNOR U19797 ( .A(n20120), .B(n20117), .Z(n20119) );
  XOR U19798 ( .A(n20121), .B(n20122), .Z(n1009) );
  AND U19799 ( .A(n20123), .B(n20124), .Z(n20122) );
  XOR U19800 ( .A(n20121), .B(n16488), .Z(n20124) );
  XOR U19801 ( .A(n20125), .B(n20126), .Z(n16488) );
  AND U19802 ( .A(n847), .B(n20127), .Z(n20126) );
  XOR U19803 ( .A(n20128), .B(n20125), .Z(n20127) );
  XNOR U19804 ( .A(n16485), .B(n20121), .Z(n20123) );
  XOR U19805 ( .A(n20129), .B(n20130), .Z(n16485) );
  AND U19806 ( .A(n844), .B(n20131), .Z(n20130) );
  XOR U19807 ( .A(n20132), .B(n20129), .Z(n20131) );
  XOR U19808 ( .A(n20133), .B(n20134), .Z(n20121) );
  AND U19809 ( .A(n20135), .B(n20136), .Z(n20134) );
  XOR U19810 ( .A(n20133), .B(n16500), .Z(n20136) );
  XOR U19811 ( .A(n20137), .B(n20138), .Z(n16500) );
  AND U19812 ( .A(n847), .B(n20139), .Z(n20138) );
  XOR U19813 ( .A(n20140), .B(n20137), .Z(n20139) );
  XNOR U19814 ( .A(n16497), .B(n20133), .Z(n20135) );
  XOR U19815 ( .A(n20141), .B(n20142), .Z(n16497) );
  AND U19816 ( .A(n844), .B(n20143), .Z(n20142) );
  XOR U19817 ( .A(n20144), .B(n20141), .Z(n20143) );
  XOR U19818 ( .A(n20145), .B(n20146), .Z(n20133) );
  AND U19819 ( .A(n20147), .B(n20148), .Z(n20146) );
  XOR U19820 ( .A(n20145), .B(n16512), .Z(n20148) );
  XOR U19821 ( .A(n20149), .B(n20150), .Z(n16512) );
  AND U19822 ( .A(n847), .B(n20151), .Z(n20150) );
  XOR U19823 ( .A(n20152), .B(n20149), .Z(n20151) );
  XNOR U19824 ( .A(n16509), .B(n20145), .Z(n20147) );
  XOR U19825 ( .A(n20153), .B(n20154), .Z(n16509) );
  AND U19826 ( .A(n844), .B(n20155), .Z(n20154) );
  XOR U19827 ( .A(n20156), .B(n20153), .Z(n20155) );
  XOR U19828 ( .A(n20157), .B(n20158), .Z(n20145) );
  AND U19829 ( .A(n20159), .B(n20160), .Z(n20158) );
  XOR U19830 ( .A(n20157), .B(n16524), .Z(n20160) );
  XOR U19831 ( .A(n20161), .B(n20162), .Z(n16524) );
  AND U19832 ( .A(n847), .B(n20163), .Z(n20162) );
  XOR U19833 ( .A(n20164), .B(n20161), .Z(n20163) );
  XNOR U19834 ( .A(n16521), .B(n20157), .Z(n20159) );
  XOR U19835 ( .A(n20165), .B(n20166), .Z(n16521) );
  AND U19836 ( .A(n844), .B(n20167), .Z(n20166) );
  XOR U19837 ( .A(n20168), .B(n20165), .Z(n20167) );
  XOR U19838 ( .A(n20169), .B(n20170), .Z(n20157) );
  AND U19839 ( .A(n20171), .B(n20172), .Z(n20170) );
  XOR U19840 ( .A(n20169), .B(n16536), .Z(n20172) );
  XOR U19841 ( .A(n20173), .B(n20174), .Z(n16536) );
  AND U19842 ( .A(n847), .B(n20175), .Z(n20174) );
  XOR U19843 ( .A(n20176), .B(n20173), .Z(n20175) );
  XNOR U19844 ( .A(n16533), .B(n20169), .Z(n20171) );
  XOR U19845 ( .A(n20177), .B(n20178), .Z(n16533) );
  AND U19846 ( .A(n844), .B(n20179), .Z(n20178) );
  XOR U19847 ( .A(n20180), .B(n20177), .Z(n20179) );
  XOR U19848 ( .A(n20181), .B(n20182), .Z(n20169) );
  AND U19849 ( .A(n20183), .B(n20184), .Z(n20182) );
  XOR U19850 ( .A(n20181), .B(n16548), .Z(n20184) );
  XOR U19851 ( .A(n20185), .B(n20186), .Z(n16548) );
  AND U19852 ( .A(n847), .B(n20187), .Z(n20186) );
  XOR U19853 ( .A(n20188), .B(n20185), .Z(n20187) );
  XNOR U19854 ( .A(n16545), .B(n20181), .Z(n20183) );
  XOR U19855 ( .A(n20189), .B(n20190), .Z(n16545) );
  AND U19856 ( .A(n844), .B(n20191), .Z(n20190) );
  XOR U19857 ( .A(n20192), .B(n20189), .Z(n20191) );
  XOR U19858 ( .A(n20193), .B(n20194), .Z(n20181) );
  AND U19859 ( .A(n20195), .B(n20196), .Z(n20194) );
  XOR U19860 ( .A(n20193), .B(n16560), .Z(n20196) );
  XOR U19861 ( .A(n20197), .B(n20198), .Z(n16560) );
  AND U19862 ( .A(n847), .B(n20199), .Z(n20198) );
  XOR U19863 ( .A(n20200), .B(n20197), .Z(n20199) );
  XNOR U19864 ( .A(n16557), .B(n20193), .Z(n20195) );
  XOR U19865 ( .A(n20201), .B(n20202), .Z(n16557) );
  AND U19866 ( .A(n844), .B(n20203), .Z(n20202) );
  XOR U19867 ( .A(n20204), .B(n20201), .Z(n20203) );
  XOR U19868 ( .A(n20205), .B(n20206), .Z(n20193) );
  AND U19869 ( .A(n20207), .B(n20208), .Z(n20206) );
  XOR U19870 ( .A(n20205), .B(n16572), .Z(n20208) );
  XOR U19871 ( .A(n20209), .B(n20210), .Z(n16572) );
  AND U19872 ( .A(n847), .B(n20211), .Z(n20210) );
  XOR U19873 ( .A(n20212), .B(n20209), .Z(n20211) );
  XNOR U19874 ( .A(n16569), .B(n20205), .Z(n20207) );
  XOR U19875 ( .A(n20213), .B(n20214), .Z(n16569) );
  AND U19876 ( .A(n844), .B(n20215), .Z(n20214) );
  XOR U19877 ( .A(n20216), .B(n20213), .Z(n20215) );
  XOR U19878 ( .A(n20217), .B(n20218), .Z(n20205) );
  AND U19879 ( .A(n20219), .B(n20220), .Z(n20218) );
  XOR U19880 ( .A(n20217), .B(n16584), .Z(n20220) );
  XOR U19881 ( .A(n20221), .B(n20222), .Z(n16584) );
  AND U19882 ( .A(n847), .B(n20223), .Z(n20222) );
  XOR U19883 ( .A(n20224), .B(n20221), .Z(n20223) );
  XNOR U19884 ( .A(n16581), .B(n20217), .Z(n20219) );
  XOR U19885 ( .A(n20225), .B(n20226), .Z(n16581) );
  AND U19886 ( .A(n844), .B(n20227), .Z(n20226) );
  XOR U19887 ( .A(n20228), .B(n20225), .Z(n20227) );
  XOR U19888 ( .A(n20229), .B(n20230), .Z(n20217) );
  AND U19889 ( .A(n20231), .B(n20232), .Z(n20230) );
  XOR U19890 ( .A(n20229), .B(n16596), .Z(n20232) );
  XOR U19891 ( .A(n20233), .B(n20234), .Z(n16596) );
  AND U19892 ( .A(n847), .B(n20235), .Z(n20234) );
  XOR U19893 ( .A(n20236), .B(n20233), .Z(n20235) );
  XNOR U19894 ( .A(n16593), .B(n20229), .Z(n20231) );
  XOR U19895 ( .A(n20237), .B(n20238), .Z(n16593) );
  AND U19896 ( .A(n844), .B(n20239), .Z(n20238) );
  XOR U19897 ( .A(n20240), .B(n20237), .Z(n20239) );
  XOR U19898 ( .A(n20241), .B(n20242), .Z(n20229) );
  AND U19899 ( .A(n20243), .B(n20244), .Z(n20242) );
  XOR U19900 ( .A(n20241), .B(n16608), .Z(n20244) );
  XOR U19901 ( .A(n20245), .B(n20246), .Z(n16608) );
  AND U19902 ( .A(n847), .B(n20247), .Z(n20246) );
  XOR U19903 ( .A(n20248), .B(n20245), .Z(n20247) );
  XNOR U19904 ( .A(n16605), .B(n20241), .Z(n20243) );
  XOR U19905 ( .A(n20249), .B(n20250), .Z(n16605) );
  AND U19906 ( .A(n844), .B(n20251), .Z(n20250) );
  XOR U19907 ( .A(n20252), .B(n20249), .Z(n20251) );
  XOR U19908 ( .A(n20253), .B(n20254), .Z(n20241) );
  AND U19909 ( .A(n20255), .B(n20256), .Z(n20254) );
  XOR U19910 ( .A(n20253), .B(n16620), .Z(n20256) );
  XOR U19911 ( .A(n20257), .B(n20258), .Z(n16620) );
  AND U19912 ( .A(n847), .B(n20259), .Z(n20258) );
  XOR U19913 ( .A(n20260), .B(n20257), .Z(n20259) );
  XNOR U19914 ( .A(n16617), .B(n20253), .Z(n20255) );
  XOR U19915 ( .A(n20261), .B(n20262), .Z(n16617) );
  AND U19916 ( .A(n844), .B(n20263), .Z(n20262) );
  XOR U19917 ( .A(n20264), .B(n20261), .Z(n20263) );
  XOR U19918 ( .A(n20265), .B(n20266), .Z(n20253) );
  AND U19919 ( .A(n20267), .B(n20268), .Z(n20266) );
  XOR U19920 ( .A(n20265), .B(n16632), .Z(n20268) );
  XOR U19921 ( .A(n20269), .B(n20270), .Z(n16632) );
  AND U19922 ( .A(n847), .B(n20271), .Z(n20270) );
  XOR U19923 ( .A(n20272), .B(n20269), .Z(n20271) );
  XNOR U19924 ( .A(n16629), .B(n20265), .Z(n20267) );
  XOR U19925 ( .A(n20273), .B(n20274), .Z(n16629) );
  AND U19926 ( .A(n844), .B(n20275), .Z(n20274) );
  XOR U19927 ( .A(n20276), .B(n20273), .Z(n20275) );
  XOR U19928 ( .A(n20277), .B(n20278), .Z(n20265) );
  AND U19929 ( .A(n20279), .B(n20280), .Z(n20278) );
  XOR U19930 ( .A(n20277), .B(n16644), .Z(n20280) );
  XOR U19931 ( .A(n20281), .B(n20282), .Z(n16644) );
  AND U19932 ( .A(n847), .B(n20283), .Z(n20282) );
  XOR U19933 ( .A(n20284), .B(n20281), .Z(n20283) );
  XNOR U19934 ( .A(n16641), .B(n20277), .Z(n20279) );
  XOR U19935 ( .A(n20285), .B(n20286), .Z(n16641) );
  AND U19936 ( .A(n844), .B(n20287), .Z(n20286) );
  XOR U19937 ( .A(n20288), .B(n20285), .Z(n20287) );
  XOR U19938 ( .A(n20289), .B(n20290), .Z(n20277) );
  AND U19939 ( .A(n20291), .B(n20292), .Z(n20290) );
  XOR U19940 ( .A(n20289), .B(n16656), .Z(n20292) );
  XOR U19941 ( .A(n20293), .B(n20294), .Z(n16656) );
  AND U19942 ( .A(n847), .B(n20295), .Z(n20294) );
  XOR U19943 ( .A(n20296), .B(n20293), .Z(n20295) );
  XNOR U19944 ( .A(n16653), .B(n20289), .Z(n20291) );
  XOR U19945 ( .A(n20297), .B(n20298), .Z(n16653) );
  AND U19946 ( .A(n844), .B(n20299), .Z(n20298) );
  XOR U19947 ( .A(n20300), .B(n20297), .Z(n20299) );
  XOR U19948 ( .A(n20301), .B(n20302), .Z(n20289) );
  AND U19949 ( .A(n20303), .B(n20304), .Z(n20302) );
  XOR U19950 ( .A(n20301), .B(n16668), .Z(n20304) );
  XOR U19951 ( .A(n20305), .B(n20306), .Z(n16668) );
  AND U19952 ( .A(n847), .B(n20307), .Z(n20306) );
  XOR U19953 ( .A(n20308), .B(n20305), .Z(n20307) );
  XNOR U19954 ( .A(n16665), .B(n20301), .Z(n20303) );
  XOR U19955 ( .A(n20309), .B(n20310), .Z(n16665) );
  AND U19956 ( .A(n844), .B(n20311), .Z(n20310) );
  XOR U19957 ( .A(n20312), .B(n20309), .Z(n20311) );
  XOR U19958 ( .A(n20313), .B(n20314), .Z(n20301) );
  AND U19959 ( .A(n20315), .B(n20316), .Z(n20314) );
  XOR U19960 ( .A(n20313), .B(n16680), .Z(n20316) );
  XOR U19961 ( .A(n20317), .B(n20318), .Z(n16680) );
  AND U19962 ( .A(n847), .B(n20319), .Z(n20318) );
  XOR U19963 ( .A(n20320), .B(n20317), .Z(n20319) );
  XNOR U19964 ( .A(n16677), .B(n20313), .Z(n20315) );
  XOR U19965 ( .A(n20321), .B(n20322), .Z(n16677) );
  AND U19966 ( .A(n844), .B(n20323), .Z(n20322) );
  XOR U19967 ( .A(n20324), .B(n20321), .Z(n20323) );
  XOR U19968 ( .A(n20325), .B(n20326), .Z(n20313) );
  AND U19969 ( .A(n20327), .B(n20328), .Z(n20326) );
  XOR U19970 ( .A(n20325), .B(n16692), .Z(n20328) );
  XOR U19971 ( .A(n20329), .B(n20330), .Z(n16692) );
  AND U19972 ( .A(n847), .B(n20331), .Z(n20330) );
  XOR U19973 ( .A(n20332), .B(n20329), .Z(n20331) );
  XNOR U19974 ( .A(n16689), .B(n20325), .Z(n20327) );
  XOR U19975 ( .A(n20333), .B(n20334), .Z(n16689) );
  AND U19976 ( .A(n844), .B(n20335), .Z(n20334) );
  XOR U19977 ( .A(n20336), .B(n20333), .Z(n20335) );
  XOR U19978 ( .A(n20337), .B(n20338), .Z(n20325) );
  AND U19979 ( .A(n20339), .B(n20340), .Z(n20338) );
  XOR U19980 ( .A(n20337), .B(n16704), .Z(n20340) );
  XOR U19981 ( .A(n20341), .B(n20342), .Z(n16704) );
  AND U19982 ( .A(n847), .B(n20343), .Z(n20342) );
  XOR U19983 ( .A(n20344), .B(n20341), .Z(n20343) );
  XNOR U19984 ( .A(n16701), .B(n20337), .Z(n20339) );
  XOR U19985 ( .A(n20345), .B(n20346), .Z(n16701) );
  AND U19986 ( .A(n844), .B(n20347), .Z(n20346) );
  XOR U19987 ( .A(n20348), .B(n20345), .Z(n20347) );
  XOR U19988 ( .A(n20349), .B(n20350), .Z(n20337) );
  AND U19989 ( .A(n20351), .B(n20352), .Z(n20350) );
  XOR U19990 ( .A(n20349), .B(n16716), .Z(n20352) );
  XOR U19991 ( .A(n20353), .B(n20354), .Z(n16716) );
  AND U19992 ( .A(n847), .B(n20355), .Z(n20354) );
  XOR U19993 ( .A(n20356), .B(n20353), .Z(n20355) );
  XNOR U19994 ( .A(n16713), .B(n20349), .Z(n20351) );
  XOR U19995 ( .A(n20357), .B(n20358), .Z(n16713) );
  AND U19996 ( .A(n844), .B(n20359), .Z(n20358) );
  XOR U19997 ( .A(n20360), .B(n20357), .Z(n20359) );
  XOR U19998 ( .A(n20361), .B(n20362), .Z(n20349) );
  AND U19999 ( .A(n20363), .B(n20364), .Z(n20362) );
  XOR U20000 ( .A(n20361), .B(n16728), .Z(n20364) );
  XOR U20001 ( .A(n20365), .B(n20366), .Z(n16728) );
  AND U20002 ( .A(n847), .B(n20367), .Z(n20366) );
  XOR U20003 ( .A(n20368), .B(n20365), .Z(n20367) );
  XNOR U20004 ( .A(n16725), .B(n20361), .Z(n20363) );
  XOR U20005 ( .A(n20369), .B(n20370), .Z(n16725) );
  AND U20006 ( .A(n844), .B(n20371), .Z(n20370) );
  XOR U20007 ( .A(n20372), .B(n20369), .Z(n20371) );
  XOR U20008 ( .A(n20373), .B(n20374), .Z(n20361) );
  AND U20009 ( .A(n20375), .B(n20376), .Z(n20374) );
  XOR U20010 ( .A(n20373), .B(n16740), .Z(n20376) );
  XOR U20011 ( .A(n20377), .B(n20378), .Z(n16740) );
  AND U20012 ( .A(n847), .B(n20379), .Z(n20378) );
  XOR U20013 ( .A(n20380), .B(n20377), .Z(n20379) );
  XNOR U20014 ( .A(n16737), .B(n20373), .Z(n20375) );
  XOR U20015 ( .A(n20381), .B(n20382), .Z(n16737) );
  AND U20016 ( .A(n844), .B(n20383), .Z(n20382) );
  XOR U20017 ( .A(n20384), .B(n20381), .Z(n20383) );
  XOR U20018 ( .A(n20385), .B(n20386), .Z(n20373) );
  AND U20019 ( .A(n20387), .B(n20388), .Z(n20386) );
  XOR U20020 ( .A(n20385), .B(n16752), .Z(n20388) );
  XOR U20021 ( .A(n20389), .B(n20390), .Z(n16752) );
  AND U20022 ( .A(n847), .B(n20391), .Z(n20390) );
  XOR U20023 ( .A(n20392), .B(n20389), .Z(n20391) );
  XNOR U20024 ( .A(n16749), .B(n20385), .Z(n20387) );
  XOR U20025 ( .A(n20393), .B(n20394), .Z(n16749) );
  AND U20026 ( .A(n844), .B(n20395), .Z(n20394) );
  XOR U20027 ( .A(n20396), .B(n20393), .Z(n20395) );
  XOR U20028 ( .A(n20397), .B(n20398), .Z(n20385) );
  AND U20029 ( .A(n20399), .B(n20400), .Z(n20398) );
  XOR U20030 ( .A(n20397), .B(n16764), .Z(n20400) );
  XOR U20031 ( .A(n20401), .B(n20402), .Z(n16764) );
  AND U20032 ( .A(n847), .B(n20403), .Z(n20402) );
  XOR U20033 ( .A(n20404), .B(n20401), .Z(n20403) );
  XNOR U20034 ( .A(n16761), .B(n20397), .Z(n20399) );
  XOR U20035 ( .A(n20405), .B(n20406), .Z(n16761) );
  AND U20036 ( .A(n844), .B(n20407), .Z(n20406) );
  XOR U20037 ( .A(n20408), .B(n20405), .Z(n20407) );
  XOR U20038 ( .A(n20409), .B(n20410), .Z(n20397) );
  AND U20039 ( .A(n20411), .B(n20412), .Z(n20410) );
  XOR U20040 ( .A(n20409), .B(n16776), .Z(n20412) );
  XOR U20041 ( .A(n20413), .B(n20414), .Z(n16776) );
  AND U20042 ( .A(n847), .B(n20415), .Z(n20414) );
  XOR U20043 ( .A(n20416), .B(n20413), .Z(n20415) );
  XNOR U20044 ( .A(n16773), .B(n20409), .Z(n20411) );
  XOR U20045 ( .A(n20417), .B(n20418), .Z(n16773) );
  AND U20046 ( .A(n844), .B(n20419), .Z(n20418) );
  XOR U20047 ( .A(n20420), .B(n20417), .Z(n20419) );
  XOR U20048 ( .A(n20421), .B(n20422), .Z(n20409) );
  AND U20049 ( .A(n20423), .B(n20424), .Z(n20422) );
  XOR U20050 ( .A(n20421), .B(n16788), .Z(n20424) );
  XOR U20051 ( .A(n20425), .B(n20426), .Z(n16788) );
  AND U20052 ( .A(n847), .B(n20427), .Z(n20426) );
  XOR U20053 ( .A(n20428), .B(n20425), .Z(n20427) );
  XNOR U20054 ( .A(n16785), .B(n20421), .Z(n20423) );
  XOR U20055 ( .A(n20429), .B(n20430), .Z(n16785) );
  AND U20056 ( .A(n844), .B(n20431), .Z(n20430) );
  XOR U20057 ( .A(n20432), .B(n20429), .Z(n20431) );
  XOR U20058 ( .A(n20433), .B(n20434), .Z(n20421) );
  AND U20059 ( .A(n20435), .B(n20436), .Z(n20434) );
  XOR U20060 ( .A(n20433), .B(n16800), .Z(n20436) );
  XOR U20061 ( .A(n20437), .B(n20438), .Z(n16800) );
  AND U20062 ( .A(n847), .B(n20439), .Z(n20438) );
  XOR U20063 ( .A(n20440), .B(n20437), .Z(n20439) );
  XNOR U20064 ( .A(n16797), .B(n20433), .Z(n20435) );
  XOR U20065 ( .A(n20441), .B(n20442), .Z(n16797) );
  AND U20066 ( .A(n844), .B(n20443), .Z(n20442) );
  XOR U20067 ( .A(n20444), .B(n20441), .Z(n20443) );
  XOR U20068 ( .A(n20445), .B(n20446), .Z(n20433) );
  AND U20069 ( .A(n20447), .B(n20448), .Z(n20446) );
  XOR U20070 ( .A(n20445), .B(n16812), .Z(n20448) );
  XOR U20071 ( .A(n20449), .B(n20450), .Z(n16812) );
  AND U20072 ( .A(n847), .B(n20451), .Z(n20450) );
  XOR U20073 ( .A(n20452), .B(n20449), .Z(n20451) );
  XNOR U20074 ( .A(n16809), .B(n20445), .Z(n20447) );
  XOR U20075 ( .A(n20453), .B(n20454), .Z(n16809) );
  AND U20076 ( .A(n844), .B(n20455), .Z(n20454) );
  XOR U20077 ( .A(n20456), .B(n20453), .Z(n20455) );
  XOR U20078 ( .A(n20457), .B(n20458), .Z(n20445) );
  AND U20079 ( .A(n20459), .B(n20460), .Z(n20458) );
  XOR U20080 ( .A(n20457), .B(n16824), .Z(n20460) );
  XOR U20081 ( .A(n20461), .B(n20462), .Z(n16824) );
  AND U20082 ( .A(n847), .B(n20463), .Z(n20462) );
  XOR U20083 ( .A(n20464), .B(n20461), .Z(n20463) );
  XNOR U20084 ( .A(n16821), .B(n20457), .Z(n20459) );
  XOR U20085 ( .A(n20465), .B(n20466), .Z(n16821) );
  AND U20086 ( .A(n844), .B(n20467), .Z(n20466) );
  XOR U20087 ( .A(n20468), .B(n20465), .Z(n20467) );
  XOR U20088 ( .A(n20469), .B(n20470), .Z(n20457) );
  AND U20089 ( .A(n20471), .B(n20472), .Z(n20470) );
  XOR U20090 ( .A(n20469), .B(n16836), .Z(n20472) );
  XOR U20091 ( .A(n20473), .B(n20474), .Z(n16836) );
  AND U20092 ( .A(n847), .B(n20475), .Z(n20474) );
  XOR U20093 ( .A(n20476), .B(n20473), .Z(n20475) );
  XNOR U20094 ( .A(n16833), .B(n20469), .Z(n20471) );
  XOR U20095 ( .A(n20477), .B(n20478), .Z(n16833) );
  AND U20096 ( .A(n844), .B(n20479), .Z(n20478) );
  XOR U20097 ( .A(n20480), .B(n20477), .Z(n20479) );
  XOR U20098 ( .A(n20481), .B(n20482), .Z(n20469) );
  AND U20099 ( .A(n20483), .B(n20484), .Z(n20482) );
  XNOR U20100 ( .A(n20485), .B(n16849), .Z(n20484) );
  XOR U20101 ( .A(n20486), .B(n20487), .Z(n16849) );
  AND U20102 ( .A(n847), .B(n20488), .Z(n20487) );
  XOR U20103 ( .A(n20486), .B(n20489), .Z(n20488) );
  XNOR U20104 ( .A(n16846), .B(n20481), .Z(n20483) );
  XOR U20105 ( .A(n20490), .B(n20491), .Z(n16846) );
  AND U20106 ( .A(n844), .B(n20492), .Z(n20491) );
  XOR U20107 ( .A(n20490), .B(n20493), .Z(n20492) );
  IV U20108 ( .A(n20485), .Z(n20481) );
  AND U20109 ( .A(n20117), .B(n20120), .Z(n20485) );
  XNOR U20110 ( .A(n20494), .B(n20495), .Z(n20120) );
  AND U20111 ( .A(n847), .B(n20496), .Z(n20495) );
  XNOR U20112 ( .A(n20497), .B(n20494), .Z(n20496) );
  XOR U20113 ( .A(n20498), .B(n20499), .Z(n847) );
  AND U20114 ( .A(n20500), .B(n20501), .Z(n20499) );
  XOR U20115 ( .A(n20498), .B(n20128), .Z(n20501) );
  XNOR U20116 ( .A(n20502), .B(n20503), .Z(n20128) );
  AND U20117 ( .A(n20504), .B(n511), .Z(n20503) );
  AND U20118 ( .A(n20502), .B(n20505), .Z(n20504) );
  XNOR U20119 ( .A(n20125), .B(n20498), .Z(n20500) );
  XOR U20120 ( .A(n20506), .B(n20507), .Z(n20125) );
  AND U20121 ( .A(n20508), .B(n509), .Z(n20507) );
  NOR U20122 ( .A(n20506), .B(n20509), .Z(n20508) );
  XOR U20123 ( .A(n20510), .B(n20511), .Z(n20498) );
  AND U20124 ( .A(n20512), .B(n20513), .Z(n20511) );
  XOR U20125 ( .A(n20510), .B(n20140), .Z(n20513) );
  XOR U20126 ( .A(n20514), .B(n20515), .Z(n20140) );
  AND U20127 ( .A(n511), .B(n20516), .Z(n20515) );
  XOR U20128 ( .A(n20517), .B(n20514), .Z(n20516) );
  XNOR U20129 ( .A(n20137), .B(n20510), .Z(n20512) );
  XOR U20130 ( .A(n20518), .B(n20519), .Z(n20137) );
  AND U20131 ( .A(n509), .B(n20520), .Z(n20519) );
  XOR U20132 ( .A(n20521), .B(n20518), .Z(n20520) );
  XOR U20133 ( .A(n20522), .B(n20523), .Z(n20510) );
  AND U20134 ( .A(n20524), .B(n20525), .Z(n20523) );
  XOR U20135 ( .A(n20522), .B(n20152), .Z(n20525) );
  XOR U20136 ( .A(n20526), .B(n20527), .Z(n20152) );
  AND U20137 ( .A(n511), .B(n20528), .Z(n20527) );
  XOR U20138 ( .A(n20529), .B(n20526), .Z(n20528) );
  XNOR U20139 ( .A(n20149), .B(n20522), .Z(n20524) );
  XOR U20140 ( .A(n20530), .B(n20531), .Z(n20149) );
  AND U20141 ( .A(n509), .B(n20532), .Z(n20531) );
  XOR U20142 ( .A(n20533), .B(n20530), .Z(n20532) );
  XOR U20143 ( .A(n20534), .B(n20535), .Z(n20522) );
  AND U20144 ( .A(n20536), .B(n20537), .Z(n20535) );
  XOR U20145 ( .A(n20534), .B(n20164), .Z(n20537) );
  XOR U20146 ( .A(n20538), .B(n20539), .Z(n20164) );
  AND U20147 ( .A(n511), .B(n20540), .Z(n20539) );
  XOR U20148 ( .A(n20541), .B(n20538), .Z(n20540) );
  XNOR U20149 ( .A(n20161), .B(n20534), .Z(n20536) );
  XOR U20150 ( .A(n20542), .B(n20543), .Z(n20161) );
  AND U20151 ( .A(n509), .B(n20544), .Z(n20543) );
  XOR U20152 ( .A(n20545), .B(n20542), .Z(n20544) );
  XOR U20153 ( .A(n20546), .B(n20547), .Z(n20534) );
  AND U20154 ( .A(n20548), .B(n20549), .Z(n20547) );
  XOR U20155 ( .A(n20546), .B(n20176), .Z(n20549) );
  XOR U20156 ( .A(n20550), .B(n20551), .Z(n20176) );
  AND U20157 ( .A(n511), .B(n20552), .Z(n20551) );
  XOR U20158 ( .A(n20553), .B(n20550), .Z(n20552) );
  XNOR U20159 ( .A(n20173), .B(n20546), .Z(n20548) );
  XOR U20160 ( .A(n20554), .B(n20555), .Z(n20173) );
  AND U20161 ( .A(n509), .B(n20556), .Z(n20555) );
  XOR U20162 ( .A(n20557), .B(n20554), .Z(n20556) );
  XOR U20163 ( .A(n20558), .B(n20559), .Z(n20546) );
  AND U20164 ( .A(n20560), .B(n20561), .Z(n20559) );
  XOR U20165 ( .A(n20558), .B(n20188), .Z(n20561) );
  XOR U20166 ( .A(n20562), .B(n20563), .Z(n20188) );
  AND U20167 ( .A(n511), .B(n20564), .Z(n20563) );
  XOR U20168 ( .A(n20565), .B(n20562), .Z(n20564) );
  XNOR U20169 ( .A(n20185), .B(n20558), .Z(n20560) );
  XOR U20170 ( .A(n20566), .B(n20567), .Z(n20185) );
  AND U20171 ( .A(n509), .B(n20568), .Z(n20567) );
  XOR U20172 ( .A(n20569), .B(n20566), .Z(n20568) );
  XOR U20173 ( .A(n20570), .B(n20571), .Z(n20558) );
  AND U20174 ( .A(n20572), .B(n20573), .Z(n20571) );
  XOR U20175 ( .A(n20570), .B(n20200), .Z(n20573) );
  XOR U20176 ( .A(n20574), .B(n20575), .Z(n20200) );
  AND U20177 ( .A(n511), .B(n20576), .Z(n20575) );
  XOR U20178 ( .A(n20577), .B(n20574), .Z(n20576) );
  XNOR U20179 ( .A(n20197), .B(n20570), .Z(n20572) );
  XOR U20180 ( .A(n20578), .B(n20579), .Z(n20197) );
  AND U20181 ( .A(n509), .B(n20580), .Z(n20579) );
  XOR U20182 ( .A(n20581), .B(n20578), .Z(n20580) );
  XOR U20183 ( .A(n20582), .B(n20583), .Z(n20570) );
  AND U20184 ( .A(n20584), .B(n20585), .Z(n20583) );
  XOR U20185 ( .A(n20582), .B(n20212), .Z(n20585) );
  XOR U20186 ( .A(n20586), .B(n20587), .Z(n20212) );
  AND U20187 ( .A(n511), .B(n20588), .Z(n20587) );
  XOR U20188 ( .A(n20589), .B(n20586), .Z(n20588) );
  XNOR U20189 ( .A(n20209), .B(n20582), .Z(n20584) );
  XOR U20190 ( .A(n20590), .B(n20591), .Z(n20209) );
  AND U20191 ( .A(n509), .B(n20592), .Z(n20591) );
  XOR U20192 ( .A(n20593), .B(n20590), .Z(n20592) );
  XOR U20193 ( .A(n20594), .B(n20595), .Z(n20582) );
  AND U20194 ( .A(n20596), .B(n20597), .Z(n20595) );
  XOR U20195 ( .A(n20594), .B(n20224), .Z(n20597) );
  XOR U20196 ( .A(n20598), .B(n20599), .Z(n20224) );
  AND U20197 ( .A(n511), .B(n20600), .Z(n20599) );
  XOR U20198 ( .A(n20601), .B(n20598), .Z(n20600) );
  XNOR U20199 ( .A(n20221), .B(n20594), .Z(n20596) );
  XOR U20200 ( .A(n20602), .B(n20603), .Z(n20221) );
  AND U20201 ( .A(n509), .B(n20604), .Z(n20603) );
  XOR U20202 ( .A(n20605), .B(n20602), .Z(n20604) );
  XOR U20203 ( .A(n20606), .B(n20607), .Z(n20594) );
  AND U20204 ( .A(n20608), .B(n20609), .Z(n20607) );
  XOR U20205 ( .A(n20606), .B(n20236), .Z(n20609) );
  XOR U20206 ( .A(n20610), .B(n20611), .Z(n20236) );
  AND U20207 ( .A(n511), .B(n20612), .Z(n20611) );
  XOR U20208 ( .A(n20613), .B(n20610), .Z(n20612) );
  XNOR U20209 ( .A(n20233), .B(n20606), .Z(n20608) );
  XOR U20210 ( .A(n20614), .B(n20615), .Z(n20233) );
  AND U20211 ( .A(n509), .B(n20616), .Z(n20615) );
  XOR U20212 ( .A(n20617), .B(n20614), .Z(n20616) );
  XOR U20213 ( .A(n20618), .B(n20619), .Z(n20606) );
  AND U20214 ( .A(n20620), .B(n20621), .Z(n20619) );
  XOR U20215 ( .A(n20618), .B(n20248), .Z(n20621) );
  XOR U20216 ( .A(n20622), .B(n20623), .Z(n20248) );
  AND U20217 ( .A(n511), .B(n20624), .Z(n20623) );
  XOR U20218 ( .A(n20625), .B(n20622), .Z(n20624) );
  XNOR U20219 ( .A(n20245), .B(n20618), .Z(n20620) );
  XOR U20220 ( .A(n20626), .B(n20627), .Z(n20245) );
  AND U20221 ( .A(n509), .B(n20628), .Z(n20627) );
  XOR U20222 ( .A(n20629), .B(n20626), .Z(n20628) );
  XOR U20223 ( .A(n20630), .B(n20631), .Z(n20618) );
  AND U20224 ( .A(n20632), .B(n20633), .Z(n20631) );
  XOR U20225 ( .A(n20630), .B(n20260), .Z(n20633) );
  XOR U20226 ( .A(n20634), .B(n20635), .Z(n20260) );
  AND U20227 ( .A(n511), .B(n20636), .Z(n20635) );
  XOR U20228 ( .A(n20637), .B(n20634), .Z(n20636) );
  XNOR U20229 ( .A(n20257), .B(n20630), .Z(n20632) );
  XOR U20230 ( .A(n20638), .B(n20639), .Z(n20257) );
  AND U20231 ( .A(n509), .B(n20640), .Z(n20639) );
  XOR U20232 ( .A(n20641), .B(n20638), .Z(n20640) );
  XOR U20233 ( .A(n20642), .B(n20643), .Z(n20630) );
  AND U20234 ( .A(n20644), .B(n20645), .Z(n20643) );
  XOR U20235 ( .A(n20642), .B(n20272), .Z(n20645) );
  XOR U20236 ( .A(n20646), .B(n20647), .Z(n20272) );
  AND U20237 ( .A(n511), .B(n20648), .Z(n20647) );
  XOR U20238 ( .A(n20649), .B(n20646), .Z(n20648) );
  XNOR U20239 ( .A(n20269), .B(n20642), .Z(n20644) );
  XOR U20240 ( .A(n20650), .B(n20651), .Z(n20269) );
  AND U20241 ( .A(n509), .B(n20652), .Z(n20651) );
  XOR U20242 ( .A(n20653), .B(n20650), .Z(n20652) );
  XOR U20243 ( .A(n20654), .B(n20655), .Z(n20642) );
  AND U20244 ( .A(n20656), .B(n20657), .Z(n20655) );
  XOR U20245 ( .A(n20654), .B(n20284), .Z(n20657) );
  XOR U20246 ( .A(n20658), .B(n20659), .Z(n20284) );
  AND U20247 ( .A(n511), .B(n20660), .Z(n20659) );
  XOR U20248 ( .A(n20661), .B(n20658), .Z(n20660) );
  XNOR U20249 ( .A(n20281), .B(n20654), .Z(n20656) );
  XOR U20250 ( .A(n20662), .B(n20663), .Z(n20281) );
  AND U20251 ( .A(n509), .B(n20664), .Z(n20663) );
  XOR U20252 ( .A(n20665), .B(n20662), .Z(n20664) );
  XOR U20253 ( .A(n20666), .B(n20667), .Z(n20654) );
  AND U20254 ( .A(n20668), .B(n20669), .Z(n20667) );
  XOR U20255 ( .A(n20666), .B(n20296), .Z(n20669) );
  XOR U20256 ( .A(n20670), .B(n20671), .Z(n20296) );
  AND U20257 ( .A(n511), .B(n20672), .Z(n20671) );
  XOR U20258 ( .A(n20673), .B(n20670), .Z(n20672) );
  XNOR U20259 ( .A(n20293), .B(n20666), .Z(n20668) );
  XOR U20260 ( .A(n20674), .B(n20675), .Z(n20293) );
  AND U20261 ( .A(n509), .B(n20676), .Z(n20675) );
  XOR U20262 ( .A(n20677), .B(n20674), .Z(n20676) );
  XOR U20263 ( .A(n20678), .B(n20679), .Z(n20666) );
  AND U20264 ( .A(n20680), .B(n20681), .Z(n20679) );
  XOR U20265 ( .A(n20678), .B(n20308), .Z(n20681) );
  XOR U20266 ( .A(n20682), .B(n20683), .Z(n20308) );
  AND U20267 ( .A(n511), .B(n20684), .Z(n20683) );
  XOR U20268 ( .A(n20685), .B(n20682), .Z(n20684) );
  XNOR U20269 ( .A(n20305), .B(n20678), .Z(n20680) );
  XOR U20270 ( .A(n20686), .B(n20687), .Z(n20305) );
  AND U20271 ( .A(n509), .B(n20688), .Z(n20687) );
  XOR U20272 ( .A(n20689), .B(n20686), .Z(n20688) );
  XOR U20273 ( .A(n20690), .B(n20691), .Z(n20678) );
  AND U20274 ( .A(n20692), .B(n20693), .Z(n20691) );
  XOR U20275 ( .A(n20690), .B(n20320), .Z(n20693) );
  XOR U20276 ( .A(n20694), .B(n20695), .Z(n20320) );
  AND U20277 ( .A(n511), .B(n20696), .Z(n20695) );
  XOR U20278 ( .A(n20697), .B(n20694), .Z(n20696) );
  XNOR U20279 ( .A(n20317), .B(n20690), .Z(n20692) );
  XOR U20280 ( .A(n20698), .B(n20699), .Z(n20317) );
  AND U20281 ( .A(n509), .B(n20700), .Z(n20699) );
  XOR U20282 ( .A(n20701), .B(n20698), .Z(n20700) );
  XOR U20283 ( .A(n20702), .B(n20703), .Z(n20690) );
  AND U20284 ( .A(n20704), .B(n20705), .Z(n20703) );
  XOR U20285 ( .A(n20702), .B(n20332), .Z(n20705) );
  XOR U20286 ( .A(n20706), .B(n20707), .Z(n20332) );
  AND U20287 ( .A(n511), .B(n20708), .Z(n20707) );
  XOR U20288 ( .A(n20709), .B(n20706), .Z(n20708) );
  XNOR U20289 ( .A(n20329), .B(n20702), .Z(n20704) );
  XOR U20290 ( .A(n20710), .B(n20711), .Z(n20329) );
  AND U20291 ( .A(n509), .B(n20712), .Z(n20711) );
  XOR U20292 ( .A(n20713), .B(n20710), .Z(n20712) );
  XOR U20293 ( .A(n20714), .B(n20715), .Z(n20702) );
  AND U20294 ( .A(n20716), .B(n20717), .Z(n20715) );
  XOR U20295 ( .A(n20714), .B(n20344), .Z(n20717) );
  XOR U20296 ( .A(n20718), .B(n20719), .Z(n20344) );
  AND U20297 ( .A(n511), .B(n20720), .Z(n20719) );
  XOR U20298 ( .A(n20721), .B(n20718), .Z(n20720) );
  XNOR U20299 ( .A(n20341), .B(n20714), .Z(n20716) );
  XOR U20300 ( .A(n20722), .B(n20723), .Z(n20341) );
  AND U20301 ( .A(n509), .B(n20724), .Z(n20723) );
  XOR U20302 ( .A(n20725), .B(n20722), .Z(n20724) );
  XOR U20303 ( .A(n20726), .B(n20727), .Z(n20714) );
  AND U20304 ( .A(n20728), .B(n20729), .Z(n20727) );
  XOR U20305 ( .A(n20726), .B(n20356), .Z(n20729) );
  XOR U20306 ( .A(n20730), .B(n20731), .Z(n20356) );
  AND U20307 ( .A(n511), .B(n20732), .Z(n20731) );
  XOR U20308 ( .A(n20733), .B(n20730), .Z(n20732) );
  XNOR U20309 ( .A(n20353), .B(n20726), .Z(n20728) );
  XOR U20310 ( .A(n20734), .B(n20735), .Z(n20353) );
  AND U20311 ( .A(n509), .B(n20736), .Z(n20735) );
  XOR U20312 ( .A(n20737), .B(n20734), .Z(n20736) );
  XOR U20313 ( .A(n20738), .B(n20739), .Z(n20726) );
  AND U20314 ( .A(n20740), .B(n20741), .Z(n20739) );
  XOR U20315 ( .A(n20738), .B(n20368), .Z(n20741) );
  XOR U20316 ( .A(n20742), .B(n20743), .Z(n20368) );
  AND U20317 ( .A(n511), .B(n20744), .Z(n20743) );
  XOR U20318 ( .A(n20745), .B(n20742), .Z(n20744) );
  XNOR U20319 ( .A(n20365), .B(n20738), .Z(n20740) );
  XOR U20320 ( .A(n20746), .B(n20747), .Z(n20365) );
  AND U20321 ( .A(n509), .B(n20748), .Z(n20747) );
  XOR U20322 ( .A(n20749), .B(n20746), .Z(n20748) );
  XOR U20323 ( .A(n20750), .B(n20751), .Z(n20738) );
  AND U20324 ( .A(n20752), .B(n20753), .Z(n20751) );
  XOR U20325 ( .A(n20750), .B(n20380), .Z(n20753) );
  XOR U20326 ( .A(n20754), .B(n20755), .Z(n20380) );
  AND U20327 ( .A(n511), .B(n20756), .Z(n20755) );
  XOR U20328 ( .A(n20757), .B(n20754), .Z(n20756) );
  XNOR U20329 ( .A(n20377), .B(n20750), .Z(n20752) );
  XOR U20330 ( .A(n20758), .B(n20759), .Z(n20377) );
  AND U20331 ( .A(n509), .B(n20760), .Z(n20759) );
  XOR U20332 ( .A(n20761), .B(n20758), .Z(n20760) );
  XOR U20333 ( .A(n20762), .B(n20763), .Z(n20750) );
  AND U20334 ( .A(n20764), .B(n20765), .Z(n20763) );
  XOR U20335 ( .A(n20762), .B(n20392), .Z(n20765) );
  XOR U20336 ( .A(n20766), .B(n20767), .Z(n20392) );
  AND U20337 ( .A(n511), .B(n20768), .Z(n20767) );
  XOR U20338 ( .A(n20769), .B(n20766), .Z(n20768) );
  XNOR U20339 ( .A(n20389), .B(n20762), .Z(n20764) );
  XOR U20340 ( .A(n20770), .B(n20771), .Z(n20389) );
  AND U20341 ( .A(n509), .B(n20772), .Z(n20771) );
  XOR U20342 ( .A(n20773), .B(n20770), .Z(n20772) );
  XOR U20343 ( .A(n20774), .B(n20775), .Z(n20762) );
  AND U20344 ( .A(n20776), .B(n20777), .Z(n20775) );
  XOR U20345 ( .A(n20774), .B(n20404), .Z(n20777) );
  XOR U20346 ( .A(n20778), .B(n20779), .Z(n20404) );
  AND U20347 ( .A(n511), .B(n20780), .Z(n20779) );
  XOR U20348 ( .A(n20781), .B(n20778), .Z(n20780) );
  XNOR U20349 ( .A(n20401), .B(n20774), .Z(n20776) );
  XOR U20350 ( .A(n20782), .B(n20783), .Z(n20401) );
  AND U20351 ( .A(n509), .B(n20784), .Z(n20783) );
  XOR U20352 ( .A(n20785), .B(n20782), .Z(n20784) );
  XOR U20353 ( .A(n20786), .B(n20787), .Z(n20774) );
  AND U20354 ( .A(n20788), .B(n20789), .Z(n20787) );
  XOR U20355 ( .A(n20786), .B(n20416), .Z(n20789) );
  XOR U20356 ( .A(n20790), .B(n20791), .Z(n20416) );
  AND U20357 ( .A(n511), .B(n20792), .Z(n20791) );
  XOR U20358 ( .A(n20793), .B(n20790), .Z(n20792) );
  XNOR U20359 ( .A(n20413), .B(n20786), .Z(n20788) );
  XOR U20360 ( .A(n20794), .B(n20795), .Z(n20413) );
  AND U20361 ( .A(n509), .B(n20796), .Z(n20795) );
  XOR U20362 ( .A(n20797), .B(n20794), .Z(n20796) );
  XOR U20363 ( .A(n20798), .B(n20799), .Z(n20786) );
  AND U20364 ( .A(n20800), .B(n20801), .Z(n20799) );
  XOR U20365 ( .A(n20798), .B(n20428), .Z(n20801) );
  XOR U20366 ( .A(n20802), .B(n20803), .Z(n20428) );
  AND U20367 ( .A(n511), .B(n20804), .Z(n20803) );
  XOR U20368 ( .A(n20805), .B(n20802), .Z(n20804) );
  XNOR U20369 ( .A(n20425), .B(n20798), .Z(n20800) );
  XOR U20370 ( .A(n20806), .B(n20807), .Z(n20425) );
  AND U20371 ( .A(n509), .B(n20808), .Z(n20807) );
  XOR U20372 ( .A(n20809), .B(n20806), .Z(n20808) );
  XOR U20373 ( .A(n20810), .B(n20811), .Z(n20798) );
  AND U20374 ( .A(n20812), .B(n20813), .Z(n20811) );
  XOR U20375 ( .A(n20810), .B(n20440), .Z(n20813) );
  XOR U20376 ( .A(n20814), .B(n20815), .Z(n20440) );
  AND U20377 ( .A(n511), .B(n20816), .Z(n20815) );
  XOR U20378 ( .A(n20817), .B(n20814), .Z(n20816) );
  XNOR U20379 ( .A(n20437), .B(n20810), .Z(n20812) );
  XOR U20380 ( .A(n20818), .B(n20819), .Z(n20437) );
  AND U20381 ( .A(n509), .B(n20820), .Z(n20819) );
  XOR U20382 ( .A(n20821), .B(n20818), .Z(n20820) );
  XOR U20383 ( .A(n20822), .B(n20823), .Z(n20810) );
  AND U20384 ( .A(n20824), .B(n20825), .Z(n20823) );
  XOR U20385 ( .A(n20822), .B(n20452), .Z(n20825) );
  XOR U20386 ( .A(n20826), .B(n20827), .Z(n20452) );
  AND U20387 ( .A(n511), .B(n20828), .Z(n20827) );
  XOR U20388 ( .A(n20829), .B(n20826), .Z(n20828) );
  XNOR U20389 ( .A(n20449), .B(n20822), .Z(n20824) );
  XOR U20390 ( .A(n20830), .B(n20831), .Z(n20449) );
  AND U20391 ( .A(n509), .B(n20832), .Z(n20831) );
  XOR U20392 ( .A(n20833), .B(n20830), .Z(n20832) );
  XOR U20393 ( .A(n20834), .B(n20835), .Z(n20822) );
  AND U20394 ( .A(n20836), .B(n20837), .Z(n20835) );
  XOR U20395 ( .A(n20834), .B(n20464), .Z(n20837) );
  XOR U20396 ( .A(n20838), .B(n20839), .Z(n20464) );
  AND U20397 ( .A(n511), .B(n20840), .Z(n20839) );
  XOR U20398 ( .A(n20841), .B(n20838), .Z(n20840) );
  XNOR U20399 ( .A(n20461), .B(n20834), .Z(n20836) );
  XOR U20400 ( .A(n20842), .B(n20843), .Z(n20461) );
  AND U20401 ( .A(n509), .B(n20844), .Z(n20843) );
  XOR U20402 ( .A(n20845), .B(n20842), .Z(n20844) );
  XOR U20403 ( .A(n20846), .B(n20847), .Z(n20834) );
  AND U20404 ( .A(n20848), .B(n20849), .Z(n20847) );
  XOR U20405 ( .A(n20846), .B(n20476), .Z(n20849) );
  XOR U20406 ( .A(n20850), .B(n20851), .Z(n20476) );
  AND U20407 ( .A(n511), .B(n20852), .Z(n20851) );
  XOR U20408 ( .A(n20853), .B(n20850), .Z(n20852) );
  XNOR U20409 ( .A(n20473), .B(n20846), .Z(n20848) );
  XOR U20410 ( .A(n20854), .B(n20855), .Z(n20473) );
  AND U20411 ( .A(n509), .B(n20856), .Z(n20855) );
  XOR U20412 ( .A(n20857), .B(n20854), .Z(n20856) );
  XOR U20413 ( .A(n20858), .B(n20859), .Z(n20846) );
  AND U20414 ( .A(n20860), .B(n20861), .Z(n20859) );
  XNOR U20415 ( .A(n20862), .B(n20489), .Z(n20861) );
  XOR U20416 ( .A(n20863), .B(n20864), .Z(n20489) );
  AND U20417 ( .A(n511), .B(n20865), .Z(n20864) );
  XOR U20418 ( .A(n20863), .B(n20866), .Z(n20865) );
  XNOR U20419 ( .A(n20486), .B(n20858), .Z(n20860) );
  XOR U20420 ( .A(n20867), .B(n20868), .Z(n20486) );
  AND U20421 ( .A(n509), .B(n20869), .Z(n20868) );
  XOR U20422 ( .A(n20867), .B(n20870), .Z(n20869) );
  IV U20423 ( .A(n20862), .Z(n20858) );
  AND U20424 ( .A(n20494), .B(n20497), .Z(n20862) );
  XNOR U20425 ( .A(n20871), .B(n20872), .Z(n20497) );
  AND U20426 ( .A(n511), .B(n20873), .Z(n20872) );
  XNOR U20427 ( .A(n20874), .B(n20871), .Z(n20873) );
  XOR U20428 ( .A(n20875), .B(n20876), .Z(n511) );
  AND U20429 ( .A(n20877), .B(n20878), .Z(n20876) );
  XOR U20430 ( .A(n20505), .B(n20875), .Z(n20878) );
  IV U20431 ( .A(n20879), .Z(n20505) );
  AND U20432 ( .A(p_input[5631]), .B(p_input[5599]), .Z(n20879) );
  XOR U20433 ( .A(n20875), .B(n20502), .Z(n20877) );
  AND U20434 ( .A(p_input[5535]), .B(p_input[5567]), .Z(n20502) );
  XOR U20435 ( .A(n20880), .B(n20881), .Z(n20875) );
  AND U20436 ( .A(n20882), .B(n20883), .Z(n20881) );
  XOR U20437 ( .A(n20880), .B(n20517), .Z(n20883) );
  XNOR U20438 ( .A(p_input[5598]), .B(n20884), .Z(n20517) );
  AND U20439 ( .A(n339), .B(n20885), .Z(n20884) );
  XOR U20440 ( .A(p_input[5630]), .B(p_input[5598]), .Z(n20885) );
  XNOR U20441 ( .A(n20514), .B(n20880), .Z(n20882) );
  XOR U20442 ( .A(n20886), .B(n20887), .Z(n20514) );
  AND U20443 ( .A(n337), .B(n20888), .Z(n20887) );
  XOR U20444 ( .A(p_input[5566]), .B(p_input[5534]), .Z(n20888) );
  XOR U20445 ( .A(n20889), .B(n20890), .Z(n20880) );
  AND U20446 ( .A(n20891), .B(n20892), .Z(n20890) );
  XOR U20447 ( .A(n20889), .B(n20529), .Z(n20892) );
  XNOR U20448 ( .A(p_input[5597]), .B(n20893), .Z(n20529) );
  AND U20449 ( .A(n339), .B(n20894), .Z(n20893) );
  XOR U20450 ( .A(p_input[5629]), .B(p_input[5597]), .Z(n20894) );
  XNOR U20451 ( .A(n20526), .B(n20889), .Z(n20891) );
  XOR U20452 ( .A(n20895), .B(n20896), .Z(n20526) );
  AND U20453 ( .A(n337), .B(n20897), .Z(n20896) );
  XOR U20454 ( .A(p_input[5565]), .B(p_input[5533]), .Z(n20897) );
  XOR U20455 ( .A(n20898), .B(n20899), .Z(n20889) );
  AND U20456 ( .A(n20900), .B(n20901), .Z(n20899) );
  XOR U20457 ( .A(n20898), .B(n20541), .Z(n20901) );
  XNOR U20458 ( .A(p_input[5596]), .B(n20902), .Z(n20541) );
  AND U20459 ( .A(n339), .B(n20903), .Z(n20902) );
  XOR U20460 ( .A(p_input[5628]), .B(p_input[5596]), .Z(n20903) );
  XNOR U20461 ( .A(n20538), .B(n20898), .Z(n20900) );
  XOR U20462 ( .A(n20904), .B(n20905), .Z(n20538) );
  AND U20463 ( .A(n337), .B(n20906), .Z(n20905) );
  XOR U20464 ( .A(p_input[5564]), .B(p_input[5532]), .Z(n20906) );
  XOR U20465 ( .A(n20907), .B(n20908), .Z(n20898) );
  AND U20466 ( .A(n20909), .B(n20910), .Z(n20908) );
  XOR U20467 ( .A(n20907), .B(n20553), .Z(n20910) );
  XNOR U20468 ( .A(p_input[5595]), .B(n20911), .Z(n20553) );
  AND U20469 ( .A(n339), .B(n20912), .Z(n20911) );
  XOR U20470 ( .A(p_input[5627]), .B(p_input[5595]), .Z(n20912) );
  XNOR U20471 ( .A(n20550), .B(n20907), .Z(n20909) );
  XOR U20472 ( .A(n20913), .B(n20914), .Z(n20550) );
  AND U20473 ( .A(n337), .B(n20915), .Z(n20914) );
  XOR U20474 ( .A(p_input[5563]), .B(p_input[5531]), .Z(n20915) );
  XOR U20475 ( .A(n20916), .B(n20917), .Z(n20907) );
  AND U20476 ( .A(n20918), .B(n20919), .Z(n20917) );
  XOR U20477 ( .A(n20916), .B(n20565), .Z(n20919) );
  XNOR U20478 ( .A(p_input[5594]), .B(n20920), .Z(n20565) );
  AND U20479 ( .A(n339), .B(n20921), .Z(n20920) );
  XOR U20480 ( .A(p_input[5626]), .B(p_input[5594]), .Z(n20921) );
  XNOR U20481 ( .A(n20562), .B(n20916), .Z(n20918) );
  XOR U20482 ( .A(n20922), .B(n20923), .Z(n20562) );
  AND U20483 ( .A(n337), .B(n20924), .Z(n20923) );
  XOR U20484 ( .A(p_input[5562]), .B(p_input[5530]), .Z(n20924) );
  XOR U20485 ( .A(n20925), .B(n20926), .Z(n20916) );
  AND U20486 ( .A(n20927), .B(n20928), .Z(n20926) );
  XOR U20487 ( .A(n20925), .B(n20577), .Z(n20928) );
  XNOR U20488 ( .A(p_input[5593]), .B(n20929), .Z(n20577) );
  AND U20489 ( .A(n339), .B(n20930), .Z(n20929) );
  XOR U20490 ( .A(p_input[5625]), .B(p_input[5593]), .Z(n20930) );
  XNOR U20491 ( .A(n20574), .B(n20925), .Z(n20927) );
  XOR U20492 ( .A(n20931), .B(n20932), .Z(n20574) );
  AND U20493 ( .A(n337), .B(n20933), .Z(n20932) );
  XOR U20494 ( .A(p_input[5561]), .B(p_input[5529]), .Z(n20933) );
  XOR U20495 ( .A(n20934), .B(n20935), .Z(n20925) );
  AND U20496 ( .A(n20936), .B(n20937), .Z(n20935) );
  XOR U20497 ( .A(n20934), .B(n20589), .Z(n20937) );
  XNOR U20498 ( .A(p_input[5592]), .B(n20938), .Z(n20589) );
  AND U20499 ( .A(n339), .B(n20939), .Z(n20938) );
  XOR U20500 ( .A(p_input[5624]), .B(p_input[5592]), .Z(n20939) );
  XNOR U20501 ( .A(n20586), .B(n20934), .Z(n20936) );
  XOR U20502 ( .A(n20940), .B(n20941), .Z(n20586) );
  AND U20503 ( .A(n337), .B(n20942), .Z(n20941) );
  XOR U20504 ( .A(p_input[5560]), .B(p_input[5528]), .Z(n20942) );
  XOR U20505 ( .A(n20943), .B(n20944), .Z(n20934) );
  AND U20506 ( .A(n20945), .B(n20946), .Z(n20944) );
  XOR U20507 ( .A(n20943), .B(n20601), .Z(n20946) );
  XNOR U20508 ( .A(p_input[5591]), .B(n20947), .Z(n20601) );
  AND U20509 ( .A(n339), .B(n20948), .Z(n20947) );
  XOR U20510 ( .A(p_input[5623]), .B(p_input[5591]), .Z(n20948) );
  XNOR U20511 ( .A(n20598), .B(n20943), .Z(n20945) );
  XOR U20512 ( .A(n20949), .B(n20950), .Z(n20598) );
  AND U20513 ( .A(n337), .B(n20951), .Z(n20950) );
  XOR U20514 ( .A(p_input[5559]), .B(p_input[5527]), .Z(n20951) );
  XOR U20515 ( .A(n20952), .B(n20953), .Z(n20943) );
  AND U20516 ( .A(n20954), .B(n20955), .Z(n20953) );
  XOR U20517 ( .A(n20952), .B(n20613), .Z(n20955) );
  XNOR U20518 ( .A(p_input[5590]), .B(n20956), .Z(n20613) );
  AND U20519 ( .A(n339), .B(n20957), .Z(n20956) );
  XOR U20520 ( .A(p_input[5622]), .B(p_input[5590]), .Z(n20957) );
  XNOR U20521 ( .A(n20610), .B(n20952), .Z(n20954) );
  XOR U20522 ( .A(n20958), .B(n20959), .Z(n20610) );
  AND U20523 ( .A(n337), .B(n20960), .Z(n20959) );
  XOR U20524 ( .A(p_input[5558]), .B(p_input[5526]), .Z(n20960) );
  XOR U20525 ( .A(n20961), .B(n20962), .Z(n20952) );
  AND U20526 ( .A(n20963), .B(n20964), .Z(n20962) );
  XOR U20527 ( .A(n20961), .B(n20625), .Z(n20964) );
  XNOR U20528 ( .A(p_input[5589]), .B(n20965), .Z(n20625) );
  AND U20529 ( .A(n339), .B(n20966), .Z(n20965) );
  XOR U20530 ( .A(p_input[5621]), .B(p_input[5589]), .Z(n20966) );
  XNOR U20531 ( .A(n20622), .B(n20961), .Z(n20963) );
  XOR U20532 ( .A(n20967), .B(n20968), .Z(n20622) );
  AND U20533 ( .A(n337), .B(n20969), .Z(n20968) );
  XOR U20534 ( .A(p_input[5557]), .B(p_input[5525]), .Z(n20969) );
  XOR U20535 ( .A(n20970), .B(n20971), .Z(n20961) );
  AND U20536 ( .A(n20972), .B(n20973), .Z(n20971) );
  XOR U20537 ( .A(n20970), .B(n20637), .Z(n20973) );
  XNOR U20538 ( .A(p_input[5588]), .B(n20974), .Z(n20637) );
  AND U20539 ( .A(n339), .B(n20975), .Z(n20974) );
  XOR U20540 ( .A(p_input[5620]), .B(p_input[5588]), .Z(n20975) );
  XNOR U20541 ( .A(n20634), .B(n20970), .Z(n20972) );
  XOR U20542 ( .A(n20976), .B(n20977), .Z(n20634) );
  AND U20543 ( .A(n337), .B(n20978), .Z(n20977) );
  XOR U20544 ( .A(p_input[5556]), .B(p_input[5524]), .Z(n20978) );
  XOR U20545 ( .A(n20979), .B(n20980), .Z(n20970) );
  AND U20546 ( .A(n20981), .B(n20982), .Z(n20980) );
  XOR U20547 ( .A(n20979), .B(n20649), .Z(n20982) );
  XNOR U20548 ( .A(p_input[5587]), .B(n20983), .Z(n20649) );
  AND U20549 ( .A(n339), .B(n20984), .Z(n20983) );
  XOR U20550 ( .A(p_input[5619]), .B(p_input[5587]), .Z(n20984) );
  XNOR U20551 ( .A(n20646), .B(n20979), .Z(n20981) );
  XOR U20552 ( .A(n20985), .B(n20986), .Z(n20646) );
  AND U20553 ( .A(n337), .B(n20987), .Z(n20986) );
  XOR U20554 ( .A(p_input[5555]), .B(p_input[5523]), .Z(n20987) );
  XOR U20555 ( .A(n20988), .B(n20989), .Z(n20979) );
  AND U20556 ( .A(n20990), .B(n20991), .Z(n20989) );
  XOR U20557 ( .A(n20988), .B(n20661), .Z(n20991) );
  XNOR U20558 ( .A(p_input[5586]), .B(n20992), .Z(n20661) );
  AND U20559 ( .A(n339), .B(n20993), .Z(n20992) );
  XOR U20560 ( .A(p_input[5618]), .B(p_input[5586]), .Z(n20993) );
  XNOR U20561 ( .A(n20658), .B(n20988), .Z(n20990) );
  XOR U20562 ( .A(n20994), .B(n20995), .Z(n20658) );
  AND U20563 ( .A(n337), .B(n20996), .Z(n20995) );
  XOR U20564 ( .A(p_input[5554]), .B(p_input[5522]), .Z(n20996) );
  XOR U20565 ( .A(n20997), .B(n20998), .Z(n20988) );
  AND U20566 ( .A(n20999), .B(n21000), .Z(n20998) );
  XOR U20567 ( .A(n20997), .B(n20673), .Z(n21000) );
  XNOR U20568 ( .A(p_input[5585]), .B(n21001), .Z(n20673) );
  AND U20569 ( .A(n339), .B(n21002), .Z(n21001) );
  XOR U20570 ( .A(p_input[5617]), .B(p_input[5585]), .Z(n21002) );
  XNOR U20571 ( .A(n20670), .B(n20997), .Z(n20999) );
  XOR U20572 ( .A(n21003), .B(n21004), .Z(n20670) );
  AND U20573 ( .A(n337), .B(n21005), .Z(n21004) );
  XOR U20574 ( .A(p_input[5553]), .B(p_input[5521]), .Z(n21005) );
  XOR U20575 ( .A(n21006), .B(n21007), .Z(n20997) );
  AND U20576 ( .A(n21008), .B(n21009), .Z(n21007) );
  XOR U20577 ( .A(n21006), .B(n20685), .Z(n21009) );
  XNOR U20578 ( .A(p_input[5584]), .B(n21010), .Z(n20685) );
  AND U20579 ( .A(n339), .B(n21011), .Z(n21010) );
  XOR U20580 ( .A(p_input[5616]), .B(p_input[5584]), .Z(n21011) );
  XNOR U20581 ( .A(n20682), .B(n21006), .Z(n21008) );
  XOR U20582 ( .A(n21012), .B(n21013), .Z(n20682) );
  AND U20583 ( .A(n337), .B(n21014), .Z(n21013) );
  XOR U20584 ( .A(p_input[5552]), .B(p_input[5520]), .Z(n21014) );
  XOR U20585 ( .A(n21015), .B(n21016), .Z(n21006) );
  AND U20586 ( .A(n21017), .B(n21018), .Z(n21016) );
  XOR U20587 ( .A(n21015), .B(n20697), .Z(n21018) );
  XNOR U20588 ( .A(p_input[5583]), .B(n21019), .Z(n20697) );
  AND U20589 ( .A(n339), .B(n21020), .Z(n21019) );
  XOR U20590 ( .A(p_input[5615]), .B(p_input[5583]), .Z(n21020) );
  XNOR U20591 ( .A(n20694), .B(n21015), .Z(n21017) );
  XOR U20592 ( .A(n21021), .B(n21022), .Z(n20694) );
  AND U20593 ( .A(n337), .B(n21023), .Z(n21022) );
  XOR U20594 ( .A(p_input[5551]), .B(p_input[5519]), .Z(n21023) );
  XOR U20595 ( .A(n21024), .B(n21025), .Z(n21015) );
  AND U20596 ( .A(n21026), .B(n21027), .Z(n21025) );
  XOR U20597 ( .A(n21024), .B(n20709), .Z(n21027) );
  XNOR U20598 ( .A(p_input[5582]), .B(n21028), .Z(n20709) );
  AND U20599 ( .A(n339), .B(n21029), .Z(n21028) );
  XOR U20600 ( .A(p_input[5614]), .B(p_input[5582]), .Z(n21029) );
  XNOR U20601 ( .A(n20706), .B(n21024), .Z(n21026) );
  XOR U20602 ( .A(n21030), .B(n21031), .Z(n20706) );
  AND U20603 ( .A(n337), .B(n21032), .Z(n21031) );
  XOR U20604 ( .A(p_input[5550]), .B(p_input[5518]), .Z(n21032) );
  XOR U20605 ( .A(n21033), .B(n21034), .Z(n21024) );
  AND U20606 ( .A(n21035), .B(n21036), .Z(n21034) );
  XOR U20607 ( .A(n21033), .B(n20721), .Z(n21036) );
  XNOR U20608 ( .A(p_input[5581]), .B(n21037), .Z(n20721) );
  AND U20609 ( .A(n339), .B(n21038), .Z(n21037) );
  XOR U20610 ( .A(p_input[5613]), .B(p_input[5581]), .Z(n21038) );
  XNOR U20611 ( .A(n20718), .B(n21033), .Z(n21035) );
  XOR U20612 ( .A(n21039), .B(n21040), .Z(n20718) );
  AND U20613 ( .A(n337), .B(n21041), .Z(n21040) );
  XOR U20614 ( .A(p_input[5549]), .B(p_input[5517]), .Z(n21041) );
  XOR U20615 ( .A(n21042), .B(n21043), .Z(n21033) );
  AND U20616 ( .A(n21044), .B(n21045), .Z(n21043) );
  XOR U20617 ( .A(n21042), .B(n20733), .Z(n21045) );
  XNOR U20618 ( .A(p_input[5580]), .B(n21046), .Z(n20733) );
  AND U20619 ( .A(n339), .B(n21047), .Z(n21046) );
  XOR U20620 ( .A(p_input[5612]), .B(p_input[5580]), .Z(n21047) );
  XNOR U20621 ( .A(n20730), .B(n21042), .Z(n21044) );
  XOR U20622 ( .A(n21048), .B(n21049), .Z(n20730) );
  AND U20623 ( .A(n337), .B(n21050), .Z(n21049) );
  XOR U20624 ( .A(p_input[5548]), .B(p_input[5516]), .Z(n21050) );
  XOR U20625 ( .A(n21051), .B(n21052), .Z(n21042) );
  AND U20626 ( .A(n21053), .B(n21054), .Z(n21052) );
  XOR U20627 ( .A(n21051), .B(n20745), .Z(n21054) );
  XNOR U20628 ( .A(p_input[5579]), .B(n21055), .Z(n20745) );
  AND U20629 ( .A(n339), .B(n21056), .Z(n21055) );
  XOR U20630 ( .A(p_input[5611]), .B(p_input[5579]), .Z(n21056) );
  XNOR U20631 ( .A(n20742), .B(n21051), .Z(n21053) );
  XOR U20632 ( .A(n21057), .B(n21058), .Z(n20742) );
  AND U20633 ( .A(n337), .B(n21059), .Z(n21058) );
  XOR U20634 ( .A(p_input[5547]), .B(p_input[5515]), .Z(n21059) );
  XOR U20635 ( .A(n21060), .B(n21061), .Z(n21051) );
  AND U20636 ( .A(n21062), .B(n21063), .Z(n21061) );
  XOR U20637 ( .A(n21060), .B(n20757), .Z(n21063) );
  XNOR U20638 ( .A(p_input[5578]), .B(n21064), .Z(n20757) );
  AND U20639 ( .A(n339), .B(n21065), .Z(n21064) );
  XOR U20640 ( .A(p_input[5610]), .B(p_input[5578]), .Z(n21065) );
  XNOR U20641 ( .A(n20754), .B(n21060), .Z(n21062) );
  XOR U20642 ( .A(n21066), .B(n21067), .Z(n20754) );
  AND U20643 ( .A(n337), .B(n21068), .Z(n21067) );
  XOR U20644 ( .A(p_input[5546]), .B(p_input[5514]), .Z(n21068) );
  XOR U20645 ( .A(n21069), .B(n21070), .Z(n21060) );
  AND U20646 ( .A(n21071), .B(n21072), .Z(n21070) );
  XOR U20647 ( .A(n21069), .B(n20769), .Z(n21072) );
  XNOR U20648 ( .A(p_input[5577]), .B(n21073), .Z(n20769) );
  AND U20649 ( .A(n339), .B(n21074), .Z(n21073) );
  XOR U20650 ( .A(p_input[5609]), .B(p_input[5577]), .Z(n21074) );
  XNOR U20651 ( .A(n20766), .B(n21069), .Z(n21071) );
  XOR U20652 ( .A(n21075), .B(n21076), .Z(n20766) );
  AND U20653 ( .A(n337), .B(n21077), .Z(n21076) );
  XOR U20654 ( .A(p_input[5545]), .B(p_input[5513]), .Z(n21077) );
  XOR U20655 ( .A(n21078), .B(n21079), .Z(n21069) );
  AND U20656 ( .A(n21080), .B(n21081), .Z(n21079) );
  XOR U20657 ( .A(n21078), .B(n20781), .Z(n21081) );
  XNOR U20658 ( .A(p_input[5576]), .B(n21082), .Z(n20781) );
  AND U20659 ( .A(n339), .B(n21083), .Z(n21082) );
  XOR U20660 ( .A(p_input[5608]), .B(p_input[5576]), .Z(n21083) );
  XNOR U20661 ( .A(n20778), .B(n21078), .Z(n21080) );
  XOR U20662 ( .A(n21084), .B(n21085), .Z(n20778) );
  AND U20663 ( .A(n337), .B(n21086), .Z(n21085) );
  XOR U20664 ( .A(p_input[5544]), .B(p_input[5512]), .Z(n21086) );
  XOR U20665 ( .A(n21087), .B(n21088), .Z(n21078) );
  AND U20666 ( .A(n21089), .B(n21090), .Z(n21088) );
  XOR U20667 ( .A(n21087), .B(n20793), .Z(n21090) );
  XNOR U20668 ( .A(p_input[5575]), .B(n21091), .Z(n20793) );
  AND U20669 ( .A(n339), .B(n21092), .Z(n21091) );
  XOR U20670 ( .A(p_input[5607]), .B(p_input[5575]), .Z(n21092) );
  XNOR U20671 ( .A(n20790), .B(n21087), .Z(n21089) );
  XOR U20672 ( .A(n21093), .B(n21094), .Z(n20790) );
  AND U20673 ( .A(n337), .B(n21095), .Z(n21094) );
  XOR U20674 ( .A(p_input[5543]), .B(p_input[5511]), .Z(n21095) );
  XOR U20675 ( .A(n21096), .B(n21097), .Z(n21087) );
  AND U20676 ( .A(n21098), .B(n21099), .Z(n21097) );
  XOR U20677 ( .A(n21096), .B(n20805), .Z(n21099) );
  XNOR U20678 ( .A(p_input[5574]), .B(n21100), .Z(n20805) );
  AND U20679 ( .A(n339), .B(n21101), .Z(n21100) );
  XOR U20680 ( .A(p_input[5606]), .B(p_input[5574]), .Z(n21101) );
  XNOR U20681 ( .A(n20802), .B(n21096), .Z(n21098) );
  XOR U20682 ( .A(n21102), .B(n21103), .Z(n20802) );
  AND U20683 ( .A(n337), .B(n21104), .Z(n21103) );
  XOR U20684 ( .A(p_input[5542]), .B(p_input[5510]), .Z(n21104) );
  XOR U20685 ( .A(n21105), .B(n21106), .Z(n21096) );
  AND U20686 ( .A(n21107), .B(n21108), .Z(n21106) );
  XOR U20687 ( .A(n21105), .B(n20817), .Z(n21108) );
  XNOR U20688 ( .A(p_input[5573]), .B(n21109), .Z(n20817) );
  AND U20689 ( .A(n339), .B(n21110), .Z(n21109) );
  XOR U20690 ( .A(p_input[5605]), .B(p_input[5573]), .Z(n21110) );
  XNOR U20691 ( .A(n20814), .B(n21105), .Z(n21107) );
  XOR U20692 ( .A(n21111), .B(n21112), .Z(n20814) );
  AND U20693 ( .A(n337), .B(n21113), .Z(n21112) );
  XOR U20694 ( .A(p_input[5541]), .B(p_input[5509]), .Z(n21113) );
  XOR U20695 ( .A(n21114), .B(n21115), .Z(n21105) );
  AND U20696 ( .A(n21116), .B(n21117), .Z(n21115) );
  XOR U20697 ( .A(n21114), .B(n20829), .Z(n21117) );
  XNOR U20698 ( .A(p_input[5572]), .B(n21118), .Z(n20829) );
  AND U20699 ( .A(n339), .B(n21119), .Z(n21118) );
  XOR U20700 ( .A(p_input[5604]), .B(p_input[5572]), .Z(n21119) );
  XNOR U20701 ( .A(n20826), .B(n21114), .Z(n21116) );
  XOR U20702 ( .A(n21120), .B(n21121), .Z(n20826) );
  AND U20703 ( .A(n337), .B(n21122), .Z(n21121) );
  XOR U20704 ( .A(p_input[5540]), .B(p_input[5508]), .Z(n21122) );
  XOR U20705 ( .A(n21123), .B(n21124), .Z(n21114) );
  AND U20706 ( .A(n21125), .B(n21126), .Z(n21124) );
  XOR U20707 ( .A(n21123), .B(n20841), .Z(n21126) );
  XNOR U20708 ( .A(p_input[5571]), .B(n21127), .Z(n20841) );
  AND U20709 ( .A(n339), .B(n21128), .Z(n21127) );
  XOR U20710 ( .A(p_input[5603]), .B(p_input[5571]), .Z(n21128) );
  XNOR U20711 ( .A(n20838), .B(n21123), .Z(n21125) );
  XOR U20712 ( .A(n21129), .B(n21130), .Z(n20838) );
  AND U20713 ( .A(n337), .B(n21131), .Z(n21130) );
  XOR U20714 ( .A(p_input[5539]), .B(p_input[5507]), .Z(n21131) );
  XOR U20715 ( .A(n21132), .B(n21133), .Z(n21123) );
  AND U20716 ( .A(n21134), .B(n21135), .Z(n21133) );
  XOR U20717 ( .A(n21132), .B(n20853), .Z(n21135) );
  XNOR U20718 ( .A(p_input[5570]), .B(n21136), .Z(n20853) );
  AND U20719 ( .A(n339), .B(n21137), .Z(n21136) );
  XOR U20720 ( .A(p_input[5602]), .B(p_input[5570]), .Z(n21137) );
  XNOR U20721 ( .A(n20850), .B(n21132), .Z(n21134) );
  XOR U20722 ( .A(n21138), .B(n21139), .Z(n20850) );
  AND U20723 ( .A(n337), .B(n21140), .Z(n21139) );
  XOR U20724 ( .A(p_input[5538]), .B(p_input[5506]), .Z(n21140) );
  XOR U20725 ( .A(n21141), .B(n21142), .Z(n21132) );
  AND U20726 ( .A(n21143), .B(n21144), .Z(n21142) );
  XNOR U20727 ( .A(n21145), .B(n20866), .Z(n21144) );
  XNOR U20728 ( .A(p_input[5569]), .B(n21146), .Z(n20866) );
  AND U20729 ( .A(n339), .B(n21147), .Z(n21146) );
  XNOR U20730 ( .A(p_input[5601]), .B(n21148), .Z(n21147) );
  IV U20731 ( .A(p_input[5569]), .Z(n21148) );
  XNOR U20732 ( .A(n20863), .B(n21141), .Z(n21143) );
  XNOR U20733 ( .A(p_input[5505]), .B(n21149), .Z(n20863) );
  AND U20734 ( .A(n337), .B(n21150), .Z(n21149) );
  XOR U20735 ( .A(p_input[5537]), .B(p_input[5505]), .Z(n21150) );
  IV U20736 ( .A(n21145), .Z(n21141) );
  AND U20737 ( .A(n20871), .B(n20874), .Z(n21145) );
  XOR U20738 ( .A(p_input[5568]), .B(n21151), .Z(n20874) );
  AND U20739 ( .A(n339), .B(n21152), .Z(n21151) );
  XOR U20740 ( .A(p_input[5600]), .B(p_input[5568]), .Z(n21152) );
  XOR U20741 ( .A(n21153), .B(n21154), .Z(n339) );
  AND U20742 ( .A(n21155), .B(n21156), .Z(n21154) );
  XNOR U20743 ( .A(p_input[5631]), .B(n21153), .Z(n21156) );
  XOR U20744 ( .A(n21153), .B(p_input[5599]), .Z(n21155) );
  XOR U20745 ( .A(n21157), .B(n21158), .Z(n21153) );
  AND U20746 ( .A(n21159), .B(n21160), .Z(n21158) );
  XNOR U20747 ( .A(p_input[5630]), .B(n21157), .Z(n21160) );
  XOR U20748 ( .A(n21157), .B(p_input[5598]), .Z(n21159) );
  XOR U20749 ( .A(n21161), .B(n21162), .Z(n21157) );
  AND U20750 ( .A(n21163), .B(n21164), .Z(n21162) );
  XNOR U20751 ( .A(p_input[5629]), .B(n21161), .Z(n21164) );
  XOR U20752 ( .A(n21161), .B(p_input[5597]), .Z(n21163) );
  XOR U20753 ( .A(n21165), .B(n21166), .Z(n21161) );
  AND U20754 ( .A(n21167), .B(n21168), .Z(n21166) );
  XNOR U20755 ( .A(p_input[5628]), .B(n21165), .Z(n21168) );
  XOR U20756 ( .A(n21165), .B(p_input[5596]), .Z(n21167) );
  XOR U20757 ( .A(n21169), .B(n21170), .Z(n21165) );
  AND U20758 ( .A(n21171), .B(n21172), .Z(n21170) );
  XNOR U20759 ( .A(p_input[5627]), .B(n21169), .Z(n21172) );
  XOR U20760 ( .A(n21169), .B(p_input[5595]), .Z(n21171) );
  XOR U20761 ( .A(n21173), .B(n21174), .Z(n21169) );
  AND U20762 ( .A(n21175), .B(n21176), .Z(n21174) );
  XNOR U20763 ( .A(p_input[5626]), .B(n21173), .Z(n21176) );
  XOR U20764 ( .A(n21173), .B(p_input[5594]), .Z(n21175) );
  XOR U20765 ( .A(n21177), .B(n21178), .Z(n21173) );
  AND U20766 ( .A(n21179), .B(n21180), .Z(n21178) );
  XNOR U20767 ( .A(p_input[5625]), .B(n21177), .Z(n21180) );
  XOR U20768 ( .A(n21177), .B(p_input[5593]), .Z(n21179) );
  XOR U20769 ( .A(n21181), .B(n21182), .Z(n21177) );
  AND U20770 ( .A(n21183), .B(n21184), .Z(n21182) );
  XNOR U20771 ( .A(p_input[5624]), .B(n21181), .Z(n21184) );
  XOR U20772 ( .A(n21181), .B(p_input[5592]), .Z(n21183) );
  XOR U20773 ( .A(n21185), .B(n21186), .Z(n21181) );
  AND U20774 ( .A(n21187), .B(n21188), .Z(n21186) );
  XNOR U20775 ( .A(p_input[5623]), .B(n21185), .Z(n21188) );
  XOR U20776 ( .A(n21185), .B(p_input[5591]), .Z(n21187) );
  XOR U20777 ( .A(n21189), .B(n21190), .Z(n21185) );
  AND U20778 ( .A(n21191), .B(n21192), .Z(n21190) );
  XNOR U20779 ( .A(p_input[5622]), .B(n21189), .Z(n21192) );
  XOR U20780 ( .A(n21189), .B(p_input[5590]), .Z(n21191) );
  XOR U20781 ( .A(n21193), .B(n21194), .Z(n21189) );
  AND U20782 ( .A(n21195), .B(n21196), .Z(n21194) );
  XNOR U20783 ( .A(p_input[5621]), .B(n21193), .Z(n21196) );
  XOR U20784 ( .A(n21193), .B(p_input[5589]), .Z(n21195) );
  XOR U20785 ( .A(n21197), .B(n21198), .Z(n21193) );
  AND U20786 ( .A(n21199), .B(n21200), .Z(n21198) );
  XNOR U20787 ( .A(p_input[5620]), .B(n21197), .Z(n21200) );
  XOR U20788 ( .A(n21197), .B(p_input[5588]), .Z(n21199) );
  XOR U20789 ( .A(n21201), .B(n21202), .Z(n21197) );
  AND U20790 ( .A(n21203), .B(n21204), .Z(n21202) );
  XNOR U20791 ( .A(p_input[5619]), .B(n21201), .Z(n21204) );
  XOR U20792 ( .A(n21201), .B(p_input[5587]), .Z(n21203) );
  XOR U20793 ( .A(n21205), .B(n21206), .Z(n21201) );
  AND U20794 ( .A(n21207), .B(n21208), .Z(n21206) );
  XNOR U20795 ( .A(p_input[5618]), .B(n21205), .Z(n21208) );
  XOR U20796 ( .A(n21205), .B(p_input[5586]), .Z(n21207) );
  XOR U20797 ( .A(n21209), .B(n21210), .Z(n21205) );
  AND U20798 ( .A(n21211), .B(n21212), .Z(n21210) );
  XNOR U20799 ( .A(p_input[5617]), .B(n21209), .Z(n21212) );
  XOR U20800 ( .A(n21209), .B(p_input[5585]), .Z(n21211) );
  XOR U20801 ( .A(n21213), .B(n21214), .Z(n21209) );
  AND U20802 ( .A(n21215), .B(n21216), .Z(n21214) );
  XNOR U20803 ( .A(p_input[5616]), .B(n21213), .Z(n21216) );
  XOR U20804 ( .A(n21213), .B(p_input[5584]), .Z(n21215) );
  XOR U20805 ( .A(n21217), .B(n21218), .Z(n21213) );
  AND U20806 ( .A(n21219), .B(n21220), .Z(n21218) );
  XNOR U20807 ( .A(p_input[5615]), .B(n21217), .Z(n21220) );
  XOR U20808 ( .A(n21217), .B(p_input[5583]), .Z(n21219) );
  XOR U20809 ( .A(n21221), .B(n21222), .Z(n21217) );
  AND U20810 ( .A(n21223), .B(n21224), .Z(n21222) );
  XNOR U20811 ( .A(p_input[5614]), .B(n21221), .Z(n21224) );
  XOR U20812 ( .A(n21221), .B(p_input[5582]), .Z(n21223) );
  XOR U20813 ( .A(n21225), .B(n21226), .Z(n21221) );
  AND U20814 ( .A(n21227), .B(n21228), .Z(n21226) );
  XNOR U20815 ( .A(p_input[5613]), .B(n21225), .Z(n21228) );
  XOR U20816 ( .A(n21225), .B(p_input[5581]), .Z(n21227) );
  XOR U20817 ( .A(n21229), .B(n21230), .Z(n21225) );
  AND U20818 ( .A(n21231), .B(n21232), .Z(n21230) );
  XNOR U20819 ( .A(p_input[5612]), .B(n21229), .Z(n21232) );
  XOR U20820 ( .A(n21229), .B(p_input[5580]), .Z(n21231) );
  XOR U20821 ( .A(n21233), .B(n21234), .Z(n21229) );
  AND U20822 ( .A(n21235), .B(n21236), .Z(n21234) );
  XNOR U20823 ( .A(p_input[5611]), .B(n21233), .Z(n21236) );
  XOR U20824 ( .A(n21233), .B(p_input[5579]), .Z(n21235) );
  XOR U20825 ( .A(n21237), .B(n21238), .Z(n21233) );
  AND U20826 ( .A(n21239), .B(n21240), .Z(n21238) );
  XNOR U20827 ( .A(p_input[5610]), .B(n21237), .Z(n21240) );
  XOR U20828 ( .A(n21237), .B(p_input[5578]), .Z(n21239) );
  XOR U20829 ( .A(n21241), .B(n21242), .Z(n21237) );
  AND U20830 ( .A(n21243), .B(n21244), .Z(n21242) );
  XNOR U20831 ( .A(p_input[5609]), .B(n21241), .Z(n21244) );
  XOR U20832 ( .A(n21241), .B(p_input[5577]), .Z(n21243) );
  XOR U20833 ( .A(n21245), .B(n21246), .Z(n21241) );
  AND U20834 ( .A(n21247), .B(n21248), .Z(n21246) );
  XNOR U20835 ( .A(p_input[5608]), .B(n21245), .Z(n21248) );
  XOR U20836 ( .A(n21245), .B(p_input[5576]), .Z(n21247) );
  XOR U20837 ( .A(n21249), .B(n21250), .Z(n21245) );
  AND U20838 ( .A(n21251), .B(n21252), .Z(n21250) );
  XNOR U20839 ( .A(p_input[5607]), .B(n21249), .Z(n21252) );
  XOR U20840 ( .A(n21249), .B(p_input[5575]), .Z(n21251) );
  XOR U20841 ( .A(n21253), .B(n21254), .Z(n21249) );
  AND U20842 ( .A(n21255), .B(n21256), .Z(n21254) );
  XNOR U20843 ( .A(p_input[5606]), .B(n21253), .Z(n21256) );
  XOR U20844 ( .A(n21253), .B(p_input[5574]), .Z(n21255) );
  XOR U20845 ( .A(n21257), .B(n21258), .Z(n21253) );
  AND U20846 ( .A(n21259), .B(n21260), .Z(n21258) );
  XNOR U20847 ( .A(p_input[5605]), .B(n21257), .Z(n21260) );
  XOR U20848 ( .A(n21257), .B(p_input[5573]), .Z(n21259) );
  XOR U20849 ( .A(n21261), .B(n21262), .Z(n21257) );
  AND U20850 ( .A(n21263), .B(n21264), .Z(n21262) );
  XNOR U20851 ( .A(p_input[5604]), .B(n21261), .Z(n21264) );
  XOR U20852 ( .A(n21261), .B(p_input[5572]), .Z(n21263) );
  XOR U20853 ( .A(n21265), .B(n21266), .Z(n21261) );
  AND U20854 ( .A(n21267), .B(n21268), .Z(n21266) );
  XNOR U20855 ( .A(p_input[5603]), .B(n21265), .Z(n21268) );
  XOR U20856 ( .A(n21265), .B(p_input[5571]), .Z(n21267) );
  XOR U20857 ( .A(n21269), .B(n21270), .Z(n21265) );
  AND U20858 ( .A(n21271), .B(n21272), .Z(n21270) );
  XNOR U20859 ( .A(p_input[5602]), .B(n21269), .Z(n21272) );
  XOR U20860 ( .A(n21269), .B(p_input[5570]), .Z(n21271) );
  XNOR U20861 ( .A(n21273), .B(n21274), .Z(n21269) );
  AND U20862 ( .A(n21275), .B(n21276), .Z(n21274) );
  XOR U20863 ( .A(p_input[5601]), .B(n21273), .Z(n21276) );
  XNOR U20864 ( .A(p_input[5569]), .B(n21273), .Z(n21275) );
  AND U20865 ( .A(p_input[5600]), .B(n21277), .Z(n21273) );
  IV U20866 ( .A(p_input[5568]), .Z(n21277) );
  XNOR U20867 ( .A(p_input[5504]), .B(n21278), .Z(n20871) );
  AND U20868 ( .A(n337), .B(n21279), .Z(n21278) );
  XOR U20869 ( .A(p_input[5536]), .B(p_input[5504]), .Z(n21279) );
  XOR U20870 ( .A(n21280), .B(n21281), .Z(n337) );
  AND U20871 ( .A(n21282), .B(n21283), .Z(n21281) );
  XNOR U20872 ( .A(p_input[5567]), .B(n21280), .Z(n21283) );
  XOR U20873 ( .A(n21280), .B(p_input[5535]), .Z(n21282) );
  XOR U20874 ( .A(n21284), .B(n21285), .Z(n21280) );
  AND U20875 ( .A(n21286), .B(n21287), .Z(n21285) );
  XNOR U20876 ( .A(p_input[5566]), .B(n21284), .Z(n21287) );
  XNOR U20877 ( .A(n21284), .B(n20886), .Z(n21286) );
  IV U20878 ( .A(p_input[5534]), .Z(n20886) );
  XOR U20879 ( .A(n21288), .B(n21289), .Z(n21284) );
  AND U20880 ( .A(n21290), .B(n21291), .Z(n21289) );
  XNOR U20881 ( .A(p_input[5565]), .B(n21288), .Z(n21291) );
  XNOR U20882 ( .A(n21288), .B(n20895), .Z(n21290) );
  IV U20883 ( .A(p_input[5533]), .Z(n20895) );
  XOR U20884 ( .A(n21292), .B(n21293), .Z(n21288) );
  AND U20885 ( .A(n21294), .B(n21295), .Z(n21293) );
  XNOR U20886 ( .A(p_input[5564]), .B(n21292), .Z(n21295) );
  XNOR U20887 ( .A(n21292), .B(n20904), .Z(n21294) );
  IV U20888 ( .A(p_input[5532]), .Z(n20904) );
  XOR U20889 ( .A(n21296), .B(n21297), .Z(n21292) );
  AND U20890 ( .A(n21298), .B(n21299), .Z(n21297) );
  XNOR U20891 ( .A(p_input[5563]), .B(n21296), .Z(n21299) );
  XNOR U20892 ( .A(n21296), .B(n20913), .Z(n21298) );
  IV U20893 ( .A(p_input[5531]), .Z(n20913) );
  XOR U20894 ( .A(n21300), .B(n21301), .Z(n21296) );
  AND U20895 ( .A(n21302), .B(n21303), .Z(n21301) );
  XNOR U20896 ( .A(p_input[5562]), .B(n21300), .Z(n21303) );
  XNOR U20897 ( .A(n21300), .B(n20922), .Z(n21302) );
  IV U20898 ( .A(p_input[5530]), .Z(n20922) );
  XOR U20899 ( .A(n21304), .B(n21305), .Z(n21300) );
  AND U20900 ( .A(n21306), .B(n21307), .Z(n21305) );
  XNOR U20901 ( .A(p_input[5561]), .B(n21304), .Z(n21307) );
  XNOR U20902 ( .A(n21304), .B(n20931), .Z(n21306) );
  IV U20903 ( .A(p_input[5529]), .Z(n20931) );
  XOR U20904 ( .A(n21308), .B(n21309), .Z(n21304) );
  AND U20905 ( .A(n21310), .B(n21311), .Z(n21309) );
  XNOR U20906 ( .A(p_input[5560]), .B(n21308), .Z(n21311) );
  XNOR U20907 ( .A(n21308), .B(n20940), .Z(n21310) );
  IV U20908 ( .A(p_input[5528]), .Z(n20940) );
  XOR U20909 ( .A(n21312), .B(n21313), .Z(n21308) );
  AND U20910 ( .A(n21314), .B(n21315), .Z(n21313) );
  XNOR U20911 ( .A(p_input[5559]), .B(n21312), .Z(n21315) );
  XNOR U20912 ( .A(n21312), .B(n20949), .Z(n21314) );
  IV U20913 ( .A(p_input[5527]), .Z(n20949) );
  XOR U20914 ( .A(n21316), .B(n21317), .Z(n21312) );
  AND U20915 ( .A(n21318), .B(n21319), .Z(n21317) );
  XNOR U20916 ( .A(p_input[5558]), .B(n21316), .Z(n21319) );
  XNOR U20917 ( .A(n21316), .B(n20958), .Z(n21318) );
  IV U20918 ( .A(p_input[5526]), .Z(n20958) );
  XOR U20919 ( .A(n21320), .B(n21321), .Z(n21316) );
  AND U20920 ( .A(n21322), .B(n21323), .Z(n21321) );
  XNOR U20921 ( .A(p_input[5557]), .B(n21320), .Z(n21323) );
  XNOR U20922 ( .A(n21320), .B(n20967), .Z(n21322) );
  IV U20923 ( .A(p_input[5525]), .Z(n20967) );
  XOR U20924 ( .A(n21324), .B(n21325), .Z(n21320) );
  AND U20925 ( .A(n21326), .B(n21327), .Z(n21325) );
  XNOR U20926 ( .A(p_input[5556]), .B(n21324), .Z(n21327) );
  XNOR U20927 ( .A(n21324), .B(n20976), .Z(n21326) );
  IV U20928 ( .A(p_input[5524]), .Z(n20976) );
  XOR U20929 ( .A(n21328), .B(n21329), .Z(n21324) );
  AND U20930 ( .A(n21330), .B(n21331), .Z(n21329) );
  XNOR U20931 ( .A(p_input[5555]), .B(n21328), .Z(n21331) );
  XNOR U20932 ( .A(n21328), .B(n20985), .Z(n21330) );
  IV U20933 ( .A(p_input[5523]), .Z(n20985) );
  XOR U20934 ( .A(n21332), .B(n21333), .Z(n21328) );
  AND U20935 ( .A(n21334), .B(n21335), .Z(n21333) );
  XNOR U20936 ( .A(p_input[5554]), .B(n21332), .Z(n21335) );
  XNOR U20937 ( .A(n21332), .B(n20994), .Z(n21334) );
  IV U20938 ( .A(p_input[5522]), .Z(n20994) );
  XOR U20939 ( .A(n21336), .B(n21337), .Z(n21332) );
  AND U20940 ( .A(n21338), .B(n21339), .Z(n21337) );
  XNOR U20941 ( .A(p_input[5553]), .B(n21336), .Z(n21339) );
  XNOR U20942 ( .A(n21336), .B(n21003), .Z(n21338) );
  IV U20943 ( .A(p_input[5521]), .Z(n21003) );
  XOR U20944 ( .A(n21340), .B(n21341), .Z(n21336) );
  AND U20945 ( .A(n21342), .B(n21343), .Z(n21341) );
  XNOR U20946 ( .A(p_input[5552]), .B(n21340), .Z(n21343) );
  XNOR U20947 ( .A(n21340), .B(n21012), .Z(n21342) );
  IV U20948 ( .A(p_input[5520]), .Z(n21012) );
  XOR U20949 ( .A(n21344), .B(n21345), .Z(n21340) );
  AND U20950 ( .A(n21346), .B(n21347), .Z(n21345) );
  XNOR U20951 ( .A(p_input[5551]), .B(n21344), .Z(n21347) );
  XNOR U20952 ( .A(n21344), .B(n21021), .Z(n21346) );
  IV U20953 ( .A(p_input[5519]), .Z(n21021) );
  XOR U20954 ( .A(n21348), .B(n21349), .Z(n21344) );
  AND U20955 ( .A(n21350), .B(n21351), .Z(n21349) );
  XNOR U20956 ( .A(p_input[5550]), .B(n21348), .Z(n21351) );
  XNOR U20957 ( .A(n21348), .B(n21030), .Z(n21350) );
  IV U20958 ( .A(p_input[5518]), .Z(n21030) );
  XOR U20959 ( .A(n21352), .B(n21353), .Z(n21348) );
  AND U20960 ( .A(n21354), .B(n21355), .Z(n21353) );
  XNOR U20961 ( .A(p_input[5549]), .B(n21352), .Z(n21355) );
  XNOR U20962 ( .A(n21352), .B(n21039), .Z(n21354) );
  IV U20963 ( .A(p_input[5517]), .Z(n21039) );
  XOR U20964 ( .A(n21356), .B(n21357), .Z(n21352) );
  AND U20965 ( .A(n21358), .B(n21359), .Z(n21357) );
  XNOR U20966 ( .A(p_input[5548]), .B(n21356), .Z(n21359) );
  XNOR U20967 ( .A(n21356), .B(n21048), .Z(n21358) );
  IV U20968 ( .A(p_input[5516]), .Z(n21048) );
  XOR U20969 ( .A(n21360), .B(n21361), .Z(n21356) );
  AND U20970 ( .A(n21362), .B(n21363), .Z(n21361) );
  XNOR U20971 ( .A(p_input[5547]), .B(n21360), .Z(n21363) );
  XNOR U20972 ( .A(n21360), .B(n21057), .Z(n21362) );
  IV U20973 ( .A(p_input[5515]), .Z(n21057) );
  XOR U20974 ( .A(n21364), .B(n21365), .Z(n21360) );
  AND U20975 ( .A(n21366), .B(n21367), .Z(n21365) );
  XNOR U20976 ( .A(p_input[5546]), .B(n21364), .Z(n21367) );
  XNOR U20977 ( .A(n21364), .B(n21066), .Z(n21366) );
  IV U20978 ( .A(p_input[5514]), .Z(n21066) );
  XOR U20979 ( .A(n21368), .B(n21369), .Z(n21364) );
  AND U20980 ( .A(n21370), .B(n21371), .Z(n21369) );
  XNOR U20981 ( .A(p_input[5545]), .B(n21368), .Z(n21371) );
  XNOR U20982 ( .A(n21368), .B(n21075), .Z(n21370) );
  IV U20983 ( .A(p_input[5513]), .Z(n21075) );
  XOR U20984 ( .A(n21372), .B(n21373), .Z(n21368) );
  AND U20985 ( .A(n21374), .B(n21375), .Z(n21373) );
  XNOR U20986 ( .A(p_input[5544]), .B(n21372), .Z(n21375) );
  XNOR U20987 ( .A(n21372), .B(n21084), .Z(n21374) );
  IV U20988 ( .A(p_input[5512]), .Z(n21084) );
  XOR U20989 ( .A(n21376), .B(n21377), .Z(n21372) );
  AND U20990 ( .A(n21378), .B(n21379), .Z(n21377) );
  XNOR U20991 ( .A(p_input[5543]), .B(n21376), .Z(n21379) );
  XNOR U20992 ( .A(n21376), .B(n21093), .Z(n21378) );
  IV U20993 ( .A(p_input[5511]), .Z(n21093) );
  XOR U20994 ( .A(n21380), .B(n21381), .Z(n21376) );
  AND U20995 ( .A(n21382), .B(n21383), .Z(n21381) );
  XNOR U20996 ( .A(p_input[5542]), .B(n21380), .Z(n21383) );
  XNOR U20997 ( .A(n21380), .B(n21102), .Z(n21382) );
  IV U20998 ( .A(p_input[5510]), .Z(n21102) );
  XOR U20999 ( .A(n21384), .B(n21385), .Z(n21380) );
  AND U21000 ( .A(n21386), .B(n21387), .Z(n21385) );
  XNOR U21001 ( .A(p_input[5541]), .B(n21384), .Z(n21387) );
  XNOR U21002 ( .A(n21384), .B(n21111), .Z(n21386) );
  IV U21003 ( .A(p_input[5509]), .Z(n21111) );
  XOR U21004 ( .A(n21388), .B(n21389), .Z(n21384) );
  AND U21005 ( .A(n21390), .B(n21391), .Z(n21389) );
  XNOR U21006 ( .A(p_input[5540]), .B(n21388), .Z(n21391) );
  XNOR U21007 ( .A(n21388), .B(n21120), .Z(n21390) );
  IV U21008 ( .A(p_input[5508]), .Z(n21120) );
  XOR U21009 ( .A(n21392), .B(n21393), .Z(n21388) );
  AND U21010 ( .A(n21394), .B(n21395), .Z(n21393) );
  XNOR U21011 ( .A(p_input[5539]), .B(n21392), .Z(n21395) );
  XNOR U21012 ( .A(n21392), .B(n21129), .Z(n21394) );
  IV U21013 ( .A(p_input[5507]), .Z(n21129) );
  XOR U21014 ( .A(n21396), .B(n21397), .Z(n21392) );
  AND U21015 ( .A(n21398), .B(n21399), .Z(n21397) );
  XNOR U21016 ( .A(p_input[5538]), .B(n21396), .Z(n21399) );
  XNOR U21017 ( .A(n21396), .B(n21138), .Z(n21398) );
  IV U21018 ( .A(p_input[5506]), .Z(n21138) );
  XNOR U21019 ( .A(n21400), .B(n21401), .Z(n21396) );
  AND U21020 ( .A(n21402), .B(n21403), .Z(n21401) );
  XOR U21021 ( .A(p_input[5537]), .B(n21400), .Z(n21403) );
  XNOR U21022 ( .A(p_input[5505]), .B(n21400), .Z(n21402) );
  AND U21023 ( .A(p_input[5536]), .B(n21404), .Z(n21400) );
  IV U21024 ( .A(p_input[5504]), .Z(n21404) );
  XOR U21025 ( .A(n21405), .B(n21406), .Z(n20494) );
  AND U21026 ( .A(n509), .B(n21407), .Z(n21406) );
  XNOR U21027 ( .A(n21408), .B(n21405), .Z(n21407) );
  XOR U21028 ( .A(n21409), .B(n21410), .Z(n509) );
  AND U21029 ( .A(n21411), .B(n21412), .Z(n21410) );
  XNOR U21030 ( .A(n20509), .B(n21409), .Z(n21412) );
  AND U21031 ( .A(p_input[5503]), .B(p_input[5471]), .Z(n20509) );
  XNOR U21032 ( .A(n21409), .B(n20506), .Z(n21411) );
  IV U21033 ( .A(n21413), .Z(n20506) );
  AND U21034 ( .A(p_input[5407]), .B(p_input[5439]), .Z(n21413) );
  XOR U21035 ( .A(n21414), .B(n21415), .Z(n21409) );
  AND U21036 ( .A(n21416), .B(n21417), .Z(n21415) );
  XOR U21037 ( .A(n21414), .B(n20521), .Z(n21417) );
  XNOR U21038 ( .A(p_input[5470]), .B(n21418), .Z(n20521) );
  AND U21039 ( .A(n343), .B(n21419), .Z(n21418) );
  XOR U21040 ( .A(p_input[5502]), .B(p_input[5470]), .Z(n21419) );
  XNOR U21041 ( .A(n20518), .B(n21414), .Z(n21416) );
  XOR U21042 ( .A(n21420), .B(n21421), .Z(n20518) );
  AND U21043 ( .A(n340), .B(n21422), .Z(n21421) );
  XOR U21044 ( .A(p_input[5438]), .B(p_input[5406]), .Z(n21422) );
  XOR U21045 ( .A(n21423), .B(n21424), .Z(n21414) );
  AND U21046 ( .A(n21425), .B(n21426), .Z(n21424) );
  XOR U21047 ( .A(n21423), .B(n20533), .Z(n21426) );
  XNOR U21048 ( .A(p_input[5469]), .B(n21427), .Z(n20533) );
  AND U21049 ( .A(n343), .B(n21428), .Z(n21427) );
  XOR U21050 ( .A(p_input[5501]), .B(p_input[5469]), .Z(n21428) );
  XNOR U21051 ( .A(n20530), .B(n21423), .Z(n21425) );
  XOR U21052 ( .A(n21429), .B(n21430), .Z(n20530) );
  AND U21053 ( .A(n340), .B(n21431), .Z(n21430) );
  XOR U21054 ( .A(p_input[5437]), .B(p_input[5405]), .Z(n21431) );
  XOR U21055 ( .A(n21432), .B(n21433), .Z(n21423) );
  AND U21056 ( .A(n21434), .B(n21435), .Z(n21433) );
  XOR U21057 ( .A(n21432), .B(n20545), .Z(n21435) );
  XNOR U21058 ( .A(p_input[5468]), .B(n21436), .Z(n20545) );
  AND U21059 ( .A(n343), .B(n21437), .Z(n21436) );
  XOR U21060 ( .A(p_input[5500]), .B(p_input[5468]), .Z(n21437) );
  XNOR U21061 ( .A(n20542), .B(n21432), .Z(n21434) );
  XOR U21062 ( .A(n21438), .B(n21439), .Z(n20542) );
  AND U21063 ( .A(n340), .B(n21440), .Z(n21439) );
  XOR U21064 ( .A(p_input[5436]), .B(p_input[5404]), .Z(n21440) );
  XOR U21065 ( .A(n21441), .B(n21442), .Z(n21432) );
  AND U21066 ( .A(n21443), .B(n21444), .Z(n21442) );
  XOR U21067 ( .A(n21441), .B(n20557), .Z(n21444) );
  XNOR U21068 ( .A(p_input[5467]), .B(n21445), .Z(n20557) );
  AND U21069 ( .A(n343), .B(n21446), .Z(n21445) );
  XOR U21070 ( .A(p_input[5499]), .B(p_input[5467]), .Z(n21446) );
  XNOR U21071 ( .A(n20554), .B(n21441), .Z(n21443) );
  XOR U21072 ( .A(n21447), .B(n21448), .Z(n20554) );
  AND U21073 ( .A(n340), .B(n21449), .Z(n21448) );
  XOR U21074 ( .A(p_input[5435]), .B(p_input[5403]), .Z(n21449) );
  XOR U21075 ( .A(n21450), .B(n21451), .Z(n21441) );
  AND U21076 ( .A(n21452), .B(n21453), .Z(n21451) );
  XOR U21077 ( .A(n21450), .B(n20569), .Z(n21453) );
  XNOR U21078 ( .A(p_input[5466]), .B(n21454), .Z(n20569) );
  AND U21079 ( .A(n343), .B(n21455), .Z(n21454) );
  XOR U21080 ( .A(p_input[5498]), .B(p_input[5466]), .Z(n21455) );
  XNOR U21081 ( .A(n20566), .B(n21450), .Z(n21452) );
  XOR U21082 ( .A(n21456), .B(n21457), .Z(n20566) );
  AND U21083 ( .A(n340), .B(n21458), .Z(n21457) );
  XOR U21084 ( .A(p_input[5434]), .B(p_input[5402]), .Z(n21458) );
  XOR U21085 ( .A(n21459), .B(n21460), .Z(n21450) );
  AND U21086 ( .A(n21461), .B(n21462), .Z(n21460) );
  XOR U21087 ( .A(n21459), .B(n20581), .Z(n21462) );
  XNOR U21088 ( .A(p_input[5465]), .B(n21463), .Z(n20581) );
  AND U21089 ( .A(n343), .B(n21464), .Z(n21463) );
  XOR U21090 ( .A(p_input[5497]), .B(p_input[5465]), .Z(n21464) );
  XNOR U21091 ( .A(n20578), .B(n21459), .Z(n21461) );
  XOR U21092 ( .A(n21465), .B(n21466), .Z(n20578) );
  AND U21093 ( .A(n340), .B(n21467), .Z(n21466) );
  XOR U21094 ( .A(p_input[5433]), .B(p_input[5401]), .Z(n21467) );
  XOR U21095 ( .A(n21468), .B(n21469), .Z(n21459) );
  AND U21096 ( .A(n21470), .B(n21471), .Z(n21469) );
  XOR U21097 ( .A(n21468), .B(n20593), .Z(n21471) );
  XNOR U21098 ( .A(p_input[5464]), .B(n21472), .Z(n20593) );
  AND U21099 ( .A(n343), .B(n21473), .Z(n21472) );
  XOR U21100 ( .A(p_input[5496]), .B(p_input[5464]), .Z(n21473) );
  XNOR U21101 ( .A(n20590), .B(n21468), .Z(n21470) );
  XOR U21102 ( .A(n21474), .B(n21475), .Z(n20590) );
  AND U21103 ( .A(n340), .B(n21476), .Z(n21475) );
  XOR U21104 ( .A(p_input[5432]), .B(p_input[5400]), .Z(n21476) );
  XOR U21105 ( .A(n21477), .B(n21478), .Z(n21468) );
  AND U21106 ( .A(n21479), .B(n21480), .Z(n21478) );
  XOR U21107 ( .A(n21477), .B(n20605), .Z(n21480) );
  XNOR U21108 ( .A(p_input[5463]), .B(n21481), .Z(n20605) );
  AND U21109 ( .A(n343), .B(n21482), .Z(n21481) );
  XOR U21110 ( .A(p_input[5495]), .B(p_input[5463]), .Z(n21482) );
  XNOR U21111 ( .A(n20602), .B(n21477), .Z(n21479) );
  XOR U21112 ( .A(n21483), .B(n21484), .Z(n20602) );
  AND U21113 ( .A(n340), .B(n21485), .Z(n21484) );
  XOR U21114 ( .A(p_input[5431]), .B(p_input[5399]), .Z(n21485) );
  XOR U21115 ( .A(n21486), .B(n21487), .Z(n21477) );
  AND U21116 ( .A(n21488), .B(n21489), .Z(n21487) );
  XOR U21117 ( .A(n21486), .B(n20617), .Z(n21489) );
  XNOR U21118 ( .A(p_input[5462]), .B(n21490), .Z(n20617) );
  AND U21119 ( .A(n343), .B(n21491), .Z(n21490) );
  XOR U21120 ( .A(p_input[5494]), .B(p_input[5462]), .Z(n21491) );
  XNOR U21121 ( .A(n20614), .B(n21486), .Z(n21488) );
  XOR U21122 ( .A(n21492), .B(n21493), .Z(n20614) );
  AND U21123 ( .A(n340), .B(n21494), .Z(n21493) );
  XOR U21124 ( .A(p_input[5430]), .B(p_input[5398]), .Z(n21494) );
  XOR U21125 ( .A(n21495), .B(n21496), .Z(n21486) );
  AND U21126 ( .A(n21497), .B(n21498), .Z(n21496) );
  XOR U21127 ( .A(n21495), .B(n20629), .Z(n21498) );
  XNOR U21128 ( .A(p_input[5461]), .B(n21499), .Z(n20629) );
  AND U21129 ( .A(n343), .B(n21500), .Z(n21499) );
  XOR U21130 ( .A(p_input[5493]), .B(p_input[5461]), .Z(n21500) );
  XNOR U21131 ( .A(n20626), .B(n21495), .Z(n21497) );
  XOR U21132 ( .A(n21501), .B(n21502), .Z(n20626) );
  AND U21133 ( .A(n340), .B(n21503), .Z(n21502) );
  XOR U21134 ( .A(p_input[5429]), .B(p_input[5397]), .Z(n21503) );
  XOR U21135 ( .A(n21504), .B(n21505), .Z(n21495) );
  AND U21136 ( .A(n21506), .B(n21507), .Z(n21505) );
  XOR U21137 ( .A(n21504), .B(n20641), .Z(n21507) );
  XNOR U21138 ( .A(p_input[5460]), .B(n21508), .Z(n20641) );
  AND U21139 ( .A(n343), .B(n21509), .Z(n21508) );
  XOR U21140 ( .A(p_input[5492]), .B(p_input[5460]), .Z(n21509) );
  XNOR U21141 ( .A(n20638), .B(n21504), .Z(n21506) );
  XOR U21142 ( .A(n21510), .B(n21511), .Z(n20638) );
  AND U21143 ( .A(n340), .B(n21512), .Z(n21511) );
  XOR U21144 ( .A(p_input[5428]), .B(p_input[5396]), .Z(n21512) );
  XOR U21145 ( .A(n21513), .B(n21514), .Z(n21504) );
  AND U21146 ( .A(n21515), .B(n21516), .Z(n21514) );
  XOR U21147 ( .A(n21513), .B(n20653), .Z(n21516) );
  XNOR U21148 ( .A(p_input[5459]), .B(n21517), .Z(n20653) );
  AND U21149 ( .A(n343), .B(n21518), .Z(n21517) );
  XOR U21150 ( .A(p_input[5491]), .B(p_input[5459]), .Z(n21518) );
  XNOR U21151 ( .A(n20650), .B(n21513), .Z(n21515) );
  XOR U21152 ( .A(n21519), .B(n21520), .Z(n20650) );
  AND U21153 ( .A(n340), .B(n21521), .Z(n21520) );
  XOR U21154 ( .A(p_input[5427]), .B(p_input[5395]), .Z(n21521) );
  XOR U21155 ( .A(n21522), .B(n21523), .Z(n21513) );
  AND U21156 ( .A(n21524), .B(n21525), .Z(n21523) );
  XOR U21157 ( .A(n21522), .B(n20665), .Z(n21525) );
  XNOR U21158 ( .A(p_input[5458]), .B(n21526), .Z(n20665) );
  AND U21159 ( .A(n343), .B(n21527), .Z(n21526) );
  XOR U21160 ( .A(p_input[5490]), .B(p_input[5458]), .Z(n21527) );
  XNOR U21161 ( .A(n20662), .B(n21522), .Z(n21524) );
  XOR U21162 ( .A(n21528), .B(n21529), .Z(n20662) );
  AND U21163 ( .A(n340), .B(n21530), .Z(n21529) );
  XOR U21164 ( .A(p_input[5426]), .B(p_input[5394]), .Z(n21530) );
  XOR U21165 ( .A(n21531), .B(n21532), .Z(n21522) );
  AND U21166 ( .A(n21533), .B(n21534), .Z(n21532) );
  XOR U21167 ( .A(n21531), .B(n20677), .Z(n21534) );
  XNOR U21168 ( .A(p_input[5457]), .B(n21535), .Z(n20677) );
  AND U21169 ( .A(n343), .B(n21536), .Z(n21535) );
  XOR U21170 ( .A(p_input[5489]), .B(p_input[5457]), .Z(n21536) );
  XNOR U21171 ( .A(n20674), .B(n21531), .Z(n21533) );
  XOR U21172 ( .A(n21537), .B(n21538), .Z(n20674) );
  AND U21173 ( .A(n340), .B(n21539), .Z(n21538) );
  XOR U21174 ( .A(p_input[5425]), .B(p_input[5393]), .Z(n21539) );
  XOR U21175 ( .A(n21540), .B(n21541), .Z(n21531) );
  AND U21176 ( .A(n21542), .B(n21543), .Z(n21541) );
  XOR U21177 ( .A(n21540), .B(n20689), .Z(n21543) );
  XNOR U21178 ( .A(p_input[5456]), .B(n21544), .Z(n20689) );
  AND U21179 ( .A(n343), .B(n21545), .Z(n21544) );
  XOR U21180 ( .A(p_input[5488]), .B(p_input[5456]), .Z(n21545) );
  XNOR U21181 ( .A(n20686), .B(n21540), .Z(n21542) );
  XOR U21182 ( .A(n21546), .B(n21547), .Z(n20686) );
  AND U21183 ( .A(n340), .B(n21548), .Z(n21547) );
  XOR U21184 ( .A(p_input[5424]), .B(p_input[5392]), .Z(n21548) );
  XOR U21185 ( .A(n21549), .B(n21550), .Z(n21540) );
  AND U21186 ( .A(n21551), .B(n21552), .Z(n21550) );
  XOR U21187 ( .A(n21549), .B(n20701), .Z(n21552) );
  XNOR U21188 ( .A(p_input[5455]), .B(n21553), .Z(n20701) );
  AND U21189 ( .A(n343), .B(n21554), .Z(n21553) );
  XOR U21190 ( .A(p_input[5487]), .B(p_input[5455]), .Z(n21554) );
  XNOR U21191 ( .A(n20698), .B(n21549), .Z(n21551) );
  XOR U21192 ( .A(n21555), .B(n21556), .Z(n20698) );
  AND U21193 ( .A(n340), .B(n21557), .Z(n21556) );
  XOR U21194 ( .A(p_input[5423]), .B(p_input[5391]), .Z(n21557) );
  XOR U21195 ( .A(n21558), .B(n21559), .Z(n21549) );
  AND U21196 ( .A(n21560), .B(n21561), .Z(n21559) );
  XOR U21197 ( .A(n21558), .B(n20713), .Z(n21561) );
  XNOR U21198 ( .A(p_input[5454]), .B(n21562), .Z(n20713) );
  AND U21199 ( .A(n343), .B(n21563), .Z(n21562) );
  XOR U21200 ( .A(p_input[5486]), .B(p_input[5454]), .Z(n21563) );
  XNOR U21201 ( .A(n20710), .B(n21558), .Z(n21560) );
  XOR U21202 ( .A(n21564), .B(n21565), .Z(n20710) );
  AND U21203 ( .A(n340), .B(n21566), .Z(n21565) );
  XOR U21204 ( .A(p_input[5422]), .B(p_input[5390]), .Z(n21566) );
  XOR U21205 ( .A(n21567), .B(n21568), .Z(n21558) );
  AND U21206 ( .A(n21569), .B(n21570), .Z(n21568) );
  XOR U21207 ( .A(n21567), .B(n20725), .Z(n21570) );
  XNOR U21208 ( .A(p_input[5453]), .B(n21571), .Z(n20725) );
  AND U21209 ( .A(n343), .B(n21572), .Z(n21571) );
  XOR U21210 ( .A(p_input[5485]), .B(p_input[5453]), .Z(n21572) );
  XNOR U21211 ( .A(n20722), .B(n21567), .Z(n21569) );
  XOR U21212 ( .A(n21573), .B(n21574), .Z(n20722) );
  AND U21213 ( .A(n340), .B(n21575), .Z(n21574) );
  XOR U21214 ( .A(p_input[5421]), .B(p_input[5389]), .Z(n21575) );
  XOR U21215 ( .A(n21576), .B(n21577), .Z(n21567) );
  AND U21216 ( .A(n21578), .B(n21579), .Z(n21577) );
  XOR U21217 ( .A(n21576), .B(n20737), .Z(n21579) );
  XNOR U21218 ( .A(p_input[5452]), .B(n21580), .Z(n20737) );
  AND U21219 ( .A(n343), .B(n21581), .Z(n21580) );
  XOR U21220 ( .A(p_input[5484]), .B(p_input[5452]), .Z(n21581) );
  XNOR U21221 ( .A(n20734), .B(n21576), .Z(n21578) );
  XOR U21222 ( .A(n21582), .B(n21583), .Z(n20734) );
  AND U21223 ( .A(n340), .B(n21584), .Z(n21583) );
  XOR U21224 ( .A(p_input[5420]), .B(p_input[5388]), .Z(n21584) );
  XOR U21225 ( .A(n21585), .B(n21586), .Z(n21576) );
  AND U21226 ( .A(n21587), .B(n21588), .Z(n21586) );
  XOR U21227 ( .A(n21585), .B(n20749), .Z(n21588) );
  XNOR U21228 ( .A(p_input[5451]), .B(n21589), .Z(n20749) );
  AND U21229 ( .A(n343), .B(n21590), .Z(n21589) );
  XOR U21230 ( .A(p_input[5483]), .B(p_input[5451]), .Z(n21590) );
  XNOR U21231 ( .A(n20746), .B(n21585), .Z(n21587) );
  XOR U21232 ( .A(n21591), .B(n21592), .Z(n20746) );
  AND U21233 ( .A(n340), .B(n21593), .Z(n21592) );
  XOR U21234 ( .A(p_input[5419]), .B(p_input[5387]), .Z(n21593) );
  XOR U21235 ( .A(n21594), .B(n21595), .Z(n21585) );
  AND U21236 ( .A(n21596), .B(n21597), .Z(n21595) );
  XOR U21237 ( .A(n21594), .B(n20761), .Z(n21597) );
  XNOR U21238 ( .A(p_input[5450]), .B(n21598), .Z(n20761) );
  AND U21239 ( .A(n343), .B(n21599), .Z(n21598) );
  XOR U21240 ( .A(p_input[5482]), .B(p_input[5450]), .Z(n21599) );
  XNOR U21241 ( .A(n20758), .B(n21594), .Z(n21596) );
  XOR U21242 ( .A(n21600), .B(n21601), .Z(n20758) );
  AND U21243 ( .A(n340), .B(n21602), .Z(n21601) );
  XOR U21244 ( .A(p_input[5418]), .B(p_input[5386]), .Z(n21602) );
  XOR U21245 ( .A(n21603), .B(n21604), .Z(n21594) );
  AND U21246 ( .A(n21605), .B(n21606), .Z(n21604) );
  XOR U21247 ( .A(n21603), .B(n20773), .Z(n21606) );
  XNOR U21248 ( .A(p_input[5449]), .B(n21607), .Z(n20773) );
  AND U21249 ( .A(n343), .B(n21608), .Z(n21607) );
  XOR U21250 ( .A(p_input[5481]), .B(p_input[5449]), .Z(n21608) );
  XNOR U21251 ( .A(n20770), .B(n21603), .Z(n21605) );
  XOR U21252 ( .A(n21609), .B(n21610), .Z(n20770) );
  AND U21253 ( .A(n340), .B(n21611), .Z(n21610) );
  XOR U21254 ( .A(p_input[5417]), .B(p_input[5385]), .Z(n21611) );
  XOR U21255 ( .A(n21612), .B(n21613), .Z(n21603) );
  AND U21256 ( .A(n21614), .B(n21615), .Z(n21613) );
  XOR U21257 ( .A(n21612), .B(n20785), .Z(n21615) );
  XNOR U21258 ( .A(p_input[5448]), .B(n21616), .Z(n20785) );
  AND U21259 ( .A(n343), .B(n21617), .Z(n21616) );
  XOR U21260 ( .A(p_input[5480]), .B(p_input[5448]), .Z(n21617) );
  XNOR U21261 ( .A(n20782), .B(n21612), .Z(n21614) );
  XOR U21262 ( .A(n21618), .B(n21619), .Z(n20782) );
  AND U21263 ( .A(n340), .B(n21620), .Z(n21619) );
  XOR U21264 ( .A(p_input[5416]), .B(p_input[5384]), .Z(n21620) );
  XOR U21265 ( .A(n21621), .B(n21622), .Z(n21612) );
  AND U21266 ( .A(n21623), .B(n21624), .Z(n21622) );
  XOR U21267 ( .A(n21621), .B(n20797), .Z(n21624) );
  XNOR U21268 ( .A(p_input[5447]), .B(n21625), .Z(n20797) );
  AND U21269 ( .A(n343), .B(n21626), .Z(n21625) );
  XOR U21270 ( .A(p_input[5479]), .B(p_input[5447]), .Z(n21626) );
  XNOR U21271 ( .A(n20794), .B(n21621), .Z(n21623) );
  XOR U21272 ( .A(n21627), .B(n21628), .Z(n20794) );
  AND U21273 ( .A(n340), .B(n21629), .Z(n21628) );
  XOR U21274 ( .A(p_input[5415]), .B(p_input[5383]), .Z(n21629) );
  XOR U21275 ( .A(n21630), .B(n21631), .Z(n21621) );
  AND U21276 ( .A(n21632), .B(n21633), .Z(n21631) );
  XOR U21277 ( .A(n21630), .B(n20809), .Z(n21633) );
  XNOR U21278 ( .A(p_input[5446]), .B(n21634), .Z(n20809) );
  AND U21279 ( .A(n343), .B(n21635), .Z(n21634) );
  XOR U21280 ( .A(p_input[5478]), .B(p_input[5446]), .Z(n21635) );
  XNOR U21281 ( .A(n20806), .B(n21630), .Z(n21632) );
  XOR U21282 ( .A(n21636), .B(n21637), .Z(n20806) );
  AND U21283 ( .A(n340), .B(n21638), .Z(n21637) );
  XOR U21284 ( .A(p_input[5414]), .B(p_input[5382]), .Z(n21638) );
  XOR U21285 ( .A(n21639), .B(n21640), .Z(n21630) );
  AND U21286 ( .A(n21641), .B(n21642), .Z(n21640) );
  XOR U21287 ( .A(n21639), .B(n20821), .Z(n21642) );
  XNOR U21288 ( .A(p_input[5445]), .B(n21643), .Z(n20821) );
  AND U21289 ( .A(n343), .B(n21644), .Z(n21643) );
  XOR U21290 ( .A(p_input[5477]), .B(p_input[5445]), .Z(n21644) );
  XNOR U21291 ( .A(n20818), .B(n21639), .Z(n21641) );
  XOR U21292 ( .A(n21645), .B(n21646), .Z(n20818) );
  AND U21293 ( .A(n340), .B(n21647), .Z(n21646) );
  XOR U21294 ( .A(p_input[5413]), .B(p_input[5381]), .Z(n21647) );
  XOR U21295 ( .A(n21648), .B(n21649), .Z(n21639) );
  AND U21296 ( .A(n21650), .B(n21651), .Z(n21649) );
  XOR U21297 ( .A(n21648), .B(n20833), .Z(n21651) );
  XNOR U21298 ( .A(p_input[5444]), .B(n21652), .Z(n20833) );
  AND U21299 ( .A(n343), .B(n21653), .Z(n21652) );
  XOR U21300 ( .A(p_input[5476]), .B(p_input[5444]), .Z(n21653) );
  XNOR U21301 ( .A(n20830), .B(n21648), .Z(n21650) );
  XOR U21302 ( .A(n21654), .B(n21655), .Z(n20830) );
  AND U21303 ( .A(n340), .B(n21656), .Z(n21655) );
  XOR U21304 ( .A(p_input[5412]), .B(p_input[5380]), .Z(n21656) );
  XOR U21305 ( .A(n21657), .B(n21658), .Z(n21648) );
  AND U21306 ( .A(n21659), .B(n21660), .Z(n21658) );
  XOR U21307 ( .A(n21657), .B(n20845), .Z(n21660) );
  XNOR U21308 ( .A(p_input[5443]), .B(n21661), .Z(n20845) );
  AND U21309 ( .A(n343), .B(n21662), .Z(n21661) );
  XOR U21310 ( .A(p_input[5475]), .B(p_input[5443]), .Z(n21662) );
  XNOR U21311 ( .A(n20842), .B(n21657), .Z(n21659) );
  XOR U21312 ( .A(n21663), .B(n21664), .Z(n20842) );
  AND U21313 ( .A(n340), .B(n21665), .Z(n21664) );
  XOR U21314 ( .A(p_input[5411]), .B(p_input[5379]), .Z(n21665) );
  XOR U21315 ( .A(n21666), .B(n21667), .Z(n21657) );
  AND U21316 ( .A(n21668), .B(n21669), .Z(n21667) );
  XOR U21317 ( .A(n21666), .B(n20857), .Z(n21669) );
  XNOR U21318 ( .A(p_input[5442]), .B(n21670), .Z(n20857) );
  AND U21319 ( .A(n343), .B(n21671), .Z(n21670) );
  XOR U21320 ( .A(p_input[5474]), .B(p_input[5442]), .Z(n21671) );
  XNOR U21321 ( .A(n20854), .B(n21666), .Z(n21668) );
  XOR U21322 ( .A(n21672), .B(n21673), .Z(n20854) );
  AND U21323 ( .A(n340), .B(n21674), .Z(n21673) );
  XOR U21324 ( .A(p_input[5410]), .B(p_input[5378]), .Z(n21674) );
  XOR U21325 ( .A(n21675), .B(n21676), .Z(n21666) );
  AND U21326 ( .A(n21677), .B(n21678), .Z(n21676) );
  XNOR U21327 ( .A(n21679), .B(n20870), .Z(n21678) );
  XNOR U21328 ( .A(p_input[5441]), .B(n21680), .Z(n20870) );
  AND U21329 ( .A(n343), .B(n21681), .Z(n21680) );
  XNOR U21330 ( .A(p_input[5473]), .B(n21682), .Z(n21681) );
  IV U21331 ( .A(p_input[5441]), .Z(n21682) );
  XNOR U21332 ( .A(n20867), .B(n21675), .Z(n21677) );
  XNOR U21333 ( .A(p_input[5377]), .B(n21683), .Z(n20867) );
  AND U21334 ( .A(n340), .B(n21684), .Z(n21683) );
  XOR U21335 ( .A(p_input[5409]), .B(p_input[5377]), .Z(n21684) );
  IV U21336 ( .A(n21679), .Z(n21675) );
  AND U21337 ( .A(n21405), .B(n21408), .Z(n21679) );
  XOR U21338 ( .A(p_input[5440]), .B(n21685), .Z(n21408) );
  AND U21339 ( .A(n343), .B(n21686), .Z(n21685) );
  XOR U21340 ( .A(p_input[5472]), .B(p_input[5440]), .Z(n21686) );
  XOR U21341 ( .A(n21687), .B(n21688), .Z(n343) );
  AND U21342 ( .A(n21689), .B(n21690), .Z(n21688) );
  XNOR U21343 ( .A(p_input[5503]), .B(n21687), .Z(n21690) );
  XOR U21344 ( .A(n21687), .B(p_input[5471]), .Z(n21689) );
  XOR U21345 ( .A(n21691), .B(n21692), .Z(n21687) );
  AND U21346 ( .A(n21693), .B(n21694), .Z(n21692) );
  XNOR U21347 ( .A(p_input[5502]), .B(n21691), .Z(n21694) );
  XOR U21348 ( .A(n21691), .B(p_input[5470]), .Z(n21693) );
  XOR U21349 ( .A(n21695), .B(n21696), .Z(n21691) );
  AND U21350 ( .A(n21697), .B(n21698), .Z(n21696) );
  XNOR U21351 ( .A(p_input[5501]), .B(n21695), .Z(n21698) );
  XOR U21352 ( .A(n21695), .B(p_input[5469]), .Z(n21697) );
  XOR U21353 ( .A(n21699), .B(n21700), .Z(n21695) );
  AND U21354 ( .A(n21701), .B(n21702), .Z(n21700) );
  XNOR U21355 ( .A(p_input[5500]), .B(n21699), .Z(n21702) );
  XOR U21356 ( .A(n21699), .B(p_input[5468]), .Z(n21701) );
  XOR U21357 ( .A(n21703), .B(n21704), .Z(n21699) );
  AND U21358 ( .A(n21705), .B(n21706), .Z(n21704) );
  XNOR U21359 ( .A(p_input[5499]), .B(n21703), .Z(n21706) );
  XOR U21360 ( .A(n21703), .B(p_input[5467]), .Z(n21705) );
  XOR U21361 ( .A(n21707), .B(n21708), .Z(n21703) );
  AND U21362 ( .A(n21709), .B(n21710), .Z(n21708) );
  XNOR U21363 ( .A(p_input[5498]), .B(n21707), .Z(n21710) );
  XOR U21364 ( .A(n21707), .B(p_input[5466]), .Z(n21709) );
  XOR U21365 ( .A(n21711), .B(n21712), .Z(n21707) );
  AND U21366 ( .A(n21713), .B(n21714), .Z(n21712) );
  XNOR U21367 ( .A(p_input[5497]), .B(n21711), .Z(n21714) );
  XOR U21368 ( .A(n21711), .B(p_input[5465]), .Z(n21713) );
  XOR U21369 ( .A(n21715), .B(n21716), .Z(n21711) );
  AND U21370 ( .A(n21717), .B(n21718), .Z(n21716) );
  XNOR U21371 ( .A(p_input[5496]), .B(n21715), .Z(n21718) );
  XOR U21372 ( .A(n21715), .B(p_input[5464]), .Z(n21717) );
  XOR U21373 ( .A(n21719), .B(n21720), .Z(n21715) );
  AND U21374 ( .A(n21721), .B(n21722), .Z(n21720) );
  XNOR U21375 ( .A(p_input[5495]), .B(n21719), .Z(n21722) );
  XOR U21376 ( .A(n21719), .B(p_input[5463]), .Z(n21721) );
  XOR U21377 ( .A(n21723), .B(n21724), .Z(n21719) );
  AND U21378 ( .A(n21725), .B(n21726), .Z(n21724) );
  XNOR U21379 ( .A(p_input[5494]), .B(n21723), .Z(n21726) );
  XOR U21380 ( .A(n21723), .B(p_input[5462]), .Z(n21725) );
  XOR U21381 ( .A(n21727), .B(n21728), .Z(n21723) );
  AND U21382 ( .A(n21729), .B(n21730), .Z(n21728) );
  XNOR U21383 ( .A(p_input[5493]), .B(n21727), .Z(n21730) );
  XOR U21384 ( .A(n21727), .B(p_input[5461]), .Z(n21729) );
  XOR U21385 ( .A(n21731), .B(n21732), .Z(n21727) );
  AND U21386 ( .A(n21733), .B(n21734), .Z(n21732) );
  XNOR U21387 ( .A(p_input[5492]), .B(n21731), .Z(n21734) );
  XOR U21388 ( .A(n21731), .B(p_input[5460]), .Z(n21733) );
  XOR U21389 ( .A(n21735), .B(n21736), .Z(n21731) );
  AND U21390 ( .A(n21737), .B(n21738), .Z(n21736) );
  XNOR U21391 ( .A(p_input[5491]), .B(n21735), .Z(n21738) );
  XOR U21392 ( .A(n21735), .B(p_input[5459]), .Z(n21737) );
  XOR U21393 ( .A(n21739), .B(n21740), .Z(n21735) );
  AND U21394 ( .A(n21741), .B(n21742), .Z(n21740) );
  XNOR U21395 ( .A(p_input[5490]), .B(n21739), .Z(n21742) );
  XOR U21396 ( .A(n21739), .B(p_input[5458]), .Z(n21741) );
  XOR U21397 ( .A(n21743), .B(n21744), .Z(n21739) );
  AND U21398 ( .A(n21745), .B(n21746), .Z(n21744) );
  XNOR U21399 ( .A(p_input[5489]), .B(n21743), .Z(n21746) );
  XOR U21400 ( .A(n21743), .B(p_input[5457]), .Z(n21745) );
  XOR U21401 ( .A(n21747), .B(n21748), .Z(n21743) );
  AND U21402 ( .A(n21749), .B(n21750), .Z(n21748) );
  XNOR U21403 ( .A(p_input[5488]), .B(n21747), .Z(n21750) );
  XOR U21404 ( .A(n21747), .B(p_input[5456]), .Z(n21749) );
  XOR U21405 ( .A(n21751), .B(n21752), .Z(n21747) );
  AND U21406 ( .A(n21753), .B(n21754), .Z(n21752) );
  XNOR U21407 ( .A(p_input[5487]), .B(n21751), .Z(n21754) );
  XOR U21408 ( .A(n21751), .B(p_input[5455]), .Z(n21753) );
  XOR U21409 ( .A(n21755), .B(n21756), .Z(n21751) );
  AND U21410 ( .A(n21757), .B(n21758), .Z(n21756) );
  XNOR U21411 ( .A(p_input[5486]), .B(n21755), .Z(n21758) );
  XOR U21412 ( .A(n21755), .B(p_input[5454]), .Z(n21757) );
  XOR U21413 ( .A(n21759), .B(n21760), .Z(n21755) );
  AND U21414 ( .A(n21761), .B(n21762), .Z(n21760) );
  XNOR U21415 ( .A(p_input[5485]), .B(n21759), .Z(n21762) );
  XOR U21416 ( .A(n21759), .B(p_input[5453]), .Z(n21761) );
  XOR U21417 ( .A(n21763), .B(n21764), .Z(n21759) );
  AND U21418 ( .A(n21765), .B(n21766), .Z(n21764) );
  XNOR U21419 ( .A(p_input[5484]), .B(n21763), .Z(n21766) );
  XOR U21420 ( .A(n21763), .B(p_input[5452]), .Z(n21765) );
  XOR U21421 ( .A(n21767), .B(n21768), .Z(n21763) );
  AND U21422 ( .A(n21769), .B(n21770), .Z(n21768) );
  XNOR U21423 ( .A(p_input[5483]), .B(n21767), .Z(n21770) );
  XOR U21424 ( .A(n21767), .B(p_input[5451]), .Z(n21769) );
  XOR U21425 ( .A(n21771), .B(n21772), .Z(n21767) );
  AND U21426 ( .A(n21773), .B(n21774), .Z(n21772) );
  XNOR U21427 ( .A(p_input[5482]), .B(n21771), .Z(n21774) );
  XOR U21428 ( .A(n21771), .B(p_input[5450]), .Z(n21773) );
  XOR U21429 ( .A(n21775), .B(n21776), .Z(n21771) );
  AND U21430 ( .A(n21777), .B(n21778), .Z(n21776) );
  XNOR U21431 ( .A(p_input[5481]), .B(n21775), .Z(n21778) );
  XOR U21432 ( .A(n21775), .B(p_input[5449]), .Z(n21777) );
  XOR U21433 ( .A(n21779), .B(n21780), .Z(n21775) );
  AND U21434 ( .A(n21781), .B(n21782), .Z(n21780) );
  XNOR U21435 ( .A(p_input[5480]), .B(n21779), .Z(n21782) );
  XOR U21436 ( .A(n21779), .B(p_input[5448]), .Z(n21781) );
  XOR U21437 ( .A(n21783), .B(n21784), .Z(n21779) );
  AND U21438 ( .A(n21785), .B(n21786), .Z(n21784) );
  XNOR U21439 ( .A(p_input[5479]), .B(n21783), .Z(n21786) );
  XOR U21440 ( .A(n21783), .B(p_input[5447]), .Z(n21785) );
  XOR U21441 ( .A(n21787), .B(n21788), .Z(n21783) );
  AND U21442 ( .A(n21789), .B(n21790), .Z(n21788) );
  XNOR U21443 ( .A(p_input[5478]), .B(n21787), .Z(n21790) );
  XOR U21444 ( .A(n21787), .B(p_input[5446]), .Z(n21789) );
  XOR U21445 ( .A(n21791), .B(n21792), .Z(n21787) );
  AND U21446 ( .A(n21793), .B(n21794), .Z(n21792) );
  XNOR U21447 ( .A(p_input[5477]), .B(n21791), .Z(n21794) );
  XOR U21448 ( .A(n21791), .B(p_input[5445]), .Z(n21793) );
  XOR U21449 ( .A(n21795), .B(n21796), .Z(n21791) );
  AND U21450 ( .A(n21797), .B(n21798), .Z(n21796) );
  XNOR U21451 ( .A(p_input[5476]), .B(n21795), .Z(n21798) );
  XOR U21452 ( .A(n21795), .B(p_input[5444]), .Z(n21797) );
  XOR U21453 ( .A(n21799), .B(n21800), .Z(n21795) );
  AND U21454 ( .A(n21801), .B(n21802), .Z(n21800) );
  XNOR U21455 ( .A(p_input[5475]), .B(n21799), .Z(n21802) );
  XOR U21456 ( .A(n21799), .B(p_input[5443]), .Z(n21801) );
  XOR U21457 ( .A(n21803), .B(n21804), .Z(n21799) );
  AND U21458 ( .A(n21805), .B(n21806), .Z(n21804) );
  XNOR U21459 ( .A(p_input[5474]), .B(n21803), .Z(n21806) );
  XOR U21460 ( .A(n21803), .B(p_input[5442]), .Z(n21805) );
  XNOR U21461 ( .A(n21807), .B(n21808), .Z(n21803) );
  AND U21462 ( .A(n21809), .B(n21810), .Z(n21808) );
  XOR U21463 ( .A(p_input[5473]), .B(n21807), .Z(n21810) );
  XNOR U21464 ( .A(p_input[5441]), .B(n21807), .Z(n21809) );
  AND U21465 ( .A(p_input[5472]), .B(n21811), .Z(n21807) );
  IV U21466 ( .A(p_input[5440]), .Z(n21811) );
  XNOR U21467 ( .A(p_input[5376]), .B(n21812), .Z(n21405) );
  AND U21468 ( .A(n340), .B(n21813), .Z(n21812) );
  XOR U21469 ( .A(p_input[5408]), .B(p_input[5376]), .Z(n21813) );
  XOR U21470 ( .A(n21814), .B(n21815), .Z(n340) );
  AND U21471 ( .A(n21816), .B(n21817), .Z(n21815) );
  XNOR U21472 ( .A(p_input[5439]), .B(n21814), .Z(n21817) );
  XOR U21473 ( .A(n21814), .B(p_input[5407]), .Z(n21816) );
  XOR U21474 ( .A(n21818), .B(n21819), .Z(n21814) );
  AND U21475 ( .A(n21820), .B(n21821), .Z(n21819) );
  XNOR U21476 ( .A(p_input[5438]), .B(n21818), .Z(n21821) );
  XNOR U21477 ( .A(n21818), .B(n21420), .Z(n21820) );
  IV U21478 ( .A(p_input[5406]), .Z(n21420) );
  XOR U21479 ( .A(n21822), .B(n21823), .Z(n21818) );
  AND U21480 ( .A(n21824), .B(n21825), .Z(n21823) );
  XNOR U21481 ( .A(p_input[5437]), .B(n21822), .Z(n21825) );
  XNOR U21482 ( .A(n21822), .B(n21429), .Z(n21824) );
  IV U21483 ( .A(p_input[5405]), .Z(n21429) );
  XOR U21484 ( .A(n21826), .B(n21827), .Z(n21822) );
  AND U21485 ( .A(n21828), .B(n21829), .Z(n21827) );
  XNOR U21486 ( .A(p_input[5436]), .B(n21826), .Z(n21829) );
  XNOR U21487 ( .A(n21826), .B(n21438), .Z(n21828) );
  IV U21488 ( .A(p_input[5404]), .Z(n21438) );
  XOR U21489 ( .A(n21830), .B(n21831), .Z(n21826) );
  AND U21490 ( .A(n21832), .B(n21833), .Z(n21831) );
  XNOR U21491 ( .A(p_input[5435]), .B(n21830), .Z(n21833) );
  XNOR U21492 ( .A(n21830), .B(n21447), .Z(n21832) );
  IV U21493 ( .A(p_input[5403]), .Z(n21447) );
  XOR U21494 ( .A(n21834), .B(n21835), .Z(n21830) );
  AND U21495 ( .A(n21836), .B(n21837), .Z(n21835) );
  XNOR U21496 ( .A(p_input[5434]), .B(n21834), .Z(n21837) );
  XNOR U21497 ( .A(n21834), .B(n21456), .Z(n21836) );
  IV U21498 ( .A(p_input[5402]), .Z(n21456) );
  XOR U21499 ( .A(n21838), .B(n21839), .Z(n21834) );
  AND U21500 ( .A(n21840), .B(n21841), .Z(n21839) );
  XNOR U21501 ( .A(p_input[5433]), .B(n21838), .Z(n21841) );
  XNOR U21502 ( .A(n21838), .B(n21465), .Z(n21840) );
  IV U21503 ( .A(p_input[5401]), .Z(n21465) );
  XOR U21504 ( .A(n21842), .B(n21843), .Z(n21838) );
  AND U21505 ( .A(n21844), .B(n21845), .Z(n21843) );
  XNOR U21506 ( .A(p_input[5432]), .B(n21842), .Z(n21845) );
  XNOR U21507 ( .A(n21842), .B(n21474), .Z(n21844) );
  IV U21508 ( .A(p_input[5400]), .Z(n21474) );
  XOR U21509 ( .A(n21846), .B(n21847), .Z(n21842) );
  AND U21510 ( .A(n21848), .B(n21849), .Z(n21847) );
  XNOR U21511 ( .A(p_input[5431]), .B(n21846), .Z(n21849) );
  XNOR U21512 ( .A(n21846), .B(n21483), .Z(n21848) );
  IV U21513 ( .A(p_input[5399]), .Z(n21483) );
  XOR U21514 ( .A(n21850), .B(n21851), .Z(n21846) );
  AND U21515 ( .A(n21852), .B(n21853), .Z(n21851) );
  XNOR U21516 ( .A(p_input[5430]), .B(n21850), .Z(n21853) );
  XNOR U21517 ( .A(n21850), .B(n21492), .Z(n21852) );
  IV U21518 ( .A(p_input[5398]), .Z(n21492) );
  XOR U21519 ( .A(n21854), .B(n21855), .Z(n21850) );
  AND U21520 ( .A(n21856), .B(n21857), .Z(n21855) );
  XNOR U21521 ( .A(p_input[5429]), .B(n21854), .Z(n21857) );
  XNOR U21522 ( .A(n21854), .B(n21501), .Z(n21856) );
  IV U21523 ( .A(p_input[5397]), .Z(n21501) );
  XOR U21524 ( .A(n21858), .B(n21859), .Z(n21854) );
  AND U21525 ( .A(n21860), .B(n21861), .Z(n21859) );
  XNOR U21526 ( .A(p_input[5428]), .B(n21858), .Z(n21861) );
  XNOR U21527 ( .A(n21858), .B(n21510), .Z(n21860) );
  IV U21528 ( .A(p_input[5396]), .Z(n21510) );
  XOR U21529 ( .A(n21862), .B(n21863), .Z(n21858) );
  AND U21530 ( .A(n21864), .B(n21865), .Z(n21863) );
  XNOR U21531 ( .A(p_input[5427]), .B(n21862), .Z(n21865) );
  XNOR U21532 ( .A(n21862), .B(n21519), .Z(n21864) );
  IV U21533 ( .A(p_input[5395]), .Z(n21519) );
  XOR U21534 ( .A(n21866), .B(n21867), .Z(n21862) );
  AND U21535 ( .A(n21868), .B(n21869), .Z(n21867) );
  XNOR U21536 ( .A(p_input[5426]), .B(n21866), .Z(n21869) );
  XNOR U21537 ( .A(n21866), .B(n21528), .Z(n21868) );
  IV U21538 ( .A(p_input[5394]), .Z(n21528) );
  XOR U21539 ( .A(n21870), .B(n21871), .Z(n21866) );
  AND U21540 ( .A(n21872), .B(n21873), .Z(n21871) );
  XNOR U21541 ( .A(p_input[5425]), .B(n21870), .Z(n21873) );
  XNOR U21542 ( .A(n21870), .B(n21537), .Z(n21872) );
  IV U21543 ( .A(p_input[5393]), .Z(n21537) );
  XOR U21544 ( .A(n21874), .B(n21875), .Z(n21870) );
  AND U21545 ( .A(n21876), .B(n21877), .Z(n21875) );
  XNOR U21546 ( .A(p_input[5424]), .B(n21874), .Z(n21877) );
  XNOR U21547 ( .A(n21874), .B(n21546), .Z(n21876) );
  IV U21548 ( .A(p_input[5392]), .Z(n21546) );
  XOR U21549 ( .A(n21878), .B(n21879), .Z(n21874) );
  AND U21550 ( .A(n21880), .B(n21881), .Z(n21879) );
  XNOR U21551 ( .A(p_input[5423]), .B(n21878), .Z(n21881) );
  XNOR U21552 ( .A(n21878), .B(n21555), .Z(n21880) );
  IV U21553 ( .A(p_input[5391]), .Z(n21555) );
  XOR U21554 ( .A(n21882), .B(n21883), .Z(n21878) );
  AND U21555 ( .A(n21884), .B(n21885), .Z(n21883) );
  XNOR U21556 ( .A(p_input[5422]), .B(n21882), .Z(n21885) );
  XNOR U21557 ( .A(n21882), .B(n21564), .Z(n21884) );
  IV U21558 ( .A(p_input[5390]), .Z(n21564) );
  XOR U21559 ( .A(n21886), .B(n21887), .Z(n21882) );
  AND U21560 ( .A(n21888), .B(n21889), .Z(n21887) );
  XNOR U21561 ( .A(p_input[5421]), .B(n21886), .Z(n21889) );
  XNOR U21562 ( .A(n21886), .B(n21573), .Z(n21888) );
  IV U21563 ( .A(p_input[5389]), .Z(n21573) );
  XOR U21564 ( .A(n21890), .B(n21891), .Z(n21886) );
  AND U21565 ( .A(n21892), .B(n21893), .Z(n21891) );
  XNOR U21566 ( .A(p_input[5420]), .B(n21890), .Z(n21893) );
  XNOR U21567 ( .A(n21890), .B(n21582), .Z(n21892) );
  IV U21568 ( .A(p_input[5388]), .Z(n21582) );
  XOR U21569 ( .A(n21894), .B(n21895), .Z(n21890) );
  AND U21570 ( .A(n21896), .B(n21897), .Z(n21895) );
  XNOR U21571 ( .A(p_input[5419]), .B(n21894), .Z(n21897) );
  XNOR U21572 ( .A(n21894), .B(n21591), .Z(n21896) );
  IV U21573 ( .A(p_input[5387]), .Z(n21591) );
  XOR U21574 ( .A(n21898), .B(n21899), .Z(n21894) );
  AND U21575 ( .A(n21900), .B(n21901), .Z(n21899) );
  XNOR U21576 ( .A(p_input[5418]), .B(n21898), .Z(n21901) );
  XNOR U21577 ( .A(n21898), .B(n21600), .Z(n21900) );
  IV U21578 ( .A(p_input[5386]), .Z(n21600) );
  XOR U21579 ( .A(n21902), .B(n21903), .Z(n21898) );
  AND U21580 ( .A(n21904), .B(n21905), .Z(n21903) );
  XNOR U21581 ( .A(p_input[5417]), .B(n21902), .Z(n21905) );
  XNOR U21582 ( .A(n21902), .B(n21609), .Z(n21904) );
  IV U21583 ( .A(p_input[5385]), .Z(n21609) );
  XOR U21584 ( .A(n21906), .B(n21907), .Z(n21902) );
  AND U21585 ( .A(n21908), .B(n21909), .Z(n21907) );
  XNOR U21586 ( .A(p_input[5416]), .B(n21906), .Z(n21909) );
  XNOR U21587 ( .A(n21906), .B(n21618), .Z(n21908) );
  IV U21588 ( .A(p_input[5384]), .Z(n21618) );
  XOR U21589 ( .A(n21910), .B(n21911), .Z(n21906) );
  AND U21590 ( .A(n21912), .B(n21913), .Z(n21911) );
  XNOR U21591 ( .A(p_input[5415]), .B(n21910), .Z(n21913) );
  XNOR U21592 ( .A(n21910), .B(n21627), .Z(n21912) );
  IV U21593 ( .A(p_input[5383]), .Z(n21627) );
  XOR U21594 ( .A(n21914), .B(n21915), .Z(n21910) );
  AND U21595 ( .A(n21916), .B(n21917), .Z(n21915) );
  XNOR U21596 ( .A(p_input[5414]), .B(n21914), .Z(n21917) );
  XNOR U21597 ( .A(n21914), .B(n21636), .Z(n21916) );
  IV U21598 ( .A(p_input[5382]), .Z(n21636) );
  XOR U21599 ( .A(n21918), .B(n21919), .Z(n21914) );
  AND U21600 ( .A(n21920), .B(n21921), .Z(n21919) );
  XNOR U21601 ( .A(p_input[5413]), .B(n21918), .Z(n21921) );
  XNOR U21602 ( .A(n21918), .B(n21645), .Z(n21920) );
  IV U21603 ( .A(p_input[5381]), .Z(n21645) );
  XOR U21604 ( .A(n21922), .B(n21923), .Z(n21918) );
  AND U21605 ( .A(n21924), .B(n21925), .Z(n21923) );
  XNOR U21606 ( .A(p_input[5412]), .B(n21922), .Z(n21925) );
  XNOR U21607 ( .A(n21922), .B(n21654), .Z(n21924) );
  IV U21608 ( .A(p_input[5380]), .Z(n21654) );
  XOR U21609 ( .A(n21926), .B(n21927), .Z(n21922) );
  AND U21610 ( .A(n21928), .B(n21929), .Z(n21927) );
  XNOR U21611 ( .A(p_input[5411]), .B(n21926), .Z(n21929) );
  XNOR U21612 ( .A(n21926), .B(n21663), .Z(n21928) );
  IV U21613 ( .A(p_input[5379]), .Z(n21663) );
  XOR U21614 ( .A(n21930), .B(n21931), .Z(n21926) );
  AND U21615 ( .A(n21932), .B(n21933), .Z(n21931) );
  XNOR U21616 ( .A(p_input[5410]), .B(n21930), .Z(n21933) );
  XNOR U21617 ( .A(n21930), .B(n21672), .Z(n21932) );
  IV U21618 ( .A(p_input[5378]), .Z(n21672) );
  XNOR U21619 ( .A(n21934), .B(n21935), .Z(n21930) );
  AND U21620 ( .A(n21936), .B(n21937), .Z(n21935) );
  XOR U21621 ( .A(p_input[5409]), .B(n21934), .Z(n21937) );
  XNOR U21622 ( .A(p_input[5377]), .B(n21934), .Z(n21936) );
  AND U21623 ( .A(p_input[5408]), .B(n21938), .Z(n21934) );
  IV U21624 ( .A(p_input[5376]), .Z(n21938) );
  XOR U21625 ( .A(n21939), .B(n21940), .Z(n20117) );
  AND U21626 ( .A(n844), .B(n21941), .Z(n21940) );
  XNOR U21627 ( .A(n21942), .B(n21939), .Z(n21941) );
  XOR U21628 ( .A(n21943), .B(n21944), .Z(n844) );
  AND U21629 ( .A(n21945), .B(n21946), .Z(n21944) );
  XOR U21630 ( .A(n21943), .B(n20132), .Z(n21946) );
  XNOR U21631 ( .A(n21947), .B(n21948), .Z(n20132) );
  AND U21632 ( .A(n21949), .B(n515), .Z(n21948) );
  AND U21633 ( .A(n21947), .B(n21950), .Z(n21949) );
  XNOR U21634 ( .A(n20129), .B(n21943), .Z(n21945) );
  XOR U21635 ( .A(n21951), .B(n21952), .Z(n20129) );
  AND U21636 ( .A(n21953), .B(n512), .Z(n21952) );
  NOR U21637 ( .A(n21951), .B(n21954), .Z(n21953) );
  XOR U21638 ( .A(n21955), .B(n21956), .Z(n21943) );
  AND U21639 ( .A(n21957), .B(n21958), .Z(n21956) );
  XOR U21640 ( .A(n21955), .B(n20144), .Z(n21958) );
  XOR U21641 ( .A(n21959), .B(n21960), .Z(n20144) );
  AND U21642 ( .A(n515), .B(n21961), .Z(n21960) );
  XOR U21643 ( .A(n21962), .B(n21959), .Z(n21961) );
  XNOR U21644 ( .A(n20141), .B(n21955), .Z(n21957) );
  XOR U21645 ( .A(n21963), .B(n21964), .Z(n20141) );
  AND U21646 ( .A(n512), .B(n21965), .Z(n21964) );
  XOR U21647 ( .A(n21966), .B(n21963), .Z(n21965) );
  XOR U21648 ( .A(n21967), .B(n21968), .Z(n21955) );
  AND U21649 ( .A(n21969), .B(n21970), .Z(n21968) );
  XOR U21650 ( .A(n21967), .B(n20156), .Z(n21970) );
  XOR U21651 ( .A(n21971), .B(n21972), .Z(n20156) );
  AND U21652 ( .A(n515), .B(n21973), .Z(n21972) );
  XOR U21653 ( .A(n21974), .B(n21971), .Z(n21973) );
  XNOR U21654 ( .A(n20153), .B(n21967), .Z(n21969) );
  XOR U21655 ( .A(n21975), .B(n21976), .Z(n20153) );
  AND U21656 ( .A(n512), .B(n21977), .Z(n21976) );
  XOR U21657 ( .A(n21978), .B(n21975), .Z(n21977) );
  XOR U21658 ( .A(n21979), .B(n21980), .Z(n21967) );
  AND U21659 ( .A(n21981), .B(n21982), .Z(n21980) );
  XOR U21660 ( .A(n21979), .B(n20168), .Z(n21982) );
  XOR U21661 ( .A(n21983), .B(n21984), .Z(n20168) );
  AND U21662 ( .A(n515), .B(n21985), .Z(n21984) );
  XOR U21663 ( .A(n21986), .B(n21983), .Z(n21985) );
  XNOR U21664 ( .A(n20165), .B(n21979), .Z(n21981) );
  XOR U21665 ( .A(n21987), .B(n21988), .Z(n20165) );
  AND U21666 ( .A(n512), .B(n21989), .Z(n21988) );
  XOR U21667 ( .A(n21990), .B(n21987), .Z(n21989) );
  XOR U21668 ( .A(n21991), .B(n21992), .Z(n21979) );
  AND U21669 ( .A(n21993), .B(n21994), .Z(n21992) );
  XOR U21670 ( .A(n21991), .B(n20180), .Z(n21994) );
  XOR U21671 ( .A(n21995), .B(n21996), .Z(n20180) );
  AND U21672 ( .A(n515), .B(n21997), .Z(n21996) );
  XOR U21673 ( .A(n21998), .B(n21995), .Z(n21997) );
  XNOR U21674 ( .A(n20177), .B(n21991), .Z(n21993) );
  XOR U21675 ( .A(n21999), .B(n22000), .Z(n20177) );
  AND U21676 ( .A(n512), .B(n22001), .Z(n22000) );
  XOR U21677 ( .A(n22002), .B(n21999), .Z(n22001) );
  XOR U21678 ( .A(n22003), .B(n22004), .Z(n21991) );
  AND U21679 ( .A(n22005), .B(n22006), .Z(n22004) );
  XOR U21680 ( .A(n22003), .B(n20192), .Z(n22006) );
  XOR U21681 ( .A(n22007), .B(n22008), .Z(n20192) );
  AND U21682 ( .A(n515), .B(n22009), .Z(n22008) );
  XOR U21683 ( .A(n22010), .B(n22007), .Z(n22009) );
  XNOR U21684 ( .A(n20189), .B(n22003), .Z(n22005) );
  XOR U21685 ( .A(n22011), .B(n22012), .Z(n20189) );
  AND U21686 ( .A(n512), .B(n22013), .Z(n22012) );
  XOR U21687 ( .A(n22014), .B(n22011), .Z(n22013) );
  XOR U21688 ( .A(n22015), .B(n22016), .Z(n22003) );
  AND U21689 ( .A(n22017), .B(n22018), .Z(n22016) );
  XOR U21690 ( .A(n22015), .B(n20204), .Z(n22018) );
  XOR U21691 ( .A(n22019), .B(n22020), .Z(n20204) );
  AND U21692 ( .A(n515), .B(n22021), .Z(n22020) );
  XOR U21693 ( .A(n22022), .B(n22019), .Z(n22021) );
  XNOR U21694 ( .A(n20201), .B(n22015), .Z(n22017) );
  XOR U21695 ( .A(n22023), .B(n22024), .Z(n20201) );
  AND U21696 ( .A(n512), .B(n22025), .Z(n22024) );
  XOR U21697 ( .A(n22026), .B(n22023), .Z(n22025) );
  XOR U21698 ( .A(n22027), .B(n22028), .Z(n22015) );
  AND U21699 ( .A(n22029), .B(n22030), .Z(n22028) );
  XOR U21700 ( .A(n22027), .B(n20216), .Z(n22030) );
  XOR U21701 ( .A(n22031), .B(n22032), .Z(n20216) );
  AND U21702 ( .A(n515), .B(n22033), .Z(n22032) );
  XOR U21703 ( .A(n22034), .B(n22031), .Z(n22033) );
  XNOR U21704 ( .A(n20213), .B(n22027), .Z(n22029) );
  XOR U21705 ( .A(n22035), .B(n22036), .Z(n20213) );
  AND U21706 ( .A(n512), .B(n22037), .Z(n22036) );
  XOR U21707 ( .A(n22038), .B(n22035), .Z(n22037) );
  XOR U21708 ( .A(n22039), .B(n22040), .Z(n22027) );
  AND U21709 ( .A(n22041), .B(n22042), .Z(n22040) );
  XOR U21710 ( .A(n22039), .B(n20228), .Z(n22042) );
  XOR U21711 ( .A(n22043), .B(n22044), .Z(n20228) );
  AND U21712 ( .A(n515), .B(n22045), .Z(n22044) );
  XOR U21713 ( .A(n22046), .B(n22043), .Z(n22045) );
  XNOR U21714 ( .A(n20225), .B(n22039), .Z(n22041) );
  XOR U21715 ( .A(n22047), .B(n22048), .Z(n20225) );
  AND U21716 ( .A(n512), .B(n22049), .Z(n22048) );
  XOR U21717 ( .A(n22050), .B(n22047), .Z(n22049) );
  XOR U21718 ( .A(n22051), .B(n22052), .Z(n22039) );
  AND U21719 ( .A(n22053), .B(n22054), .Z(n22052) );
  XOR U21720 ( .A(n22051), .B(n20240), .Z(n22054) );
  XOR U21721 ( .A(n22055), .B(n22056), .Z(n20240) );
  AND U21722 ( .A(n515), .B(n22057), .Z(n22056) );
  XOR U21723 ( .A(n22058), .B(n22055), .Z(n22057) );
  XNOR U21724 ( .A(n20237), .B(n22051), .Z(n22053) );
  XOR U21725 ( .A(n22059), .B(n22060), .Z(n20237) );
  AND U21726 ( .A(n512), .B(n22061), .Z(n22060) );
  XOR U21727 ( .A(n22062), .B(n22059), .Z(n22061) );
  XOR U21728 ( .A(n22063), .B(n22064), .Z(n22051) );
  AND U21729 ( .A(n22065), .B(n22066), .Z(n22064) );
  XOR U21730 ( .A(n22063), .B(n20252), .Z(n22066) );
  XOR U21731 ( .A(n22067), .B(n22068), .Z(n20252) );
  AND U21732 ( .A(n515), .B(n22069), .Z(n22068) );
  XOR U21733 ( .A(n22070), .B(n22067), .Z(n22069) );
  XNOR U21734 ( .A(n20249), .B(n22063), .Z(n22065) );
  XOR U21735 ( .A(n22071), .B(n22072), .Z(n20249) );
  AND U21736 ( .A(n512), .B(n22073), .Z(n22072) );
  XOR U21737 ( .A(n22074), .B(n22071), .Z(n22073) );
  XOR U21738 ( .A(n22075), .B(n22076), .Z(n22063) );
  AND U21739 ( .A(n22077), .B(n22078), .Z(n22076) );
  XOR U21740 ( .A(n22075), .B(n20264), .Z(n22078) );
  XOR U21741 ( .A(n22079), .B(n22080), .Z(n20264) );
  AND U21742 ( .A(n515), .B(n22081), .Z(n22080) );
  XOR U21743 ( .A(n22082), .B(n22079), .Z(n22081) );
  XNOR U21744 ( .A(n20261), .B(n22075), .Z(n22077) );
  XOR U21745 ( .A(n22083), .B(n22084), .Z(n20261) );
  AND U21746 ( .A(n512), .B(n22085), .Z(n22084) );
  XOR U21747 ( .A(n22086), .B(n22083), .Z(n22085) );
  XOR U21748 ( .A(n22087), .B(n22088), .Z(n22075) );
  AND U21749 ( .A(n22089), .B(n22090), .Z(n22088) );
  XOR U21750 ( .A(n22087), .B(n20276), .Z(n22090) );
  XOR U21751 ( .A(n22091), .B(n22092), .Z(n20276) );
  AND U21752 ( .A(n515), .B(n22093), .Z(n22092) );
  XOR U21753 ( .A(n22094), .B(n22091), .Z(n22093) );
  XNOR U21754 ( .A(n20273), .B(n22087), .Z(n22089) );
  XOR U21755 ( .A(n22095), .B(n22096), .Z(n20273) );
  AND U21756 ( .A(n512), .B(n22097), .Z(n22096) );
  XOR U21757 ( .A(n22098), .B(n22095), .Z(n22097) );
  XOR U21758 ( .A(n22099), .B(n22100), .Z(n22087) );
  AND U21759 ( .A(n22101), .B(n22102), .Z(n22100) );
  XOR U21760 ( .A(n22099), .B(n20288), .Z(n22102) );
  XOR U21761 ( .A(n22103), .B(n22104), .Z(n20288) );
  AND U21762 ( .A(n515), .B(n22105), .Z(n22104) );
  XOR U21763 ( .A(n22106), .B(n22103), .Z(n22105) );
  XNOR U21764 ( .A(n20285), .B(n22099), .Z(n22101) );
  XOR U21765 ( .A(n22107), .B(n22108), .Z(n20285) );
  AND U21766 ( .A(n512), .B(n22109), .Z(n22108) );
  XOR U21767 ( .A(n22110), .B(n22107), .Z(n22109) );
  XOR U21768 ( .A(n22111), .B(n22112), .Z(n22099) );
  AND U21769 ( .A(n22113), .B(n22114), .Z(n22112) );
  XOR U21770 ( .A(n22111), .B(n20300), .Z(n22114) );
  XOR U21771 ( .A(n22115), .B(n22116), .Z(n20300) );
  AND U21772 ( .A(n515), .B(n22117), .Z(n22116) );
  XOR U21773 ( .A(n22118), .B(n22115), .Z(n22117) );
  XNOR U21774 ( .A(n20297), .B(n22111), .Z(n22113) );
  XOR U21775 ( .A(n22119), .B(n22120), .Z(n20297) );
  AND U21776 ( .A(n512), .B(n22121), .Z(n22120) );
  XOR U21777 ( .A(n22122), .B(n22119), .Z(n22121) );
  XOR U21778 ( .A(n22123), .B(n22124), .Z(n22111) );
  AND U21779 ( .A(n22125), .B(n22126), .Z(n22124) );
  XOR U21780 ( .A(n22123), .B(n20312), .Z(n22126) );
  XOR U21781 ( .A(n22127), .B(n22128), .Z(n20312) );
  AND U21782 ( .A(n515), .B(n22129), .Z(n22128) );
  XOR U21783 ( .A(n22130), .B(n22127), .Z(n22129) );
  XNOR U21784 ( .A(n20309), .B(n22123), .Z(n22125) );
  XOR U21785 ( .A(n22131), .B(n22132), .Z(n20309) );
  AND U21786 ( .A(n512), .B(n22133), .Z(n22132) );
  XOR U21787 ( .A(n22134), .B(n22131), .Z(n22133) );
  XOR U21788 ( .A(n22135), .B(n22136), .Z(n22123) );
  AND U21789 ( .A(n22137), .B(n22138), .Z(n22136) );
  XOR U21790 ( .A(n22135), .B(n20324), .Z(n22138) );
  XOR U21791 ( .A(n22139), .B(n22140), .Z(n20324) );
  AND U21792 ( .A(n515), .B(n22141), .Z(n22140) );
  XOR U21793 ( .A(n22142), .B(n22139), .Z(n22141) );
  XNOR U21794 ( .A(n20321), .B(n22135), .Z(n22137) );
  XOR U21795 ( .A(n22143), .B(n22144), .Z(n20321) );
  AND U21796 ( .A(n512), .B(n22145), .Z(n22144) );
  XOR U21797 ( .A(n22146), .B(n22143), .Z(n22145) );
  XOR U21798 ( .A(n22147), .B(n22148), .Z(n22135) );
  AND U21799 ( .A(n22149), .B(n22150), .Z(n22148) );
  XOR U21800 ( .A(n22147), .B(n20336), .Z(n22150) );
  XOR U21801 ( .A(n22151), .B(n22152), .Z(n20336) );
  AND U21802 ( .A(n515), .B(n22153), .Z(n22152) );
  XOR U21803 ( .A(n22154), .B(n22151), .Z(n22153) );
  XNOR U21804 ( .A(n20333), .B(n22147), .Z(n22149) );
  XOR U21805 ( .A(n22155), .B(n22156), .Z(n20333) );
  AND U21806 ( .A(n512), .B(n22157), .Z(n22156) );
  XOR U21807 ( .A(n22158), .B(n22155), .Z(n22157) );
  XOR U21808 ( .A(n22159), .B(n22160), .Z(n22147) );
  AND U21809 ( .A(n22161), .B(n22162), .Z(n22160) );
  XOR U21810 ( .A(n22159), .B(n20348), .Z(n22162) );
  XOR U21811 ( .A(n22163), .B(n22164), .Z(n20348) );
  AND U21812 ( .A(n515), .B(n22165), .Z(n22164) );
  XOR U21813 ( .A(n22166), .B(n22163), .Z(n22165) );
  XNOR U21814 ( .A(n20345), .B(n22159), .Z(n22161) );
  XOR U21815 ( .A(n22167), .B(n22168), .Z(n20345) );
  AND U21816 ( .A(n512), .B(n22169), .Z(n22168) );
  XOR U21817 ( .A(n22170), .B(n22167), .Z(n22169) );
  XOR U21818 ( .A(n22171), .B(n22172), .Z(n22159) );
  AND U21819 ( .A(n22173), .B(n22174), .Z(n22172) );
  XOR U21820 ( .A(n22171), .B(n20360), .Z(n22174) );
  XOR U21821 ( .A(n22175), .B(n22176), .Z(n20360) );
  AND U21822 ( .A(n515), .B(n22177), .Z(n22176) );
  XOR U21823 ( .A(n22178), .B(n22175), .Z(n22177) );
  XNOR U21824 ( .A(n20357), .B(n22171), .Z(n22173) );
  XOR U21825 ( .A(n22179), .B(n22180), .Z(n20357) );
  AND U21826 ( .A(n512), .B(n22181), .Z(n22180) );
  XOR U21827 ( .A(n22182), .B(n22179), .Z(n22181) );
  XOR U21828 ( .A(n22183), .B(n22184), .Z(n22171) );
  AND U21829 ( .A(n22185), .B(n22186), .Z(n22184) );
  XOR U21830 ( .A(n22183), .B(n20372), .Z(n22186) );
  XOR U21831 ( .A(n22187), .B(n22188), .Z(n20372) );
  AND U21832 ( .A(n515), .B(n22189), .Z(n22188) );
  XOR U21833 ( .A(n22190), .B(n22187), .Z(n22189) );
  XNOR U21834 ( .A(n20369), .B(n22183), .Z(n22185) );
  XOR U21835 ( .A(n22191), .B(n22192), .Z(n20369) );
  AND U21836 ( .A(n512), .B(n22193), .Z(n22192) );
  XOR U21837 ( .A(n22194), .B(n22191), .Z(n22193) );
  XOR U21838 ( .A(n22195), .B(n22196), .Z(n22183) );
  AND U21839 ( .A(n22197), .B(n22198), .Z(n22196) );
  XOR U21840 ( .A(n22195), .B(n20384), .Z(n22198) );
  XOR U21841 ( .A(n22199), .B(n22200), .Z(n20384) );
  AND U21842 ( .A(n515), .B(n22201), .Z(n22200) );
  XOR U21843 ( .A(n22202), .B(n22199), .Z(n22201) );
  XNOR U21844 ( .A(n20381), .B(n22195), .Z(n22197) );
  XOR U21845 ( .A(n22203), .B(n22204), .Z(n20381) );
  AND U21846 ( .A(n512), .B(n22205), .Z(n22204) );
  XOR U21847 ( .A(n22206), .B(n22203), .Z(n22205) );
  XOR U21848 ( .A(n22207), .B(n22208), .Z(n22195) );
  AND U21849 ( .A(n22209), .B(n22210), .Z(n22208) );
  XOR U21850 ( .A(n22207), .B(n20396), .Z(n22210) );
  XOR U21851 ( .A(n22211), .B(n22212), .Z(n20396) );
  AND U21852 ( .A(n515), .B(n22213), .Z(n22212) );
  XOR U21853 ( .A(n22214), .B(n22211), .Z(n22213) );
  XNOR U21854 ( .A(n20393), .B(n22207), .Z(n22209) );
  XOR U21855 ( .A(n22215), .B(n22216), .Z(n20393) );
  AND U21856 ( .A(n512), .B(n22217), .Z(n22216) );
  XOR U21857 ( .A(n22218), .B(n22215), .Z(n22217) );
  XOR U21858 ( .A(n22219), .B(n22220), .Z(n22207) );
  AND U21859 ( .A(n22221), .B(n22222), .Z(n22220) );
  XOR U21860 ( .A(n22219), .B(n20408), .Z(n22222) );
  XOR U21861 ( .A(n22223), .B(n22224), .Z(n20408) );
  AND U21862 ( .A(n515), .B(n22225), .Z(n22224) );
  XOR U21863 ( .A(n22226), .B(n22223), .Z(n22225) );
  XNOR U21864 ( .A(n20405), .B(n22219), .Z(n22221) );
  XOR U21865 ( .A(n22227), .B(n22228), .Z(n20405) );
  AND U21866 ( .A(n512), .B(n22229), .Z(n22228) );
  XOR U21867 ( .A(n22230), .B(n22227), .Z(n22229) );
  XOR U21868 ( .A(n22231), .B(n22232), .Z(n22219) );
  AND U21869 ( .A(n22233), .B(n22234), .Z(n22232) );
  XOR U21870 ( .A(n22231), .B(n20420), .Z(n22234) );
  XOR U21871 ( .A(n22235), .B(n22236), .Z(n20420) );
  AND U21872 ( .A(n515), .B(n22237), .Z(n22236) );
  XOR U21873 ( .A(n22238), .B(n22235), .Z(n22237) );
  XNOR U21874 ( .A(n20417), .B(n22231), .Z(n22233) );
  XOR U21875 ( .A(n22239), .B(n22240), .Z(n20417) );
  AND U21876 ( .A(n512), .B(n22241), .Z(n22240) );
  XOR U21877 ( .A(n22242), .B(n22239), .Z(n22241) );
  XOR U21878 ( .A(n22243), .B(n22244), .Z(n22231) );
  AND U21879 ( .A(n22245), .B(n22246), .Z(n22244) );
  XOR U21880 ( .A(n22243), .B(n20432), .Z(n22246) );
  XOR U21881 ( .A(n22247), .B(n22248), .Z(n20432) );
  AND U21882 ( .A(n515), .B(n22249), .Z(n22248) );
  XOR U21883 ( .A(n22250), .B(n22247), .Z(n22249) );
  XNOR U21884 ( .A(n20429), .B(n22243), .Z(n22245) );
  XOR U21885 ( .A(n22251), .B(n22252), .Z(n20429) );
  AND U21886 ( .A(n512), .B(n22253), .Z(n22252) );
  XOR U21887 ( .A(n22254), .B(n22251), .Z(n22253) );
  XOR U21888 ( .A(n22255), .B(n22256), .Z(n22243) );
  AND U21889 ( .A(n22257), .B(n22258), .Z(n22256) );
  XOR U21890 ( .A(n22255), .B(n20444), .Z(n22258) );
  XOR U21891 ( .A(n22259), .B(n22260), .Z(n20444) );
  AND U21892 ( .A(n515), .B(n22261), .Z(n22260) );
  XOR U21893 ( .A(n22262), .B(n22259), .Z(n22261) );
  XNOR U21894 ( .A(n20441), .B(n22255), .Z(n22257) );
  XOR U21895 ( .A(n22263), .B(n22264), .Z(n20441) );
  AND U21896 ( .A(n512), .B(n22265), .Z(n22264) );
  XOR U21897 ( .A(n22266), .B(n22263), .Z(n22265) );
  XOR U21898 ( .A(n22267), .B(n22268), .Z(n22255) );
  AND U21899 ( .A(n22269), .B(n22270), .Z(n22268) );
  XOR U21900 ( .A(n22267), .B(n20456), .Z(n22270) );
  XOR U21901 ( .A(n22271), .B(n22272), .Z(n20456) );
  AND U21902 ( .A(n515), .B(n22273), .Z(n22272) );
  XOR U21903 ( .A(n22274), .B(n22271), .Z(n22273) );
  XNOR U21904 ( .A(n20453), .B(n22267), .Z(n22269) );
  XOR U21905 ( .A(n22275), .B(n22276), .Z(n20453) );
  AND U21906 ( .A(n512), .B(n22277), .Z(n22276) );
  XOR U21907 ( .A(n22278), .B(n22275), .Z(n22277) );
  XOR U21908 ( .A(n22279), .B(n22280), .Z(n22267) );
  AND U21909 ( .A(n22281), .B(n22282), .Z(n22280) );
  XOR U21910 ( .A(n22279), .B(n20468), .Z(n22282) );
  XOR U21911 ( .A(n22283), .B(n22284), .Z(n20468) );
  AND U21912 ( .A(n515), .B(n22285), .Z(n22284) );
  XOR U21913 ( .A(n22286), .B(n22283), .Z(n22285) );
  XNOR U21914 ( .A(n20465), .B(n22279), .Z(n22281) );
  XOR U21915 ( .A(n22287), .B(n22288), .Z(n20465) );
  AND U21916 ( .A(n512), .B(n22289), .Z(n22288) );
  XOR U21917 ( .A(n22290), .B(n22287), .Z(n22289) );
  XOR U21918 ( .A(n22291), .B(n22292), .Z(n22279) );
  AND U21919 ( .A(n22293), .B(n22294), .Z(n22292) );
  XOR U21920 ( .A(n22291), .B(n20480), .Z(n22294) );
  XOR U21921 ( .A(n22295), .B(n22296), .Z(n20480) );
  AND U21922 ( .A(n515), .B(n22297), .Z(n22296) );
  XOR U21923 ( .A(n22298), .B(n22295), .Z(n22297) );
  XNOR U21924 ( .A(n20477), .B(n22291), .Z(n22293) );
  XOR U21925 ( .A(n22299), .B(n22300), .Z(n20477) );
  AND U21926 ( .A(n512), .B(n22301), .Z(n22300) );
  XOR U21927 ( .A(n22302), .B(n22299), .Z(n22301) );
  XOR U21928 ( .A(n22303), .B(n22304), .Z(n22291) );
  AND U21929 ( .A(n22305), .B(n22306), .Z(n22304) );
  XNOR U21930 ( .A(n22307), .B(n20493), .Z(n22306) );
  XOR U21931 ( .A(n22308), .B(n22309), .Z(n20493) );
  AND U21932 ( .A(n515), .B(n22310), .Z(n22309) );
  XOR U21933 ( .A(n22308), .B(n22311), .Z(n22310) );
  XNOR U21934 ( .A(n20490), .B(n22303), .Z(n22305) );
  XOR U21935 ( .A(n22312), .B(n22313), .Z(n20490) );
  AND U21936 ( .A(n512), .B(n22314), .Z(n22313) );
  XOR U21937 ( .A(n22312), .B(n22315), .Z(n22314) );
  IV U21938 ( .A(n22307), .Z(n22303) );
  AND U21939 ( .A(n21939), .B(n21942), .Z(n22307) );
  XNOR U21940 ( .A(n22316), .B(n22317), .Z(n21942) );
  AND U21941 ( .A(n515), .B(n22318), .Z(n22317) );
  XNOR U21942 ( .A(n22319), .B(n22316), .Z(n22318) );
  XOR U21943 ( .A(n22320), .B(n22321), .Z(n515) );
  AND U21944 ( .A(n22322), .B(n22323), .Z(n22321) );
  XOR U21945 ( .A(n21950), .B(n22320), .Z(n22323) );
  IV U21946 ( .A(n22324), .Z(n21950) );
  AND U21947 ( .A(p_input[5375]), .B(p_input[5343]), .Z(n22324) );
  XOR U21948 ( .A(n22320), .B(n21947), .Z(n22322) );
  AND U21949 ( .A(p_input[5279]), .B(p_input[5311]), .Z(n21947) );
  XOR U21950 ( .A(n22325), .B(n22326), .Z(n22320) );
  AND U21951 ( .A(n22327), .B(n22328), .Z(n22326) );
  XOR U21952 ( .A(n22325), .B(n21962), .Z(n22328) );
  XNOR U21953 ( .A(p_input[5342]), .B(n22329), .Z(n21962) );
  AND U21954 ( .A(n351), .B(n22330), .Z(n22329) );
  XOR U21955 ( .A(p_input[5374]), .B(p_input[5342]), .Z(n22330) );
  XNOR U21956 ( .A(n21959), .B(n22325), .Z(n22327) );
  XOR U21957 ( .A(n22331), .B(n22332), .Z(n21959) );
  AND U21958 ( .A(n349), .B(n22333), .Z(n22332) );
  XOR U21959 ( .A(p_input[5310]), .B(p_input[5278]), .Z(n22333) );
  XOR U21960 ( .A(n22334), .B(n22335), .Z(n22325) );
  AND U21961 ( .A(n22336), .B(n22337), .Z(n22335) );
  XOR U21962 ( .A(n22334), .B(n21974), .Z(n22337) );
  XNOR U21963 ( .A(p_input[5341]), .B(n22338), .Z(n21974) );
  AND U21964 ( .A(n351), .B(n22339), .Z(n22338) );
  XOR U21965 ( .A(p_input[5373]), .B(p_input[5341]), .Z(n22339) );
  XNOR U21966 ( .A(n21971), .B(n22334), .Z(n22336) );
  XOR U21967 ( .A(n22340), .B(n22341), .Z(n21971) );
  AND U21968 ( .A(n349), .B(n22342), .Z(n22341) );
  XOR U21969 ( .A(p_input[5309]), .B(p_input[5277]), .Z(n22342) );
  XOR U21970 ( .A(n22343), .B(n22344), .Z(n22334) );
  AND U21971 ( .A(n22345), .B(n22346), .Z(n22344) );
  XOR U21972 ( .A(n22343), .B(n21986), .Z(n22346) );
  XNOR U21973 ( .A(p_input[5340]), .B(n22347), .Z(n21986) );
  AND U21974 ( .A(n351), .B(n22348), .Z(n22347) );
  XOR U21975 ( .A(p_input[5372]), .B(p_input[5340]), .Z(n22348) );
  XNOR U21976 ( .A(n21983), .B(n22343), .Z(n22345) );
  XOR U21977 ( .A(n22349), .B(n22350), .Z(n21983) );
  AND U21978 ( .A(n349), .B(n22351), .Z(n22350) );
  XOR U21979 ( .A(p_input[5308]), .B(p_input[5276]), .Z(n22351) );
  XOR U21980 ( .A(n22352), .B(n22353), .Z(n22343) );
  AND U21981 ( .A(n22354), .B(n22355), .Z(n22353) );
  XOR U21982 ( .A(n22352), .B(n21998), .Z(n22355) );
  XNOR U21983 ( .A(p_input[5339]), .B(n22356), .Z(n21998) );
  AND U21984 ( .A(n351), .B(n22357), .Z(n22356) );
  XOR U21985 ( .A(p_input[5371]), .B(p_input[5339]), .Z(n22357) );
  XNOR U21986 ( .A(n21995), .B(n22352), .Z(n22354) );
  XOR U21987 ( .A(n22358), .B(n22359), .Z(n21995) );
  AND U21988 ( .A(n349), .B(n22360), .Z(n22359) );
  XOR U21989 ( .A(p_input[5307]), .B(p_input[5275]), .Z(n22360) );
  XOR U21990 ( .A(n22361), .B(n22362), .Z(n22352) );
  AND U21991 ( .A(n22363), .B(n22364), .Z(n22362) );
  XOR U21992 ( .A(n22361), .B(n22010), .Z(n22364) );
  XNOR U21993 ( .A(p_input[5338]), .B(n22365), .Z(n22010) );
  AND U21994 ( .A(n351), .B(n22366), .Z(n22365) );
  XOR U21995 ( .A(p_input[5370]), .B(p_input[5338]), .Z(n22366) );
  XNOR U21996 ( .A(n22007), .B(n22361), .Z(n22363) );
  XOR U21997 ( .A(n22367), .B(n22368), .Z(n22007) );
  AND U21998 ( .A(n349), .B(n22369), .Z(n22368) );
  XOR U21999 ( .A(p_input[5306]), .B(p_input[5274]), .Z(n22369) );
  XOR U22000 ( .A(n22370), .B(n22371), .Z(n22361) );
  AND U22001 ( .A(n22372), .B(n22373), .Z(n22371) );
  XOR U22002 ( .A(n22370), .B(n22022), .Z(n22373) );
  XNOR U22003 ( .A(p_input[5337]), .B(n22374), .Z(n22022) );
  AND U22004 ( .A(n351), .B(n22375), .Z(n22374) );
  XOR U22005 ( .A(p_input[5369]), .B(p_input[5337]), .Z(n22375) );
  XNOR U22006 ( .A(n22019), .B(n22370), .Z(n22372) );
  XOR U22007 ( .A(n22376), .B(n22377), .Z(n22019) );
  AND U22008 ( .A(n349), .B(n22378), .Z(n22377) );
  XOR U22009 ( .A(p_input[5305]), .B(p_input[5273]), .Z(n22378) );
  XOR U22010 ( .A(n22379), .B(n22380), .Z(n22370) );
  AND U22011 ( .A(n22381), .B(n22382), .Z(n22380) );
  XOR U22012 ( .A(n22379), .B(n22034), .Z(n22382) );
  XNOR U22013 ( .A(p_input[5336]), .B(n22383), .Z(n22034) );
  AND U22014 ( .A(n351), .B(n22384), .Z(n22383) );
  XOR U22015 ( .A(p_input[5368]), .B(p_input[5336]), .Z(n22384) );
  XNOR U22016 ( .A(n22031), .B(n22379), .Z(n22381) );
  XOR U22017 ( .A(n22385), .B(n22386), .Z(n22031) );
  AND U22018 ( .A(n349), .B(n22387), .Z(n22386) );
  XOR U22019 ( .A(p_input[5304]), .B(p_input[5272]), .Z(n22387) );
  XOR U22020 ( .A(n22388), .B(n22389), .Z(n22379) );
  AND U22021 ( .A(n22390), .B(n22391), .Z(n22389) );
  XOR U22022 ( .A(n22388), .B(n22046), .Z(n22391) );
  XNOR U22023 ( .A(p_input[5335]), .B(n22392), .Z(n22046) );
  AND U22024 ( .A(n351), .B(n22393), .Z(n22392) );
  XOR U22025 ( .A(p_input[5367]), .B(p_input[5335]), .Z(n22393) );
  XNOR U22026 ( .A(n22043), .B(n22388), .Z(n22390) );
  XOR U22027 ( .A(n22394), .B(n22395), .Z(n22043) );
  AND U22028 ( .A(n349), .B(n22396), .Z(n22395) );
  XOR U22029 ( .A(p_input[5303]), .B(p_input[5271]), .Z(n22396) );
  XOR U22030 ( .A(n22397), .B(n22398), .Z(n22388) );
  AND U22031 ( .A(n22399), .B(n22400), .Z(n22398) );
  XOR U22032 ( .A(n22397), .B(n22058), .Z(n22400) );
  XNOR U22033 ( .A(p_input[5334]), .B(n22401), .Z(n22058) );
  AND U22034 ( .A(n351), .B(n22402), .Z(n22401) );
  XOR U22035 ( .A(p_input[5366]), .B(p_input[5334]), .Z(n22402) );
  XNOR U22036 ( .A(n22055), .B(n22397), .Z(n22399) );
  XOR U22037 ( .A(n22403), .B(n22404), .Z(n22055) );
  AND U22038 ( .A(n349), .B(n22405), .Z(n22404) );
  XOR U22039 ( .A(p_input[5302]), .B(p_input[5270]), .Z(n22405) );
  XOR U22040 ( .A(n22406), .B(n22407), .Z(n22397) );
  AND U22041 ( .A(n22408), .B(n22409), .Z(n22407) );
  XOR U22042 ( .A(n22406), .B(n22070), .Z(n22409) );
  XNOR U22043 ( .A(p_input[5333]), .B(n22410), .Z(n22070) );
  AND U22044 ( .A(n351), .B(n22411), .Z(n22410) );
  XOR U22045 ( .A(p_input[5365]), .B(p_input[5333]), .Z(n22411) );
  XNOR U22046 ( .A(n22067), .B(n22406), .Z(n22408) );
  XOR U22047 ( .A(n22412), .B(n22413), .Z(n22067) );
  AND U22048 ( .A(n349), .B(n22414), .Z(n22413) );
  XOR U22049 ( .A(p_input[5301]), .B(p_input[5269]), .Z(n22414) );
  XOR U22050 ( .A(n22415), .B(n22416), .Z(n22406) );
  AND U22051 ( .A(n22417), .B(n22418), .Z(n22416) );
  XOR U22052 ( .A(n22415), .B(n22082), .Z(n22418) );
  XNOR U22053 ( .A(p_input[5332]), .B(n22419), .Z(n22082) );
  AND U22054 ( .A(n351), .B(n22420), .Z(n22419) );
  XOR U22055 ( .A(p_input[5364]), .B(p_input[5332]), .Z(n22420) );
  XNOR U22056 ( .A(n22079), .B(n22415), .Z(n22417) );
  XOR U22057 ( .A(n22421), .B(n22422), .Z(n22079) );
  AND U22058 ( .A(n349), .B(n22423), .Z(n22422) );
  XOR U22059 ( .A(p_input[5300]), .B(p_input[5268]), .Z(n22423) );
  XOR U22060 ( .A(n22424), .B(n22425), .Z(n22415) );
  AND U22061 ( .A(n22426), .B(n22427), .Z(n22425) );
  XOR U22062 ( .A(n22424), .B(n22094), .Z(n22427) );
  XNOR U22063 ( .A(p_input[5331]), .B(n22428), .Z(n22094) );
  AND U22064 ( .A(n351), .B(n22429), .Z(n22428) );
  XOR U22065 ( .A(p_input[5363]), .B(p_input[5331]), .Z(n22429) );
  XNOR U22066 ( .A(n22091), .B(n22424), .Z(n22426) );
  XOR U22067 ( .A(n22430), .B(n22431), .Z(n22091) );
  AND U22068 ( .A(n349), .B(n22432), .Z(n22431) );
  XOR U22069 ( .A(p_input[5299]), .B(p_input[5267]), .Z(n22432) );
  XOR U22070 ( .A(n22433), .B(n22434), .Z(n22424) );
  AND U22071 ( .A(n22435), .B(n22436), .Z(n22434) );
  XOR U22072 ( .A(n22433), .B(n22106), .Z(n22436) );
  XNOR U22073 ( .A(p_input[5330]), .B(n22437), .Z(n22106) );
  AND U22074 ( .A(n351), .B(n22438), .Z(n22437) );
  XOR U22075 ( .A(p_input[5362]), .B(p_input[5330]), .Z(n22438) );
  XNOR U22076 ( .A(n22103), .B(n22433), .Z(n22435) );
  XOR U22077 ( .A(n22439), .B(n22440), .Z(n22103) );
  AND U22078 ( .A(n349), .B(n22441), .Z(n22440) );
  XOR U22079 ( .A(p_input[5298]), .B(p_input[5266]), .Z(n22441) );
  XOR U22080 ( .A(n22442), .B(n22443), .Z(n22433) );
  AND U22081 ( .A(n22444), .B(n22445), .Z(n22443) );
  XOR U22082 ( .A(n22442), .B(n22118), .Z(n22445) );
  XNOR U22083 ( .A(p_input[5329]), .B(n22446), .Z(n22118) );
  AND U22084 ( .A(n351), .B(n22447), .Z(n22446) );
  XOR U22085 ( .A(p_input[5361]), .B(p_input[5329]), .Z(n22447) );
  XNOR U22086 ( .A(n22115), .B(n22442), .Z(n22444) );
  XOR U22087 ( .A(n22448), .B(n22449), .Z(n22115) );
  AND U22088 ( .A(n349), .B(n22450), .Z(n22449) );
  XOR U22089 ( .A(p_input[5297]), .B(p_input[5265]), .Z(n22450) );
  XOR U22090 ( .A(n22451), .B(n22452), .Z(n22442) );
  AND U22091 ( .A(n22453), .B(n22454), .Z(n22452) );
  XOR U22092 ( .A(n22451), .B(n22130), .Z(n22454) );
  XNOR U22093 ( .A(p_input[5328]), .B(n22455), .Z(n22130) );
  AND U22094 ( .A(n351), .B(n22456), .Z(n22455) );
  XOR U22095 ( .A(p_input[5360]), .B(p_input[5328]), .Z(n22456) );
  XNOR U22096 ( .A(n22127), .B(n22451), .Z(n22453) );
  XOR U22097 ( .A(n22457), .B(n22458), .Z(n22127) );
  AND U22098 ( .A(n349), .B(n22459), .Z(n22458) );
  XOR U22099 ( .A(p_input[5296]), .B(p_input[5264]), .Z(n22459) );
  XOR U22100 ( .A(n22460), .B(n22461), .Z(n22451) );
  AND U22101 ( .A(n22462), .B(n22463), .Z(n22461) );
  XOR U22102 ( .A(n22460), .B(n22142), .Z(n22463) );
  XNOR U22103 ( .A(p_input[5327]), .B(n22464), .Z(n22142) );
  AND U22104 ( .A(n351), .B(n22465), .Z(n22464) );
  XOR U22105 ( .A(p_input[5359]), .B(p_input[5327]), .Z(n22465) );
  XNOR U22106 ( .A(n22139), .B(n22460), .Z(n22462) );
  XOR U22107 ( .A(n22466), .B(n22467), .Z(n22139) );
  AND U22108 ( .A(n349), .B(n22468), .Z(n22467) );
  XOR U22109 ( .A(p_input[5295]), .B(p_input[5263]), .Z(n22468) );
  XOR U22110 ( .A(n22469), .B(n22470), .Z(n22460) );
  AND U22111 ( .A(n22471), .B(n22472), .Z(n22470) );
  XOR U22112 ( .A(n22469), .B(n22154), .Z(n22472) );
  XNOR U22113 ( .A(p_input[5326]), .B(n22473), .Z(n22154) );
  AND U22114 ( .A(n351), .B(n22474), .Z(n22473) );
  XOR U22115 ( .A(p_input[5358]), .B(p_input[5326]), .Z(n22474) );
  XNOR U22116 ( .A(n22151), .B(n22469), .Z(n22471) );
  XOR U22117 ( .A(n22475), .B(n22476), .Z(n22151) );
  AND U22118 ( .A(n349), .B(n22477), .Z(n22476) );
  XOR U22119 ( .A(p_input[5294]), .B(p_input[5262]), .Z(n22477) );
  XOR U22120 ( .A(n22478), .B(n22479), .Z(n22469) );
  AND U22121 ( .A(n22480), .B(n22481), .Z(n22479) );
  XOR U22122 ( .A(n22478), .B(n22166), .Z(n22481) );
  XNOR U22123 ( .A(p_input[5325]), .B(n22482), .Z(n22166) );
  AND U22124 ( .A(n351), .B(n22483), .Z(n22482) );
  XOR U22125 ( .A(p_input[5357]), .B(p_input[5325]), .Z(n22483) );
  XNOR U22126 ( .A(n22163), .B(n22478), .Z(n22480) );
  XOR U22127 ( .A(n22484), .B(n22485), .Z(n22163) );
  AND U22128 ( .A(n349), .B(n22486), .Z(n22485) );
  XOR U22129 ( .A(p_input[5293]), .B(p_input[5261]), .Z(n22486) );
  XOR U22130 ( .A(n22487), .B(n22488), .Z(n22478) );
  AND U22131 ( .A(n22489), .B(n22490), .Z(n22488) );
  XOR U22132 ( .A(n22487), .B(n22178), .Z(n22490) );
  XNOR U22133 ( .A(p_input[5324]), .B(n22491), .Z(n22178) );
  AND U22134 ( .A(n351), .B(n22492), .Z(n22491) );
  XOR U22135 ( .A(p_input[5356]), .B(p_input[5324]), .Z(n22492) );
  XNOR U22136 ( .A(n22175), .B(n22487), .Z(n22489) );
  XOR U22137 ( .A(n22493), .B(n22494), .Z(n22175) );
  AND U22138 ( .A(n349), .B(n22495), .Z(n22494) );
  XOR U22139 ( .A(p_input[5292]), .B(p_input[5260]), .Z(n22495) );
  XOR U22140 ( .A(n22496), .B(n22497), .Z(n22487) );
  AND U22141 ( .A(n22498), .B(n22499), .Z(n22497) );
  XOR U22142 ( .A(n22496), .B(n22190), .Z(n22499) );
  XNOR U22143 ( .A(p_input[5323]), .B(n22500), .Z(n22190) );
  AND U22144 ( .A(n351), .B(n22501), .Z(n22500) );
  XOR U22145 ( .A(p_input[5355]), .B(p_input[5323]), .Z(n22501) );
  XNOR U22146 ( .A(n22187), .B(n22496), .Z(n22498) );
  XOR U22147 ( .A(n22502), .B(n22503), .Z(n22187) );
  AND U22148 ( .A(n349), .B(n22504), .Z(n22503) );
  XOR U22149 ( .A(p_input[5291]), .B(p_input[5259]), .Z(n22504) );
  XOR U22150 ( .A(n22505), .B(n22506), .Z(n22496) );
  AND U22151 ( .A(n22507), .B(n22508), .Z(n22506) );
  XOR U22152 ( .A(n22505), .B(n22202), .Z(n22508) );
  XNOR U22153 ( .A(p_input[5322]), .B(n22509), .Z(n22202) );
  AND U22154 ( .A(n351), .B(n22510), .Z(n22509) );
  XOR U22155 ( .A(p_input[5354]), .B(p_input[5322]), .Z(n22510) );
  XNOR U22156 ( .A(n22199), .B(n22505), .Z(n22507) );
  XOR U22157 ( .A(n22511), .B(n22512), .Z(n22199) );
  AND U22158 ( .A(n349), .B(n22513), .Z(n22512) );
  XOR U22159 ( .A(p_input[5290]), .B(p_input[5258]), .Z(n22513) );
  XOR U22160 ( .A(n22514), .B(n22515), .Z(n22505) );
  AND U22161 ( .A(n22516), .B(n22517), .Z(n22515) );
  XOR U22162 ( .A(n22514), .B(n22214), .Z(n22517) );
  XNOR U22163 ( .A(p_input[5321]), .B(n22518), .Z(n22214) );
  AND U22164 ( .A(n351), .B(n22519), .Z(n22518) );
  XOR U22165 ( .A(p_input[5353]), .B(p_input[5321]), .Z(n22519) );
  XNOR U22166 ( .A(n22211), .B(n22514), .Z(n22516) );
  XOR U22167 ( .A(n22520), .B(n22521), .Z(n22211) );
  AND U22168 ( .A(n349), .B(n22522), .Z(n22521) );
  XOR U22169 ( .A(p_input[5289]), .B(p_input[5257]), .Z(n22522) );
  XOR U22170 ( .A(n22523), .B(n22524), .Z(n22514) );
  AND U22171 ( .A(n22525), .B(n22526), .Z(n22524) );
  XOR U22172 ( .A(n22523), .B(n22226), .Z(n22526) );
  XNOR U22173 ( .A(p_input[5320]), .B(n22527), .Z(n22226) );
  AND U22174 ( .A(n351), .B(n22528), .Z(n22527) );
  XOR U22175 ( .A(p_input[5352]), .B(p_input[5320]), .Z(n22528) );
  XNOR U22176 ( .A(n22223), .B(n22523), .Z(n22525) );
  XOR U22177 ( .A(n22529), .B(n22530), .Z(n22223) );
  AND U22178 ( .A(n349), .B(n22531), .Z(n22530) );
  XOR U22179 ( .A(p_input[5288]), .B(p_input[5256]), .Z(n22531) );
  XOR U22180 ( .A(n22532), .B(n22533), .Z(n22523) );
  AND U22181 ( .A(n22534), .B(n22535), .Z(n22533) );
  XOR U22182 ( .A(n22532), .B(n22238), .Z(n22535) );
  XNOR U22183 ( .A(p_input[5319]), .B(n22536), .Z(n22238) );
  AND U22184 ( .A(n351), .B(n22537), .Z(n22536) );
  XOR U22185 ( .A(p_input[5351]), .B(p_input[5319]), .Z(n22537) );
  XNOR U22186 ( .A(n22235), .B(n22532), .Z(n22534) );
  XOR U22187 ( .A(n22538), .B(n22539), .Z(n22235) );
  AND U22188 ( .A(n349), .B(n22540), .Z(n22539) );
  XOR U22189 ( .A(p_input[5287]), .B(p_input[5255]), .Z(n22540) );
  XOR U22190 ( .A(n22541), .B(n22542), .Z(n22532) );
  AND U22191 ( .A(n22543), .B(n22544), .Z(n22542) );
  XOR U22192 ( .A(n22541), .B(n22250), .Z(n22544) );
  XNOR U22193 ( .A(p_input[5318]), .B(n22545), .Z(n22250) );
  AND U22194 ( .A(n351), .B(n22546), .Z(n22545) );
  XOR U22195 ( .A(p_input[5350]), .B(p_input[5318]), .Z(n22546) );
  XNOR U22196 ( .A(n22247), .B(n22541), .Z(n22543) );
  XOR U22197 ( .A(n22547), .B(n22548), .Z(n22247) );
  AND U22198 ( .A(n349), .B(n22549), .Z(n22548) );
  XOR U22199 ( .A(p_input[5286]), .B(p_input[5254]), .Z(n22549) );
  XOR U22200 ( .A(n22550), .B(n22551), .Z(n22541) );
  AND U22201 ( .A(n22552), .B(n22553), .Z(n22551) );
  XOR U22202 ( .A(n22550), .B(n22262), .Z(n22553) );
  XNOR U22203 ( .A(p_input[5317]), .B(n22554), .Z(n22262) );
  AND U22204 ( .A(n351), .B(n22555), .Z(n22554) );
  XOR U22205 ( .A(p_input[5349]), .B(p_input[5317]), .Z(n22555) );
  XNOR U22206 ( .A(n22259), .B(n22550), .Z(n22552) );
  XOR U22207 ( .A(n22556), .B(n22557), .Z(n22259) );
  AND U22208 ( .A(n349), .B(n22558), .Z(n22557) );
  XOR U22209 ( .A(p_input[5285]), .B(p_input[5253]), .Z(n22558) );
  XOR U22210 ( .A(n22559), .B(n22560), .Z(n22550) );
  AND U22211 ( .A(n22561), .B(n22562), .Z(n22560) );
  XOR U22212 ( .A(n22559), .B(n22274), .Z(n22562) );
  XNOR U22213 ( .A(p_input[5316]), .B(n22563), .Z(n22274) );
  AND U22214 ( .A(n351), .B(n22564), .Z(n22563) );
  XOR U22215 ( .A(p_input[5348]), .B(p_input[5316]), .Z(n22564) );
  XNOR U22216 ( .A(n22271), .B(n22559), .Z(n22561) );
  XOR U22217 ( .A(n22565), .B(n22566), .Z(n22271) );
  AND U22218 ( .A(n349), .B(n22567), .Z(n22566) );
  XOR U22219 ( .A(p_input[5284]), .B(p_input[5252]), .Z(n22567) );
  XOR U22220 ( .A(n22568), .B(n22569), .Z(n22559) );
  AND U22221 ( .A(n22570), .B(n22571), .Z(n22569) );
  XOR U22222 ( .A(n22568), .B(n22286), .Z(n22571) );
  XNOR U22223 ( .A(p_input[5315]), .B(n22572), .Z(n22286) );
  AND U22224 ( .A(n351), .B(n22573), .Z(n22572) );
  XOR U22225 ( .A(p_input[5347]), .B(p_input[5315]), .Z(n22573) );
  XNOR U22226 ( .A(n22283), .B(n22568), .Z(n22570) );
  XOR U22227 ( .A(n22574), .B(n22575), .Z(n22283) );
  AND U22228 ( .A(n349), .B(n22576), .Z(n22575) );
  XOR U22229 ( .A(p_input[5283]), .B(p_input[5251]), .Z(n22576) );
  XOR U22230 ( .A(n22577), .B(n22578), .Z(n22568) );
  AND U22231 ( .A(n22579), .B(n22580), .Z(n22578) );
  XOR U22232 ( .A(n22577), .B(n22298), .Z(n22580) );
  XNOR U22233 ( .A(p_input[5314]), .B(n22581), .Z(n22298) );
  AND U22234 ( .A(n351), .B(n22582), .Z(n22581) );
  XOR U22235 ( .A(p_input[5346]), .B(p_input[5314]), .Z(n22582) );
  XNOR U22236 ( .A(n22295), .B(n22577), .Z(n22579) );
  XOR U22237 ( .A(n22583), .B(n22584), .Z(n22295) );
  AND U22238 ( .A(n349), .B(n22585), .Z(n22584) );
  XOR U22239 ( .A(p_input[5282]), .B(p_input[5250]), .Z(n22585) );
  XOR U22240 ( .A(n22586), .B(n22587), .Z(n22577) );
  AND U22241 ( .A(n22588), .B(n22589), .Z(n22587) );
  XNOR U22242 ( .A(n22590), .B(n22311), .Z(n22589) );
  XNOR U22243 ( .A(p_input[5313]), .B(n22591), .Z(n22311) );
  AND U22244 ( .A(n351), .B(n22592), .Z(n22591) );
  XNOR U22245 ( .A(p_input[5345]), .B(n22593), .Z(n22592) );
  IV U22246 ( .A(p_input[5313]), .Z(n22593) );
  XNOR U22247 ( .A(n22308), .B(n22586), .Z(n22588) );
  XNOR U22248 ( .A(p_input[5249]), .B(n22594), .Z(n22308) );
  AND U22249 ( .A(n349), .B(n22595), .Z(n22594) );
  XOR U22250 ( .A(p_input[5281]), .B(p_input[5249]), .Z(n22595) );
  IV U22251 ( .A(n22590), .Z(n22586) );
  AND U22252 ( .A(n22316), .B(n22319), .Z(n22590) );
  XOR U22253 ( .A(p_input[5312]), .B(n22596), .Z(n22319) );
  AND U22254 ( .A(n351), .B(n22597), .Z(n22596) );
  XOR U22255 ( .A(p_input[5344]), .B(p_input[5312]), .Z(n22597) );
  XOR U22256 ( .A(n22598), .B(n22599), .Z(n351) );
  AND U22257 ( .A(n22600), .B(n22601), .Z(n22599) );
  XNOR U22258 ( .A(p_input[5375]), .B(n22598), .Z(n22601) );
  XOR U22259 ( .A(n22598), .B(p_input[5343]), .Z(n22600) );
  XOR U22260 ( .A(n22602), .B(n22603), .Z(n22598) );
  AND U22261 ( .A(n22604), .B(n22605), .Z(n22603) );
  XNOR U22262 ( .A(p_input[5374]), .B(n22602), .Z(n22605) );
  XOR U22263 ( .A(n22602), .B(p_input[5342]), .Z(n22604) );
  XOR U22264 ( .A(n22606), .B(n22607), .Z(n22602) );
  AND U22265 ( .A(n22608), .B(n22609), .Z(n22607) );
  XNOR U22266 ( .A(p_input[5373]), .B(n22606), .Z(n22609) );
  XOR U22267 ( .A(n22606), .B(p_input[5341]), .Z(n22608) );
  XOR U22268 ( .A(n22610), .B(n22611), .Z(n22606) );
  AND U22269 ( .A(n22612), .B(n22613), .Z(n22611) );
  XNOR U22270 ( .A(p_input[5372]), .B(n22610), .Z(n22613) );
  XOR U22271 ( .A(n22610), .B(p_input[5340]), .Z(n22612) );
  XOR U22272 ( .A(n22614), .B(n22615), .Z(n22610) );
  AND U22273 ( .A(n22616), .B(n22617), .Z(n22615) );
  XNOR U22274 ( .A(p_input[5371]), .B(n22614), .Z(n22617) );
  XOR U22275 ( .A(n22614), .B(p_input[5339]), .Z(n22616) );
  XOR U22276 ( .A(n22618), .B(n22619), .Z(n22614) );
  AND U22277 ( .A(n22620), .B(n22621), .Z(n22619) );
  XNOR U22278 ( .A(p_input[5370]), .B(n22618), .Z(n22621) );
  XOR U22279 ( .A(n22618), .B(p_input[5338]), .Z(n22620) );
  XOR U22280 ( .A(n22622), .B(n22623), .Z(n22618) );
  AND U22281 ( .A(n22624), .B(n22625), .Z(n22623) );
  XNOR U22282 ( .A(p_input[5369]), .B(n22622), .Z(n22625) );
  XOR U22283 ( .A(n22622), .B(p_input[5337]), .Z(n22624) );
  XOR U22284 ( .A(n22626), .B(n22627), .Z(n22622) );
  AND U22285 ( .A(n22628), .B(n22629), .Z(n22627) );
  XNOR U22286 ( .A(p_input[5368]), .B(n22626), .Z(n22629) );
  XOR U22287 ( .A(n22626), .B(p_input[5336]), .Z(n22628) );
  XOR U22288 ( .A(n22630), .B(n22631), .Z(n22626) );
  AND U22289 ( .A(n22632), .B(n22633), .Z(n22631) );
  XNOR U22290 ( .A(p_input[5367]), .B(n22630), .Z(n22633) );
  XOR U22291 ( .A(n22630), .B(p_input[5335]), .Z(n22632) );
  XOR U22292 ( .A(n22634), .B(n22635), .Z(n22630) );
  AND U22293 ( .A(n22636), .B(n22637), .Z(n22635) );
  XNOR U22294 ( .A(p_input[5366]), .B(n22634), .Z(n22637) );
  XOR U22295 ( .A(n22634), .B(p_input[5334]), .Z(n22636) );
  XOR U22296 ( .A(n22638), .B(n22639), .Z(n22634) );
  AND U22297 ( .A(n22640), .B(n22641), .Z(n22639) );
  XNOR U22298 ( .A(p_input[5365]), .B(n22638), .Z(n22641) );
  XOR U22299 ( .A(n22638), .B(p_input[5333]), .Z(n22640) );
  XOR U22300 ( .A(n22642), .B(n22643), .Z(n22638) );
  AND U22301 ( .A(n22644), .B(n22645), .Z(n22643) );
  XNOR U22302 ( .A(p_input[5364]), .B(n22642), .Z(n22645) );
  XOR U22303 ( .A(n22642), .B(p_input[5332]), .Z(n22644) );
  XOR U22304 ( .A(n22646), .B(n22647), .Z(n22642) );
  AND U22305 ( .A(n22648), .B(n22649), .Z(n22647) );
  XNOR U22306 ( .A(p_input[5363]), .B(n22646), .Z(n22649) );
  XOR U22307 ( .A(n22646), .B(p_input[5331]), .Z(n22648) );
  XOR U22308 ( .A(n22650), .B(n22651), .Z(n22646) );
  AND U22309 ( .A(n22652), .B(n22653), .Z(n22651) );
  XNOR U22310 ( .A(p_input[5362]), .B(n22650), .Z(n22653) );
  XOR U22311 ( .A(n22650), .B(p_input[5330]), .Z(n22652) );
  XOR U22312 ( .A(n22654), .B(n22655), .Z(n22650) );
  AND U22313 ( .A(n22656), .B(n22657), .Z(n22655) );
  XNOR U22314 ( .A(p_input[5361]), .B(n22654), .Z(n22657) );
  XOR U22315 ( .A(n22654), .B(p_input[5329]), .Z(n22656) );
  XOR U22316 ( .A(n22658), .B(n22659), .Z(n22654) );
  AND U22317 ( .A(n22660), .B(n22661), .Z(n22659) );
  XNOR U22318 ( .A(p_input[5360]), .B(n22658), .Z(n22661) );
  XOR U22319 ( .A(n22658), .B(p_input[5328]), .Z(n22660) );
  XOR U22320 ( .A(n22662), .B(n22663), .Z(n22658) );
  AND U22321 ( .A(n22664), .B(n22665), .Z(n22663) );
  XNOR U22322 ( .A(p_input[5359]), .B(n22662), .Z(n22665) );
  XOR U22323 ( .A(n22662), .B(p_input[5327]), .Z(n22664) );
  XOR U22324 ( .A(n22666), .B(n22667), .Z(n22662) );
  AND U22325 ( .A(n22668), .B(n22669), .Z(n22667) );
  XNOR U22326 ( .A(p_input[5358]), .B(n22666), .Z(n22669) );
  XOR U22327 ( .A(n22666), .B(p_input[5326]), .Z(n22668) );
  XOR U22328 ( .A(n22670), .B(n22671), .Z(n22666) );
  AND U22329 ( .A(n22672), .B(n22673), .Z(n22671) );
  XNOR U22330 ( .A(p_input[5357]), .B(n22670), .Z(n22673) );
  XOR U22331 ( .A(n22670), .B(p_input[5325]), .Z(n22672) );
  XOR U22332 ( .A(n22674), .B(n22675), .Z(n22670) );
  AND U22333 ( .A(n22676), .B(n22677), .Z(n22675) );
  XNOR U22334 ( .A(p_input[5356]), .B(n22674), .Z(n22677) );
  XOR U22335 ( .A(n22674), .B(p_input[5324]), .Z(n22676) );
  XOR U22336 ( .A(n22678), .B(n22679), .Z(n22674) );
  AND U22337 ( .A(n22680), .B(n22681), .Z(n22679) );
  XNOR U22338 ( .A(p_input[5355]), .B(n22678), .Z(n22681) );
  XOR U22339 ( .A(n22678), .B(p_input[5323]), .Z(n22680) );
  XOR U22340 ( .A(n22682), .B(n22683), .Z(n22678) );
  AND U22341 ( .A(n22684), .B(n22685), .Z(n22683) );
  XNOR U22342 ( .A(p_input[5354]), .B(n22682), .Z(n22685) );
  XOR U22343 ( .A(n22682), .B(p_input[5322]), .Z(n22684) );
  XOR U22344 ( .A(n22686), .B(n22687), .Z(n22682) );
  AND U22345 ( .A(n22688), .B(n22689), .Z(n22687) );
  XNOR U22346 ( .A(p_input[5353]), .B(n22686), .Z(n22689) );
  XOR U22347 ( .A(n22686), .B(p_input[5321]), .Z(n22688) );
  XOR U22348 ( .A(n22690), .B(n22691), .Z(n22686) );
  AND U22349 ( .A(n22692), .B(n22693), .Z(n22691) );
  XNOR U22350 ( .A(p_input[5352]), .B(n22690), .Z(n22693) );
  XOR U22351 ( .A(n22690), .B(p_input[5320]), .Z(n22692) );
  XOR U22352 ( .A(n22694), .B(n22695), .Z(n22690) );
  AND U22353 ( .A(n22696), .B(n22697), .Z(n22695) );
  XNOR U22354 ( .A(p_input[5351]), .B(n22694), .Z(n22697) );
  XOR U22355 ( .A(n22694), .B(p_input[5319]), .Z(n22696) );
  XOR U22356 ( .A(n22698), .B(n22699), .Z(n22694) );
  AND U22357 ( .A(n22700), .B(n22701), .Z(n22699) );
  XNOR U22358 ( .A(p_input[5350]), .B(n22698), .Z(n22701) );
  XOR U22359 ( .A(n22698), .B(p_input[5318]), .Z(n22700) );
  XOR U22360 ( .A(n22702), .B(n22703), .Z(n22698) );
  AND U22361 ( .A(n22704), .B(n22705), .Z(n22703) );
  XNOR U22362 ( .A(p_input[5349]), .B(n22702), .Z(n22705) );
  XOR U22363 ( .A(n22702), .B(p_input[5317]), .Z(n22704) );
  XOR U22364 ( .A(n22706), .B(n22707), .Z(n22702) );
  AND U22365 ( .A(n22708), .B(n22709), .Z(n22707) );
  XNOR U22366 ( .A(p_input[5348]), .B(n22706), .Z(n22709) );
  XOR U22367 ( .A(n22706), .B(p_input[5316]), .Z(n22708) );
  XOR U22368 ( .A(n22710), .B(n22711), .Z(n22706) );
  AND U22369 ( .A(n22712), .B(n22713), .Z(n22711) );
  XNOR U22370 ( .A(p_input[5347]), .B(n22710), .Z(n22713) );
  XOR U22371 ( .A(n22710), .B(p_input[5315]), .Z(n22712) );
  XOR U22372 ( .A(n22714), .B(n22715), .Z(n22710) );
  AND U22373 ( .A(n22716), .B(n22717), .Z(n22715) );
  XNOR U22374 ( .A(p_input[5346]), .B(n22714), .Z(n22717) );
  XOR U22375 ( .A(n22714), .B(p_input[5314]), .Z(n22716) );
  XNOR U22376 ( .A(n22718), .B(n22719), .Z(n22714) );
  AND U22377 ( .A(n22720), .B(n22721), .Z(n22719) );
  XOR U22378 ( .A(p_input[5345]), .B(n22718), .Z(n22721) );
  XNOR U22379 ( .A(p_input[5313]), .B(n22718), .Z(n22720) );
  AND U22380 ( .A(p_input[5344]), .B(n22722), .Z(n22718) );
  IV U22381 ( .A(p_input[5312]), .Z(n22722) );
  XNOR U22382 ( .A(p_input[5248]), .B(n22723), .Z(n22316) );
  AND U22383 ( .A(n349), .B(n22724), .Z(n22723) );
  XOR U22384 ( .A(p_input[5280]), .B(p_input[5248]), .Z(n22724) );
  XOR U22385 ( .A(n22725), .B(n22726), .Z(n349) );
  AND U22386 ( .A(n22727), .B(n22728), .Z(n22726) );
  XNOR U22387 ( .A(p_input[5311]), .B(n22725), .Z(n22728) );
  XOR U22388 ( .A(n22725), .B(p_input[5279]), .Z(n22727) );
  XOR U22389 ( .A(n22729), .B(n22730), .Z(n22725) );
  AND U22390 ( .A(n22731), .B(n22732), .Z(n22730) );
  XNOR U22391 ( .A(p_input[5310]), .B(n22729), .Z(n22732) );
  XNOR U22392 ( .A(n22729), .B(n22331), .Z(n22731) );
  IV U22393 ( .A(p_input[5278]), .Z(n22331) );
  XOR U22394 ( .A(n22733), .B(n22734), .Z(n22729) );
  AND U22395 ( .A(n22735), .B(n22736), .Z(n22734) );
  XNOR U22396 ( .A(p_input[5309]), .B(n22733), .Z(n22736) );
  XNOR U22397 ( .A(n22733), .B(n22340), .Z(n22735) );
  IV U22398 ( .A(p_input[5277]), .Z(n22340) );
  XOR U22399 ( .A(n22737), .B(n22738), .Z(n22733) );
  AND U22400 ( .A(n22739), .B(n22740), .Z(n22738) );
  XNOR U22401 ( .A(p_input[5308]), .B(n22737), .Z(n22740) );
  XNOR U22402 ( .A(n22737), .B(n22349), .Z(n22739) );
  IV U22403 ( .A(p_input[5276]), .Z(n22349) );
  XOR U22404 ( .A(n22741), .B(n22742), .Z(n22737) );
  AND U22405 ( .A(n22743), .B(n22744), .Z(n22742) );
  XNOR U22406 ( .A(p_input[5307]), .B(n22741), .Z(n22744) );
  XNOR U22407 ( .A(n22741), .B(n22358), .Z(n22743) );
  IV U22408 ( .A(p_input[5275]), .Z(n22358) );
  XOR U22409 ( .A(n22745), .B(n22746), .Z(n22741) );
  AND U22410 ( .A(n22747), .B(n22748), .Z(n22746) );
  XNOR U22411 ( .A(p_input[5306]), .B(n22745), .Z(n22748) );
  XNOR U22412 ( .A(n22745), .B(n22367), .Z(n22747) );
  IV U22413 ( .A(p_input[5274]), .Z(n22367) );
  XOR U22414 ( .A(n22749), .B(n22750), .Z(n22745) );
  AND U22415 ( .A(n22751), .B(n22752), .Z(n22750) );
  XNOR U22416 ( .A(p_input[5305]), .B(n22749), .Z(n22752) );
  XNOR U22417 ( .A(n22749), .B(n22376), .Z(n22751) );
  IV U22418 ( .A(p_input[5273]), .Z(n22376) );
  XOR U22419 ( .A(n22753), .B(n22754), .Z(n22749) );
  AND U22420 ( .A(n22755), .B(n22756), .Z(n22754) );
  XNOR U22421 ( .A(p_input[5304]), .B(n22753), .Z(n22756) );
  XNOR U22422 ( .A(n22753), .B(n22385), .Z(n22755) );
  IV U22423 ( .A(p_input[5272]), .Z(n22385) );
  XOR U22424 ( .A(n22757), .B(n22758), .Z(n22753) );
  AND U22425 ( .A(n22759), .B(n22760), .Z(n22758) );
  XNOR U22426 ( .A(p_input[5303]), .B(n22757), .Z(n22760) );
  XNOR U22427 ( .A(n22757), .B(n22394), .Z(n22759) );
  IV U22428 ( .A(p_input[5271]), .Z(n22394) );
  XOR U22429 ( .A(n22761), .B(n22762), .Z(n22757) );
  AND U22430 ( .A(n22763), .B(n22764), .Z(n22762) );
  XNOR U22431 ( .A(p_input[5302]), .B(n22761), .Z(n22764) );
  XNOR U22432 ( .A(n22761), .B(n22403), .Z(n22763) );
  IV U22433 ( .A(p_input[5270]), .Z(n22403) );
  XOR U22434 ( .A(n22765), .B(n22766), .Z(n22761) );
  AND U22435 ( .A(n22767), .B(n22768), .Z(n22766) );
  XNOR U22436 ( .A(p_input[5301]), .B(n22765), .Z(n22768) );
  XNOR U22437 ( .A(n22765), .B(n22412), .Z(n22767) );
  IV U22438 ( .A(p_input[5269]), .Z(n22412) );
  XOR U22439 ( .A(n22769), .B(n22770), .Z(n22765) );
  AND U22440 ( .A(n22771), .B(n22772), .Z(n22770) );
  XNOR U22441 ( .A(p_input[5300]), .B(n22769), .Z(n22772) );
  XNOR U22442 ( .A(n22769), .B(n22421), .Z(n22771) );
  IV U22443 ( .A(p_input[5268]), .Z(n22421) );
  XOR U22444 ( .A(n22773), .B(n22774), .Z(n22769) );
  AND U22445 ( .A(n22775), .B(n22776), .Z(n22774) );
  XNOR U22446 ( .A(p_input[5299]), .B(n22773), .Z(n22776) );
  XNOR U22447 ( .A(n22773), .B(n22430), .Z(n22775) );
  IV U22448 ( .A(p_input[5267]), .Z(n22430) );
  XOR U22449 ( .A(n22777), .B(n22778), .Z(n22773) );
  AND U22450 ( .A(n22779), .B(n22780), .Z(n22778) );
  XNOR U22451 ( .A(p_input[5298]), .B(n22777), .Z(n22780) );
  XNOR U22452 ( .A(n22777), .B(n22439), .Z(n22779) );
  IV U22453 ( .A(p_input[5266]), .Z(n22439) );
  XOR U22454 ( .A(n22781), .B(n22782), .Z(n22777) );
  AND U22455 ( .A(n22783), .B(n22784), .Z(n22782) );
  XNOR U22456 ( .A(p_input[5297]), .B(n22781), .Z(n22784) );
  XNOR U22457 ( .A(n22781), .B(n22448), .Z(n22783) );
  IV U22458 ( .A(p_input[5265]), .Z(n22448) );
  XOR U22459 ( .A(n22785), .B(n22786), .Z(n22781) );
  AND U22460 ( .A(n22787), .B(n22788), .Z(n22786) );
  XNOR U22461 ( .A(p_input[5296]), .B(n22785), .Z(n22788) );
  XNOR U22462 ( .A(n22785), .B(n22457), .Z(n22787) );
  IV U22463 ( .A(p_input[5264]), .Z(n22457) );
  XOR U22464 ( .A(n22789), .B(n22790), .Z(n22785) );
  AND U22465 ( .A(n22791), .B(n22792), .Z(n22790) );
  XNOR U22466 ( .A(p_input[5295]), .B(n22789), .Z(n22792) );
  XNOR U22467 ( .A(n22789), .B(n22466), .Z(n22791) );
  IV U22468 ( .A(p_input[5263]), .Z(n22466) );
  XOR U22469 ( .A(n22793), .B(n22794), .Z(n22789) );
  AND U22470 ( .A(n22795), .B(n22796), .Z(n22794) );
  XNOR U22471 ( .A(p_input[5294]), .B(n22793), .Z(n22796) );
  XNOR U22472 ( .A(n22793), .B(n22475), .Z(n22795) );
  IV U22473 ( .A(p_input[5262]), .Z(n22475) );
  XOR U22474 ( .A(n22797), .B(n22798), .Z(n22793) );
  AND U22475 ( .A(n22799), .B(n22800), .Z(n22798) );
  XNOR U22476 ( .A(p_input[5293]), .B(n22797), .Z(n22800) );
  XNOR U22477 ( .A(n22797), .B(n22484), .Z(n22799) );
  IV U22478 ( .A(p_input[5261]), .Z(n22484) );
  XOR U22479 ( .A(n22801), .B(n22802), .Z(n22797) );
  AND U22480 ( .A(n22803), .B(n22804), .Z(n22802) );
  XNOR U22481 ( .A(p_input[5292]), .B(n22801), .Z(n22804) );
  XNOR U22482 ( .A(n22801), .B(n22493), .Z(n22803) );
  IV U22483 ( .A(p_input[5260]), .Z(n22493) );
  XOR U22484 ( .A(n22805), .B(n22806), .Z(n22801) );
  AND U22485 ( .A(n22807), .B(n22808), .Z(n22806) );
  XNOR U22486 ( .A(p_input[5291]), .B(n22805), .Z(n22808) );
  XNOR U22487 ( .A(n22805), .B(n22502), .Z(n22807) );
  IV U22488 ( .A(p_input[5259]), .Z(n22502) );
  XOR U22489 ( .A(n22809), .B(n22810), .Z(n22805) );
  AND U22490 ( .A(n22811), .B(n22812), .Z(n22810) );
  XNOR U22491 ( .A(p_input[5290]), .B(n22809), .Z(n22812) );
  XNOR U22492 ( .A(n22809), .B(n22511), .Z(n22811) );
  IV U22493 ( .A(p_input[5258]), .Z(n22511) );
  XOR U22494 ( .A(n22813), .B(n22814), .Z(n22809) );
  AND U22495 ( .A(n22815), .B(n22816), .Z(n22814) );
  XNOR U22496 ( .A(p_input[5289]), .B(n22813), .Z(n22816) );
  XNOR U22497 ( .A(n22813), .B(n22520), .Z(n22815) );
  IV U22498 ( .A(p_input[5257]), .Z(n22520) );
  XOR U22499 ( .A(n22817), .B(n22818), .Z(n22813) );
  AND U22500 ( .A(n22819), .B(n22820), .Z(n22818) );
  XNOR U22501 ( .A(p_input[5288]), .B(n22817), .Z(n22820) );
  XNOR U22502 ( .A(n22817), .B(n22529), .Z(n22819) );
  IV U22503 ( .A(p_input[5256]), .Z(n22529) );
  XOR U22504 ( .A(n22821), .B(n22822), .Z(n22817) );
  AND U22505 ( .A(n22823), .B(n22824), .Z(n22822) );
  XNOR U22506 ( .A(p_input[5287]), .B(n22821), .Z(n22824) );
  XNOR U22507 ( .A(n22821), .B(n22538), .Z(n22823) );
  IV U22508 ( .A(p_input[5255]), .Z(n22538) );
  XOR U22509 ( .A(n22825), .B(n22826), .Z(n22821) );
  AND U22510 ( .A(n22827), .B(n22828), .Z(n22826) );
  XNOR U22511 ( .A(p_input[5286]), .B(n22825), .Z(n22828) );
  XNOR U22512 ( .A(n22825), .B(n22547), .Z(n22827) );
  IV U22513 ( .A(p_input[5254]), .Z(n22547) );
  XOR U22514 ( .A(n22829), .B(n22830), .Z(n22825) );
  AND U22515 ( .A(n22831), .B(n22832), .Z(n22830) );
  XNOR U22516 ( .A(p_input[5285]), .B(n22829), .Z(n22832) );
  XNOR U22517 ( .A(n22829), .B(n22556), .Z(n22831) );
  IV U22518 ( .A(p_input[5253]), .Z(n22556) );
  XOR U22519 ( .A(n22833), .B(n22834), .Z(n22829) );
  AND U22520 ( .A(n22835), .B(n22836), .Z(n22834) );
  XNOR U22521 ( .A(p_input[5284]), .B(n22833), .Z(n22836) );
  XNOR U22522 ( .A(n22833), .B(n22565), .Z(n22835) );
  IV U22523 ( .A(p_input[5252]), .Z(n22565) );
  XOR U22524 ( .A(n22837), .B(n22838), .Z(n22833) );
  AND U22525 ( .A(n22839), .B(n22840), .Z(n22838) );
  XNOR U22526 ( .A(p_input[5283]), .B(n22837), .Z(n22840) );
  XNOR U22527 ( .A(n22837), .B(n22574), .Z(n22839) );
  IV U22528 ( .A(p_input[5251]), .Z(n22574) );
  XOR U22529 ( .A(n22841), .B(n22842), .Z(n22837) );
  AND U22530 ( .A(n22843), .B(n22844), .Z(n22842) );
  XNOR U22531 ( .A(p_input[5282]), .B(n22841), .Z(n22844) );
  XNOR U22532 ( .A(n22841), .B(n22583), .Z(n22843) );
  IV U22533 ( .A(p_input[5250]), .Z(n22583) );
  XNOR U22534 ( .A(n22845), .B(n22846), .Z(n22841) );
  AND U22535 ( .A(n22847), .B(n22848), .Z(n22846) );
  XOR U22536 ( .A(p_input[5281]), .B(n22845), .Z(n22848) );
  XNOR U22537 ( .A(p_input[5249]), .B(n22845), .Z(n22847) );
  AND U22538 ( .A(p_input[5280]), .B(n22849), .Z(n22845) );
  IV U22539 ( .A(p_input[5248]), .Z(n22849) );
  XOR U22540 ( .A(n22850), .B(n22851), .Z(n21939) );
  AND U22541 ( .A(n512), .B(n22852), .Z(n22851) );
  XNOR U22542 ( .A(n22853), .B(n22850), .Z(n22852) );
  XOR U22543 ( .A(n22854), .B(n22855), .Z(n512) );
  AND U22544 ( .A(n22856), .B(n22857), .Z(n22855) );
  XNOR U22545 ( .A(n21954), .B(n22854), .Z(n22857) );
  AND U22546 ( .A(p_input[5247]), .B(p_input[5215]), .Z(n21954) );
  XNOR U22547 ( .A(n22854), .B(n21951), .Z(n22856) );
  IV U22548 ( .A(n22858), .Z(n21951) );
  AND U22549 ( .A(p_input[5151]), .B(p_input[5183]), .Z(n22858) );
  XOR U22550 ( .A(n22859), .B(n22860), .Z(n22854) );
  AND U22551 ( .A(n22861), .B(n22862), .Z(n22860) );
  XOR U22552 ( .A(n22859), .B(n21966), .Z(n22862) );
  XNOR U22553 ( .A(p_input[5214]), .B(n22863), .Z(n21966) );
  AND U22554 ( .A(n355), .B(n22864), .Z(n22863) );
  XOR U22555 ( .A(p_input[5246]), .B(p_input[5214]), .Z(n22864) );
  XNOR U22556 ( .A(n21963), .B(n22859), .Z(n22861) );
  XOR U22557 ( .A(n22865), .B(n22866), .Z(n21963) );
  AND U22558 ( .A(n352), .B(n22867), .Z(n22866) );
  XOR U22559 ( .A(p_input[5182]), .B(p_input[5150]), .Z(n22867) );
  XOR U22560 ( .A(n22868), .B(n22869), .Z(n22859) );
  AND U22561 ( .A(n22870), .B(n22871), .Z(n22869) );
  XOR U22562 ( .A(n22868), .B(n21978), .Z(n22871) );
  XNOR U22563 ( .A(p_input[5213]), .B(n22872), .Z(n21978) );
  AND U22564 ( .A(n355), .B(n22873), .Z(n22872) );
  XOR U22565 ( .A(p_input[5245]), .B(p_input[5213]), .Z(n22873) );
  XNOR U22566 ( .A(n21975), .B(n22868), .Z(n22870) );
  XOR U22567 ( .A(n22874), .B(n22875), .Z(n21975) );
  AND U22568 ( .A(n352), .B(n22876), .Z(n22875) );
  XOR U22569 ( .A(p_input[5181]), .B(p_input[5149]), .Z(n22876) );
  XOR U22570 ( .A(n22877), .B(n22878), .Z(n22868) );
  AND U22571 ( .A(n22879), .B(n22880), .Z(n22878) );
  XOR U22572 ( .A(n22877), .B(n21990), .Z(n22880) );
  XNOR U22573 ( .A(p_input[5212]), .B(n22881), .Z(n21990) );
  AND U22574 ( .A(n355), .B(n22882), .Z(n22881) );
  XOR U22575 ( .A(p_input[5244]), .B(p_input[5212]), .Z(n22882) );
  XNOR U22576 ( .A(n21987), .B(n22877), .Z(n22879) );
  XOR U22577 ( .A(n22883), .B(n22884), .Z(n21987) );
  AND U22578 ( .A(n352), .B(n22885), .Z(n22884) );
  XOR U22579 ( .A(p_input[5180]), .B(p_input[5148]), .Z(n22885) );
  XOR U22580 ( .A(n22886), .B(n22887), .Z(n22877) );
  AND U22581 ( .A(n22888), .B(n22889), .Z(n22887) );
  XOR U22582 ( .A(n22886), .B(n22002), .Z(n22889) );
  XNOR U22583 ( .A(p_input[5211]), .B(n22890), .Z(n22002) );
  AND U22584 ( .A(n355), .B(n22891), .Z(n22890) );
  XOR U22585 ( .A(p_input[5243]), .B(p_input[5211]), .Z(n22891) );
  XNOR U22586 ( .A(n21999), .B(n22886), .Z(n22888) );
  XOR U22587 ( .A(n22892), .B(n22893), .Z(n21999) );
  AND U22588 ( .A(n352), .B(n22894), .Z(n22893) );
  XOR U22589 ( .A(p_input[5179]), .B(p_input[5147]), .Z(n22894) );
  XOR U22590 ( .A(n22895), .B(n22896), .Z(n22886) );
  AND U22591 ( .A(n22897), .B(n22898), .Z(n22896) );
  XOR U22592 ( .A(n22895), .B(n22014), .Z(n22898) );
  XNOR U22593 ( .A(p_input[5210]), .B(n22899), .Z(n22014) );
  AND U22594 ( .A(n355), .B(n22900), .Z(n22899) );
  XOR U22595 ( .A(p_input[5242]), .B(p_input[5210]), .Z(n22900) );
  XNOR U22596 ( .A(n22011), .B(n22895), .Z(n22897) );
  XOR U22597 ( .A(n22901), .B(n22902), .Z(n22011) );
  AND U22598 ( .A(n352), .B(n22903), .Z(n22902) );
  XOR U22599 ( .A(p_input[5178]), .B(p_input[5146]), .Z(n22903) );
  XOR U22600 ( .A(n22904), .B(n22905), .Z(n22895) );
  AND U22601 ( .A(n22906), .B(n22907), .Z(n22905) );
  XOR U22602 ( .A(n22904), .B(n22026), .Z(n22907) );
  XNOR U22603 ( .A(p_input[5209]), .B(n22908), .Z(n22026) );
  AND U22604 ( .A(n355), .B(n22909), .Z(n22908) );
  XOR U22605 ( .A(p_input[5241]), .B(p_input[5209]), .Z(n22909) );
  XNOR U22606 ( .A(n22023), .B(n22904), .Z(n22906) );
  XOR U22607 ( .A(n22910), .B(n22911), .Z(n22023) );
  AND U22608 ( .A(n352), .B(n22912), .Z(n22911) );
  XOR U22609 ( .A(p_input[5177]), .B(p_input[5145]), .Z(n22912) );
  XOR U22610 ( .A(n22913), .B(n22914), .Z(n22904) );
  AND U22611 ( .A(n22915), .B(n22916), .Z(n22914) );
  XOR U22612 ( .A(n22913), .B(n22038), .Z(n22916) );
  XNOR U22613 ( .A(p_input[5208]), .B(n22917), .Z(n22038) );
  AND U22614 ( .A(n355), .B(n22918), .Z(n22917) );
  XOR U22615 ( .A(p_input[5240]), .B(p_input[5208]), .Z(n22918) );
  XNOR U22616 ( .A(n22035), .B(n22913), .Z(n22915) );
  XOR U22617 ( .A(n22919), .B(n22920), .Z(n22035) );
  AND U22618 ( .A(n352), .B(n22921), .Z(n22920) );
  XOR U22619 ( .A(p_input[5176]), .B(p_input[5144]), .Z(n22921) );
  XOR U22620 ( .A(n22922), .B(n22923), .Z(n22913) );
  AND U22621 ( .A(n22924), .B(n22925), .Z(n22923) );
  XOR U22622 ( .A(n22922), .B(n22050), .Z(n22925) );
  XNOR U22623 ( .A(p_input[5207]), .B(n22926), .Z(n22050) );
  AND U22624 ( .A(n355), .B(n22927), .Z(n22926) );
  XOR U22625 ( .A(p_input[5239]), .B(p_input[5207]), .Z(n22927) );
  XNOR U22626 ( .A(n22047), .B(n22922), .Z(n22924) );
  XOR U22627 ( .A(n22928), .B(n22929), .Z(n22047) );
  AND U22628 ( .A(n352), .B(n22930), .Z(n22929) );
  XOR U22629 ( .A(p_input[5175]), .B(p_input[5143]), .Z(n22930) );
  XOR U22630 ( .A(n22931), .B(n22932), .Z(n22922) );
  AND U22631 ( .A(n22933), .B(n22934), .Z(n22932) );
  XOR U22632 ( .A(n22931), .B(n22062), .Z(n22934) );
  XNOR U22633 ( .A(p_input[5206]), .B(n22935), .Z(n22062) );
  AND U22634 ( .A(n355), .B(n22936), .Z(n22935) );
  XOR U22635 ( .A(p_input[5238]), .B(p_input[5206]), .Z(n22936) );
  XNOR U22636 ( .A(n22059), .B(n22931), .Z(n22933) );
  XOR U22637 ( .A(n22937), .B(n22938), .Z(n22059) );
  AND U22638 ( .A(n352), .B(n22939), .Z(n22938) );
  XOR U22639 ( .A(p_input[5174]), .B(p_input[5142]), .Z(n22939) );
  XOR U22640 ( .A(n22940), .B(n22941), .Z(n22931) );
  AND U22641 ( .A(n22942), .B(n22943), .Z(n22941) );
  XOR U22642 ( .A(n22940), .B(n22074), .Z(n22943) );
  XNOR U22643 ( .A(p_input[5205]), .B(n22944), .Z(n22074) );
  AND U22644 ( .A(n355), .B(n22945), .Z(n22944) );
  XOR U22645 ( .A(p_input[5237]), .B(p_input[5205]), .Z(n22945) );
  XNOR U22646 ( .A(n22071), .B(n22940), .Z(n22942) );
  XOR U22647 ( .A(n22946), .B(n22947), .Z(n22071) );
  AND U22648 ( .A(n352), .B(n22948), .Z(n22947) );
  XOR U22649 ( .A(p_input[5173]), .B(p_input[5141]), .Z(n22948) );
  XOR U22650 ( .A(n22949), .B(n22950), .Z(n22940) );
  AND U22651 ( .A(n22951), .B(n22952), .Z(n22950) );
  XOR U22652 ( .A(n22949), .B(n22086), .Z(n22952) );
  XNOR U22653 ( .A(p_input[5204]), .B(n22953), .Z(n22086) );
  AND U22654 ( .A(n355), .B(n22954), .Z(n22953) );
  XOR U22655 ( .A(p_input[5236]), .B(p_input[5204]), .Z(n22954) );
  XNOR U22656 ( .A(n22083), .B(n22949), .Z(n22951) );
  XOR U22657 ( .A(n22955), .B(n22956), .Z(n22083) );
  AND U22658 ( .A(n352), .B(n22957), .Z(n22956) );
  XOR U22659 ( .A(p_input[5172]), .B(p_input[5140]), .Z(n22957) );
  XOR U22660 ( .A(n22958), .B(n22959), .Z(n22949) );
  AND U22661 ( .A(n22960), .B(n22961), .Z(n22959) );
  XOR U22662 ( .A(n22958), .B(n22098), .Z(n22961) );
  XNOR U22663 ( .A(p_input[5203]), .B(n22962), .Z(n22098) );
  AND U22664 ( .A(n355), .B(n22963), .Z(n22962) );
  XOR U22665 ( .A(p_input[5235]), .B(p_input[5203]), .Z(n22963) );
  XNOR U22666 ( .A(n22095), .B(n22958), .Z(n22960) );
  XOR U22667 ( .A(n22964), .B(n22965), .Z(n22095) );
  AND U22668 ( .A(n352), .B(n22966), .Z(n22965) );
  XOR U22669 ( .A(p_input[5171]), .B(p_input[5139]), .Z(n22966) );
  XOR U22670 ( .A(n22967), .B(n22968), .Z(n22958) );
  AND U22671 ( .A(n22969), .B(n22970), .Z(n22968) );
  XOR U22672 ( .A(n22967), .B(n22110), .Z(n22970) );
  XNOR U22673 ( .A(p_input[5202]), .B(n22971), .Z(n22110) );
  AND U22674 ( .A(n355), .B(n22972), .Z(n22971) );
  XOR U22675 ( .A(p_input[5234]), .B(p_input[5202]), .Z(n22972) );
  XNOR U22676 ( .A(n22107), .B(n22967), .Z(n22969) );
  XOR U22677 ( .A(n22973), .B(n22974), .Z(n22107) );
  AND U22678 ( .A(n352), .B(n22975), .Z(n22974) );
  XOR U22679 ( .A(p_input[5170]), .B(p_input[5138]), .Z(n22975) );
  XOR U22680 ( .A(n22976), .B(n22977), .Z(n22967) );
  AND U22681 ( .A(n22978), .B(n22979), .Z(n22977) );
  XOR U22682 ( .A(n22976), .B(n22122), .Z(n22979) );
  XNOR U22683 ( .A(p_input[5201]), .B(n22980), .Z(n22122) );
  AND U22684 ( .A(n355), .B(n22981), .Z(n22980) );
  XOR U22685 ( .A(p_input[5233]), .B(p_input[5201]), .Z(n22981) );
  XNOR U22686 ( .A(n22119), .B(n22976), .Z(n22978) );
  XOR U22687 ( .A(n22982), .B(n22983), .Z(n22119) );
  AND U22688 ( .A(n352), .B(n22984), .Z(n22983) );
  XOR U22689 ( .A(p_input[5169]), .B(p_input[5137]), .Z(n22984) );
  XOR U22690 ( .A(n22985), .B(n22986), .Z(n22976) );
  AND U22691 ( .A(n22987), .B(n22988), .Z(n22986) );
  XOR U22692 ( .A(n22985), .B(n22134), .Z(n22988) );
  XNOR U22693 ( .A(p_input[5200]), .B(n22989), .Z(n22134) );
  AND U22694 ( .A(n355), .B(n22990), .Z(n22989) );
  XOR U22695 ( .A(p_input[5232]), .B(p_input[5200]), .Z(n22990) );
  XNOR U22696 ( .A(n22131), .B(n22985), .Z(n22987) );
  XOR U22697 ( .A(n22991), .B(n22992), .Z(n22131) );
  AND U22698 ( .A(n352), .B(n22993), .Z(n22992) );
  XOR U22699 ( .A(p_input[5168]), .B(p_input[5136]), .Z(n22993) );
  XOR U22700 ( .A(n22994), .B(n22995), .Z(n22985) );
  AND U22701 ( .A(n22996), .B(n22997), .Z(n22995) );
  XOR U22702 ( .A(n22994), .B(n22146), .Z(n22997) );
  XNOR U22703 ( .A(p_input[5199]), .B(n22998), .Z(n22146) );
  AND U22704 ( .A(n355), .B(n22999), .Z(n22998) );
  XOR U22705 ( .A(p_input[5231]), .B(p_input[5199]), .Z(n22999) );
  XNOR U22706 ( .A(n22143), .B(n22994), .Z(n22996) );
  XOR U22707 ( .A(n23000), .B(n23001), .Z(n22143) );
  AND U22708 ( .A(n352), .B(n23002), .Z(n23001) );
  XOR U22709 ( .A(p_input[5167]), .B(p_input[5135]), .Z(n23002) );
  XOR U22710 ( .A(n23003), .B(n23004), .Z(n22994) );
  AND U22711 ( .A(n23005), .B(n23006), .Z(n23004) );
  XOR U22712 ( .A(n23003), .B(n22158), .Z(n23006) );
  XNOR U22713 ( .A(p_input[5198]), .B(n23007), .Z(n22158) );
  AND U22714 ( .A(n355), .B(n23008), .Z(n23007) );
  XOR U22715 ( .A(p_input[5230]), .B(p_input[5198]), .Z(n23008) );
  XNOR U22716 ( .A(n22155), .B(n23003), .Z(n23005) );
  XOR U22717 ( .A(n23009), .B(n23010), .Z(n22155) );
  AND U22718 ( .A(n352), .B(n23011), .Z(n23010) );
  XOR U22719 ( .A(p_input[5166]), .B(p_input[5134]), .Z(n23011) );
  XOR U22720 ( .A(n23012), .B(n23013), .Z(n23003) );
  AND U22721 ( .A(n23014), .B(n23015), .Z(n23013) );
  XOR U22722 ( .A(n23012), .B(n22170), .Z(n23015) );
  XNOR U22723 ( .A(p_input[5197]), .B(n23016), .Z(n22170) );
  AND U22724 ( .A(n355), .B(n23017), .Z(n23016) );
  XOR U22725 ( .A(p_input[5229]), .B(p_input[5197]), .Z(n23017) );
  XNOR U22726 ( .A(n22167), .B(n23012), .Z(n23014) );
  XOR U22727 ( .A(n23018), .B(n23019), .Z(n22167) );
  AND U22728 ( .A(n352), .B(n23020), .Z(n23019) );
  XOR U22729 ( .A(p_input[5165]), .B(p_input[5133]), .Z(n23020) );
  XOR U22730 ( .A(n23021), .B(n23022), .Z(n23012) );
  AND U22731 ( .A(n23023), .B(n23024), .Z(n23022) );
  XOR U22732 ( .A(n23021), .B(n22182), .Z(n23024) );
  XNOR U22733 ( .A(p_input[5196]), .B(n23025), .Z(n22182) );
  AND U22734 ( .A(n355), .B(n23026), .Z(n23025) );
  XOR U22735 ( .A(p_input[5228]), .B(p_input[5196]), .Z(n23026) );
  XNOR U22736 ( .A(n22179), .B(n23021), .Z(n23023) );
  XOR U22737 ( .A(n23027), .B(n23028), .Z(n22179) );
  AND U22738 ( .A(n352), .B(n23029), .Z(n23028) );
  XOR U22739 ( .A(p_input[5164]), .B(p_input[5132]), .Z(n23029) );
  XOR U22740 ( .A(n23030), .B(n23031), .Z(n23021) );
  AND U22741 ( .A(n23032), .B(n23033), .Z(n23031) );
  XOR U22742 ( .A(n23030), .B(n22194), .Z(n23033) );
  XNOR U22743 ( .A(p_input[5195]), .B(n23034), .Z(n22194) );
  AND U22744 ( .A(n355), .B(n23035), .Z(n23034) );
  XOR U22745 ( .A(p_input[5227]), .B(p_input[5195]), .Z(n23035) );
  XNOR U22746 ( .A(n22191), .B(n23030), .Z(n23032) );
  XOR U22747 ( .A(n23036), .B(n23037), .Z(n22191) );
  AND U22748 ( .A(n352), .B(n23038), .Z(n23037) );
  XOR U22749 ( .A(p_input[5163]), .B(p_input[5131]), .Z(n23038) );
  XOR U22750 ( .A(n23039), .B(n23040), .Z(n23030) );
  AND U22751 ( .A(n23041), .B(n23042), .Z(n23040) );
  XOR U22752 ( .A(n23039), .B(n22206), .Z(n23042) );
  XNOR U22753 ( .A(p_input[5194]), .B(n23043), .Z(n22206) );
  AND U22754 ( .A(n355), .B(n23044), .Z(n23043) );
  XOR U22755 ( .A(p_input[5226]), .B(p_input[5194]), .Z(n23044) );
  XNOR U22756 ( .A(n22203), .B(n23039), .Z(n23041) );
  XOR U22757 ( .A(n23045), .B(n23046), .Z(n22203) );
  AND U22758 ( .A(n352), .B(n23047), .Z(n23046) );
  XOR U22759 ( .A(p_input[5162]), .B(p_input[5130]), .Z(n23047) );
  XOR U22760 ( .A(n23048), .B(n23049), .Z(n23039) );
  AND U22761 ( .A(n23050), .B(n23051), .Z(n23049) );
  XOR U22762 ( .A(n23048), .B(n22218), .Z(n23051) );
  XNOR U22763 ( .A(p_input[5193]), .B(n23052), .Z(n22218) );
  AND U22764 ( .A(n355), .B(n23053), .Z(n23052) );
  XOR U22765 ( .A(p_input[5225]), .B(p_input[5193]), .Z(n23053) );
  XNOR U22766 ( .A(n22215), .B(n23048), .Z(n23050) );
  XOR U22767 ( .A(n23054), .B(n23055), .Z(n22215) );
  AND U22768 ( .A(n352), .B(n23056), .Z(n23055) );
  XOR U22769 ( .A(p_input[5161]), .B(p_input[5129]), .Z(n23056) );
  XOR U22770 ( .A(n23057), .B(n23058), .Z(n23048) );
  AND U22771 ( .A(n23059), .B(n23060), .Z(n23058) );
  XOR U22772 ( .A(n23057), .B(n22230), .Z(n23060) );
  XNOR U22773 ( .A(p_input[5192]), .B(n23061), .Z(n22230) );
  AND U22774 ( .A(n355), .B(n23062), .Z(n23061) );
  XOR U22775 ( .A(p_input[5224]), .B(p_input[5192]), .Z(n23062) );
  XNOR U22776 ( .A(n22227), .B(n23057), .Z(n23059) );
  XOR U22777 ( .A(n23063), .B(n23064), .Z(n22227) );
  AND U22778 ( .A(n352), .B(n23065), .Z(n23064) );
  XOR U22779 ( .A(p_input[5160]), .B(p_input[5128]), .Z(n23065) );
  XOR U22780 ( .A(n23066), .B(n23067), .Z(n23057) );
  AND U22781 ( .A(n23068), .B(n23069), .Z(n23067) );
  XOR U22782 ( .A(n23066), .B(n22242), .Z(n23069) );
  XNOR U22783 ( .A(p_input[5191]), .B(n23070), .Z(n22242) );
  AND U22784 ( .A(n355), .B(n23071), .Z(n23070) );
  XOR U22785 ( .A(p_input[5223]), .B(p_input[5191]), .Z(n23071) );
  XNOR U22786 ( .A(n22239), .B(n23066), .Z(n23068) );
  XOR U22787 ( .A(n23072), .B(n23073), .Z(n22239) );
  AND U22788 ( .A(n352), .B(n23074), .Z(n23073) );
  XOR U22789 ( .A(p_input[5159]), .B(p_input[5127]), .Z(n23074) );
  XOR U22790 ( .A(n23075), .B(n23076), .Z(n23066) );
  AND U22791 ( .A(n23077), .B(n23078), .Z(n23076) );
  XOR U22792 ( .A(n23075), .B(n22254), .Z(n23078) );
  XNOR U22793 ( .A(p_input[5190]), .B(n23079), .Z(n22254) );
  AND U22794 ( .A(n355), .B(n23080), .Z(n23079) );
  XOR U22795 ( .A(p_input[5222]), .B(p_input[5190]), .Z(n23080) );
  XNOR U22796 ( .A(n22251), .B(n23075), .Z(n23077) );
  XOR U22797 ( .A(n23081), .B(n23082), .Z(n22251) );
  AND U22798 ( .A(n352), .B(n23083), .Z(n23082) );
  XOR U22799 ( .A(p_input[5158]), .B(p_input[5126]), .Z(n23083) );
  XOR U22800 ( .A(n23084), .B(n23085), .Z(n23075) );
  AND U22801 ( .A(n23086), .B(n23087), .Z(n23085) );
  XOR U22802 ( .A(n23084), .B(n22266), .Z(n23087) );
  XNOR U22803 ( .A(p_input[5189]), .B(n23088), .Z(n22266) );
  AND U22804 ( .A(n355), .B(n23089), .Z(n23088) );
  XOR U22805 ( .A(p_input[5221]), .B(p_input[5189]), .Z(n23089) );
  XNOR U22806 ( .A(n22263), .B(n23084), .Z(n23086) );
  XOR U22807 ( .A(n23090), .B(n23091), .Z(n22263) );
  AND U22808 ( .A(n352), .B(n23092), .Z(n23091) );
  XOR U22809 ( .A(p_input[5157]), .B(p_input[5125]), .Z(n23092) );
  XOR U22810 ( .A(n23093), .B(n23094), .Z(n23084) );
  AND U22811 ( .A(n23095), .B(n23096), .Z(n23094) );
  XOR U22812 ( .A(n23093), .B(n22278), .Z(n23096) );
  XNOR U22813 ( .A(p_input[5188]), .B(n23097), .Z(n22278) );
  AND U22814 ( .A(n355), .B(n23098), .Z(n23097) );
  XOR U22815 ( .A(p_input[5220]), .B(p_input[5188]), .Z(n23098) );
  XNOR U22816 ( .A(n22275), .B(n23093), .Z(n23095) );
  XOR U22817 ( .A(n23099), .B(n23100), .Z(n22275) );
  AND U22818 ( .A(n352), .B(n23101), .Z(n23100) );
  XOR U22819 ( .A(p_input[5156]), .B(p_input[5124]), .Z(n23101) );
  XOR U22820 ( .A(n23102), .B(n23103), .Z(n23093) );
  AND U22821 ( .A(n23104), .B(n23105), .Z(n23103) );
  XOR U22822 ( .A(n23102), .B(n22290), .Z(n23105) );
  XNOR U22823 ( .A(p_input[5187]), .B(n23106), .Z(n22290) );
  AND U22824 ( .A(n355), .B(n23107), .Z(n23106) );
  XOR U22825 ( .A(p_input[5219]), .B(p_input[5187]), .Z(n23107) );
  XNOR U22826 ( .A(n22287), .B(n23102), .Z(n23104) );
  XOR U22827 ( .A(n23108), .B(n23109), .Z(n22287) );
  AND U22828 ( .A(n352), .B(n23110), .Z(n23109) );
  XOR U22829 ( .A(p_input[5155]), .B(p_input[5123]), .Z(n23110) );
  XOR U22830 ( .A(n23111), .B(n23112), .Z(n23102) );
  AND U22831 ( .A(n23113), .B(n23114), .Z(n23112) );
  XOR U22832 ( .A(n23111), .B(n22302), .Z(n23114) );
  XNOR U22833 ( .A(p_input[5186]), .B(n23115), .Z(n22302) );
  AND U22834 ( .A(n355), .B(n23116), .Z(n23115) );
  XOR U22835 ( .A(p_input[5218]), .B(p_input[5186]), .Z(n23116) );
  XNOR U22836 ( .A(n22299), .B(n23111), .Z(n23113) );
  XOR U22837 ( .A(n23117), .B(n23118), .Z(n22299) );
  AND U22838 ( .A(n352), .B(n23119), .Z(n23118) );
  XOR U22839 ( .A(p_input[5154]), .B(p_input[5122]), .Z(n23119) );
  XOR U22840 ( .A(n23120), .B(n23121), .Z(n23111) );
  AND U22841 ( .A(n23122), .B(n23123), .Z(n23121) );
  XNOR U22842 ( .A(n23124), .B(n22315), .Z(n23123) );
  XNOR U22843 ( .A(p_input[5185]), .B(n23125), .Z(n22315) );
  AND U22844 ( .A(n355), .B(n23126), .Z(n23125) );
  XNOR U22845 ( .A(p_input[5217]), .B(n23127), .Z(n23126) );
  IV U22846 ( .A(p_input[5185]), .Z(n23127) );
  XNOR U22847 ( .A(n22312), .B(n23120), .Z(n23122) );
  XNOR U22848 ( .A(p_input[5121]), .B(n23128), .Z(n22312) );
  AND U22849 ( .A(n352), .B(n23129), .Z(n23128) );
  XOR U22850 ( .A(p_input[5153]), .B(p_input[5121]), .Z(n23129) );
  IV U22851 ( .A(n23124), .Z(n23120) );
  AND U22852 ( .A(n22850), .B(n22853), .Z(n23124) );
  XOR U22853 ( .A(p_input[5184]), .B(n23130), .Z(n22853) );
  AND U22854 ( .A(n355), .B(n23131), .Z(n23130) );
  XOR U22855 ( .A(p_input[5216]), .B(p_input[5184]), .Z(n23131) );
  XOR U22856 ( .A(n23132), .B(n23133), .Z(n355) );
  AND U22857 ( .A(n23134), .B(n23135), .Z(n23133) );
  XNOR U22858 ( .A(p_input[5247]), .B(n23132), .Z(n23135) );
  XOR U22859 ( .A(n23132), .B(p_input[5215]), .Z(n23134) );
  XOR U22860 ( .A(n23136), .B(n23137), .Z(n23132) );
  AND U22861 ( .A(n23138), .B(n23139), .Z(n23137) );
  XNOR U22862 ( .A(p_input[5246]), .B(n23136), .Z(n23139) );
  XOR U22863 ( .A(n23136), .B(p_input[5214]), .Z(n23138) );
  XOR U22864 ( .A(n23140), .B(n23141), .Z(n23136) );
  AND U22865 ( .A(n23142), .B(n23143), .Z(n23141) );
  XNOR U22866 ( .A(p_input[5245]), .B(n23140), .Z(n23143) );
  XOR U22867 ( .A(n23140), .B(p_input[5213]), .Z(n23142) );
  XOR U22868 ( .A(n23144), .B(n23145), .Z(n23140) );
  AND U22869 ( .A(n23146), .B(n23147), .Z(n23145) );
  XNOR U22870 ( .A(p_input[5244]), .B(n23144), .Z(n23147) );
  XOR U22871 ( .A(n23144), .B(p_input[5212]), .Z(n23146) );
  XOR U22872 ( .A(n23148), .B(n23149), .Z(n23144) );
  AND U22873 ( .A(n23150), .B(n23151), .Z(n23149) );
  XNOR U22874 ( .A(p_input[5243]), .B(n23148), .Z(n23151) );
  XOR U22875 ( .A(n23148), .B(p_input[5211]), .Z(n23150) );
  XOR U22876 ( .A(n23152), .B(n23153), .Z(n23148) );
  AND U22877 ( .A(n23154), .B(n23155), .Z(n23153) );
  XNOR U22878 ( .A(p_input[5242]), .B(n23152), .Z(n23155) );
  XOR U22879 ( .A(n23152), .B(p_input[5210]), .Z(n23154) );
  XOR U22880 ( .A(n23156), .B(n23157), .Z(n23152) );
  AND U22881 ( .A(n23158), .B(n23159), .Z(n23157) );
  XNOR U22882 ( .A(p_input[5241]), .B(n23156), .Z(n23159) );
  XOR U22883 ( .A(n23156), .B(p_input[5209]), .Z(n23158) );
  XOR U22884 ( .A(n23160), .B(n23161), .Z(n23156) );
  AND U22885 ( .A(n23162), .B(n23163), .Z(n23161) );
  XNOR U22886 ( .A(p_input[5240]), .B(n23160), .Z(n23163) );
  XOR U22887 ( .A(n23160), .B(p_input[5208]), .Z(n23162) );
  XOR U22888 ( .A(n23164), .B(n23165), .Z(n23160) );
  AND U22889 ( .A(n23166), .B(n23167), .Z(n23165) );
  XNOR U22890 ( .A(p_input[5239]), .B(n23164), .Z(n23167) );
  XOR U22891 ( .A(n23164), .B(p_input[5207]), .Z(n23166) );
  XOR U22892 ( .A(n23168), .B(n23169), .Z(n23164) );
  AND U22893 ( .A(n23170), .B(n23171), .Z(n23169) );
  XNOR U22894 ( .A(p_input[5238]), .B(n23168), .Z(n23171) );
  XOR U22895 ( .A(n23168), .B(p_input[5206]), .Z(n23170) );
  XOR U22896 ( .A(n23172), .B(n23173), .Z(n23168) );
  AND U22897 ( .A(n23174), .B(n23175), .Z(n23173) );
  XNOR U22898 ( .A(p_input[5237]), .B(n23172), .Z(n23175) );
  XOR U22899 ( .A(n23172), .B(p_input[5205]), .Z(n23174) );
  XOR U22900 ( .A(n23176), .B(n23177), .Z(n23172) );
  AND U22901 ( .A(n23178), .B(n23179), .Z(n23177) );
  XNOR U22902 ( .A(p_input[5236]), .B(n23176), .Z(n23179) );
  XOR U22903 ( .A(n23176), .B(p_input[5204]), .Z(n23178) );
  XOR U22904 ( .A(n23180), .B(n23181), .Z(n23176) );
  AND U22905 ( .A(n23182), .B(n23183), .Z(n23181) );
  XNOR U22906 ( .A(p_input[5235]), .B(n23180), .Z(n23183) );
  XOR U22907 ( .A(n23180), .B(p_input[5203]), .Z(n23182) );
  XOR U22908 ( .A(n23184), .B(n23185), .Z(n23180) );
  AND U22909 ( .A(n23186), .B(n23187), .Z(n23185) );
  XNOR U22910 ( .A(p_input[5234]), .B(n23184), .Z(n23187) );
  XOR U22911 ( .A(n23184), .B(p_input[5202]), .Z(n23186) );
  XOR U22912 ( .A(n23188), .B(n23189), .Z(n23184) );
  AND U22913 ( .A(n23190), .B(n23191), .Z(n23189) );
  XNOR U22914 ( .A(p_input[5233]), .B(n23188), .Z(n23191) );
  XOR U22915 ( .A(n23188), .B(p_input[5201]), .Z(n23190) );
  XOR U22916 ( .A(n23192), .B(n23193), .Z(n23188) );
  AND U22917 ( .A(n23194), .B(n23195), .Z(n23193) );
  XNOR U22918 ( .A(p_input[5232]), .B(n23192), .Z(n23195) );
  XOR U22919 ( .A(n23192), .B(p_input[5200]), .Z(n23194) );
  XOR U22920 ( .A(n23196), .B(n23197), .Z(n23192) );
  AND U22921 ( .A(n23198), .B(n23199), .Z(n23197) );
  XNOR U22922 ( .A(p_input[5231]), .B(n23196), .Z(n23199) );
  XOR U22923 ( .A(n23196), .B(p_input[5199]), .Z(n23198) );
  XOR U22924 ( .A(n23200), .B(n23201), .Z(n23196) );
  AND U22925 ( .A(n23202), .B(n23203), .Z(n23201) );
  XNOR U22926 ( .A(p_input[5230]), .B(n23200), .Z(n23203) );
  XOR U22927 ( .A(n23200), .B(p_input[5198]), .Z(n23202) );
  XOR U22928 ( .A(n23204), .B(n23205), .Z(n23200) );
  AND U22929 ( .A(n23206), .B(n23207), .Z(n23205) );
  XNOR U22930 ( .A(p_input[5229]), .B(n23204), .Z(n23207) );
  XOR U22931 ( .A(n23204), .B(p_input[5197]), .Z(n23206) );
  XOR U22932 ( .A(n23208), .B(n23209), .Z(n23204) );
  AND U22933 ( .A(n23210), .B(n23211), .Z(n23209) );
  XNOR U22934 ( .A(p_input[5228]), .B(n23208), .Z(n23211) );
  XOR U22935 ( .A(n23208), .B(p_input[5196]), .Z(n23210) );
  XOR U22936 ( .A(n23212), .B(n23213), .Z(n23208) );
  AND U22937 ( .A(n23214), .B(n23215), .Z(n23213) );
  XNOR U22938 ( .A(p_input[5227]), .B(n23212), .Z(n23215) );
  XOR U22939 ( .A(n23212), .B(p_input[5195]), .Z(n23214) );
  XOR U22940 ( .A(n23216), .B(n23217), .Z(n23212) );
  AND U22941 ( .A(n23218), .B(n23219), .Z(n23217) );
  XNOR U22942 ( .A(p_input[5226]), .B(n23216), .Z(n23219) );
  XOR U22943 ( .A(n23216), .B(p_input[5194]), .Z(n23218) );
  XOR U22944 ( .A(n23220), .B(n23221), .Z(n23216) );
  AND U22945 ( .A(n23222), .B(n23223), .Z(n23221) );
  XNOR U22946 ( .A(p_input[5225]), .B(n23220), .Z(n23223) );
  XOR U22947 ( .A(n23220), .B(p_input[5193]), .Z(n23222) );
  XOR U22948 ( .A(n23224), .B(n23225), .Z(n23220) );
  AND U22949 ( .A(n23226), .B(n23227), .Z(n23225) );
  XNOR U22950 ( .A(p_input[5224]), .B(n23224), .Z(n23227) );
  XOR U22951 ( .A(n23224), .B(p_input[5192]), .Z(n23226) );
  XOR U22952 ( .A(n23228), .B(n23229), .Z(n23224) );
  AND U22953 ( .A(n23230), .B(n23231), .Z(n23229) );
  XNOR U22954 ( .A(p_input[5223]), .B(n23228), .Z(n23231) );
  XOR U22955 ( .A(n23228), .B(p_input[5191]), .Z(n23230) );
  XOR U22956 ( .A(n23232), .B(n23233), .Z(n23228) );
  AND U22957 ( .A(n23234), .B(n23235), .Z(n23233) );
  XNOR U22958 ( .A(p_input[5222]), .B(n23232), .Z(n23235) );
  XOR U22959 ( .A(n23232), .B(p_input[5190]), .Z(n23234) );
  XOR U22960 ( .A(n23236), .B(n23237), .Z(n23232) );
  AND U22961 ( .A(n23238), .B(n23239), .Z(n23237) );
  XNOR U22962 ( .A(p_input[5221]), .B(n23236), .Z(n23239) );
  XOR U22963 ( .A(n23236), .B(p_input[5189]), .Z(n23238) );
  XOR U22964 ( .A(n23240), .B(n23241), .Z(n23236) );
  AND U22965 ( .A(n23242), .B(n23243), .Z(n23241) );
  XNOR U22966 ( .A(p_input[5220]), .B(n23240), .Z(n23243) );
  XOR U22967 ( .A(n23240), .B(p_input[5188]), .Z(n23242) );
  XOR U22968 ( .A(n23244), .B(n23245), .Z(n23240) );
  AND U22969 ( .A(n23246), .B(n23247), .Z(n23245) );
  XNOR U22970 ( .A(p_input[5219]), .B(n23244), .Z(n23247) );
  XOR U22971 ( .A(n23244), .B(p_input[5187]), .Z(n23246) );
  XOR U22972 ( .A(n23248), .B(n23249), .Z(n23244) );
  AND U22973 ( .A(n23250), .B(n23251), .Z(n23249) );
  XNOR U22974 ( .A(p_input[5218]), .B(n23248), .Z(n23251) );
  XOR U22975 ( .A(n23248), .B(p_input[5186]), .Z(n23250) );
  XNOR U22976 ( .A(n23252), .B(n23253), .Z(n23248) );
  AND U22977 ( .A(n23254), .B(n23255), .Z(n23253) );
  XOR U22978 ( .A(p_input[5217]), .B(n23252), .Z(n23255) );
  XNOR U22979 ( .A(p_input[5185]), .B(n23252), .Z(n23254) );
  AND U22980 ( .A(p_input[5216]), .B(n23256), .Z(n23252) );
  IV U22981 ( .A(p_input[5184]), .Z(n23256) );
  XNOR U22982 ( .A(p_input[5120]), .B(n23257), .Z(n22850) );
  AND U22983 ( .A(n352), .B(n23258), .Z(n23257) );
  XOR U22984 ( .A(p_input[5152]), .B(p_input[5120]), .Z(n23258) );
  XOR U22985 ( .A(n23259), .B(n23260), .Z(n352) );
  AND U22986 ( .A(n23261), .B(n23262), .Z(n23260) );
  XNOR U22987 ( .A(p_input[5183]), .B(n23259), .Z(n23262) );
  XOR U22988 ( .A(n23259), .B(p_input[5151]), .Z(n23261) );
  XOR U22989 ( .A(n23263), .B(n23264), .Z(n23259) );
  AND U22990 ( .A(n23265), .B(n23266), .Z(n23264) );
  XNOR U22991 ( .A(p_input[5182]), .B(n23263), .Z(n23266) );
  XNOR U22992 ( .A(n23263), .B(n22865), .Z(n23265) );
  IV U22993 ( .A(p_input[5150]), .Z(n22865) );
  XOR U22994 ( .A(n23267), .B(n23268), .Z(n23263) );
  AND U22995 ( .A(n23269), .B(n23270), .Z(n23268) );
  XNOR U22996 ( .A(p_input[5181]), .B(n23267), .Z(n23270) );
  XNOR U22997 ( .A(n23267), .B(n22874), .Z(n23269) );
  IV U22998 ( .A(p_input[5149]), .Z(n22874) );
  XOR U22999 ( .A(n23271), .B(n23272), .Z(n23267) );
  AND U23000 ( .A(n23273), .B(n23274), .Z(n23272) );
  XNOR U23001 ( .A(p_input[5180]), .B(n23271), .Z(n23274) );
  XNOR U23002 ( .A(n23271), .B(n22883), .Z(n23273) );
  IV U23003 ( .A(p_input[5148]), .Z(n22883) );
  XOR U23004 ( .A(n23275), .B(n23276), .Z(n23271) );
  AND U23005 ( .A(n23277), .B(n23278), .Z(n23276) );
  XNOR U23006 ( .A(p_input[5179]), .B(n23275), .Z(n23278) );
  XNOR U23007 ( .A(n23275), .B(n22892), .Z(n23277) );
  IV U23008 ( .A(p_input[5147]), .Z(n22892) );
  XOR U23009 ( .A(n23279), .B(n23280), .Z(n23275) );
  AND U23010 ( .A(n23281), .B(n23282), .Z(n23280) );
  XNOR U23011 ( .A(p_input[5178]), .B(n23279), .Z(n23282) );
  XNOR U23012 ( .A(n23279), .B(n22901), .Z(n23281) );
  IV U23013 ( .A(p_input[5146]), .Z(n22901) );
  XOR U23014 ( .A(n23283), .B(n23284), .Z(n23279) );
  AND U23015 ( .A(n23285), .B(n23286), .Z(n23284) );
  XNOR U23016 ( .A(p_input[5177]), .B(n23283), .Z(n23286) );
  XNOR U23017 ( .A(n23283), .B(n22910), .Z(n23285) );
  IV U23018 ( .A(p_input[5145]), .Z(n22910) );
  XOR U23019 ( .A(n23287), .B(n23288), .Z(n23283) );
  AND U23020 ( .A(n23289), .B(n23290), .Z(n23288) );
  XNOR U23021 ( .A(p_input[5176]), .B(n23287), .Z(n23290) );
  XNOR U23022 ( .A(n23287), .B(n22919), .Z(n23289) );
  IV U23023 ( .A(p_input[5144]), .Z(n22919) );
  XOR U23024 ( .A(n23291), .B(n23292), .Z(n23287) );
  AND U23025 ( .A(n23293), .B(n23294), .Z(n23292) );
  XNOR U23026 ( .A(p_input[5175]), .B(n23291), .Z(n23294) );
  XNOR U23027 ( .A(n23291), .B(n22928), .Z(n23293) );
  IV U23028 ( .A(p_input[5143]), .Z(n22928) );
  XOR U23029 ( .A(n23295), .B(n23296), .Z(n23291) );
  AND U23030 ( .A(n23297), .B(n23298), .Z(n23296) );
  XNOR U23031 ( .A(p_input[5174]), .B(n23295), .Z(n23298) );
  XNOR U23032 ( .A(n23295), .B(n22937), .Z(n23297) );
  IV U23033 ( .A(p_input[5142]), .Z(n22937) );
  XOR U23034 ( .A(n23299), .B(n23300), .Z(n23295) );
  AND U23035 ( .A(n23301), .B(n23302), .Z(n23300) );
  XNOR U23036 ( .A(p_input[5173]), .B(n23299), .Z(n23302) );
  XNOR U23037 ( .A(n23299), .B(n22946), .Z(n23301) );
  IV U23038 ( .A(p_input[5141]), .Z(n22946) );
  XOR U23039 ( .A(n23303), .B(n23304), .Z(n23299) );
  AND U23040 ( .A(n23305), .B(n23306), .Z(n23304) );
  XNOR U23041 ( .A(p_input[5172]), .B(n23303), .Z(n23306) );
  XNOR U23042 ( .A(n23303), .B(n22955), .Z(n23305) );
  IV U23043 ( .A(p_input[5140]), .Z(n22955) );
  XOR U23044 ( .A(n23307), .B(n23308), .Z(n23303) );
  AND U23045 ( .A(n23309), .B(n23310), .Z(n23308) );
  XNOR U23046 ( .A(p_input[5171]), .B(n23307), .Z(n23310) );
  XNOR U23047 ( .A(n23307), .B(n22964), .Z(n23309) );
  IV U23048 ( .A(p_input[5139]), .Z(n22964) );
  XOR U23049 ( .A(n23311), .B(n23312), .Z(n23307) );
  AND U23050 ( .A(n23313), .B(n23314), .Z(n23312) );
  XNOR U23051 ( .A(p_input[5170]), .B(n23311), .Z(n23314) );
  XNOR U23052 ( .A(n23311), .B(n22973), .Z(n23313) );
  IV U23053 ( .A(p_input[5138]), .Z(n22973) );
  XOR U23054 ( .A(n23315), .B(n23316), .Z(n23311) );
  AND U23055 ( .A(n23317), .B(n23318), .Z(n23316) );
  XNOR U23056 ( .A(p_input[5169]), .B(n23315), .Z(n23318) );
  XNOR U23057 ( .A(n23315), .B(n22982), .Z(n23317) );
  IV U23058 ( .A(p_input[5137]), .Z(n22982) );
  XOR U23059 ( .A(n23319), .B(n23320), .Z(n23315) );
  AND U23060 ( .A(n23321), .B(n23322), .Z(n23320) );
  XNOR U23061 ( .A(p_input[5168]), .B(n23319), .Z(n23322) );
  XNOR U23062 ( .A(n23319), .B(n22991), .Z(n23321) );
  IV U23063 ( .A(p_input[5136]), .Z(n22991) );
  XOR U23064 ( .A(n23323), .B(n23324), .Z(n23319) );
  AND U23065 ( .A(n23325), .B(n23326), .Z(n23324) );
  XNOR U23066 ( .A(p_input[5167]), .B(n23323), .Z(n23326) );
  XNOR U23067 ( .A(n23323), .B(n23000), .Z(n23325) );
  IV U23068 ( .A(p_input[5135]), .Z(n23000) );
  XOR U23069 ( .A(n23327), .B(n23328), .Z(n23323) );
  AND U23070 ( .A(n23329), .B(n23330), .Z(n23328) );
  XNOR U23071 ( .A(p_input[5166]), .B(n23327), .Z(n23330) );
  XNOR U23072 ( .A(n23327), .B(n23009), .Z(n23329) );
  IV U23073 ( .A(p_input[5134]), .Z(n23009) );
  XOR U23074 ( .A(n23331), .B(n23332), .Z(n23327) );
  AND U23075 ( .A(n23333), .B(n23334), .Z(n23332) );
  XNOR U23076 ( .A(p_input[5165]), .B(n23331), .Z(n23334) );
  XNOR U23077 ( .A(n23331), .B(n23018), .Z(n23333) );
  IV U23078 ( .A(p_input[5133]), .Z(n23018) );
  XOR U23079 ( .A(n23335), .B(n23336), .Z(n23331) );
  AND U23080 ( .A(n23337), .B(n23338), .Z(n23336) );
  XNOR U23081 ( .A(p_input[5164]), .B(n23335), .Z(n23338) );
  XNOR U23082 ( .A(n23335), .B(n23027), .Z(n23337) );
  IV U23083 ( .A(p_input[5132]), .Z(n23027) );
  XOR U23084 ( .A(n23339), .B(n23340), .Z(n23335) );
  AND U23085 ( .A(n23341), .B(n23342), .Z(n23340) );
  XNOR U23086 ( .A(p_input[5163]), .B(n23339), .Z(n23342) );
  XNOR U23087 ( .A(n23339), .B(n23036), .Z(n23341) );
  IV U23088 ( .A(p_input[5131]), .Z(n23036) );
  XOR U23089 ( .A(n23343), .B(n23344), .Z(n23339) );
  AND U23090 ( .A(n23345), .B(n23346), .Z(n23344) );
  XNOR U23091 ( .A(p_input[5162]), .B(n23343), .Z(n23346) );
  XNOR U23092 ( .A(n23343), .B(n23045), .Z(n23345) );
  IV U23093 ( .A(p_input[5130]), .Z(n23045) );
  XOR U23094 ( .A(n23347), .B(n23348), .Z(n23343) );
  AND U23095 ( .A(n23349), .B(n23350), .Z(n23348) );
  XNOR U23096 ( .A(p_input[5161]), .B(n23347), .Z(n23350) );
  XNOR U23097 ( .A(n23347), .B(n23054), .Z(n23349) );
  IV U23098 ( .A(p_input[5129]), .Z(n23054) );
  XOR U23099 ( .A(n23351), .B(n23352), .Z(n23347) );
  AND U23100 ( .A(n23353), .B(n23354), .Z(n23352) );
  XNOR U23101 ( .A(p_input[5160]), .B(n23351), .Z(n23354) );
  XNOR U23102 ( .A(n23351), .B(n23063), .Z(n23353) );
  IV U23103 ( .A(p_input[5128]), .Z(n23063) );
  XOR U23104 ( .A(n23355), .B(n23356), .Z(n23351) );
  AND U23105 ( .A(n23357), .B(n23358), .Z(n23356) );
  XNOR U23106 ( .A(p_input[5159]), .B(n23355), .Z(n23358) );
  XNOR U23107 ( .A(n23355), .B(n23072), .Z(n23357) );
  IV U23108 ( .A(p_input[5127]), .Z(n23072) );
  XOR U23109 ( .A(n23359), .B(n23360), .Z(n23355) );
  AND U23110 ( .A(n23361), .B(n23362), .Z(n23360) );
  XNOR U23111 ( .A(p_input[5158]), .B(n23359), .Z(n23362) );
  XNOR U23112 ( .A(n23359), .B(n23081), .Z(n23361) );
  IV U23113 ( .A(p_input[5126]), .Z(n23081) );
  XOR U23114 ( .A(n23363), .B(n23364), .Z(n23359) );
  AND U23115 ( .A(n23365), .B(n23366), .Z(n23364) );
  XNOR U23116 ( .A(p_input[5157]), .B(n23363), .Z(n23366) );
  XNOR U23117 ( .A(n23363), .B(n23090), .Z(n23365) );
  IV U23118 ( .A(p_input[5125]), .Z(n23090) );
  XOR U23119 ( .A(n23367), .B(n23368), .Z(n23363) );
  AND U23120 ( .A(n23369), .B(n23370), .Z(n23368) );
  XNOR U23121 ( .A(p_input[5156]), .B(n23367), .Z(n23370) );
  XNOR U23122 ( .A(n23367), .B(n23099), .Z(n23369) );
  IV U23123 ( .A(p_input[5124]), .Z(n23099) );
  XOR U23124 ( .A(n23371), .B(n23372), .Z(n23367) );
  AND U23125 ( .A(n23373), .B(n23374), .Z(n23372) );
  XNOR U23126 ( .A(p_input[5155]), .B(n23371), .Z(n23374) );
  XNOR U23127 ( .A(n23371), .B(n23108), .Z(n23373) );
  IV U23128 ( .A(p_input[5123]), .Z(n23108) );
  XOR U23129 ( .A(n23375), .B(n23376), .Z(n23371) );
  AND U23130 ( .A(n23377), .B(n23378), .Z(n23376) );
  XNOR U23131 ( .A(p_input[5154]), .B(n23375), .Z(n23378) );
  XNOR U23132 ( .A(n23375), .B(n23117), .Z(n23377) );
  IV U23133 ( .A(p_input[5122]), .Z(n23117) );
  XNOR U23134 ( .A(n23379), .B(n23380), .Z(n23375) );
  AND U23135 ( .A(n23381), .B(n23382), .Z(n23380) );
  XOR U23136 ( .A(p_input[5153]), .B(n23379), .Z(n23382) );
  XNOR U23137 ( .A(p_input[5121]), .B(n23379), .Z(n23381) );
  AND U23138 ( .A(p_input[5152]), .B(n23383), .Z(n23379) );
  IV U23139 ( .A(p_input[5120]), .Z(n23383) );
  XOR U23140 ( .A(n23384), .B(n23385), .Z(n16096) );
  AND U23141 ( .A(n1088), .B(n23386), .Z(n23385) );
  XNOR U23142 ( .A(n23387), .B(n23384), .Z(n23386) );
  XOR U23143 ( .A(n23388), .B(n23389), .Z(n1088) );
  AND U23144 ( .A(n23390), .B(n23391), .Z(n23389) );
  XOR U23145 ( .A(n23388), .B(n16111), .Z(n23391) );
  XOR U23146 ( .A(n23392), .B(n23393), .Z(n16111) );
  AND U23147 ( .A(n1015), .B(n23394), .Z(n23393) );
  XOR U23148 ( .A(n23395), .B(n23392), .Z(n23394) );
  XNOR U23149 ( .A(n16108), .B(n23388), .Z(n23390) );
  XOR U23150 ( .A(n23396), .B(n23397), .Z(n16108) );
  AND U23151 ( .A(n1012), .B(n23398), .Z(n23397) );
  XOR U23152 ( .A(n23399), .B(n23396), .Z(n23398) );
  XOR U23153 ( .A(n23400), .B(n23401), .Z(n23388) );
  AND U23154 ( .A(n23402), .B(n23403), .Z(n23401) );
  XOR U23155 ( .A(n23400), .B(n16123), .Z(n23403) );
  XOR U23156 ( .A(n23404), .B(n23405), .Z(n16123) );
  AND U23157 ( .A(n1015), .B(n23406), .Z(n23405) );
  XOR U23158 ( .A(n23407), .B(n23404), .Z(n23406) );
  XNOR U23159 ( .A(n16120), .B(n23400), .Z(n23402) );
  XOR U23160 ( .A(n23408), .B(n23409), .Z(n16120) );
  AND U23161 ( .A(n1012), .B(n23410), .Z(n23409) );
  XOR U23162 ( .A(n23411), .B(n23408), .Z(n23410) );
  XOR U23163 ( .A(n23412), .B(n23413), .Z(n23400) );
  AND U23164 ( .A(n23414), .B(n23415), .Z(n23413) );
  XOR U23165 ( .A(n23412), .B(n16135), .Z(n23415) );
  XOR U23166 ( .A(n23416), .B(n23417), .Z(n16135) );
  AND U23167 ( .A(n1015), .B(n23418), .Z(n23417) );
  XOR U23168 ( .A(n23419), .B(n23416), .Z(n23418) );
  XNOR U23169 ( .A(n16132), .B(n23412), .Z(n23414) );
  XOR U23170 ( .A(n23420), .B(n23421), .Z(n16132) );
  AND U23171 ( .A(n1012), .B(n23422), .Z(n23421) );
  XOR U23172 ( .A(n23423), .B(n23420), .Z(n23422) );
  XOR U23173 ( .A(n23424), .B(n23425), .Z(n23412) );
  AND U23174 ( .A(n23426), .B(n23427), .Z(n23425) );
  XOR U23175 ( .A(n23424), .B(n16147), .Z(n23427) );
  XOR U23176 ( .A(n23428), .B(n23429), .Z(n16147) );
  AND U23177 ( .A(n1015), .B(n23430), .Z(n23429) );
  XOR U23178 ( .A(n23431), .B(n23428), .Z(n23430) );
  XNOR U23179 ( .A(n16144), .B(n23424), .Z(n23426) );
  XOR U23180 ( .A(n23432), .B(n23433), .Z(n16144) );
  AND U23181 ( .A(n1012), .B(n23434), .Z(n23433) );
  XOR U23182 ( .A(n23435), .B(n23432), .Z(n23434) );
  XOR U23183 ( .A(n23436), .B(n23437), .Z(n23424) );
  AND U23184 ( .A(n23438), .B(n23439), .Z(n23437) );
  XOR U23185 ( .A(n23436), .B(n16159), .Z(n23439) );
  XOR U23186 ( .A(n23440), .B(n23441), .Z(n16159) );
  AND U23187 ( .A(n1015), .B(n23442), .Z(n23441) );
  XOR U23188 ( .A(n23443), .B(n23440), .Z(n23442) );
  XNOR U23189 ( .A(n16156), .B(n23436), .Z(n23438) );
  XOR U23190 ( .A(n23444), .B(n23445), .Z(n16156) );
  AND U23191 ( .A(n1012), .B(n23446), .Z(n23445) );
  XOR U23192 ( .A(n23447), .B(n23444), .Z(n23446) );
  XOR U23193 ( .A(n23448), .B(n23449), .Z(n23436) );
  AND U23194 ( .A(n23450), .B(n23451), .Z(n23449) );
  XOR U23195 ( .A(n23448), .B(n16171), .Z(n23451) );
  XOR U23196 ( .A(n23452), .B(n23453), .Z(n16171) );
  AND U23197 ( .A(n1015), .B(n23454), .Z(n23453) );
  XOR U23198 ( .A(n23455), .B(n23452), .Z(n23454) );
  XNOR U23199 ( .A(n16168), .B(n23448), .Z(n23450) );
  XOR U23200 ( .A(n23456), .B(n23457), .Z(n16168) );
  AND U23201 ( .A(n1012), .B(n23458), .Z(n23457) );
  XOR U23202 ( .A(n23459), .B(n23456), .Z(n23458) );
  XOR U23203 ( .A(n23460), .B(n23461), .Z(n23448) );
  AND U23204 ( .A(n23462), .B(n23463), .Z(n23461) );
  XOR U23205 ( .A(n23460), .B(n16183), .Z(n23463) );
  XOR U23206 ( .A(n23464), .B(n23465), .Z(n16183) );
  AND U23207 ( .A(n1015), .B(n23466), .Z(n23465) );
  XOR U23208 ( .A(n23467), .B(n23464), .Z(n23466) );
  XNOR U23209 ( .A(n16180), .B(n23460), .Z(n23462) );
  XOR U23210 ( .A(n23468), .B(n23469), .Z(n16180) );
  AND U23211 ( .A(n1012), .B(n23470), .Z(n23469) );
  XOR U23212 ( .A(n23471), .B(n23468), .Z(n23470) );
  XOR U23213 ( .A(n23472), .B(n23473), .Z(n23460) );
  AND U23214 ( .A(n23474), .B(n23475), .Z(n23473) );
  XOR U23215 ( .A(n23472), .B(n16195), .Z(n23475) );
  XOR U23216 ( .A(n23476), .B(n23477), .Z(n16195) );
  AND U23217 ( .A(n1015), .B(n23478), .Z(n23477) );
  XOR U23218 ( .A(n23479), .B(n23476), .Z(n23478) );
  XNOR U23219 ( .A(n16192), .B(n23472), .Z(n23474) );
  XOR U23220 ( .A(n23480), .B(n23481), .Z(n16192) );
  AND U23221 ( .A(n1012), .B(n23482), .Z(n23481) );
  XOR U23222 ( .A(n23483), .B(n23480), .Z(n23482) );
  XOR U23223 ( .A(n23484), .B(n23485), .Z(n23472) );
  AND U23224 ( .A(n23486), .B(n23487), .Z(n23485) );
  XOR U23225 ( .A(n23484), .B(n16207), .Z(n23487) );
  XOR U23226 ( .A(n23488), .B(n23489), .Z(n16207) );
  AND U23227 ( .A(n1015), .B(n23490), .Z(n23489) );
  XOR U23228 ( .A(n23491), .B(n23488), .Z(n23490) );
  XNOR U23229 ( .A(n16204), .B(n23484), .Z(n23486) );
  XOR U23230 ( .A(n23492), .B(n23493), .Z(n16204) );
  AND U23231 ( .A(n1012), .B(n23494), .Z(n23493) );
  XOR U23232 ( .A(n23495), .B(n23492), .Z(n23494) );
  XOR U23233 ( .A(n23496), .B(n23497), .Z(n23484) );
  AND U23234 ( .A(n23498), .B(n23499), .Z(n23497) );
  XOR U23235 ( .A(n23496), .B(n16219), .Z(n23499) );
  XOR U23236 ( .A(n23500), .B(n23501), .Z(n16219) );
  AND U23237 ( .A(n1015), .B(n23502), .Z(n23501) );
  XOR U23238 ( .A(n23503), .B(n23500), .Z(n23502) );
  XNOR U23239 ( .A(n16216), .B(n23496), .Z(n23498) );
  XOR U23240 ( .A(n23504), .B(n23505), .Z(n16216) );
  AND U23241 ( .A(n1012), .B(n23506), .Z(n23505) );
  XOR U23242 ( .A(n23507), .B(n23504), .Z(n23506) );
  XOR U23243 ( .A(n23508), .B(n23509), .Z(n23496) );
  AND U23244 ( .A(n23510), .B(n23511), .Z(n23509) );
  XOR U23245 ( .A(n23508), .B(n16231), .Z(n23511) );
  XOR U23246 ( .A(n23512), .B(n23513), .Z(n16231) );
  AND U23247 ( .A(n1015), .B(n23514), .Z(n23513) );
  XOR U23248 ( .A(n23515), .B(n23512), .Z(n23514) );
  XNOR U23249 ( .A(n16228), .B(n23508), .Z(n23510) );
  XOR U23250 ( .A(n23516), .B(n23517), .Z(n16228) );
  AND U23251 ( .A(n1012), .B(n23518), .Z(n23517) );
  XOR U23252 ( .A(n23519), .B(n23516), .Z(n23518) );
  XOR U23253 ( .A(n23520), .B(n23521), .Z(n23508) );
  AND U23254 ( .A(n23522), .B(n23523), .Z(n23521) );
  XOR U23255 ( .A(n23520), .B(n16243), .Z(n23523) );
  XOR U23256 ( .A(n23524), .B(n23525), .Z(n16243) );
  AND U23257 ( .A(n1015), .B(n23526), .Z(n23525) );
  XOR U23258 ( .A(n23527), .B(n23524), .Z(n23526) );
  XNOR U23259 ( .A(n16240), .B(n23520), .Z(n23522) );
  XOR U23260 ( .A(n23528), .B(n23529), .Z(n16240) );
  AND U23261 ( .A(n1012), .B(n23530), .Z(n23529) );
  XOR U23262 ( .A(n23531), .B(n23528), .Z(n23530) );
  XOR U23263 ( .A(n23532), .B(n23533), .Z(n23520) );
  AND U23264 ( .A(n23534), .B(n23535), .Z(n23533) );
  XOR U23265 ( .A(n23532), .B(n16255), .Z(n23535) );
  XOR U23266 ( .A(n23536), .B(n23537), .Z(n16255) );
  AND U23267 ( .A(n1015), .B(n23538), .Z(n23537) );
  XOR U23268 ( .A(n23539), .B(n23536), .Z(n23538) );
  XNOR U23269 ( .A(n16252), .B(n23532), .Z(n23534) );
  XOR U23270 ( .A(n23540), .B(n23541), .Z(n16252) );
  AND U23271 ( .A(n1012), .B(n23542), .Z(n23541) );
  XOR U23272 ( .A(n23543), .B(n23540), .Z(n23542) );
  XOR U23273 ( .A(n23544), .B(n23545), .Z(n23532) );
  AND U23274 ( .A(n23546), .B(n23547), .Z(n23545) );
  XOR U23275 ( .A(n23544), .B(n16267), .Z(n23547) );
  XOR U23276 ( .A(n23548), .B(n23549), .Z(n16267) );
  AND U23277 ( .A(n1015), .B(n23550), .Z(n23549) );
  XOR U23278 ( .A(n23551), .B(n23548), .Z(n23550) );
  XNOR U23279 ( .A(n16264), .B(n23544), .Z(n23546) );
  XOR U23280 ( .A(n23552), .B(n23553), .Z(n16264) );
  AND U23281 ( .A(n1012), .B(n23554), .Z(n23553) );
  XOR U23282 ( .A(n23555), .B(n23552), .Z(n23554) );
  XOR U23283 ( .A(n23556), .B(n23557), .Z(n23544) );
  AND U23284 ( .A(n23558), .B(n23559), .Z(n23557) );
  XOR U23285 ( .A(n23556), .B(n16279), .Z(n23559) );
  XOR U23286 ( .A(n23560), .B(n23561), .Z(n16279) );
  AND U23287 ( .A(n1015), .B(n23562), .Z(n23561) );
  XOR U23288 ( .A(n23563), .B(n23560), .Z(n23562) );
  XNOR U23289 ( .A(n16276), .B(n23556), .Z(n23558) );
  XOR U23290 ( .A(n23564), .B(n23565), .Z(n16276) );
  AND U23291 ( .A(n1012), .B(n23566), .Z(n23565) );
  XOR U23292 ( .A(n23567), .B(n23564), .Z(n23566) );
  XOR U23293 ( .A(n23568), .B(n23569), .Z(n23556) );
  AND U23294 ( .A(n23570), .B(n23571), .Z(n23569) );
  XOR U23295 ( .A(n23568), .B(n16291), .Z(n23571) );
  XOR U23296 ( .A(n23572), .B(n23573), .Z(n16291) );
  AND U23297 ( .A(n1015), .B(n23574), .Z(n23573) );
  XOR U23298 ( .A(n23575), .B(n23572), .Z(n23574) );
  XNOR U23299 ( .A(n16288), .B(n23568), .Z(n23570) );
  XOR U23300 ( .A(n23576), .B(n23577), .Z(n16288) );
  AND U23301 ( .A(n1012), .B(n23578), .Z(n23577) );
  XOR U23302 ( .A(n23579), .B(n23576), .Z(n23578) );
  XOR U23303 ( .A(n23580), .B(n23581), .Z(n23568) );
  AND U23304 ( .A(n23582), .B(n23583), .Z(n23581) );
  XOR U23305 ( .A(n23580), .B(n16303), .Z(n23583) );
  XOR U23306 ( .A(n23584), .B(n23585), .Z(n16303) );
  AND U23307 ( .A(n1015), .B(n23586), .Z(n23585) );
  XOR U23308 ( .A(n23587), .B(n23584), .Z(n23586) );
  XNOR U23309 ( .A(n16300), .B(n23580), .Z(n23582) );
  XOR U23310 ( .A(n23588), .B(n23589), .Z(n16300) );
  AND U23311 ( .A(n1012), .B(n23590), .Z(n23589) );
  XOR U23312 ( .A(n23591), .B(n23588), .Z(n23590) );
  XOR U23313 ( .A(n23592), .B(n23593), .Z(n23580) );
  AND U23314 ( .A(n23594), .B(n23595), .Z(n23593) );
  XOR U23315 ( .A(n23592), .B(n16315), .Z(n23595) );
  XOR U23316 ( .A(n23596), .B(n23597), .Z(n16315) );
  AND U23317 ( .A(n1015), .B(n23598), .Z(n23597) );
  XOR U23318 ( .A(n23599), .B(n23596), .Z(n23598) );
  XNOR U23319 ( .A(n16312), .B(n23592), .Z(n23594) );
  XOR U23320 ( .A(n23600), .B(n23601), .Z(n16312) );
  AND U23321 ( .A(n1012), .B(n23602), .Z(n23601) );
  XOR U23322 ( .A(n23603), .B(n23600), .Z(n23602) );
  XOR U23323 ( .A(n23604), .B(n23605), .Z(n23592) );
  AND U23324 ( .A(n23606), .B(n23607), .Z(n23605) );
  XOR U23325 ( .A(n23604), .B(n16327), .Z(n23607) );
  XOR U23326 ( .A(n23608), .B(n23609), .Z(n16327) );
  AND U23327 ( .A(n1015), .B(n23610), .Z(n23609) );
  XOR U23328 ( .A(n23611), .B(n23608), .Z(n23610) );
  XNOR U23329 ( .A(n16324), .B(n23604), .Z(n23606) );
  XOR U23330 ( .A(n23612), .B(n23613), .Z(n16324) );
  AND U23331 ( .A(n1012), .B(n23614), .Z(n23613) );
  XOR U23332 ( .A(n23615), .B(n23612), .Z(n23614) );
  XOR U23333 ( .A(n23616), .B(n23617), .Z(n23604) );
  AND U23334 ( .A(n23618), .B(n23619), .Z(n23617) );
  XOR U23335 ( .A(n23616), .B(n16339), .Z(n23619) );
  XOR U23336 ( .A(n23620), .B(n23621), .Z(n16339) );
  AND U23337 ( .A(n1015), .B(n23622), .Z(n23621) );
  XOR U23338 ( .A(n23623), .B(n23620), .Z(n23622) );
  XNOR U23339 ( .A(n16336), .B(n23616), .Z(n23618) );
  XOR U23340 ( .A(n23624), .B(n23625), .Z(n16336) );
  AND U23341 ( .A(n1012), .B(n23626), .Z(n23625) );
  XOR U23342 ( .A(n23627), .B(n23624), .Z(n23626) );
  XOR U23343 ( .A(n23628), .B(n23629), .Z(n23616) );
  AND U23344 ( .A(n23630), .B(n23631), .Z(n23629) );
  XOR U23345 ( .A(n23628), .B(n16351), .Z(n23631) );
  XOR U23346 ( .A(n23632), .B(n23633), .Z(n16351) );
  AND U23347 ( .A(n1015), .B(n23634), .Z(n23633) );
  XOR U23348 ( .A(n23635), .B(n23632), .Z(n23634) );
  XNOR U23349 ( .A(n16348), .B(n23628), .Z(n23630) );
  XOR U23350 ( .A(n23636), .B(n23637), .Z(n16348) );
  AND U23351 ( .A(n1012), .B(n23638), .Z(n23637) );
  XOR U23352 ( .A(n23639), .B(n23636), .Z(n23638) );
  XOR U23353 ( .A(n23640), .B(n23641), .Z(n23628) );
  AND U23354 ( .A(n23642), .B(n23643), .Z(n23641) );
  XOR U23355 ( .A(n23640), .B(n16363), .Z(n23643) );
  XOR U23356 ( .A(n23644), .B(n23645), .Z(n16363) );
  AND U23357 ( .A(n1015), .B(n23646), .Z(n23645) );
  XOR U23358 ( .A(n23647), .B(n23644), .Z(n23646) );
  XNOR U23359 ( .A(n16360), .B(n23640), .Z(n23642) );
  XOR U23360 ( .A(n23648), .B(n23649), .Z(n16360) );
  AND U23361 ( .A(n1012), .B(n23650), .Z(n23649) );
  XOR U23362 ( .A(n23651), .B(n23648), .Z(n23650) );
  XOR U23363 ( .A(n23652), .B(n23653), .Z(n23640) );
  AND U23364 ( .A(n23654), .B(n23655), .Z(n23653) );
  XOR U23365 ( .A(n23652), .B(n16375), .Z(n23655) );
  XOR U23366 ( .A(n23656), .B(n23657), .Z(n16375) );
  AND U23367 ( .A(n1015), .B(n23658), .Z(n23657) );
  XOR U23368 ( .A(n23659), .B(n23656), .Z(n23658) );
  XNOR U23369 ( .A(n16372), .B(n23652), .Z(n23654) );
  XOR U23370 ( .A(n23660), .B(n23661), .Z(n16372) );
  AND U23371 ( .A(n1012), .B(n23662), .Z(n23661) );
  XOR U23372 ( .A(n23663), .B(n23660), .Z(n23662) );
  XOR U23373 ( .A(n23664), .B(n23665), .Z(n23652) );
  AND U23374 ( .A(n23666), .B(n23667), .Z(n23665) );
  XOR U23375 ( .A(n23664), .B(n16387), .Z(n23667) );
  XOR U23376 ( .A(n23668), .B(n23669), .Z(n16387) );
  AND U23377 ( .A(n1015), .B(n23670), .Z(n23669) );
  XOR U23378 ( .A(n23671), .B(n23668), .Z(n23670) );
  XNOR U23379 ( .A(n16384), .B(n23664), .Z(n23666) );
  XOR U23380 ( .A(n23672), .B(n23673), .Z(n16384) );
  AND U23381 ( .A(n1012), .B(n23674), .Z(n23673) );
  XOR U23382 ( .A(n23675), .B(n23672), .Z(n23674) );
  XOR U23383 ( .A(n23676), .B(n23677), .Z(n23664) );
  AND U23384 ( .A(n23678), .B(n23679), .Z(n23677) );
  XOR U23385 ( .A(n23676), .B(n16399), .Z(n23679) );
  XOR U23386 ( .A(n23680), .B(n23681), .Z(n16399) );
  AND U23387 ( .A(n1015), .B(n23682), .Z(n23681) );
  XOR U23388 ( .A(n23683), .B(n23680), .Z(n23682) );
  XNOR U23389 ( .A(n16396), .B(n23676), .Z(n23678) );
  XOR U23390 ( .A(n23684), .B(n23685), .Z(n16396) );
  AND U23391 ( .A(n1012), .B(n23686), .Z(n23685) );
  XOR U23392 ( .A(n23687), .B(n23684), .Z(n23686) );
  XOR U23393 ( .A(n23688), .B(n23689), .Z(n23676) );
  AND U23394 ( .A(n23690), .B(n23691), .Z(n23689) );
  XOR U23395 ( .A(n23688), .B(n16411), .Z(n23691) );
  XOR U23396 ( .A(n23692), .B(n23693), .Z(n16411) );
  AND U23397 ( .A(n1015), .B(n23694), .Z(n23693) );
  XOR U23398 ( .A(n23695), .B(n23692), .Z(n23694) );
  XNOR U23399 ( .A(n16408), .B(n23688), .Z(n23690) );
  XOR U23400 ( .A(n23696), .B(n23697), .Z(n16408) );
  AND U23401 ( .A(n1012), .B(n23698), .Z(n23697) );
  XOR U23402 ( .A(n23699), .B(n23696), .Z(n23698) );
  XOR U23403 ( .A(n23700), .B(n23701), .Z(n23688) );
  AND U23404 ( .A(n23702), .B(n23703), .Z(n23701) );
  XOR U23405 ( .A(n23700), .B(n16423), .Z(n23703) );
  XOR U23406 ( .A(n23704), .B(n23705), .Z(n16423) );
  AND U23407 ( .A(n1015), .B(n23706), .Z(n23705) );
  XOR U23408 ( .A(n23707), .B(n23704), .Z(n23706) );
  XNOR U23409 ( .A(n16420), .B(n23700), .Z(n23702) );
  XOR U23410 ( .A(n23708), .B(n23709), .Z(n16420) );
  AND U23411 ( .A(n1012), .B(n23710), .Z(n23709) );
  XOR U23412 ( .A(n23711), .B(n23708), .Z(n23710) );
  XOR U23413 ( .A(n23712), .B(n23713), .Z(n23700) );
  AND U23414 ( .A(n23714), .B(n23715), .Z(n23713) );
  XOR U23415 ( .A(n23712), .B(n16435), .Z(n23715) );
  XOR U23416 ( .A(n23716), .B(n23717), .Z(n16435) );
  AND U23417 ( .A(n1015), .B(n23718), .Z(n23717) );
  XOR U23418 ( .A(n23719), .B(n23716), .Z(n23718) );
  XNOR U23419 ( .A(n16432), .B(n23712), .Z(n23714) );
  XOR U23420 ( .A(n23720), .B(n23721), .Z(n16432) );
  AND U23421 ( .A(n1012), .B(n23722), .Z(n23721) );
  XOR U23422 ( .A(n23723), .B(n23720), .Z(n23722) );
  XOR U23423 ( .A(n23724), .B(n23725), .Z(n23712) );
  AND U23424 ( .A(n23726), .B(n23727), .Z(n23725) );
  XOR U23425 ( .A(n23724), .B(n16447), .Z(n23727) );
  XOR U23426 ( .A(n23728), .B(n23729), .Z(n16447) );
  AND U23427 ( .A(n1015), .B(n23730), .Z(n23729) );
  XOR U23428 ( .A(n23731), .B(n23728), .Z(n23730) );
  XNOR U23429 ( .A(n16444), .B(n23724), .Z(n23726) );
  XOR U23430 ( .A(n23732), .B(n23733), .Z(n16444) );
  AND U23431 ( .A(n1012), .B(n23734), .Z(n23733) );
  XOR U23432 ( .A(n23735), .B(n23732), .Z(n23734) );
  XOR U23433 ( .A(n23736), .B(n23737), .Z(n23724) );
  AND U23434 ( .A(n23738), .B(n23739), .Z(n23737) );
  XOR U23435 ( .A(n23736), .B(n16459), .Z(n23739) );
  XOR U23436 ( .A(n23740), .B(n23741), .Z(n16459) );
  AND U23437 ( .A(n1015), .B(n23742), .Z(n23741) );
  XOR U23438 ( .A(n23743), .B(n23740), .Z(n23742) );
  XNOR U23439 ( .A(n16456), .B(n23736), .Z(n23738) );
  XOR U23440 ( .A(n23744), .B(n23745), .Z(n16456) );
  AND U23441 ( .A(n1012), .B(n23746), .Z(n23745) );
  XOR U23442 ( .A(n23747), .B(n23744), .Z(n23746) );
  XOR U23443 ( .A(n23748), .B(n23749), .Z(n23736) );
  AND U23444 ( .A(n23750), .B(n23751), .Z(n23749) );
  XNOR U23445 ( .A(n23752), .B(n16472), .Z(n23751) );
  XOR U23446 ( .A(n23753), .B(n23754), .Z(n16472) );
  AND U23447 ( .A(n1015), .B(n23755), .Z(n23754) );
  XOR U23448 ( .A(n23753), .B(n23756), .Z(n23755) );
  XNOR U23449 ( .A(n16469), .B(n23748), .Z(n23750) );
  XOR U23450 ( .A(n23757), .B(n23758), .Z(n16469) );
  AND U23451 ( .A(n1012), .B(n23759), .Z(n23758) );
  XOR U23452 ( .A(n23757), .B(n23760), .Z(n23759) );
  IV U23453 ( .A(n23752), .Z(n23748) );
  AND U23454 ( .A(n23384), .B(n23387), .Z(n23752) );
  XNOR U23455 ( .A(n23761), .B(n23762), .Z(n23387) );
  AND U23456 ( .A(n1015), .B(n23763), .Z(n23762) );
  XNOR U23457 ( .A(n23764), .B(n23761), .Z(n23763) );
  XOR U23458 ( .A(n23765), .B(n23766), .Z(n1015) );
  AND U23459 ( .A(n23767), .B(n23768), .Z(n23766) );
  XOR U23460 ( .A(n23765), .B(n23395), .Z(n23768) );
  XOR U23461 ( .A(n23769), .B(n23770), .Z(n23395) );
  AND U23462 ( .A(n855), .B(n23771), .Z(n23770) );
  XOR U23463 ( .A(n23772), .B(n23769), .Z(n23771) );
  XNOR U23464 ( .A(n23392), .B(n23765), .Z(n23767) );
  XOR U23465 ( .A(n23773), .B(n23774), .Z(n23392) );
  AND U23466 ( .A(n853), .B(n23775), .Z(n23774) );
  XOR U23467 ( .A(n23776), .B(n23773), .Z(n23775) );
  XOR U23468 ( .A(n23777), .B(n23778), .Z(n23765) );
  AND U23469 ( .A(n23779), .B(n23780), .Z(n23778) );
  XOR U23470 ( .A(n23777), .B(n23407), .Z(n23780) );
  XOR U23471 ( .A(n23781), .B(n23782), .Z(n23407) );
  AND U23472 ( .A(n855), .B(n23783), .Z(n23782) );
  XOR U23473 ( .A(n23784), .B(n23781), .Z(n23783) );
  XNOR U23474 ( .A(n23404), .B(n23777), .Z(n23779) );
  XOR U23475 ( .A(n23785), .B(n23786), .Z(n23404) );
  AND U23476 ( .A(n853), .B(n23787), .Z(n23786) );
  XOR U23477 ( .A(n23788), .B(n23785), .Z(n23787) );
  XOR U23478 ( .A(n23789), .B(n23790), .Z(n23777) );
  AND U23479 ( .A(n23791), .B(n23792), .Z(n23790) );
  XOR U23480 ( .A(n23789), .B(n23419), .Z(n23792) );
  XOR U23481 ( .A(n23793), .B(n23794), .Z(n23419) );
  AND U23482 ( .A(n855), .B(n23795), .Z(n23794) );
  XOR U23483 ( .A(n23796), .B(n23793), .Z(n23795) );
  XNOR U23484 ( .A(n23416), .B(n23789), .Z(n23791) );
  XOR U23485 ( .A(n23797), .B(n23798), .Z(n23416) );
  AND U23486 ( .A(n853), .B(n23799), .Z(n23798) );
  XOR U23487 ( .A(n23800), .B(n23797), .Z(n23799) );
  XOR U23488 ( .A(n23801), .B(n23802), .Z(n23789) );
  AND U23489 ( .A(n23803), .B(n23804), .Z(n23802) );
  XOR U23490 ( .A(n23801), .B(n23431), .Z(n23804) );
  XOR U23491 ( .A(n23805), .B(n23806), .Z(n23431) );
  AND U23492 ( .A(n855), .B(n23807), .Z(n23806) );
  XOR U23493 ( .A(n23808), .B(n23805), .Z(n23807) );
  XNOR U23494 ( .A(n23428), .B(n23801), .Z(n23803) );
  XOR U23495 ( .A(n23809), .B(n23810), .Z(n23428) );
  AND U23496 ( .A(n853), .B(n23811), .Z(n23810) );
  XOR U23497 ( .A(n23812), .B(n23809), .Z(n23811) );
  XOR U23498 ( .A(n23813), .B(n23814), .Z(n23801) );
  AND U23499 ( .A(n23815), .B(n23816), .Z(n23814) );
  XOR U23500 ( .A(n23813), .B(n23443), .Z(n23816) );
  XOR U23501 ( .A(n23817), .B(n23818), .Z(n23443) );
  AND U23502 ( .A(n855), .B(n23819), .Z(n23818) );
  XOR U23503 ( .A(n23820), .B(n23817), .Z(n23819) );
  XNOR U23504 ( .A(n23440), .B(n23813), .Z(n23815) );
  XOR U23505 ( .A(n23821), .B(n23822), .Z(n23440) );
  AND U23506 ( .A(n853), .B(n23823), .Z(n23822) );
  XOR U23507 ( .A(n23824), .B(n23821), .Z(n23823) );
  XOR U23508 ( .A(n23825), .B(n23826), .Z(n23813) );
  AND U23509 ( .A(n23827), .B(n23828), .Z(n23826) );
  XOR U23510 ( .A(n23825), .B(n23455), .Z(n23828) );
  XOR U23511 ( .A(n23829), .B(n23830), .Z(n23455) );
  AND U23512 ( .A(n855), .B(n23831), .Z(n23830) );
  XOR U23513 ( .A(n23832), .B(n23829), .Z(n23831) );
  XNOR U23514 ( .A(n23452), .B(n23825), .Z(n23827) );
  XOR U23515 ( .A(n23833), .B(n23834), .Z(n23452) );
  AND U23516 ( .A(n853), .B(n23835), .Z(n23834) );
  XOR U23517 ( .A(n23836), .B(n23833), .Z(n23835) );
  XOR U23518 ( .A(n23837), .B(n23838), .Z(n23825) );
  AND U23519 ( .A(n23839), .B(n23840), .Z(n23838) );
  XOR U23520 ( .A(n23837), .B(n23467), .Z(n23840) );
  XOR U23521 ( .A(n23841), .B(n23842), .Z(n23467) );
  AND U23522 ( .A(n855), .B(n23843), .Z(n23842) );
  XOR U23523 ( .A(n23844), .B(n23841), .Z(n23843) );
  XNOR U23524 ( .A(n23464), .B(n23837), .Z(n23839) );
  XOR U23525 ( .A(n23845), .B(n23846), .Z(n23464) );
  AND U23526 ( .A(n853), .B(n23847), .Z(n23846) );
  XOR U23527 ( .A(n23848), .B(n23845), .Z(n23847) );
  XOR U23528 ( .A(n23849), .B(n23850), .Z(n23837) );
  AND U23529 ( .A(n23851), .B(n23852), .Z(n23850) );
  XOR U23530 ( .A(n23849), .B(n23479), .Z(n23852) );
  XOR U23531 ( .A(n23853), .B(n23854), .Z(n23479) );
  AND U23532 ( .A(n855), .B(n23855), .Z(n23854) );
  XOR U23533 ( .A(n23856), .B(n23853), .Z(n23855) );
  XNOR U23534 ( .A(n23476), .B(n23849), .Z(n23851) );
  XOR U23535 ( .A(n23857), .B(n23858), .Z(n23476) );
  AND U23536 ( .A(n853), .B(n23859), .Z(n23858) );
  XOR U23537 ( .A(n23860), .B(n23857), .Z(n23859) );
  XOR U23538 ( .A(n23861), .B(n23862), .Z(n23849) );
  AND U23539 ( .A(n23863), .B(n23864), .Z(n23862) );
  XOR U23540 ( .A(n23861), .B(n23491), .Z(n23864) );
  XOR U23541 ( .A(n23865), .B(n23866), .Z(n23491) );
  AND U23542 ( .A(n855), .B(n23867), .Z(n23866) );
  XOR U23543 ( .A(n23868), .B(n23865), .Z(n23867) );
  XNOR U23544 ( .A(n23488), .B(n23861), .Z(n23863) );
  XOR U23545 ( .A(n23869), .B(n23870), .Z(n23488) );
  AND U23546 ( .A(n853), .B(n23871), .Z(n23870) );
  XOR U23547 ( .A(n23872), .B(n23869), .Z(n23871) );
  XOR U23548 ( .A(n23873), .B(n23874), .Z(n23861) );
  AND U23549 ( .A(n23875), .B(n23876), .Z(n23874) );
  XOR U23550 ( .A(n23873), .B(n23503), .Z(n23876) );
  XOR U23551 ( .A(n23877), .B(n23878), .Z(n23503) );
  AND U23552 ( .A(n855), .B(n23879), .Z(n23878) );
  XOR U23553 ( .A(n23880), .B(n23877), .Z(n23879) );
  XNOR U23554 ( .A(n23500), .B(n23873), .Z(n23875) );
  XOR U23555 ( .A(n23881), .B(n23882), .Z(n23500) );
  AND U23556 ( .A(n853), .B(n23883), .Z(n23882) );
  XOR U23557 ( .A(n23884), .B(n23881), .Z(n23883) );
  XOR U23558 ( .A(n23885), .B(n23886), .Z(n23873) );
  AND U23559 ( .A(n23887), .B(n23888), .Z(n23886) );
  XOR U23560 ( .A(n23885), .B(n23515), .Z(n23888) );
  XOR U23561 ( .A(n23889), .B(n23890), .Z(n23515) );
  AND U23562 ( .A(n855), .B(n23891), .Z(n23890) );
  XOR U23563 ( .A(n23892), .B(n23889), .Z(n23891) );
  XNOR U23564 ( .A(n23512), .B(n23885), .Z(n23887) );
  XOR U23565 ( .A(n23893), .B(n23894), .Z(n23512) );
  AND U23566 ( .A(n853), .B(n23895), .Z(n23894) );
  XOR U23567 ( .A(n23896), .B(n23893), .Z(n23895) );
  XOR U23568 ( .A(n23897), .B(n23898), .Z(n23885) );
  AND U23569 ( .A(n23899), .B(n23900), .Z(n23898) );
  XOR U23570 ( .A(n23897), .B(n23527), .Z(n23900) );
  XOR U23571 ( .A(n23901), .B(n23902), .Z(n23527) );
  AND U23572 ( .A(n855), .B(n23903), .Z(n23902) );
  XOR U23573 ( .A(n23904), .B(n23901), .Z(n23903) );
  XNOR U23574 ( .A(n23524), .B(n23897), .Z(n23899) );
  XOR U23575 ( .A(n23905), .B(n23906), .Z(n23524) );
  AND U23576 ( .A(n853), .B(n23907), .Z(n23906) );
  XOR U23577 ( .A(n23908), .B(n23905), .Z(n23907) );
  XOR U23578 ( .A(n23909), .B(n23910), .Z(n23897) );
  AND U23579 ( .A(n23911), .B(n23912), .Z(n23910) );
  XOR U23580 ( .A(n23909), .B(n23539), .Z(n23912) );
  XOR U23581 ( .A(n23913), .B(n23914), .Z(n23539) );
  AND U23582 ( .A(n855), .B(n23915), .Z(n23914) );
  XOR U23583 ( .A(n23916), .B(n23913), .Z(n23915) );
  XNOR U23584 ( .A(n23536), .B(n23909), .Z(n23911) );
  XOR U23585 ( .A(n23917), .B(n23918), .Z(n23536) );
  AND U23586 ( .A(n853), .B(n23919), .Z(n23918) );
  XOR U23587 ( .A(n23920), .B(n23917), .Z(n23919) );
  XOR U23588 ( .A(n23921), .B(n23922), .Z(n23909) );
  AND U23589 ( .A(n23923), .B(n23924), .Z(n23922) );
  XOR U23590 ( .A(n23921), .B(n23551), .Z(n23924) );
  XOR U23591 ( .A(n23925), .B(n23926), .Z(n23551) );
  AND U23592 ( .A(n855), .B(n23927), .Z(n23926) );
  XOR U23593 ( .A(n23928), .B(n23925), .Z(n23927) );
  XNOR U23594 ( .A(n23548), .B(n23921), .Z(n23923) );
  XOR U23595 ( .A(n23929), .B(n23930), .Z(n23548) );
  AND U23596 ( .A(n853), .B(n23931), .Z(n23930) );
  XOR U23597 ( .A(n23932), .B(n23929), .Z(n23931) );
  XOR U23598 ( .A(n23933), .B(n23934), .Z(n23921) );
  AND U23599 ( .A(n23935), .B(n23936), .Z(n23934) );
  XOR U23600 ( .A(n23933), .B(n23563), .Z(n23936) );
  XOR U23601 ( .A(n23937), .B(n23938), .Z(n23563) );
  AND U23602 ( .A(n855), .B(n23939), .Z(n23938) );
  XOR U23603 ( .A(n23940), .B(n23937), .Z(n23939) );
  XNOR U23604 ( .A(n23560), .B(n23933), .Z(n23935) );
  XOR U23605 ( .A(n23941), .B(n23942), .Z(n23560) );
  AND U23606 ( .A(n853), .B(n23943), .Z(n23942) );
  XOR U23607 ( .A(n23944), .B(n23941), .Z(n23943) );
  XOR U23608 ( .A(n23945), .B(n23946), .Z(n23933) );
  AND U23609 ( .A(n23947), .B(n23948), .Z(n23946) );
  XOR U23610 ( .A(n23945), .B(n23575), .Z(n23948) );
  XOR U23611 ( .A(n23949), .B(n23950), .Z(n23575) );
  AND U23612 ( .A(n855), .B(n23951), .Z(n23950) );
  XOR U23613 ( .A(n23952), .B(n23949), .Z(n23951) );
  XNOR U23614 ( .A(n23572), .B(n23945), .Z(n23947) );
  XOR U23615 ( .A(n23953), .B(n23954), .Z(n23572) );
  AND U23616 ( .A(n853), .B(n23955), .Z(n23954) );
  XOR U23617 ( .A(n23956), .B(n23953), .Z(n23955) );
  XOR U23618 ( .A(n23957), .B(n23958), .Z(n23945) );
  AND U23619 ( .A(n23959), .B(n23960), .Z(n23958) );
  XOR U23620 ( .A(n23957), .B(n23587), .Z(n23960) );
  XOR U23621 ( .A(n23961), .B(n23962), .Z(n23587) );
  AND U23622 ( .A(n855), .B(n23963), .Z(n23962) );
  XOR U23623 ( .A(n23964), .B(n23961), .Z(n23963) );
  XNOR U23624 ( .A(n23584), .B(n23957), .Z(n23959) );
  XOR U23625 ( .A(n23965), .B(n23966), .Z(n23584) );
  AND U23626 ( .A(n853), .B(n23967), .Z(n23966) );
  XOR U23627 ( .A(n23968), .B(n23965), .Z(n23967) );
  XOR U23628 ( .A(n23969), .B(n23970), .Z(n23957) );
  AND U23629 ( .A(n23971), .B(n23972), .Z(n23970) );
  XOR U23630 ( .A(n23969), .B(n23599), .Z(n23972) );
  XOR U23631 ( .A(n23973), .B(n23974), .Z(n23599) );
  AND U23632 ( .A(n855), .B(n23975), .Z(n23974) );
  XOR U23633 ( .A(n23976), .B(n23973), .Z(n23975) );
  XNOR U23634 ( .A(n23596), .B(n23969), .Z(n23971) );
  XOR U23635 ( .A(n23977), .B(n23978), .Z(n23596) );
  AND U23636 ( .A(n853), .B(n23979), .Z(n23978) );
  XOR U23637 ( .A(n23980), .B(n23977), .Z(n23979) );
  XOR U23638 ( .A(n23981), .B(n23982), .Z(n23969) );
  AND U23639 ( .A(n23983), .B(n23984), .Z(n23982) );
  XOR U23640 ( .A(n23981), .B(n23611), .Z(n23984) );
  XOR U23641 ( .A(n23985), .B(n23986), .Z(n23611) );
  AND U23642 ( .A(n855), .B(n23987), .Z(n23986) );
  XOR U23643 ( .A(n23988), .B(n23985), .Z(n23987) );
  XNOR U23644 ( .A(n23608), .B(n23981), .Z(n23983) );
  XOR U23645 ( .A(n23989), .B(n23990), .Z(n23608) );
  AND U23646 ( .A(n853), .B(n23991), .Z(n23990) );
  XOR U23647 ( .A(n23992), .B(n23989), .Z(n23991) );
  XOR U23648 ( .A(n23993), .B(n23994), .Z(n23981) );
  AND U23649 ( .A(n23995), .B(n23996), .Z(n23994) );
  XOR U23650 ( .A(n23993), .B(n23623), .Z(n23996) );
  XOR U23651 ( .A(n23997), .B(n23998), .Z(n23623) );
  AND U23652 ( .A(n855), .B(n23999), .Z(n23998) );
  XOR U23653 ( .A(n24000), .B(n23997), .Z(n23999) );
  XNOR U23654 ( .A(n23620), .B(n23993), .Z(n23995) );
  XOR U23655 ( .A(n24001), .B(n24002), .Z(n23620) );
  AND U23656 ( .A(n853), .B(n24003), .Z(n24002) );
  XOR U23657 ( .A(n24004), .B(n24001), .Z(n24003) );
  XOR U23658 ( .A(n24005), .B(n24006), .Z(n23993) );
  AND U23659 ( .A(n24007), .B(n24008), .Z(n24006) );
  XOR U23660 ( .A(n24005), .B(n23635), .Z(n24008) );
  XOR U23661 ( .A(n24009), .B(n24010), .Z(n23635) );
  AND U23662 ( .A(n855), .B(n24011), .Z(n24010) );
  XOR U23663 ( .A(n24012), .B(n24009), .Z(n24011) );
  XNOR U23664 ( .A(n23632), .B(n24005), .Z(n24007) );
  XOR U23665 ( .A(n24013), .B(n24014), .Z(n23632) );
  AND U23666 ( .A(n853), .B(n24015), .Z(n24014) );
  XOR U23667 ( .A(n24016), .B(n24013), .Z(n24015) );
  XOR U23668 ( .A(n24017), .B(n24018), .Z(n24005) );
  AND U23669 ( .A(n24019), .B(n24020), .Z(n24018) );
  XOR U23670 ( .A(n24017), .B(n23647), .Z(n24020) );
  XOR U23671 ( .A(n24021), .B(n24022), .Z(n23647) );
  AND U23672 ( .A(n855), .B(n24023), .Z(n24022) );
  XOR U23673 ( .A(n24024), .B(n24021), .Z(n24023) );
  XNOR U23674 ( .A(n23644), .B(n24017), .Z(n24019) );
  XOR U23675 ( .A(n24025), .B(n24026), .Z(n23644) );
  AND U23676 ( .A(n853), .B(n24027), .Z(n24026) );
  XOR U23677 ( .A(n24028), .B(n24025), .Z(n24027) );
  XOR U23678 ( .A(n24029), .B(n24030), .Z(n24017) );
  AND U23679 ( .A(n24031), .B(n24032), .Z(n24030) );
  XOR U23680 ( .A(n24029), .B(n23659), .Z(n24032) );
  XOR U23681 ( .A(n24033), .B(n24034), .Z(n23659) );
  AND U23682 ( .A(n855), .B(n24035), .Z(n24034) );
  XOR U23683 ( .A(n24036), .B(n24033), .Z(n24035) );
  XNOR U23684 ( .A(n23656), .B(n24029), .Z(n24031) );
  XOR U23685 ( .A(n24037), .B(n24038), .Z(n23656) );
  AND U23686 ( .A(n853), .B(n24039), .Z(n24038) );
  XOR U23687 ( .A(n24040), .B(n24037), .Z(n24039) );
  XOR U23688 ( .A(n24041), .B(n24042), .Z(n24029) );
  AND U23689 ( .A(n24043), .B(n24044), .Z(n24042) );
  XOR U23690 ( .A(n24041), .B(n23671), .Z(n24044) );
  XOR U23691 ( .A(n24045), .B(n24046), .Z(n23671) );
  AND U23692 ( .A(n855), .B(n24047), .Z(n24046) );
  XOR U23693 ( .A(n24048), .B(n24045), .Z(n24047) );
  XNOR U23694 ( .A(n23668), .B(n24041), .Z(n24043) );
  XOR U23695 ( .A(n24049), .B(n24050), .Z(n23668) );
  AND U23696 ( .A(n853), .B(n24051), .Z(n24050) );
  XOR U23697 ( .A(n24052), .B(n24049), .Z(n24051) );
  XOR U23698 ( .A(n24053), .B(n24054), .Z(n24041) );
  AND U23699 ( .A(n24055), .B(n24056), .Z(n24054) );
  XOR U23700 ( .A(n24053), .B(n23683), .Z(n24056) );
  XOR U23701 ( .A(n24057), .B(n24058), .Z(n23683) );
  AND U23702 ( .A(n855), .B(n24059), .Z(n24058) );
  XOR U23703 ( .A(n24060), .B(n24057), .Z(n24059) );
  XNOR U23704 ( .A(n23680), .B(n24053), .Z(n24055) );
  XOR U23705 ( .A(n24061), .B(n24062), .Z(n23680) );
  AND U23706 ( .A(n853), .B(n24063), .Z(n24062) );
  XOR U23707 ( .A(n24064), .B(n24061), .Z(n24063) );
  XOR U23708 ( .A(n24065), .B(n24066), .Z(n24053) );
  AND U23709 ( .A(n24067), .B(n24068), .Z(n24066) );
  XOR U23710 ( .A(n24065), .B(n23695), .Z(n24068) );
  XOR U23711 ( .A(n24069), .B(n24070), .Z(n23695) );
  AND U23712 ( .A(n855), .B(n24071), .Z(n24070) );
  XOR U23713 ( .A(n24072), .B(n24069), .Z(n24071) );
  XNOR U23714 ( .A(n23692), .B(n24065), .Z(n24067) );
  XOR U23715 ( .A(n24073), .B(n24074), .Z(n23692) );
  AND U23716 ( .A(n853), .B(n24075), .Z(n24074) );
  XOR U23717 ( .A(n24076), .B(n24073), .Z(n24075) );
  XOR U23718 ( .A(n24077), .B(n24078), .Z(n24065) );
  AND U23719 ( .A(n24079), .B(n24080), .Z(n24078) );
  XOR U23720 ( .A(n24077), .B(n23707), .Z(n24080) );
  XOR U23721 ( .A(n24081), .B(n24082), .Z(n23707) );
  AND U23722 ( .A(n855), .B(n24083), .Z(n24082) );
  XOR U23723 ( .A(n24084), .B(n24081), .Z(n24083) );
  XNOR U23724 ( .A(n23704), .B(n24077), .Z(n24079) );
  XOR U23725 ( .A(n24085), .B(n24086), .Z(n23704) );
  AND U23726 ( .A(n853), .B(n24087), .Z(n24086) );
  XOR U23727 ( .A(n24088), .B(n24085), .Z(n24087) );
  XOR U23728 ( .A(n24089), .B(n24090), .Z(n24077) );
  AND U23729 ( .A(n24091), .B(n24092), .Z(n24090) );
  XOR U23730 ( .A(n24089), .B(n23719), .Z(n24092) );
  XOR U23731 ( .A(n24093), .B(n24094), .Z(n23719) );
  AND U23732 ( .A(n855), .B(n24095), .Z(n24094) );
  XOR U23733 ( .A(n24096), .B(n24093), .Z(n24095) );
  XNOR U23734 ( .A(n23716), .B(n24089), .Z(n24091) );
  XOR U23735 ( .A(n24097), .B(n24098), .Z(n23716) );
  AND U23736 ( .A(n853), .B(n24099), .Z(n24098) );
  XOR U23737 ( .A(n24100), .B(n24097), .Z(n24099) );
  XOR U23738 ( .A(n24101), .B(n24102), .Z(n24089) );
  AND U23739 ( .A(n24103), .B(n24104), .Z(n24102) );
  XOR U23740 ( .A(n24101), .B(n23731), .Z(n24104) );
  XOR U23741 ( .A(n24105), .B(n24106), .Z(n23731) );
  AND U23742 ( .A(n855), .B(n24107), .Z(n24106) );
  XOR U23743 ( .A(n24108), .B(n24105), .Z(n24107) );
  XNOR U23744 ( .A(n23728), .B(n24101), .Z(n24103) );
  XOR U23745 ( .A(n24109), .B(n24110), .Z(n23728) );
  AND U23746 ( .A(n853), .B(n24111), .Z(n24110) );
  XOR U23747 ( .A(n24112), .B(n24109), .Z(n24111) );
  XOR U23748 ( .A(n24113), .B(n24114), .Z(n24101) );
  AND U23749 ( .A(n24115), .B(n24116), .Z(n24114) );
  XOR U23750 ( .A(n24113), .B(n23743), .Z(n24116) );
  XOR U23751 ( .A(n24117), .B(n24118), .Z(n23743) );
  AND U23752 ( .A(n855), .B(n24119), .Z(n24118) );
  XOR U23753 ( .A(n24120), .B(n24117), .Z(n24119) );
  XNOR U23754 ( .A(n23740), .B(n24113), .Z(n24115) );
  XOR U23755 ( .A(n24121), .B(n24122), .Z(n23740) );
  AND U23756 ( .A(n853), .B(n24123), .Z(n24122) );
  XOR U23757 ( .A(n24124), .B(n24121), .Z(n24123) );
  XOR U23758 ( .A(n24125), .B(n24126), .Z(n24113) );
  AND U23759 ( .A(n24127), .B(n24128), .Z(n24126) );
  XNOR U23760 ( .A(n24129), .B(n23756), .Z(n24128) );
  XOR U23761 ( .A(n24130), .B(n24131), .Z(n23756) );
  AND U23762 ( .A(n855), .B(n24132), .Z(n24131) );
  XOR U23763 ( .A(n24130), .B(n24133), .Z(n24132) );
  XNOR U23764 ( .A(n23753), .B(n24125), .Z(n24127) );
  XOR U23765 ( .A(n24134), .B(n24135), .Z(n23753) );
  AND U23766 ( .A(n853), .B(n24136), .Z(n24135) );
  XOR U23767 ( .A(n24134), .B(n24137), .Z(n24136) );
  IV U23768 ( .A(n24129), .Z(n24125) );
  AND U23769 ( .A(n23761), .B(n23764), .Z(n24129) );
  XNOR U23770 ( .A(n24138), .B(n24139), .Z(n23764) );
  AND U23771 ( .A(n855), .B(n24140), .Z(n24139) );
  XNOR U23772 ( .A(n24141), .B(n24138), .Z(n24140) );
  XOR U23773 ( .A(n24142), .B(n24143), .Z(n855) );
  AND U23774 ( .A(n24144), .B(n24145), .Z(n24143) );
  XOR U23775 ( .A(n24142), .B(n23772), .Z(n24145) );
  XNOR U23776 ( .A(n24146), .B(n24147), .Z(n23772) );
  AND U23777 ( .A(n24148), .B(n527), .Z(n24147) );
  AND U23778 ( .A(n24146), .B(n24149), .Z(n24148) );
  XNOR U23779 ( .A(n23769), .B(n24142), .Z(n24144) );
  XOR U23780 ( .A(n24150), .B(n24151), .Z(n23769) );
  AND U23781 ( .A(n24152), .B(n525), .Z(n24151) );
  NOR U23782 ( .A(n24150), .B(n24153), .Z(n24152) );
  XOR U23783 ( .A(n24154), .B(n24155), .Z(n24142) );
  AND U23784 ( .A(n24156), .B(n24157), .Z(n24155) );
  XOR U23785 ( .A(n24154), .B(n23784), .Z(n24157) );
  XOR U23786 ( .A(n24158), .B(n24159), .Z(n23784) );
  AND U23787 ( .A(n527), .B(n24160), .Z(n24159) );
  XOR U23788 ( .A(n24161), .B(n24158), .Z(n24160) );
  XNOR U23789 ( .A(n23781), .B(n24154), .Z(n24156) );
  XOR U23790 ( .A(n24162), .B(n24163), .Z(n23781) );
  AND U23791 ( .A(n525), .B(n24164), .Z(n24163) );
  XOR U23792 ( .A(n24165), .B(n24162), .Z(n24164) );
  XOR U23793 ( .A(n24166), .B(n24167), .Z(n24154) );
  AND U23794 ( .A(n24168), .B(n24169), .Z(n24167) );
  XOR U23795 ( .A(n24166), .B(n23796), .Z(n24169) );
  XOR U23796 ( .A(n24170), .B(n24171), .Z(n23796) );
  AND U23797 ( .A(n527), .B(n24172), .Z(n24171) );
  XOR U23798 ( .A(n24173), .B(n24170), .Z(n24172) );
  XNOR U23799 ( .A(n23793), .B(n24166), .Z(n24168) );
  XOR U23800 ( .A(n24174), .B(n24175), .Z(n23793) );
  AND U23801 ( .A(n525), .B(n24176), .Z(n24175) );
  XOR U23802 ( .A(n24177), .B(n24174), .Z(n24176) );
  XOR U23803 ( .A(n24178), .B(n24179), .Z(n24166) );
  AND U23804 ( .A(n24180), .B(n24181), .Z(n24179) );
  XOR U23805 ( .A(n24178), .B(n23808), .Z(n24181) );
  XOR U23806 ( .A(n24182), .B(n24183), .Z(n23808) );
  AND U23807 ( .A(n527), .B(n24184), .Z(n24183) );
  XOR U23808 ( .A(n24185), .B(n24182), .Z(n24184) );
  XNOR U23809 ( .A(n23805), .B(n24178), .Z(n24180) );
  XOR U23810 ( .A(n24186), .B(n24187), .Z(n23805) );
  AND U23811 ( .A(n525), .B(n24188), .Z(n24187) );
  XOR U23812 ( .A(n24189), .B(n24186), .Z(n24188) );
  XOR U23813 ( .A(n24190), .B(n24191), .Z(n24178) );
  AND U23814 ( .A(n24192), .B(n24193), .Z(n24191) );
  XOR U23815 ( .A(n24190), .B(n23820), .Z(n24193) );
  XOR U23816 ( .A(n24194), .B(n24195), .Z(n23820) );
  AND U23817 ( .A(n527), .B(n24196), .Z(n24195) );
  XOR U23818 ( .A(n24197), .B(n24194), .Z(n24196) );
  XNOR U23819 ( .A(n23817), .B(n24190), .Z(n24192) );
  XOR U23820 ( .A(n24198), .B(n24199), .Z(n23817) );
  AND U23821 ( .A(n525), .B(n24200), .Z(n24199) );
  XOR U23822 ( .A(n24201), .B(n24198), .Z(n24200) );
  XOR U23823 ( .A(n24202), .B(n24203), .Z(n24190) );
  AND U23824 ( .A(n24204), .B(n24205), .Z(n24203) );
  XOR U23825 ( .A(n24202), .B(n23832), .Z(n24205) );
  XOR U23826 ( .A(n24206), .B(n24207), .Z(n23832) );
  AND U23827 ( .A(n527), .B(n24208), .Z(n24207) );
  XOR U23828 ( .A(n24209), .B(n24206), .Z(n24208) );
  XNOR U23829 ( .A(n23829), .B(n24202), .Z(n24204) );
  XOR U23830 ( .A(n24210), .B(n24211), .Z(n23829) );
  AND U23831 ( .A(n525), .B(n24212), .Z(n24211) );
  XOR U23832 ( .A(n24213), .B(n24210), .Z(n24212) );
  XOR U23833 ( .A(n24214), .B(n24215), .Z(n24202) );
  AND U23834 ( .A(n24216), .B(n24217), .Z(n24215) );
  XOR U23835 ( .A(n24214), .B(n23844), .Z(n24217) );
  XOR U23836 ( .A(n24218), .B(n24219), .Z(n23844) );
  AND U23837 ( .A(n527), .B(n24220), .Z(n24219) );
  XOR U23838 ( .A(n24221), .B(n24218), .Z(n24220) );
  XNOR U23839 ( .A(n23841), .B(n24214), .Z(n24216) );
  XOR U23840 ( .A(n24222), .B(n24223), .Z(n23841) );
  AND U23841 ( .A(n525), .B(n24224), .Z(n24223) );
  XOR U23842 ( .A(n24225), .B(n24222), .Z(n24224) );
  XOR U23843 ( .A(n24226), .B(n24227), .Z(n24214) );
  AND U23844 ( .A(n24228), .B(n24229), .Z(n24227) );
  XOR U23845 ( .A(n24226), .B(n23856), .Z(n24229) );
  XOR U23846 ( .A(n24230), .B(n24231), .Z(n23856) );
  AND U23847 ( .A(n527), .B(n24232), .Z(n24231) );
  XOR U23848 ( .A(n24233), .B(n24230), .Z(n24232) );
  XNOR U23849 ( .A(n23853), .B(n24226), .Z(n24228) );
  XOR U23850 ( .A(n24234), .B(n24235), .Z(n23853) );
  AND U23851 ( .A(n525), .B(n24236), .Z(n24235) );
  XOR U23852 ( .A(n24237), .B(n24234), .Z(n24236) );
  XOR U23853 ( .A(n24238), .B(n24239), .Z(n24226) );
  AND U23854 ( .A(n24240), .B(n24241), .Z(n24239) );
  XOR U23855 ( .A(n24238), .B(n23868), .Z(n24241) );
  XOR U23856 ( .A(n24242), .B(n24243), .Z(n23868) );
  AND U23857 ( .A(n527), .B(n24244), .Z(n24243) );
  XOR U23858 ( .A(n24245), .B(n24242), .Z(n24244) );
  XNOR U23859 ( .A(n23865), .B(n24238), .Z(n24240) );
  XOR U23860 ( .A(n24246), .B(n24247), .Z(n23865) );
  AND U23861 ( .A(n525), .B(n24248), .Z(n24247) );
  XOR U23862 ( .A(n24249), .B(n24246), .Z(n24248) );
  XOR U23863 ( .A(n24250), .B(n24251), .Z(n24238) );
  AND U23864 ( .A(n24252), .B(n24253), .Z(n24251) );
  XOR U23865 ( .A(n24250), .B(n23880), .Z(n24253) );
  XOR U23866 ( .A(n24254), .B(n24255), .Z(n23880) );
  AND U23867 ( .A(n527), .B(n24256), .Z(n24255) );
  XOR U23868 ( .A(n24257), .B(n24254), .Z(n24256) );
  XNOR U23869 ( .A(n23877), .B(n24250), .Z(n24252) );
  XOR U23870 ( .A(n24258), .B(n24259), .Z(n23877) );
  AND U23871 ( .A(n525), .B(n24260), .Z(n24259) );
  XOR U23872 ( .A(n24261), .B(n24258), .Z(n24260) );
  XOR U23873 ( .A(n24262), .B(n24263), .Z(n24250) );
  AND U23874 ( .A(n24264), .B(n24265), .Z(n24263) );
  XOR U23875 ( .A(n24262), .B(n23892), .Z(n24265) );
  XOR U23876 ( .A(n24266), .B(n24267), .Z(n23892) );
  AND U23877 ( .A(n527), .B(n24268), .Z(n24267) );
  XOR U23878 ( .A(n24269), .B(n24266), .Z(n24268) );
  XNOR U23879 ( .A(n23889), .B(n24262), .Z(n24264) );
  XOR U23880 ( .A(n24270), .B(n24271), .Z(n23889) );
  AND U23881 ( .A(n525), .B(n24272), .Z(n24271) );
  XOR U23882 ( .A(n24273), .B(n24270), .Z(n24272) );
  XOR U23883 ( .A(n24274), .B(n24275), .Z(n24262) );
  AND U23884 ( .A(n24276), .B(n24277), .Z(n24275) );
  XOR U23885 ( .A(n24274), .B(n23904), .Z(n24277) );
  XOR U23886 ( .A(n24278), .B(n24279), .Z(n23904) );
  AND U23887 ( .A(n527), .B(n24280), .Z(n24279) );
  XOR U23888 ( .A(n24281), .B(n24278), .Z(n24280) );
  XNOR U23889 ( .A(n23901), .B(n24274), .Z(n24276) );
  XOR U23890 ( .A(n24282), .B(n24283), .Z(n23901) );
  AND U23891 ( .A(n525), .B(n24284), .Z(n24283) );
  XOR U23892 ( .A(n24285), .B(n24282), .Z(n24284) );
  XOR U23893 ( .A(n24286), .B(n24287), .Z(n24274) );
  AND U23894 ( .A(n24288), .B(n24289), .Z(n24287) );
  XOR U23895 ( .A(n24286), .B(n23916), .Z(n24289) );
  XOR U23896 ( .A(n24290), .B(n24291), .Z(n23916) );
  AND U23897 ( .A(n527), .B(n24292), .Z(n24291) );
  XOR U23898 ( .A(n24293), .B(n24290), .Z(n24292) );
  XNOR U23899 ( .A(n23913), .B(n24286), .Z(n24288) );
  XOR U23900 ( .A(n24294), .B(n24295), .Z(n23913) );
  AND U23901 ( .A(n525), .B(n24296), .Z(n24295) );
  XOR U23902 ( .A(n24297), .B(n24294), .Z(n24296) );
  XOR U23903 ( .A(n24298), .B(n24299), .Z(n24286) );
  AND U23904 ( .A(n24300), .B(n24301), .Z(n24299) );
  XOR U23905 ( .A(n24298), .B(n23928), .Z(n24301) );
  XOR U23906 ( .A(n24302), .B(n24303), .Z(n23928) );
  AND U23907 ( .A(n527), .B(n24304), .Z(n24303) );
  XOR U23908 ( .A(n24305), .B(n24302), .Z(n24304) );
  XNOR U23909 ( .A(n23925), .B(n24298), .Z(n24300) );
  XOR U23910 ( .A(n24306), .B(n24307), .Z(n23925) );
  AND U23911 ( .A(n525), .B(n24308), .Z(n24307) );
  XOR U23912 ( .A(n24309), .B(n24306), .Z(n24308) );
  XOR U23913 ( .A(n24310), .B(n24311), .Z(n24298) );
  AND U23914 ( .A(n24312), .B(n24313), .Z(n24311) );
  XOR U23915 ( .A(n24310), .B(n23940), .Z(n24313) );
  XOR U23916 ( .A(n24314), .B(n24315), .Z(n23940) );
  AND U23917 ( .A(n527), .B(n24316), .Z(n24315) );
  XOR U23918 ( .A(n24317), .B(n24314), .Z(n24316) );
  XNOR U23919 ( .A(n23937), .B(n24310), .Z(n24312) );
  XOR U23920 ( .A(n24318), .B(n24319), .Z(n23937) );
  AND U23921 ( .A(n525), .B(n24320), .Z(n24319) );
  XOR U23922 ( .A(n24321), .B(n24318), .Z(n24320) );
  XOR U23923 ( .A(n24322), .B(n24323), .Z(n24310) );
  AND U23924 ( .A(n24324), .B(n24325), .Z(n24323) );
  XOR U23925 ( .A(n24322), .B(n23952), .Z(n24325) );
  XOR U23926 ( .A(n24326), .B(n24327), .Z(n23952) );
  AND U23927 ( .A(n527), .B(n24328), .Z(n24327) );
  XOR U23928 ( .A(n24329), .B(n24326), .Z(n24328) );
  XNOR U23929 ( .A(n23949), .B(n24322), .Z(n24324) );
  XOR U23930 ( .A(n24330), .B(n24331), .Z(n23949) );
  AND U23931 ( .A(n525), .B(n24332), .Z(n24331) );
  XOR U23932 ( .A(n24333), .B(n24330), .Z(n24332) );
  XOR U23933 ( .A(n24334), .B(n24335), .Z(n24322) );
  AND U23934 ( .A(n24336), .B(n24337), .Z(n24335) );
  XOR U23935 ( .A(n24334), .B(n23964), .Z(n24337) );
  XOR U23936 ( .A(n24338), .B(n24339), .Z(n23964) );
  AND U23937 ( .A(n527), .B(n24340), .Z(n24339) );
  XOR U23938 ( .A(n24341), .B(n24338), .Z(n24340) );
  XNOR U23939 ( .A(n23961), .B(n24334), .Z(n24336) );
  XOR U23940 ( .A(n24342), .B(n24343), .Z(n23961) );
  AND U23941 ( .A(n525), .B(n24344), .Z(n24343) );
  XOR U23942 ( .A(n24345), .B(n24342), .Z(n24344) );
  XOR U23943 ( .A(n24346), .B(n24347), .Z(n24334) );
  AND U23944 ( .A(n24348), .B(n24349), .Z(n24347) );
  XOR U23945 ( .A(n24346), .B(n23976), .Z(n24349) );
  XOR U23946 ( .A(n24350), .B(n24351), .Z(n23976) );
  AND U23947 ( .A(n527), .B(n24352), .Z(n24351) );
  XOR U23948 ( .A(n24353), .B(n24350), .Z(n24352) );
  XNOR U23949 ( .A(n23973), .B(n24346), .Z(n24348) );
  XOR U23950 ( .A(n24354), .B(n24355), .Z(n23973) );
  AND U23951 ( .A(n525), .B(n24356), .Z(n24355) );
  XOR U23952 ( .A(n24357), .B(n24354), .Z(n24356) );
  XOR U23953 ( .A(n24358), .B(n24359), .Z(n24346) );
  AND U23954 ( .A(n24360), .B(n24361), .Z(n24359) );
  XOR U23955 ( .A(n24358), .B(n23988), .Z(n24361) );
  XOR U23956 ( .A(n24362), .B(n24363), .Z(n23988) );
  AND U23957 ( .A(n527), .B(n24364), .Z(n24363) );
  XOR U23958 ( .A(n24365), .B(n24362), .Z(n24364) );
  XNOR U23959 ( .A(n23985), .B(n24358), .Z(n24360) );
  XOR U23960 ( .A(n24366), .B(n24367), .Z(n23985) );
  AND U23961 ( .A(n525), .B(n24368), .Z(n24367) );
  XOR U23962 ( .A(n24369), .B(n24366), .Z(n24368) );
  XOR U23963 ( .A(n24370), .B(n24371), .Z(n24358) );
  AND U23964 ( .A(n24372), .B(n24373), .Z(n24371) );
  XOR U23965 ( .A(n24370), .B(n24000), .Z(n24373) );
  XOR U23966 ( .A(n24374), .B(n24375), .Z(n24000) );
  AND U23967 ( .A(n527), .B(n24376), .Z(n24375) );
  XOR U23968 ( .A(n24377), .B(n24374), .Z(n24376) );
  XNOR U23969 ( .A(n23997), .B(n24370), .Z(n24372) );
  XOR U23970 ( .A(n24378), .B(n24379), .Z(n23997) );
  AND U23971 ( .A(n525), .B(n24380), .Z(n24379) );
  XOR U23972 ( .A(n24381), .B(n24378), .Z(n24380) );
  XOR U23973 ( .A(n24382), .B(n24383), .Z(n24370) );
  AND U23974 ( .A(n24384), .B(n24385), .Z(n24383) );
  XOR U23975 ( .A(n24382), .B(n24012), .Z(n24385) );
  XOR U23976 ( .A(n24386), .B(n24387), .Z(n24012) );
  AND U23977 ( .A(n527), .B(n24388), .Z(n24387) );
  XOR U23978 ( .A(n24389), .B(n24386), .Z(n24388) );
  XNOR U23979 ( .A(n24009), .B(n24382), .Z(n24384) );
  XOR U23980 ( .A(n24390), .B(n24391), .Z(n24009) );
  AND U23981 ( .A(n525), .B(n24392), .Z(n24391) );
  XOR U23982 ( .A(n24393), .B(n24390), .Z(n24392) );
  XOR U23983 ( .A(n24394), .B(n24395), .Z(n24382) );
  AND U23984 ( .A(n24396), .B(n24397), .Z(n24395) );
  XOR U23985 ( .A(n24394), .B(n24024), .Z(n24397) );
  XOR U23986 ( .A(n24398), .B(n24399), .Z(n24024) );
  AND U23987 ( .A(n527), .B(n24400), .Z(n24399) );
  XOR U23988 ( .A(n24401), .B(n24398), .Z(n24400) );
  XNOR U23989 ( .A(n24021), .B(n24394), .Z(n24396) );
  XOR U23990 ( .A(n24402), .B(n24403), .Z(n24021) );
  AND U23991 ( .A(n525), .B(n24404), .Z(n24403) );
  XOR U23992 ( .A(n24405), .B(n24402), .Z(n24404) );
  XOR U23993 ( .A(n24406), .B(n24407), .Z(n24394) );
  AND U23994 ( .A(n24408), .B(n24409), .Z(n24407) );
  XOR U23995 ( .A(n24406), .B(n24036), .Z(n24409) );
  XOR U23996 ( .A(n24410), .B(n24411), .Z(n24036) );
  AND U23997 ( .A(n527), .B(n24412), .Z(n24411) );
  XOR U23998 ( .A(n24413), .B(n24410), .Z(n24412) );
  XNOR U23999 ( .A(n24033), .B(n24406), .Z(n24408) );
  XOR U24000 ( .A(n24414), .B(n24415), .Z(n24033) );
  AND U24001 ( .A(n525), .B(n24416), .Z(n24415) );
  XOR U24002 ( .A(n24417), .B(n24414), .Z(n24416) );
  XOR U24003 ( .A(n24418), .B(n24419), .Z(n24406) );
  AND U24004 ( .A(n24420), .B(n24421), .Z(n24419) );
  XOR U24005 ( .A(n24418), .B(n24048), .Z(n24421) );
  XOR U24006 ( .A(n24422), .B(n24423), .Z(n24048) );
  AND U24007 ( .A(n527), .B(n24424), .Z(n24423) );
  XOR U24008 ( .A(n24425), .B(n24422), .Z(n24424) );
  XNOR U24009 ( .A(n24045), .B(n24418), .Z(n24420) );
  XOR U24010 ( .A(n24426), .B(n24427), .Z(n24045) );
  AND U24011 ( .A(n525), .B(n24428), .Z(n24427) );
  XOR U24012 ( .A(n24429), .B(n24426), .Z(n24428) );
  XOR U24013 ( .A(n24430), .B(n24431), .Z(n24418) );
  AND U24014 ( .A(n24432), .B(n24433), .Z(n24431) );
  XOR U24015 ( .A(n24430), .B(n24060), .Z(n24433) );
  XOR U24016 ( .A(n24434), .B(n24435), .Z(n24060) );
  AND U24017 ( .A(n527), .B(n24436), .Z(n24435) );
  XOR U24018 ( .A(n24437), .B(n24434), .Z(n24436) );
  XNOR U24019 ( .A(n24057), .B(n24430), .Z(n24432) );
  XOR U24020 ( .A(n24438), .B(n24439), .Z(n24057) );
  AND U24021 ( .A(n525), .B(n24440), .Z(n24439) );
  XOR U24022 ( .A(n24441), .B(n24438), .Z(n24440) );
  XOR U24023 ( .A(n24442), .B(n24443), .Z(n24430) );
  AND U24024 ( .A(n24444), .B(n24445), .Z(n24443) );
  XOR U24025 ( .A(n24442), .B(n24072), .Z(n24445) );
  XOR U24026 ( .A(n24446), .B(n24447), .Z(n24072) );
  AND U24027 ( .A(n527), .B(n24448), .Z(n24447) );
  XOR U24028 ( .A(n24449), .B(n24446), .Z(n24448) );
  XNOR U24029 ( .A(n24069), .B(n24442), .Z(n24444) );
  XOR U24030 ( .A(n24450), .B(n24451), .Z(n24069) );
  AND U24031 ( .A(n525), .B(n24452), .Z(n24451) );
  XOR U24032 ( .A(n24453), .B(n24450), .Z(n24452) );
  XOR U24033 ( .A(n24454), .B(n24455), .Z(n24442) );
  AND U24034 ( .A(n24456), .B(n24457), .Z(n24455) );
  XOR U24035 ( .A(n24454), .B(n24084), .Z(n24457) );
  XOR U24036 ( .A(n24458), .B(n24459), .Z(n24084) );
  AND U24037 ( .A(n527), .B(n24460), .Z(n24459) );
  XOR U24038 ( .A(n24461), .B(n24458), .Z(n24460) );
  XNOR U24039 ( .A(n24081), .B(n24454), .Z(n24456) );
  XOR U24040 ( .A(n24462), .B(n24463), .Z(n24081) );
  AND U24041 ( .A(n525), .B(n24464), .Z(n24463) );
  XOR U24042 ( .A(n24465), .B(n24462), .Z(n24464) );
  XOR U24043 ( .A(n24466), .B(n24467), .Z(n24454) );
  AND U24044 ( .A(n24468), .B(n24469), .Z(n24467) );
  XOR U24045 ( .A(n24466), .B(n24096), .Z(n24469) );
  XOR U24046 ( .A(n24470), .B(n24471), .Z(n24096) );
  AND U24047 ( .A(n527), .B(n24472), .Z(n24471) );
  XOR U24048 ( .A(n24473), .B(n24470), .Z(n24472) );
  XNOR U24049 ( .A(n24093), .B(n24466), .Z(n24468) );
  XOR U24050 ( .A(n24474), .B(n24475), .Z(n24093) );
  AND U24051 ( .A(n525), .B(n24476), .Z(n24475) );
  XOR U24052 ( .A(n24477), .B(n24474), .Z(n24476) );
  XOR U24053 ( .A(n24478), .B(n24479), .Z(n24466) );
  AND U24054 ( .A(n24480), .B(n24481), .Z(n24479) );
  XOR U24055 ( .A(n24478), .B(n24108), .Z(n24481) );
  XOR U24056 ( .A(n24482), .B(n24483), .Z(n24108) );
  AND U24057 ( .A(n527), .B(n24484), .Z(n24483) );
  XOR U24058 ( .A(n24485), .B(n24482), .Z(n24484) );
  XNOR U24059 ( .A(n24105), .B(n24478), .Z(n24480) );
  XOR U24060 ( .A(n24486), .B(n24487), .Z(n24105) );
  AND U24061 ( .A(n525), .B(n24488), .Z(n24487) );
  XOR U24062 ( .A(n24489), .B(n24486), .Z(n24488) );
  XOR U24063 ( .A(n24490), .B(n24491), .Z(n24478) );
  AND U24064 ( .A(n24492), .B(n24493), .Z(n24491) );
  XOR U24065 ( .A(n24490), .B(n24120), .Z(n24493) );
  XOR U24066 ( .A(n24494), .B(n24495), .Z(n24120) );
  AND U24067 ( .A(n527), .B(n24496), .Z(n24495) );
  XOR U24068 ( .A(n24497), .B(n24494), .Z(n24496) );
  XNOR U24069 ( .A(n24117), .B(n24490), .Z(n24492) );
  XOR U24070 ( .A(n24498), .B(n24499), .Z(n24117) );
  AND U24071 ( .A(n525), .B(n24500), .Z(n24499) );
  XOR U24072 ( .A(n24501), .B(n24498), .Z(n24500) );
  XOR U24073 ( .A(n24502), .B(n24503), .Z(n24490) );
  AND U24074 ( .A(n24504), .B(n24505), .Z(n24503) );
  XNOR U24075 ( .A(n24506), .B(n24133), .Z(n24505) );
  XOR U24076 ( .A(n24507), .B(n24508), .Z(n24133) );
  AND U24077 ( .A(n527), .B(n24509), .Z(n24508) );
  XOR U24078 ( .A(n24507), .B(n24510), .Z(n24509) );
  XNOR U24079 ( .A(n24130), .B(n24502), .Z(n24504) );
  XOR U24080 ( .A(n24511), .B(n24512), .Z(n24130) );
  AND U24081 ( .A(n525), .B(n24513), .Z(n24512) );
  XOR U24082 ( .A(n24511), .B(n24514), .Z(n24513) );
  IV U24083 ( .A(n24506), .Z(n24502) );
  AND U24084 ( .A(n24138), .B(n24141), .Z(n24506) );
  XNOR U24085 ( .A(n24515), .B(n24516), .Z(n24141) );
  AND U24086 ( .A(n527), .B(n24517), .Z(n24516) );
  XNOR U24087 ( .A(n24518), .B(n24515), .Z(n24517) );
  XOR U24088 ( .A(n24519), .B(n24520), .Z(n527) );
  AND U24089 ( .A(n24521), .B(n24522), .Z(n24520) );
  XOR U24090 ( .A(n24149), .B(n24519), .Z(n24522) );
  IV U24091 ( .A(n24523), .Z(n24149) );
  AND U24092 ( .A(p_input[5119]), .B(p_input[5087]), .Z(n24523) );
  XOR U24093 ( .A(n24519), .B(n24146), .Z(n24521) );
  AND U24094 ( .A(p_input[5023]), .B(p_input[5055]), .Z(n24146) );
  XOR U24095 ( .A(n24524), .B(n24525), .Z(n24519) );
  AND U24096 ( .A(n24526), .B(n24527), .Z(n24525) );
  XOR U24097 ( .A(n24524), .B(n24161), .Z(n24527) );
  XNOR U24098 ( .A(p_input[5086]), .B(n24528), .Z(n24161) );
  AND U24099 ( .A(n371), .B(n24529), .Z(n24528) );
  XOR U24100 ( .A(p_input[5118]), .B(p_input[5086]), .Z(n24529) );
  XNOR U24101 ( .A(n24158), .B(n24524), .Z(n24526) );
  XOR U24102 ( .A(n24530), .B(n24531), .Z(n24158) );
  AND U24103 ( .A(n369), .B(n24532), .Z(n24531) );
  XOR U24104 ( .A(p_input[5054]), .B(p_input[5022]), .Z(n24532) );
  XOR U24105 ( .A(n24533), .B(n24534), .Z(n24524) );
  AND U24106 ( .A(n24535), .B(n24536), .Z(n24534) );
  XOR U24107 ( .A(n24533), .B(n24173), .Z(n24536) );
  XNOR U24108 ( .A(p_input[5085]), .B(n24537), .Z(n24173) );
  AND U24109 ( .A(n371), .B(n24538), .Z(n24537) );
  XOR U24110 ( .A(p_input[5117]), .B(p_input[5085]), .Z(n24538) );
  XNOR U24111 ( .A(n24170), .B(n24533), .Z(n24535) );
  XOR U24112 ( .A(n24539), .B(n24540), .Z(n24170) );
  AND U24113 ( .A(n369), .B(n24541), .Z(n24540) );
  XOR U24114 ( .A(p_input[5053]), .B(p_input[5021]), .Z(n24541) );
  XOR U24115 ( .A(n24542), .B(n24543), .Z(n24533) );
  AND U24116 ( .A(n24544), .B(n24545), .Z(n24543) );
  XOR U24117 ( .A(n24542), .B(n24185), .Z(n24545) );
  XNOR U24118 ( .A(p_input[5084]), .B(n24546), .Z(n24185) );
  AND U24119 ( .A(n371), .B(n24547), .Z(n24546) );
  XOR U24120 ( .A(p_input[5116]), .B(p_input[5084]), .Z(n24547) );
  XNOR U24121 ( .A(n24182), .B(n24542), .Z(n24544) );
  XOR U24122 ( .A(n24548), .B(n24549), .Z(n24182) );
  AND U24123 ( .A(n369), .B(n24550), .Z(n24549) );
  XOR U24124 ( .A(p_input[5052]), .B(p_input[5020]), .Z(n24550) );
  XOR U24125 ( .A(n24551), .B(n24552), .Z(n24542) );
  AND U24126 ( .A(n24553), .B(n24554), .Z(n24552) );
  XOR U24127 ( .A(n24551), .B(n24197), .Z(n24554) );
  XNOR U24128 ( .A(p_input[5083]), .B(n24555), .Z(n24197) );
  AND U24129 ( .A(n371), .B(n24556), .Z(n24555) );
  XOR U24130 ( .A(p_input[5115]), .B(p_input[5083]), .Z(n24556) );
  XNOR U24131 ( .A(n24194), .B(n24551), .Z(n24553) );
  XOR U24132 ( .A(n24557), .B(n24558), .Z(n24194) );
  AND U24133 ( .A(n369), .B(n24559), .Z(n24558) );
  XOR U24134 ( .A(p_input[5051]), .B(p_input[5019]), .Z(n24559) );
  XOR U24135 ( .A(n24560), .B(n24561), .Z(n24551) );
  AND U24136 ( .A(n24562), .B(n24563), .Z(n24561) );
  XOR U24137 ( .A(n24560), .B(n24209), .Z(n24563) );
  XNOR U24138 ( .A(p_input[5082]), .B(n24564), .Z(n24209) );
  AND U24139 ( .A(n371), .B(n24565), .Z(n24564) );
  XOR U24140 ( .A(p_input[5114]), .B(p_input[5082]), .Z(n24565) );
  XNOR U24141 ( .A(n24206), .B(n24560), .Z(n24562) );
  XOR U24142 ( .A(n24566), .B(n24567), .Z(n24206) );
  AND U24143 ( .A(n369), .B(n24568), .Z(n24567) );
  XOR U24144 ( .A(p_input[5050]), .B(p_input[5018]), .Z(n24568) );
  XOR U24145 ( .A(n24569), .B(n24570), .Z(n24560) );
  AND U24146 ( .A(n24571), .B(n24572), .Z(n24570) );
  XOR U24147 ( .A(n24569), .B(n24221), .Z(n24572) );
  XNOR U24148 ( .A(p_input[5081]), .B(n24573), .Z(n24221) );
  AND U24149 ( .A(n371), .B(n24574), .Z(n24573) );
  XOR U24150 ( .A(p_input[5113]), .B(p_input[5081]), .Z(n24574) );
  XNOR U24151 ( .A(n24218), .B(n24569), .Z(n24571) );
  XOR U24152 ( .A(n24575), .B(n24576), .Z(n24218) );
  AND U24153 ( .A(n369), .B(n24577), .Z(n24576) );
  XOR U24154 ( .A(p_input[5049]), .B(p_input[5017]), .Z(n24577) );
  XOR U24155 ( .A(n24578), .B(n24579), .Z(n24569) );
  AND U24156 ( .A(n24580), .B(n24581), .Z(n24579) );
  XOR U24157 ( .A(n24578), .B(n24233), .Z(n24581) );
  XNOR U24158 ( .A(p_input[5080]), .B(n24582), .Z(n24233) );
  AND U24159 ( .A(n371), .B(n24583), .Z(n24582) );
  XOR U24160 ( .A(p_input[5112]), .B(p_input[5080]), .Z(n24583) );
  XNOR U24161 ( .A(n24230), .B(n24578), .Z(n24580) );
  XOR U24162 ( .A(n24584), .B(n24585), .Z(n24230) );
  AND U24163 ( .A(n369), .B(n24586), .Z(n24585) );
  XOR U24164 ( .A(p_input[5048]), .B(p_input[5016]), .Z(n24586) );
  XOR U24165 ( .A(n24587), .B(n24588), .Z(n24578) );
  AND U24166 ( .A(n24589), .B(n24590), .Z(n24588) );
  XOR U24167 ( .A(n24587), .B(n24245), .Z(n24590) );
  XNOR U24168 ( .A(p_input[5079]), .B(n24591), .Z(n24245) );
  AND U24169 ( .A(n371), .B(n24592), .Z(n24591) );
  XOR U24170 ( .A(p_input[5111]), .B(p_input[5079]), .Z(n24592) );
  XNOR U24171 ( .A(n24242), .B(n24587), .Z(n24589) );
  XOR U24172 ( .A(n24593), .B(n24594), .Z(n24242) );
  AND U24173 ( .A(n369), .B(n24595), .Z(n24594) );
  XOR U24174 ( .A(p_input[5047]), .B(p_input[5015]), .Z(n24595) );
  XOR U24175 ( .A(n24596), .B(n24597), .Z(n24587) );
  AND U24176 ( .A(n24598), .B(n24599), .Z(n24597) );
  XOR U24177 ( .A(n24596), .B(n24257), .Z(n24599) );
  XNOR U24178 ( .A(p_input[5078]), .B(n24600), .Z(n24257) );
  AND U24179 ( .A(n371), .B(n24601), .Z(n24600) );
  XOR U24180 ( .A(p_input[5110]), .B(p_input[5078]), .Z(n24601) );
  XNOR U24181 ( .A(n24254), .B(n24596), .Z(n24598) );
  XOR U24182 ( .A(n24602), .B(n24603), .Z(n24254) );
  AND U24183 ( .A(n369), .B(n24604), .Z(n24603) );
  XOR U24184 ( .A(p_input[5046]), .B(p_input[5014]), .Z(n24604) );
  XOR U24185 ( .A(n24605), .B(n24606), .Z(n24596) );
  AND U24186 ( .A(n24607), .B(n24608), .Z(n24606) );
  XOR U24187 ( .A(n24605), .B(n24269), .Z(n24608) );
  XNOR U24188 ( .A(p_input[5077]), .B(n24609), .Z(n24269) );
  AND U24189 ( .A(n371), .B(n24610), .Z(n24609) );
  XOR U24190 ( .A(p_input[5109]), .B(p_input[5077]), .Z(n24610) );
  XNOR U24191 ( .A(n24266), .B(n24605), .Z(n24607) );
  XOR U24192 ( .A(n24611), .B(n24612), .Z(n24266) );
  AND U24193 ( .A(n369), .B(n24613), .Z(n24612) );
  XOR U24194 ( .A(p_input[5045]), .B(p_input[5013]), .Z(n24613) );
  XOR U24195 ( .A(n24614), .B(n24615), .Z(n24605) );
  AND U24196 ( .A(n24616), .B(n24617), .Z(n24615) );
  XOR U24197 ( .A(n24614), .B(n24281), .Z(n24617) );
  XNOR U24198 ( .A(p_input[5076]), .B(n24618), .Z(n24281) );
  AND U24199 ( .A(n371), .B(n24619), .Z(n24618) );
  XOR U24200 ( .A(p_input[5108]), .B(p_input[5076]), .Z(n24619) );
  XNOR U24201 ( .A(n24278), .B(n24614), .Z(n24616) );
  XOR U24202 ( .A(n24620), .B(n24621), .Z(n24278) );
  AND U24203 ( .A(n369), .B(n24622), .Z(n24621) );
  XOR U24204 ( .A(p_input[5044]), .B(p_input[5012]), .Z(n24622) );
  XOR U24205 ( .A(n24623), .B(n24624), .Z(n24614) );
  AND U24206 ( .A(n24625), .B(n24626), .Z(n24624) );
  XOR U24207 ( .A(n24623), .B(n24293), .Z(n24626) );
  XNOR U24208 ( .A(p_input[5075]), .B(n24627), .Z(n24293) );
  AND U24209 ( .A(n371), .B(n24628), .Z(n24627) );
  XOR U24210 ( .A(p_input[5107]), .B(p_input[5075]), .Z(n24628) );
  XNOR U24211 ( .A(n24290), .B(n24623), .Z(n24625) );
  XOR U24212 ( .A(n24629), .B(n24630), .Z(n24290) );
  AND U24213 ( .A(n369), .B(n24631), .Z(n24630) );
  XOR U24214 ( .A(p_input[5043]), .B(p_input[5011]), .Z(n24631) );
  XOR U24215 ( .A(n24632), .B(n24633), .Z(n24623) );
  AND U24216 ( .A(n24634), .B(n24635), .Z(n24633) );
  XOR U24217 ( .A(n24632), .B(n24305), .Z(n24635) );
  XNOR U24218 ( .A(p_input[5074]), .B(n24636), .Z(n24305) );
  AND U24219 ( .A(n371), .B(n24637), .Z(n24636) );
  XOR U24220 ( .A(p_input[5106]), .B(p_input[5074]), .Z(n24637) );
  XNOR U24221 ( .A(n24302), .B(n24632), .Z(n24634) );
  XOR U24222 ( .A(n24638), .B(n24639), .Z(n24302) );
  AND U24223 ( .A(n369), .B(n24640), .Z(n24639) );
  XOR U24224 ( .A(p_input[5042]), .B(p_input[5010]), .Z(n24640) );
  XOR U24225 ( .A(n24641), .B(n24642), .Z(n24632) );
  AND U24226 ( .A(n24643), .B(n24644), .Z(n24642) );
  XOR U24227 ( .A(n24641), .B(n24317), .Z(n24644) );
  XNOR U24228 ( .A(p_input[5073]), .B(n24645), .Z(n24317) );
  AND U24229 ( .A(n371), .B(n24646), .Z(n24645) );
  XOR U24230 ( .A(p_input[5105]), .B(p_input[5073]), .Z(n24646) );
  XNOR U24231 ( .A(n24314), .B(n24641), .Z(n24643) );
  XOR U24232 ( .A(n24647), .B(n24648), .Z(n24314) );
  AND U24233 ( .A(n369), .B(n24649), .Z(n24648) );
  XOR U24234 ( .A(p_input[5041]), .B(p_input[5009]), .Z(n24649) );
  XOR U24235 ( .A(n24650), .B(n24651), .Z(n24641) );
  AND U24236 ( .A(n24652), .B(n24653), .Z(n24651) );
  XOR U24237 ( .A(n24650), .B(n24329), .Z(n24653) );
  XNOR U24238 ( .A(p_input[5072]), .B(n24654), .Z(n24329) );
  AND U24239 ( .A(n371), .B(n24655), .Z(n24654) );
  XOR U24240 ( .A(p_input[5104]), .B(p_input[5072]), .Z(n24655) );
  XNOR U24241 ( .A(n24326), .B(n24650), .Z(n24652) );
  XOR U24242 ( .A(n24656), .B(n24657), .Z(n24326) );
  AND U24243 ( .A(n369), .B(n24658), .Z(n24657) );
  XOR U24244 ( .A(p_input[5040]), .B(p_input[5008]), .Z(n24658) );
  XOR U24245 ( .A(n24659), .B(n24660), .Z(n24650) );
  AND U24246 ( .A(n24661), .B(n24662), .Z(n24660) );
  XOR U24247 ( .A(n24659), .B(n24341), .Z(n24662) );
  XNOR U24248 ( .A(p_input[5071]), .B(n24663), .Z(n24341) );
  AND U24249 ( .A(n371), .B(n24664), .Z(n24663) );
  XOR U24250 ( .A(p_input[5103]), .B(p_input[5071]), .Z(n24664) );
  XNOR U24251 ( .A(n24338), .B(n24659), .Z(n24661) );
  XOR U24252 ( .A(n24665), .B(n24666), .Z(n24338) );
  AND U24253 ( .A(n369), .B(n24667), .Z(n24666) );
  XOR U24254 ( .A(p_input[5039]), .B(p_input[5007]), .Z(n24667) );
  XOR U24255 ( .A(n24668), .B(n24669), .Z(n24659) );
  AND U24256 ( .A(n24670), .B(n24671), .Z(n24669) );
  XOR U24257 ( .A(n24668), .B(n24353), .Z(n24671) );
  XNOR U24258 ( .A(p_input[5070]), .B(n24672), .Z(n24353) );
  AND U24259 ( .A(n371), .B(n24673), .Z(n24672) );
  XOR U24260 ( .A(p_input[5102]), .B(p_input[5070]), .Z(n24673) );
  XNOR U24261 ( .A(n24350), .B(n24668), .Z(n24670) );
  XOR U24262 ( .A(n24674), .B(n24675), .Z(n24350) );
  AND U24263 ( .A(n369), .B(n24676), .Z(n24675) );
  XOR U24264 ( .A(p_input[5038]), .B(p_input[5006]), .Z(n24676) );
  XOR U24265 ( .A(n24677), .B(n24678), .Z(n24668) );
  AND U24266 ( .A(n24679), .B(n24680), .Z(n24678) );
  XOR U24267 ( .A(n24677), .B(n24365), .Z(n24680) );
  XNOR U24268 ( .A(p_input[5069]), .B(n24681), .Z(n24365) );
  AND U24269 ( .A(n371), .B(n24682), .Z(n24681) );
  XOR U24270 ( .A(p_input[5101]), .B(p_input[5069]), .Z(n24682) );
  XNOR U24271 ( .A(n24362), .B(n24677), .Z(n24679) );
  XOR U24272 ( .A(n24683), .B(n24684), .Z(n24362) );
  AND U24273 ( .A(n369), .B(n24685), .Z(n24684) );
  XOR U24274 ( .A(p_input[5037]), .B(p_input[5005]), .Z(n24685) );
  XOR U24275 ( .A(n24686), .B(n24687), .Z(n24677) );
  AND U24276 ( .A(n24688), .B(n24689), .Z(n24687) );
  XOR U24277 ( .A(n24686), .B(n24377), .Z(n24689) );
  XNOR U24278 ( .A(p_input[5068]), .B(n24690), .Z(n24377) );
  AND U24279 ( .A(n371), .B(n24691), .Z(n24690) );
  XOR U24280 ( .A(p_input[5100]), .B(p_input[5068]), .Z(n24691) );
  XNOR U24281 ( .A(n24374), .B(n24686), .Z(n24688) );
  XOR U24282 ( .A(n24692), .B(n24693), .Z(n24374) );
  AND U24283 ( .A(n369), .B(n24694), .Z(n24693) );
  XOR U24284 ( .A(p_input[5036]), .B(p_input[5004]), .Z(n24694) );
  XOR U24285 ( .A(n24695), .B(n24696), .Z(n24686) );
  AND U24286 ( .A(n24697), .B(n24698), .Z(n24696) );
  XOR U24287 ( .A(n24695), .B(n24389), .Z(n24698) );
  XNOR U24288 ( .A(p_input[5067]), .B(n24699), .Z(n24389) );
  AND U24289 ( .A(n371), .B(n24700), .Z(n24699) );
  XOR U24290 ( .A(p_input[5099]), .B(p_input[5067]), .Z(n24700) );
  XNOR U24291 ( .A(n24386), .B(n24695), .Z(n24697) );
  XOR U24292 ( .A(n24701), .B(n24702), .Z(n24386) );
  AND U24293 ( .A(n369), .B(n24703), .Z(n24702) );
  XOR U24294 ( .A(p_input[5035]), .B(p_input[5003]), .Z(n24703) );
  XOR U24295 ( .A(n24704), .B(n24705), .Z(n24695) );
  AND U24296 ( .A(n24706), .B(n24707), .Z(n24705) );
  XOR U24297 ( .A(n24704), .B(n24401), .Z(n24707) );
  XNOR U24298 ( .A(p_input[5066]), .B(n24708), .Z(n24401) );
  AND U24299 ( .A(n371), .B(n24709), .Z(n24708) );
  XOR U24300 ( .A(p_input[5098]), .B(p_input[5066]), .Z(n24709) );
  XNOR U24301 ( .A(n24398), .B(n24704), .Z(n24706) );
  XOR U24302 ( .A(n24710), .B(n24711), .Z(n24398) );
  AND U24303 ( .A(n369), .B(n24712), .Z(n24711) );
  XOR U24304 ( .A(p_input[5034]), .B(p_input[5002]), .Z(n24712) );
  XOR U24305 ( .A(n24713), .B(n24714), .Z(n24704) );
  AND U24306 ( .A(n24715), .B(n24716), .Z(n24714) );
  XOR U24307 ( .A(n24713), .B(n24413), .Z(n24716) );
  XNOR U24308 ( .A(p_input[5065]), .B(n24717), .Z(n24413) );
  AND U24309 ( .A(n371), .B(n24718), .Z(n24717) );
  XOR U24310 ( .A(p_input[5097]), .B(p_input[5065]), .Z(n24718) );
  XNOR U24311 ( .A(n24410), .B(n24713), .Z(n24715) );
  XOR U24312 ( .A(n24719), .B(n24720), .Z(n24410) );
  AND U24313 ( .A(n369), .B(n24721), .Z(n24720) );
  XOR U24314 ( .A(p_input[5033]), .B(p_input[5001]), .Z(n24721) );
  XOR U24315 ( .A(n24722), .B(n24723), .Z(n24713) );
  AND U24316 ( .A(n24724), .B(n24725), .Z(n24723) );
  XOR U24317 ( .A(n24722), .B(n24425), .Z(n24725) );
  XNOR U24318 ( .A(p_input[5064]), .B(n24726), .Z(n24425) );
  AND U24319 ( .A(n371), .B(n24727), .Z(n24726) );
  XOR U24320 ( .A(p_input[5096]), .B(p_input[5064]), .Z(n24727) );
  XNOR U24321 ( .A(n24422), .B(n24722), .Z(n24724) );
  XOR U24322 ( .A(n24728), .B(n24729), .Z(n24422) );
  AND U24323 ( .A(n369), .B(n24730), .Z(n24729) );
  XOR U24324 ( .A(p_input[5032]), .B(p_input[5000]), .Z(n24730) );
  XOR U24325 ( .A(n24731), .B(n24732), .Z(n24722) );
  AND U24326 ( .A(n24733), .B(n24734), .Z(n24732) );
  XOR U24327 ( .A(n24731), .B(n24437), .Z(n24734) );
  XNOR U24328 ( .A(p_input[5063]), .B(n24735), .Z(n24437) );
  AND U24329 ( .A(n371), .B(n24736), .Z(n24735) );
  XOR U24330 ( .A(p_input[5095]), .B(p_input[5063]), .Z(n24736) );
  XNOR U24331 ( .A(n24434), .B(n24731), .Z(n24733) );
  XOR U24332 ( .A(n24737), .B(n24738), .Z(n24434) );
  AND U24333 ( .A(n369), .B(n24739), .Z(n24738) );
  XOR U24334 ( .A(p_input[5031]), .B(p_input[4999]), .Z(n24739) );
  XOR U24335 ( .A(n24740), .B(n24741), .Z(n24731) );
  AND U24336 ( .A(n24742), .B(n24743), .Z(n24741) );
  XOR U24337 ( .A(n24740), .B(n24449), .Z(n24743) );
  XNOR U24338 ( .A(p_input[5062]), .B(n24744), .Z(n24449) );
  AND U24339 ( .A(n371), .B(n24745), .Z(n24744) );
  XOR U24340 ( .A(p_input[5094]), .B(p_input[5062]), .Z(n24745) );
  XNOR U24341 ( .A(n24446), .B(n24740), .Z(n24742) );
  XOR U24342 ( .A(n24746), .B(n24747), .Z(n24446) );
  AND U24343 ( .A(n369), .B(n24748), .Z(n24747) );
  XOR U24344 ( .A(p_input[5030]), .B(p_input[4998]), .Z(n24748) );
  XOR U24345 ( .A(n24749), .B(n24750), .Z(n24740) );
  AND U24346 ( .A(n24751), .B(n24752), .Z(n24750) );
  XOR U24347 ( .A(n24749), .B(n24461), .Z(n24752) );
  XNOR U24348 ( .A(p_input[5061]), .B(n24753), .Z(n24461) );
  AND U24349 ( .A(n371), .B(n24754), .Z(n24753) );
  XOR U24350 ( .A(p_input[5093]), .B(p_input[5061]), .Z(n24754) );
  XNOR U24351 ( .A(n24458), .B(n24749), .Z(n24751) );
  XOR U24352 ( .A(n24755), .B(n24756), .Z(n24458) );
  AND U24353 ( .A(n369), .B(n24757), .Z(n24756) );
  XOR U24354 ( .A(p_input[5029]), .B(p_input[4997]), .Z(n24757) );
  XOR U24355 ( .A(n24758), .B(n24759), .Z(n24749) );
  AND U24356 ( .A(n24760), .B(n24761), .Z(n24759) );
  XOR U24357 ( .A(n24758), .B(n24473), .Z(n24761) );
  XNOR U24358 ( .A(p_input[5060]), .B(n24762), .Z(n24473) );
  AND U24359 ( .A(n371), .B(n24763), .Z(n24762) );
  XOR U24360 ( .A(p_input[5092]), .B(p_input[5060]), .Z(n24763) );
  XNOR U24361 ( .A(n24470), .B(n24758), .Z(n24760) );
  XOR U24362 ( .A(n24764), .B(n24765), .Z(n24470) );
  AND U24363 ( .A(n369), .B(n24766), .Z(n24765) );
  XOR U24364 ( .A(p_input[5028]), .B(p_input[4996]), .Z(n24766) );
  XOR U24365 ( .A(n24767), .B(n24768), .Z(n24758) );
  AND U24366 ( .A(n24769), .B(n24770), .Z(n24768) );
  XOR U24367 ( .A(n24767), .B(n24485), .Z(n24770) );
  XNOR U24368 ( .A(p_input[5059]), .B(n24771), .Z(n24485) );
  AND U24369 ( .A(n371), .B(n24772), .Z(n24771) );
  XOR U24370 ( .A(p_input[5091]), .B(p_input[5059]), .Z(n24772) );
  XNOR U24371 ( .A(n24482), .B(n24767), .Z(n24769) );
  XOR U24372 ( .A(n24773), .B(n24774), .Z(n24482) );
  AND U24373 ( .A(n369), .B(n24775), .Z(n24774) );
  XOR U24374 ( .A(p_input[5027]), .B(p_input[4995]), .Z(n24775) );
  XOR U24375 ( .A(n24776), .B(n24777), .Z(n24767) );
  AND U24376 ( .A(n24778), .B(n24779), .Z(n24777) );
  XOR U24377 ( .A(n24776), .B(n24497), .Z(n24779) );
  XNOR U24378 ( .A(p_input[5058]), .B(n24780), .Z(n24497) );
  AND U24379 ( .A(n371), .B(n24781), .Z(n24780) );
  XOR U24380 ( .A(p_input[5090]), .B(p_input[5058]), .Z(n24781) );
  XNOR U24381 ( .A(n24494), .B(n24776), .Z(n24778) );
  XOR U24382 ( .A(n24782), .B(n24783), .Z(n24494) );
  AND U24383 ( .A(n369), .B(n24784), .Z(n24783) );
  XOR U24384 ( .A(p_input[5026]), .B(p_input[4994]), .Z(n24784) );
  XOR U24385 ( .A(n24785), .B(n24786), .Z(n24776) );
  AND U24386 ( .A(n24787), .B(n24788), .Z(n24786) );
  XNOR U24387 ( .A(n24789), .B(n24510), .Z(n24788) );
  XNOR U24388 ( .A(p_input[5057]), .B(n24790), .Z(n24510) );
  AND U24389 ( .A(n371), .B(n24791), .Z(n24790) );
  XNOR U24390 ( .A(p_input[5089]), .B(n24792), .Z(n24791) );
  IV U24391 ( .A(p_input[5057]), .Z(n24792) );
  XNOR U24392 ( .A(n24507), .B(n24785), .Z(n24787) );
  XNOR U24393 ( .A(p_input[4993]), .B(n24793), .Z(n24507) );
  AND U24394 ( .A(n369), .B(n24794), .Z(n24793) );
  XOR U24395 ( .A(p_input[5025]), .B(p_input[4993]), .Z(n24794) );
  IV U24396 ( .A(n24789), .Z(n24785) );
  AND U24397 ( .A(n24515), .B(n24518), .Z(n24789) );
  XOR U24398 ( .A(p_input[5056]), .B(n24795), .Z(n24518) );
  AND U24399 ( .A(n371), .B(n24796), .Z(n24795) );
  XOR U24400 ( .A(p_input[5088]), .B(p_input[5056]), .Z(n24796) );
  XOR U24401 ( .A(n24797), .B(n24798), .Z(n371) );
  AND U24402 ( .A(n24799), .B(n24800), .Z(n24798) );
  XNOR U24403 ( .A(p_input[5119]), .B(n24797), .Z(n24800) );
  XOR U24404 ( .A(n24797), .B(p_input[5087]), .Z(n24799) );
  XOR U24405 ( .A(n24801), .B(n24802), .Z(n24797) );
  AND U24406 ( .A(n24803), .B(n24804), .Z(n24802) );
  XNOR U24407 ( .A(p_input[5118]), .B(n24801), .Z(n24804) );
  XOR U24408 ( .A(n24801), .B(p_input[5086]), .Z(n24803) );
  XOR U24409 ( .A(n24805), .B(n24806), .Z(n24801) );
  AND U24410 ( .A(n24807), .B(n24808), .Z(n24806) );
  XNOR U24411 ( .A(p_input[5117]), .B(n24805), .Z(n24808) );
  XOR U24412 ( .A(n24805), .B(p_input[5085]), .Z(n24807) );
  XOR U24413 ( .A(n24809), .B(n24810), .Z(n24805) );
  AND U24414 ( .A(n24811), .B(n24812), .Z(n24810) );
  XNOR U24415 ( .A(p_input[5116]), .B(n24809), .Z(n24812) );
  XOR U24416 ( .A(n24809), .B(p_input[5084]), .Z(n24811) );
  XOR U24417 ( .A(n24813), .B(n24814), .Z(n24809) );
  AND U24418 ( .A(n24815), .B(n24816), .Z(n24814) );
  XNOR U24419 ( .A(p_input[5115]), .B(n24813), .Z(n24816) );
  XOR U24420 ( .A(n24813), .B(p_input[5083]), .Z(n24815) );
  XOR U24421 ( .A(n24817), .B(n24818), .Z(n24813) );
  AND U24422 ( .A(n24819), .B(n24820), .Z(n24818) );
  XNOR U24423 ( .A(p_input[5114]), .B(n24817), .Z(n24820) );
  XOR U24424 ( .A(n24817), .B(p_input[5082]), .Z(n24819) );
  XOR U24425 ( .A(n24821), .B(n24822), .Z(n24817) );
  AND U24426 ( .A(n24823), .B(n24824), .Z(n24822) );
  XNOR U24427 ( .A(p_input[5113]), .B(n24821), .Z(n24824) );
  XOR U24428 ( .A(n24821), .B(p_input[5081]), .Z(n24823) );
  XOR U24429 ( .A(n24825), .B(n24826), .Z(n24821) );
  AND U24430 ( .A(n24827), .B(n24828), .Z(n24826) );
  XNOR U24431 ( .A(p_input[5112]), .B(n24825), .Z(n24828) );
  XOR U24432 ( .A(n24825), .B(p_input[5080]), .Z(n24827) );
  XOR U24433 ( .A(n24829), .B(n24830), .Z(n24825) );
  AND U24434 ( .A(n24831), .B(n24832), .Z(n24830) );
  XNOR U24435 ( .A(p_input[5111]), .B(n24829), .Z(n24832) );
  XOR U24436 ( .A(n24829), .B(p_input[5079]), .Z(n24831) );
  XOR U24437 ( .A(n24833), .B(n24834), .Z(n24829) );
  AND U24438 ( .A(n24835), .B(n24836), .Z(n24834) );
  XNOR U24439 ( .A(p_input[5110]), .B(n24833), .Z(n24836) );
  XOR U24440 ( .A(n24833), .B(p_input[5078]), .Z(n24835) );
  XOR U24441 ( .A(n24837), .B(n24838), .Z(n24833) );
  AND U24442 ( .A(n24839), .B(n24840), .Z(n24838) );
  XNOR U24443 ( .A(p_input[5109]), .B(n24837), .Z(n24840) );
  XOR U24444 ( .A(n24837), .B(p_input[5077]), .Z(n24839) );
  XOR U24445 ( .A(n24841), .B(n24842), .Z(n24837) );
  AND U24446 ( .A(n24843), .B(n24844), .Z(n24842) );
  XNOR U24447 ( .A(p_input[5108]), .B(n24841), .Z(n24844) );
  XOR U24448 ( .A(n24841), .B(p_input[5076]), .Z(n24843) );
  XOR U24449 ( .A(n24845), .B(n24846), .Z(n24841) );
  AND U24450 ( .A(n24847), .B(n24848), .Z(n24846) );
  XNOR U24451 ( .A(p_input[5107]), .B(n24845), .Z(n24848) );
  XOR U24452 ( .A(n24845), .B(p_input[5075]), .Z(n24847) );
  XOR U24453 ( .A(n24849), .B(n24850), .Z(n24845) );
  AND U24454 ( .A(n24851), .B(n24852), .Z(n24850) );
  XNOR U24455 ( .A(p_input[5106]), .B(n24849), .Z(n24852) );
  XOR U24456 ( .A(n24849), .B(p_input[5074]), .Z(n24851) );
  XOR U24457 ( .A(n24853), .B(n24854), .Z(n24849) );
  AND U24458 ( .A(n24855), .B(n24856), .Z(n24854) );
  XNOR U24459 ( .A(p_input[5105]), .B(n24853), .Z(n24856) );
  XOR U24460 ( .A(n24853), .B(p_input[5073]), .Z(n24855) );
  XOR U24461 ( .A(n24857), .B(n24858), .Z(n24853) );
  AND U24462 ( .A(n24859), .B(n24860), .Z(n24858) );
  XNOR U24463 ( .A(p_input[5104]), .B(n24857), .Z(n24860) );
  XOR U24464 ( .A(n24857), .B(p_input[5072]), .Z(n24859) );
  XOR U24465 ( .A(n24861), .B(n24862), .Z(n24857) );
  AND U24466 ( .A(n24863), .B(n24864), .Z(n24862) );
  XNOR U24467 ( .A(p_input[5103]), .B(n24861), .Z(n24864) );
  XOR U24468 ( .A(n24861), .B(p_input[5071]), .Z(n24863) );
  XOR U24469 ( .A(n24865), .B(n24866), .Z(n24861) );
  AND U24470 ( .A(n24867), .B(n24868), .Z(n24866) );
  XNOR U24471 ( .A(p_input[5102]), .B(n24865), .Z(n24868) );
  XOR U24472 ( .A(n24865), .B(p_input[5070]), .Z(n24867) );
  XOR U24473 ( .A(n24869), .B(n24870), .Z(n24865) );
  AND U24474 ( .A(n24871), .B(n24872), .Z(n24870) );
  XNOR U24475 ( .A(p_input[5101]), .B(n24869), .Z(n24872) );
  XOR U24476 ( .A(n24869), .B(p_input[5069]), .Z(n24871) );
  XOR U24477 ( .A(n24873), .B(n24874), .Z(n24869) );
  AND U24478 ( .A(n24875), .B(n24876), .Z(n24874) );
  XNOR U24479 ( .A(p_input[5100]), .B(n24873), .Z(n24876) );
  XOR U24480 ( .A(n24873), .B(p_input[5068]), .Z(n24875) );
  XOR U24481 ( .A(n24877), .B(n24878), .Z(n24873) );
  AND U24482 ( .A(n24879), .B(n24880), .Z(n24878) );
  XNOR U24483 ( .A(p_input[5099]), .B(n24877), .Z(n24880) );
  XOR U24484 ( .A(n24877), .B(p_input[5067]), .Z(n24879) );
  XOR U24485 ( .A(n24881), .B(n24882), .Z(n24877) );
  AND U24486 ( .A(n24883), .B(n24884), .Z(n24882) );
  XNOR U24487 ( .A(p_input[5098]), .B(n24881), .Z(n24884) );
  XOR U24488 ( .A(n24881), .B(p_input[5066]), .Z(n24883) );
  XOR U24489 ( .A(n24885), .B(n24886), .Z(n24881) );
  AND U24490 ( .A(n24887), .B(n24888), .Z(n24886) );
  XNOR U24491 ( .A(p_input[5097]), .B(n24885), .Z(n24888) );
  XOR U24492 ( .A(n24885), .B(p_input[5065]), .Z(n24887) );
  XOR U24493 ( .A(n24889), .B(n24890), .Z(n24885) );
  AND U24494 ( .A(n24891), .B(n24892), .Z(n24890) );
  XNOR U24495 ( .A(p_input[5096]), .B(n24889), .Z(n24892) );
  XOR U24496 ( .A(n24889), .B(p_input[5064]), .Z(n24891) );
  XOR U24497 ( .A(n24893), .B(n24894), .Z(n24889) );
  AND U24498 ( .A(n24895), .B(n24896), .Z(n24894) );
  XNOR U24499 ( .A(p_input[5095]), .B(n24893), .Z(n24896) );
  XOR U24500 ( .A(n24893), .B(p_input[5063]), .Z(n24895) );
  XOR U24501 ( .A(n24897), .B(n24898), .Z(n24893) );
  AND U24502 ( .A(n24899), .B(n24900), .Z(n24898) );
  XNOR U24503 ( .A(p_input[5094]), .B(n24897), .Z(n24900) );
  XOR U24504 ( .A(n24897), .B(p_input[5062]), .Z(n24899) );
  XOR U24505 ( .A(n24901), .B(n24902), .Z(n24897) );
  AND U24506 ( .A(n24903), .B(n24904), .Z(n24902) );
  XNOR U24507 ( .A(p_input[5093]), .B(n24901), .Z(n24904) );
  XOR U24508 ( .A(n24901), .B(p_input[5061]), .Z(n24903) );
  XOR U24509 ( .A(n24905), .B(n24906), .Z(n24901) );
  AND U24510 ( .A(n24907), .B(n24908), .Z(n24906) );
  XNOR U24511 ( .A(p_input[5092]), .B(n24905), .Z(n24908) );
  XOR U24512 ( .A(n24905), .B(p_input[5060]), .Z(n24907) );
  XOR U24513 ( .A(n24909), .B(n24910), .Z(n24905) );
  AND U24514 ( .A(n24911), .B(n24912), .Z(n24910) );
  XNOR U24515 ( .A(p_input[5091]), .B(n24909), .Z(n24912) );
  XOR U24516 ( .A(n24909), .B(p_input[5059]), .Z(n24911) );
  XOR U24517 ( .A(n24913), .B(n24914), .Z(n24909) );
  AND U24518 ( .A(n24915), .B(n24916), .Z(n24914) );
  XNOR U24519 ( .A(p_input[5090]), .B(n24913), .Z(n24916) );
  XOR U24520 ( .A(n24913), .B(p_input[5058]), .Z(n24915) );
  XNOR U24521 ( .A(n24917), .B(n24918), .Z(n24913) );
  AND U24522 ( .A(n24919), .B(n24920), .Z(n24918) );
  XOR U24523 ( .A(p_input[5089]), .B(n24917), .Z(n24920) );
  XNOR U24524 ( .A(p_input[5057]), .B(n24917), .Z(n24919) );
  AND U24525 ( .A(p_input[5088]), .B(n24921), .Z(n24917) );
  IV U24526 ( .A(p_input[5056]), .Z(n24921) );
  XNOR U24527 ( .A(p_input[4992]), .B(n24922), .Z(n24515) );
  AND U24528 ( .A(n369), .B(n24923), .Z(n24922) );
  XOR U24529 ( .A(p_input[5024]), .B(p_input[4992]), .Z(n24923) );
  XOR U24530 ( .A(n24924), .B(n24925), .Z(n369) );
  AND U24531 ( .A(n24926), .B(n24927), .Z(n24925) );
  XNOR U24532 ( .A(p_input[5055]), .B(n24924), .Z(n24927) );
  XOR U24533 ( .A(n24924), .B(p_input[5023]), .Z(n24926) );
  XOR U24534 ( .A(n24928), .B(n24929), .Z(n24924) );
  AND U24535 ( .A(n24930), .B(n24931), .Z(n24929) );
  XNOR U24536 ( .A(p_input[5054]), .B(n24928), .Z(n24931) );
  XNOR U24537 ( .A(n24928), .B(n24530), .Z(n24930) );
  IV U24538 ( .A(p_input[5022]), .Z(n24530) );
  XOR U24539 ( .A(n24932), .B(n24933), .Z(n24928) );
  AND U24540 ( .A(n24934), .B(n24935), .Z(n24933) );
  XNOR U24541 ( .A(p_input[5053]), .B(n24932), .Z(n24935) );
  XNOR U24542 ( .A(n24932), .B(n24539), .Z(n24934) );
  IV U24543 ( .A(p_input[5021]), .Z(n24539) );
  XOR U24544 ( .A(n24936), .B(n24937), .Z(n24932) );
  AND U24545 ( .A(n24938), .B(n24939), .Z(n24937) );
  XNOR U24546 ( .A(p_input[5052]), .B(n24936), .Z(n24939) );
  XNOR U24547 ( .A(n24936), .B(n24548), .Z(n24938) );
  IV U24548 ( .A(p_input[5020]), .Z(n24548) );
  XOR U24549 ( .A(n24940), .B(n24941), .Z(n24936) );
  AND U24550 ( .A(n24942), .B(n24943), .Z(n24941) );
  XNOR U24551 ( .A(p_input[5051]), .B(n24940), .Z(n24943) );
  XNOR U24552 ( .A(n24940), .B(n24557), .Z(n24942) );
  IV U24553 ( .A(p_input[5019]), .Z(n24557) );
  XOR U24554 ( .A(n24944), .B(n24945), .Z(n24940) );
  AND U24555 ( .A(n24946), .B(n24947), .Z(n24945) );
  XNOR U24556 ( .A(p_input[5050]), .B(n24944), .Z(n24947) );
  XNOR U24557 ( .A(n24944), .B(n24566), .Z(n24946) );
  IV U24558 ( .A(p_input[5018]), .Z(n24566) );
  XOR U24559 ( .A(n24948), .B(n24949), .Z(n24944) );
  AND U24560 ( .A(n24950), .B(n24951), .Z(n24949) );
  XNOR U24561 ( .A(p_input[5049]), .B(n24948), .Z(n24951) );
  XNOR U24562 ( .A(n24948), .B(n24575), .Z(n24950) );
  IV U24563 ( .A(p_input[5017]), .Z(n24575) );
  XOR U24564 ( .A(n24952), .B(n24953), .Z(n24948) );
  AND U24565 ( .A(n24954), .B(n24955), .Z(n24953) );
  XNOR U24566 ( .A(p_input[5048]), .B(n24952), .Z(n24955) );
  XNOR U24567 ( .A(n24952), .B(n24584), .Z(n24954) );
  IV U24568 ( .A(p_input[5016]), .Z(n24584) );
  XOR U24569 ( .A(n24956), .B(n24957), .Z(n24952) );
  AND U24570 ( .A(n24958), .B(n24959), .Z(n24957) );
  XNOR U24571 ( .A(p_input[5047]), .B(n24956), .Z(n24959) );
  XNOR U24572 ( .A(n24956), .B(n24593), .Z(n24958) );
  IV U24573 ( .A(p_input[5015]), .Z(n24593) );
  XOR U24574 ( .A(n24960), .B(n24961), .Z(n24956) );
  AND U24575 ( .A(n24962), .B(n24963), .Z(n24961) );
  XNOR U24576 ( .A(p_input[5046]), .B(n24960), .Z(n24963) );
  XNOR U24577 ( .A(n24960), .B(n24602), .Z(n24962) );
  IV U24578 ( .A(p_input[5014]), .Z(n24602) );
  XOR U24579 ( .A(n24964), .B(n24965), .Z(n24960) );
  AND U24580 ( .A(n24966), .B(n24967), .Z(n24965) );
  XNOR U24581 ( .A(p_input[5045]), .B(n24964), .Z(n24967) );
  XNOR U24582 ( .A(n24964), .B(n24611), .Z(n24966) );
  IV U24583 ( .A(p_input[5013]), .Z(n24611) );
  XOR U24584 ( .A(n24968), .B(n24969), .Z(n24964) );
  AND U24585 ( .A(n24970), .B(n24971), .Z(n24969) );
  XNOR U24586 ( .A(p_input[5044]), .B(n24968), .Z(n24971) );
  XNOR U24587 ( .A(n24968), .B(n24620), .Z(n24970) );
  IV U24588 ( .A(p_input[5012]), .Z(n24620) );
  XOR U24589 ( .A(n24972), .B(n24973), .Z(n24968) );
  AND U24590 ( .A(n24974), .B(n24975), .Z(n24973) );
  XNOR U24591 ( .A(p_input[5043]), .B(n24972), .Z(n24975) );
  XNOR U24592 ( .A(n24972), .B(n24629), .Z(n24974) );
  IV U24593 ( .A(p_input[5011]), .Z(n24629) );
  XOR U24594 ( .A(n24976), .B(n24977), .Z(n24972) );
  AND U24595 ( .A(n24978), .B(n24979), .Z(n24977) );
  XNOR U24596 ( .A(p_input[5042]), .B(n24976), .Z(n24979) );
  XNOR U24597 ( .A(n24976), .B(n24638), .Z(n24978) );
  IV U24598 ( .A(p_input[5010]), .Z(n24638) );
  XOR U24599 ( .A(n24980), .B(n24981), .Z(n24976) );
  AND U24600 ( .A(n24982), .B(n24983), .Z(n24981) );
  XNOR U24601 ( .A(p_input[5041]), .B(n24980), .Z(n24983) );
  XNOR U24602 ( .A(n24980), .B(n24647), .Z(n24982) );
  IV U24603 ( .A(p_input[5009]), .Z(n24647) );
  XOR U24604 ( .A(n24984), .B(n24985), .Z(n24980) );
  AND U24605 ( .A(n24986), .B(n24987), .Z(n24985) );
  XNOR U24606 ( .A(p_input[5040]), .B(n24984), .Z(n24987) );
  XNOR U24607 ( .A(n24984), .B(n24656), .Z(n24986) );
  IV U24608 ( .A(p_input[5008]), .Z(n24656) );
  XOR U24609 ( .A(n24988), .B(n24989), .Z(n24984) );
  AND U24610 ( .A(n24990), .B(n24991), .Z(n24989) );
  XNOR U24611 ( .A(p_input[5039]), .B(n24988), .Z(n24991) );
  XNOR U24612 ( .A(n24988), .B(n24665), .Z(n24990) );
  IV U24613 ( .A(p_input[5007]), .Z(n24665) );
  XOR U24614 ( .A(n24992), .B(n24993), .Z(n24988) );
  AND U24615 ( .A(n24994), .B(n24995), .Z(n24993) );
  XNOR U24616 ( .A(p_input[5038]), .B(n24992), .Z(n24995) );
  XNOR U24617 ( .A(n24992), .B(n24674), .Z(n24994) );
  IV U24618 ( .A(p_input[5006]), .Z(n24674) );
  XOR U24619 ( .A(n24996), .B(n24997), .Z(n24992) );
  AND U24620 ( .A(n24998), .B(n24999), .Z(n24997) );
  XNOR U24621 ( .A(p_input[5037]), .B(n24996), .Z(n24999) );
  XNOR U24622 ( .A(n24996), .B(n24683), .Z(n24998) );
  IV U24623 ( .A(p_input[5005]), .Z(n24683) );
  XOR U24624 ( .A(n25000), .B(n25001), .Z(n24996) );
  AND U24625 ( .A(n25002), .B(n25003), .Z(n25001) );
  XNOR U24626 ( .A(p_input[5036]), .B(n25000), .Z(n25003) );
  XNOR U24627 ( .A(n25000), .B(n24692), .Z(n25002) );
  IV U24628 ( .A(p_input[5004]), .Z(n24692) );
  XOR U24629 ( .A(n25004), .B(n25005), .Z(n25000) );
  AND U24630 ( .A(n25006), .B(n25007), .Z(n25005) );
  XNOR U24631 ( .A(p_input[5035]), .B(n25004), .Z(n25007) );
  XNOR U24632 ( .A(n25004), .B(n24701), .Z(n25006) );
  IV U24633 ( .A(p_input[5003]), .Z(n24701) );
  XOR U24634 ( .A(n25008), .B(n25009), .Z(n25004) );
  AND U24635 ( .A(n25010), .B(n25011), .Z(n25009) );
  XNOR U24636 ( .A(p_input[5034]), .B(n25008), .Z(n25011) );
  XNOR U24637 ( .A(n25008), .B(n24710), .Z(n25010) );
  IV U24638 ( .A(p_input[5002]), .Z(n24710) );
  XOR U24639 ( .A(n25012), .B(n25013), .Z(n25008) );
  AND U24640 ( .A(n25014), .B(n25015), .Z(n25013) );
  XNOR U24641 ( .A(p_input[5033]), .B(n25012), .Z(n25015) );
  XNOR U24642 ( .A(n25012), .B(n24719), .Z(n25014) );
  IV U24643 ( .A(p_input[5001]), .Z(n24719) );
  XOR U24644 ( .A(n25016), .B(n25017), .Z(n25012) );
  AND U24645 ( .A(n25018), .B(n25019), .Z(n25017) );
  XNOR U24646 ( .A(p_input[5032]), .B(n25016), .Z(n25019) );
  XNOR U24647 ( .A(n25016), .B(n24728), .Z(n25018) );
  IV U24648 ( .A(p_input[5000]), .Z(n24728) );
  XOR U24649 ( .A(n25020), .B(n25021), .Z(n25016) );
  AND U24650 ( .A(n25022), .B(n25023), .Z(n25021) );
  XNOR U24651 ( .A(p_input[5031]), .B(n25020), .Z(n25023) );
  XNOR U24652 ( .A(n25020), .B(n24737), .Z(n25022) );
  IV U24653 ( .A(p_input[4999]), .Z(n24737) );
  XOR U24654 ( .A(n25024), .B(n25025), .Z(n25020) );
  AND U24655 ( .A(n25026), .B(n25027), .Z(n25025) );
  XNOR U24656 ( .A(p_input[5030]), .B(n25024), .Z(n25027) );
  XNOR U24657 ( .A(n25024), .B(n24746), .Z(n25026) );
  IV U24658 ( .A(p_input[4998]), .Z(n24746) );
  XOR U24659 ( .A(n25028), .B(n25029), .Z(n25024) );
  AND U24660 ( .A(n25030), .B(n25031), .Z(n25029) );
  XNOR U24661 ( .A(p_input[5029]), .B(n25028), .Z(n25031) );
  XNOR U24662 ( .A(n25028), .B(n24755), .Z(n25030) );
  IV U24663 ( .A(p_input[4997]), .Z(n24755) );
  XOR U24664 ( .A(n25032), .B(n25033), .Z(n25028) );
  AND U24665 ( .A(n25034), .B(n25035), .Z(n25033) );
  XNOR U24666 ( .A(p_input[5028]), .B(n25032), .Z(n25035) );
  XNOR U24667 ( .A(n25032), .B(n24764), .Z(n25034) );
  IV U24668 ( .A(p_input[4996]), .Z(n24764) );
  XOR U24669 ( .A(n25036), .B(n25037), .Z(n25032) );
  AND U24670 ( .A(n25038), .B(n25039), .Z(n25037) );
  XNOR U24671 ( .A(p_input[5027]), .B(n25036), .Z(n25039) );
  XNOR U24672 ( .A(n25036), .B(n24773), .Z(n25038) );
  IV U24673 ( .A(p_input[4995]), .Z(n24773) );
  XOR U24674 ( .A(n25040), .B(n25041), .Z(n25036) );
  AND U24675 ( .A(n25042), .B(n25043), .Z(n25041) );
  XNOR U24676 ( .A(p_input[5026]), .B(n25040), .Z(n25043) );
  XNOR U24677 ( .A(n25040), .B(n24782), .Z(n25042) );
  IV U24678 ( .A(p_input[4994]), .Z(n24782) );
  XNOR U24679 ( .A(n25044), .B(n25045), .Z(n25040) );
  AND U24680 ( .A(n25046), .B(n25047), .Z(n25045) );
  XOR U24681 ( .A(p_input[5025]), .B(n25044), .Z(n25047) );
  XNOR U24682 ( .A(p_input[4993]), .B(n25044), .Z(n25046) );
  AND U24683 ( .A(p_input[5024]), .B(n25048), .Z(n25044) );
  IV U24684 ( .A(p_input[4992]), .Z(n25048) );
  XOR U24685 ( .A(n25049), .B(n25050), .Z(n24138) );
  AND U24686 ( .A(n525), .B(n25051), .Z(n25050) );
  XNOR U24687 ( .A(n25052), .B(n25049), .Z(n25051) );
  XOR U24688 ( .A(n25053), .B(n25054), .Z(n525) );
  AND U24689 ( .A(n25055), .B(n25056), .Z(n25054) );
  XNOR U24690 ( .A(n24153), .B(n25053), .Z(n25056) );
  AND U24691 ( .A(p_input[4991]), .B(p_input[4959]), .Z(n24153) );
  XNOR U24692 ( .A(n25053), .B(n24150), .Z(n25055) );
  IV U24693 ( .A(n25057), .Z(n24150) );
  AND U24694 ( .A(p_input[4895]), .B(p_input[4927]), .Z(n25057) );
  XOR U24695 ( .A(n25058), .B(n25059), .Z(n25053) );
  AND U24696 ( .A(n25060), .B(n25061), .Z(n25059) );
  XOR U24697 ( .A(n25058), .B(n24165), .Z(n25061) );
  XNOR U24698 ( .A(p_input[4958]), .B(n25062), .Z(n24165) );
  AND U24699 ( .A(n375), .B(n25063), .Z(n25062) );
  XOR U24700 ( .A(p_input[4990]), .B(p_input[4958]), .Z(n25063) );
  XNOR U24701 ( .A(n24162), .B(n25058), .Z(n25060) );
  XOR U24702 ( .A(n25064), .B(n25065), .Z(n24162) );
  AND U24703 ( .A(n372), .B(n25066), .Z(n25065) );
  XOR U24704 ( .A(p_input[4926]), .B(p_input[4894]), .Z(n25066) );
  XOR U24705 ( .A(n25067), .B(n25068), .Z(n25058) );
  AND U24706 ( .A(n25069), .B(n25070), .Z(n25068) );
  XOR U24707 ( .A(n25067), .B(n24177), .Z(n25070) );
  XNOR U24708 ( .A(p_input[4957]), .B(n25071), .Z(n24177) );
  AND U24709 ( .A(n375), .B(n25072), .Z(n25071) );
  XOR U24710 ( .A(p_input[4989]), .B(p_input[4957]), .Z(n25072) );
  XNOR U24711 ( .A(n24174), .B(n25067), .Z(n25069) );
  XOR U24712 ( .A(n25073), .B(n25074), .Z(n24174) );
  AND U24713 ( .A(n372), .B(n25075), .Z(n25074) );
  XOR U24714 ( .A(p_input[4925]), .B(p_input[4893]), .Z(n25075) );
  XOR U24715 ( .A(n25076), .B(n25077), .Z(n25067) );
  AND U24716 ( .A(n25078), .B(n25079), .Z(n25077) );
  XOR U24717 ( .A(n25076), .B(n24189), .Z(n25079) );
  XNOR U24718 ( .A(p_input[4956]), .B(n25080), .Z(n24189) );
  AND U24719 ( .A(n375), .B(n25081), .Z(n25080) );
  XOR U24720 ( .A(p_input[4988]), .B(p_input[4956]), .Z(n25081) );
  XNOR U24721 ( .A(n24186), .B(n25076), .Z(n25078) );
  XOR U24722 ( .A(n25082), .B(n25083), .Z(n24186) );
  AND U24723 ( .A(n372), .B(n25084), .Z(n25083) );
  XOR U24724 ( .A(p_input[4924]), .B(p_input[4892]), .Z(n25084) );
  XOR U24725 ( .A(n25085), .B(n25086), .Z(n25076) );
  AND U24726 ( .A(n25087), .B(n25088), .Z(n25086) );
  XOR U24727 ( .A(n25085), .B(n24201), .Z(n25088) );
  XNOR U24728 ( .A(p_input[4955]), .B(n25089), .Z(n24201) );
  AND U24729 ( .A(n375), .B(n25090), .Z(n25089) );
  XOR U24730 ( .A(p_input[4987]), .B(p_input[4955]), .Z(n25090) );
  XNOR U24731 ( .A(n24198), .B(n25085), .Z(n25087) );
  XOR U24732 ( .A(n25091), .B(n25092), .Z(n24198) );
  AND U24733 ( .A(n372), .B(n25093), .Z(n25092) );
  XOR U24734 ( .A(p_input[4923]), .B(p_input[4891]), .Z(n25093) );
  XOR U24735 ( .A(n25094), .B(n25095), .Z(n25085) );
  AND U24736 ( .A(n25096), .B(n25097), .Z(n25095) );
  XOR U24737 ( .A(n25094), .B(n24213), .Z(n25097) );
  XNOR U24738 ( .A(p_input[4954]), .B(n25098), .Z(n24213) );
  AND U24739 ( .A(n375), .B(n25099), .Z(n25098) );
  XOR U24740 ( .A(p_input[4986]), .B(p_input[4954]), .Z(n25099) );
  XNOR U24741 ( .A(n24210), .B(n25094), .Z(n25096) );
  XOR U24742 ( .A(n25100), .B(n25101), .Z(n24210) );
  AND U24743 ( .A(n372), .B(n25102), .Z(n25101) );
  XOR U24744 ( .A(p_input[4922]), .B(p_input[4890]), .Z(n25102) );
  XOR U24745 ( .A(n25103), .B(n25104), .Z(n25094) );
  AND U24746 ( .A(n25105), .B(n25106), .Z(n25104) );
  XOR U24747 ( .A(n25103), .B(n24225), .Z(n25106) );
  XNOR U24748 ( .A(p_input[4953]), .B(n25107), .Z(n24225) );
  AND U24749 ( .A(n375), .B(n25108), .Z(n25107) );
  XOR U24750 ( .A(p_input[4985]), .B(p_input[4953]), .Z(n25108) );
  XNOR U24751 ( .A(n24222), .B(n25103), .Z(n25105) );
  XOR U24752 ( .A(n25109), .B(n25110), .Z(n24222) );
  AND U24753 ( .A(n372), .B(n25111), .Z(n25110) );
  XOR U24754 ( .A(p_input[4921]), .B(p_input[4889]), .Z(n25111) );
  XOR U24755 ( .A(n25112), .B(n25113), .Z(n25103) );
  AND U24756 ( .A(n25114), .B(n25115), .Z(n25113) );
  XOR U24757 ( .A(n25112), .B(n24237), .Z(n25115) );
  XNOR U24758 ( .A(p_input[4952]), .B(n25116), .Z(n24237) );
  AND U24759 ( .A(n375), .B(n25117), .Z(n25116) );
  XOR U24760 ( .A(p_input[4984]), .B(p_input[4952]), .Z(n25117) );
  XNOR U24761 ( .A(n24234), .B(n25112), .Z(n25114) );
  XOR U24762 ( .A(n25118), .B(n25119), .Z(n24234) );
  AND U24763 ( .A(n372), .B(n25120), .Z(n25119) );
  XOR U24764 ( .A(p_input[4920]), .B(p_input[4888]), .Z(n25120) );
  XOR U24765 ( .A(n25121), .B(n25122), .Z(n25112) );
  AND U24766 ( .A(n25123), .B(n25124), .Z(n25122) );
  XOR U24767 ( .A(n25121), .B(n24249), .Z(n25124) );
  XNOR U24768 ( .A(p_input[4951]), .B(n25125), .Z(n24249) );
  AND U24769 ( .A(n375), .B(n25126), .Z(n25125) );
  XOR U24770 ( .A(p_input[4983]), .B(p_input[4951]), .Z(n25126) );
  XNOR U24771 ( .A(n24246), .B(n25121), .Z(n25123) );
  XOR U24772 ( .A(n25127), .B(n25128), .Z(n24246) );
  AND U24773 ( .A(n372), .B(n25129), .Z(n25128) );
  XOR U24774 ( .A(p_input[4919]), .B(p_input[4887]), .Z(n25129) );
  XOR U24775 ( .A(n25130), .B(n25131), .Z(n25121) );
  AND U24776 ( .A(n25132), .B(n25133), .Z(n25131) );
  XOR U24777 ( .A(n25130), .B(n24261), .Z(n25133) );
  XNOR U24778 ( .A(p_input[4950]), .B(n25134), .Z(n24261) );
  AND U24779 ( .A(n375), .B(n25135), .Z(n25134) );
  XOR U24780 ( .A(p_input[4982]), .B(p_input[4950]), .Z(n25135) );
  XNOR U24781 ( .A(n24258), .B(n25130), .Z(n25132) );
  XOR U24782 ( .A(n25136), .B(n25137), .Z(n24258) );
  AND U24783 ( .A(n372), .B(n25138), .Z(n25137) );
  XOR U24784 ( .A(p_input[4918]), .B(p_input[4886]), .Z(n25138) );
  XOR U24785 ( .A(n25139), .B(n25140), .Z(n25130) );
  AND U24786 ( .A(n25141), .B(n25142), .Z(n25140) );
  XOR U24787 ( .A(n25139), .B(n24273), .Z(n25142) );
  XNOR U24788 ( .A(p_input[4949]), .B(n25143), .Z(n24273) );
  AND U24789 ( .A(n375), .B(n25144), .Z(n25143) );
  XOR U24790 ( .A(p_input[4981]), .B(p_input[4949]), .Z(n25144) );
  XNOR U24791 ( .A(n24270), .B(n25139), .Z(n25141) );
  XOR U24792 ( .A(n25145), .B(n25146), .Z(n24270) );
  AND U24793 ( .A(n372), .B(n25147), .Z(n25146) );
  XOR U24794 ( .A(p_input[4917]), .B(p_input[4885]), .Z(n25147) );
  XOR U24795 ( .A(n25148), .B(n25149), .Z(n25139) );
  AND U24796 ( .A(n25150), .B(n25151), .Z(n25149) );
  XOR U24797 ( .A(n25148), .B(n24285), .Z(n25151) );
  XNOR U24798 ( .A(p_input[4948]), .B(n25152), .Z(n24285) );
  AND U24799 ( .A(n375), .B(n25153), .Z(n25152) );
  XOR U24800 ( .A(p_input[4980]), .B(p_input[4948]), .Z(n25153) );
  XNOR U24801 ( .A(n24282), .B(n25148), .Z(n25150) );
  XOR U24802 ( .A(n25154), .B(n25155), .Z(n24282) );
  AND U24803 ( .A(n372), .B(n25156), .Z(n25155) );
  XOR U24804 ( .A(p_input[4916]), .B(p_input[4884]), .Z(n25156) );
  XOR U24805 ( .A(n25157), .B(n25158), .Z(n25148) );
  AND U24806 ( .A(n25159), .B(n25160), .Z(n25158) );
  XOR U24807 ( .A(n25157), .B(n24297), .Z(n25160) );
  XNOR U24808 ( .A(p_input[4947]), .B(n25161), .Z(n24297) );
  AND U24809 ( .A(n375), .B(n25162), .Z(n25161) );
  XOR U24810 ( .A(p_input[4979]), .B(p_input[4947]), .Z(n25162) );
  XNOR U24811 ( .A(n24294), .B(n25157), .Z(n25159) );
  XOR U24812 ( .A(n25163), .B(n25164), .Z(n24294) );
  AND U24813 ( .A(n372), .B(n25165), .Z(n25164) );
  XOR U24814 ( .A(p_input[4915]), .B(p_input[4883]), .Z(n25165) );
  XOR U24815 ( .A(n25166), .B(n25167), .Z(n25157) );
  AND U24816 ( .A(n25168), .B(n25169), .Z(n25167) );
  XOR U24817 ( .A(n25166), .B(n24309), .Z(n25169) );
  XNOR U24818 ( .A(p_input[4946]), .B(n25170), .Z(n24309) );
  AND U24819 ( .A(n375), .B(n25171), .Z(n25170) );
  XOR U24820 ( .A(p_input[4978]), .B(p_input[4946]), .Z(n25171) );
  XNOR U24821 ( .A(n24306), .B(n25166), .Z(n25168) );
  XOR U24822 ( .A(n25172), .B(n25173), .Z(n24306) );
  AND U24823 ( .A(n372), .B(n25174), .Z(n25173) );
  XOR U24824 ( .A(p_input[4914]), .B(p_input[4882]), .Z(n25174) );
  XOR U24825 ( .A(n25175), .B(n25176), .Z(n25166) );
  AND U24826 ( .A(n25177), .B(n25178), .Z(n25176) );
  XOR U24827 ( .A(n25175), .B(n24321), .Z(n25178) );
  XNOR U24828 ( .A(p_input[4945]), .B(n25179), .Z(n24321) );
  AND U24829 ( .A(n375), .B(n25180), .Z(n25179) );
  XOR U24830 ( .A(p_input[4977]), .B(p_input[4945]), .Z(n25180) );
  XNOR U24831 ( .A(n24318), .B(n25175), .Z(n25177) );
  XOR U24832 ( .A(n25181), .B(n25182), .Z(n24318) );
  AND U24833 ( .A(n372), .B(n25183), .Z(n25182) );
  XOR U24834 ( .A(p_input[4913]), .B(p_input[4881]), .Z(n25183) );
  XOR U24835 ( .A(n25184), .B(n25185), .Z(n25175) );
  AND U24836 ( .A(n25186), .B(n25187), .Z(n25185) );
  XOR U24837 ( .A(n25184), .B(n24333), .Z(n25187) );
  XNOR U24838 ( .A(p_input[4944]), .B(n25188), .Z(n24333) );
  AND U24839 ( .A(n375), .B(n25189), .Z(n25188) );
  XOR U24840 ( .A(p_input[4976]), .B(p_input[4944]), .Z(n25189) );
  XNOR U24841 ( .A(n24330), .B(n25184), .Z(n25186) );
  XOR U24842 ( .A(n25190), .B(n25191), .Z(n24330) );
  AND U24843 ( .A(n372), .B(n25192), .Z(n25191) );
  XOR U24844 ( .A(p_input[4912]), .B(p_input[4880]), .Z(n25192) );
  XOR U24845 ( .A(n25193), .B(n25194), .Z(n25184) );
  AND U24846 ( .A(n25195), .B(n25196), .Z(n25194) );
  XOR U24847 ( .A(n25193), .B(n24345), .Z(n25196) );
  XNOR U24848 ( .A(p_input[4943]), .B(n25197), .Z(n24345) );
  AND U24849 ( .A(n375), .B(n25198), .Z(n25197) );
  XOR U24850 ( .A(p_input[4975]), .B(p_input[4943]), .Z(n25198) );
  XNOR U24851 ( .A(n24342), .B(n25193), .Z(n25195) );
  XOR U24852 ( .A(n25199), .B(n25200), .Z(n24342) );
  AND U24853 ( .A(n372), .B(n25201), .Z(n25200) );
  XOR U24854 ( .A(p_input[4911]), .B(p_input[4879]), .Z(n25201) );
  XOR U24855 ( .A(n25202), .B(n25203), .Z(n25193) );
  AND U24856 ( .A(n25204), .B(n25205), .Z(n25203) );
  XOR U24857 ( .A(n25202), .B(n24357), .Z(n25205) );
  XNOR U24858 ( .A(p_input[4942]), .B(n25206), .Z(n24357) );
  AND U24859 ( .A(n375), .B(n25207), .Z(n25206) );
  XOR U24860 ( .A(p_input[4974]), .B(p_input[4942]), .Z(n25207) );
  XNOR U24861 ( .A(n24354), .B(n25202), .Z(n25204) );
  XOR U24862 ( .A(n25208), .B(n25209), .Z(n24354) );
  AND U24863 ( .A(n372), .B(n25210), .Z(n25209) );
  XOR U24864 ( .A(p_input[4910]), .B(p_input[4878]), .Z(n25210) );
  XOR U24865 ( .A(n25211), .B(n25212), .Z(n25202) );
  AND U24866 ( .A(n25213), .B(n25214), .Z(n25212) );
  XOR U24867 ( .A(n25211), .B(n24369), .Z(n25214) );
  XNOR U24868 ( .A(p_input[4941]), .B(n25215), .Z(n24369) );
  AND U24869 ( .A(n375), .B(n25216), .Z(n25215) );
  XOR U24870 ( .A(p_input[4973]), .B(p_input[4941]), .Z(n25216) );
  XNOR U24871 ( .A(n24366), .B(n25211), .Z(n25213) );
  XOR U24872 ( .A(n25217), .B(n25218), .Z(n24366) );
  AND U24873 ( .A(n372), .B(n25219), .Z(n25218) );
  XOR U24874 ( .A(p_input[4909]), .B(p_input[4877]), .Z(n25219) );
  XOR U24875 ( .A(n25220), .B(n25221), .Z(n25211) );
  AND U24876 ( .A(n25222), .B(n25223), .Z(n25221) );
  XOR U24877 ( .A(n25220), .B(n24381), .Z(n25223) );
  XNOR U24878 ( .A(p_input[4940]), .B(n25224), .Z(n24381) );
  AND U24879 ( .A(n375), .B(n25225), .Z(n25224) );
  XOR U24880 ( .A(p_input[4972]), .B(p_input[4940]), .Z(n25225) );
  XNOR U24881 ( .A(n24378), .B(n25220), .Z(n25222) );
  XOR U24882 ( .A(n25226), .B(n25227), .Z(n24378) );
  AND U24883 ( .A(n372), .B(n25228), .Z(n25227) );
  XOR U24884 ( .A(p_input[4908]), .B(p_input[4876]), .Z(n25228) );
  XOR U24885 ( .A(n25229), .B(n25230), .Z(n25220) );
  AND U24886 ( .A(n25231), .B(n25232), .Z(n25230) );
  XOR U24887 ( .A(n25229), .B(n24393), .Z(n25232) );
  XNOR U24888 ( .A(p_input[4939]), .B(n25233), .Z(n24393) );
  AND U24889 ( .A(n375), .B(n25234), .Z(n25233) );
  XOR U24890 ( .A(p_input[4971]), .B(p_input[4939]), .Z(n25234) );
  XNOR U24891 ( .A(n24390), .B(n25229), .Z(n25231) );
  XOR U24892 ( .A(n25235), .B(n25236), .Z(n24390) );
  AND U24893 ( .A(n372), .B(n25237), .Z(n25236) );
  XOR U24894 ( .A(p_input[4907]), .B(p_input[4875]), .Z(n25237) );
  XOR U24895 ( .A(n25238), .B(n25239), .Z(n25229) );
  AND U24896 ( .A(n25240), .B(n25241), .Z(n25239) );
  XOR U24897 ( .A(n25238), .B(n24405), .Z(n25241) );
  XNOR U24898 ( .A(p_input[4938]), .B(n25242), .Z(n24405) );
  AND U24899 ( .A(n375), .B(n25243), .Z(n25242) );
  XOR U24900 ( .A(p_input[4970]), .B(p_input[4938]), .Z(n25243) );
  XNOR U24901 ( .A(n24402), .B(n25238), .Z(n25240) );
  XOR U24902 ( .A(n25244), .B(n25245), .Z(n24402) );
  AND U24903 ( .A(n372), .B(n25246), .Z(n25245) );
  XOR U24904 ( .A(p_input[4906]), .B(p_input[4874]), .Z(n25246) );
  XOR U24905 ( .A(n25247), .B(n25248), .Z(n25238) );
  AND U24906 ( .A(n25249), .B(n25250), .Z(n25248) );
  XOR U24907 ( .A(n25247), .B(n24417), .Z(n25250) );
  XNOR U24908 ( .A(p_input[4937]), .B(n25251), .Z(n24417) );
  AND U24909 ( .A(n375), .B(n25252), .Z(n25251) );
  XOR U24910 ( .A(p_input[4969]), .B(p_input[4937]), .Z(n25252) );
  XNOR U24911 ( .A(n24414), .B(n25247), .Z(n25249) );
  XOR U24912 ( .A(n25253), .B(n25254), .Z(n24414) );
  AND U24913 ( .A(n372), .B(n25255), .Z(n25254) );
  XOR U24914 ( .A(p_input[4905]), .B(p_input[4873]), .Z(n25255) );
  XOR U24915 ( .A(n25256), .B(n25257), .Z(n25247) );
  AND U24916 ( .A(n25258), .B(n25259), .Z(n25257) );
  XOR U24917 ( .A(n25256), .B(n24429), .Z(n25259) );
  XNOR U24918 ( .A(p_input[4936]), .B(n25260), .Z(n24429) );
  AND U24919 ( .A(n375), .B(n25261), .Z(n25260) );
  XOR U24920 ( .A(p_input[4968]), .B(p_input[4936]), .Z(n25261) );
  XNOR U24921 ( .A(n24426), .B(n25256), .Z(n25258) );
  XOR U24922 ( .A(n25262), .B(n25263), .Z(n24426) );
  AND U24923 ( .A(n372), .B(n25264), .Z(n25263) );
  XOR U24924 ( .A(p_input[4904]), .B(p_input[4872]), .Z(n25264) );
  XOR U24925 ( .A(n25265), .B(n25266), .Z(n25256) );
  AND U24926 ( .A(n25267), .B(n25268), .Z(n25266) );
  XOR U24927 ( .A(n25265), .B(n24441), .Z(n25268) );
  XNOR U24928 ( .A(p_input[4935]), .B(n25269), .Z(n24441) );
  AND U24929 ( .A(n375), .B(n25270), .Z(n25269) );
  XOR U24930 ( .A(p_input[4967]), .B(p_input[4935]), .Z(n25270) );
  XNOR U24931 ( .A(n24438), .B(n25265), .Z(n25267) );
  XOR U24932 ( .A(n25271), .B(n25272), .Z(n24438) );
  AND U24933 ( .A(n372), .B(n25273), .Z(n25272) );
  XOR U24934 ( .A(p_input[4903]), .B(p_input[4871]), .Z(n25273) );
  XOR U24935 ( .A(n25274), .B(n25275), .Z(n25265) );
  AND U24936 ( .A(n25276), .B(n25277), .Z(n25275) );
  XOR U24937 ( .A(n25274), .B(n24453), .Z(n25277) );
  XNOR U24938 ( .A(p_input[4934]), .B(n25278), .Z(n24453) );
  AND U24939 ( .A(n375), .B(n25279), .Z(n25278) );
  XOR U24940 ( .A(p_input[4966]), .B(p_input[4934]), .Z(n25279) );
  XNOR U24941 ( .A(n24450), .B(n25274), .Z(n25276) );
  XOR U24942 ( .A(n25280), .B(n25281), .Z(n24450) );
  AND U24943 ( .A(n372), .B(n25282), .Z(n25281) );
  XOR U24944 ( .A(p_input[4902]), .B(p_input[4870]), .Z(n25282) );
  XOR U24945 ( .A(n25283), .B(n25284), .Z(n25274) );
  AND U24946 ( .A(n25285), .B(n25286), .Z(n25284) );
  XOR U24947 ( .A(n25283), .B(n24465), .Z(n25286) );
  XNOR U24948 ( .A(p_input[4933]), .B(n25287), .Z(n24465) );
  AND U24949 ( .A(n375), .B(n25288), .Z(n25287) );
  XOR U24950 ( .A(p_input[4965]), .B(p_input[4933]), .Z(n25288) );
  XNOR U24951 ( .A(n24462), .B(n25283), .Z(n25285) );
  XOR U24952 ( .A(n25289), .B(n25290), .Z(n24462) );
  AND U24953 ( .A(n372), .B(n25291), .Z(n25290) );
  XOR U24954 ( .A(p_input[4901]), .B(p_input[4869]), .Z(n25291) );
  XOR U24955 ( .A(n25292), .B(n25293), .Z(n25283) );
  AND U24956 ( .A(n25294), .B(n25295), .Z(n25293) );
  XOR U24957 ( .A(n25292), .B(n24477), .Z(n25295) );
  XNOR U24958 ( .A(p_input[4932]), .B(n25296), .Z(n24477) );
  AND U24959 ( .A(n375), .B(n25297), .Z(n25296) );
  XOR U24960 ( .A(p_input[4964]), .B(p_input[4932]), .Z(n25297) );
  XNOR U24961 ( .A(n24474), .B(n25292), .Z(n25294) );
  XOR U24962 ( .A(n25298), .B(n25299), .Z(n24474) );
  AND U24963 ( .A(n372), .B(n25300), .Z(n25299) );
  XOR U24964 ( .A(p_input[4900]), .B(p_input[4868]), .Z(n25300) );
  XOR U24965 ( .A(n25301), .B(n25302), .Z(n25292) );
  AND U24966 ( .A(n25303), .B(n25304), .Z(n25302) );
  XOR U24967 ( .A(n25301), .B(n24489), .Z(n25304) );
  XNOR U24968 ( .A(p_input[4931]), .B(n25305), .Z(n24489) );
  AND U24969 ( .A(n375), .B(n25306), .Z(n25305) );
  XOR U24970 ( .A(p_input[4963]), .B(p_input[4931]), .Z(n25306) );
  XNOR U24971 ( .A(n24486), .B(n25301), .Z(n25303) );
  XOR U24972 ( .A(n25307), .B(n25308), .Z(n24486) );
  AND U24973 ( .A(n372), .B(n25309), .Z(n25308) );
  XOR U24974 ( .A(p_input[4899]), .B(p_input[4867]), .Z(n25309) );
  XOR U24975 ( .A(n25310), .B(n25311), .Z(n25301) );
  AND U24976 ( .A(n25312), .B(n25313), .Z(n25311) );
  XOR U24977 ( .A(n25310), .B(n24501), .Z(n25313) );
  XNOR U24978 ( .A(p_input[4930]), .B(n25314), .Z(n24501) );
  AND U24979 ( .A(n375), .B(n25315), .Z(n25314) );
  XOR U24980 ( .A(p_input[4962]), .B(p_input[4930]), .Z(n25315) );
  XNOR U24981 ( .A(n24498), .B(n25310), .Z(n25312) );
  XOR U24982 ( .A(n25316), .B(n25317), .Z(n24498) );
  AND U24983 ( .A(n372), .B(n25318), .Z(n25317) );
  XOR U24984 ( .A(p_input[4898]), .B(p_input[4866]), .Z(n25318) );
  XOR U24985 ( .A(n25319), .B(n25320), .Z(n25310) );
  AND U24986 ( .A(n25321), .B(n25322), .Z(n25320) );
  XNOR U24987 ( .A(n25323), .B(n24514), .Z(n25322) );
  XNOR U24988 ( .A(p_input[4929]), .B(n25324), .Z(n24514) );
  AND U24989 ( .A(n375), .B(n25325), .Z(n25324) );
  XNOR U24990 ( .A(p_input[4961]), .B(n25326), .Z(n25325) );
  IV U24991 ( .A(p_input[4929]), .Z(n25326) );
  XNOR U24992 ( .A(n24511), .B(n25319), .Z(n25321) );
  XNOR U24993 ( .A(p_input[4865]), .B(n25327), .Z(n24511) );
  AND U24994 ( .A(n372), .B(n25328), .Z(n25327) );
  XOR U24995 ( .A(p_input[4897]), .B(p_input[4865]), .Z(n25328) );
  IV U24996 ( .A(n25323), .Z(n25319) );
  AND U24997 ( .A(n25049), .B(n25052), .Z(n25323) );
  XOR U24998 ( .A(p_input[4928]), .B(n25329), .Z(n25052) );
  AND U24999 ( .A(n375), .B(n25330), .Z(n25329) );
  XOR U25000 ( .A(p_input[4960]), .B(p_input[4928]), .Z(n25330) );
  XOR U25001 ( .A(n25331), .B(n25332), .Z(n375) );
  AND U25002 ( .A(n25333), .B(n25334), .Z(n25332) );
  XNOR U25003 ( .A(p_input[4991]), .B(n25331), .Z(n25334) );
  XOR U25004 ( .A(n25331), .B(p_input[4959]), .Z(n25333) );
  XOR U25005 ( .A(n25335), .B(n25336), .Z(n25331) );
  AND U25006 ( .A(n25337), .B(n25338), .Z(n25336) );
  XNOR U25007 ( .A(p_input[4990]), .B(n25335), .Z(n25338) );
  XOR U25008 ( .A(n25335), .B(p_input[4958]), .Z(n25337) );
  XOR U25009 ( .A(n25339), .B(n25340), .Z(n25335) );
  AND U25010 ( .A(n25341), .B(n25342), .Z(n25340) );
  XNOR U25011 ( .A(p_input[4989]), .B(n25339), .Z(n25342) );
  XOR U25012 ( .A(n25339), .B(p_input[4957]), .Z(n25341) );
  XOR U25013 ( .A(n25343), .B(n25344), .Z(n25339) );
  AND U25014 ( .A(n25345), .B(n25346), .Z(n25344) );
  XNOR U25015 ( .A(p_input[4988]), .B(n25343), .Z(n25346) );
  XOR U25016 ( .A(n25343), .B(p_input[4956]), .Z(n25345) );
  XOR U25017 ( .A(n25347), .B(n25348), .Z(n25343) );
  AND U25018 ( .A(n25349), .B(n25350), .Z(n25348) );
  XNOR U25019 ( .A(p_input[4987]), .B(n25347), .Z(n25350) );
  XOR U25020 ( .A(n25347), .B(p_input[4955]), .Z(n25349) );
  XOR U25021 ( .A(n25351), .B(n25352), .Z(n25347) );
  AND U25022 ( .A(n25353), .B(n25354), .Z(n25352) );
  XNOR U25023 ( .A(p_input[4986]), .B(n25351), .Z(n25354) );
  XOR U25024 ( .A(n25351), .B(p_input[4954]), .Z(n25353) );
  XOR U25025 ( .A(n25355), .B(n25356), .Z(n25351) );
  AND U25026 ( .A(n25357), .B(n25358), .Z(n25356) );
  XNOR U25027 ( .A(p_input[4985]), .B(n25355), .Z(n25358) );
  XOR U25028 ( .A(n25355), .B(p_input[4953]), .Z(n25357) );
  XOR U25029 ( .A(n25359), .B(n25360), .Z(n25355) );
  AND U25030 ( .A(n25361), .B(n25362), .Z(n25360) );
  XNOR U25031 ( .A(p_input[4984]), .B(n25359), .Z(n25362) );
  XOR U25032 ( .A(n25359), .B(p_input[4952]), .Z(n25361) );
  XOR U25033 ( .A(n25363), .B(n25364), .Z(n25359) );
  AND U25034 ( .A(n25365), .B(n25366), .Z(n25364) );
  XNOR U25035 ( .A(p_input[4983]), .B(n25363), .Z(n25366) );
  XOR U25036 ( .A(n25363), .B(p_input[4951]), .Z(n25365) );
  XOR U25037 ( .A(n25367), .B(n25368), .Z(n25363) );
  AND U25038 ( .A(n25369), .B(n25370), .Z(n25368) );
  XNOR U25039 ( .A(p_input[4982]), .B(n25367), .Z(n25370) );
  XOR U25040 ( .A(n25367), .B(p_input[4950]), .Z(n25369) );
  XOR U25041 ( .A(n25371), .B(n25372), .Z(n25367) );
  AND U25042 ( .A(n25373), .B(n25374), .Z(n25372) );
  XNOR U25043 ( .A(p_input[4981]), .B(n25371), .Z(n25374) );
  XOR U25044 ( .A(n25371), .B(p_input[4949]), .Z(n25373) );
  XOR U25045 ( .A(n25375), .B(n25376), .Z(n25371) );
  AND U25046 ( .A(n25377), .B(n25378), .Z(n25376) );
  XNOR U25047 ( .A(p_input[4980]), .B(n25375), .Z(n25378) );
  XOR U25048 ( .A(n25375), .B(p_input[4948]), .Z(n25377) );
  XOR U25049 ( .A(n25379), .B(n25380), .Z(n25375) );
  AND U25050 ( .A(n25381), .B(n25382), .Z(n25380) );
  XNOR U25051 ( .A(p_input[4979]), .B(n25379), .Z(n25382) );
  XOR U25052 ( .A(n25379), .B(p_input[4947]), .Z(n25381) );
  XOR U25053 ( .A(n25383), .B(n25384), .Z(n25379) );
  AND U25054 ( .A(n25385), .B(n25386), .Z(n25384) );
  XNOR U25055 ( .A(p_input[4978]), .B(n25383), .Z(n25386) );
  XOR U25056 ( .A(n25383), .B(p_input[4946]), .Z(n25385) );
  XOR U25057 ( .A(n25387), .B(n25388), .Z(n25383) );
  AND U25058 ( .A(n25389), .B(n25390), .Z(n25388) );
  XNOR U25059 ( .A(p_input[4977]), .B(n25387), .Z(n25390) );
  XOR U25060 ( .A(n25387), .B(p_input[4945]), .Z(n25389) );
  XOR U25061 ( .A(n25391), .B(n25392), .Z(n25387) );
  AND U25062 ( .A(n25393), .B(n25394), .Z(n25392) );
  XNOR U25063 ( .A(p_input[4976]), .B(n25391), .Z(n25394) );
  XOR U25064 ( .A(n25391), .B(p_input[4944]), .Z(n25393) );
  XOR U25065 ( .A(n25395), .B(n25396), .Z(n25391) );
  AND U25066 ( .A(n25397), .B(n25398), .Z(n25396) );
  XNOR U25067 ( .A(p_input[4975]), .B(n25395), .Z(n25398) );
  XOR U25068 ( .A(n25395), .B(p_input[4943]), .Z(n25397) );
  XOR U25069 ( .A(n25399), .B(n25400), .Z(n25395) );
  AND U25070 ( .A(n25401), .B(n25402), .Z(n25400) );
  XNOR U25071 ( .A(p_input[4974]), .B(n25399), .Z(n25402) );
  XOR U25072 ( .A(n25399), .B(p_input[4942]), .Z(n25401) );
  XOR U25073 ( .A(n25403), .B(n25404), .Z(n25399) );
  AND U25074 ( .A(n25405), .B(n25406), .Z(n25404) );
  XNOR U25075 ( .A(p_input[4973]), .B(n25403), .Z(n25406) );
  XOR U25076 ( .A(n25403), .B(p_input[4941]), .Z(n25405) );
  XOR U25077 ( .A(n25407), .B(n25408), .Z(n25403) );
  AND U25078 ( .A(n25409), .B(n25410), .Z(n25408) );
  XNOR U25079 ( .A(p_input[4972]), .B(n25407), .Z(n25410) );
  XOR U25080 ( .A(n25407), .B(p_input[4940]), .Z(n25409) );
  XOR U25081 ( .A(n25411), .B(n25412), .Z(n25407) );
  AND U25082 ( .A(n25413), .B(n25414), .Z(n25412) );
  XNOR U25083 ( .A(p_input[4971]), .B(n25411), .Z(n25414) );
  XOR U25084 ( .A(n25411), .B(p_input[4939]), .Z(n25413) );
  XOR U25085 ( .A(n25415), .B(n25416), .Z(n25411) );
  AND U25086 ( .A(n25417), .B(n25418), .Z(n25416) );
  XNOR U25087 ( .A(p_input[4970]), .B(n25415), .Z(n25418) );
  XOR U25088 ( .A(n25415), .B(p_input[4938]), .Z(n25417) );
  XOR U25089 ( .A(n25419), .B(n25420), .Z(n25415) );
  AND U25090 ( .A(n25421), .B(n25422), .Z(n25420) );
  XNOR U25091 ( .A(p_input[4969]), .B(n25419), .Z(n25422) );
  XOR U25092 ( .A(n25419), .B(p_input[4937]), .Z(n25421) );
  XOR U25093 ( .A(n25423), .B(n25424), .Z(n25419) );
  AND U25094 ( .A(n25425), .B(n25426), .Z(n25424) );
  XNOR U25095 ( .A(p_input[4968]), .B(n25423), .Z(n25426) );
  XOR U25096 ( .A(n25423), .B(p_input[4936]), .Z(n25425) );
  XOR U25097 ( .A(n25427), .B(n25428), .Z(n25423) );
  AND U25098 ( .A(n25429), .B(n25430), .Z(n25428) );
  XNOR U25099 ( .A(p_input[4967]), .B(n25427), .Z(n25430) );
  XOR U25100 ( .A(n25427), .B(p_input[4935]), .Z(n25429) );
  XOR U25101 ( .A(n25431), .B(n25432), .Z(n25427) );
  AND U25102 ( .A(n25433), .B(n25434), .Z(n25432) );
  XNOR U25103 ( .A(p_input[4966]), .B(n25431), .Z(n25434) );
  XOR U25104 ( .A(n25431), .B(p_input[4934]), .Z(n25433) );
  XOR U25105 ( .A(n25435), .B(n25436), .Z(n25431) );
  AND U25106 ( .A(n25437), .B(n25438), .Z(n25436) );
  XNOR U25107 ( .A(p_input[4965]), .B(n25435), .Z(n25438) );
  XOR U25108 ( .A(n25435), .B(p_input[4933]), .Z(n25437) );
  XOR U25109 ( .A(n25439), .B(n25440), .Z(n25435) );
  AND U25110 ( .A(n25441), .B(n25442), .Z(n25440) );
  XNOR U25111 ( .A(p_input[4964]), .B(n25439), .Z(n25442) );
  XOR U25112 ( .A(n25439), .B(p_input[4932]), .Z(n25441) );
  XOR U25113 ( .A(n25443), .B(n25444), .Z(n25439) );
  AND U25114 ( .A(n25445), .B(n25446), .Z(n25444) );
  XNOR U25115 ( .A(p_input[4963]), .B(n25443), .Z(n25446) );
  XOR U25116 ( .A(n25443), .B(p_input[4931]), .Z(n25445) );
  XOR U25117 ( .A(n25447), .B(n25448), .Z(n25443) );
  AND U25118 ( .A(n25449), .B(n25450), .Z(n25448) );
  XNOR U25119 ( .A(p_input[4962]), .B(n25447), .Z(n25450) );
  XOR U25120 ( .A(n25447), .B(p_input[4930]), .Z(n25449) );
  XNOR U25121 ( .A(n25451), .B(n25452), .Z(n25447) );
  AND U25122 ( .A(n25453), .B(n25454), .Z(n25452) );
  XOR U25123 ( .A(p_input[4961]), .B(n25451), .Z(n25454) );
  XNOR U25124 ( .A(p_input[4929]), .B(n25451), .Z(n25453) );
  AND U25125 ( .A(p_input[4960]), .B(n25455), .Z(n25451) );
  IV U25126 ( .A(p_input[4928]), .Z(n25455) );
  XNOR U25127 ( .A(p_input[4864]), .B(n25456), .Z(n25049) );
  AND U25128 ( .A(n372), .B(n25457), .Z(n25456) );
  XOR U25129 ( .A(p_input[4896]), .B(p_input[4864]), .Z(n25457) );
  XOR U25130 ( .A(n25458), .B(n25459), .Z(n372) );
  AND U25131 ( .A(n25460), .B(n25461), .Z(n25459) );
  XNOR U25132 ( .A(p_input[4927]), .B(n25458), .Z(n25461) );
  XOR U25133 ( .A(n25458), .B(p_input[4895]), .Z(n25460) );
  XOR U25134 ( .A(n25462), .B(n25463), .Z(n25458) );
  AND U25135 ( .A(n25464), .B(n25465), .Z(n25463) );
  XNOR U25136 ( .A(p_input[4926]), .B(n25462), .Z(n25465) );
  XNOR U25137 ( .A(n25462), .B(n25064), .Z(n25464) );
  IV U25138 ( .A(p_input[4894]), .Z(n25064) );
  XOR U25139 ( .A(n25466), .B(n25467), .Z(n25462) );
  AND U25140 ( .A(n25468), .B(n25469), .Z(n25467) );
  XNOR U25141 ( .A(p_input[4925]), .B(n25466), .Z(n25469) );
  XNOR U25142 ( .A(n25466), .B(n25073), .Z(n25468) );
  IV U25143 ( .A(p_input[4893]), .Z(n25073) );
  XOR U25144 ( .A(n25470), .B(n25471), .Z(n25466) );
  AND U25145 ( .A(n25472), .B(n25473), .Z(n25471) );
  XNOR U25146 ( .A(p_input[4924]), .B(n25470), .Z(n25473) );
  XNOR U25147 ( .A(n25470), .B(n25082), .Z(n25472) );
  IV U25148 ( .A(p_input[4892]), .Z(n25082) );
  XOR U25149 ( .A(n25474), .B(n25475), .Z(n25470) );
  AND U25150 ( .A(n25476), .B(n25477), .Z(n25475) );
  XNOR U25151 ( .A(p_input[4923]), .B(n25474), .Z(n25477) );
  XNOR U25152 ( .A(n25474), .B(n25091), .Z(n25476) );
  IV U25153 ( .A(p_input[4891]), .Z(n25091) );
  XOR U25154 ( .A(n25478), .B(n25479), .Z(n25474) );
  AND U25155 ( .A(n25480), .B(n25481), .Z(n25479) );
  XNOR U25156 ( .A(p_input[4922]), .B(n25478), .Z(n25481) );
  XNOR U25157 ( .A(n25478), .B(n25100), .Z(n25480) );
  IV U25158 ( .A(p_input[4890]), .Z(n25100) );
  XOR U25159 ( .A(n25482), .B(n25483), .Z(n25478) );
  AND U25160 ( .A(n25484), .B(n25485), .Z(n25483) );
  XNOR U25161 ( .A(p_input[4921]), .B(n25482), .Z(n25485) );
  XNOR U25162 ( .A(n25482), .B(n25109), .Z(n25484) );
  IV U25163 ( .A(p_input[4889]), .Z(n25109) );
  XOR U25164 ( .A(n25486), .B(n25487), .Z(n25482) );
  AND U25165 ( .A(n25488), .B(n25489), .Z(n25487) );
  XNOR U25166 ( .A(p_input[4920]), .B(n25486), .Z(n25489) );
  XNOR U25167 ( .A(n25486), .B(n25118), .Z(n25488) );
  IV U25168 ( .A(p_input[4888]), .Z(n25118) );
  XOR U25169 ( .A(n25490), .B(n25491), .Z(n25486) );
  AND U25170 ( .A(n25492), .B(n25493), .Z(n25491) );
  XNOR U25171 ( .A(p_input[4919]), .B(n25490), .Z(n25493) );
  XNOR U25172 ( .A(n25490), .B(n25127), .Z(n25492) );
  IV U25173 ( .A(p_input[4887]), .Z(n25127) );
  XOR U25174 ( .A(n25494), .B(n25495), .Z(n25490) );
  AND U25175 ( .A(n25496), .B(n25497), .Z(n25495) );
  XNOR U25176 ( .A(p_input[4918]), .B(n25494), .Z(n25497) );
  XNOR U25177 ( .A(n25494), .B(n25136), .Z(n25496) );
  IV U25178 ( .A(p_input[4886]), .Z(n25136) );
  XOR U25179 ( .A(n25498), .B(n25499), .Z(n25494) );
  AND U25180 ( .A(n25500), .B(n25501), .Z(n25499) );
  XNOR U25181 ( .A(p_input[4917]), .B(n25498), .Z(n25501) );
  XNOR U25182 ( .A(n25498), .B(n25145), .Z(n25500) );
  IV U25183 ( .A(p_input[4885]), .Z(n25145) );
  XOR U25184 ( .A(n25502), .B(n25503), .Z(n25498) );
  AND U25185 ( .A(n25504), .B(n25505), .Z(n25503) );
  XNOR U25186 ( .A(p_input[4916]), .B(n25502), .Z(n25505) );
  XNOR U25187 ( .A(n25502), .B(n25154), .Z(n25504) );
  IV U25188 ( .A(p_input[4884]), .Z(n25154) );
  XOR U25189 ( .A(n25506), .B(n25507), .Z(n25502) );
  AND U25190 ( .A(n25508), .B(n25509), .Z(n25507) );
  XNOR U25191 ( .A(p_input[4915]), .B(n25506), .Z(n25509) );
  XNOR U25192 ( .A(n25506), .B(n25163), .Z(n25508) );
  IV U25193 ( .A(p_input[4883]), .Z(n25163) );
  XOR U25194 ( .A(n25510), .B(n25511), .Z(n25506) );
  AND U25195 ( .A(n25512), .B(n25513), .Z(n25511) );
  XNOR U25196 ( .A(p_input[4914]), .B(n25510), .Z(n25513) );
  XNOR U25197 ( .A(n25510), .B(n25172), .Z(n25512) );
  IV U25198 ( .A(p_input[4882]), .Z(n25172) );
  XOR U25199 ( .A(n25514), .B(n25515), .Z(n25510) );
  AND U25200 ( .A(n25516), .B(n25517), .Z(n25515) );
  XNOR U25201 ( .A(p_input[4913]), .B(n25514), .Z(n25517) );
  XNOR U25202 ( .A(n25514), .B(n25181), .Z(n25516) );
  IV U25203 ( .A(p_input[4881]), .Z(n25181) );
  XOR U25204 ( .A(n25518), .B(n25519), .Z(n25514) );
  AND U25205 ( .A(n25520), .B(n25521), .Z(n25519) );
  XNOR U25206 ( .A(p_input[4912]), .B(n25518), .Z(n25521) );
  XNOR U25207 ( .A(n25518), .B(n25190), .Z(n25520) );
  IV U25208 ( .A(p_input[4880]), .Z(n25190) );
  XOR U25209 ( .A(n25522), .B(n25523), .Z(n25518) );
  AND U25210 ( .A(n25524), .B(n25525), .Z(n25523) );
  XNOR U25211 ( .A(p_input[4911]), .B(n25522), .Z(n25525) );
  XNOR U25212 ( .A(n25522), .B(n25199), .Z(n25524) );
  IV U25213 ( .A(p_input[4879]), .Z(n25199) );
  XOR U25214 ( .A(n25526), .B(n25527), .Z(n25522) );
  AND U25215 ( .A(n25528), .B(n25529), .Z(n25527) );
  XNOR U25216 ( .A(p_input[4910]), .B(n25526), .Z(n25529) );
  XNOR U25217 ( .A(n25526), .B(n25208), .Z(n25528) );
  IV U25218 ( .A(p_input[4878]), .Z(n25208) );
  XOR U25219 ( .A(n25530), .B(n25531), .Z(n25526) );
  AND U25220 ( .A(n25532), .B(n25533), .Z(n25531) );
  XNOR U25221 ( .A(p_input[4909]), .B(n25530), .Z(n25533) );
  XNOR U25222 ( .A(n25530), .B(n25217), .Z(n25532) );
  IV U25223 ( .A(p_input[4877]), .Z(n25217) );
  XOR U25224 ( .A(n25534), .B(n25535), .Z(n25530) );
  AND U25225 ( .A(n25536), .B(n25537), .Z(n25535) );
  XNOR U25226 ( .A(p_input[4908]), .B(n25534), .Z(n25537) );
  XNOR U25227 ( .A(n25534), .B(n25226), .Z(n25536) );
  IV U25228 ( .A(p_input[4876]), .Z(n25226) );
  XOR U25229 ( .A(n25538), .B(n25539), .Z(n25534) );
  AND U25230 ( .A(n25540), .B(n25541), .Z(n25539) );
  XNOR U25231 ( .A(p_input[4907]), .B(n25538), .Z(n25541) );
  XNOR U25232 ( .A(n25538), .B(n25235), .Z(n25540) );
  IV U25233 ( .A(p_input[4875]), .Z(n25235) );
  XOR U25234 ( .A(n25542), .B(n25543), .Z(n25538) );
  AND U25235 ( .A(n25544), .B(n25545), .Z(n25543) );
  XNOR U25236 ( .A(p_input[4906]), .B(n25542), .Z(n25545) );
  XNOR U25237 ( .A(n25542), .B(n25244), .Z(n25544) );
  IV U25238 ( .A(p_input[4874]), .Z(n25244) );
  XOR U25239 ( .A(n25546), .B(n25547), .Z(n25542) );
  AND U25240 ( .A(n25548), .B(n25549), .Z(n25547) );
  XNOR U25241 ( .A(p_input[4905]), .B(n25546), .Z(n25549) );
  XNOR U25242 ( .A(n25546), .B(n25253), .Z(n25548) );
  IV U25243 ( .A(p_input[4873]), .Z(n25253) );
  XOR U25244 ( .A(n25550), .B(n25551), .Z(n25546) );
  AND U25245 ( .A(n25552), .B(n25553), .Z(n25551) );
  XNOR U25246 ( .A(p_input[4904]), .B(n25550), .Z(n25553) );
  XNOR U25247 ( .A(n25550), .B(n25262), .Z(n25552) );
  IV U25248 ( .A(p_input[4872]), .Z(n25262) );
  XOR U25249 ( .A(n25554), .B(n25555), .Z(n25550) );
  AND U25250 ( .A(n25556), .B(n25557), .Z(n25555) );
  XNOR U25251 ( .A(p_input[4903]), .B(n25554), .Z(n25557) );
  XNOR U25252 ( .A(n25554), .B(n25271), .Z(n25556) );
  IV U25253 ( .A(p_input[4871]), .Z(n25271) );
  XOR U25254 ( .A(n25558), .B(n25559), .Z(n25554) );
  AND U25255 ( .A(n25560), .B(n25561), .Z(n25559) );
  XNOR U25256 ( .A(p_input[4902]), .B(n25558), .Z(n25561) );
  XNOR U25257 ( .A(n25558), .B(n25280), .Z(n25560) );
  IV U25258 ( .A(p_input[4870]), .Z(n25280) );
  XOR U25259 ( .A(n25562), .B(n25563), .Z(n25558) );
  AND U25260 ( .A(n25564), .B(n25565), .Z(n25563) );
  XNOR U25261 ( .A(p_input[4901]), .B(n25562), .Z(n25565) );
  XNOR U25262 ( .A(n25562), .B(n25289), .Z(n25564) );
  IV U25263 ( .A(p_input[4869]), .Z(n25289) );
  XOR U25264 ( .A(n25566), .B(n25567), .Z(n25562) );
  AND U25265 ( .A(n25568), .B(n25569), .Z(n25567) );
  XNOR U25266 ( .A(p_input[4900]), .B(n25566), .Z(n25569) );
  XNOR U25267 ( .A(n25566), .B(n25298), .Z(n25568) );
  IV U25268 ( .A(p_input[4868]), .Z(n25298) );
  XOR U25269 ( .A(n25570), .B(n25571), .Z(n25566) );
  AND U25270 ( .A(n25572), .B(n25573), .Z(n25571) );
  XNOR U25271 ( .A(p_input[4899]), .B(n25570), .Z(n25573) );
  XNOR U25272 ( .A(n25570), .B(n25307), .Z(n25572) );
  IV U25273 ( .A(p_input[4867]), .Z(n25307) );
  XOR U25274 ( .A(n25574), .B(n25575), .Z(n25570) );
  AND U25275 ( .A(n25576), .B(n25577), .Z(n25575) );
  XNOR U25276 ( .A(p_input[4898]), .B(n25574), .Z(n25577) );
  XNOR U25277 ( .A(n25574), .B(n25316), .Z(n25576) );
  IV U25278 ( .A(p_input[4866]), .Z(n25316) );
  XNOR U25279 ( .A(n25578), .B(n25579), .Z(n25574) );
  AND U25280 ( .A(n25580), .B(n25581), .Z(n25579) );
  XOR U25281 ( .A(p_input[4897]), .B(n25578), .Z(n25581) );
  XNOR U25282 ( .A(p_input[4865]), .B(n25578), .Z(n25580) );
  AND U25283 ( .A(p_input[4896]), .B(n25582), .Z(n25578) );
  IV U25284 ( .A(p_input[4864]), .Z(n25582) );
  XOR U25285 ( .A(n25583), .B(n25584), .Z(n23761) );
  AND U25286 ( .A(n853), .B(n25585), .Z(n25584) );
  XNOR U25287 ( .A(n25586), .B(n25583), .Z(n25585) );
  XOR U25288 ( .A(n25587), .B(n25588), .Z(n853) );
  AND U25289 ( .A(n25589), .B(n25590), .Z(n25588) );
  XOR U25290 ( .A(n25587), .B(n23776), .Z(n25590) );
  XNOR U25291 ( .A(n25591), .B(n25592), .Z(n23776) );
  AND U25292 ( .A(n25593), .B(n531), .Z(n25592) );
  AND U25293 ( .A(n25591), .B(n25594), .Z(n25593) );
  XNOR U25294 ( .A(n23773), .B(n25587), .Z(n25589) );
  XOR U25295 ( .A(n25595), .B(n25596), .Z(n23773) );
  AND U25296 ( .A(n25597), .B(n528), .Z(n25596) );
  NOR U25297 ( .A(n25595), .B(n25598), .Z(n25597) );
  XOR U25298 ( .A(n25599), .B(n25600), .Z(n25587) );
  AND U25299 ( .A(n25601), .B(n25602), .Z(n25600) );
  XOR U25300 ( .A(n25599), .B(n23788), .Z(n25602) );
  XOR U25301 ( .A(n25603), .B(n25604), .Z(n23788) );
  AND U25302 ( .A(n531), .B(n25605), .Z(n25604) );
  XOR U25303 ( .A(n25606), .B(n25603), .Z(n25605) );
  XNOR U25304 ( .A(n23785), .B(n25599), .Z(n25601) );
  XOR U25305 ( .A(n25607), .B(n25608), .Z(n23785) );
  AND U25306 ( .A(n528), .B(n25609), .Z(n25608) );
  XOR U25307 ( .A(n25610), .B(n25607), .Z(n25609) );
  XOR U25308 ( .A(n25611), .B(n25612), .Z(n25599) );
  AND U25309 ( .A(n25613), .B(n25614), .Z(n25612) );
  XOR U25310 ( .A(n25611), .B(n23800), .Z(n25614) );
  XOR U25311 ( .A(n25615), .B(n25616), .Z(n23800) );
  AND U25312 ( .A(n531), .B(n25617), .Z(n25616) );
  XOR U25313 ( .A(n25618), .B(n25615), .Z(n25617) );
  XNOR U25314 ( .A(n23797), .B(n25611), .Z(n25613) );
  XOR U25315 ( .A(n25619), .B(n25620), .Z(n23797) );
  AND U25316 ( .A(n528), .B(n25621), .Z(n25620) );
  XOR U25317 ( .A(n25622), .B(n25619), .Z(n25621) );
  XOR U25318 ( .A(n25623), .B(n25624), .Z(n25611) );
  AND U25319 ( .A(n25625), .B(n25626), .Z(n25624) );
  XOR U25320 ( .A(n25623), .B(n23812), .Z(n25626) );
  XOR U25321 ( .A(n25627), .B(n25628), .Z(n23812) );
  AND U25322 ( .A(n531), .B(n25629), .Z(n25628) );
  XOR U25323 ( .A(n25630), .B(n25627), .Z(n25629) );
  XNOR U25324 ( .A(n23809), .B(n25623), .Z(n25625) );
  XOR U25325 ( .A(n25631), .B(n25632), .Z(n23809) );
  AND U25326 ( .A(n528), .B(n25633), .Z(n25632) );
  XOR U25327 ( .A(n25634), .B(n25631), .Z(n25633) );
  XOR U25328 ( .A(n25635), .B(n25636), .Z(n25623) );
  AND U25329 ( .A(n25637), .B(n25638), .Z(n25636) );
  XOR U25330 ( .A(n25635), .B(n23824), .Z(n25638) );
  XOR U25331 ( .A(n25639), .B(n25640), .Z(n23824) );
  AND U25332 ( .A(n531), .B(n25641), .Z(n25640) );
  XOR U25333 ( .A(n25642), .B(n25639), .Z(n25641) );
  XNOR U25334 ( .A(n23821), .B(n25635), .Z(n25637) );
  XOR U25335 ( .A(n25643), .B(n25644), .Z(n23821) );
  AND U25336 ( .A(n528), .B(n25645), .Z(n25644) );
  XOR U25337 ( .A(n25646), .B(n25643), .Z(n25645) );
  XOR U25338 ( .A(n25647), .B(n25648), .Z(n25635) );
  AND U25339 ( .A(n25649), .B(n25650), .Z(n25648) );
  XOR U25340 ( .A(n25647), .B(n23836), .Z(n25650) );
  XOR U25341 ( .A(n25651), .B(n25652), .Z(n23836) );
  AND U25342 ( .A(n531), .B(n25653), .Z(n25652) );
  XOR U25343 ( .A(n25654), .B(n25651), .Z(n25653) );
  XNOR U25344 ( .A(n23833), .B(n25647), .Z(n25649) );
  XOR U25345 ( .A(n25655), .B(n25656), .Z(n23833) );
  AND U25346 ( .A(n528), .B(n25657), .Z(n25656) );
  XOR U25347 ( .A(n25658), .B(n25655), .Z(n25657) );
  XOR U25348 ( .A(n25659), .B(n25660), .Z(n25647) );
  AND U25349 ( .A(n25661), .B(n25662), .Z(n25660) );
  XOR U25350 ( .A(n25659), .B(n23848), .Z(n25662) );
  XOR U25351 ( .A(n25663), .B(n25664), .Z(n23848) );
  AND U25352 ( .A(n531), .B(n25665), .Z(n25664) );
  XOR U25353 ( .A(n25666), .B(n25663), .Z(n25665) );
  XNOR U25354 ( .A(n23845), .B(n25659), .Z(n25661) );
  XOR U25355 ( .A(n25667), .B(n25668), .Z(n23845) );
  AND U25356 ( .A(n528), .B(n25669), .Z(n25668) );
  XOR U25357 ( .A(n25670), .B(n25667), .Z(n25669) );
  XOR U25358 ( .A(n25671), .B(n25672), .Z(n25659) );
  AND U25359 ( .A(n25673), .B(n25674), .Z(n25672) );
  XOR U25360 ( .A(n25671), .B(n23860), .Z(n25674) );
  XOR U25361 ( .A(n25675), .B(n25676), .Z(n23860) );
  AND U25362 ( .A(n531), .B(n25677), .Z(n25676) );
  XOR U25363 ( .A(n25678), .B(n25675), .Z(n25677) );
  XNOR U25364 ( .A(n23857), .B(n25671), .Z(n25673) );
  XOR U25365 ( .A(n25679), .B(n25680), .Z(n23857) );
  AND U25366 ( .A(n528), .B(n25681), .Z(n25680) );
  XOR U25367 ( .A(n25682), .B(n25679), .Z(n25681) );
  XOR U25368 ( .A(n25683), .B(n25684), .Z(n25671) );
  AND U25369 ( .A(n25685), .B(n25686), .Z(n25684) );
  XOR U25370 ( .A(n25683), .B(n23872), .Z(n25686) );
  XOR U25371 ( .A(n25687), .B(n25688), .Z(n23872) );
  AND U25372 ( .A(n531), .B(n25689), .Z(n25688) );
  XOR U25373 ( .A(n25690), .B(n25687), .Z(n25689) );
  XNOR U25374 ( .A(n23869), .B(n25683), .Z(n25685) );
  XOR U25375 ( .A(n25691), .B(n25692), .Z(n23869) );
  AND U25376 ( .A(n528), .B(n25693), .Z(n25692) );
  XOR U25377 ( .A(n25694), .B(n25691), .Z(n25693) );
  XOR U25378 ( .A(n25695), .B(n25696), .Z(n25683) );
  AND U25379 ( .A(n25697), .B(n25698), .Z(n25696) );
  XOR U25380 ( .A(n25695), .B(n23884), .Z(n25698) );
  XOR U25381 ( .A(n25699), .B(n25700), .Z(n23884) );
  AND U25382 ( .A(n531), .B(n25701), .Z(n25700) );
  XOR U25383 ( .A(n25702), .B(n25699), .Z(n25701) );
  XNOR U25384 ( .A(n23881), .B(n25695), .Z(n25697) );
  XOR U25385 ( .A(n25703), .B(n25704), .Z(n23881) );
  AND U25386 ( .A(n528), .B(n25705), .Z(n25704) );
  XOR U25387 ( .A(n25706), .B(n25703), .Z(n25705) );
  XOR U25388 ( .A(n25707), .B(n25708), .Z(n25695) );
  AND U25389 ( .A(n25709), .B(n25710), .Z(n25708) );
  XOR U25390 ( .A(n25707), .B(n23896), .Z(n25710) );
  XOR U25391 ( .A(n25711), .B(n25712), .Z(n23896) );
  AND U25392 ( .A(n531), .B(n25713), .Z(n25712) );
  XOR U25393 ( .A(n25714), .B(n25711), .Z(n25713) );
  XNOR U25394 ( .A(n23893), .B(n25707), .Z(n25709) );
  XOR U25395 ( .A(n25715), .B(n25716), .Z(n23893) );
  AND U25396 ( .A(n528), .B(n25717), .Z(n25716) );
  XOR U25397 ( .A(n25718), .B(n25715), .Z(n25717) );
  XOR U25398 ( .A(n25719), .B(n25720), .Z(n25707) );
  AND U25399 ( .A(n25721), .B(n25722), .Z(n25720) );
  XOR U25400 ( .A(n25719), .B(n23908), .Z(n25722) );
  XOR U25401 ( .A(n25723), .B(n25724), .Z(n23908) );
  AND U25402 ( .A(n531), .B(n25725), .Z(n25724) );
  XOR U25403 ( .A(n25726), .B(n25723), .Z(n25725) );
  XNOR U25404 ( .A(n23905), .B(n25719), .Z(n25721) );
  XOR U25405 ( .A(n25727), .B(n25728), .Z(n23905) );
  AND U25406 ( .A(n528), .B(n25729), .Z(n25728) );
  XOR U25407 ( .A(n25730), .B(n25727), .Z(n25729) );
  XOR U25408 ( .A(n25731), .B(n25732), .Z(n25719) );
  AND U25409 ( .A(n25733), .B(n25734), .Z(n25732) );
  XOR U25410 ( .A(n25731), .B(n23920), .Z(n25734) );
  XOR U25411 ( .A(n25735), .B(n25736), .Z(n23920) );
  AND U25412 ( .A(n531), .B(n25737), .Z(n25736) );
  XOR U25413 ( .A(n25738), .B(n25735), .Z(n25737) );
  XNOR U25414 ( .A(n23917), .B(n25731), .Z(n25733) );
  XOR U25415 ( .A(n25739), .B(n25740), .Z(n23917) );
  AND U25416 ( .A(n528), .B(n25741), .Z(n25740) );
  XOR U25417 ( .A(n25742), .B(n25739), .Z(n25741) );
  XOR U25418 ( .A(n25743), .B(n25744), .Z(n25731) );
  AND U25419 ( .A(n25745), .B(n25746), .Z(n25744) );
  XOR U25420 ( .A(n25743), .B(n23932), .Z(n25746) );
  XOR U25421 ( .A(n25747), .B(n25748), .Z(n23932) );
  AND U25422 ( .A(n531), .B(n25749), .Z(n25748) );
  XOR U25423 ( .A(n25750), .B(n25747), .Z(n25749) );
  XNOR U25424 ( .A(n23929), .B(n25743), .Z(n25745) );
  XOR U25425 ( .A(n25751), .B(n25752), .Z(n23929) );
  AND U25426 ( .A(n528), .B(n25753), .Z(n25752) );
  XOR U25427 ( .A(n25754), .B(n25751), .Z(n25753) );
  XOR U25428 ( .A(n25755), .B(n25756), .Z(n25743) );
  AND U25429 ( .A(n25757), .B(n25758), .Z(n25756) );
  XOR U25430 ( .A(n25755), .B(n23944), .Z(n25758) );
  XOR U25431 ( .A(n25759), .B(n25760), .Z(n23944) );
  AND U25432 ( .A(n531), .B(n25761), .Z(n25760) );
  XOR U25433 ( .A(n25762), .B(n25759), .Z(n25761) );
  XNOR U25434 ( .A(n23941), .B(n25755), .Z(n25757) );
  XOR U25435 ( .A(n25763), .B(n25764), .Z(n23941) );
  AND U25436 ( .A(n528), .B(n25765), .Z(n25764) );
  XOR U25437 ( .A(n25766), .B(n25763), .Z(n25765) );
  XOR U25438 ( .A(n25767), .B(n25768), .Z(n25755) );
  AND U25439 ( .A(n25769), .B(n25770), .Z(n25768) );
  XOR U25440 ( .A(n25767), .B(n23956), .Z(n25770) );
  XOR U25441 ( .A(n25771), .B(n25772), .Z(n23956) );
  AND U25442 ( .A(n531), .B(n25773), .Z(n25772) );
  XOR U25443 ( .A(n25774), .B(n25771), .Z(n25773) );
  XNOR U25444 ( .A(n23953), .B(n25767), .Z(n25769) );
  XOR U25445 ( .A(n25775), .B(n25776), .Z(n23953) );
  AND U25446 ( .A(n528), .B(n25777), .Z(n25776) );
  XOR U25447 ( .A(n25778), .B(n25775), .Z(n25777) );
  XOR U25448 ( .A(n25779), .B(n25780), .Z(n25767) );
  AND U25449 ( .A(n25781), .B(n25782), .Z(n25780) );
  XOR U25450 ( .A(n25779), .B(n23968), .Z(n25782) );
  XOR U25451 ( .A(n25783), .B(n25784), .Z(n23968) );
  AND U25452 ( .A(n531), .B(n25785), .Z(n25784) );
  XOR U25453 ( .A(n25786), .B(n25783), .Z(n25785) );
  XNOR U25454 ( .A(n23965), .B(n25779), .Z(n25781) );
  XOR U25455 ( .A(n25787), .B(n25788), .Z(n23965) );
  AND U25456 ( .A(n528), .B(n25789), .Z(n25788) );
  XOR U25457 ( .A(n25790), .B(n25787), .Z(n25789) );
  XOR U25458 ( .A(n25791), .B(n25792), .Z(n25779) );
  AND U25459 ( .A(n25793), .B(n25794), .Z(n25792) );
  XOR U25460 ( .A(n25791), .B(n23980), .Z(n25794) );
  XOR U25461 ( .A(n25795), .B(n25796), .Z(n23980) );
  AND U25462 ( .A(n531), .B(n25797), .Z(n25796) );
  XOR U25463 ( .A(n25798), .B(n25795), .Z(n25797) );
  XNOR U25464 ( .A(n23977), .B(n25791), .Z(n25793) );
  XOR U25465 ( .A(n25799), .B(n25800), .Z(n23977) );
  AND U25466 ( .A(n528), .B(n25801), .Z(n25800) );
  XOR U25467 ( .A(n25802), .B(n25799), .Z(n25801) );
  XOR U25468 ( .A(n25803), .B(n25804), .Z(n25791) );
  AND U25469 ( .A(n25805), .B(n25806), .Z(n25804) );
  XOR U25470 ( .A(n25803), .B(n23992), .Z(n25806) );
  XOR U25471 ( .A(n25807), .B(n25808), .Z(n23992) );
  AND U25472 ( .A(n531), .B(n25809), .Z(n25808) );
  XOR U25473 ( .A(n25810), .B(n25807), .Z(n25809) );
  XNOR U25474 ( .A(n23989), .B(n25803), .Z(n25805) );
  XOR U25475 ( .A(n25811), .B(n25812), .Z(n23989) );
  AND U25476 ( .A(n528), .B(n25813), .Z(n25812) );
  XOR U25477 ( .A(n25814), .B(n25811), .Z(n25813) );
  XOR U25478 ( .A(n25815), .B(n25816), .Z(n25803) );
  AND U25479 ( .A(n25817), .B(n25818), .Z(n25816) );
  XOR U25480 ( .A(n25815), .B(n24004), .Z(n25818) );
  XOR U25481 ( .A(n25819), .B(n25820), .Z(n24004) );
  AND U25482 ( .A(n531), .B(n25821), .Z(n25820) );
  XOR U25483 ( .A(n25822), .B(n25819), .Z(n25821) );
  XNOR U25484 ( .A(n24001), .B(n25815), .Z(n25817) );
  XOR U25485 ( .A(n25823), .B(n25824), .Z(n24001) );
  AND U25486 ( .A(n528), .B(n25825), .Z(n25824) );
  XOR U25487 ( .A(n25826), .B(n25823), .Z(n25825) );
  XOR U25488 ( .A(n25827), .B(n25828), .Z(n25815) );
  AND U25489 ( .A(n25829), .B(n25830), .Z(n25828) );
  XOR U25490 ( .A(n25827), .B(n24016), .Z(n25830) );
  XOR U25491 ( .A(n25831), .B(n25832), .Z(n24016) );
  AND U25492 ( .A(n531), .B(n25833), .Z(n25832) );
  XOR U25493 ( .A(n25834), .B(n25831), .Z(n25833) );
  XNOR U25494 ( .A(n24013), .B(n25827), .Z(n25829) );
  XOR U25495 ( .A(n25835), .B(n25836), .Z(n24013) );
  AND U25496 ( .A(n528), .B(n25837), .Z(n25836) );
  XOR U25497 ( .A(n25838), .B(n25835), .Z(n25837) );
  XOR U25498 ( .A(n25839), .B(n25840), .Z(n25827) );
  AND U25499 ( .A(n25841), .B(n25842), .Z(n25840) );
  XOR U25500 ( .A(n25839), .B(n24028), .Z(n25842) );
  XOR U25501 ( .A(n25843), .B(n25844), .Z(n24028) );
  AND U25502 ( .A(n531), .B(n25845), .Z(n25844) );
  XOR U25503 ( .A(n25846), .B(n25843), .Z(n25845) );
  XNOR U25504 ( .A(n24025), .B(n25839), .Z(n25841) );
  XOR U25505 ( .A(n25847), .B(n25848), .Z(n24025) );
  AND U25506 ( .A(n528), .B(n25849), .Z(n25848) );
  XOR U25507 ( .A(n25850), .B(n25847), .Z(n25849) );
  XOR U25508 ( .A(n25851), .B(n25852), .Z(n25839) );
  AND U25509 ( .A(n25853), .B(n25854), .Z(n25852) );
  XOR U25510 ( .A(n25851), .B(n24040), .Z(n25854) );
  XOR U25511 ( .A(n25855), .B(n25856), .Z(n24040) );
  AND U25512 ( .A(n531), .B(n25857), .Z(n25856) );
  XOR U25513 ( .A(n25858), .B(n25855), .Z(n25857) );
  XNOR U25514 ( .A(n24037), .B(n25851), .Z(n25853) );
  XOR U25515 ( .A(n25859), .B(n25860), .Z(n24037) );
  AND U25516 ( .A(n528), .B(n25861), .Z(n25860) );
  XOR U25517 ( .A(n25862), .B(n25859), .Z(n25861) );
  XOR U25518 ( .A(n25863), .B(n25864), .Z(n25851) );
  AND U25519 ( .A(n25865), .B(n25866), .Z(n25864) );
  XOR U25520 ( .A(n25863), .B(n24052), .Z(n25866) );
  XOR U25521 ( .A(n25867), .B(n25868), .Z(n24052) );
  AND U25522 ( .A(n531), .B(n25869), .Z(n25868) );
  XOR U25523 ( .A(n25870), .B(n25867), .Z(n25869) );
  XNOR U25524 ( .A(n24049), .B(n25863), .Z(n25865) );
  XOR U25525 ( .A(n25871), .B(n25872), .Z(n24049) );
  AND U25526 ( .A(n528), .B(n25873), .Z(n25872) );
  XOR U25527 ( .A(n25874), .B(n25871), .Z(n25873) );
  XOR U25528 ( .A(n25875), .B(n25876), .Z(n25863) );
  AND U25529 ( .A(n25877), .B(n25878), .Z(n25876) );
  XOR U25530 ( .A(n25875), .B(n24064), .Z(n25878) );
  XOR U25531 ( .A(n25879), .B(n25880), .Z(n24064) );
  AND U25532 ( .A(n531), .B(n25881), .Z(n25880) );
  XOR U25533 ( .A(n25882), .B(n25879), .Z(n25881) );
  XNOR U25534 ( .A(n24061), .B(n25875), .Z(n25877) );
  XOR U25535 ( .A(n25883), .B(n25884), .Z(n24061) );
  AND U25536 ( .A(n528), .B(n25885), .Z(n25884) );
  XOR U25537 ( .A(n25886), .B(n25883), .Z(n25885) );
  XOR U25538 ( .A(n25887), .B(n25888), .Z(n25875) );
  AND U25539 ( .A(n25889), .B(n25890), .Z(n25888) );
  XOR U25540 ( .A(n25887), .B(n24076), .Z(n25890) );
  XOR U25541 ( .A(n25891), .B(n25892), .Z(n24076) );
  AND U25542 ( .A(n531), .B(n25893), .Z(n25892) );
  XOR U25543 ( .A(n25894), .B(n25891), .Z(n25893) );
  XNOR U25544 ( .A(n24073), .B(n25887), .Z(n25889) );
  XOR U25545 ( .A(n25895), .B(n25896), .Z(n24073) );
  AND U25546 ( .A(n528), .B(n25897), .Z(n25896) );
  XOR U25547 ( .A(n25898), .B(n25895), .Z(n25897) );
  XOR U25548 ( .A(n25899), .B(n25900), .Z(n25887) );
  AND U25549 ( .A(n25901), .B(n25902), .Z(n25900) );
  XOR U25550 ( .A(n25899), .B(n24088), .Z(n25902) );
  XOR U25551 ( .A(n25903), .B(n25904), .Z(n24088) );
  AND U25552 ( .A(n531), .B(n25905), .Z(n25904) );
  XOR U25553 ( .A(n25906), .B(n25903), .Z(n25905) );
  XNOR U25554 ( .A(n24085), .B(n25899), .Z(n25901) );
  XOR U25555 ( .A(n25907), .B(n25908), .Z(n24085) );
  AND U25556 ( .A(n528), .B(n25909), .Z(n25908) );
  XOR U25557 ( .A(n25910), .B(n25907), .Z(n25909) );
  XOR U25558 ( .A(n25911), .B(n25912), .Z(n25899) );
  AND U25559 ( .A(n25913), .B(n25914), .Z(n25912) );
  XOR U25560 ( .A(n25911), .B(n24100), .Z(n25914) );
  XOR U25561 ( .A(n25915), .B(n25916), .Z(n24100) );
  AND U25562 ( .A(n531), .B(n25917), .Z(n25916) );
  XOR U25563 ( .A(n25918), .B(n25915), .Z(n25917) );
  XNOR U25564 ( .A(n24097), .B(n25911), .Z(n25913) );
  XOR U25565 ( .A(n25919), .B(n25920), .Z(n24097) );
  AND U25566 ( .A(n528), .B(n25921), .Z(n25920) );
  XOR U25567 ( .A(n25922), .B(n25919), .Z(n25921) );
  XOR U25568 ( .A(n25923), .B(n25924), .Z(n25911) );
  AND U25569 ( .A(n25925), .B(n25926), .Z(n25924) );
  XOR U25570 ( .A(n25923), .B(n24112), .Z(n25926) );
  XOR U25571 ( .A(n25927), .B(n25928), .Z(n24112) );
  AND U25572 ( .A(n531), .B(n25929), .Z(n25928) );
  XOR U25573 ( .A(n25930), .B(n25927), .Z(n25929) );
  XNOR U25574 ( .A(n24109), .B(n25923), .Z(n25925) );
  XOR U25575 ( .A(n25931), .B(n25932), .Z(n24109) );
  AND U25576 ( .A(n528), .B(n25933), .Z(n25932) );
  XOR U25577 ( .A(n25934), .B(n25931), .Z(n25933) );
  XOR U25578 ( .A(n25935), .B(n25936), .Z(n25923) );
  AND U25579 ( .A(n25937), .B(n25938), .Z(n25936) );
  XOR U25580 ( .A(n25935), .B(n24124), .Z(n25938) );
  XOR U25581 ( .A(n25939), .B(n25940), .Z(n24124) );
  AND U25582 ( .A(n531), .B(n25941), .Z(n25940) );
  XOR U25583 ( .A(n25942), .B(n25939), .Z(n25941) );
  XNOR U25584 ( .A(n24121), .B(n25935), .Z(n25937) );
  XOR U25585 ( .A(n25943), .B(n25944), .Z(n24121) );
  AND U25586 ( .A(n528), .B(n25945), .Z(n25944) );
  XOR U25587 ( .A(n25946), .B(n25943), .Z(n25945) );
  XOR U25588 ( .A(n25947), .B(n25948), .Z(n25935) );
  AND U25589 ( .A(n25949), .B(n25950), .Z(n25948) );
  XNOR U25590 ( .A(n25951), .B(n24137), .Z(n25950) );
  XOR U25591 ( .A(n25952), .B(n25953), .Z(n24137) );
  AND U25592 ( .A(n531), .B(n25954), .Z(n25953) );
  XOR U25593 ( .A(n25952), .B(n25955), .Z(n25954) );
  XNOR U25594 ( .A(n24134), .B(n25947), .Z(n25949) );
  XOR U25595 ( .A(n25956), .B(n25957), .Z(n24134) );
  AND U25596 ( .A(n528), .B(n25958), .Z(n25957) );
  XOR U25597 ( .A(n25956), .B(n25959), .Z(n25958) );
  IV U25598 ( .A(n25951), .Z(n25947) );
  AND U25599 ( .A(n25583), .B(n25586), .Z(n25951) );
  XNOR U25600 ( .A(n25960), .B(n25961), .Z(n25586) );
  AND U25601 ( .A(n531), .B(n25962), .Z(n25961) );
  XNOR U25602 ( .A(n25963), .B(n25960), .Z(n25962) );
  XOR U25603 ( .A(n25964), .B(n25965), .Z(n531) );
  AND U25604 ( .A(n25966), .B(n25967), .Z(n25965) );
  XOR U25605 ( .A(n25594), .B(n25964), .Z(n25967) );
  IV U25606 ( .A(n25968), .Z(n25594) );
  AND U25607 ( .A(p_input[4863]), .B(p_input[4831]), .Z(n25968) );
  XOR U25608 ( .A(n25964), .B(n25591), .Z(n25966) );
  AND U25609 ( .A(p_input[4767]), .B(p_input[4799]), .Z(n25591) );
  XOR U25610 ( .A(n25969), .B(n25970), .Z(n25964) );
  AND U25611 ( .A(n25971), .B(n25972), .Z(n25970) );
  XOR U25612 ( .A(n25969), .B(n25606), .Z(n25972) );
  XNOR U25613 ( .A(p_input[4830]), .B(n25973), .Z(n25606) );
  AND U25614 ( .A(n383), .B(n25974), .Z(n25973) );
  XOR U25615 ( .A(p_input[4862]), .B(p_input[4830]), .Z(n25974) );
  XNOR U25616 ( .A(n25603), .B(n25969), .Z(n25971) );
  XOR U25617 ( .A(n25975), .B(n25976), .Z(n25603) );
  AND U25618 ( .A(n381), .B(n25977), .Z(n25976) );
  XOR U25619 ( .A(p_input[4798]), .B(p_input[4766]), .Z(n25977) );
  XOR U25620 ( .A(n25978), .B(n25979), .Z(n25969) );
  AND U25621 ( .A(n25980), .B(n25981), .Z(n25979) );
  XOR U25622 ( .A(n25978), .B(n25618), .Z(n25981) );
  XNOR U25623 ( .A(p_input[4829]), .B(n25982), .Z(n25618) );
  AND U25624 ( .A(n383), .B(n25983), .Z(n25982) );
  XOR U25625 ( .A(p_input[4861]), .B(p_input[4829]), .Z(n25983) );
  XNOR U25626 ( .A(n25615), .B(n25978), .Z(n25980) );
  XOR U25627 ( .A(n25984), .B(n25985), .Z(n25615) );
  AND U25628 ( .A(n381), .B(n25986), .Z(n25985) );
  XOR U25629 ( .A(p_input[4797]), .B(p_input[4765]), .Z(n25986) );
  XOR U25630 ( .A(n25987), .B(n25988), .Z(n25978) );
  AND U25631 ( .A(n25989), .B(n25990), .Z(n25988) );
  XOR U25632 ( .A(n25987), .B(n25630), .Z(n25990) );
  XNOR U25633 ( .A(p_input[4828]), .B(n25991), .Z(n25630) );
  AND U25634 ( .A(n383), .B(n25992), .Z(n25991) );
  XOR U25635 ( .A(p_input[4860]), .B(p_input[4828]), .Z(n25992) );
  XNOR U25636 ( .A(n25627), .B(n25987), .Z(n25989) );
  XOR U25637 ( .A(n25993), .B(n25994), .Z(n25627) );
  AND U25638 ( .A(n381), .B(n25995), .Z(n25994) );
  XOR U25639 ( .A(p_input[4796]), .B(p_input[4764]), .Z(n25995) );
  XOR U25640 ( .A(n25996), .B(n25997), .Z(n25987) );
  AND U25641 ( .A(n25998), .B(n25999), .Z(n25997) );
  XOR U25642 ( .A(n25996), .B(n25642), .Z(n25999) );
  XNOR U25643 ( .A(p_input[4827]), .B(n26000), .Z(n25642) );
  AND U25644 ( .A(n383), .B(n26001), .Z(n26000) );
  XOR U25645 ( .A(p_input[4859]), .B(p_input[4827]), .Z(n26001) );
  XNOR U25646 ( .A(n25639), .B(n25996), .Z(n25998) );
  XOR U25647 ( .A(n26002), .B(n26003), .Z(n25639) );
  AND U25648 ( .A(n381), .B(n26004), .Z(n26003) );
  XOR U25649 ( .A(p_input[4795]), .B(p_input[4763]), .Z(n26004) );
  XOR U25650 ( .A(n26005), .B(n26006), .Z(n25996) );
  AND U25651 ( .A(n26007), .B(n26008), .Z(n26006) );
  XOR U25652 ( .A(n26005), .B(n25654), .Z(n26008) );
  XNOR U25653 ( .A(p_input[4826]), .B(n26009), .Z(n25654) );
  AND U25654 ( .A(n383), .B(n26010), .Z(n26009) );
  XOR U25655 ( .A(p_input[4858]), .B(p_input[4826]), .Z(n26010) );
  XNOR U25656 ( .A(n25651), .B(n26005), .Z(n26007) );
  XOR U25657 ( .A(n26011), .B(n26012), .Z(n25651) );
  AND U25658 ( .A(n381), .B(n26013), .Z(n26012) );
  XOR U25659 ( .A(p_input[4794]), .B(p_input[4762]), .Z(n26013) );
  XOR U25660 ( .A(n26014), .B(n26015), .Z(n26005) );
  AND U25661 ( .A(n26016), .B(n26017), .Z(n26015) );
  XOR U25662 ( .A(n26014), .B(n25666), .Z(n26017) );
  XNOR U25663 ( .A(p_input[4825]), .B(n26018), .Z(n25666) );
  AND U25664 ( .A(n383), .B(n26019), .Z(n26018) );
  XOR U25665 ( .A(p_input[4857]), .B(p_input[4825]), .Z(n26019) );
  XNOR U25666 ( .A(n25663), .B(n26014), .Z(n26016) );
  XOR U25667 ( .A(n26020), .B(n26021), .Z(n25663) );
  AND U25668 ( .A(n381), .B(n26022), .Z(n26021) );
  XOR U25669 ( .A(p_input[4793]), .B(p_input[4761]), .Z(n26022) );
  XOR U25670 ( .A(n26023), .B(n26024), .Z(n26014) );
  AND U25671 ( .A(n26025), .B(n26026), .Z(n26024) );
  XOR U25672 ( .A(n26023), .B(n25678), .Z(n26026) );
  XNOR U25673 ( .A(p_input[4824]), .B(n26027), .Z(n25678) );
  AND U25674 ( .A(n383), .B(n26028), .Z(n26027) );
  XOR U25675 ( .A(p_input[4856]), .B(p_input[4824]), .Z(n26028) );
  XNOR U25676 ( .A(n25675), .B(n26023), .Z(n26025) );
  XOR U25677 ( .A(n26029), .B(n26030), .Z(n25675) );
  AND U25678 ( .A(n381), .B(n26031), .Z(n26030) );
  XOR U25679 ( .A(p_input[4792]), .B(p_input[4760]), .Z(n26031) );
  XOR U25680 ( .A(n26032), .B(n26033), .Z(n26023) );
  AND U25681 ( .A(n26034), .B(n26035), .Z(n26033) );
  XOR U25682 ( .A(n26032), .B(n25690), .Z(n26035) );
  XNOR U25683 ( .A(p_input[4823]), .B(n26036), .Z(n25690) );
  AND U25684 ( .A(n383), .B(n26037), .Z(n26036) );
  XOR U25685 ( .A(p_input[4855]), .B(p_input[4823]), .Z(n26037) );
  XNOR U25686 ( .A(n25687), .B(n26032), .Z(n26034) );
  XOR U25687 ( .A(n26038), .B(n26039), .Z(n25687) );
  AND U25688 ( .A(n381), .B(n26040), .Z(n26039) );
  XOR U25689 ( .A(p_input[4791]), .B(p_input[4759]), .Z(n26040) );
  XOR U25690 ( .A(n26041), .B(n26042), .Z(n26032) );
  AND U25691 ( .A(n26043), .B(n26044), .Z(n26042) );
  XOR U25692 ( .A(n26041), .B(n25702), .Z(n26044) );
  XNOR U25693 ( .A(p_input[4822]), .B(n26045), .Z(n25702) );
  AND U25694 ( .A(n383), .B(n26046), .Z(n26045) );
  XOR U25695 ( .A(p_input[4854]), .B(p_input[4822]), .Z(n26046) );
  XNOR U25696 ( .A(n25699), .B(n26041), .Z(n26043) );
  XOR U25697 ( .A(n26047), .B(n26048), .Z(n25699) );
  AND U25698 ( .A(n381), .B(n26049), .Z(n26048) );
  XOR U25699 ( .A(p_input[4790]), .B(p_input[4758]), .Z(n26049) );
  XOR U25700 ( .A(n26050), .B(n26051), .Z(n26041) );
  AND U25701 ( .A(n26052), .B(n26053), .Z(n26051) );
  XOR U25702 ( .A(n26050), .B(n25714), .Z(n26053) );
  XNOR U25703 ( .A(p_input[4821]), .B(n26054), .Z(n25714) );
  AND U25704 ( .A(n383), .B(n26055), .Z(n26054) );
  XOR U25705 ( .A(p_input[4853]), .B(p_input[4821]), .Z(n26055) );
  XNOR U25706 ( .A(n25711), .B(n26050), .Z(n26052) );
  XOR U25707 ( .A(n26056), .B(n26057), .Z(n25711) );
  AND U25708 ( .A(n381), .B(n26058), .Z(n26057) );
  XOR U25709 ( .A(p_input[4789]), .B(p_input[4757]), .Z(n26058) );
  XOR U25710 ( .A(n26059), .B(n26060), .Z(n26050) );
  AND U25711 ( .A(n26061), .B(n26062), .Z(n26060) );
  XOR U25712 ( .A(n26059), .B(n25726), .Z(n26062) );
  XNOR U25713 ( .A(p_input[4820]), .B(n26063), .Z(n25726) );
  AND U25714 ( .A(n383), .B(n26064), .Z(n26063) );
  XOR U25715 ( .A(p_input[4852]), .B(p_input[4820]), .Z(n26064) );
  XNOR U25716 ( .A(n25723), .B(n26059), .Z(n26061) );
  XOR U25717 ( .A(n26065), .B(n26066), .Z(n25723) );
  AND U25718 ( .A(n381), .B(n26067), .Z(n26066) );
  XOR U25719 ( .A(p_input[4788]), .B(p_input[4756]), .Z(n26067) );
  XOR U25720 ( .A(n26068), .B(n26069), .Z(n26059) );
  AND U25721 ( .A(n26070), .B(n26071), .Z(n26069) );
  XOR U25722 ( .A(n26068), .B(n25738), .Z(n26071) );
  XNOR U25723 ( .A(p_input[4819]), .B(n26072), .Z(n25738) );
  AND U25724 ( .A(n383), .B(n26073), .Z(n26072) );
  XOR U25725 ( .A(p_input[4851]), .B(p_input[4819]), .Z(n26073) );
  XNOR U25726 ( .A(n25735), .B(n26068), .Z(n26070) );
  XOR U25727 ( .A(n26074), .B(n26075), .Z(n25735) );
  AND U25728 ( .A(n381), .B(n26076), .Z(n26075) );
  XOR U25729 ( .A(p_input[4787]), .B(p_input[4755]), .Z(n26076) );
  XOR U25730 ( .A(n26077), .B(n26078), .Z(n26068) );
  AND U25731 ( .A(n26079), .B(n26080), .Z(n26078) );
  XOR U25732 ( .A(n26077), .B(n25750), .Z(n26080) );
  XNOR U25733 ( .A(p_input[4818]), .B(n26081), .Z(n25750) );
  AND U25734 ( .A(n383), .B(n26082), .Z(n26081) );
  XOR U25735 ( .A(p_input[4850]), .B(p_input[4818]), .Z(n26082) );
  XNOR U25736 ( .A(n25747), .B(n26077), .Z(n26079) );
  XOR U25737 ( .A(n26083), .B(n26084), .Z(n25747) );
  AND U25738 ( .A(n381), .B(n26085), .Z(n26084) );
  XOR U25739 ( .A(p_input[4786]), .B(p_input[4754]), .Z(n26085) );
  XOR U25740 ( .A(n26086), .B(n26087), .Z(n26077) );
  AND U25741 ( .A(n26088), .B(n26089), .Z(n26087) );
  XOR U25742 ( .A(n26086), .B(n25762), .Z(n26089) );
  XNOR U25743 ( .A(p_input[4817]), .B(n26090), .Z(n25762) );
  AND U25744 ( .A(n383), .B(n26091), .Z(n26090) );
  XOR U25745 ( .A(p_input[4849]), .B(p_input[4817]), .Z(n26091) );
  XNOR U25746 ( .A(n25759), .B(n26086), .Z(n26088) );
  XOR U25747 ( .A(n26092), .B(n26093), .Z(n25759) );
  AND U25748 ( .A(n381), .B(n26094), .Z(n26093) );
  XOR U25749 ( .A(p_input[4785]), .B(p_input[4753]), .Z(n26094) );
  XOR U25750 ( .A(n26095), .B(n26096), .Z(n26086) );
  AND U25751 ( .A(n26097), .B(n26098), .Z(n26096) );
  XOR U25752 ( .A(n26095), .B(n25774), .Z(n26098) );
  XNOR U25753 ( .A(p_input[4816]), .B(n26099), .Z(n25774) );
  AND U25754 ( .A(n383), .B(n26100), .Z(n26099) );
  XOR U25755 ( .A(p_input[4848]), .B(p_input[4816]), .Z(n26100) );
  XNOR U25756 ( .A(n25771), .B(n26095), .Z(n26097) );
  XOR U25757 ( .A(n26101), .B(n26102), .Z(n25771) );
  AND U25758 ( .A(n381), .B(n26103), .Z(n26102) );
  XOR U25759 ( .A(p_input[4784]), .B(p_input[4752]), .Z(n26103) );
  XOR U25760 ( .A(n26104), .B(n26105), .Z(n26095) );
  AND U25761 ( .A(n26106), .B(n26107), .Z(n26105) );
  XOR U25762 ( .A(n26104), .B(n25786), .Z(n26107) );
  XNOR U25763 ( .A(p_input[4815]), .B(n26108), .Z(n25786) );
  AND U25764 ( .A(n383), .B(n26109), .Z(n26108) );
  XOR U25765 ( .A(p_input[4847]), .B(p_input[4815]), .Z(n26109) );
  XNOR U25766 ( .A(n25783), .B(n26104), .Z(n26106) );
  XOR U25767 ( .A(n26110), .B(n26111), .Z(n25783) );
  AND U25768 ( .A(n381), .B(n26112), .Z(n26111) );
  XOR U25769 ( .A(p_input[4783]), .B(p_input[4751]), .Z(n26112) );
  XOR U25770 ( .A(n26113), .B(n26114), .Z(n26104) );
  AND U25771 ( .A(n26115), .B(n26116), .Z(n26114) );
  XOR U25772 ( .A(n26113), .B(n25798), .Z(n26116) );
  XNOR U25773 ( .A(p_input[4814]), .B(n26117), .Z(n25798) );
  AND U25774 ( .A(n383), .B(n26118), .Z(n26117) );
  XOR U25775 ( .A(p_input[4846]), .B(p_input[4814]), .Z(n26118) );
  XNOR U25776 ( .A(n25795), .B(n26113), .Z(n26115) );
  XOR U25777 ( .A(n26119), .B(n26120), .Z(n25795) );
  AND U25778 ( .A(n381), .B(n26121), .Z(n26120) );
  XOR U25779 ( .A(p_input[4782]), .B(p_input[4750]), .Z(n26121) );
  XOR U25780 ( .A(n26122), .B(n26123), .Z(n26113) );
  AND U25781 ( .A(n26124), .B(n26125), .Z(n26123) );
  XOR U25782 ( .A(n26122), .B(n25810), .Z(n26125) );
  XNOR U25783 ( .A(p_input[4813]), .B(n26126), .Z(n25810) );
  AND U25784 ( .A(n383), .B(n26127), .Z(n26126) );
  XOR U25785 ( .A(p_input[4845]), .B(p_input[4813]), .Z(n26127) );
  XNOR U25786 ( .A(n25807), .B(n26122), .Z(n26124) );
  XOR U25787 ( .A(n26128), .B(n26129), .Z(n25807) );
  AND U25788 ( .A(n381), .B(n26130), .Z(n26129) );
  XOR U25789 ( .A(p_input[4781]), .B(p_input[4749]), .Z(n26130) );
  XOR U25790 ( .A(n26131), .B(n26132), .Z(n26122) );
  AND U25791 ( .A(n26133), .B(n26134), .Z(n26132) );
  XOR U25792 ( .A(n26131), .B(n25822), .Z(n26134) );
  XNOR U25793 ( .A(p_input[4812]), .B(n26135), .Z(n25822) );
  AND U25794 ( .A(n383), .B(n26136), .Z(n26135) );
  XOR U25795 ( .A(p_input[4844]), .B(p_input[4812]), .Z(n26136) );
  XNOR U25796 ( .A(n25819), .B(n26131), .Z(n26133) );
  XOR U25797 ( .A(n26137), .B(n26138), .Z(n25819) );
  AND U25798 ( .A(n381), .B(n26139), .Z(n26138) );
  XOR U25799 ( .A(p_input[4780]), .B(p_input[4748]), .Z(n26139) );
  XOR U25800 ( .A(n26140), .B(n26141), .Z(n26131) );
  AND U25801 ( .A(n26142), .B(n26143), .Z(n26141) );
  XOR U25802 ( .A(n26140), .B(n25834), .Z(n26143) );
  XNOR U25803 ( .A(p_input[4811]), .B(n26144), .Z(n25834) );
  AND U25804 ( .A(n383), .B(n26145), .Z(n26144) );
  XOR U25805 ( .A(p_input[4843]), .B(p_input[4811]), .Z(n26145) );
  XNOR U25806 ( .A(n25831), .B(n26140), .Z(n26142) );
  XOR U25807 ( .A(n26146), .B(n26147), .Z(n25831) );
  AND U25808 ( .A(n381), .B(n26148), .Z(n26147) );
  XOR U25809 ( .A(p_input[4779]), .B(p_input[4747]), .Z(n26148) );
  XOR U25810 ( .A(n26149), .B(n26150), .Z(n26140) );
  AND U25811 ( .A(n26151), .B(n26152), .Z(n26150) );
  XOR U25812 ( .A(n26149), .B(n25846), .Z(n26152) );
  XNOR U25813 ( .A(p_input[4810]), .B(n26153), .Z(n25846) );
  AND U25814 ( .A(n383), .B(n26154), .Z(n26153) );
  XOR U25815 ( .A(p_input[4842]), .B(p_input[4810]), .Z(n26154) );
  XNOR U25816 ( .A(n25843), .B(n26149), .Z(n26151) );
  XOR U25817 ( .A(n26155), .B(n26156), .Z(n25843) );
  AND U25818 ( .A(n381), .B(n26157), .Z(n26156) );
  XOR U25819 ( .A(p_input[4778]), .B(p_input[4746]), .Z(n26157) );
  XOR U25820 ( .A(n26158), .B(n26159), .Z(n26149) );
  AND U25821 ( .A(n26160), .B(n26161), .Z(n26159) );
  XOR U25822 ( .A(n26158), .B(n25858), .Z(n26161) );
  XNOR U25823 ( .A(p_input[4809]), .B(n26162), .Z(n25858) );
  AND U25824 ( .A(n383), .B(n26163), .Z(n26162) );
  XOR U25825 ( .A(p_input[4841]), .B(p_input[4809]), .Z(n26163) );
  XNOR U25826 ( .A(n25855), .B(n26158), .Z(n26160) );
  XOR U25827 ( .A(n26164), .B(n26165), .Z(n25855) );
  AND U25828 ( .A(n381), .B(n26166), .Z(n26165) );
  XOR U25829 ( .A(p_input[4777]), .B(p_input[4745]), .Z(n26166) );
  XOR U25830 ( .A(n26167), .B(n26168), .Z(n26158) );
  AND U25831 ( .A(n26169), .B(n26170), .Z(n26168) );
  XOR U25832 ( .A(n26167), .B(n25870), .Z(n26170) );
  XNOR U25833 ( .A(p_input[4808]), .B(n26171), .Z(n25870) );
  AND U25834 ( .A(n383), .B(n26172), .Z(n26171) );
  XOR U25835 ( .A(p_input[4840]), .B(p_input[4808]), .Z(n26172) );
  XNOR U25836 ( .A(n25867), .B(n26167), .Z(n26169) );
  XOR U25837 ( .A(n26173), .B(n26174), .Z(n25867) );
  AND U25838 ( .A(n381), .B(n26175), .Z(n26174) );
  XOR U25839 ( .A(p_input[4776]), .B(p_input[4744]), .Z(n26175) );
  XOR U25840 ( .A(n26176), .B(n26177), .Z(n26167) );
  AND U25841 ( .A(n26178), .B(n26179), .Z(n26177) );
  XOR U25842 ( .A(n26176), .B(n25882), .Z(n26179) );
  XNOR U25843 ( .A(p_input[4807]), .B(n26180), .Z(n25882) );
  AND U25844 ( .A(n383), .B(n26181), .Z(n26180) );
  XOR U25845 ( .A(p_input[4839]), .B(p_input[4807]), .Z(n26181) );
  XNOR U25846 ( .A(n25879), .B(n26176), .Z(n26178) );
  XOR U25847 ( .A(n26182), .B(n26183), .Z(n25879) );
  AND U25848 ( .A(n381), .B(n26184), .Z(n26183) );
  XOR U25849 ( .A(p_input[4775]), .B(p_input[4743]), .Z(n26184) );
  XOR U25850 ( .A(n26185), .B(n26186), .Z(n26176) );
  AND U25851 ( .A(n26187), .B(n26188), .Z(n26186) );
  XOR U25852 ( .A(n26185), .B(n25894), .Z(n26188) );
  XNOR U25853 ( .A(p_input[4806]), .B(n26189), .Z(n25894) );
  AND U25854 ( .A(n383), .B(n26190), .Z(n26189) );
  XOR U25855 ( .A(p_input[4838]), .B(p_input[4806]), .Z(n26190) );
  XNOR U25856 ( .A(n25891), .B(n26185), .Z(n26187) );
  XOR U25857 ( .A(n26191), .B(n26192), .Z(n25891) );
  AND U25858 ( .A(n381), .B(n26193), .Z(n26192) );
  XOR U25859 ( .A(p_input[4774]), .B(p_input[4742]), .Z(n26193) );
  XOR U25860 ( .A(n26194), .B(n26195), .Z(n26185) );
  AND U25861 ( .A(n26196), .B(n26197), .Z(n26195) );
  XOR U25862 ( .A(n26194), .B(n25906), .Z(n26197) );
  XNOR U25863 ( .A(p_input[4805]), .B(n26198), .Z(n25906) );
  AND U25864 ( .A(n383), .B(n26199), .Z(n26198) );
  XOR U25865 ( .A(p_input[4837]), .B(p_input[4805]), .Z(n26199) );
  XNOR U25866 ( .A(n25903), .B(n26194), .Z(n26196) );
  XOR U25867 ( .A(n26200), .B(n26201), .Z(n25903) );
  AND U25868 ( .A(n381), .B(n26202), .Z(n26201) );
  XOR U25869 ( .A(p_input[4773]), .B(p_input[4741]), .Z(n26202) );
  XOR U25870 ( .A(n26203), .B(n26204), .Z(n26194) );
  AND U25871 ( .A(n26205), .B(n26206), .Z(n26204) );
  XOR U25872 ( .A(n26203), .B(n25918), .Z(n26206) );
  XNOR U25873 ( .A(p_input[4804]), .B(n26207), .Z(n25918) );
  AND U25874 ( .A(n383), .B(n26208), .Z(n26207) );
  XOR U25875 ( .A(p_input[4836]), .B(p_input[4804]), .Z(n26208) );
  XNOR U25876 ( .A(n25915), .B(n26203), .Z(n26205) );
  XOR U25877 ( .A(n26209), .B(n26210), .Z(n25915) );
  AND U25878 ( .A(n381), .B(n26211), .Z(n26210) );
  XOR U25879 ( .A(p_input[4772]), .B(p_input[4740]), .Z(n26211) );
  XOR U25880 ( .A(n26212), .B(n26213), .Z(n26203) );
  AND U25881 ( .A(n26214), .B(n26215), .Z(n26213) );
  XOR U25882 ( .A(n26212), .B(n25930), .Z(n26215) );
  XNOR U25883 ( .A(p_input[4803]), .B(n26216), .Z(n25930) );
  AND U25884 ( .A(n383), .B(n26217), .Z(n26216) );
  XOR U25885 ( .A(p_input[4835]), .B(p_input[4803]), .Z(n26217) );
  XNOR U25886 ( .A(n25927), .B(n26212), .Z(n26214) );
  XOR U25887 ( .A(n26218), .B(n26219), .Z(n25927) );
  AND U25888 ( .A(n381), .B(n26220), .Z(n26219) );
  XOR U25889 ( .A(p_input[4771]), .B(p_input[4739]), .Z(n26220) );
  XOR U25890 ( .A(n26221), .B(n26222), .Z(n26212) );
  AND U25891 ( .A(n26223), .B(n26224), .Z(n26222) );
  XOR U25892 ( .A(n26221), .B(n25942), .Z(n26224) );
  XNOR U25893 ( .A(p_input[4802]), .B(n26225), .Z(n25942) );
  AND U25894 ( .A(n383), .B(n26226), .Z(n26225) );
  XOR U25895 ( .A(p_input[4834]), .B(p_input[4802]), .Z(n26226) );
  XNOR U25896 ( .A(n25939), .B(n26221), .Z(n26223) );
  XOR U25897 ( .A(n26227), .B(n26228), .Z(n25939) );
  AND U25898 ( .A(n381), .B(n26229), .Z(n26228) );
  XOR U25899 ( .A(p_input[4770]), .B(p_input[4738]), .Z(n26229) );
  XOR U25900 ( .A(n26230), .B(n26231), .Z(n26221) );
  AND U25901 ( .A(n26232), .B(n26233), .Z(n26231) );
  XNOR U25902 ( .A(n26234), .B(n25955), .Z(n26233) );
  XNOR U25903 ( .A(p_input[4801]), .B(n26235), .Z(n25955) );
  AND U25904 ( .A(n383), .B(n26236), .Z(n26235) );
  XNOR U25905 ( .A(p_input[4833]), .B(n26237), .Z(n26236) );
  IV U25906 ( .A(p_input[4801]), .Z(n26237) );
  XNOR U25907 ( .A(n25952), .B(n26230), .Z(n26232) );
  XNOR U25908 ( .A(p_input[4737]), .B(n26238), .Z(n25952) );
  AND U25909 ( .A(n381), .B(n26239), .Z(n26238) );
  XOR U25910 ( .A(p_input[4769]), .B(p_input[4737]), .Z(n26239) );
  IV U25911 ( .A(n26234), .Z(n26230) );
  AND U25912 ( .A(n25960), .B(n25963), .Z(n26234) );
  XOR U25913 ( .A(p_input[4800]), .B(n26240), .Z(n25963) );
  AND U25914 ( .A(n383), .B(n26241), .Z(n26240) );
  XOR U25915 ( .A(p_input[4832]), .B(p_input[4800]), .Z(n26241) );
  XOR U25916 ( .A(n26242), .B(n26243), .Z(n383) );
  AND U25917 ( .A(n26244), .B(n26245), .Z(n26243) );
  XNOR U25918 ( .A(p_input[4863]), .B(n26242), .Z(n26245) );
  XOR U25919 ( .A(n26242), .B(p_input[4831]), .Z(n26244) );
  XOR U25920 ( .A(n26246), .B(n26247), .Z(n26242) );
  AND U25921 ( .A(n26248), .B(n26249), .Z(n26247) );
  XNOR U25922 ( .A(p_input[4862]), .B(n26246), .Z(n26249) );
  XOR U25923 ( .A(n26246), .B(p_input[4830]), .Z(n26248) );
  XOR U25924 ( .A(n26250), .B(n26251), .Z(n26246) );
  AND U25925 ( .A(n26252), .B(n26253), .Z(n26251) );
  XNOR U25926 ( .A(p_input[4861]), .B(n26250), .Z(n26253) );
  XOR U25927 ( .A(n26250), .B(p_input[4829]), .Z(n26252) );
  XOR U25928 ( .A(n26254), .B(n26255), .Z(n26250) );
  AND U25929 ( .A(n26256), .B(n26257), .Z(n26255) );
  XNOR U25930 ( .A(p_input[4860]), .B(n26254), .Z(n26257) );
  XOR U25931 ( .A(n26254), .B(p_input[4828]), .Z(n26256) );
  XOR U25932 ( .A(n26258), .B(n26259), .Z(n26254) );
  AND U25933 ( .A(n26260), .B(n26261), .Z(n26259) );
  XNOR U25934 ( .A(p_input[4859]), .B(n26258), .Z(n26261) );
  XOR U25935 ( .A(n26258), .B(p_input[4827]), .Z(n26260) );
  XOR U25936 ( .A(n26262), .B(n26263), .Z(n26258) );
  AND U25937 ( .A(n26264), .B(n26265), .Z(n26263) );
  XNOR U25938 ( .A(p_input[4858]), .B(n26262), .Z(n26265) );
  XOR U25939 ( .A(n26262), .B(p_input[4826]), .Z(n26264) );
  XOR U25940 ( .A(n26266), .B(n26267), .Z(n26262) );
  AND U25941 ( .A(n26268), .B(n26269), .Z(n26267) );
  XNOR U25942 ( .A(p_input[4857]), .B(n26266), .Z(n26269) );
  XOR U25943 ( .A(n26266), .B(p_input[4825]), .Z(n26268) );
  XOR U25944 ( .A(n26270), .B(n26271), .Z(n26266) );
  AND U25945 ( .A(n26272), .B(n26273), .Z(n26271) );
  XNOR U25946 ( .A(p_input[4856]), .B(n26270), .Z(n26273) );
  XOR U25947 ( .A(n26270), .B(p_input[4824]), .Z(n26272) );
  XOR U25948 ( .A(n26274), .B(n26275), .Z(n26270) );
  AND U25949 ( .A(n26276), .B(n26277), .Z(n26275) );
  XNOR U25950 ( .A(p_input[4855]), .B(n26274), .Z(n26277) );
  XOR U25951 ( .A(n26274), .B(p_input[4823]), .Z(n26276) );
  XOR U25952 ( .A(n26278), .B(n26279), .Z(n26274) );
  AND U25953 ( .A(n26280), .B(n26281), .Z(n26279) );
  XNOR U25954 ( .A(p_input[4854]), .B(n26278), .Z(n26281) );
  XOR U25955 ( .A(n26278), .B(p_input[4822]), .Z(n26280) );
  XOR U25956 ( .A(n26282), .B(n26283), .Z(n26278) );
  AND U25957 ( .A(n26284), .B(n26285), .Z(n26283) );
  XNOR U25958 ( .A(p_input[4853]), .B(n26282), .Z(n26285) );
  XOR U25959 ( .A(n26282), .B(p_input[4821]), .Z(n26284) );
  XOR U25960 ( .A(n26286), .B(n26287), .Z(n26282) );
  AND U25961 ( .A(n26288), .B(n26289), .Z(n26287) );
  XNOR U25962 ( .A(p_input[4852]), .B(n26286), .Z(n26289) );
  XOR U25963 ( .A(n26286), .B(p_input[4820]), .Z(n26288) );
  XOR U25964 ( .A(n26290), .B(n26291), .Z(n26286) );
  AND U25965 ( .A(n26292), .B(n26293), .Z(n26291) );
  XNOR U25966 ( .A(p_input[4851]), .B(n26290), .Z(n26293) );
  XOR U25967 ( .A(n26290), .B(p_input[4819]), .Z(n26292) );
  XOR U25968 ( .A(n26294), .B(n26295), .Z(n26290) );
  AND U25969 ( .A(n26296), .B(n26297), .Z(n26295) );
  XNOR U25970 ( .A(p_input[4850]), .B(n26294), .Z(n26297) );
  XOR U25971 ( .A(n26294), .B(p_input[4818]), .Z(n26296) );
  XOR U25972 ( .A(n26298), .B(n26299), .Z(n26294) );
  AND U25973 ( .A(n26300), .B(n26301), .Z(n26299) );
  XNOR U25974 ( .A(p_input[4849]), .B(n26298), .Z(n26301) );
  XOR U25975 ( .A(n26298), .B(p_input[4817]), .Z(n26300) );
  XOR U25976 ( .A(n26302), .B(n26303), .Z(n26298) );
  AND U25977 ( .A(n26304), .B(n26305), .Z(n26303) );
  XNOR U25978 ( .A(p_input[4848]), .B(n26302), .Z(n26305) );
  XOR U25979 ( .A(n26302), .B(p_input[4816]), .Z(n26304) );
  XOR U25980 ( .A(n26306), .B(n26307), .Z(n26302) );
  AND U25981 ( .A(n26308), .B(n26309), .Z(n26307) );
  XNOR U25982 ( .A(p_input[4847]), .B(n26306), .Z(n26309) );
  XOR U25983 ( .A(n26306), .B(p_input[4815]), .Z(n26308) );
  XOR U25984 ( .A(n26310), .B(n26311), .Z(n26306) );
  AND U25985 ( .A(n26312), .B(n26313), .Z(n26311) );
  XNOR U25986 ( .A(p_input[4846]), .B(n26310), .Z(n26313) );
  XOR U25987 ( .A(n26310), .B(p_input[4814]), .Z(n26312) );
  XOR U25988 ( .A(n26314), .B(n26315), .Z(n26310) );
  AND U25989 ( .A(n26316), .B(n26317), .Z(n26315) );
  XNOR U25990 ( .A(p_input[4845]), .B(n26314), .Z(n26317) );
  XOR U25991 ( .A(n26314), .B(p_input[4813]), .Z(n26316) );
  XOR U25992 ( .A(n26318), .B(n26319), .Z(n26314) );
  AND U25993 ( .A(n26320), .B(n26321), .Z(n26319) );
  XNOR U25994 ( .A(p_input[4844]), .B(n26318), .Z(n26321) );
  XOR U25995 ( .A(n26318), .B(p_input[4812]), .Z(n26320) );
  XOR U25996 ( .A(n26322), .B(n26323), .Z(n26318) );
  AND U25997 ( .A(n26324), .B(n26325), .Z(n26323) );
  XNOR U25998 ( .A(p_input[4843]), .B(n26322), .Z(n26325) );
  XOR U25999 ( .A(n26322), .B(p_input[4811]), .Z(n26324) );
  XOR U26000 ( .A(n26326), .B(n26327), .Z(n26322) );
  AND U26001 ( .A(n26328), .B(n26329), .Z(n26327) );
  XNOR U26002 ( .A(p_input[4842]), .B(n26326), .Z(n26329) );
  XOR U26003 ( .A(n26326), .B(p_input[4810]), .Z(n26328) );
  XOR U26004 ( .A(n26330), .B(n26331), .Z(n26326) );
  AND U26005 ( .A(n26332), .B(n26333), .Z(n26331) );
  XNOR U26006 ( .A(p_input[4841]), .B(n26330), .Z(n26333) );
  XOR U26007 ( .A(n26330), .B(p_input[4809]), .Z(n26332) );
  XOR U26008 ( .A(n26334), .B(n26335), .Z(n26330) );
  AND U26009 ( .A(n26336), .B(n26337), .Z(n26335) );
  XNOR U26010 ( .A(p_input[4840]), .B(n26334), .Z(n26337) );
  XOR U26011 ( .A(n26334), .B(p_input[4808]), .Z(n26336) );
  XOR U26012 ( .A(n26338), .B(n26339), .Z(n26334) );
  AND U26013 ( .A(n26340), .B(n26341), .Z(n26339) );
  XNOR U26014 ( .A(p_input[4839]), .B(n26338), .Z(n26341) );
  XOR U26015 ( .A(n26338), .B(p_input[4807]), .Z(n26340) );
  XOR U26016 ( .A(n26342), .B(n26343), .Z(n26338) );
  AND U26017 ( .A(n26344), .B(n26345), .Z(n26343) );
  XNOR U26018 ( .A(p_input[4838]), .B(n26342), .Z(n26345) );
  XOR U26019 ( .A(n26342), .B(p_input[4806]), .Z(n26344) );
  XOR U26020 ( .A(n26346), .B(n26347), .Z(n26342) );
  AND U26021 ( .A(n26348), .B(n26349), .Z(n26347) );
  XNOR U26022 ( .A(p_input[4837]), .B(n26346), .Z(n26349) );
  XOR U26023 ( .A(n26346), .B(p_input[4805]), .Z(n26348) );
  XOR U26024 ( .A(n26350), .B(n26351), .Z(n26346) );
  AND U26025 ( .A(n26352), .B(n26353), .Z(n26351) );
  XNOR U26026 ( .A(p_input[4836]), .B(n26350), .Z(n26353) );
  XOR U26027 ( .A(n26350), .B(p_input[4804]), .Z(n26352) );
  XOR U26028 ( .A(n26354), .B(n26355), .Z(n26350) );
  AND U26029 ( .A(n26356), .B(n26357), .Z(n26355) );
  XNOR U26030 ( .A(p_input[4835]), .B(n26354), .Z(n26357) );
  XOR U26031 ( .A(n26354), .B(p_input[4803]), .Z(n26356) );
  XOR U26032 ( .A(n26358), .B(n26359), .Z(n26354) );
  AND U26033 ( .A(n26360), .B(n26361), .Z(n26359) );
  XNOR U26034 ( .A(p_input[4834]), .B(n26358), .Z(n26361) );
  XOR U26035 ( .A(n26358), .B(p_input[4802]), .Z(n26360) );
  XNOR U26036 ( .A(n26362), .B(n26363), .Z(n26358) );
  AND U26037 ( .A(n26364), .B(n26365), .Z(n26363) );
  XOR U26038 ( .A(p_input[4833]), .B(n26362), .Z(n26365) );
  XNOR U26039 ( .A(p_input[4801]), .B(n26362), .Z(n26364) );
  AND U26040 ( .A(p_input[4832]), .B(n26366), .Z(n26362) );
  IV U26041 ( .A(p_input[4800]), .Z(n26366) );
  XNOR U26042 ( .A(p_input[4736]), .B(n26367), .Z(n25960) );
  AND U26043 ( .A(n381), .B(n26368), .Z(n26367) );
  XOR U26044 ( .A(p_input[4768]), .B(p_input[4736]), .Z(n26368) );
  XOR U26045 ( .A(n26369), .B(n26370), .Z(n381) );
  AND U26046 ( .A(n26371), .B(n26372), .Z(n26370) );
  XNOR U26047 ( .A(p_input[4799]), .B(n26369), .Z(n26372) );
  XOR U26048 ( .A(n26369), .B(p_input[4767]), .Z(n26371) );
  XOR U26049 ( .A(n26373), .B(n26374), .Z(n26369) );
  AND U26050 ( .A(n26375), .B(n26376), .Z(n26374) );
  XNOR U26051 ( .A(p_input[4798]), .B(n26373), .Z(n26376) );
  XNOR U26052 ( .A(n26373), .B(n25975), .Z(n26375) );
  IV U26053 ( .A(p_input[4766]), .Z(n25975) );
  XOR U26054 ( .A(n26377), .B(n26378), .Z(n26373) );
  AND U26055 ( .A(n26379), .B(n26380), .Z(n26378) );
  XNOR U26056 ( .A(p_input[4797]), .B(n26377), .Z(n26380) );
  XNOR U26057 ( .A(n26377), .B(n25984), .Z(n26379) );
  IV U26058 ( .A(p_input[4765]), .Z(n25984) );
  XOR U26059 ( .A(n26381), .B(n26382), .Z(n26377) );
  AND U26060 ( .A(n26383), .B(n26384), .Z(n26382) );
  XNOR U26061 ( .A(p_input[4796]), .B(n26381), .Z(n26384) );
  XNOR U26062 ( .A(n26381), .B(n25993), .Z(n26383) );
  IV U26063 ( .A(p_input[4764]), .Z(n25993) );
  XOR U26064 ( .A(n26385), .B(n26386), .Z(n26381) );
  AND U26065 ( .A(n26387), .B(n26388), .Z(n26386) );
  XNOR U26066 ( .A(p_input[4795]), .B(n26385), .Z(n26388) );
  XNOR U26067 ( .A(n26385), .B(n26002), .Z(n26387) );
  IV U26068 ( .A(p_input[4763]), .Z(n26002) );
  XOR U26069 ( .A(n26389), .B(n26390), .Z(n26385) );
  AND U26070 ( .A(n26391), .B(n26392), .Z(n26390) );
  XNOR U26071 ( .A(p_input[4794]), .B(n26389), .Z(n26392) );
  XNOR U26072 ( .A(n26389), .B(n26011), .Z(n26391) );
  IV U26073 ( .A(p_input[4762]), .Z(n26011) );
  XOR U26074 ( .A(n26393), .B(n26394), .Z(n26389) );
  AND U26075 ( .A(n26395), .B(n26396), .Z(n26394) );
  XNOR U26076 ( .A(p_input[4793]), .B(n26393), .Z(n26396) );
  XNOR U26077 ( .A(n26393), .B(n26020), .Z(n26395) );
  IV U26078 ( .A(p_input[4761]), .Z(n26020) );
  XOR U26079 ( .A(n26397), .B(n26398), .Z(n26393) );
  AND U26080 ( .A(n26399), .B(n26400), .Z(n26398) );
  XNOR U26081 ( .A(p_input[4792]), .B(n26397), .Z(n26400) );
  XNOR U26082 ( .A(n26397), .B(n26029), .Z(n26399) );
  IV U26083 ( .A(p_input[4760]), .Z(n26029) );
  XOR U26084 ( .A(n26401), .B(n26402), .Z(n26397) );
  AND U26085 ( .A(n26403), .B(n26404), .Z(n26402) );
  XNOR U26086 ( .A(p_input[4791]), .B(n26401), .Z(n26404) );
  XNOR U26087 ( .A(n26401), .B(n26038), .Z(n26403) );
  IV U26088 ( .A(p_input[4759]), .Z(n26038) );
  XOR U26089 ( .A(n26405), .B(n26406), .Z(n26401) );
  AND U26090 ( .A(n26407), .B(n26408), .Z(n26406) );
  XNOR U26091 ( .A(p_input[4790]), .B(n26405), .Z(n26408) );
  XNOR U26092 ( .A(n26405), .B(n26047), .Z(n26407) );
  IV U26093 ( .A(p_input[4758]), .Z(n26047) );
  XOR U26094 ( .A(n26409), .B(n26410), .Z(n26405) );
  AND U26095 ( .A(n26411), .B(n26412), .Z(n26410) );
  XNOR U26096 ( .A(p_input[4789]), .B(n26409), .Z(n26412) );
  XNOR U26097 ( .A(n26409), .B(n26056), .Z(n26411) );
  IV U26098 ( .A(p_input[4757]), .Z(n26056) );
  XOR U26099 ( .A(n26413), .B(n26414), .Z(n26409) );
  AND U26100 ( .A(n26415), .B(n26416), .Z(n26414) );
  XNOR U26101 ( .A(p_input[4788]), .B(n26413), .Z(n26416) );
  XNOR U26102 ( .A(n26413), .B(n26065), .Z(n26415) );
  IV U26103 ( .A(p_input[4756]), .Z(n26065) );
  XOR U26104 ( .A(n26417), .B(n26418), .Z(n26413) );
  AND U26105 ( .A(n26419), .B(n26420), .Z(n26418) );
  XNOR U26106 ( .A(p_input[4787]), .B(n26417), .Z(n26420) );
  XNOR U26107 ( .A(n26417), .B(n26074), .Z(n26419) );
  IV U26108 ( .A(p_input[4755]), .Z(n26074) );
  XOR U26109 ( .A(n26421), .B(n26422), .Z(n26417) );
  AND U26110 ( .A(n26423), .B(n26424), .Z(n26422) );
  XNOR U26111 ( .A(p_input[4786]), .B(n26421), .Z(n26424) );
  XNOR U26112 ( .A(n26421), .B(n26083), .Z(n26423) );
  IV U26113 ( .A(p_input[4754]), .Z(n26083) );
  XOR U26114 ( .A(n26425), .B(n26426), .Z(n26421) );
  AND U26115 ( .A(n26427), .B(n26428), .Z(n26426) );
  XNOR U26116 ( .A(p_input[4785]), .B(n26425), .Z(n26428) );
  XNOR U26117 ( .A(n26425), .B(n26092), .Z(n26427) );
  IV U26118 ( .A(p_input[4753]), .Z(n26092) );
  XOR U26119 ( .A(n26429), .B(n26430), .Z(n26425) );
  AND U26120 ( .A(n26431), .B(n26432), .Z(n26430) );
  XNOR U26121 ( .A(p_input[4784]), .B(n26429), .Z(n26432) );
  XNOR U26122 ( .A(n26429), .B(n26101), .Z(n26431) );
  IV U26123 ( .A(p_input[4752]), .Z(n26101) );
  XOR U26124 ( .A(n26433), .B(n26434), .Z(n26429) );
  AND U26125 ( .A(n26435), .B(n26436), .Z(n26434) );
  XNOR U26126 ( .A(p_input[4783]), .B(n26433), .Z(n26436) );
  XNOR U26127 ( .A(n26433), .B(n26110), .Z(n26435) );
  IV U26128 ( .A(p_input[4751]), .Z(n26110) );
  XOR U26129 ( .A(n26437), .B(n26438), .Z(n26433) );
  AND U26130 ( .A(n26439), .B(n26440), .Z(n26438) );
  XNOR U26131 ( .A(p_input[4782]), .B(n26437), .Z(n26440) );
  XNOR U26132 ( .A(n26437), .B(n26119), .Z(n26439) );
  IV U26133 ( .A(p_input[4750]), .Z(n26119) );
  XOR U26134 ( .A(n26441), .B(n26442), .Z(n26437) );
  AND U26135 ( .A(n26443), .B(n26444), .Z(n26442) );
  XNOR U26136 ( .A(p_input[4781]), .B(n26441), .Z(n26444) );
  XNOR U26137 ( .A(n26441), .B(n26128), .Z(n26443) );
  IV U26138 ( .A(p_input[4749]), .Z(n26128) );
  XOR U26139 ( .A(n26445), .B(n26446), .Z(n26441) );
  AND U26140 ( .A(n26447), .B(n26448), .Z(n26446) );
  XNOR U26141 ( .A(p_input[4780]), .B(n26445), .Z(n26448) );
  XNOR U26142 ( .A(n26445), .B(n26137), .Z(n26447) );
  IV U26143 ( .A(p_input[4748]), .Z(n26137) );
  XOR U26144 ( .A(n26449), .B(n26450), .Z(n26445) );
  AND U26145 ( .A(n26451), .B(n26452), .Z(n26450) );
  XNOR U26146 ( .A(p_input[4779]), .B(n26449), .Z(n26452) );
  XNOR U26147 ( .A(n26449), .B(n26146), .Z(n26451) );
  IV U26148 ( .A(p_input[4747]), .Z(n26146) );
  XOR U26149 ( .A(n26453), .B(n26454), .Z(n26449) );
  AND U26150 ( .A(n26455), .B(n26456), .Z(n26454) );
  XNOR U26151 ( .A(p_input[4778]), .B(n26453), .Z(n26456) );
  XNOR U26152 ( .A(n26453), .B(n26155), .Z(n26455) );
  IV U26153 ( .A(p_input[4746]), .Z(n26155) );
  XOR U26154 ( .A(n26457), .B(n26458), .Z(n26453) );
  AND U26155 ( .A(n26459), .B(n26460), .Z(n26458) );
  XNOR U26156 ( .A(p_input[4777]), .B(n26457), .Z(n26460) );
  XNOR U26157 ( .A(n26457), .B(n26164), .Z(n26459) );
  IV U26158 ( .A(p_input[4745]), .Z(n26164) );
  XOR U26159 ( .A(n26461), .B(n26462), .Z(n26457) );
  AND U26160 ( .A(n26463), .B(n26464), .Z(n26462) );
  XNOR U26161 ( .A(p_input[4776]), .B(n26461), .Z(n26464) );
  XNOR U26162 ( .A(n26461), .B(n26173), .Z(n26463) );
  IV U26163 ( .A(p_input[4744]), .Z(n26173) );
  XOR U26164 ( .A(n26465), .B(n26466), .Z(n26461) );
  AND U26165 ( .A(n26467), .B(n26468), .Z(n26466) );
  XNOR U26166 ( .A(p_input[4775]), .B(n26465), .Z(n26468) );
  XNOR U26167 ( .A(n26465), .B(n26182), .Z(n26467) );
  IV U26168 ( .A(p_input[4743]), .Z(n26182) );
  XOR U26169 ( .A(n26469), .B(n26470), .Z(n26465) );
  AND U26170 ( .A(n26471), .B(n26472), .Z(n26470) );
  XNOR U26171 ( .A(p_input[4774]), .B(n26469), .Z(n26472) );
  XNOR U26172 ( .A(n26469), .B(n26191), .Z(n26471) );
  IV U26173 ( .A(p_input[4742]), .Z(n26191) );
  XOR U26174 ( .A(n26473), .B(n26474), .Z(n26469) );
  AND U26175 ( .A(n26475), .B(n26476), .Z(n26474) );
  XNOR U26176 ( .A(p_input[4773]), .B(n26473), .Z(n26476) );
  XNOR U26177 ( .A(n26473), .B(n26200), .Z(n26475) );
  IV U26178 ( .A(p_input[4741]), .Z(n26200) );
  XOR U26179 ( .A(n26477), .B(n26478), .Z(n26473) );
  AND U26180 ( .A(n26479), .B(n26480), .Z(n26478) );
  XNOR U26181 ( .A(p_input[4772]), .B(n26477), .Z(n26480) );
  XNOR U26182 ( .A(n26477), .B(n26209), .Z(n26479) );
  IV U26183 ( .A(p_input[4740]), .Z(n26209) );
  XOR U26184 ( .A(n26481), .B(n26482), .Z(n26477) );
  AND U26185 ( .A(n26483), .B(n26484), .Z(n26482) );
  XNOR U26186 ( .A(p_input[4771]), .B(n26481), .Z(n26484) );
  XNOR U26187 ( .A(n26481), .B(n26218), .Z(n26483) );
  IV U26188 ( .A(p_input[4739]), .Z(n26218) );
  XOR U26189 ( .A(n26485), .B(n26486), .Z(n26481) );
  AND U26190 ( .A(n26487), .B(n26488), .Z(n26486) );
  XNOR U26191 ( .A(p_input[4770]), .B(n26485), .Z(n26488) );
  XNOR U26192 ( .A(n26485), .B(n26227), .Z(n26487) );
  IV U26193 ( .A(p_input[4738]), .Z(n26227) );
  XNOR U26194 ( .A(n26489), .B(n26490), .Z(n26485) );
  AND U26195 ( .A(n26491), .B(n26492), .Z(n26490) );
  XOR U26196 ( .A(p_input[4769]), .B(n26489), .Z(n26492) );
  XNOR U26197 ( .A(p_input[4737]), .B(n26489), .Z(n26491) );
  AND U26198 ( .A(p_input[4768]), .B(n26493), .Z(n26489) );
  IV U26199 ( .A(p_input[4736]), .Z(n26493) );
  XOR U26200 ( .A(n26494), .B(n26495), .Z(n25583) );
  AND U26201 ( .A(n528), .B(n26496), .Z(n26495) );
  XNOR U26202 ( .A(n26497), .B(n26494), .Z(n26496) );
  XOR U26203 ( .A(n26498), .B(n26499), .Z(n528) );
  AND U26204 ( .A(n26500), .B(n26501), .Z(n26499) );
  XNOR U26205 ( .A(n25598), .B(n26498), .Z(n26501) );
  AND U26206 ( .A(p_input[4735]), .B(p_input[4703]), .Z(n25598) );
  XNOR U26207 ( .A(n26498), .B(n25595), .Z(n26500) );
  IV U26208 ( .A(n26502), .Z(n25595) );
  AND U26209 ( .A(p_input[4639]), .B(p_input[4671]), .Z(n26502) );
  XOR U26210 ( .A(n26503), .B(n26504), .Z(n26498) );
  AND U26211 ( .A(n26505), .B(n26506), .Z(n26504) );
  XOR U26212 ( .A(n26503), .B(n25610), .Z(n26506) );
  XNOR U26213 ( .A(p_input[4702]), .B(n26507), .Z(n25610) );
  AND U26214 ( .A(n387), .B(n26508), .Z(n26507) );
  XOR U26215 ( .A(p_input[4734]), .B(p_input[4702]), .Z(n26508) );
  XNOR U26216 ( .A(n25607), .B(n26503), .Z(n26505) );
  XOR U26217 ( .A(n26509), .B(n26510), .Z(n25607) );
  AND U26218 ( .A(n384), .B(n26511), .Z(n26510) );
  XOR U26219 ( .A(p_input[4670]), .B(p_input[4638]), .Z(n26511) );
  XOR U26220 ( .A(n26512), .B(n26513), .Z(n26503) );
  AND U26221 ( .A(n26514), .B(n26515), .Z(n26513) );
  XOR U26222 ( .A(n26512), .B(n25622), .Z(n26515) );
  XNOR U26223 ( .A(p_input[4701]), .B(n26516), .Z(n25622) );
  AND U26224 ( .A(n387), .B(n26517), .Z(n26516) );
  XOR U26225 ( .A(p_input[4733]), .B(p_input[4701]), .Z(n26517) );
  XNOR U26226 ( .A(n25619), .B(n26512), .Z(n26514) );
  XOR U26227 ( .A(n26518), .B(n26519), .Z(n25619) );
  AND U26228 ( .A(n384), .B(n26520), .Z(n26519) );
  XOR U26229 ( .A(p_input[4669]), .B(p_input[4637]), .Z(n26520) );
  XOR U26230 ( .A(n26521), .B(n26522), .Z(n26512) );
  AND U26231 ( .A(n26523), .B(n26524), .Z(n26522) );
  XOR U26232 ( .A(n26521), .B(n25634), .Z(n26524) );
  XNOR U26233 ( .A(p_input[4700]), .B(n26525), .Z(n25634) );
  AND U26234 ( .A(n387), .B(n26526), .Z(n26525) );
  XOR U26235 ( .A(p_input[4732]), .B(p_input[4700]), .Z(n26526) );
  XNOR U26236 ( .A(n25631), .B(n26521), .Z(n26523) );
  XOR U26237 ( .A(n26527), .B(n26528), .Z(n25631) );
  AND U26238 ( .A(n384), .B(n26529), .Z(n26528) );
  XOR U26239 ( .A(p_input[4668]), .B(p_input[4636]), .Z(n26529) );
  XOR U26240 ( .A(n26530), .B(n26531), .Z(n26521) );
  AND U26241 ( .A(n26532), .B(n26533), .Z(n26531) );
  XOR U26242 ( .A(n26530), .B(n25646), .Z(n26533) );
  XNOR U26243 ( .A(p_input[4699]), .B(n26534), .Z(n25646) );
  AND U26244 ( .A(n387), .B(n26535), .Z(n26534) );
  XOR U26245 ( .A(p_input[4731]), .B(p_input[4699]), .Z(n26535) );
  XNOR U26246 ( .A(n25643), .B(n26530), .Z(n26532) );
  XOR U26247 ( .A(n26536), .B(n26537), .Z(n25643) );
  AND U26248 ( .A(n384), .B(n26538), .Z(n26537) );
  XOR U26249 ( .A(p_input[4667]), .B(p_input[4635]), .Z(n26538) );
  XOR U26250 ( .A(n26539), .B(n26540), .Z(n26530) );
  AND U26251 ( .A(n26541), .B(n26542), .Z(n26540) );
  XOR U26252 ( .A(n26539), .B(n25658), .Z(n26542) );
  XNOR U26253 ( .A(p_input[4698]), .B(n26543), .Z(n25658) );
  AND U26254 ( .A(n387), .B(n26544), .Z(n26543) );
  XOR U26255 ( .A(p_input[4730]), .B(p_input[4698]), .Z(n26544) );
  XNOR U26256 ( .A(n25655), .B(n26539), .Z(n26541) );
  XOR U26257 ( .A(n26545), .B(n26546), .Z(n25655) );
  AND U26258 ( .A(n384), .B(n26547), .Z(n26546) );
  XOR U26259 ( .A(p_input[4666]), .B(p_input[4634]), .Z(n26547) );
  XOR U26260 ( .A(n26548), .B(n26549), .Z(n26539) );
  AND U26261 ( .A(n26550), .B(n26551), .Z(n26549) );
  XOR U26262 ( .A(n26548), .B(n25670), .Z(n26551) );
  XNOR U26263 ( .A(p_input[4697]), .B(n26552), .Z(n25670) );
  AND U26264 ( .A(n387), .B(n26553), .Z(n26552) );
  XOR U26265 ( .A(p_input[4729]), .B(p_input[4697]), .Z(n26553) );
  XNOR U26266 ( .A(n25667), .B(n26548), .Z(n26550) );
  XOR U26267 ( .A(n26554), .B(n26555), .Z(n25667) );
  AND U26268 ( .A(n384), .B(n26556), .Z(n26555) );
  XOR U26269 ( .A(p_input[4665]), .B(p_input[4633]), .Z(n26556) );
  XOR U26270 ( .A(n26557), .B(n26558), .Z(n26548) );
  AND U26271 ( .A(n26559), .B(n26560), .Z(n26558) );
  XOR U26272 ( .A(n26557), .B(n25682), .Z(n26560) );
  XNOR U26273 ( .A(p_input[4696]), .B(n26561), .Z(n25682) );
  AND U26274 ( .A(n387), .B(n26562), .Z(n26561) );
  XOR U26275 ( .A(p_input[4728]), .B(p_input[4696]), .Z(n26562) );
  XNOR U26276 ( .A(n25679), .B(n26557), .Z(n26559) );
  XOR U26277 ( .A(n26563), .B(n26564), .Z(n25679) );
  AND U26278 ( .A(n384), .B(n26565), .Z(n26564) );
  XOR U26279 ( .A(p_input[4664]), .B(p_input[4632]), .Z(n26565) );
  XOR U26280 ( .A(n26566), .B(n26567), .Z(n26557) );
  AND U26281 ( .A(n26568), .B(n26569), .Z(n26567) );
  XOR U26282 ( .A(n26566), .B(n25694), .Z(n26569) );
  XNOR U26283 ( .A(p_input[4695]), .B(n26570), .Z(n25694) );
  AND U26284 ( .A(n387), .B(n26571), .Z(n26570) );
  XOR U26285 ( .A(p_input[4727]), .B(p_input[4695]), .Z(n26571) );
  XNOR U26286 ( .A(n25691), .B(n26566), .Z(n26568) );
  XOR U26287 ( .A(n26572), .B(n26573), .Z(n25691) );
  AND U26288 ( .A(n384), .B(n26574), .Z(n26573) );
  XOR U26289 ( .A(p_input[4663]), .B(p_input[4631]), .Z(n26574) );
  XOR U26290 ( .A(n26575), .B(n26576), .Z(n26566) );
  AND U26291 ( .A(n26577), .B(n26578), .Z(n26576) );
  XOR U26292 ( .A(n26575), .B(n25706), .Z(n26578) );
  XNOR U26293 ( .A(p_input[4694]), .B(n26579), .Z(n25706) );
  AND U26294 ( .A(n387), .B(n26580), .Z(n26579) );
  XOR U26295 ( .A(p_input[4726]), .B(p_input[4694]), .Z(n26580) );
  XNOR U26296 ( .A(n25703), .B(n26575), .Z(n26577) );
  XOR U26297 ( .A(n26581), .B(n26582), .Z(n25703) );
  AND U26298 ( .A(n384), .B(n26583), .Z(n26582) );
  XOR U26299 ( .A(p_input[4662]), .B(p_input[4630]), .Z(n26583) );
  XOR U26300 ( .A(n26584), .B(n26585), .Z(n26575) );
  AND U26301 ( .A(n26586), .B(n26587), .Z(n26585) );
  XOR U26302 ( .A(n26584), .B(n25718), .Z(n26587) );
  XNOR U26303 ( .A(p_input[4693]), .B(n26588), .Z(n25718) );
  AND U26304 ( .A(n387), .B(n26589), .Z(n26588) );
  XOR U26305 ( .A(p_input[4725]), .B(p_input[4693]), .Z(n26589) );
  XNOR U26306 ( .A(n25715), .B(n26584), .Z(n26586) );
  XOR U26307 ( .A(n26590), .B(n26591), .Z(n25715) );
  AND U26308 ( .A(n384), .B(n26592), .Z(n26591) );
  XOR U26309 ( .A(p_input[4661]), .B(p_input[4629]), .Z(n26592) );
  XOR U26310 ( .A(n26593), .B(n26594), .Z(n26584) );
  AND U26311 ( .A(n26595), .B(n26596), .Z(n26594) );
  XOR U26312 ( .A(n26593), .B(n25730), .Z(n26596) );
  XNOR U26313 ( .A(p_input[4692]), .B(n26597), .Z(n25730) );
  AND U26314 ( .A(n387), .B(n26598), .Z(n26597) );
  XOR U26315 ( .A(p_input[4724]), .B(p_input[4692]), .Z(n26598) );
  XNOR U26316 ( .A(n25727), .B(n26593), .Z(n26595) );
  XOR U26317 ( .A(n26599), .B(n26600), .Z(n25727) );
  AND U26318 ( .A(n384), .B(n26601), .Z(n26600) );
  XOR U26319 ( .A(p_input[4660]), .B(p_input[4628]), .Z(n26601) );
  XOR U26320 ( .A(n26602), .B(n26603), .Z(n26593) );
  AND U26321 ( .A(n26604), .B(n26605), .Z(n26603) );
  XOR U26322 ( .A(n26602), .B(n25742), .Z(n26605) );
  XNOR U26323 ( .A(p_input[4691]), .B(n26606), .Z(n25742) );
  AND U26324 ( .A(n387), .B(n26607), .Z(n26606) );
  XOR U26325 ( .A(p_input[4723]), .B(p_input[4691]), .Z(n26607) );
  XNOR U26326 ( .A(n25739), .B(n26602), .Z(n26604) );
  XOR U26327 ( .A(n26608), .B(n26609), .Z(n25739) );
  AND U26328 ( .A(n384), .B(n26610), .Z(n26609) );
  XOR U26329 ( .A(p_input[4659]), .B(p_input[4627]), .Z(n26610) );
  XOR U26330 ( .A(n26611), .B(n26612), .Z(n26602) );
  AND U26331 ( .A(n26613), .B(n26614), .Z(n26612) );
  XOR U26332 ( .A(n26611), .B(n25754), .Z(n26614) );
  XNOR U26333 ( .A(p_input[4690]), .B(n26615), .Z(n25754) );
  AND U26334 ( .A(n387), .B(n26616), .Z(n26615) );
  XOR U26335 ( .A(p_input[4722]), .B(p_input[4690]), .Z(n26616) );
  XNOR U26336 ( .A(n25751), .B(n26611), .Z(n26613) );
  XOR U26337 ( .A(n26617), .B(n26618), .Z(n25751) );
  AND U26338 ( .A(n384), .B(n26619), .Z(n26618) );
  XOR U26339 ( .A(p_input[4658]), .B(p_input[4626]), .Z(n26619) );
  XOR U26340 ( .A(n26620), .B(n26621), .Z(n26611) );
  AND U26341 ( .A(n26622), .B(n26623), .Z(n26621) );
  XOR U26342 ( .A(n26620), .B(n25766), .Z(n26623) );
  XNOR U26343 ( .A(p_input[4689]), .B(n26624), .Z(n25766) );
  AND U26344 ( .A(n387), .B(n26625), .Z(n26624) );
  XOR U26345 ( .A(p_input[4721]), .B(p_input[4689]), .Z(n26625) );
  XNOR U26346 ( .A(n25763), .B(n26620), .Z(n26622) );
  XOR U26347 ( .A(n26626), .B(n26627), .Z(n25763) );
  AND U26348 ( .A(n384), .B(n26628), .Z(n26627) );
  XOR U26349 ( .A(p_input[4657]), .B(p_input[4625]), .Z(n26628) );
  XOR U26350 ( .A(n26629), .B(n26630), .Z(n26620) );
  AND U26351 ( .A(n26631), .B(n26632), .Z(n26630) );
  XOR U26352 ( .A(n26629), .B(n25778), .Z(n26632) );
  XNOR U26353 ( .A(p_input[4688]), .B(n26633), .Z(n25778) );
  AND U26354 ( .A(n387), .B(n26634), .Z(n26633) );
  XOR U26355 ( .A(p_input[4720]), .B(p_input[4688]), .Z(n26634) );
  XNOR U26356 ( .A(n25775), .B(n26629), .Z(n26631) );
  XOR U26357 ( .A(n26635), .B(n26636), .Z(n25775) );
  AND U26358 ( .A(n384), .B(n26637), .Z(n26636) );
  XOR U26359 ( .A(p_input[4656]), .B(p_input[4624]), .Z(n26637) );
  XOR U26360 ( .A(n26638), .B(n26639), .Z(n26629) );
  AND U26361 ( .A(n26640), .B(n26641), .Z(n26639) );
  XOR U26362 ( .A(n26638), .B(n25790), .Z(n26641) );
  XNOR U26363 ( .A(p_input[4687]), .B(n26642), .Z(n25790) );
  AND U26364 ( .A(n387), .B(n26643), .Z(n26642) );
  XOR U26365 ( .A(p_input[4719]), .B(p_input[4687]), .Z(n26643) );
  XNOR U26366 ( .A(n25787), .B(n26638), .Z(n26640) );
  XOR U26367 ( .A(n26644), .B(n26645), .Z(n25787) );
  AND U26368 ( .A(n384), .B(n26646), .Z(n26645) );
  XOR U26369 ( .A(p_input[4655]), .B(p_input[4623]), .Z(n26646) );
  XOR U26370 ( .A(n26647), .B(n26648), .Z(n26638) );
  AND U26371 ( .A(n26649), .B(n26650), .Z(n26648) );
  XOR U26372 ( .A(n26647), .B(n25802), .Z(n26650) );
  XNOR U26373 ( .A(p_input[4686]), .B(n26651), .Z(n25802) );
  AND U26374 ( .A(n387), .B(n26652), .Z(n26651) );
  XOR U26375 ( .A(p_input[4718]), .B(p_input[4686]), .Z(n26652) );
  XNOR U26376 ( .A(n25799), .B(n26647), .Z(n26649) );
  XOR U26377 ( .A(n26653), .B(n26654), .Z(n25799) );
  AND U26378 ( .A(n384), .B(n26655), .Z(n26654) );
  XOR U26379 ( .A(p_input[4654]), .B(p_input[4622]), .Z(n26655) );
  XOR U26380 ( .A(n26656), .B(n26657), .Z(n26647) );
  AND U26381 ( .A(n26658), .B(n26659), .Z(n26657) );
  XOR U26382 ( .A(n26656), .B(n25814), .Z(n26659) );
  XNOR U26383 ( .A(p_input[4685]), .B(n26660), .Z(n25814) );
  AND U26384 ( .A(n387), .B(n26661), .Z(n26660) );
  XOR U26385 ( .A(p_input[4717]), .B(p_input[4685]), .Z(n26661) );
  XNOR U26386 ( .A(n25811), .B(n26656), .Z(n26658) );
  XOR U26387 ( .A(n26662), .B(n26663), .Z(n25811) );
  AND U26388 ( .A(n384), .B(n26664), .Z(n26663) );
  XOR U26389 ( .A(p_input[4653]), .B(p_input[4621]), .Z(n26664) );
  XOR U26390 ( .A(n26665), .B(n26666), .Z(n26656) );
  AND U26391 ( .A(n26667), .B(n26668), .Z(n26666) );
  XOR U26392 ( .A(n26665), .B(n25826), .Z(n26668) );
  XNOR U26393 ( .A(p_input[4684]), .B(n26669), .Z(n25826) );
  AND U26394 ( .A(n387), .B(n26670), .Z(n26669) );
  XOR U26395 ( .A(p_input[4716]), .B(p_input[4684]), .Z(n26670) );
  XNOR U26396 ( .A(n25823), .B(n26665), .Z(n26667) );
  XOR U26397 ( .A(n26671), .B(n26672), .Z(n25823) );
  AND U26398 ( .A(n384), .B(n26673), .Z(n26672) );
  XOR U26399 ( .A(p_input[4652]), .B(p_input[4620]), .Z(n26673) );
  XOR U26400 ( .A(n26674), .B(n26675), .Z(n26665) );
  AND U26401 ( .A(n26676), .B(n26677), .Z(n26675) );
  XOR U26402 ( .A(n26674), .B(n25838), .Z(n26677) );
  XNOR U26403 ( .A(p_input[4683]), .B(n26678), .Z(n25838) );
  AND U26404 ( .A(n387), .B(n26679), .Z(n26678) );
  XOR U26405 ( .A(p_input[4715]), .B(p_input[4683]), .Z(n26679) );
  XNOR U26406 ( .A(n25835), .B(n26674), .Z(n26676) );
  XOR U26407 ( .A(n26680), .B(n26681), .Z(n25835) );
  AND U26408 ( .A(n384), .B(n26682), .Z(n26681) );
  XOR U26409 ( .A(p_input[4651]), .B(p_input[4619]), .Z(n26682) );
  XOR U26410 ( .A(n26683), .B(n26684), .Z(n26674) );
  AND U26411 ( .A(n26685), .B(n26686), .Z(n26684) );
  XOR U26412 ( .A(n26683), .B(n25850), .Z(n26686) );
  XNOR U26413 ( .A(p_input[4682]), .B(n26687), .Z(n25850) );
  AND U26414 ( .A(n387), .B(n26688), .Z(n26687) );
  XOR U26415 ( .A(p_input[4714]), .B(p_input[4682]), .Z(n26688) );
  XNOR U26416 ( .A(n25847), .B(n26683), .Z(n26685) );
  XOR U26417 ( .A(n26689), .B(n26690), .Z(n25847) );
  AND U26418 ( .A(n384), .B(n26691), .Z(n26690) );
  XOR U26419 ( .A(p_input[4650]), .B(p_input[4618]), .Z(n26691) );
  XOR U26420 ( .A(n26692), .B(n26693), .Z(n26683) );
  AND U26421 ( .A(n26694), .B(n26695), .Z(n26693) );
  XOR U26422 ( .A(n26692), .B(n25862), .Z(n26695) );
  XNOR U26423 ( .A(p_input[4681]), .B(n26696), .Z(n25862) );
  AND U26424 ( .A(n387), .B(n26697), .Z(n26696) );
  XOR U26425 ( .A(p_input[4713]), .B(p_input[4681]), .Z(n26697) );
  XNOR U26426 ( .A(n25859), .B(n26692), .Z(n26694) );
  XOR U26427 ( .A(n26698), .B(n26699), .Z(n25859) );
  AND U26428 ( .A(n384), .B(n26700), .Z(n26699) );
  XOR U26429 ( .A(p_input[4649]), .B(p_input[4617]), .Z(n26700) );
  XOR U26430 ( .A(n26701), .B(n26702), .Z(n26692) );
  AND U26431 ( .A(n26703), .B(n26704), .Z(n26702) );
  XOR U26432 ( .A(n26701), .B(n25874), .Z(n26704) );
  XNOR U26433 ( .A(p_input[4680]), .B(n26705), .Z(n25874) );
  AND U26434 ( .A(n387), .B(n26706), .Z(n26705) );
  XOR U26435 ( .A(p_input[4712]), .B(p_input[4680]), .Z(n26706) );
  XNOR U26436 ( .A(n25871), .B(n26701), .Z(n26703) );
  XOR U26437 ( .A(n26707), .B(n26708), .Z(n25871) );
  AND U26438 ( .A(n384), .B(n26709), .Z(n26708) );
  XOR U26439 ( .A(p_input[4648]), .B(p_input[4616]), .Z(n26709) );
  XOR U26440 ( .A(n26710), .B(n26711), .Z(n26701) );
  AND U26441 ( .A(n26712), .B(n26713), .Z(n26711) );
  XOR U26442 ( .A(n26710), .B(n25886), .Z(n26713) );
  XNOR U26443 ( .A(p_input[4679]), .B(n26714), .Z(n25886) );
  AND U26444 ( .A(n387), .B(n26715), .Z(n26714) );
  XOR U26445 ( .A(p_input[4711]), .B(p_input[4679]), .Z(n26715) );
  XNOR U26446 ( .A(n25883), .B(n26710), .Z(n26712) );
  XOR U26447 ( .A(n26716), .B(n26717), .Z(n25883) );
  AND U26448 ( .A(n384), .B(n26718), .Z(n26717) );
  XOR U26449 ( .A(p_input[4647]), .B(p_input[4615]), .Z(n26718) );
  XOR U26450 ( .A(n26719), .B(n26720), .Z(n26710) );
  AND U26451 ( .A(n26721), .B(n26722), .Z(n26720) );
  XOR U26452 ( .A(n26719), .B(n25898), .Z(n26722) );
  XNOR U26453 ( .A(p_input[4678]), .B(n26723), .Z(n25898) );
  AND U26454 ( .A(n387), .B(n26724), .Z(n26723) );
  XOR U26455 ( .A(p_input[4710]), .B(p_input[4678]), .Z(n26724) );
  XNOR U26456 ( .A(n25895), .B(n26719), .Z(n26721) );
  XOR U26457 ( .A(n26725), .B(n26726), .Z(n25895) );
  AND U26458 ( .A(n384), .B(n26727), .Z(n26726) );
  XOR U26459 ( .A(p_input[4646]), .B(p_input[4614]), .Z(n26727) );
  XOR U26460 ( .A(n26728), .B(n26729), .Z(n26719) );
  AND U26461 ( .A(n26730), .B(n26731), .Z(n26729) );
  XOR U26462 ( .A(n26728), .B(n25910), .Z(n26731) );
  XNOR U26463 ( .A(p_input[4677]), .B(n26732), .Z(n25910) );
  AND U26464 ( .A(n387), .B(n26733), .Z(n26732) );
  XOR U26465 ( .A(p_input[4709]), .B(p_input[4677]), .Z(n26733) );
  XNOR U26466 ( .A(n25907), .B(n26728), .Z(n26730) );
  XOR U26467 ( .A(n26734), .B(n26735), .Z(n25907) );
  AND U26468 ( .A(n384), .B(n26736), .Z(n26735) );
  XOR U26469 ( .A(p_input[4645]), .B(p_input[4613]), .Z(n26736) );
  XOR U26470 ( .A(n26737), .B(n26738), .Z(n26728) );
  AND U26471 ( .A(n26739), .B(n26740), .Z(n26738) );
  XOR U26472 ( .A(n26737), .B(n25922), .Z(n26740) );
  XNOR U26473 ( .A(p_input[4676]), .B(n26741), .Z(n25922) );
  AND U26474 ( .A(n387), .B(n26742), .Z(n26741) );
  XOR U26475 ( .A(p_input[4708]), .B(p_input[4676]), .Z(n26742) );
  XNOR U26476 ( .A(n25919), .B(n26737), .Z(n26739) );
  XOR U26477 ( .A(n26743), .B(n26744), .Z(n25919) );
  AND U26478 ( .A(n384), .B(n26745), .Z(n26744) );
  XOR U26479 ( .A(p_input[4644]), .B(p_input[4612]), .Z(n26745) );
  XOR U26480 ( .A(n26746), .B(n26747), .Z(n26737) );
  AND U26481 ( .A(n26748), .B(n26749), .Z(n26747) );
  XOR U26482 ( .A(n26746), .B(n25934), .Z(n26749) );
  XNOR U26483 ( .A(p_input[4675]), .B(n26750), .Z(n25934) );
  AND U26484 ( .A(n387), .B(n26751), .Z(n26750) );
  XOR U26485 ( .A(p_input[4707]), .B(p_input[4675]), .Z(n26751) );
  XNOR U26486 ( .A(n25931), .B(n26746), .Z(n26748) );
  XOR U26487 ( .A(n26752), .B(n26753), .Z(n25931) );
  AND U26488 ( .A(n384), .B(n26754), .Z(n26753) );
  XOR U26489 ( .A(p_input[4643]), .B(p_input[4611]), .Z(n26754) );
  XOR U26490 ( .A(n26755), .B(n26756), .Z(n26746) );
  AND U26491 ( .A(n26757), .B(n26758), .Z(n26756) );
  XOR U26492 ( .A(n26755), .B(n25946), .Z(n26758) );
  XNOR U26493 ( .A(p_input[4674]), .B(n26759), .Z(n25946) );
  AND U26494 ( .A(n387), .B(n26760), .Z(n26759) );
  XOR U26495 ( .A(p_input[4706]), .B(p_input[4674]), .Z(n26760) );
  XNOR U26496 ( .A(n25943), .B(n26755), .Z(n26757) );
  XOR U26497 ( .A(n26761), .B(n26762), .Z(n25943) );
  AND U26498 ( .A(n384), .B(n26763), .Z(n26762) );
  XOR U26499 ( .A(p_input[4642]), .B(p_input[4610]), .Z(n26763) );
  XOR U26500 ( .A(n26764), .B(n26765), .Z(n26755) );
  AND U26501 ( .A(n26766), .B(n26767), .Z(n26765) );
  XNOR U26502 ( .A(n26768), .B(n25959), .Z(n26767) );
  XNOR U26503 ( .A(p_input[4673]), .B(n26769), .Z(n25959) );
  AND U26504 ( .A(n387), .B(n26770), .Z(n26769) );
  XNOR U26505 ( .A(p_input[4705]), .B(n26771), .Z(n26770) );
  IV U26506 ( .A(p_input[4673]), .Z(n26771) );
  XNOR U26507 ( .A(n25956), .B(n26764), .Z(n26766) );
  XNOR U26508 ( .A(p_input[4609]), .B(n26772), .Z(n25956) );
  AND U26509 ( .A(n384), .B(n26773), .Z(n26772) );
  XOR U26510 ( .A(p_input[4641]), .B(p_input[4609]), .Z(n26773) );
  IV U26511 ( .A(n26768), .Z(n26764) );
  AND U26512 ( .A(n26494), .B(n26497), .Z(n26768) );
  XOR U26513 ( .A(p_input[4672]), .B(n26774), .Z(n26497) );
  AND U26514 ( .A(n387), .B(n26775), .Z(n26774) );
  XOR U26515 ( .A(p_input[4704]), .B(p_input[4672]), .Z(n26775) );
  XOR U26516 ( .A(n26776), .B(n26777), .Z(n387) );
  AND U26517 ( .A(n26778), .B(n26779), .Z(n26777) );
  XNOR U26518 ( .A(p_input[4735]), .B(n26776), .Z(n26779) );
  XOR U26519 ( .A(n26776), .B(p_input[4703]), .Z(n26778) );
  XOR U26520 ( .A(n26780), .B(n26781), .Z(n26776) );
  AND U26521 ( .A(n26782), .B(n26783), .Z(n26781) );
  XNOR U26522 ( .A(p_input[4734]), .B(n26780), .Z(n26783) );
  XOR U26523 ( .A(n26780), .B(p_input[4702]), .Z(n26782) );
  XOR U26524 ( .A(n26784), .B(n26785), .Z(n26780) );
  AND U26525 ( .A(n26786), .B(n26787), .Z(n26785) );
  XNOR U26526 ( .A(p_input[4733]), .B(n26784), .Z(n26787) );
  XOR U26527 ( .A(n26784), .B(p_input[4701]), .Z(n26786) );
  XOR U26528 ( .A(n26788), .B(n26789), .Z(n26784) );
  AND U26529 ( .A(n26790), .B(n26791), .Z(n26789) );
  XNOR U26530 ( .A(p_input[4732]), .B(n26788), .Z(n26791) );
  XOR U26531 ( .A(n26788), .B(p_input[4700]), .Z(n26790) );
  XOR U26532 ( .A(n26792), .B(n26793), .Z(n26788) );
  AND U26533 ( .A(n26794), .B(n26795), .Z(n26793) );
  XNOR U26534 ( .A(p_input[4731]), .B(n26792), .Z(n26795) );
  XOR U26535 ( .A(n26792), .B(p_input[4699]), .Z(n26794) );
  XOR U26536 ( .A(n26796), .B(n26797), .Z(n26792) );
  AND U26537 ( .A(n26798), .B(n26799), .Z(n26797) );
  XNOR U26538 ( .A(p_input[4730]), .B(n26796), .Z(n26799) );
  XOR U26539 ( .A(n26796), .B(p_input[4698]), .Z(n26798) );
  XOR U26540 ( .A(n26800), .B(n26801), .Z(n26796) );
  AND U26541 ( .A(n26802), .B(n26803), .Z(n26801) );
  XNOR U26542 ( .A(p_input[4729]), .B(n26800), .Z(n26803) );
  XOR U26543 ( .A(n26800), .B(p_input[4697]), .Z(n26802) );
  XOR U26544 ( .A(n26804), .B(n26805), .Z(n26800) );
  AND U26545 ( .A(n26806), .B(n26807), .Z(n26805) );
  XNOR U26546 ( .A(p_input[4728]), .B(n26804), .Z(n26807) );
  XOR U26547 ( .A(n26804), .B(p_input[4696]), .Z(n26806) );
  XOR U26548 ( .A(n26808), .B(n26809), .Z(n26804) );
  AND U26549 ( .A(n26810), .B(n26811), .Z(n26809) );
  XNOR U26550 ( .A(p_input[4727]), .B(n26808), .Z(n26811) );
  XOR U26551 ( .A(n26808), .B(p_input[4695]), .Z(n26810) );
  XOR U26552 ( .A(n26812), .B(n26813), .Z(n26808) );
  AND U26553 ( .A(n26814), .B(n26815), .Z(n26813) );
  XNOR U26554 ( .A(p_input[4726]), .B(n26812), .Z(n26815) );
  XOR U26555 ( .A(n26812), .B(p_input[4694]), .Z(n26814) );
  XOR U26556 ( .A(n26816), .B(n26817), .Z(n26812) );
  AND U26557 ( .A(n26818), .B(n26819), .Z(n26817) );
  XNOR U26558 ( .A(p_input[4725]), .B(n26816), .Z(n26819) );
  XOR U26559 ( .A(n26816), .B(p_input[4693]), .Z(n26818) );
  XOR U26560 ( .A(n26820), .B(n26821), .Z(n26816) );
  AND U26561 ( .A(n26822), .B(n26823), .Z(n26821) );
  XNOR U26562 ( .A(p_input[4724]), .B(n26820), .Z(n26823) );
  XOR U26563 ( .A(n26820), .B(p_input[4692]), .Z(n26822) );
  XOR U26564 ( .A(n26824), .B(n26825), .Z(n26820) );
  AND U26565 ( .A(n26826), .B(n26827), .Z(n26825) );
  XNOR U26566 ( .A(p_input[4723]), .B(n26824), .Z(n26827) );
  XOR U26567 ( .A(n26824), .B(p_input[4691]), .Z(n26826) );
  XOR U26568 ( .A(n26828), .B(n26829), .Z(n26824) );
  AND U26569 ( .A(n26830), .B(n26831), .Z(n26829) );
  XNOR U26570 ( .A(p_input[4722]), .B(n26828), .Z(n26831) );
  XOR U26571 ( .A(n26828), .B(p_input[4690]), .Z(n26830) );
  XOR U26572 ( .A(n26832), .B(n26833), .Z(n26828) );
  AND U26573 ( .A(n26834), .B(n26835), .Z(n26833) );
  XNOR U26574 ( .A(p_input[4721]), .B(n26832), .Z(n26835) );
  XOR U26575 ( .A(n26832), .B(p_input[4689]), .Z(n26834) );
  XOR U26576 ( .A(n26836), .B(n26837), .Z(n26832) );
  AND U26577 ( .A(n26838), .B(n26839), .Z(n26837) );
  XNOR U26578 ( .A(p_input[4720]), .B(n26836), .Z(n26839) );
  XOR U26579 ( .A(n26836), .B(p_input[4688]), .Z(n26838) );
  XOR U26580 ( .A(n26840), .B(n26841), .Z(n26836) );
  AND U26581 ( .A(n26842), .B(n26843), .Z(n26841) );
  XNOR U26582 ( .A(p_input[4719]), .B(n26840), .Z(n26843) );
  XOR U26583 ( .A(n26840), .B(p_input[4687]), .Z(n26842) );
  XOR U26584 ( .A(n26844), .B(n26845), .Z(n26840) );
  AND U26585 ( .A(n26846), .B(n26847), .Z(n26845) );
  XNOR U26586 ( .A(p_input[4718]), .B(n26844), .Z(n26847) );
  XOR U26587 ( .A(n26844), .B(p_input[4686]), .Z(n26846) );
  XOR U26588 ( .A(n26848), .B(n26849), .Z(n26844) );
  AND U26589 ( .A(n26850), .B(n26851), .Z(n26849) );
  XNOR U26590 ( .A(p_input[4717]), .B(n26848), .Z(n26851) );
  XOR U26591 ( .A(n26848), .B(p_input[4685]), .Z(n26850) );
  XOR U26592 ( .A(n26852), .B(n26853), .Z(n26848) );
  AND U26593 ( .A(n26854), .B(n26855), .Z(n26853) );
  XNOR U26594 ( .A(p_input[4716]), .B(n26852), .Z(n26855) );
  XOR U26595 ( .A(n26852), .B(p_input[4684]), .Z(n26854) );
  XOR U26596 ( .A(n26856), .B(n26857), .Z(n26852) );
  AND U26597 ( .A(n26858), .B(n26859), .Z(n26857) );
  XNOR U26598 ( .A(p_input[4715]), .B(n26856), .Z(n26859) );
  XOR U26599 ( .A(n26856), .B(p_input[4683]), .Z(n26858) );
  XOR U26600 ( .A(n26860), .B(n26861), .Z(n26856) );
  AND U26601 ( .A(n26862), .B(n26863), .Z(n26861) );
  XNOR U26602 ( .A(p_input[4714]), .B(n26860), .Z(n26863) );
  XOR U26603 ( .A(n26860), .B(p_input[4682]), .Z(n26862) );
  XOR U26604 ( .A(n26864), .B(n26865), .Z(n26860) );
  AND U26605 ( .A(n26866), .B(n26867), .Z(n26865) );
  XNOR U26606 ( .A(p_input[4713]), .B(n26864), .Z(n26867) );
  XOR U26607 ( .A(n26864), .B(p_input[4681]), .Z(n26866) );
  XOR U26608 ( .A(n26868), .B(n26869), .Z(n26864) );
  AND U26609 ( .A(n26870), .B(n26871), .Z(n26869) );
  XNOR U26610 ( .A(p_input[4712]), .B(n26868), .Z(n26871) );
  XOR U26611 ( .A(n26868), .B(p_input[4680]), .Z(n26870) );
  XOR U26612 ( .A(n26872), .B(n26873), .Z(n26868) );
  AND U26613 ( .A(n26874), .B(n26875), .Z(n26873) );
  XNOR U26614 ( .A(p_input[4711]), .B(n26872), .Z(n26875) );
  XOR U26615 ( .A(n26872), .B(p_input[4679]), .Z(n26874) );
  XOR U26616 ( .A(n26876), .B(n26877), .Z(n26872) );
  AND U26617 ( .A(n26878), .B(n26879), .Z(n26877) );
  XNOR U26618 ( .A(p_input[4710]), .B(n26876), .Z(n26879) );
  XOR U26619 ( .A(n26876), .B(p_input[4678]), .Z(n26878) );
  XOR U26620 ( .A(n26880), .B(n26881), .Z(n26876) );
  AND U26621 ( .A(n26882), .B(n26883), .Z(n26881) );
  XNOR U26622 ( .A(p_input[4709]), .B(n26880), .Z(n26883) );
  XOR U26623 ( .A(n26880), .B(p_input[4677]), .Z(n26882) );
  XOR U26624 ( .A(n26884), .B(n26885), .Z(n26880) );
  AND U26625 ( .A(n26886), .B(n26887), .Z(n26885) );
  XNOR U26626 ( .A(p_input[4708]), .B(n26884), .Z(n26887) );
  XOR U26627 ( .A(n26884), .B(p_input[4676]), .Z(n26886) );
  XOR U26628 ( .A(n26888), .B(n26889), .Z(n26884) );
  AND U26629 ( .A(n26890), .B(n26891), .Z(n26889) );
  XNOR U26630 ( .A(p_input[4707]), .B(n26888), .Z(n26891) );
  XOR U26631 ( .A(n26888), .B(p_input[4675]), .Z(n26890) );
  XOR U26632 ( .A(n26892), .B(n26893), .Z(n26888) );
  AND U26633 ( .A(n26894), .B(n26895), .Z(n26893) );
  XNOR U26634 ( .A(p_input[4706]), .B(n26892), .Z(n26895) );
  XOR U26635 ( .A(n26892), .B(p_input[4674]), .Z(n26894) );
  XNOR U26636 ( .A(n26896), .B(n26897), .Z(n26892) );
  AND U26637 ( .A(n26898), .B(n26899), .Z(n26897) );
  XOR U26638 ( .A(p_input[4705]), .B(n26896), .Z(n26899) );
  XNOR U26639 ( .A(p_input[4673]), .B(n26896), .Z(n26898) );
  AND U26640 ( .A(p_input[4704]), .B(n26900), .Z(n26896) );
  IV U26641 ( .A(p_input[4672]), .Z(n26900) );
  XNOR U26642 ( .A(p_input[4608]), .B(n26901), .Z(n26494) );
  AND U26643 ( .A(n384), .B(n26902), .Z(n26901) );
  XOR U26644 ( .A(p_input[4640]), .B(p_input[4608]), .Z(n26902) );
  XOR U26645 ( .A(n26903), .B(n26904), .Z(n384) );
  AND U26646 ( .A(n26905), .B(n26906), .Z(n26904) );
  XNOR U26647 ( .A(p_input[4671]), .B(n26903), .Z(n26906) );
  XOR U26648 ( .A(n26903), .B(p_input[4639]), .Z(n26905) );
  XOR U26649 ( .A(n26907), .B(n26908), .Z(n26903) );
  AND U26650 ( .A(n26909), .B(n26910), .Z(n26908) );
  XNOR U26651 ( .A(p_input[4670]), .B(n26907), .Z(n26910) );
  XNOR U26652 ( .A(n26907), .B(n26509), .Z(n26909) );
  IV U26653 ( .A(p_input[4638]), .Z(n26509) );
  XOR U26654 ( .A(n26911), .B(n26912), .Z(n26907) );
  AND U26655 ( .A(n26913), .B(n26914), .Z(n26912) );
  XNOR U26656 ( .A(p_input[4669]), .B(n26911), .Z(n26914) );
  XNOR U26657 ( .A(n26911), .B(n26518), .Z(n26913) );
  IV U26658 ( .A(p_input[4637]), .Z(n26518) );
  XOR U26659 ( .A(n26915), .B(n26916), .Z(n26911) );
  AND U26660 ( .A(n26917), .B(n26918), .Z(n26916) );
  XNOR U26661 ( .A(p_input[4668]), .B(n26915), .Z(n26918) );
  XNOR U26662 ( .A(n26915), .B(n26527), .Z(n26917) );
  IV U26663 ( .A(p_input[4636]), .Z(n26527) );
  XOR U26664 ( .A(n26919), .B(n26920), .Z(n26915) );
  AND U26665 ( .A(n26921), .B(n26922), .Z(n26920) );
  XNOR U26666 ( .A(p_input[4667]), .B(n26919), .Z(n26922) );
  XNOR U26667 ( .A(n26919), .B(n26536), .Z(n26921) );
  IV U26668 ( .A(p_input[4635]), .Z(n26536) );
  XOR U26669 ( .A(n26923), .B(n26924), .Z(n26919) );
  AND U26670 ( .A(n26925), .B(n26926), .Z(n26924) );
  XNOR U26671 ( .A(p_input[4666]), .B(n26923), .Z(n26926) );
  XNOR U26672 ( .A(n26923), .B(n26545), .Z(n26925) );
  IV U26673 ( .A(p_input[4634]), .Z(n26545) );
  XOR U26674 ( .A(n26927), .B(n26928), .Z(n26923) );
  AND U26675 ( .A(n26929), .B(n26930), .Z(n26928) );
  XNOR U26676 ( .A(p_input[4665]), .B(n26927), .Z(n26930) );
  XNOR U26677 ( .A(n26927), .B(n26554), .Z(n26929) );
  IV U26678 ( .A(p_input[4633]), .Z(n26554) );
  XOR U26679 ( .A(n26931), .B(n26932), .Z(n26927) );
  AND U26680 ( .A(n26933), .B(n26934), .Z(n26932) );
  XNOR U26681 ( .A(p_input[4664]), .B(n26931), .Z(n26934) );
  XNOR U26682 ( .A(n26931), .B(n26563), .Z(n26933) );
  IV U26683 ( .A(p_input[4632]), .Z(n26563) );
  XOR U26684 ( .A(n26935), .B(n26936), .Z(n26931) );
  AND U26685 ( .A(n26937), .B(n26938), .Z(n26936) );
  XNOR U26686 ( .A(p_input[4663]), .B(n26935), .Z(n26938) );
  XNOR U26687 ( .A(n26935), .B(n26572), .Z(n26937) );
  IV U26688 ( .A(p_input[4631]), .Z(n26572) );
  XOR U26689 ( .A(n26939), .B(n26940), .Z(n26935) );
  AND U26690 ( .A(n26941), .B(n26942), .Z(n26940) );
  XNOR U26691 ( .A(p_input[4662]), .B(n26939), .Z(n26942) );
  XNOR U26692 ( .A(n26939), .B(n26581), .Z(n26941) );
  IV U26693 ( .A(p_input[4630]), .Z(n26581) );
  XOR U26694 ( .A(n26943), .B(n26944), .Z(n26939) );
  AND U26695 ( .A(n26945), .B(n26946), .Z(n26944) );
  XNOR U26696 ( .A(p_input[4661]), .B(n26943), .Z(n26946) );
  XNOR U26697 ( .A(n26943), .B(n26590), .Z(n26945) );
  IV U26698 ( .A(p_input[4629]), .Z(n26590) );
  XOR U26699 ( .A(n26947), .B(n26948), .Z(n26943) );
  AND U26700 ( .A(n26949), .B(n26950), .Z(n26948) );
  XNOR U26701 ( .A(p_input[4660]), .B(n26947), .Z(n26950) );
  XNOR U26702 ( .A(n26947), .B(n26599), .Z(n26949) );
  IV U26703 ( .A(p_input[4628]), .Z(n26599) );
  XOR U26704 ( .A(n26951), .B(n26952), .Z(n26947) );
  AND U26705 ( .A(n26953), .B(n26954), .Z(n26952) );
  XNOR U26706 ( .A(p_input[4659]), .B(n26951), .Z(n26954) );
  XNOR U26707 ( .A(n26951), .B(n26608), .Z(n26953) );
  IV U26708 ( .A(p_input[4627]), .Z(n26608) );
  XOR U26709 ( .A(n26955), .B(n26956), .Z(n26951) );
  AND U26710 ( .A(n26957), .B(n26958), .Z(n26956) );
  XNOR U26711 ( .A(p_input[4658]), .B(n26955), .Z(n26958) );
  XNOR U26712 ( .A(n26955), .B(n26617), .Z(n26957) );
  IV U26713 ( .A(p_input[4626]), .Z(n26617) );
  XOR U26714 ( .A(n26959), .B(n26960), .Z(n26955) );
  AND U26715 ( .A(n26961), .B(n26962), .Z(n26960) );
  XNOR U26716 ( .A(p_input[4657]), .B(n26959), .Z(n26962) );
  XNOR U26717 ( .A(n26959), .B(n26626), .Z(n26961) );
  IV U26718 ( .A(p_input[4625]), .Z(n26626) );
  XOR U26719 ( .A(n26963), .B(n26964), .Z(n26959) );
  AND U26720 ( .A(n26965), .B(n26966), .Z(n26964) );
  XNOR U26721 ( .A(p_input[4656]), .B(n26963), .Z(n26966) );
  XNOR U26722 ( .A(n26963), .B(n26635), .Z(n26965) );
  IV U26723 ( .A(p_input[4624]), .Z(n26635) );
  XOR U26724 ( .A(n26967), .B(n26968), .Z(n26963) );
  AND U26725 ( .A(n26969), .B(n26970), .Z(n26968) );
  XNOR U26726 ( .A(p_input[4655]), .B(n26967), .Z(n26970) );
  XNOR U26727 ( .A(n26967), .B(n26644), .Z(n26969) );
  IV U26728 ( .A(p_input[4623]), .Z(n26644) );
  XOR U26729 ( .A(n26971), .B(n26972), .Z(n26967) );
  AND U26730 ( .A(n26973), .B(n26974), .Z(n26972) );
  XNOR U26731 ( .A(p_input[4654]), .B(n26971), .Z(n26974) );
  XNOR U26732 ( .A(n26971), .B(n26653), .Z(n26973) );
  IV U26733 ( .A(p_input[4622]), .Z(n26653) );
  XOR U26734 ( .A(n26975), .B(n26976), .Z(n26971) );
  AND U26735 ( .A(n26977), .B(n26978), .Z(n26976) );
  XNOR U26736 ( .A(p_input[4653]), .B(n26975), .Z(n26978) );
  XNOR U26737 ( .A(n26975), .B(n26662), .Z(n26977) );
  IV U26738 ( .A(p_input[4621]), .Z(n26662) );
  XOR U26739 ( .A(n26979), .B(n26980), .Z(n26975) );
  AND U26740 ( .A(n26981), .B(n26982), .Z(n26980) );
  XNOR U26741 ( .A(p_input[4652]), .B(n26979), .Z(n26982) );
  XNOR U26742 ( .A(n26979), .B(n26671), .Z(n26981) );
  IV U26743 ( .A(p_input[4620]), .Z(n26671) );
  XOR U26744 ( .A(n26983), .B(n26984), .Z(n26979) );
  AND U26745 ( .A(n26985), .B(n26986), .Z(n26984) );
  XNOR U26746 ( .A(p_input[4651]), .B(n26983), .Z(n26986) );
  XNOR U26747 ( .A(n26983), .B(n26680), .Z(n26985) );
  IV U26748 ( .A(p_input[4619]), .Z(n26680) );
  XOR U26749 ( .A(n26987), .B(n26988), .Z(n26983) );
  AND U26750 ( .A(n26989), .B(n26990), .Z(n26988) );
  XNOR U26751 ( .A(p_input[4650]), .B(n26987), .Z(n26990) );
  XNOR U26752 ( .A(n26987), .B(n26689), .Z(n26989) );
  IV U26753 ( .A(p_input[4618]), .Z(n26689) );
  XOR U26754 ( .A(n26991), .B(n26992), .Z(n26987) );
  AND U26755 ( .A(n26993), .B(n26994), .Z(n26992) );
  XNOR U26756 ( .A(p_input[4649]), .B(n26991), .Z(n26994) );
  XNOR U26757 ( .A(n26991), .B(n26698), .Z(n26993) );
  IV U26758 ( .A(p_input[4617]), .Z(n26698) );
  XOR U26759 ( .A(n26995), .B(n26996), .Z(n26991) );
  AND U26760 ( .A(n26997), .B(n26998), .Z(n26996) );
  XNOR U26761 ( .A(p_input[4648]), .B(n26995), .Z(n26998) );
  XNOR U26762 ( .A(n26995), .B(n26707), .Z(n26997) );
  IV U26763 ( .A(p_input[4616]), .Z(n26707) );
  XOR U26764 ( .A(n26999), .B(n27000), .Z(n26995) );
  AND U26765 ( .A(n27001), .B(n27002), .Z(n27000) );
  XNOR U26766 ( .A(p_input[4647]), .B(n26999), .Z(n27002) );
  XNOR U26767 ( .A(n26999), .B(n26716), .Z(n27001) );
  IV U26768 ( .A(p_input[4615]), .Z(n26716) );
  XOR U26769 ( .A(n27003), .B(n27004), .Z(n26999) );
  AND U26770 ( .A(n27005), .B(n27006), .Z(n27004) );
  XNOR U26771 ( .A(p_input[4646]), .B(n27003), .Z(n27006) );
  XNOR U26772 ( .A(n27003), .B(n26725), .Z(n27005) );
  IV U26773 ( .A(p_input[4614]), .Z(n26725) );
  XOR U26774 ( .A(n27007), .B(n27008), .Z(n27003) );
  AND U26775 ( .A(n27009), .B(n27010), .Z(n27008) );
  XNOR U26776 ( .A(p_input[4645]), .B(n27007), .Z(n27010) );
  XNOR U26777 ( .A(n27007), .B(n26734), .Z(n27009) );
  IV U26778 ( .A(p_input[4613]), .Z(n26734) );
  XOR U26779 ( .A(n27011), .B(n27012), .Z(n27007) );
  AND U26780 ( .A(n27013), .B(n27014), .Z(n27012) );
  XNOR U26781 ( .A(p_input[4644]), .B(n27011), .Z(n27014) );
  XNOR U26782 ( .A(n27011), .B(n26743), .Z(n27013) );
  IV U26783 ( .A(p_input[4612]), .Z(n26743) );
  XOR U26784 ( .A(n27015), .B(n27016), .Z(n27011) );
  AND U26785 ( .A(n27017), .B(n27018), .Z(n27016) );
  XNOR U26786 ( .A(p_input[4643]), .B(n27015), .Z(n27018) );
  XNOR U26787 ( .A(n27015), .B(n26752), .Z(n27017) );
  IV U26788 ( .A(p_input[4611]), .Z(n26752) );
  XOR U26789 ( .A(n27019), .B(n27020), .Z(n27015) );
  AND U26790 ( .A(n27021), .B(n27022), .Z(n27020) );
  XNOR U26791 ( .A(p_input[4642]), .B(n27019), .Z(n27022) );
  XNOR U26792 ( .A(n27019), .B(n26761), .Z(n27021) );
  IV U26793 ( .A(p_input[4610]), .Z(n26761) );
  XNOR U26794 ( .A(n27023), .B(n27024), .Z(n27019) );
  AND U26795 ( .A(n27025), .B(n27026), .Z(n27024) );
  XOR U26796 ( .A(p_input[4641]), .B(n27023), .Z(n27026) );
  XNOR U26797 ( .A(p_input[4609]), .B(n27023), .Z(n27025) );
  AND U26798 ( .A(p_input[4640]), .B(n27027), .Z(n27023) );
  IV U26799 ( .A(p_input[4608]), .Z(n27027) );
  XOR U26800 ( .A(n27028), .B(n27029), .Z(n23384) );
  AND U26801 ( .A(n1012), .B(n27030), .Z(n27029) );
  XNOR U26802 ( .A(n27031), .B(n27028), .Z(n27030) );
  XOR U26803 ( .A(n27032), .B(n27033), .Z(n1012) );
  AND U26804 ( .A(n27034), .B(n27035), .Z(n27033) );
  XOR U26805 ( .A(n27032), .B(n23399), .Z(n27035) );
  XOR U26806 ( .A(n27036), .B(n27037), .Z(n23399) );
  AND U26807 ( .A(n859), .B(n27038), .Z(n27037) );
  XOR U26808 ( .A(n27039), .B(n27036), .Z(n27038) );
  XNOR U26809 ( .A(n23396), .B(n27032), .Z(n27034) );
  XOR U26810 ( .A(n27040), .B(n27041), .Z(n23396) );
  AND U26811 ( .A(n856), .B(n27042), .Z(n27041) );
  XOR U26812 ( .A(n27043), .B(n27040), .Z(n27042) );
  XOR U26813 ( .A(n27044), .B(n27045), .Z(n27032) );
  AND U26814 ( .A(n27046), .B(n27047), .Z(n27045) );
  XOR U26815 ( .A(n27044), .B(n23411), .Z(n27047) );
  XOR U26816 ( .A(n27048), .B(n27049), .Z(n23411) );
  AND U26817 ( .A(n859), .B(n27050), .Z(n27049) );
  XOR U26818 ( .A(n27051), .B(n27048), .Z(n27050) );
  XNOR U26819 ( .A(n23408), .B(n27044), .Z(n27046) );
  XOR U26820 ( .A(n27052), .B(n27053), .Z(n23408) );
  AND U26821 ( .A(n856), .B(n27054), .Z(n27053) );
  XOR U26822 ( .A(n27055), .B(n27052), .Z(n27054) );
  XOR U26823 ( .A(n27056), .B(n27057), .Z(n27044) );
  AND U26824 ( .A(n27058), .B(n27059), .Z(n27057) );
  XOR U26825 ( .A(n27056), .B(n23423), .Z(n27059) );
  XOR U26826 ( .A(n27060), .B(n27061), .Z(n23423) );
  AND U26827 ( .A(n859), .B(n27062), .Z(n27061) );
  XOR U26828 ( .A(n27063), .B(n27060), .Z(n27062) );
  XNOR U26829 ( .A(n23420), .B(n27056), .Z(n27058) );
  XOR U26830 ( .A(n27064), .B(n27065), .Z(n23420) );
  AND U26831 ( .A(n856), .B(n27066), .Z(n27065) );
  XOR U26832 ( .A(n27067), .B(n27064), .Z(n27066) );
  XOR U26833 ( .A(n27068), .B(n27069), .Z(n27056) );
  AND U26834 ( .A(n27070), .B(n27071), .Z(n27069) );
  XOR U26835 ( .A(n27068), .B(n23435), .Z(n27071) );
  XOR U26836 ( .A(n27072), .B(n27073), .Z(n23435) );
  AND U26837 ( .A(n859), .B(n27074), .Z(n27073) );
  XOR U26838 ( .A(n27075), .B(n27072), .Z(n27074) );
  XNOR U26839 ( .A(n23432), .B(n27068), .Z(n27070) );
  XOR U26840 ( .A(n27076), .B(n27077), .Z(n23432) );
  AND U26841 ( .A(n856), .B(n27078), .Z(n27077) );
  XOR U26842 ( .A(n27079), .B(n27076), .Z(n27078) );
  XOR U26843 ( .A(n27080), .B(n27081), .Z(n27068) );
  AND U26844 ( .A(n27082), .B(n27083), .Z(n27081) );
  XOR U26845 ( .A(n27080), .B(n23447), .Z(n27083) );
  XOR U26846 ( .A(n27084), .B(n27085), .Z(n23447) );
  AND U26847 ( .A(n859), .B(n27086), .Z(n27085) );
  XOR U26848 ( .A(n27087), .B(n27084), .Z(n27086) );
  XNOR U26849 ( .A(n23444), .B(n27080), .Z(n27082) );
  XOR U26850 ( .A(n27088), .B(n27089), .Z(n23444) );
  AND U26851 ( .A(n856), .B(n27090), .Z(n27089) );
  XOR U26852 ( .A(n27091), .B(n27088), .Z(n27090) );
  XOR U26853 ( .A(n27092), .B(n27093), .Z(n27080) );
  AND U26854 ( .A(n27094), .B(n27095), .Z(n27093) );
  XOR U26855 ( .A(n27092), .B(n23459), .Z(n27095) );
  XOR U26856 ( .A(n27096), .B(n27097), .Z(n23459) );
  AND U26857 ( .A(n859), .B(n27098), .Z(n27097) );
  XOR U26858 ( .A(n27099), .B(n27096), .Z(n27098) );
  XNOR U26859 ( .A(n23456), .B(n27092), .Z(n27094) );
  XOR U26860 ( .A(n27100), .B(n27101), .Z(n23456) );
  AND U26861 ( .A(n856), .B(n27102), .Z(n27101) );
  XOR U26862 ( .A(n27103), .B(n27100), .Z(n27102) );
  XOR U26863 ( .A(n27104), .B(n27105), .Z(n27092) );
  AND U26864 ( .A(n27106), .B(n27107), .Z(n27105) );
  XOR U26865 ( .A(n27104), .B(n23471), .Z(n27107) );
  XOR U26866 ( .A(n27108), .B(n27109), .Z(n23471) );
  AND U26867 ( .A(n859), .B(n27110), .Z(n27109) );
  XOR U26868 ( .A(n27111), .B(n27108), .Z(n27110) );
  XNOR U26869 ( .A(n23468), .B(n27104), .Z(n27106) );
  XOR U26870 ( .A(n27112), .B(n27113), .Z(n23468) );
  AND U26871 ( .A(n856), .B(n27114), .Z(n27113) );
  XOR U26872 ( .A(n27115), .B(n27112), .Z(n27114) );
  XOR U26873 ( .A(n27116), .B(n27117), .Z(n27104) );
  AND U26874 ( .A(n27118), .B(n27119), .Z(n27117) );
  XOR U26875 ( .A(n27116), .B(n23483), .Z(n27119) );
  XOR U26876 ( .A(n27120), .B(n27121), .Z(n23483) );
  AND U26877 ( .A(n859), .B(n27122), .Z(n27121) );
  XOR U26878 ( .A(n27123), .B(n27120), .Z(n27122) );
  XNOR U26879 ( .A(n23480), .B(n27116), .Z(n27118) );
  XOR U26880 ( .A(n27124), .B(n27125), .Z(n23480) );
  AND U26881 ( .A(n856), .B(n27126), .Z(n27125) );
  XOR U26882 ( .A(n27127), .B(n27124), .Z(n27126) );
  XOR U26883 ( .A(n27128), .B(n27129), .Z(n27116) );
  AND U26884 ( .A(n27130), .B(n27131), .Z(n27129) );
  XOR U26885 ( .A(n27128), .B(n23495), .Z(n27131) );
  XOR U26886 ( .A(n27132), .B(n27133), .Z(n23495) );
  AND U26887 ( .A(n859), .B(n27134), .Z(n27133) );
  XOR U26888 ( .A(n27135), .B(n27132), .Z(n27134) );
  XNOR U26889 ( .A(n23492), .B(n27128), .Z(n27130) );
  XOR U26890 ( .A(n27136), .B(n27137), .Z(n23492) );
  AND U26891 ( .A(n856), .B(n27138), .Z(n27137) );
  XOR U26892 ( .A(n27139), .B(n27136), .Z(n27138) );
  XOR U26893 ( .A(n27140), .B(n27141), .Z(n27128) );
  AND U26894 ( .A(n27142), .B(n27143), .Z(n27141) );
  XOR U26895 ( .A(n27140), .B(n23507), .Z(n27143) );
  XOR U26896 ( .A(n27144), .B(n27145), .Z(n23507) );
  AND U26897 ( .A(n859), .B(n27146), .Z(n27145) );
  XOR U26898 ( .A(n27147), .B(n27144), .Z(n27146) );
  XNOR U26899 ( .A(n23504), .B(n27140), .Z(n27142) );
  XOR U26900 ( .A(n27148), .B(n27149), .Z(n23504) );
  AND U26901 ( .A(n856), .B(n27150), .Z(n27149) );
  XOR U26902 ( .A(n27151), .B(n27148), .Z(n27150) );
  XOR U26903 ( .A(n27152), .B(n27153), .Z(n27140) );
  AND U26904 ( .A(n27154), .B(n27155), .Z(n27153) );
  XOR U26905 ( .A(n27152), .B(n23519), .Z(n27155) );
  XOR U26906 ( .A(n27156), .B(n27157), .Z(n23519) );
  AND U26907 ( .A(n859), .B(n27158), .Z(n27157) );
  XOR U26908 ( .A(n27159), .B(n27156), .Z(n27158) );
  XNOR U26909 ( .A(n23516), .B(n27152), .Z(n27154) );
  XOR U26910 ( .A(n27160), .B(n27161), .Z(n23516) );
  AND U26911 ( .A(n856), .B(n27162), .Z(n27161) );
  XOR U26912 ( .A(n27163), .B(n27160), .Z(n27162) );
  XOR U26913 ( .A(n27164), .B(n27165), .Z(n27152) );
  AND U26914 ( .A(n27166), .B(n27167), .Z(n27165) );
  XOR U26915 ( .A(n27164), .B(n23531), .Z(n27167) );
  XOR U26916 ( .A(n27168), .B(n27169), .Z(n23531) );
  AND U26917 ( .A(n859), .B(n27170), .Z(n27169) );
  XOR U26918 ( .A(n27171), .B(n27168), .Z(n27170) );
  XNOR U26919 ( .A(n23528), .B(n27164), .Z(n27166) );
  XOR U26920 ( .A(n27172), .B(n27173), .Z(n23528) );
  AND U26921 ( .A(n856), .B(n27174), .Z(n27173) );
  XOR U26922 ( .A(n27175), .B(n27172), .Z(n27174) );
  XOR U26923 ( .A(n27176), .B(n27177), .Z(n27164) );
  AND U26924 ( .A(n27178), .B(n27179), .Z(n27177) );
  XOR U26925 ( .A(n27176), .B(n23543), .Z(n27179) );
  XOR U26926 ( .A(n27180), .B(n27181), .Z(n23543) );
  AND U26927 ( .A(n859), .B(n27182), .Z(n27181) );
  XOR U26928 ( .A(n27183), .B(n27180), .Z(n27182) );
  XNOR U26929 ( .A(n23540), .B(n27176), .Z(n27178) );
  XOR U26930 ( .A(n27184), .B(n27185), .Z(n23540) );
  AND U26931 ( .A(n856), .B(n27186), .Z(n27185) );
  XOR U26932 ( .A(n27187), .B(n27184), .Z(n27186) );
  XOR U26933 ( .A(n27188), .B(n27189), .Z(n27176) );
  AND U26934 ( .A(n27190), .B(n27191), .Z(n27189) );
  XOR U26935 ( .A(n27188), .B(n23555), .Z(n27191) );
  XOR U26936 ( .A(n27192), .B(n27193), .Z(n23555) );
  AND U26937 ( .A(n859), .B(n27194), .Z(n27193) );
  XOR U26938 ( .A(n27195), .B(n27192), .Z(n27194) );
  XNOR U26939 ( .A(n23552), .B(n27188), .Z(n27190) );
  XOR U26940 ( .A(n27196), .B(n27197), .Z(n23552) );
  AND U26941 ( .A(n856), .B(n27198), .Z(n27197) );
  XOR U26942 ( .A(n27199), .B(n27196), .Z(n27198) );
  XOR U26943 ( .A(n27200), .B(n27201), .Z(n27188) );
  AND U26944 ( .A(n27202), .B(n27203), .Z(n27201) );
  XOR U26945 ( .A(n27200), .B(n23567), .Z(n27203) );
  XOR U26946 ( .A(n27204), .B(n27205), .Z(n23567) );
  AND U26947 ( .A(n859), .B(n27206), .Z(n27205) );
  XOR U26948 ( .A(n27207), .B(n27204), .Z(n27206) );
  XNOR U26949 ( .A(n23564), .B(n27200), .Z(n27202) );
  XOR U26950 ( .A(n27208), .B(n27209), .Z(n23564) );
  AND U26951 ( .A(n856), .B(n27210), .Z(n27209) );
  XOR U26952 ( .A(n27211), .B(n27208), .Z(n27210) );
  XOR U26953 ( .A(n27212), .B(n27213), .Z(n27200) );
  AND U26954 ( .A(n27214), .B(n27215), .Z(n27213) );
  XOR U26955 ( .A(n27212), .B(n23579), .Z(n27215) );
  XOR U26956 ( .A(n27216), .B(n27217), .Z(n23579) );
  AND U26957 ( .A(n859), .B(n27218), .Z(n27217) );
  XOR U26958 ( .A(n27219), .B(n27216), .Z(n27218) );
  XNOR U26959 ( .A(n23576), .B(n27212), .Z(n27214) );
  XOR U26960 ( .A(n27220), .B(n27221), .Z(n23576) );
  AND U26961 ( .A(n856), .B(n27222), .Z(n27221) );
  XOR U26962 ( .A(n27223), .B(n27220), .Z(n27222) );
  XOR U26963 ( .A(n27224), .B(n27225), .Z(n27212) );
  AND U26964 ( .A(n27226), .B(n27227), .Z(n27225) );
  XOR U26965 ( .A(n27224), .B(n23591), .Z(n27227) );
  XOR U26966 ( .A(n27228), .B(n27229), .Z(n23591) );
  AND U26967 ( .A(n859), .B(n27230), .Z(n27229) );
  XOR U26968 ( .A(n27231), .B(n27228), .Z(n27230) );
  XNOR U26969 ( .A(n23588), .B(n27224), .Z(n27226) );
  XOR U26970 ( .A(n27232), .B(n27233), .Z(n23588) );
  AND U26971 ( .A(n856), .B(n27234), .Z(n27233) );
  XOR U26972 ( .A(n27235), .B(n27232), .Z(n27234) );
  XOR U26973 ( .A(n27236), .B(n27237), .Z(n27224) );
  AND U26974 ( .A(n27238), .B(n27239), .Z(n27237) );
  XOR U26975 ( .A(n27236), .B(n23603), .Z(n27239) );
  XOR U26976 ( .A(n27240), .B(n27241), .Z(n23603) );
  AND U26977 ( .A(n859), .B(n27242), .Z(n27241) );
  XOR U26978 ( .A(n27243), .B(n27240), .Z(n27242) );
  XNOR U26979 ( .A(n23600), .B(n27236), .Z(n27238) );
  XOR U26980 ( .A(n27244), .B(n27245), .Z(n23600) );
  AND U26981 ( .A(n856), .B(n27246), .Z(n27245) );
  XOR U26982 ( .A(n27247), .B(n27244), .Z(n27246) );
  XOR U26983 ( .A(n27248), .B(n27249), .Z(n27236) );
  AND U26984 ( .A(n27250), .B(n27251), .Z(n27249) );
  XOR U26985 ( .A(n27248), .B(n23615), .Z(n27251) );
  XOR U26986 ( .A(n27252), .B(n27253), .Z(n23615) );
  AND U26987 ( .A(n859), .B(n27254), .Z(n27253) );
  XOR U26988 ( .A(n27255), .B(n27252), .Z(n27254) );
  XNOR U26989 ( .A(n23612), .B(n27248), .Z(n27250) );
  XOR U26990 ( .A(n27256), .B(n27257), .Z(n23612) );
  AND U26991 ( .A(n856), .B(n27258), .Z(n27257) );
  XOR U26992 ( .A(n27259), .B(n27256), .Z(n27258) );
  XOR U26993 ( .A(n27260), .B(n27261), .Z(n27248) );
  AND U26994 ( .A(n27262), .B(n27263), .Z(n27261) );
  XOR U26995 ( .A(n27260), .B(n23627), .Z(n27263) );
  XOR U26996 ( .A(n27264), .B(n27265), .Z(n23627) );
  AND U26997 ( .A(n859), .B(n27266), .Z(n27265) );
  XOR U26998 ( .A(n27267), .B(n27264), .Z(n27266) );
  XNOR U26999 ( .A(n23624), .B(n27260), .Z(n27262) );
  XOR U27000 ( .A(n27268), .B(n27269), .Z(n23624) );
  AND U27001 ( .A(n856), .B(n27270), .Z(n27269) );
  XOR U27002 ( .A(n27271), .B(n27268), .Z(n27270) );
  XOR U27003 ( .A(n27272), .B(n27273), .Z(n27260) );
  AND U27004 ( .A(n27274), .B(n27275), .Z(n27273) );
  XOR U27005 ( .A(n27272), .B(n23639), .Z(n27275) );
  XOR U27006 ( .A(n27276), .B(n27277), .Z(n23639) );
  AND U27007 ( .A(n859), .B(n27278), .Z(n27277) );
  XOR U27008 ( .A(n27279), .B(n27276), .Z(n27278) );
  XNOR U27009 ( .A(n23636), .B(n27272), .Z(n27274) );
  XOR U27010 ( .A(n27280), .B(n27281), .Z(n23636) );
  AND U27011 ( .A(n856), .B(n27282), .Z(n27281) );
  XOR U27012 ( .A(n27283), .B(n27280), .Z(n27282) );
  XOR U27013 ( .A(n27284), .B(n27285), .Z(n27272) );
  AND U27014 ( .A(n27286), .B(n27287), .Z(n27285) );
  XOR U27015 ( .A(n27284), .B(n23651), .Z(n27287) );
  XOR U27016 ( .A(n27288), .B(n27289), .Z(n23651) );
  AND U27017 ( .A(n859), .B(n27290), .Z(n27289) );
  XOR U27018 ( .A(n27291), .B(n27288), .Z(n27290) );
  XNOR U27019 ( .A(n23648), .B(n27284), .Z(n27286) );
  XOR U27020 ( .A(n27292), .B(n27293), .Z(n23648) );
  AND U27021 ( .A(n856), .B(n27294), .Z(n27293) );
  XOR U27022 ( .A(n27295), .B(n27292), .Z(n27294) );
  XOR U27023 ( .A(n27296), .B(n27297), .Z(n27284) );
  AND U27024 ( .A(n27298), .B(n27299), .Z(n27297) );
  XOR U27025 ( .A(n27296), .B(n23663), .Z(n27299) );
  XOR U27026 ( .A(n27300), .B(n27301), .Z(n23663) );
  AND U27027 ( .A(n859), .B(n27302), .Z(n27301) );
  XOR U27028 ( .A(n27303), .B(n27300), .Z(n27302) );
  XNOR U27029 ( .A(n23660), .B(n27296), .Z(n27298) );
  XOR U27030 ( .A(n27304), .B(n27305), .Z(n23660) );
  AND U27031 ( .A(n856), .B(n27306), .Z(n27305) );
  XOR U27032 ( .A(n27307), .B(n27304), .Z(n27306) );
  XOR U27033 ( .A(n27308), .B(n27309), .Z(n27296) );
  AND U27034 ( .A(n27310), .B(n27311), .Z(n27309) );
  XOR U27035 ( .A(n27308), .B(n23675), .Z(n27311) );
  XOR U27036 ( .A(n27312), .B(n27313), .Z(n23675) );
  AND U27037 ( .A(n859), .B(n27314), .Z(n27313) );
  XOR U27038 ( .A(n27315), .B(n27312), .Z(n27314) );
  XNOR U27039 ( .A(n23672), .B(n27308), .Z(n27310) );
  XOR U27040 ( .A(n27316), .B(n27317), .Z(n23672) );
  AND U27041 ( .A(n856), .B(n27318), .Z(n27317) );
  XOR U27042 ( .A(n27319), .B(n27316), .Z(n27318) );
  XOR U27043 ( .A(n27320), .B(n27321), .Z(n27308) );
  AND U27044 ( .A(n27322), .B(n27323), .Z(n27321) );
  XOR U27045 ( .A(n27320), .B(n23687), .Z(n27323) );
  XOR U27046 ( .A(n27324), .B(n27325), .Z(n23687) );
  AND U27047 ( .A(n859), .B(n27326), .Z(n27325) );
  XOR U27048 ( .A(n27327), .B(n27324), .Z(n27326) );
  XNOR U27049 ( .A(n23684), .B(n27320), .Z(n27322) );
  XOR U27050 ( .A(n27328), .B(n27329), .Z(n23684) );
  AND U27051 ( .A(n856), .B(n27330), .Z(n27329) );
  XOR U27052 ( .A(n27331), .B(n27328), .Z(n27330) );
  XOR U27053 ( .A(n27332), .B(n27333), .Z(n27320) );
  AND U27054 ( .A(n27334), .B(n27335), .Z(n27333) );
  XOR U27055 ( .A(n27332), .B(n23699), .Z(n27335) );
  XOR U27056 ( .A(n27336), .B(n27337), .Z(n23699) );
  AND U27057 ( .A(n859), .B(n27338), .Z(n27337) );
  XOR U27058 ( .A(n27339), .B(n27336), .Z(n27338) );
  XNOR U27059 ( .A(n23696), .B(n27332), .Z(n27334) );
  XOR U27060 ( .A(n27340), .B(n27341), .Z(n23696) );
  AND U27061 ( .A(n856), .B(n27342), .Z(n27341) );
  XOR U27062 ( .A(n27343), .B(n27340), .Z(n27342) );
  XOR U27063 ( .A(n27344), .B(n27345), .Z(n27332) );
  AND U27064 ( .A(n27346), .B(n27347), .Z(n27345) );
  XOR U27065 ( .A(n27344), .B(n23711), .Z(n27347) );
  XOR U27066 ( .A(n27348), .B(n27349), .Z(n23711) );
  AND U27067 ( .A(n859), .B(n27350), .Z(n27349) );
  XOR U27068 ( .A(n27351), .B(n27348), .Z(n27350) );
  XNOR U27069 ( .A(n23708), .B(n27344), .Z(n27346) );
  XOR U27070 ( .A(n27352), .B(n27353), .Z(n23708) );
  AND U27071 ( .A(n856), .B(n27354), .Z(n27353) );
  XOR U27072 ( .A(n27355), .B(n27352), .Z(n27354) );
  XOR U27073 ( .A(n27356), .B(n27357), .Z(n27344) );
  AND U27074 ( .A(n27358), .B(n27359), .Z(n27357) );
  XOR U27075 ( .A(n27356), .B(n23723), .Z(n27359) );
  XOR U27076 ( .A(n27360), .B(n27361), .Z(n23723) );
  AND U27077 ( .A(n859), .B(n27362), .Z(n27361) );
  XOR U27078 ( .A(n27363), .B(n27360), .Z(n27362) );
  XNOR U27079 ( .A(n23720), .B(n27356), .Z(n27358) );
  XOR U27080 ( .A(n27364), .B(n27365), .Z(n23720) );
  AND U27081 ( .A(n856), .B(n27366), .Z(n27365) );
  XOR U27082 ( .A(n27367), .B(n27364), .Z(n27366) );
  XOR U27083 ( .A(n27368), .B(n27369), .Z(n27356) );
  AND U27084 ( .A(n27370), .B(n27371), .Z(n27369) );
  XOR U27085 ( .A(n27368), .B(n23735), .Z(n27371) );
  XOR U27086 ( .A(n27372), .B(n27373), .Z(n23735) );
  AND U27087 ( .A(n859), .B(n27374), .Z(n27373) );
  XOR U27088 ( .A(n27375), .B(n27372), .Z(n27374) );
  XNOR U27089 ( .A(n23732), .B(n27368), .Z(n27370) );
  XOR U27090 ( .A(n27376), .B(n27377), .Z(n23732) );
  AND U27091 ( .A(n856), .B(n27378), .Z(n27377) );
  XOR U27092 ( .A(n27379), .B(n27376), .Z(n27378) );
  XOR U27093 ( .A(n27380), .B(n27381), .Z(n27368) );
  AND U27094 ( .A(n27382), .B(n27383), .Z(n27381) );
  XOR U27095 ( .A(n27380), .B(n23747), .Z(n27383) );
  XOR U27096 ( .A(n27384), .B(n27385), .Z(n23747) );
  AND U27097 ( .A(n859), .B(n27386), .Z(n27385) );
  XOR U27098 ( .A(n27387), .B(n27384), .Z(n27386) );
  XNOR U27099 ( .A(n23744), .B(n27380), .Z(n27382) );
  XOR U27100 ( .A(n27388), .B(n27389), .Z(n23744) );
  AND U27101 ( .A(n856), .B(n27390), .Z(n27389) );
  XOR U27102 ( .A(n27391), .B(n27388), .Z(n27390) );
  XOR U27103 ( .A(n27392), .B(n27393), .Z(n27380) );
  AND U27104 ( .A(n27394), .B(n27395), .Z(n27393) );
  XNOR U27105 ( .A(n27396), .B(n23760), .Z(n27395) );
  XOR U27106 ( .A(n27397), .B(n27398), .Z(n23760) );
  AND U27107 ( .A(n859), .B(n27399), .Z(n27398) );
  XOR U27108 ( .A(n27397), .B(n27400), .Z(n27399) );
  XNOR U27109 ( .A(n23757), .B(n27392), .Z(n27394) );
  XOR U27110 ( .A(n27401), .B(n27402), .Z(n23757) );
  AND U27111 ( .A(n856), .B(n27403), .Z(n27402) );
  XOR U27112 ( .A(n27401), .B(n27404), .Z(n27403) );
  IV U27113 ( .A(n27396), .Z(n27392) );
  AND U27114 ( .A(n27028), .B(n27031), .Z(n27396) );
  XNOR U27115 ( .A(n27405), .B(n27406), .Z(n27031) );
  AND U27116 ( .A(n859), .B(n27407), .Z(n27406) );
  XNOR U27117 ( .A(n27408), .B(n27405), .Z(n27407) );
  XOR U27118 ( .A(n27409), .B(n27410), .Z(n859) );
  AND U27119 ( .A(n27411), .B(n27412), .Z(n27410) );
  XOR U27120 ( .A(n27409), .B(n27039), .Z(n27412) );
  XNOR U27121 ( .A(n27413), .B(n27414), .Z(n27039) );
  AND U27122 ( .A(n27415), .B(n539), .Z(n27414) );
  AND U27123 ( .A(n27413), .B(n27416), .Z(n27415) );
  XNOR U27124 ( .A(n27036), .B(n27409), .Z(n27411) );
  XOR U27125 ( .A(n27417), .B(n27418), .Z(n27036) );
  AND U27126 ( .A(n27419), .B(n537), .Z(n27418) );
  NOR U27127 ( .A(n27417), .B(n27420), .Z(n27419) );
  XOR U27128 ( .A(n27421), .B(n27422), .Z(n27409) );
  AND U27129 ( .A(n27423), .B(n27424), .Z(n27422) );
  XOR U27130 ( .A(n27421), .B(n27051), .Z(n27424) );
  XOR U27131 ( .A(n27425), .B(n27426), .Z(n27051) );
  AND U27132 ( .A(n539), .B(n27427), .Z(n27426) );
  XOR U27133 ( .A(n27428), .B(n27425), .Z(n27427) );
  XNOR U27134 ( .A(n27048), .B(n27421), .Z(n27423) );
  XOR U27135 ( .A(n27429), .B(n27430), .Z(n27048) );
  AND U27136 ( .A(n537), .B(n27431), .Z(n27430) );
  XOR U27137 ( .A(n27432), .B(n27429), .Z(n27431) );
  XOR U27138 ( .A(n27433), .B(n27434), .Z(n27421) );
  AND U27139 ( .A(n27435), .B(n27436), .Z(n27434) );
  XOR U27140 ( .A(n27433), .B(n27063), .Z(n27436) );
  XOR U27141 ( .A(n27437), .B(n27438), .Z(n27063) );
  AND U27142 ( .A(n539), .B(n27439), .Z(n27438) );
  XOR U27143 ( .A(n27440), .B(n27437), .Z(n27439) );
  XNOR U27144 ( .A(n27060), .B(n27433), .Z(n27435) );
  XOR U27145 ( .A(n27441), .B(n27442), .Z(n27060) );
  AND U27146 ( .A(n537), .B(n27443), .Z(n27442) );
  XOR U27147 ( .A(n27444), .B(n27441), .Z(n27443) );
  XOR U27148 ( .A(n27445), .B(n27446), .Z(n27433) );
  AND U27149 ( .A(n27447), .B(n27448), .Z(n27446) );
  XOR U27150 ( .A(n27445), .B(n27075), .Z(n27448) );
  XOR U27151 ( .A(n27449), .B(n27450), .Z(n27075) );
  AND U27152 ( .A(n539), .B(n27451), .Z(n27450) );
  XOR U27153 ( .A(n27452), .B(n27449), .Z(n27451) );
  XNOR U27154 ( .A(n27072), .B(n27445), .Z(n27447) );
  XOR U27155 ( .A(n27453), .B(n27454), .Z(n27072) );
  AND U27156 ( .A(n537), .B(n27455), .Z(n27454) );
  XOR U27157 ( .A(n27456), .B(n27453), .Z(n27455) );
  XOR U27158 ( .A(n27457), .B(n27458), .Z(n27445) );
  AND U27159 ( .A(n27459), .B(n27460), .Z(n27458) );
  XOR U27160 ( .A(n27457), .B(n27087), .Z(n27460) );
  XOR U27161 ( .A(n27461), .B(n27462), .Z(n27087) );
  AND U27162 ( .A(n539), .B(n27463), .Z(n27462) );
  XOR U27163 ( .A(n27464), .B(n27461), .Z(n27463) );
  XNOR U27164 ( .A(n27084), .B(n27457), .Z(n27459) );
  XOR U27165 ( .A(n27465), .B(n27466), .Z(n27084) );
  AND U27166 ( .A(n537), .B(n27467), .Z(n27466) );
  XOR U27167 ( .A(n27468), .B(n27465), .Z(n27467) );
  XOR U27168 ( .A(n27469), .B(n27470), .Z(n27457) );
  AND U27169 ( .A(n27471), .B(n27472), .Z(n27470) );
  XOR U27170 ( .A(n27469), .B(n27099), .Z(n27472) );
  XOR U27171 ( .A(n27473), .B(n27474), .Z(n27099) );
  AND U27172 ( .A(n539), .B(n27475), .Z(n27474) );
  XOR U27173 ( .A(n27476), .B(n27473), .Z(n27475) );
  XNOR U27174 ( .A(n27096), .B(n27469), .Z(n27471) );
  XOR U27175 ( .A(n27477), .B(n27478), .Z(n27096) );
  AND U27176 ( .A(n537), .B(n27479), .Z(n27478) );
  XOR U27177 ( .A(n27480), .B(n27477), .Z(n27479) );
  XOR U27178 ( .A(n27481), .B(n27482), .Z(n27469) );
  AND U27179 ( .A(n27483), .B(n27484), .Z(n27482) );
  XOR U27180 ( .A(n27481), .B(n27111), .Z(n27484) );
  XOR U27181 ( .A(n27485), .B(n27486), .Z(n27111) );
  AND U27182 ( .A(n539), .B(n27487), .Z(n27486) );
  XOR U27183 ( .A(n27488), .B(n27485), .Z(n27487) );
  XNOR U27184 ( .A(n27108), .B(n27481), .Z(n27483) );
  XOR U27185 ( .A(n27489), .B(n27490), .Z(n27108) );
  AND U27186 ( .A(n537), .B(n27491), .Z(n27490) );
  XOR U27187 ( .A(n27492), .B(n27489), .Z(n27491) );
  XOR U27188 ( .A(n27493), .B(n27494), .Z(n27481) );
  AND U27189 ( .A(n27495), .B(n27496), .Z(n27494) );
  XOR U27190 ( .A(n27493), .B(n27123), .Z(n27496) );
  XOR U27191 ( .A(n27497), .B(n27498), .Z(n27123) );
  AND U27192 ( .A(n539), .B(n27499), .Z(n27498) );
  XOR U27193 ( .A(n27500), .B(n27497), .Z(n27499) );
  XNOR U27194 ( .A(n27120), .B(n27493), .Z(n27495) );
  XOR U27195 ( .A(n27501), .B(n27502), .Z(n27120) );
  AND U27196 ( .A(n537), .B(n27503), .Z(n27502) );
  XOR U27197 ( .A(n27504), .B(n27501), .Z(n27503) );
  XOR U27198 ( .A(n27505), .B(n27506), .Z(n27493) );
  AND U27199 ( .A(n27507), .B(n27508), .Z(n27506) );
  XOR U27200 ( .A(n27505), .B(n27135), .Z(n27508) );
  XOR U27201 ( .A(n27509), .B(n27510), .Z(n27135) );
  AND U27202 ( .A(n539), .B(n27511), .Z(n27510) );
  XOR U27203 ( .A(n27512), .B(n27509), .Z(n27511) );
  XNOR U27204 ( .A(n27132), .B(n27505), .Z(n27507) );
  XOR U27205 ( .A(n27513), .B(n27514), .Z(n27132) );
  AND U27206 ( .A(n537), .B(n27515), .Z(n27514) );
  XOR U27207 ( .A(n27516), .B(n27513), .Z(n27515) );
  XOR U27208 ( .A(n27517), .B(n27518), .Z(n27505) );
  AND U27209 ( .A(n27519), .B(n27520), .Z(n27518) );
  XOR U27210 ( .A(n27517), .B(n27147), .Z(n27520) );
  XOR U27211 ( .A(n27521), .B(n27522), .Z(n27147) );
  AND U27212 ( .A(n539), .B(n27523), .Z(n27522) );
  XOR U27213 ( .A(n27524), .B(n27521), .Z(n27523) );
  XNOR U27214 ( .A(n27144), .B(n27517), .Z(n27519) );
  XOR U27215 ( .A(n27525), .B(n27526), .Z(n27144) );
  AND U27216 ( .A(n537), .B(n27527), .Z(n27526) );
  XOR U27217 ( .A(n27528), .B(n27525), .Z(n27527) );
  XOR U27218 ( .A(n27529), .B(n27530), .Z(n27517) );
  AND U27219 ( .A(n27531), .B(n27532), .Z(n27530) );
  XOR U27220 ( .A(n27529), .B(n27159), .Z(n27532) );
  XOR U27221 ( .A(n27533), .B(n27534), .Z(n27159) );
  AND U27222 ( .A(n539), .B(n27535), .Z(n27534) );
  XOR U27223 ( .A(n27536), .B(n27533), .Z(n27535) );
  XNOR U27224 ( .A(n27156), .B(n27529), .Z(n27531) );
  XOR U27225 ( .A(n27537), .B(n27538), .Z(n27156) );
  AND U27226 ( .A(n537), .B(n27539), .Z(n27538) );
  XOR U27227 ( .A(n27540), .B(n27537), .Z(n27539) );
  XOR U27228 ( .A(n27541), .B(n27542), .Z(n27529) );
  AND U27229 ( .A(n27543), .B(n27544), .Z(n27542) );
  XOR U27230 ( .A(n27541), .B(n27171), .Z(n27544) );
  XOR U27231 ( .A(n27545), .B(n27546), .Z(n27171) );
  AND U27232 ( .A(n539), .B(n27547), .Z(n27546) );
  XOR U27233 ( .A(n27548), .B(n27545), .Z(n27547) );
  XNOR U27234 ( .A(n27168), .B(n27541), .Z(n27543) );
  XOR U27235 ( .A(n27549), .B(n27550), .Z(n27168) );
  AND U27236 ( .A(n537), .B(n27551), .Z(n27550) );
  XOR U27237 ( .A(n27552), .B(n27549), .Z(n27551) );
  XOR U27238 ( .A(n27553), .B(n27554), .Z(n27541) );
  AND U27239 ( .A(n27555), .B(n27556), .Z(n27554) );
  XOR U27240 ( .A(n27553), .B(n27183), .Z(n27556) );
  XOR U27241 ( .A(n27557), .B(n27558), .Z(n27183) );
  AND U27242 ( .A(n539), .B(n27559), .Z(n27558) );
  XOR U27243 ( .A(n27560), .B(n27557), .Z(n27559) );
  XNOR U27244 ( .A(n27180), .B(n27553), .Z(n27555) );
  XOR U27245 ( .A(n27561), .B(n27562), .Z(n27180) );
  AND U27246 ( .A(n537), .B(n27563), .Z(n27562) );
  XOR U27247 ( .A(n27564), .B(n27561), .Z(n27563) );
  XOR U27248 ( .A(n27565), .B(n27566), .Z(n27553) );
  AND U27249 ( .A(n27567), .B(n27568), .Z(n27566) );
  XOR U27250 ( .A(n27565), .B(n27195), .Z(n27568) );
  XOR U27251 ( .A(n27569), .B(n27570), .Z(n27195) );
  AND U27252 ( .A(n539), .B(n27571), .Z(n27570) );
  XOR U27253 ( .A(n27572), .B(n27569), .Z(n27571) );
  XNOR U27254 ( .A(n27192), .B(n27565), .Z(n27567) );
  XOR U27255 ( .A(n27573), .B(n27574), .Z(n27192) );
  AND U27256 ( .A(n537), .B(n27575), .Z(n27574) );
  XOR U27257 ( .A(n27576), .B(n27573), .Z(n27575) );
  XOR U27258 ( .A(n27577), .B(n27578), .Z(n27565) );
  AND U27259 ( .A(n27579), .B(n27580), .Z(n27578) );
  XOR U27260 ( .A(n27577), .B(n27207), .Z(n27580) );
  XOR U27261 ( .A(n27581), .B(n27582), .Z(n27207) );
  AND U27262 ( .A(n539), .B(n27583), .Z(n27582) );
  XOR U27263 ( .A(n27584), .B(n27581), .Z(n27583) );
  XNOR U27264 ( .A(n27204), .B(n27577), .Z(n27579) );
  XOR U27265 ( .A(n27585), .B(n27586), .Z(n27204) );
  AND U27266 ( .A(n537), .B(n27587), .Z(n27586) );
  XOR U27267 ( .A(n27588), .B(n27585), .Z(n27587) );
  XOR U27268 ( .A(n27589), .B(n27590), .Z(n27577) );
  AND U27269 ( .A(n27591), .B(n27592), .Z(n27590) );
  XOR U27270 ( .A(n27589), .B(n27219), .Z(n27592) );
  XOR U27271 ( .A(n27593), .B(n27594), .Z(n27219) );
  AND U27272 ( .A(n539), .B(n27595), .Z(n27594) );
  XOR U27273 ( .A(n27596), .B(n27593), .Z(n27595) );
  XNOR U27274 ( .A(n27216), .B(n27589), .Z(n27591) );
  XOR U27275 ( .A(n27597), .B(n27598), .Z(n27216) );
  AND U27276 ( .A(n537), .B(n27599), .Z(n27598) );
  XOR U27277 ( .A(n27600), .B(n27597), .Z(n27599) );
  XOR U27278 ( .A(n27601), .B(n27602), .Z(n27589) );
  AND U27279 ( .A(n27603), .B(n27604), .Z(n27602) );
  XOR U27280 ( .A(n27601), .B(n27231), .Z(n27604) );
  XOR U27281 ( .A(n27605), .B(n27606), .Z(n27231) );
  AND U27282 ( .A(n539), .B(n27607), .Z(n27606) );
  XOR U27283 ( .A(n27608), .B(n27605), .Z(n27607) );
  XNOR U27284 ( .A(n27228), .B(n27601), .Z(n27603) );
  XOR U27285 ( .A(n27609), .B(n27610), .Z(n27228) );
  AND U27286 ( .A(n537), .B(n27611), .Z(n27610) );
  XOR U27287 ( .A(n27612), .B(n27609), .Z(n27611) );
  XOR U27288 ( .A(n27613), .B(n27614), .Z(n27601) );
  AND U27289 ( .A(n27615), .B(n27616), .Z(n27614) );
  XOR U27290 ( .A(n27613), .B(n27243), .Z(n27616) );
  XOR U27291 ( .A(n27617), .B(n27618), .Z(n27243) );
  AND U27292 ( .A(n539), .B(n27619), .Z(n27618) );
  XOR U27293 ( .A(n27620), .B(n27617), .Z(n27619) );
  XNOR U27294 ( .A(n27240), .B(n27613), .Z(n27615) );
  XOR U27295 ( .A(n27621), .B(n27622), .Z(n27240) );
  AND U27296 ( .A(n537), .B(n27623), .Z(n27622) );
  XOR U27297 ( .A(n27624), .B(n27621), .Z(n27623) );
  XOR U27298 ( .A(n27625), .B(n27626), .Z(n27613) );
  AND U27299 ( .A(n27627), .B(n27628), .Z(n27626) );
  XOR U27300 ( .A(n27625), .B(n27255), .Z(n27628) );
  XOR U27301 ( .A(n27629), .B(n27630), .Z(n27255) );
  AND U27302 ( .A(n539), .B(n27631), .Z(n27630) );
  XOR U27303 ( .A(n27632), .B(n27629), .Z(n27631) );
  XNOR U27304 ( .A(n27252), .B(n27625), .Z(n27627) );
  XOR U27305 ( .A(n27633), .B(n27634), .Z(n27252) );
  AND U27306 ( .A(n537), .B(n27635), .Z(n27634) );
  XOR U27307 ( .A(n27636), .B(n27633), .Z(n27635) );
  XOR U27308 ( .A(n27637), .B(n27638), .Z(n27625) );
  AND U27309 ( .A(n27639), .B(n27640), .Z(n27638) );
  XOR U27310 ( .A(n27637), .B(n27267), .Z(n27640) );
  XOR U27311 ( .A(n27641), .B(n27642), .Z(n27267) );
  AND U27312 ( .A(n539), .B(n27643), .Z(n27642) );
  XOR U27313 ( .A(n27644), .B(n27641), .Z(n27643) );
  XNOR U27314 ( .A(n27264), .B(n27637), .Z(n27639) );
  XOR U27315 ( .A(n27645), .B(n27646), .Z(n27264) );
  AND U27316 ( .A(n537), .B(n27647), .Z(n27646) );
  XOR U27317 ( .A(n27648), .B(n27645), .Z(n27647) );
  XOR U27318 ( .A(n27649), .B(n27650), .Z(n27637) );
  AND U27319 ( .A(n27651), .B(n27652), .Z(n27650) );
  XOR U27320 ( .A(n27649), .B(n27279), .Z(n27652) );
  XOR U27321 ( .A(n27653), .B(n27654), .Z(n27279) );
  AND U27322 ( .A(n539), .B(n27655), .Z(n27654) );
  XOR U27323 ( .A(n27656), .B(n27653), .Z(n27655) );
  XNOR U27324 ( .A(n27276), .B(n27649), .Z(n27651) );
  XOR U27325 ( .A(n27657), .B(n27658), .Z(n27276) );
  AND U27326 ( .A(n537), .B(n27659), .Z(n27658) );
  XOR U27327 ( .A(n27660), .B(n27657), .Z(n27659) );
  XOR U27328 ( .A(n27661), .B(n27662), .Z(n27649) );
  AND U27329 ( .A(n27663), .B(n27664), .Z(n27662) );
  XOR U27330 ( .A(n27661), .B(n27291), .Z(n27664) );
  XOR U27331 ( .A(n27665), .B(n27666), .Z(n27291) );
  AND U27332 ( .A(n539), .B(n27667), .Z(n27666) );
  XOR U27333 ( .A(n27668), .B(n27665), .Z(n27667) );
  XNOR U27334 ( .A(n27288), .B(n27661), .Z(n27663) );
  XOR U27335 ( .A(n27669), .B(n27670), .Z(n27288) );
  AND U27336 ( .A(n537), .B(n27671), .Z(n27670) );
  XOR U27337 ( .A(n27672), .B(n27669), .Z(n27671) );
  XOR U27338 ( .A(n27673), .B(n27674), .Z(n27661) );
  AND U27339 ( .A(n27675), .B(n27676), .Z(n27674) );
  XOR U27340 ( .A(n27673), .B(n27303), .Z(n27676) );
  XOR U27341 ( .A(n27677), .B(n27678), .Z(n27303) );
  AND U27342 ( .A(n539), .B(n27679), .Z(n27678) );
  XOR U27343 ( .A(n27680), .B(n27677), .Z(n27679) );
  XNOR U27344 ( .A(n27300), .B(n27673), .Z(n27675) );
  XOR U27345 ( .A(n27681), .B(n27682), .Z(n27300) );
  AND U27346 ( .A(n537), .B(n27683), .Z(n27682) );
  XOR U27347 ( .A(n27684), .B(n27681), .Z(n27683) );
  XOR U27348 ( .A(n27685), .B(n27686), .Z(n27673) );
  AND U27349 ( .A(n27687), .B(n27688), .Z(n27686) );
  XOR U27350 ( .A(n27685), .B(n27315), .Z(n27688) );
  XOR U27351 ( .A(n27689), .B(n27690), .Z(n27315) );
  AND U27352 ( .A(n539), .B(n27691), .Z(n27690) );
  XOR U27353 ( .A(n27692), .B(n27689), .Z(n27691) );
  XNOR U27354 ( .A(n27312), .B(n27685), .Z(n27687) );
  XOR U27355 ( .A(n27693), .B(n27694), .Z(n27312) );
  AND U27356 ( .A(n537), .B(n27695), .Z(n27694) );
  XOR U27357 ( .A(n27696), .B(n27693), .Z(n27695) );
  XOR U27358 ( .A(n27697), .B(n27698), .Z(n27685) );
  AND U27359 ( .A(n27699), .B(n27700), .Z(n27698) );
  XOR U27360 ( .A(n27697), .B(n27327), .Z(n27700) );
  XOR U27361 ( .A(n27701), .B(n27702), .Z(n27327) );
  AND U27362 ( .A(n539), .B(n27703), .Z(n27702) );
  XOR U27363 ( .A(n27704), .B(n27701), .Z(n27703) );
  XNOR U27364 ( .A(n27324), .B(n27697), .Z(n27699) );
  XOR U27365 ( .A(n27705), .B(n27706), .Z(n27324) );
  AND U27366 ( .A(n537), .B(n27707), .Z(n27706) );
  XOR U27367 ( .A(n27708), .B(n27705), .Z(n27707) );
  XOR U27368 ( .A(n27709), .B(n27710), .Z(n27697) );
  AND U27369 ( .A(n27711), .B(n27712), .Z(n27710) );
  XOR U27370 ( .A(n27709), .B(n27339), .Z(n27712) );
  XOR U27371 ( .A(n27713), .B(n27714), .Z(n27339) );
  AND U27372 ( .A(n539), .B(n27715), .Z(n27714) );
  XOR U27373 ( .A(n27716), .B(n27713), .Z(n27715) );
  XNOR U27374 ( .A(n27336), .B(n27709), .Z(n27711) );
  XOR U27375 ( .A(n27717), .B(n27718), .Z(n27336) );
  AND U27376 ( .A(n537), .B(n27719), .Z(n27718) );
  XOR U27377 ( .A(n27720), .B(n27717), .Z(n27719) );
  XOR U27378 ( .A(n27721), .B(n27722), .Z(n27709) );
  AND U27379 ( .A(n27723), .B(n27724), .Z(n27722) );
  XOR U27380 ( .A(n27721), .B(n27351), .Z(n27724) );
  XOR U27381 ( .A(n27725), .B(n27726), .Z(n27351) );
  AND U27382 ( .A(n539), .B(n27727), .Z(n27726) );
  XOR U27383 ( .A(n27728), .B(n27725), .Z(n27727) );
  XNOR U27384 ( .A(n27348), .B(n27721), .Z(n27723) );
  XOR U27385 ( .A(n27729), .B(n27730), .Z(n27348) );
  AND U27386 ( .A(n537), .B(n27731), .Z(n27730) );
  XOR U27387 ( .A(n27732), .B(n27729), .Z(n27731) );
  XOR U27388 ( .A(n27733), .B(n27734), .Z(n27721) );
  AND U27389 ( .A(n27735), .B(n27736), .Z(n27734) );
  XOR U27390 ( .A(n27733), .B(n27363), .Z(n27736) );
  XOR U27391 ( .A(n27737), .B(n27738), .Z(n27363) );
  AND U27392 ( .A(n539), .B(n27739), .Z(n27738) );
  XOR U27393 ( .A(n27740), .B(n27737), .Z(n27739) );
  XNOR U27394 ( .A(n27360), .B(n27733), .Z(n27735) );
  XOR U27395 ( .A(n27741), .B(n27742), .Z(n27360) );
  AND U27396 ( .A(n537), .B(n27743), .Z(n27742) );
  XOR U27397 ( .A(n27744), .B(n27741), .Z(n27743) );
  XOR U27398 ( .A(n27745), .B(n27746), .Z(n27733) );
  AND U27399 ( .A(n27747), .B(n27748), .Z(n27746) );
  XOR U27400 ( .A(n27745), .B(n27375), .Z(n27748) );
  XOR U27401 ( .A(n27749), .B(n27750), .Z(n27375) );
  AND U27402 ( .A(n539), .B(n27751), .Z(n27750) );
  XOR U27403 ( .A(n27752), .B(n27749), .Z(n27751) );
  XNOR U27404 ( .A(n27372), .B(n27745), .Z(n27747) );
  XOR U27405 ( .A(n27753), .B(n27754), .Z(n27372) );
  AND U27406 ( .A(n537), .B(n27755), .Z(n27754) );
  XOR U27407 ( .A(n27756), .B(n27753), .Z(n27755) );
  XOR U27408 ( .A(n27757), .B(n27758), .Z(n27745) );
  AND U27409 ( .A(n27759), .B(n27760), .Z(n27758) );
  XOR U27410 ( .A(n27757), .B(n27387), .Z(n27760) );
  XOR U27411 ( .A(n27761), .B(n27762), .Z(n27387) );
  AND U27412 ( .A(n539), .B(n27763), .Z(n27762) );
  XOR U27413 ( .A(n27764), .B(n27761), .Z(n27763) );
  XNOR U27414 ( .A(n27384), .B(n27757), .Z(n27759) );
  XOR U27415 ( .A(n27765), .B(n27766), .Z(n27384) );
  AND U27416 ( .A(n537), .B(n27767), .Z(n27766) );
  XOR U27417 ( .A(n27768), .B(n27765), .Z(n27767) );
  XOR U27418 ( .A(n27769), .B(n27770), .Z(n27757) );
  AND U27419 ( .A(n27771), .B(n27772), .Z(n27770) );
  XNOR U27420 ( .A(n27773), .B(n27400), .Z(n27772) );
  XOR U27421 ( .A(n27774), .B(n27775), .Z(n27400) );
  AND U27422 ( .A(n539), .B(n27776), .Z(n27775) );
  XOR U27423 ( .A(n27774), .B(n27777), .Z(n27776) );
  XNOR U27424 ( .A(n27397), .B(n27769), .Z(n27771) );
  XOR U27425 ( .A(n27778), .B(n27779), .Z(n27397) );
  AND U27426 ( .A(n537), .B(n27780), .Z(n27779) );
  XOR U27427 ( .A(n27778), .B(n27781), .Z(n27780) );
  IV U27428 ( .A(n27773), .Z(n27769) );
  AND U27429 ( .A(n27405), .B(n27408), .Z(n27773) );
  XNOR U27430 ( .A(n27782), .B(n27783), .Z(n27408) );
  AND U27431 ( .A(n539), .B(n27784), .Z(n27783) );
  XNOR U27432 ( .A(n27785), .B(n27782), .Z(n27784) );
  XOR U27433 ( .A(n27786), .B(n27787), .Z(n539) );
  AND U27434 ( .A(n27788), .B(n27789), .Z(n27787) );
  XOR U27435 ( .A(n27416), .B(n27786), .Z(n27789) );
  IV U27436 ( .A(n27790), .Z(n27416) );
  AND U27437 ( .A(p_input[4607]), .B(p_input[4575]), .Z(n27790) );
  XOR U27438 ( .A(n27786), .B(n27413), .Z(n27788) );
  AND U27439 ( .A(p_input[4511]), .B(p_input[4543]), .Z(n27413) );
  XOR U27440 ( .A(n27791), .B(n27792), .Z(n27786) );
  AND U27441 ( .A(n27793), .B(n27794), .Z(n27792) );
  XOR U27442 ( .A(n27791), .B(n27428), .Z(n27794) );
  XNOR U27443 ( .A(p_input[4574]), .B(n27795), .Z(n27428) );
  AND U27444 ( .A(n399), .B(n27796), .Z(n27795) );
  XOR U27445 ( .A(p_input[4606]), .B(p_input[4574]), .Z(n27796) );
  XNOR U27446 ( .A(n27425), .B(n27791), .Z(n27793) );
  XOR U27447 ( .A(n27797), .B(n27798), .Z(n27425) );
  AND U27448 ( .A(n397), .B(n27799), .Z(n27798) );
  XOR U27449 ( .A(p_input[4542]), .B(p_input[4510]), .Z(n27799) );
  XOR U27450 ( .A(n27800), .B(n27801), .Z(n27791) );
  AND U27451 ( .A(n27802), .B(n27803), .Z(n27801) );
  XOR U27452 ( .A(n27800), .B(n27440), .Z(n27803) );
  XNOR U27453 ( .A(p_input[4573]), .B(n27804), .Z(n27440) );
  AND U27454 ( .A(n399), .B(n27805), .Z(n27804) );
  XOR U27455 ( .A(p_input[4605]), .B(p_input[4573]), .Z(n27805) );
  XNOR U27456 ( .A(n27437), .B(n27800), .Z(n27802) );
  XOR U27457 ( .A(n27806), .B(n27807), .Z(n27437) );
  AND U27458 ( .A(n397), .B(n27808), .Z(n27807) );
  XOR U27459 ( .A(p_input[4541]), .B(p_input[4509]), .Z(n27808) );
  XOR U27460 ( .A(n27809), .B(n27810), .Z(n27800) );
  AND U27461 ( .A(n27811), .B(n27812), .Z(n27810) );
  XOR U27462 ( .A(n27809), .B(n27452), .Z(n27812) );
  XNOR U27463 ( .A(p_input[4572]), .B(n27813), .Z(n27452) );
  AND U27464 ( .A(n399), .B(n27814), .Z(n27813) );
  XOR U27465 ( .A(p_input[4604]), .B(p_input[4572]), .Z(n27814) );
  XNOR U27466 ( .A(n27449), .B(n27809), .Z(n27811) );
  XOR U27467 ( .A(n27815), .B(n27816), .Z(n27449) );
  AND U27468 ( .A(n397), .B(n27817), .Z(n27816) );
  XOR U27469 ( .A(p_input[4540]), .B(p_input[4508]), .Z(n27817) );
  XOR U27470 ( .A(n27818), .B(n27819), .Z(n27809) );
  AND U27471 ( .A(n27820), .B(n27821), .Z(n27819) );
  XOR U27472 ( .A(n27818), .B(n27464), .Z(n27821) );
  XNOR U27473 ( .A(p_input[4571]), .B(n27822), .Z(n27464) );
  AND U27474 ( .A(n399), .B(n27823), .Z(n27822) );
  XOR U27475 ( .A(p_input[4603]), .B(p_input[4571]), .Z(n27823) );
  XNOR U27476 ( .A(n27461), .B(n27818), .Z(n27820) );
  XOR U27477 ( .A(n27824), .B(n27825), .Z(n27461) );
  AND U27478 ( .A(n397), .B(n27826), .Z(n27825) );
  XOR U27479 ( .A(p_input[4539]), .B(p_input[4507]), .Z(n27826) );
  XOR U27480 ( .A(n27827), .B(n27828), .Z(n27818) );
  AND U27481 ( .A(n27829), .B(n27830), .Z(n27828) );
  XOR U27482 ( .A(n27827), .B(n27476), .Z(n27830) );
  XNOR U27483 ( .A(p_input[4570]), .B(n27831), .Z(n27476) );
  AND U27484 ( .A(n399), .B(n27832), .Z(n27831) );
  XOR U27485 ( .A(p_input[4602]), .B(p_input[4570]), .Z(n27832) );
  XNOR U27486 ( .A(n27473), .B(n27827), .Z(n27829) );
  XOR U27487 ( .A(n27833), .B(n27834), .Z(n27473) );
  AND U27488 ( .A(n397), .B(n27835), .Z(n27834) );
  XOR U27489 ( .A(p_input[4538]), .B(p_input[4506]), .Z(n27835) );
  XOR U27490 ( .A(n27836), .B(n27837), .Z(n27827) );
  AND U27491 ( .A(n27838), .B(n27839), .Z(n27837) );
  XOR U27492 ( .A(n27836), .B(n27488), .Z(n27839) );
  XNOR U27493 ( .A(p_input[4569]), .B(n27840), .Z(n27488) );
  AND U27494 ( .A(n399), .B(n27841), .Z(n27840) );
  XOR U27495 ( .A(p_input[4601]), .B(p_input[4569]), .Z(n27841) );
  XNOR U27496 ( .A(n27485), .B(n27836), .Z(n27838) );
  XOR U27497 ( .A(n27842), .B(n27843), .Z(n27485) );
  AND U27498 ( .A(n397), .B(n27844), .Z(n27843) );
  XOR U27499 ( .A(p_input[4537]), .B(p_input[4505]), .Z(n27844) );
  XOR U27500 ( .A(n27845), .B(n27846), .Z(n27836) );
  AND U27501 ( .A(n27847), .B(n27848), .Z(n27846) );
  XOR U27502 ( .A(n27845), .B(n27500), .Z(n27848) );
  XNOR U27503 ( .A(p_input[4568]), .B(n27849), .Z(n27500) );
  AND U27504 ( .A(n399), .B(n27850), .Z(n27849) );
  XOR U27505 ( .A(p_input[4600]), .B(p_input[4568]), .Z(n27850) );
  XNOR U27506 ( .A(n27497), .B(n27845), .Z(n27847) );
  XOR U27507 ( .A(n27851), .B(n27852), .Z(n27497) );
  AND U27508 ( .A(n397), .B(n27853), .Z(n27852) );
  XOR U27509 ( .A(p_input[4536]), .B(p_input[4504]), .Z(n27853) );
  XOR U27510 ( .A(n27854), .B(n27855), .Z(n27845) );
  AND U27511 ( .A(n27856), .B(n27857), .Z(n27855) );
  XOR U27512 ( .A(n27854), .B(n27512), .Z(n27857) );
  XNOR U27513 ( .A(p_input[4567]), .B(n27858), .Z(n27512) );
  AND U27514 ( .A(n399), .B(n27859), .Z(n27858) );
  XOR U27515 ( .A(p_input[4599]), .B(p_input[4567]), .Z(n27859) );
  XNOR U27516 ( .A(n27509), .B(n27854), .Z(n27856) );
  XOR U27517 ( .A(n27860), .B(n27861), .Z(n27509) );
  AND U27518 ( .A(n397), .B(n27862), .Z(n27861) );
  XOR U27519 ( .A(p_input[4535]), .B(p_input[4503]), .Z(n27862) );
  XOR U27520 ( .A(n27863), .B(n27864), .Z(n27854) );
  AND U27521 ( .A(n27865), .B(n27866), .Z(n27864) );
  XOR U27522 ( .A(n27863), .B(n27524), .Z(n27866) );
  XNOR U27523 ( .A(p_input[4566]), .B(n27867), .Z(n27524) );
  AND U27524 ( .A(n399), .B(n27868), .Z(n27867) );
  XOR U27525 ( .A(p_input[4598]), .B(p_input[4566]), .Z(n27868) );
  XNOR U27526 ( .A(n27521), .B(n27863), .Z(n27865) );
  XOR U27527 ( .A(n27869), .B(n27870), .Z(n27521) );
  AND U27528 ( .A(n397), .B(n27871), .Z(n27870) );
  XOR U27529 ( .A(p_input[4534]), .B(p_input[4502]), .Z(n27871) );
  XOR U27530 ( .A(n27872), .B(n27873), .Z(n27863) );
  AND U27531 ( .A(n27874), .B(n27875), .Z(n27873) );
  XOR U27532 ( .A(n27872), .B(n27536), .Z(n27875) );
  XNOR U27533 ( .A(p_input[4565]), .B(n27876), .Z(n27536) );
  AND U27534 ( .A(n399), .B(n27877), .Z(n27876) );
  XOR U27535 ( .A(p_input[4597]), .B(p_input[4565]), .Z(n27877) );
  XNOR U27536 ( .A(n27533), .B(n27872), .Z(n27874) );
  XOR U27537 ( .A(n27878), .B(n27879), .Z(n27533) );
  AND U27538 ( .A(n397), .B(n27880), .Z(n27879) );
  XOR U27539 ( .A(p_input[4533]), .B(p_input[4501]), .Z(n27880) );
  XOR U27540 ( .A(n27881), .B(n27882), .Z(n27872) );
  AND U27541 ( .A(n27883), .B(n27884), .Z(n27882) );
  XOR U27542 ( .A(n27881), .B(n27548), .Z(n27884) );
  XNOR U27543 ( .A(p_input[4564]), .B(n27885), .Z(n27548) );
  AND U27544 ( .A(n399), .B(n27886), .Z(n27885) );
  XOR U27545 ( .A(p_input[4596]), .B(p_input[4564]), .Z(n27886) );
  XNOR U27546 ( .A(n27545), .B(n27881), .Z(n27883) );
  XOR U27547 ( .A(n27887), .B(n27888), .Z(n27545) );
  AND U27548 ( .A(n397), .B(n27889), .Z(n27888) );
  XOR U27549 ( .A(p_input[4532]), .B(p_input[4500]), .Z(n27889) );
  XOR U27550 ( .A(n27890), .B(n27891), .Z(n27881) );
  AND U27551 ( .A(n27892), .B(n27893), .Z(n27891) );
  XOR U27552 ( .A(n27890), .B(n27560), .Z(n27893) );
  XNOR U27553 ( .A(p_input[4563]), .B(n27894), .Z(n27560) );
  AND U27554 ( .A(n399), .B(n27895), .Z(n27894) );
  XOR U27555 ( .A(p_input[4595]), .B(p_input[4563]), .Z(n27895) );
  XNOR U27556 ( .A(n27557), .B(n27890), .Z(n27892) );
  XOR U27557 ( .A(n27896), .B(n27897), .Z(n27557) );
  AND U27558 ( .A(n397), .B(n27898), .Z(n27897) );
  XOR U27559 ( .A(p_input[4531]), .B(p_input[4499]), .Z(n27898) );
  XOR U27560 ( .A(n27899), .B(n27900), .Z(n27890) );
  AND U27561 ( .A(n27901), .B(n27902), .Z(n27900) );
  XOR U27562 ( .A(n27899), .B(n27572), .Z(n27902) );
  XNOR U27563 ( .A(p_input[4562]), .B(n27903), .Z(n27572) );
  AND U27564 ( .A(n399), .B(n27904), .Z(n27903) );
  XOR U27565 ( .A(p_input[4594]), .B(p_input[4562]), .Z(n27904) );
  XNOR U27566 ( .A(n27569), .B(n27899), .Z(n27901) );
  XOR U27567 ( .A(n27905), .B(n27906), .Z(n27569) );
  AND U27568 ( .A(n397), .B(n27907), .Z(n27906) );
  XOR U27569 ( .A(p_input[4530]), .B(p_input[4498]), .Z(n27907) );
  XOR U27570 ( .A(n27908), .B(n27909), .Z(n27899) );
  AND U27571 ( .A(n27910), .B(n27911), .Z(n27909) );
  XOR U27572 ( .A(n27908), .B(n27584), .Z(n27911) );
  XNOR U27573 ( .A(p_input[4561]), .B(n27912), .Z(n27584) );
  AND U27574 ( .A(n399), .B(n27913), .Z(n27912) );
  XOR U27575 ( .A(p_input[4593]), .B(p_input[4561]), .Z(n27913) );
  XNOR U27576 ( .A(n27581), .B(n27908), .Z(n27910) );
  XOR U27577 ( .A(n27914), .B(n27915), .Z(n27581) );
  AND U27578 ( .A(n397), .B(n27916), .Z(n27915) );
  XOR U27579 ( .A(p_input[4529]), .B(p_input[4497]), .Z(n27916) );
  XOR U27580 ( .A(n27917), .B(n27918), .Z(n27908) );
  AND U27581 ( .A(n27919), .B(n27920), .Z(n27918) );
  XOR U27582 ( .A(n27917), .B(n27596), .Z(n27920) );
  XNOR U27583 ( .A(p_input[4560]), .B(n27921), .Z(n27596) );
  AND U27584 ( .A(n399), .B(n27922), .Z(n27921) );
  XOR U27585 ( .A(p_input[4592]), .B(p_input[4560]), .Z(n27922) );
  XNOR U27586 ( .A(n27593), .B(n27917), .Z(n27919) );
  XOR U27587 ( .A(n27923), .B(n27924), .Z(n27593) );
  AND U27588 ( .A(n397), .B(n27925), .Z(n27924) );
  XOR U27589 ( .A(p_input[4528]), .B(p_input[4496]), .Z(n27925) );
  XOR U27590 ( .A(n27926), .B(n27927), .Z(n27917) );
  AND U27591 ( .A(n27928), .B(n27929), .Z(n27927) );
  XOR U27592 ( .A(n27926), .B(n27608), .Z(n27929) );
  XNOR U27593 ( .A(p_input[4559]), .B(n27930), .Z(n27608) );
  AND U27594 ( .A(n399), .B(n27931), .Z(n27930) );
  XOR U27595 ( .A(p_input[4591]), .B(p_input[4559]), .Z(n27931) );
  XNOR U27596 ( .A(n27605), .B(n27926), .Z(n27928) );
  XOR U27597 ( .A(n27932), .B(n27933), .Z(n27605) );
  AND U27598 ( .A(n397), .B(n27934), .Z(n27933) );
  XOR U27599 ( .A(p_input[4527]), .B(p_input[4495]), .Z(n27934) );
  XOR U27600 ( .A(n27935), .B(n27936), .Z(n27926) );
  AND U27601 ( .A(n27937), .B(n27938), .Z(n27936) );
  XOR U27602 ( .A(n27935), .B(n27620), .Z(n27938) );
  XNOR U27603 ( .A(p_input[4558]), .B(n27939), .Z(n27620) );
  AND U27604 ( .A(n399), .B(n27940), .Z(n27939) );
  XOR U27605 ( .A(p_input[4590]), .B(p_input[4558]), .Z(n27940) );
  XNOR U27606 ( .A(n27617), .B(n27935), .Z(n27937) );
  XOR U27607 ( .A(n27941), .B(n27942), .Z(n27617) );
  AND U27608 ( .A(n397), .B(n27943), .Z(n27942) );
  XOR U27609 ( .A(p_input[4526]), .B(p_input[4494]), .Z(n27943) );
  XOR U27610 ( .A(n27944), .B(n27945), .Z(n27935) );
  AND U27611 ( .A(n27946), .B(n27947), .Z(n27945) );
  XOR U27612 ( .A(n27944), .B(n27632), .Z(n27947) );
  XNOR U27613 ( .A(p_input[4557]), .B(n27948), .Z(n27632) );
  AND U27614 ( .A(n399), .B(n27949), .Z(n27948) );
  XOR U27615 ( .A(p_input[4589]), .B(p_input[4557]), .Z(n27949) );
  XNOR U27616 ( .A(n27629), .B(n27944), .Z(n27946) );
  XOR U27617 ( .A(n27950), .B(n27951), .Z(n27629) );
  AND U27618 ( .A(n397), .B(n27952), .Z(n27951) );
  XOR U27619 ( .A(p_input[4525]), .B(p_input[4493]), .Z(n27952) );
  XOR U27620 ( .A(n27953), .B(n27954), .Z(n27944) );
  AND U27621 ( .A(n27955), .B(n27956), .Z(n27954) );
  XOR U27622 ( .A(n27953), .B(n27644), .Z(n27956) );
  XNOR U27623 ( .A(p_input[4556]), .B(n27957), .Z(n27644) );
  AND U27624 ( .A(n399), .B(n27958), .Z(n27957) );
  XOR U27625 ( .A(p_input[4588]), .B(p_input[4556]), .Z(n27958) );
  XNOR U27626 ( .A(n27641), .B(n27953), .Z(n27955) );
  XOR U27627 ( .A(n27959), .B(n27960), .Z(n27641) );
  AND U27628 ( .A(n397), .B(n27961), .Z(n27960) );
  XOR U27629 ( .A(p_input[4524]), .B(p_input[4492]), .Z(n27961) );
  XOR U27630 ( .A(n27962), .B(n27963), .Z(n27953) );
  AND U27631 ( .A(n27964), .B(n27965), .Z(n27963) );
  XOR U27632 ( .A(n27962), .B(n27656), .Z(n27965) );
  XNOR U27633 ( .A(p_input[4555]), .B(n27966), .Z(n27656) );
  AND U27634 ( .A(n399), .B(n27967), .Z(n27966) );
  XOR U27635 ( .A(p_input[4587]), .B(p_input[4555]), .Z(n27967) );
  XNOR U27636 ( .A(n27653), .B(n27962), .Z(n27964) );
  XOR U27637 ( .A(n27968), .B(n27969), .Z(n27653) );
  AND U27638 ( .A(n397), .B(n27970), .Z(n27969) );
  XOR U27639 ( .A(p_input[4523]), .B(p_input[4491]), .Z(n27970) );
  XOR U27640 ( .A(n27971), .B(n27972), .Z(n27962) );
  AND U27641 ( .A(n27973), .B(n27974), .Z(n27972) );
  XOR U27642 ( .A(n27971), .B(n27668), .Z(n27974) );
  XNOR U27643 ( .A(p_input[4554]), .B(n27975), .Z(n27668) );
  AND U27644 ( .A(n399), .B(n27976), .Z(n27975) );
  XOR U27645 ( .A(p_input[4586]), .B(p_input[4554]), .Z(n27976) );
  XNOR U27646 ( .A(n27665), .B(n27971), .Z(n27973) );
  XOR U27647 ( .A(n27977), .B(n27978), .Z(n27665) );
  AND U27648 ( .A(n397), .B(n27979), .Z(n27978) );
  XOR U27649 ( .A(p_input[4522]), .B(p_input[4490]), .Z(n27979) );
  XOR U27650 ( .A(n27980), .B(n27981), .Z(n27971) );
  AND U27651 ( .A(n27982), .B(n27983), .Z(n27981) );
  XOR U27652 ( .A(n27980), .B(n27680), .Z(n27983) );
  XNOR U27653 ( .A(p_input[4553]), .B(n27984), .Z(n27680) );
  AND U27654 ( .A(n399), .B(n27985), .Z(n27984) );
  XOR U27655 ( .A(p_input[4585]), .B(p_input[4553]), .Z(n27985) );
  XNOR U27656 ( .A(n27677), .B(n27980), .Z(n27982) );
  XOR U27657 ( .A(n27986), .B(n27987), .Z(n27677) );
  AND U27658 ( .A(n397), .B(n27988), .Z(n27987) );
  XOR U27659 ( .A(p_input[4521]), .B(p_input[4489]), .Z(n27988) );
  XOR U27660 ( .A(n27989), .B(n27990), .Z(n27980) );
  AND U27661 ( .A(n27991), .B(n27992), .Z(n27990) );
  XOR U27662 ( .A(n27989), .B(n27692), .Z(n27992) );
  XNOR U27663 ( .A(p_input[4552]), .B(n27993), .Z(n27692) );
  AND U27664 ( .A(n399), .B(n27994), .Z(n27993) );
  XOR U27665 ( .A(p_input[4584]), .B(p_input[4552]), .Z(n27994) );
  XNOR U27666 ( .A(n27689), .B(n27989), .Z(n27991) );
  XOR U27667 ( .A(n27995), .B(n27996), .Z(n27689) );
  AND U27668 ( .A(n397), .B(n27997), .Z(n27996) );
  XOR U27669 ( .A(p_input[4520]), .B(p_input[4488]), .Z(n27997) );
  XOR U27670 ( .A(n27998), .B(n27999), .Z(n27989) );
  AND U27671 ( .A(n28000), .B(n28001), .Z(n27999) );
  XOR U27672 ( .A(n27998), .B(n27704), .Z(n28001) );
  XNOR U27673 ( .A(p_input[4551]), .B(n28002), .Z(n27704) );
  AND U27674 ( .A(n399), .B(n28003), .Z(n28002) );
  XOR U27675 ( .A(p_input[4583]), .B(p_input[4551]), .Z(n28003) );
  XNOR U27676 ( .A(n27701), .B(n27998), .Z(n28000) );
  XOR U27677 ( .A(n28004), .B(n28005), .Z(n27701) );
  AND U27678 ( .A(n397), .B(n28006), .Z(n28005) );
  XOR U27679 ( .A(p_input[4519]), .B(p_input[4487]), .Z(n28006) );
  XOR U27680 ( .A(n28007), .B(n28008), .Z(n27998) );
  AND U27681 ( .A(n28009), .B(n28010), .Z(n28008) );
  XOR U27682 ( .A(n28007), .B(n27716), .Z(n28010) );
  XNOR U27683 ( .A(p_input[4550]), .B(n28011), .Z(n27716) );
  AND U27684 ( .A(n399), .B(n28012), .Z(n28011) );
  XOR U27685 ( .A(p_input[4582]), .B(p_input[4550]), .Z(n28012) );
  XNOR U27686 ( .A(n27713), .B(n28007), .Z(n28009) );
  XOR U27687 ( .A(n28013), .B(n28014), .Z(n27713) );
  AND U27688 ( .A(n397), .B(n28015), .Z(n28014) );
  XOR U27689 ( .A(p_input[4518]), .B(p_input[4486]), .Z(n28015) );
  XOR U27690 ( .A(n28016), .B(n28017), .Z(n28007) );
  AND U27691 ( .A(n28018), .B(n28019), .Z(n28017) );
  XOR U27692 ( .A(n28016), .B(n27728), .Z(n28019) );
  XNOR U27693 ( .A(p_input[4549]), .B(n28020), .Z(n27728) );
  AND U27694 ( .A(n399), .B(n28021), .Z(n28020) );
  XOR U27695 ( .A(p_input[4581]), .B(p_input[4549]), .Z(n28021) );
  XNOR U27696 ( .A(n27725), .B(n28016), .Z(n28018) );
  XOR U27697 ( .A(n28022), .B(n28023), .Z(n27725) );
  AND U27698 ( .A(n397), .B(n28024), .Z(n28023) );
  XOR U27699 ( .A(p_input[4517]), .B(p_input[4485]), .Z(n28024) );
  XOR U27700 ( .A(n28025), .B(n28026), .Z(n28016) );
  AND U27701 ( .A(n28027), .B(n28028), .Z(n28026) );
  XOR U27702 ( .A(n28025), .B(n27740), .Z(n28028) );
  XNOR U27703 ( .A(p_input[4548]), .B(n28029), .Z(n27740) );
  AND U27704 ( .A(n399), .B(n28030), .Z(n28029) );
  XOR U27705 ( .A(p_input[4580]), .B(p_input[4548]), .Z(n28030) );
  XNOR U27706 ( .A(n27737), .B(n28025), .Z(n28027) );
  XOR U27707 ( .A(n28031), .B(n28032), .Z(n27737) );
  AND U27708 ( .A(n397), .B(n28033), .Z(n28032) );
  XOR U27709 ( .A(p_input[4516]), .B(p_input[4484]), .Z(n28033) );
  XOR U27710 ( .A(n28034), .B(n28035), .Z(n28025) );
  AND U27711 ( .A(n28036), .B(n28037), .Z(n28035) );
  XOR U27712 ( .A(n28034), .B(n27752), .Z(n28037) );
  XNOR U27713 ( .A(p_input[4547]), .B(n28038), .Z(n27752) );
  AND U27714 ( .A(n399), .B(n28039), .Z(n28038) );
  XOR U27715 ( .A(p_input[4579]), .B(p_input[4547]), .Z(n28039) );
  XNOR U27716 ( .A(n27749), .B(n28034), .Z(n28036) );
  XOR U27717 ( .A(n28040), .B(n28041), .Z(n27749) );
  AND U27718 ( .A(n397), .B(n28042), .Z(n28041) );
  XOR U27719 ( .A(p_input[4515]), .B(p_input[4483]), .Z(n28042) );
  XOR U27720 ( .A(n28043), .B(n28044), .Z(n28034) );
  AND U27721 ( .A(n28045), .B(n28046), .Z(n28044) );
  XOR U27722 ( .A(n28043), .B(n27764), .Z(n28046) );
  XNOR U27723 ( .A(p_input[4546]), .B(n28047), .Z(n27764) );
  AND U27724 ( .A(n399), .B(n28048), .Z(n28047) );
  XOR U27725 ( .A(p_input[4578]), .B(p_input[4546]), .Z(n28048) );
  XNOR U27726 ( .A(n27761), .B(n28043), .Z(n28045) );
  XOR U27727 ( .A(n28049), .B(n28050), .Z(n27761) );
  AND U27728 ( .A(n397), .B(n28051), .Z(n28050) );
  XOR U27729 ( .A(p_input[4514]), .B(p_input[4482]), .Z(n28051) );
  XOR U27730 ( .A(n28052), .B(n28053), .Z(n28043) );
  AND U27731 ( .A(n28054), .B(n28055), .Z(n28053) );
  XNOR U27732 ( .A(n28056), .B(n27777), .Z(n28055) );
  XNOR U27733 ( .A(p_input[4545]), .B(n28057), .Z(n27777) );
  AND U27734 ( .A(n399), .B(n28058), .Z(n28057) );
  XNOR U27735 ( .A(p_input[4577]), .B(n28059), .Z(n28058) );
  IV U27736 ( .A(p_input[4545]), .Z(n28059) );
  XNOR U27737 ( .A(n27774), .B(n28052), .Z(n28054) );
  XNOR U27738 ( .A(p_input[4481]), .B(n28060), .Z(n27774) );
  AND U27739 ( .A(n397), .B(n28061), .Z(n28060) );
  XOR U27740 ( .A(p_input[4513]), .B(p_input[4481]), .Z(n28061) );
  IV U27741 ( .A(n28056), .Z(n28052) );
  AND U27742 ( .A(n27782), .B(n27785), .Z(n28056) );
  XOR U27743 ( .A(p_input[4544]), .B(n28062), .Z(n27785) );
  AND U27744 ( .A(n399), .B(n28063), .Z(n28062) );
  XOR U27745 ( .A(p_input[4576]), .B(p_input[4544]), .Z(n28063) );
  XOR U27746 ( .A(n28064), .B(n28065), .Z(n399) );
  AND U27747 ( .A(n28066), .B(n28067), .Z(n28065) );
  XNOR U27748 ( .A(p_input[4607]), .B(n28064), .Z(n28067) );
  XOR U27749 ( .A(n28064), .B(p_input[4575]), .Z(n28066) );
  XOR U27750 ( .A(n28068), .B(n28069), .Z(n28064) );
  AND U27751 ( .A(n28070), .B(n28071), .Z(n28069) );
  XNOR U27752 ( .A(p_input[4606]), .B(n28068), .Z(n28071) );
  XOR U27753 ( .A(n28068), .B(p_input[4574]), .Z(n28070) );
  XOR U27754 ( .A(n28072), .B(n28073), .Z(n28068) );
  AND U27755 ( .A(n28074), .B(n28075), .Z(n28073) );
  XNOR U27756 ( .A(p_input[4605]), .B(n28072), .Z(n28075) );
  XOR U27757 ( .A(n28072), .B(p_input[4573]), .Z(n28074) );
  XOR U27758 ( .A(n28076), .B(n28077), .Z(n28072) );
  AND U27759 ( .A(n28078), .B(n28079), .Z(n28077) );
  XNOR U27760 ( .A(p_input[4604]), .B(n28076), .Z(n28079) );
  XOR U27761 ( .A(n28076), .B(p_input[4572]), .Z(n28078) );
  XOR U27762 ( .A(n28080), .B(n28081), .Z(n28076) );
  AND U27763 ( .A(n28082), .B(n28083), .Z(n28081) );
  XNOR U27764 ( .A(p_input[4603]), .B(n28080), .Z(n28083) );
  XOR U27765 ( .A(n28080), .B(p_input[4571]), .Z(n28082) );
  XOR U27766 ( .A(n28084), .B(n28085), .Z(n28080) );
  AND U27767 ( .A(n28086), .B(n28087), .Z(n28085) );
  XNOR U27768 ( .A(p_input[4602]), .B(n28084), .Z(n28087) );
  XOR U27769 ( .A(n28084), .B(p_input[4570]), .Z(n28086) );
  XOR U27770 ( .A(n28088), .B(n28089), .Z(n28084) );
  AND U27771 ( .A(n28090), .B(n28091), .Z(n28089) );
  XNOR U27772 ( .A(p_input[4601]), .B(n28088), .Z(n28091) );
  XOR U27773 ( .A(n28088), .B(p_input[4569]), .Z(n28090) );
  XOR U27774 ( .A(n28092), .B(n28093), .Z(n28088) );
  AND U27775 ( .A(n28094), .B(n28095), .Z(n28093) );
  XNOR U27776 ( .A(p_input[4600]), .B(n28092), .Z(n28095) );
  XOR U27777 ( .A(n28092), .B(p_input[4568]), .Z(n28094) );
  XOR U27778 ( .A(n28096), .B(n28097), .Z(n28092) );
  AND U27779 ( .A(n28098), .B(n28099), .Z(n28097) );
  XNOR U27780 ( .A(p_input[4599]), .B(n28096), .Z(n28099) );
  XOR U27781 ( .A(n28096), .B(p_input[4567]), .Z(n28098) );
  XOR U27782 ( .A(n28100), .B(n28101), .Z(n28096) );
  AND U27783 ( .A(n28102), .B(n28103), .Z(n28101) );
  XNOR U27784 ( .A(p_input[4598]), .B(n28100), .Z(n28103) );
  XOR U27785 ( .A(n28100), .B(p_input[4566]), .Z(n28102) );
  XOR U27786 ( .A(n28104), .B(n28105), .Z(n28100) );
  AND U27787 ( .A(n28106), .B(n28107), .Z(n28105) );
  XNOR U27788 ( .A(p_input[4597]), .B(n28104), .Z(n28107) );
  XOR U27789 ( .A(n28104), .B(p_input[4565]), .Z(n28106) );
  XOR U27790 ( .A(n28108), .B(n28109), .Z(n28104) );
  AND U27791 ( .A(n28110), .B(n28111), .Z(n28109) );
  XNOR U27792 ( .A(p_input[4596]), .B(n28108), .Z(n28111) );
  XOR U27793 ( .A(n28108), .B(p_input[4564]), .Z(n28110) );
  XOR U27794 ( .A(n28112), .B(n28113), .Z(n28108) );
  AND U27795 ( .A(n28114), .B(n28115), .Z(n28113) );
  XNOR U27796 ( .A(p_input[4595]), .B(n28112), .Z(n28115) );
  XOR U27797 ( .A(n28112), .B(p_input[4563]), .Z(n28114) );
  XOR U27798 ( .A(n28116), .B(n28117), .Z(n28112) );
  AND U27799 ( .A(n28118), .B(n28119), .Z(n28117) );
  XNOR U27800 ( .A(p_input[4594]), .B(n28116), .Z(n28119) );
  XOR U27801 ( .A(n28116), .B(p_input[4562]), .Z(n28118) );
  XOR U27802 ( .A(n28120), .B(n28121), .Z(n28116) );
  AND U27803 ( .A(n28122), .B(n28123), .Z(n28121) );
  XNOR U27804 ( .A(p_input[4593]), .B(n28120), .Z(n28123) );
  XOR U27805 ( .A(n28120), .B(p_input[4561]), .Z(n28122) );
  XOR U27806 ( .A(n28124), .B(n28125), .Z(n28120) );
  AND U27807 ( .A(n28126), .B(n28127), .Z(n28125) );
  XNOR U27808 ( .A(p_input[4592]), .B(n28124), .Z(n28127) );
  XOR U27809 ( .A(n28124), .B(p_input[4560]), .Z(n28126) );
  XOR U27810 ( .A(n28128), .B(n28129), .Z(n28124) );
  AND U27811 ( .A(n28130), .B(n28131), .Z(n28129) );
  XNOR U27812 ( .A(p_input[4591]), .B(n28128), .Z(n28131) );
  XOR U27813 ( .A(n28128), .B(p_input[4559]), .Z(n28130) );
  XOR U27814 ( .A(n28132), .B(n28133), .Z(n28128) );
  AND U27815 ( .A(n28134), .B(n28135), .Z(n28133) );
  XNOR U27816 ( .A(p_input[4590]), .B(n28132), .Z(n28135) );
  XOR U27817 ( .A(n28132), .B(p_input[4558]), .Z(n28134) );
  XOR U27818 ( .A(n28136), .B(n28137), .Z(n28132) );
  AND U27819 ( .A(n28138), .B(n28139), .Z(n28137) );
  XNOR U27820 ( .A(p_input[4589]), .B(n28136), .Z(n28139) );
  XOR U27821 ( .A(n28136), .B(p_input[4557]), .Z(n28138) );
  XOR U27822 ( .A(n28140), .B(n28141), .Z(n28136) );
  AND U27823 ( .A(n28142), .B(n28143), .Z(n28141) );
  XNOR U27824 ( .A(p_input[4588]), .B(n28140), .Z(n28143) );
  XOR U27825 ( .A(n28140), .B(p_input[4556]), .Z(n28142) );
  XOR U27826 ( .A(n28144), .B(n28145), .Z(n28140) );
  AND U27827 ( .A(n28146), .B(n28147), .Z(n28145) );
  XNOR U27828 ( .A(p_input[4587]), .B(n28144), .Z(n28147) );
  XOR U27829 ( .A(n28144), .B(p_input[4555]), .Z(n28146) );
  XOR U27830 ( .A(n28148), .B(n28149), .Z(n28144) );
  AND U27831 ( .A(n28150), .B(n28151), .Z(n28149) );
  XNOR U27832 ( .A(p_input[4586]), .B(n28148), .Z(n28151) );
  XOR U27833 ( .A(n28148), .B(p_input[4554]), .Z(n28150) );
  XOR U27834 ( .A(n28152), .B(n28153), .Z(n28148) );
  AND U27835 ( .A(n28154), .B(n28155), .Z(n28153) );
  XNOR U27836 ( .A(p_input[4585]), .B(n28152), .Z(n28155) );
  XOR U27837 ( .A(n28152), .B(p_input[4553]), .Z(n28154) );
  XOR U27838 ( .A(n28156), .B(n28157), .Z(n28152) );
  AND U27839 ( .A(n28158), .B(n28159), .Z(n28157) );
  XNOR U27840 ( .A(p_input[4584]), .B(n28156), .Z(n28159) );
  XOR U27841 ( .A(n28156), .B(p_input[4552]), .Z(n28158) );
  XOR U27842 ( .A(n28160), .B(n28161), .Z(n28156) );
  AND U27843 ( .A(n28162), .B(n28163), .Z(n28161) );
  XNOR U27844 ( .A(p_input[4583]), .B(n28160), .Z(n28163) );
  XOR U27845 ( .A(n28160), .B(p_input[4551]), .Z(n28162) );
  XOR U27846 ( .A(n28164), .B(n28165), .Z(n28160) );
  AND U27847 ( .A(n28166), .B(n28167), .Z(n28165) );
  XNOR U27848 ( .A(p_input[4582]), .B(n28164), .Z(n28167) );
  XOR U27849 ( .A(n28164), .B(p_input[4550]), .Z(n28166) );
  XOR U27850 ( .A(n28168), .B(n28169), .Z(n28164) );
  AND U27851 ( .A(n28170), .B(n28171), .Z(n28169) );
  XNOR U27852 ( .A(p_input[4581]), .B(n28168), .Z(n28171) );
  XOR U27853 ( .A(n28168), .B(p_input[4549]), .Z(n28170) );
  XOR U27854 ( .A(n28172), .B(n28173), .Z(n28168) );
  AND U27855 ( .A(n28174), .B(n28175), .Z(n28173) );
  XNOR U27856 ( .A(p_input[4580]), .B(n28172), .Z(n28175) );
  XOR U27857 ( .A(n28172), .B(p_input[4548]), .Z(n28174) );
  XOR U27858 ( .A(n28176), .B(n28177), .Z(n28172) );
  AND U27859 ( .A(n28178), .B(n28179), .Z(n28177) );
  XNOR U27860 ( .A(p_input[4579]), .B(n28176), .Z(n28179) );
  XOR U27861 ( .A(n28176), .B(p_input[4547]), .Z(n28178) );
  XOR U27862 ( .A(n28180), .B(n28181), .Z(n28176) );
  AND U27863 ( .A(n28182), .B(n28183), .Z(n28181) );
  XNOR U27864 ( .A(p_input[4578]), .B(n28180), .Z(n28183) );
  XOR U27865 ( .A(n28180), .B(p_input[4546]), .Z(n28182) );
  XNOR U27866 ( .A(n28184), .B(n28185), .Z(n28180) );
  AND U27867 ( .A(n28186), .B(n28187), .Z(n28185) );
  XOR U27868 ( .A(p_input[4577]), .B(n28184), .Z(n28187) );
  XNOR U27869 ( .A(p_input[4545]), .B(n28184), .Z(n28186) );
  AND U27870 ( .A(p_input[4576]), .B(n28188), .Z(n28184) );
  IV U27871 ( .A(p_input[4544]), .Z(n28188) );
  XNOR U27872 ( .A(p_input[4480]), .B(n28189), .Z(n27782) );
  AND U27873 ( .A(n397), .B(n28190), .Z(n28189) );
  XOR U27874 ( .A(p_input[4512]), .B(p_input[4480]), .Z(n28190) );
  XOR U27875 ( .A(n28191), .B(n28192), .Z(n397) );
  AND U27876 ( .A(n28193), .B(n28194), .Z(n28192) );
  XNOR U27877 ( .A(p_input[4543]), .B(n28191), .Z(n28194) );
  XOR U27878 ( .A(n28191), .B(p_input[4511]), .Z(n28193) );
  XOR U27879 ( .A(n28195), .B(n28196), .Z(n28191) );
  AND U27880 ( .A(n28197), .B(n28198), .Z(n28196) );
  XNOR U27881 ( .A(p_input[4542]), .B(n28195), .Z(n28198) );
  XNOR U27882 ( .A(n28195), .B(n27797), .Z(n28197) );
  IV U27883 ( .A(p_input[4510]), .Z(n27797) );
  XOR U27884 ( .A(n28199), .B(n28200), .Z(n28195) );
  AND U27885 ( .A(n28201), .B(n28202), .Z(n28200) );
  XNOR U27886 ( .A(p_input[4541]), .B(n28199), .Z(n28202) );
  XNOR U27887 ( .A(n28199), .B(n27806), .Z(n28201) );
  IV U27888 ( .A(p_input[4509]), .Z(n27806) );
  XOR U27889 ( .A(n28203), .B(n28204), .Z(n28199) );
  AND U27890 ( .A(n28205), .B(n28206), .Z(n28204) );
  XNOR U27891 ( .A(p_input[4540]), .B(n28203), .Z(n28206) );
  XNOR U27892 ( .A(n28203), .B(n27815), .Z(n28205) );
  IV U27893 ( .A(p_input[4508]), .Z(n27815) );
  XOR U27894 ( .A(n28207), .B(n28208), .Z(n28203) );
  AND U27895 ( .A(n28209), .B(n28210), .Z(n28208) );
  XNOR U27896 ( .A(p_input[4539]), .B(n28207), .Z(n28210) );
  XNOR U27897 ( .A(n28207), .B(n27824), .Z(n28209) );
  IV U27898 ( .A(p_input[4507]), .Z(n27824) );
  XOR U27899 ( .A(n28211), .B(n28212), .Z(n28207) );
  AND U27900 ( .A(n28213), .B(n28214), .Z(n28212) );
  XNOR U27901 ( .A(p_input[4538]), .B(n28211), .Z(n28214) );
  XNOR U27902 ( .A(n28211), .B(n27833), .Z(n28213) );
  IV U27903 ( .A(p_input[4506]), .Z(n27833) );
  XOR U27904 ( .A(n28215), .B(n28216), .Z(n28211) );
  AND U27905 ( .A(n28217), .B(n28218), .Z(n28216) );
  XNOR U27906 ( .A(p_input[4537]), .B(n28215), .Z(n28218) );
  XNOR U27907 ( .A(n28215), .B(n27842), .Z(n28217) );
  IV U27908 ( .A(p_input[4505]), .Z(n27842) );
  XOR U27909 ( .A(n28219), .B(n28220), .Z(n28215) );
  AND U27910 ( .A(n28221), .B(n28222), .Z(n28220) );
  XNOR U27911 ( .A(p_input[4536]), .B(n28219), .Z(n28222) );
  XNOR U27912 ( .A(n28219), .B(n27851), .Z(n28221) );
  IV U27913 ( .A(p_input[4504]), .Z(n27851) );
  XOR U27914 ( .A(n28223), .B(n28224), .Z(n28219) );
  AND U27915 ( .A(n28225), .B(n28226), .Z(n28224) );
  XNOR U27916 ( .A(p_input[4535]), .B(n28223), .Z(n28226) );
  XNOR U27917 ( .A(n28223), .B(n27860), .Z(n28225) );
  IV U27918 ( .A(p_input[4503]), .Z(n27860) );
  XOR U27919 ( .A(n28227), .B(n28228), .Z(n28223) );
  AND U27920 ( .A(n28229), .B(n28230), .Z(n28228) );
  XNOR U27921 ( .A(p_input[4534]), .B(n28227), .Z(n28230) );
  XNOR U27922 ( .A(n28227), .B(n27869), .Z(n28229) );
  IV U27923 ( .A(p_input[4502]), .Z(n27869) );
  XOR U27924 ( .A(n28231), .B(n28232), .Z(n28227) );
  AND U27925 ( .A(n28233), .B(n28234), .Z(n28232) );
  XNOR U27926 ( .A(p_input[4533]), .B(n28231), .Z(n28234) );
  XNOR U27927 ( .A(n28231), .B(n27878), .Z(n28233) );
  IV U27928 ( .A(p_input[4501]), .Z(n27878) );
  XOR U27929 ( .A(n28235), .B(n28236), .Z(n28231) );
  AND U27930 ( .A(n28237), .B(n28238), .Z(n28236) );
  XNOR U27931 ( .A(p_input[4532]), .B(n28235), .Z(n28238) );
  XNOR U27932 ( .A(n28235), .B(n27887), .Z(n28237) );
  IV U27933 ( .A(p_input[4500]), .Z(n27887) );
  XOR U27934 ( .A(n28239), .B(n28240), .Z(n28235) );
  AND U27935 ( .A(n28241), .B(n28242), .Z(n28240) );
  XNOR U27936 ( .A(p_input[4531]), .B(n28239), .Z(n28242) );
  XNOR U27937 ( .A(n28239), .B(n27896), .Z(n28241) );
  IV U27938 ( .A(p_input[4499]), .Z(n27896) );
  XOR U27939 ( .A(n28243), .B(n28244), .Z(n28239) );
  AND U27940 ( .A(n28245), .B(n28246), .Z(n28244) );
  XNOR U27941 ( .A(p_input[4530]), .B(n28243), .Z(n28246) );
  XNOR U27942 ( .A(n28243), .B(n27905), .Z(n28245) );
  IV U27943 ( .A(p_input[4498]), .Z(n27905) );
  XOR U27944 ( .A(n28247), .B(n28248), .Z(n28243) );
  AND U27945 ( .A(n28249), .B(n28250), .Z(n28248) );
  XNOR U27946 ( .A(p_input[4529]), .B(n28247), .Z(n28250) );
  XNOR U27947 ( .A(n28247), .B(n27914), .Z(n28249) );
  IV U27948 ( .A(p_input[4497]), .Z(n27914) );
  XOR U27949 ( .A(n28251), .B(n28252), .Z(n28247) );
  AND U27950 ( .A(n28253), .B(n28254), .Z(n28252) );
  XNOR U27951 ( .A(p_input[4528]), .B(n28251), .Z(n28254) );
  XNOR U27952 ( .A(n28251), .B(n27923), .Z(n28253) );
  IV U27953 ( .A(p_input[4496]), .Z(n27923) );
  XOR U27954 ( .A(n28255), .B(n28256), .Z(n28251) );
  AND U27955 ( .A(n28257), .B(n28258), .Z(n28256) );
  XNOR U27956 ( .A(p_input[4527]), .B(n28255), .Z(n28258) );
  XNOR U27957 ( .A(n28255), .B(n27932), .Z(n28257) );
  IV U27958 ( .A(p_input[4495]), .Z(n27932) );
  XOR U27959 ( .A(n28259), .B(n28260), .Z(n28255) );
  AND U27960 ( .A(n28261), .B(n28262), .Z(n28260) );
  XNOR U27961 ( .A(p_input[4526]), .B(n28259), .Z(n28262) );
  XNOR U27962 ( .A(n28259), .B(n27941), .Z(n28261) );
  IV U27963 ( .A(p_input[4494]), .Z(n27941) );
  XOR U27964 ( .A(n28263), .B(n28264), .Z(n28259) );
  AND U27965 ( .A(n28265), .B(n28266), .Z(n28264) );
  XNOR U27966 ( .A(p_input[4525]), .B(n28263), .Z(n28266) );
  XNOR U27967 ( .A(n28263), .B(n27950), .Z(n28265) );
  IV U27968 ( .A(p_input[4493]), .Z(n27950) );
  XOR U27969 ( .A(n28267), .B(n28268), .Z(n28263) );
  AND U27970 ( .A(n28269), .B(n28270), .Z(n28268) );
  XNOR U27971 ( .A(p_input[4524]), .B(n28267), .Z(n28270) );
  XNOR U27972 ( .A(n28267), .B(n27959), .Z(n28269) );
  IV U27973 ( .A(p_input[4492]), .Z(n27959) );
  XOR U27974 ( .A(n28271), .B(n28272), .Z(n28267) );
  AND U27975 ( .A(n28273), .B(n28274), .Z(n28272) );
  XNOR U27976 ( .A(p_input[4523]), .B(n28271), .Z(n28274) );
  XNOR U27977 ( .A(n28271), .B(n27968), .Z(n28273) );
  IV U27978 ( .A(p_input[4491]), .Z(n27968) );
  XOR U27979 ( .A(n28275), .B(n28276), .Z(n28271) );
  AND U27980 ( .A(n28277), .B(n28278), .Z(n28276) );
  XNOR U27981 ( .A(p_input[4522]), .B(n28275), .Z(n28278) );
  XNOR U27982 ( .A(n28275), .B(n27977), .Z(n28277) );
  IV U27983 ( .A(p_input[4490]), .Z(n27977) );
  XOR U27984 ( .A(n28279), .B(n28280), .Z(n28275) );
  AND U27985 ( .A(n28281), .B(n28282), .Z(n28280) );
  XNOR U27986 ( .A(p_input[4521]), .B(n28279), .Z(n28282) );
  XNOR U27987 ( .A(n28279), .B(n27986), .Z(n28281) );
  IV U27988 ( .A(p_input[4489]), .Z(n27986) );
  XOR U27989 ( .A(n28283), .B(n28284), .Z(n28279) );
  AND U27990 ( .A(n28285), .B(n28286), .Z(n28284) );
  XNOR U27991 ( .A(p_input[4520]), .B(n28283), .Z(n28286) );
  XNOR U27992 ( .A(n28283), .B(n27995), .Z(n28285) );
  IV U27993 ( .A(p_input[4488]), .Z(n27995) );
  XOR U27994 ( .A(n28287), .B(n28288), .Z(n28283) );
  AND U27995 ( .A(n28289), .B(n28290), .Z(n28288) );
  XNOR U27996 ( .A(p_input[4519]), .B(n28287), .Z(n28290) );
  XNOR U27997 ( .A(n28287), .B(n28004), .Z(n28289) );
  IV U27998 ( .A(p_input[4487]), .Z(n28004) );
  XOR U27999 ( .A(n28291), .B(n28292), .Z(n28287) );
  AND U28000 ( .A(n28293), .B(n28294), .Z(n28292) );
  XNOR U28001 ( .A(p_input[4518]), .B(n28291), .Z(n28294) );
  XNOR U28002 ( .A(n28291), .B(n28013), .Z(n28293) );
  IV U28003 ( .A(p_input[4486]), .Z(n28013) );
  XOR U28004 ( .A(n28295), .B(n28296), .Z(n28291) );
  AND U28005 ( .A(n28297), .B(n28298), .Z(n28296) );
  XNOR U28006 ( .A(p_input[4517]), .B(n28295), .Z(n28298) );
  XNOR U28007 ( .A(n28295), .B(n28022), .Z(n28297) );
  IV U28008 ( .A(p_input[4485]), .Z(n28022) );
  XOR U28009 ( .A(n28299), .B(n28300), .Z(n28295) );
  AND U28010 ( .A(n28301), .B(n28302), .Z(n28300) );
  XNOR U28011 ( .A(p_input[4516]), .B(n28299), .Z(n28302) );
  XNOR U28012 ( .A(n28299), .B(n28031), .Z(n28301) );
  IV U28013 ( .A(p_input[4484]), .Z(n28031) );
  XOR U28014 ( .A(n28303), .B(n28304), .Z(n28299) );
  AND U28015 ( .A(n28305), .B(n28306), .Z(n28304) );
  XNOR U28016 ( .A(p_input[4515]), .B(n28303), .Z(n28306) );
  XNOR U28017 ( .A(n28303), .B(n28040), .Z(n28305) );
  IV U28018 ( .A(p_input[4483]), .Z(n28040) );
  XOR U28019 ( .A(n28307), .B(n28308), .Z(n28303) );
  AND U28020 ( .A(n28309), .B(n28310), .Z(n28308) );
  XNOR U28021 ( .A(p_input[4514]), .B(n28307), .Z(n28310) );
  XNOR U28022 ( .A(n28307), .B(n28049), .Z(n28309) );
  IV U28023 ( .A(p_input[4482]), .Z(n28049) );
  XNOR U28024 ( .A(n28311), .B(n28312), .Z(n28307) );
  AND U28025 ( .A(n28313), .B(n28314), .Z(n28312) );
  XOR U28026 ( .A(p_input[4513]), .B(n28311), .Z(n28314) );
  XNOR U28027 ( .A(p_input[4481]), .B(n28311), .Z(n28313) );
  AND U28028 ( .A(p_input[4512]), .B(n28315), .Z(n28311) );
  IV U28029 ( .A(p_input[4480]), .Z(n28315) );
  XOR U28030 ( .A(n28316), .B(n28317), .Z(n27405) );
  AND U28031 ( .A(n537), .B(n28318), .Z(n28317) );
  XNOR U28032 ( .A(n28319), .B(n28316), .Z(n28318) );
  XOR U28033 ( .A(n28320), .B(n28321), .Z(n537) );
  AND U28034 ( .A(n28322), .B(n28323), .Z(n28321) );
  XNOR U28035 ( .A(n27420), .B(n28320), .Z(n28323) );
  AND U28036 ( .A(p_input[4479]), .B(p_input[4447]), .Z(n27420) );
  XNOR U28037 ( .A(n28320), .B(n27417), .Z(n28322) );
  IV U28038 ( .A(n28324), .Z(n27417) );
  AND U28039 ( .A(p_input[4383]), .B(p_input[4415]), .Z(n28324) );
  XOR U28040 ( .A(n28325), .B(n28326), .Z(n28320) );
  AND U28041 ( .A(n28327), .B(n28328), .Z(n28326) );
  XOR U28042 ( .A(n28325), .B(n27432), .Z(n28328) );
  XNOR U28043 ( .A(p_input[4446]), .B(n28329), .Z(n27432) );
  AND U28044 ( .A(n403), .B(n28330), .Z(n28329) );
  XOR U28045 ( .A(p_input[4478]), .B(p_input[4446]), .Z(n28330) );
  XNOR U28046 ( .A(n27429), .B(n28325), .Z(n28327) );
  XOR U28047 ( .A(n28331), .B(n28332), .Z(n27429) );
  AND U28048 ( .A(n400), .B(n28333), .Z(n28332) );
  XOR U28049 ( .A(p_input[4414]), .B(p_input[4382]), .Z(n28333) );
  XOR U28050 ( .A(n28334), .B(n28335), .Z(n28325) );
  AND U28051 ( .A(n28336), .B(n28337), .Z(n28335) );
  XOR U28052 ( .A(n28334), .B(n27444), .Z(n28337) );
  XNOR U28053 ( .A(p_input[4445]), .B(n28338), .Z(n27444) );
  AND U28054 ( .A(n403), .B(n28339), .Z(n28338) );
  XOR U28055 ( .A(p_input[4477]), .B(p_input[4445]), .Z(n28339) );
  XNOR U28056 ( .A(n27441), .B(n28334), .Z(n28336) );
  XOR U28057 ( .A(n28340), .B(n28341), .Z(n27441) );
  AND U28058 ( .A(n400), .B(n28342), .Z(n28341) );
  XOR U28059 ( .A(p_input[4413]), .B(p_input[4381]), .Z(n28342) );
  XOR U28060 ( .A(n28343), .B(n28344), .Z(n28334) );
  AND U28061 ( .A(n28345), .B(n28346), .Z(n28344) );
  XOR U28062 ( .A(n28343), .B(n27456), .Z(n28346) );
  XNOR U28063 ( .A(p_input[4444]), .B(n28347), .Z(n27456) );
  AND U28064 ( .A(n403), .B(n28348), .Z(n28347) );
  XOR U28065 ( .A(p_input[4476]), .B(p_input[4444]), .Z(n28348) );
  XNOR U28066 ( .A(n27453), .B(n28343), .Z(n28345) );
  XOR U28067 ( .A(n28349), .B(n28350), .Z(n27453) );
  AND U28068 ( .A(n400), .B(n28351), .Z(n28350) );
  XOR U28069 ( .A(p_input[4412]), .B(p_input[4380]), .Z(n28351) );
  XOR U28070 ( .A(n28352), .B(n28353), .Z(n28343) );
  AND U28071 ( .A(n28354), .B(n28355), .Z(n28353) );
  XOR U28072 ( .A(n28352), .B(n27468), .Z(n28355) );
  XNOR U28073 ( .A(p_input[4443]), .B(n28356), .Z(n27468) );
  AND U28074 ( .A(n403), .B(n28357), .Z(n28356) );
  XOR U28075 ( .A(p_input[4475]), .B(p_input[4443]), .Z(n28357) );
  XNOR U28076 ( .A(n27465), .B(n28352), .Z(n28354) );
  XOR U28077 ( .A(n28358), .B(n28359), .Z(n27465) );
  AND U28078 ( .A(n400), .B(n28360), .Z(n28359) );
  XOR U28079 ( .A(p_input[4411]), .B(p_input[4379]), .Z(n28360) );
  XOR U28080 ( .A(n28361), .B(n28362), .Z(n28352) );
  AND U28081 ( .A(n28363), .B(n28364), .Z(n28362) );
  XOR U28082 ( .A(n28361), .B(n27480), .Z(n28364) );
  XNOR U28083 ( .A(p_input[4442]), .B(n28365), .Z(n27480) );
  AND U28084 ( .A(n403), .B(n28366), .Z(n28365) );
  XOR U28085 ( .A(p_input[4474]), .B(p_input[4442]), .Z(n28366) );
  XNOR U28086 ( .A(n27477), .B(n28361), .Z(n28363) );
  XOR U28087 ( .A(n28367), .B(n28368), .Z(n27477) );
  AND U28088 ( .A(n400), .B(n28369), .Z(n28368) );
  XOR U28089 ( .A(p_input[4410]), .B(p_input[4378]), .Z(n28369) );
  XOR U28090 ( .A(n28370), .B(n28371), .Z(n28361) );
  AND U28091 ( .A(n28372), .B(n28373), .Z(n28371) );
  XOR U28092 ( .A(n28370), .B(n27492), .Z(n28373) );
  XNOR U28093 ( .A(p_input[4441]), .B(n28374), .Z(n27492) );
  AND U28094 ( .A(n403), .B(n28375), .Z(n28374) );
  XOR U28095 ( .A(p_input[4473]), .B(p_input[4441]), .Z(n28375) );
  XNOR U28096 ( .A(n27489), .B(n28370), .Z(n28372) );
  XOR U28097 ( .A(n28376), .B(n28377), .Z(n27489) );
  AND U28098 ( .A(n400), .B(n28378), .Z(n28377) );
  XOR U28099 ( .A(p_input[4409]), .B(p_input[4377]), .Z(n28378) );
  XOR U28100 ( .A(n28379), .B(n28380), .Z(n28370) );
  AND U28101 ( .A(n28381), .B(n28382), .Z(n28380) );
  XOR U28102 ( .A(n28379), .B(n27504), .Z(n28382) );
  XNOR U28103 ( .A(p_input[4440]), .B(n28383), .Z(n27504) );
  AND U28104 ( .A(n403), .B(n28384), .Z(n28383) );
  XOR U28105 ( .A(p_input[4472]), .B(p_input[4440]), .Z(n28384) );
  XNOR U28106 ( .A(n27501), .B(n28379), .Z(n28381) );
  XOR U28107 ( .A(n28385), .B(n28386), .Z(n27501) );
  AND U28108 ( .A(n400), .B(n28387), .Z(n28386) );
  XOR U28109 ( .A(p_input[4408]), .B(p_input[4376]), .Z(n28387) );
  XOR U28110 ( .A(n28388), .B(n28389), .Z(n28379) );
  AND U28111 ( .A(n28390), .B(n28391), .Z(n28389) );
  XOR U28112 ( .A(n28388), .B(n27516), .Z(n28391) );
  XNOR U28113 ( .A(p_input[4439]), .B(n28392), .Z(n27516) );
  AND U28114 ( .A(n403), .B(n28393), .Z(n28392) );
  XOR U28115 ( .A(p_input[4471]), .B(p_input[4439]), .Z(n28393) );
  XNOR U28116 ( .A(n27513), .B(n28388), .Z(n28390) );
  XOR U28117 ( .A(n28394), .B(n28395), .Z(n27513) );
  AND U28118 ( .A(n400), .B(n28396), .Z(n28395) );
  XOR U28119 ( .A(p_input[4407]), .B(p_input[4375]), .Z(n28396) );
  XOR U28120 ( .A(n28397), .B(n28398), .Z(n28388) );
  AND U28121 ( .A(n28399), .B(n28400), .Z(n28398) );
  XOR U28122 ( .A(n28397), .B(n27528), .Z(n28400) );
  XNOR U28123 ( .A(p_input[4438]), .B(n28401), .Z(n27528) );
  AND U28124 ( .A(n403), .B(n28402), .Z(n28401) );
  XOR U28125 ( .A(p_input[4470]), .B(p_input[4438]), .Z(n28402) );
  XNOR U28126 ( .A(n27525), .B(n28397), .Z(n28399) );
  XOR U28127 ( .A(n28403), .B(n28404), .Z(n27525) );
  AND U28128 ( .A(n400), .B(n28405), .Z(n28404) );
  XOR U28129 ( .A(p_input[4406]), .B(p_input[4374]), .Z(n28405) );
  XOR U28130 ( .A(n28406), .B(n28407), .Z(n28397) );
  AND U28131 ( .A(n28408), .B(n28409), .Z(n28407) );
  XOR U28132 ( .A(n28406), .B(n27540), .Z(n28409) );
  XNOR U28133 ( .A(p_input[4437]), .B(n28410), .Z(n27540) );
  AND U28134 ( .A(n403), .B(n28411), .Z(n28410) );
  XOR U28135 ( .A(p_input[4469]), .B(p_input[4437]), .Z(n28411) );
  XNOR U28136 ( .A(n27537), .B(n28406), .Z(n28408) );
  XOR U28137 ( .A(n28412), .B(n28413), .Z(n27537) );
  AND U28138 ( .A(n400), .B(n28414), .Z(n28413) );
  XOR U28139 ( .A(p_input[4405]), .B(p_input[4373]), .Z(n28414) );
  XOR U28140 ( .A(n28415), .B(n28416), .Z(n28406) );
  AND U28141 ( .A(n28417), .B(n28418), .Z(n28416) );
  XOR U28142 ( .A(n28415), .B(n27552), .Z(n28418) );
  XNOR U28143 ( .A(p_input[4436]), .B(n28419), .Z(n27552) );
  AND U28144 ( .A(n403), .B(n28420), .Z(n28419) );
  XOR U28145 ( .A(p_input[4468]), .B(p_input[4436]), .Z(n28420) );
  XNOR U28146 ( .A(n27549), .B(n28415), .Z(n28417) );
  XOR U28147 ( .A(n28421), .B(n28422), .Z(n27549) );
  AND U28148 ( .A(n400), .B(n28423), .Z(n28422) );
  XOR U28149 ( .A(p_input[4404]), .B(p_input[4372]), .Z(n28423) );
  XOR U28150 ( .A(n28424), .B(n28425), .Z(n28415) );
  AND U28151 ( .A(n28426), .B(n28427), .Z(n28425) );
  XOR U28152 ( .A(n28424), .B(n27564), .Z(n28427) );
  XNOR U28153 ( .A(p_input[4435]), .B(n28428), .Z(n27564) );
  AND U28154 ( .A(n403), .B(n28429), .Z(n28428) );
  XOR U28155 ( .A(p_input[4467]), .B(p_input[4435]), .Z(n28429) );
  XNOR U28156 ( .A(n27561), .B(n28424), .Z(n28426) );
  XOR U28157 ( .A(n28430), .B(n28431), .Z(n27561) );
  AND U28158 ( .A(n400), .B(n28432), .Z(n28431) );
  XOR U28159 ( .A(p_input[4403]), .B(p_input[4371]), .Z(n28432) );
  XOR U28160 ( .A(n28433), .B(n28434), .Z(n28424) );
  AND U28161 ( .A(n28435), .B(n28436), .Z(n28434) );
  XOR U28162 ( .A(n28433), .B(n27576), .Z(n28436) );
  XNOR U28163 ( .A(p_input[4434]), .B(n28437), .Z(n27576) );
  AND U28164 ( .A(n403), .B(n28438), .Z(n28437) );
  XOR U28165 ( .A(p_input[4466]), .B(p_input[4434]), .Z(n28438) );
  XNOR U28166 ( .A(n27573), .B(n28433), .Z(n28435) );
  XOR U28167 ( .A(n28439), .B(n28440), .Z(n27573) );
  AND U28168 ( .A(n400), .B(n28441), .Z(n28440) );
  XOR U28169 ( .A(p_input[4402]), .B(p_input[4370]), .Z(n28441) );
  XOR U28170 ( .A(n28442), .B(n28443), .Z(n28433) );
  AND U28171 ( .A(n28444), .B(n28445), .Z(n28443) );
  XOR U28172 ( .A(n28442), .B(n27588), .Z(n28445) );
  XNOR U28173 ( .A(p_input[4433]), .B(n28446), .Z(n27588) );
  AND U28174 ( .A(n403), .B(n28447), .Z(n28446) );
  XOR U28175 ( .A(p_input[4465]), .B(p_input[4433]), .Z(n28447) );
  XNOR U28176 ( .A(n27585), .B(n28442), .Z(n28444) );
  XOR U28177 ( .A(n28448), .B(n28449), .Z(n27585) );
  AND U28178 ( .A(n400), .B(n28450), .Z(n28449) );
  XOR U28179 ( .A(p_input[4401]), .B(p_input[4369]), .Z(n28450) );
  XOR U28180 ( .A(n28451), .B(n28452), .Z(n28442) );
  AND U28181 ( .A(n28453), .B(n28454), .Z(n28452) );
  XOR U28182 ( .A(n28451), .B(n27600), .Z(n28454) );
  XNOR U28183 ( .A(p_input[4432]), .B(n28455), .Z(n27600) );
  AND U28184 ( .A(n403), .B(n28456), .Z(n28455) );
  XOR U28185 ( .A(p_input[4464]), .B(p_input[4432]), .Z(n28456) );
  XNOR U28186 ( .A(n27597), .B(n28451), .Z(n28453) );
  XOR U28187 ( .A(n28457), .B(n28458), .Z(n27597) );
  AND U28188 ( .A(n400), .B(n28459), .Z(n28458) );
  XOR U28189 ( .A(p_input[4400]), .B(p_input[4368]), .Z(n28459) );
  XOR U28190 ( .A(n28460), .B(n28461), .Z(n28451) );
  AND U28191 ( .A(n28462), .B(n28463), .Z(n28461) );
  XOR U28192 ( .A(n28460), .B(n27612), .Z(n28463) );
  XNOR U28193 ( .A(p_input[4431]), .B(n28464), .Z(n27612) );
  AND U28194 ( .A(n403), .B(n28465), .Z(n28464) );
  XOR U28195 ( .A(p_input[4463]), .B(p_input[4431]), .Z(n28465) );
  XNOR U28196 ( .A(n27609), .B(n28460), .Z(n28462) );
  XOR U28197 ( .A(n28466), .B(n28467), .Z(n27609) );
  AND U28198 ( .A(n400), .B(n28468), .Z(n28467) );
  XOR U28199 ( .A(p_input[4399]), .B(p_input[4367]), .Z(n28468) );
  XOR U28200 ( .A(n28469), .B(n28470), .Z(n28460) );
  AND U28201 ( .A(n28471), .B(n28472), .Z(n28470) );
  XOR U28202 ( .A(n28469), .B(n27624), .Z(n28472) );
  XNOR U28203 ( .A(p_input[4430]), .B(n28473), .Z(n27624) );
  AND U28204 ( .A(n403), .B(n28474), .Z(n28473) );
  XOR U28205 ( .A(p_input[4462]), .B(p_input[4430]), .Z(n28474) );
  XNOR U28206 ( .A(n27621), .B(n28469), .Z(n28471) );
  XOR U28207 ( .A(n28475), .B(n28476), .Z(n27621) );
  AND U28208 ( .A(n400), .B(n28477), .Z(n28476) );
  XOR U28209 ( .A(p_input[4398]), .B(p_input[4366]), .Z(n28477) );
  XOR U28210 ( .A(n28478), .B(n28479), .Z(n28469) );
  AND U28211 ( .A(n28480), .B(n28481), .Z(n28479) );
  XOR U28212 ( .A(n28478), .B(n27636), .Z(n28481) );
  XNOR U28213 ( .A(p_input[4429]), .B(n28482), .Z(n27636) );
  AND U28214 ( .A(n403), .B(n28483), .Z(n28482) );
  XOR U28215 ( .A(p_input[4461]), .B(p_input[4429]), .Z(n28483) );
  XNOR U28216 ( .A(n27633), .B(n28478), .Z(n28480) );
  XOR U28217 ( .A(n28484), .B(n28485), .Z(n27633) );
  AND U28218 ( .A(n400), .B(n28486), .Z(n28485) );
  XOR U28219 ( .A(p_input[4397]), .B(p_input[4365]), .Z(n28486) );
  XOR U28220 ( .A(n28487), .B(n28488), .Z(n28478) );
  AND U28221 ( .A(n28489), .B(n28490), .Z(n28488) );
  XOR U28222 ( .A(n28487), .B(n27648), .Z(n28490) );
  XNOR U28223 ( .A(p_input[4428]), .B(n28491), .Z(n27648) );
  AND U28224 ( .A(n403), .B(n28492), .Z(n28491) );
  XOR U28225 ( .A(p_input[4460]), .B(p_input[4428]), .Z(n28492) );
  XNOR U28226 ( .A(n27645), .B(n28487), .Z(n28489) );
  XOR U28227 ( .A(n28493), .B(n28494), .Z(n27645) );
  AND U28228 ( .A(n400), .B(n28495), .Z(n28494) );
  XOR U28229 ( .A(p_input[4396]), .B(p_input[4364]), .Z(n28495) );
  XOR U28230 ( .A(n28496), .B(n28497), .Z(n28487) );
  AND U28231 ( .A(n28498), .B(n28499), .Z(n28497) );
  XOR U28232 ( .A(n28496), .B(n27660), .Z(n28499) );
  XNOR U28233 ( .A(p_input[4427]), .B(n28500), .Z(n27660) );
  AND U28234 ( .A(n403), .B(n28501), .Z(n28500) );
  XOR U28235 ( .A(p_input[4459]), .B(p_input[4427]), .Z(n28501) );
  XNOR U28236 ( .A(n27657), .B(n28496), .Z(n28498) );
  XOR U28237 ( .A(n28502), .B(n28503), .Z(n27657) );
  AND U28238 ( .A(n400), .B(n28504), .Z(n28503) );
  XOR U28239 ( .A(p_input[4395]), .B(p_input[4363]), .Z(n28504) );
  XOR U28240 ( .A(n28505), .B(n28506), .Z(n28496) );
  AND U28241 ( .A(n28507), .B(n28508), .Z(n28506) );
  XOR U28242 ( .A(n28505), .B(n27672), .Z(n28508) );
  XNOR U28243 ( .A(p_input[4426]), .B(n28509), .Z(n27672) );
  AND U28244 ( .A(n403), .B(n28510), .Z(n28509) );
  XOR U28245 ( .A(p_input[4458]), .B(p_input[4426]), .Z(n28510) );
  XNOR U28246 ( .A(n27669), .B(n28505), .Z(n28507) );
  XOR U28247 ( .A(n28511), .B(n28512), .Z(n27669) );
  AND U28248 ( .A(n400), .B(n28513), .Z(n28512) );
  XOR U28249 ( .A(p_input[4394]), .B(p_input[4362]), .Z(n28513) );
  XOR U28250 ( .A(n28514), .B(n28515), .Z(n28505) );
  AND U28251 ( .A(n28516), .B(n28517), .Z(n28515) );
  XOR U28252 ( .A(n28514), .B(n27684), .Z(n28517) );
  XNOR U28253 ( .A(p_input[4425]), .B(n28518), .Z(n27684) );
  AND U28254 ( .A(n403), .B(n28519), .Z(n28518) );
  XOR U28255 ( .A(p_input[4457]), .B(p_input[4425]), .Z(n28519) );
  XNOR U28256 ( .A(n27681), .B(n28514), .Z(n28516) );
  XOR U28257 ( .A(n28520), .B(n28521), .Z(n27681) );
  AND U28258 ( .A(n400), .B(n28522), .Z(n28521) );
  XOR U28259 ( .A(p_input[4393]), .B(p_input[4361]), .Z(n28522) );
  XOR U28260 ( .A(n28523), .B(n28524), .Z(n28514) );
  AND U28261 ( .A(n28525), .B(n28526), .Z(n28524) );
  XOR U28262 ( .A(n28523), .B(n27696), .Z(n28526) );
  XNOR U28263 ( .A(p_input[4424]), .B(n28527), .Z(n27696) );
  AND U28264 ( .A(n403), .B(n28528), .Z(n28527) );
  XOR U28265 ( .A(p_input[4456]), .B(p_input[4424]), .Z(n28528) );
  XNOR U28266 ( .A(n27693), .B(n28523), .Z(n28525) );
  XOR U28267 ( .A(n28529), .B(n28530), .Z(n27693) );
  AND U28268 ( .A(n400), .B(n28531), .Z(n28530) );
  XOR U28269 ( .A(p_input[4392]), .B(p_input[4360]), .Z(n28531) );
  XOR U28270 ( .A(n28532), .B(n28533), .Z(n28523) );
  AND U28271 ( .A(n28534), .B(n28535), .Z(n28533) );
  XOR U28272 ( .A(n28532), .B(n27708), .Z(n28535) );
  XNOR U28273 ( .A(p_input[4423]), .B(n28536), .Z(n27708) );
  AND U28274 ( .A(n403), .B(n28537), .Z(n28536) );
  XOR U28275 ( .A(p_input[4455]), .B(p_input[4423]), .Z(n28537) );
  XNOR U28276 ( .A(n27705), .B(n28532), .Z(n28534) );
  XOR U28277 ( .A(n28538), .B(n28539), .Z(n27705) );
  AND U28278 ( .A(n400), .B(n28540), .Z(n28539) );
  XOR U28279 ( .A(p_input[4391]), .B(p_input[4359]), .Z(n28540) );
  XOR U28280 ( .A(n28541), .B(n28542), .Z(n28532) );
  AND U28281 ( .A(n28543), .B(n28544), .Z(n28542) );
  XOR U28282 ( .A(n28541), .B(n27720), .Z(n28544) );
  XNOR U28283 ( .A(p_input[4422]), .B(n28545), .Z(n27720) );
  AND U28284 ( .A(n403), .B(n28546), .Z(n28545) );
  XOR U28285 ( .A(p_input[4454]), .B(p_input[4422]), .Z(n28546) );
  XNOR U28286 ( .A(n27717), .B(n28541), .Z(n28543) );
  XOR U28287 ( .A(n28547), .B(n28548), .Z(n27717) );
  AND U28288 ( .A(n400), .B(n28549), .Z(n28548) );
  XOR U28289 ( .A(p_input[4390]), .B(p_input[4358]), .Z(n28549) );
  XOR U28290 ( .A(n28550), .B(n28551), .Z(n28541) );
  AND U28291 ( .A(n28552), .B(n28553), .Z(n28551) );
  XOR U28292 ( .A(n28550), .B(n27732), .Z(n28553) );
  XNOR U28293 ( .A(p_input[4421]), .B(n28554), .Z(n27732) );
  AND U28294 ( .A(n403), .B(n28555), .Z(n28554) );
  XOR U28295 ( .A(p_input[4453]), .B(p_input[4421]), .Z(n28555) );
  XNOR U28296 ( .A(n27729), .B(n28550), .Z(n28552) );
  XOR U28297 ( .A(n28556), .B(n28557), .Z(n27729) );
  AND U28298 ( .A(n400), .B(n28558), .Z(n28557) );
  XOR U28299 ( .A(p_input[4389]), .B(p_input[4357]), .Z(n28558) );
  XOR U28300 ( .A(n28559), .B(n28560), .Z(n28550) );
  AND U28301 ( .A(n28561), .B(n28562), .Z(n28560) );
  XOR U28302 ( .A(n28559), .B(n27744), .Z(n28562) );
  XNOR U28303 ( .A(p_input[4420]), .B(n28563), .Z(n27744) );
  AND U28304 ( .A(n403), .B(n28564), .Z(n28563) );
  XOR U28305 ( .A(p_input[4452]), .B(p_input[4420]), .Z(n28564) );
  XNOR U28306 ( .A(n27741), .B(n28559), .Z(n28561) );
  XOR U28307 ( .A(n28565), .B(n28566), .Z(n27741) );
  AND U28308 ( .A(n400), .B(n28567), .Z(n28566) );
  XOR U28309 ( .A(p_input[4388]), .B(p_input[4356]), .Z(n28567) );
  XOR U28310 ( .A(n28568), .B(n28569), .Z(n28559) );
  AND U28311 ( .A(n28570), .B(n28571), .Z(n28569) );
  XOR U28312 ( .A(n28568), .B(n27756), .Z(n28571) );
  XNOR U28313 ( .A(p_input[4419]), .B(n28572), .Z(n27756) );
  AND U28314 ( .A(n403), .B(n28573), .Z(n28572) );
  XOR U28315 ( .A(p_input[4451]), .B(p_input[4419]), .Z(n28573) );
  XNOR U28316 ( .A(n27753), .B(n28568), .Z(n28570) );
  XOR U28317 ( .A(n28574), .B(n28575), .Z(n27753) );
  AND U28318 ( .A(n400), .B(n28576), .Z(n28575) );
  XOR U28319 ( .A(p_input[4387]), .B(p_input[4355]), .Z(n28576) );
  XOR U28320 ( .A(n28577), .B(n28578), .Z(n28568) );
  AND U28321 ( .A(n28579), .B(n28580), .Z(n28578) );
  XOR U28322 ( .A(n28577), .B(n27768), .Z(n28580) );
  XNOR U28323 ( .A(p_input[4418]), .B(n28581), .Z(n27768) );
  AND U28324 ( .A(n403), .B(n28582), .Z(n28581) );
  XOR U28325 ( .A(p_input[4450]), .B(p_input[4418]), .Z(n28582) );
  XNOR U28326 ( .A(n27765), .B(n28577), .Z(n28579) );
  XOR U28327 ( .A(n28583), .B(n28584), .Z(n27765) );
  AND U28328 ( .A(n400), .B(n28585), .Z(n28584) );
  XOR U28329 ( .A(p_input[4386]), .B(p_input[4354]), .Z(n28585) );
  XOR U28330 ( .A(n28586), .B(n28587), .Z(n28577) );
  AND U28331 ( .A(n28588), .B(n28589), .Z(n28587) );
  XNOR U28332 ( .A(n28590), .B(n27781), .Z(n28589) );
  XNOR U28333 ( .A(p_input[4417]), .B(n28591), .Z(n27781) );
  AND U28334 ( .A(n403), .B(n28592), .Z(n28591) );
  XNOR U28335 ( .A(p_input[4449]), .B(n28593), .Z(n28592) );
  IV U28336 ( .A(p_input[4417]), .Z(n28593) );
  XNOR U28337 ( .A(n27778), .B(n28586), .Z(n28588) );
  XNOR U28338 ( .A(p_input[4353]), .B(n28594), .Z(n27778) );
  AND U28339 ( .A(n400), .B(n28595), .Z(n28594) );
  XOR U28340 ( .A(p_input[4385]), .B(p_input[4353]), .Z(n28595) );
  IV U28341 ( .A(n28590), .Z(n28586) );
  AND U28342 ( .A(n28316), .B(n28319), .Z(n28590) );
  XOR U28343 ( .A(p_input[4416]), .B(n28596), .Z(n28319) );
  AND U28344 ( .A(n403), .B(n28597), .Z(n28596) );
  XOR U28345 ( .A(p_input[4448]), .B(p_input[4416]), .Z(n28597) );
  XOR U28346 ( .A(n28598), .B(n28599), .Z(n403) );
  AND U28347 ( .A(n28600), .B(n28601), .Z(n28599) );
  XNOR U28348 ( .A(p_input[4479]), .B(n28598), .Z(n28601) );
  XOR U28349 ( .A(n28598), .B(p_input[4447]), .Z(n28600) );
  XOR U28350 ( .A(n28602), .B(n28603), .Z(n28598) );
  AND U28351 ( .A(n28604), .B(n28605), .Z(n28603) );
  XNOR U28352 ( .A(p_input[4478]), .B(n28602), .Z(n28605) );
  XOR U28353 ( .A(n28602), .B(p_input[4446]), .Z(n28604) );
  XOR U28354 ( .A(n28606), .B(n28607), .Z(n28602) );
  AND U28355 ( .A(n28608), .B(n28609), .Z(n28607) );
  XNOR U28356 ( .A(p_input[4477]), .B(n28606), .Z(n28609) );
  XOR U28357 ( .A(n28606), .B(p_input[4445]), .Z(n28608) );
  XOR U28358 ( .A(n28610), .B(n28611), .Z(n28606) );
  AND U28359 ( .A(n28612), .B(n28613), .Z(n28611) );
  XNOR U28360 ( .A(p_input[4476]), .B(n28610), .Z(n28613) );
  XOR U28361 ( .A(n28610), .B(p_input[4444]), .Z(n28612) );
  XOR U28362 ( .A(n28614), .B(n28615), .Z(n28610) );
  AND U28363 ( .A(n28616), .B(n28617), .Z(n28615) );
  XNOR U28364 ( .A(p_input[4475]), .B(n28614), .Z(n28617) );
  XOR U28365 ( .A(n28614), .B(p_input[4443]), .Z(n28616) );
  XOR U28366 ( .A(n28618), .B(n28619), .Z(n28614) );
  AND U28367 ( .A(n28620), .B(n28621), .Z(n28619) );
  XNOR U28368 ( .A(p_input[4474]), .B(n28618), .Z(n28621) );
  XOR U28369 ( .A(n28618), .B(p_input[4442]), .Z(n28620) );
  XOR U28370 ( .A(n28622), .B(n28623), .Z(n28618) );
  AND U28371 ( .A(n28624), .B(n28625), .Z(n28623) );
  XNOR U28372 ( .A(p_input[4473]), .B(n28622), .Z(n28625) );
  XOR U28373 ( .A(n28622), .B(p_input[4441]), .Z(n28624) );
  XOR U28374 ( .A(n28626), .B(n28627), .Z(n28622) );
  AND U28375 ( .A(n28628), .B(n28629), .Z(n28627) );
  XNOR U28376 ( .A(p_input[4472]), .B(n28626), .Z(n28629) );
  XOR U28377 ( .A(n28626), .B(p_input[4440]), .Z(n28628) );
  XOR U28378 ( .A(n28630), .B(n28631), .Z(n28626) );
  AND U28379 ( .A(n28632), .B(n28633), .Z(n28631) );
  XNOR U28380 ( .A(p_input[4471]), .B(n28630), .Z(n28633) );
  XOR U28381 ( .A(n28630), .B(p_input[4439]), .Z(n28632) );
  XOR U28382 ( .A(n28634), .B(n28635), .Z(n28630) );
  AND U28383 ( .A(n28636), .B(n28637), .Z(n28635) );
  XNOR U28384 ( .A(p_input[4470]), .B(n28634), .Z(n28637) );
  XOR U28385 ( .A(n28634), .B(p_input[4438]), .Z(n28636) );
  XOR U28386 ( .A(n28638), .B(n28639), .Z(n28634) );
  AND U28387 ( .A(n28640), .B(n28641), .Z(n28639) );
  XNOR U28388 ( .A(p_input[4469]), .B(n28638), .Z(n28641) );
  XOR U28389 ( .A(n28638), .B(p_input[4437]), .Z(n28640) );
  XOR U28390 ( .A(n28642), .B(n28643), .Z(n28638) );
  AND U28391 ( .A(n28644), .B(n28645), .Z(n28643) );
  XNOR U28392 ( .A(p_input[4468]), .B(n28642), .Z(n28645) );
  XOR U28393 ( .A(n28642), .B(p_input[4436]), .Z(n28644) );
  XOR U28394 ( .A(n28646), .B(n28647), .Z(n28642) );
  AND U28395 ( .A(n28648), .B(n28649), .Z(n28647) );
  XNOR U28396 ( .A(p_input[4467]), .B(n28646), .Z(n28649) );
  XOR U28397 ( .A(n28646), .B(p_input[4435]), .Z(n28648) );
  XOR U28398 ( .A(n28650), .B(n28651), .Z(n28646) );
  AND U28399 ( .A(n28652), .B(n28653), .Z(n28651) );
  XNOR U28400 ( .A(p_input[4466]), .B(n28650), .Z(n28653) );
  XOR U28401 ( .A(n28650), .B(p_input[4434]), .Z(n28652) );
  XOR U28402 ( .A(n28654), .B(n28655), .Z(n28650) );
  AND U28403 ( .A(n28656), .B(n28657), .Z(n28655) );
  XNOR U28404 ( .A(p_input[4465]), .B(n28654), .Z(n28657) );
  XOR U28405 ( .A(n28654), .B(p_input[4433]), .Z(n28656) );
  XOR U28406 ( .A(n28658), .B(n28659), .Z(n28654) );
  AND U28407 ( .A(n28660), .B(n28661), .Z(n28659) );
  XNOR U28408 ( .A(p_input[4464]), .B(n28658), .Z(n28661) );
  XOR U28409 ( .A(n28658), .B(p_input[4432]), .Z(n28660) );
  XOR U28410 ( .A(n28662), .B(n28663), .Z(n28658) );
  AND U28411 ( .A(n28664), .B(n28665), .Z(n28663) );
  XNOR U28412 ( .A(p_input[4463]), .B(n28662), .Z(n28665) );
  XOR U28413 ( .A(n28662), .B(p_input[4431]), .Z(n28664) );
  XOR U28414 ( .A(n28666), .B(n28667), .Z(n28662) );
  AND U28415 ( .A(n28668), .B(n28669), .Z(n28667) );
  XNOR U28416 ( .A(p_input[4462]), .B(n28666), .Z(n28669) );
  XOR U28417 ( .A(n28666), .B(p_input[4430]), .Z(n28668) );
  XOR U28418 ( .A(n28670), .B(n28671), .Z(n28666) );
  AND U28419 ( .A(n28672), .B(n28673), .Z(n28671) );
  XNOR U28420 ( .A(p_input[4461]), .B(n28670), .Z(n28673) );
  XOR U28421 ( .A(n28670), .B(p_input[4429]), .Z(n28672) );
  XOR U28422 ( .A(n28674), .B(n28675), .Z(n28670) );
  AND U28423 ( .A(n28676), .B(n28677), .Z(n28675) );
  XNOR U28424 ( .A(p_input[4460]), .B(n28674), .Z(n28677) );
  XOR U28425 ( .A(n28674), .B(p_input[4428]), .Z(n28676) );
  XOR U28426 ( .A(n28678), .B(n28679), .Z(n28674) );
  AND U28427 ( .A(n28680), .B(n28681), .Z(n28679) );
  XNOR U28428 ( .A(p_input[4459]), .B(n28678), .Z(n28681) );
  XOR U28429 ( .A(n28678), .B(p_input[4427]), .Z(n28680) );
  XOR U28430 ( .A(n28682), .B(n28683), .Z(n28678) );
  AND U28431 ( .A(n28684), .B(n28685), .Z(n28683) );
  XNOR U28432 ( .A(p_input[4458]), .B(n28682), .Z(n28685) );
  XOR U28433 ( .A(n28682), .B(p_input[4426]), .Z(n28684) );
  XOR U28434 ( .A(n28686), .B(n28687), .Z(n28682) );
  AND U28435 ( .A(n28688), .B(n28689), .Z(n28687) );
  XNOR U28436 ( .A(p_input[4457]), .B(n28686), .Z(n28689) );
  XOR U28437 ( .A(n28686), .B(p_input[4425]), .Z(n28688) );
  XOR U28438 ( .A(n28690), .B(n28691), .Z(n28686) );
  AND U28439 ( .A(n28692), .B(n28693), .Z(n28691) );
  XNOR U28440 ( .A(p_input[4456]), .B(n28690), .Z(n28693) );
  XOR U28441 ( .A(n28690), .B(p_input[4424]), .Z(n28692) );
  XOR U28442 ( .A(n28694), .B(n28695), .Z(n28690) );
  AND U28443 ( .A(n28696), .B(n28697), .Z(n28695) );
  XNOR U28444 ( .A(p_input[4455]), .B(n28694), .Z(n28697) );
  XOR U28445 ( .A(n28694), .B(p_input[4423]), .Z(n28696) );
  XOR U28446 ( .A(n28698), .B(n28699), .Z(n28694) );
  AND U28447 ( .A(n28700), .B(n28701), .Z(n28699) );
  XNOR U28448 ( .A(p_input[4454]), .B(n28698), .Z(n28701) );
  XOR U28449 ( .A(n28698), .B(p_input[4422]), .Z(n28700) );
  XOR U28450 ( .A(n28702), .B(n28703), .Z(n28698) );
  AND U28451 ( .A(n28704), .B(n28705), .Z(n28703) );
  XNOR U28452 ( .A(p_input[4453]), .B(n28702), .Z(n28705) );
  XOR U28453 ( .A(n28702), .B(p_input[4421]), .Z(n28704) );
  XOR U28454 ( .A(n28706), .B(n28707), .Z(n28702) );
  AND U28455 ( .A(n28708), .B(n28709), .Z(n28707) );
  XNOR U28456 ( .A(p_input[4452]), .B(n28706), .Z(n28709) );
  XOR U28457 ( .A(n28706), .B(p_input[4420]), .Z(n28708) );
  XOR U28458 ( .A(n28710), .B(n28711), .Z(n28706) );
  AND U28459 ( .A(n28712), .B(n28713), .Z(n28711) );
  XNOR U28460 ( .A(p_input[4451]), .B(n28710), .Z(n28713) );
  XOR U28461 ( .A(n28710), .B(p_input[4419]), .Z(n28712) );
  XOR U28462 ( .A(n28714), .B(n28715), .Z(n28710) );
  AND U28463 ( .A(n28716), .B(n28717), .Z(n28715) );
  XNOR U28464 ( .A(p_input[4450]), .B(n28714), .Z(n28717) );
  XOR U28465 ( .A(n28714), .B(p_input[4418]), .Z(n28716) );
  XNOR U28466 ( .A(n28718), .B(n28719), .Z(n28714) );
  AND U28467 ( .A(n28720), .B(n28721), .Z(n28719) );
  XOR U28468 ( .A(p_input[4449]), .B(n28718), .Z(n28721) );
  XNOR U28469 ( .A(p_input[4417]), .B(n28718), .Z(n28720) );
  AND U28470 ( .A(p_input[4448]), .B(n28722), .Z(n28718) );
  IV U28471 ( .A(p_input[4416]), .Z(n28722) );
  XNOR U28472 ( .A(p_input[4352]), .B(n28723), .Z(n28316) );
  AND U28473 ( .A(n400), .B(n28724), .Z(n28723) );
  XOR U28474 ( .A(p_input[4384]), .B(p_input[4352]), .Z(n28724) );
  XOR U28475 ( .A(n28725), .B(n28726), .Z(n400) );
  AND U28476 ( .A(n28727), .B(n28728), .Z(n28726) );
  XNOR U28477 ( .A(p_input[4415]), .B(n28725), .Z(n28728) );
  XOR U28478 ( .A(n28725), .B(p_input[4383]), .Z(n28727) );
  XOR U28479 ( .A(n28729), .B(n28730), .Z(n28725) );
  AND U28480 ( .A(n28731), .B(n28732), .Z(n28730) );
  XNOR U28481 ( .A(p_input[4414]), .B(n28729), .Z(n28732) );
  XNOR U28482 ( .A(n28729), .B(n28331), .Z(n28731) );
  IV U28483 ( .A(p_input[4382]), .Z(n28331) );
  XOR U28484 ( .A(n28733), .B(n28734), .Z(n28729) );
  AND U28485 ( .A(n28735), .B(n28736), .Z(n28734) );
  XNOR U28486 ( .A(p_input[4413]), .B(n28733), .Z(n28736) );
  XNOR U28487 ( .A(n28733), .B(n28340), .Z(n28735) );
  IV U28488 ( .A(p_input[4381]), .Z(n28340) );
  XOR U28489 ( .A(n28737), .B(n28738), .Z(n28733) );
  AND U28490 ( .A(n28739), .B(n28740), .Z(n28738) );
  XNOR U28491 ( .A(p_input[4412]), .B(n28737), .Z(n28740) );
  XNOR U28492 ( .A(n28737), .B(n28349), .Z(n28739) );
  IV U28493 ( .A(p_input[4380]), .Z(n28349) );
  XOR U28494 ( .A(n28741), .B(n28742), .Z(n28737) );
  AND U28495 ( .A(n28743), .B(n28744), .Z(n28742) );
  XNOR U28496 ( .A(p_input[4411]), .B(n28741), .Z(n28744) );
  XNOR U28497 ( .A(n28741), .B(n28358), .Z(n28743) );
  IV U28498 ( .A(p_input[4379]), .Z(n28358) );
  XOR U28499 ( .A(n28745), .B(n28746), .Z(n28741) );
  AND U28500 ( .A(n28747), .B(n28748), .Z(n28746) );
  XNOR U28501 ( .A(p_input[4410]), .B(n28745), .Z(n28748) );
  XNOR U28502 ( .A(n28745), .B(n28367), .Z(n28747) );
  IV U28503 ( .A(p_input[4378]), .Z(n28367) );
  XOR U28504 ( .A(n28749), .B(n28750), .Z(n28745) );
  AND U28505 ( .A(n28751), .B(n28752), .Z(n28750) );
  XNOR U28506 ( .A(p_input[4409]), .B(n28749), .Z(n28752) );
  XNOR U28507 ( .A(n28749), .B(n28376), .Z(n28751) );
  IV U28508 ( .A(p_input[4377]), .Z(n28376) );
  XOR U28509 ( .A(n28753), .B(n28754), .Z(n28749) );
  AND U28510 ( .A(n28755), .B(n28756), .Z(n28754) );
  XNOR U28511 ( .A(p_input[4408]), .B(n28753), .Z(n28756) );
  XNOR U28512 ( .A(n28753), .B(n28385), .Z(n28755) );
  IV U28513 ( .A(p_input[4376]), .Z(n28385) );
  XOR U28514 ( .A(n28757), .B(n28758), .Z(n28753) );
  AND U28515 ( .A(n28759), .B(n28760), .Z(n28758) );
  XNOR U28516 ( .A(p_input[4407]), .B(n28757), .Z(n28760) );
  XNOR U28517 ( .A(n28757), .B(n28394), .Z(n28759) );
  IV U28518 ( .A(p_input[4375]), .Z(n28394) );
  XOR U28519 ( .A(n28761), .B(n28762), .Z(n28757) );
  AND U28520 ( .A(n28763), .B(n28764), .Z(n28762) );
  XNOR U28521 ( .A(p_input[4406]), .B(n28761), .Z(n28764) );
  XNOR U28522 ( .A(n28761), .B(n28403), .Z(n28763) );
  IV U28523 ( .A(p_input[4374]), .Z(n28403) );
  XOR U28524 ( .A(n28765), .B(n28766), .Z(n28761) );
  AND U28525 ( .A(n28767), .B(n28768), .Z(n28766) );
  XNOR U28526 ( .A(p_input[4405]), .B(n28765), .Z(n28768) );
  XNOR U28527 ( .A(n28765), .B(n28412), .Z(n28767) );
  IV U28528 ( .A(p_input[4373]), .Z(n28412) );
  XOR U28529 ( .A(n28769), .B(n28770), .Z(n28765) );
  AND U28530 ( .A(n28771), .B(n28772), .Z(n28770) );
  XNOR U28531 ( .A(p_input[4404]), .B(n28769), .Z(n28772) );
  XNOR U28532 ( .A(n28769), .B(n28421), .Z(n28771) );
  IV U28533 ( .A(p_input[4372]), .Z(n28421) );
  XOR U28534 ( .A(n28773), .B(n28774), .Z(n28769) );
  AND U28535 ( .A(n28775), .B(n28776), .Z(n28774) );
  XNOR U28536 ( .A(p_input[4403]), .B(n28773), .Z(n28776) );
  XNOR U28537 ( .A(n28773), .B(n28430), .Z(n28775) );
  IV U28538 ( .A(p_input[4371]), .Z(n28430) );
  XOR U28539 ( .A(n28777), .B(n28778), .Z(n28773) );
  AND U28540 ( .A(n28779), .B(n28780), .Z(n28778) );
  XNOR U28541 ( .A(p_input[4402]), .B(n28777), .Z(n28780) );
  XNOR U28542 ( .A(n28777), .B(n28439), .Z(n28779) );
  IV U28543 ( .A(p_input[4370]), .Z(n28439) );
  XOR U28544 ( .A(n28781), .B(n28782), .Z(n28777) );
  AND U28545 ( .A(n28783), .B(n28784), .Z(n28782) );
  XNOR U28546 ( .A(p_input[4401]), .B(n28781), .Z(n28784) );
  XNOR U28547 ( .A(n28781), .B(n28448), .Z(n28783) );
  IV U28548 ( .A(p_input[4369]), .Z(n28448) );
  XOR U28549 ( .A(n28785), .B(n28786), .Z(n28781) );
  AND U28550 ( .A(n28787), .B(n28788), .Z(n28786) );
  XNOR U28551 ( .A(p_input[4400]), .B(n28785), .Z(n28788) );
  XNOR U28552 ( .A(n28785), .B(n28457), .Z(n28787) );
  IV U28553 ( .A(p_input[4368]), .Z(n28457) );
  XOR U28554 ( .A(n28789), .B(n28790), .Z(n28785) );
  AND U28555 ( .A(n28791), .B(n28792), .Z(n28790) );
  XNOR U28556 ( .A(p_input[4399]), .B(n28789), .Z(n28792) );
  XNOR U28557 ( .A(n28789), .B(n28466), .Z(n28791) );
  IV U28558 ( .A(p_input[4367]), .Z(n28466) );
  XOR U28559 ( .A(n28793), .B(n28794), .Z(n28789) );
  AND U28560 ( .A(n28795), .B(n28796), .Z(n28794) );
  XNOR U28561 ( .A(p_input[4398]), .B(n28793), .Z(n28796) );
  XNOR U28562 ( .A(n28793), .B(n28475), .Z(n28795) );
  IV U28563 ( .A(p_input[4366]), .Z(n28475) );
  XOR U28564 ( .A(n28797), .B(n28798), .Z(n28793) );
  AND U28565 ( .A(n28799), .B(n28800), .Z(n28798) );
  XNOR U28566 ( .A(p_input[4397]), .B(n28797), .Z(n28800) );
  XNOR U28567 ( .A(n28797), .B(n28484), .Z(n28799) );
  IV U28568 ( .A(p_input[4365]), .Z(n28484) );
  XOR U28569 ( .A(n28801), .B(n28802), .Z(n28797) );
  AND U28570 ( .A(n28803), .B(n28804), .Z(n28802) );
  XNOR U28571 ( .A(p_input[4396]), .B(n28801), .Z(n28804) );
  XNOR U28572 ( .A(n28801), .B(n28493), .Z(n28803) );
  IV U28573 ( .A(p_input[4364]), .Z(n28493) );
  XOR U28574 ( .A(n28805), .B(n28806), .Z(n28801) );
  AND U28575 ( .A(n28807), .B(n28808), .Z(n28806) );
  XNOR U28576 ( .A(p_input[4395]), .B(n28805), .Z(n28808) );
  XNOR U28577 ( .A(n28805), .B(n28502), .Z(n28807) );
  IV U28578 ( .A(p_input[4363]), .Z(n28502) );
  XOR U28579 ( .A(n28809), .B(n28810), .Z(n28805) );
  AND U28580 ( .A(n28811), .B(n28812), .Z(n28810) );
  XNOR U28581 ( .A(p_input[4394]), .B(n28809), .Z(n28812) );
  XNOR U28582 ( .A(n28809), .B(n28511), .Z(n28811) );
  IV U28583 ( .A(p_input[4362]), .Z(n28511) );
  XOR U28584 ( .A(n28813), .B(n28814), .Z(n28809) );
  AND U28585 ( .A(n28815), .B(n28816), .Z(n28814) );
  XNOR U28586 ( .A(p_input[4393]), .B(n28813), .Z(n28816) );
  XNOR U28587 ( .A(n28813), .B(n28520), .Z(n28815) );
  IV U28588 ( .A(p_input[4361]), .Z(n28520) );
  XOR U28589 ( .A(n28817), .B(n28818), .Z(n28813) );
  AND U28590 ( .A(n28819), .B(n28820), .Z(n28818) );
  XNOR U28591 ( .A(p_input[4392]), .B(n28817), .Z(n28820) );
  XNOR U28592 ( .A(n28817), .B(n28529), .Z(n28819) );
  IV U28593 ( .A(p_input[4360]), .Z(n28529) );
  XOR U28594 ( .A(n28821), .B(n28822), .Z(n28817) );
  AND U28595 ( .A(n28823), .B(n28824), .Z(n28822) );
  XNOR U28596 ( .A(p_input[4391]), .B(n28821), .Z(n28824) );
  XNOR U28597 ( .A(n28821), .B(n28538), .Z(n28823) );
  IV U28598 ( .A(p_input[4359]), .Z(n28538) );
  XOR U28599 ( .A(n28825), .B(n28826), .Z(n28821) );
  AND U28600 ( .A(n28827), .B(n28828), .Z(n28826) );
  XNOR U28601 ( .A(p_input[4390]), .B(n28825), .Z(n28828) );
  XNOR U28602 ( .A(n28825), .B(n28547), .Z(n28827) );
  IV U28603 ( .A(p_input[4358]), .Z(n28547) );
  XOR U28604 ( .A(n28829), .B(n28830), .Z(n28825) );
  AND U28605 ( .A(n28831), .B(n28832), .Z(n28830) );
  XNOR U28606 ( .A(p_input[4389]), .B(n28829), .Z(n28832) );
  XNOR U28607 ( .A(n28829), .B(n28556), .Z(n28831) );
  IV U28608 ( .A(p_input[4357]), .Z(n28556) );
  XOR U28609 ( .A(n28833), .B(n28834), .Z(n28829) );
  AND U28610 ( .A(n28835), .B(n28836), .Z(n28834) );
  XNOR U28611 ( .A(p_input[4388]), .B(n28833), .Z(n28836) );
  XNOR U28612 ( .A(n28833), .B(n28565), .Z(n28835) );
  IV U28613 ( .A(p_input[4356]), .Z(n28565) );
  XOR U28614 ( .A(n28837), .B(n28838), .Z(n28833) );
  AND U28615 ( .A(n28839), .B(n28840), .Z(n28838) );
  XNOR U28616 ( .A(p_input[4387]), .B(n28837), .Z(n28840) );
  XNOR U28617 ( .A(n28837), .B(n28574), .Z(n28839) );
  IV U28618 ( .A(p_input[4355]), .Z(n28574) );
  XOR U28619 ( .A(n28841), .B(n28842), .Z(n28837) );
  AND U28620 ( .A(n28843), .B(n28844), .Z(n28842) );
  XNOR U28621 ( .A(p_input[4386]), .B(n28841), .Z(n28844) );
  XNOR U28622 ( .A(n28841), .B(n28583), .Z(n28843) );
  IV U28623 ( .A(p_input[4354]), .Z(n28583) );
  XNOR U28624 ( .A(n28845), .B(n28846), .Z(n28841) );
  AND U28625 ( .A(n28847), .B(n28848), .Z(n28846) );
  XOR U28626 ( .A(p_input[4385]), .B(n28845), .Z(n28848) );
  XNOR U28627 ( .A(p_input[4353]), .B(n28845), .Z(n28847) );
  AND U28628 ( .A(p_input[4384]), .B(n28849), .Z(n28845) );
  IV U28629 ( .A(p_input[4352]), .Z(n28849) );
  XOR U28630 ( .A(n28850), .B(n28851), .Z(n27028) );
  AND U28631 ( .A(n856), .B(n28852), .Z(n28851) );
  XNOR U28632 ( .A(n28853), .B(n28850), .Z(n28852) );
  XOR U28633 ( .A(n28854), .B(n28855), .Z(n856) );
  AND U28634 ( .A(n28856), .B(n28857), .Z(n28855) );
  XOR U28635 ( .A(n28854), .B(n27043), .Z(n28857) );
  XNOR U28636 ( .A(n28858), .B(n28859), .Z(n27043) );
  AND U28637 ( .A(n28860), .B(n543), .Z(n28859) );
  AND U28638 ( .A(n28858), .B(n28861), .Z(n28860) );
  XNOR U28639 ( .A(n27040), .B(n28854), .Z(n28856) );
  XOR U28640 ( .A(n28862), .B(n28863), .Z(n27040) );
  AND U28641 ( .A(n28864), .B(n540), .Z(n28863) );
  NOR U28642 ( .A(n28862), .B(n28865), .Z(n28864) );
  XOR U28643 ( .A(n28866), .B(n28867), .Z(n28854) );
  AND U28644 ( .A(n28868), .B(n28869), .Z(n28867) );
  XOR U28645 ( .A(n28866), .B(n27055), .Z(n28869) );
  XOR U28646 ( .A(n28870), .B(n28871), .Z(n27055) );
  AND U28647 ( .A(n543), .B(n28872), .Z(n28871) );
  XOR U28648 ( .A(n28873), .B(n28870), .Z(n28872) );
  XNOR U28649 ( .A(n27052), .B(n28866), .Z(n28868) );
  XOR U28650 ( .A(n28874), .B(n28875), .Z(n27052) );
  AND U28651 ( .A(n540), .B(n28876), .Z(n28875) );
  XOR U28652 ( .A(n28877), .B(n28874), .Z(n28876) );
  XOR U28653 ( .A(n28878), .B(n28879), .Z(n28866) );
  AND U28654 ( .A(n28880), .B(n28881), .Z(n28879) );
  XOR U28655 ( .A(n28878), .B(n27067), .Z(n28881) );
  XOR U28656 ( .A(n28882), .B(n28883), .Z(n27067) );
  AND U28657 ( .A(n543), .B(n28884), .Z(n28883) );
  XOR U28658 ( .A(n28885), .B(n28882), .Z(n28884) );
  XNOR U28659 ( .A(n27064), .B(n28878), .Z(n28880) );
  XOR U28660 ( .A(n28886), .B(n28887), .Z(n27064) );
  AND U28661 ( .A(n540), .B(n28888), .Z(n28887) );
  XOR U28662 ( .A(n28889), .B(n28886), .Z(n28888) );
  XOR U28663 ( .A(n28890), .B(n28891), .Z(n28878) );
  AND U28664 ( .A(n28892), .B(n28893), .Z(n28891) );
  XOR U28665 ( .A(n28890), .B(n27079), .Z(n28893) );
  XOR U28666 ( .A(n28894), .B(n28895), .Z(n27079) );
  AND U28667 ( .A(n543), .B(n28896), .Z(n28895) );
  XOR U28668 ( .A(n28897), .B(n28894), .Z(n28896) );
  XNOR U28669 ( .A(n27076), .B(n28890), .Z(n28892) );
  XOR U28670 ( .A(n28898), .B(n28899), .Z(n27076) );
  AND U28671 ( .A(n540), .B(n28900), .Z(n28899) );
  XOR U28672 ( .A(n28901), .B(n28898), .Z(n28900) );
  XOR U28673 ( .A(n28902), .B(n28903), .Z(n28890) );
  AND U28674 ( .A(n28904), .B(n28905), .Z(n28903) );
  XOR U28675 ( .A(n28902), .B(n27091), .Z(n28905) );
  XOR U28676 ( .A(n28906), .B(n28907), .Z(n27091) );
  AND U28677 ( .A(n543), .B(n28908), .Z(n28907) );
  XOR U28678 ( .A(n28909), .B(n28906), .Z(n28908) );
  XNOR U28679 ( .A(n27088), .B(n28902), .Z(n28904) );
  XOR U28680 ( .A(n28910), .B(n28911), .Z(n27088) );
  AND U28681 ( .A(n540), .B(n28912), .Z(n28911) );
  XOR U28682 ( .A(n28913), .B(n28910), .Z(n28912) );
  XOR U28683 ( .A(n28914), .B(n28915), .Z(n28902) );
  AND U28684 ( .A(n28916), .B(n28917), .Z(n28915) );
  XOR U28685 ( .A(n28914), .B(n27103), .Z(n28917) );
  XOR U28686 ( .A(n28918), .B(n28919), .Z(n27103) );
  AND U28687 ( .A(n543), .B(n28920), .Z(n28919) );
  XOR U28688 ( .A(n28921), .B(n28918), .Z(n28920) );
  XNOR U28689 ( .A(n27100), .B(n28914), .Z(n28916) );
  XOR U28690 ( .A(n28922), .B(n28923), .Z(n27100) );
  AND U28691 ( .A(n540), .B(n28924), .Z(n28923) );
  XOR U28692 ( .A(n28925), .B(n28922), .Z(n28924) );
  XOR U28693 ( .A(n28926), .B(n28927), .Z(n28914) );
  AND U28694 ( .A(n28928), .B(n28929), .Z(n28927) );
  XOR U28695 ( .A(n28926), .B(n27115), .Z(n28929) );
  XOR U28696 ( .A(n28930), .B(n28931), .Z(n27115) );
  AND U28697 ( .A(n543), .B(n28932), .Z(n28931) );
  XOR U28698 ( .A(n28933), .B(n28930), .Z(n28932) );
  XNOR U28699 ( .A(n27112), .B(n28926), .Z(n28928) );
  XOR U28700 ( .A(n28934), .B(n28935), .Z(n27112) );
  AND U28701 ( .A(n540), .B(n28936), .Z(n28935) );
  XOR U28702 ( .A(n28937), .B(n28934), .Z(n28936) );
  XOR U28703 ( .A(n28938), .B(n28939), .Z(n28926) );
  AND U28704 ( .A(n28940), .B(n28941), .Z(n28939) );
  XOR U28705 ( .A(n28938), .B(n27127), .Z(n28941) );
  XOR U28706 ( .A(n28942), .B(n28943), .Z(n27127) );
  AND U28707 ( .A(n543), .B(n28944), .Z(n28943) );
  XOR U28708 ( .A(n28945), .B(n28942), .Z(n28944) );
  XNOR U28709 ( .A(n27124), .B(n28938), .Z(n28940) );
  XOR U28710 ( .A(n28946), .B(n28947), .Z(n27124) );
  AND U28711 ( .A(n540), .B(n28948), .Z(n28947) );
  XOR U28712 ( .A(n28949), .B(n28946), .Z(n28948) );
  XOR U28713 ( .A(n28950), .B(n28951), .Z(n28938) );
  AND U28714 ( .A(n28952), .B(n28953), .Z(n28951) );
  XOR U28715 ( .A(n28950), .B(n27139), .Z(n28953) );
  XOR U28716 ( .A(n28954), .B(n28955), .Z(n27139) );
  AND U28717 ( .A(n543), .B(n28956), .Z(n28955) );
  XOR U28718 ( .A(n28957), .B(n28954), .Z(n28956) );
  XNOR U28719 ( .A(n27136), .B(n28950), .Z(n28952) );
  XOR U28720 ( .A(n28958), .B(n28959), .Z(n27136) );
  AND U28721 ( .A(n540), .B(n28960), .Z(n28959) );
  XOR U28722 ( .A(n28961), .B(n28958), .Z(n28960) );
  XOR U28723 ( .A(n28962), .B(n28963), .Z(n28950) );
  AND U28724 ( .A(n28964), .B(n28965), .Z(n28963) );
  XOR U28725 ( .A(n28962), .B(n27151), .Z(n28965) );
  XOR U28726 ( .A(n28966), .B(n28967), .Z(n27151) );
  AND U28727 ( .A(n543), .B(n28968), .Z(n28967) );
  XOR U28728 ( .A(n28969), .B(n28966), .Z(n28968) );
  XNOR U28729 ( .A(n27148), .B(n28962), .Z(n28964) );
  XOR U28730 ( .A(n28970), .B(n28971), .Z(n27148) );
  AND U28731 ( .A(n540), .B(n28972), .Z(n28971) );
  XOR U28732 ( .A(n28973), .B(n28970), .Z(n28972) );
  XOR U28733 ( .A(n28974), .B(n28975), .Z(n28962) );
  AND U28734 ( .A(n28976), .B(n28977), .Z(n28975) );
  XOR U28735 ( .A(n28974), .B(n27163), .Z(n28977) );
  XOR U28736 ( .A(n28978), .B(n28979), .Z(n27163) );
  AND U28737 ( .A(n543), .B(n28980), .Z(n28979) );
  XOR U28738 ( .A(n28981), .B(n28978), .Z(n28980) );
  XNOR U28739 ( .A(n27160), .B(n28974), .Z(n28976) );
  XOR U28740 ( .A(n28982), .B(n28983), .Z(n27160) );
  AND U28741 ( .A(n540), .B(n28984), .Z(n28983) );
  XOR U28742 ( .A(n28985), .B(n28982), .Z(n28984) );
  XOR U28743 ( .A(n28986), .B(n28987), .Z(n28974) );
  AND U28744 ( .A(n28988), .B(n28989), .Z(n28987) );
  XOR U28745 ( .A(n28986), .B(n27175), .Z(n28989) );
  XOR U28746 ( .A(n28990), .B(n28991), .Z(n27175) );
  AND U28747 ( .A(n543), .B(n28992), .Z(n28991) );
  XOR U28748 ( .A(n28993), .B(n28990), .Z(n28992) );
  XNOR U28749 ( .A(n27172), .B(n28986), .Z(n28988) );
  XOR U28750 ( .A(n28994), .B(n28995), .Z(n27172) );
  AND U28751 ( .A(n540), .B(n28996), .Z(n28995) );
  XOR U28752 ( .A(n28997), .B(n28994), .Z(n28996) );
  XOR U28753 ( .A(n28998), .B(n28999), .Z(n28986) );
  AND U28754 ( .A(n29000), .B(n29001), .Z(n28999) );
  XOR U28755 ( .A(n28998), .B(n27187), .Z(n29001) );
  XOR U28756 ( .A(n29002), .B(n29003), .Z(n27187) );
  AND U28757 ( .A(n543), .B(n29004), .Z(n29003) );
  XOR U28758 ( .A(n29005), .B(n29002), .Z(n29004) );
  XNOR U28759 ( .A(n27184), .B(n28998), .Z(n29000) );
  XOR U28760 ( .A(n29006), .B(n29007), .Z(n27184) );
  AND U28761 ( .A(n540), .B(n29008), .Z(n29007) );
  XOR U28762 ( .A(n29009), .B(n29006), .Z(n29008) );
  XOR U28763 ( .A(n29010), .B(n29011), .Z(n28998) );
  AND U28764 ( .A(n29012), .B(n29013), .Z(n29011) );
  XOR U28765 ( .A(n29010), .B(n27199), .Z(n29013) );
  XOR U28766 ( .A(n29014), .B(n29015), .Z(n27199) );
  AND U28767 ( .A(n543), .B(n29016), .Z(n29015) );
  XOR U28768 ( .A(n29017), .B(n29014), .Z(n29016) );
  XNOR U28769 ( .A(n27196), .B(n29010), .Z(n29012) );
  XOR U28770 ( .A(n29018), .B(n29019), .Z(n27196) );
  AND U28771 ( .A(n540), .B(n29020), .Z(n29019) );
  XOR U28772 ( .A(n29021), .B(n29018), .Z(n29020) );
  XOR U28773 ( .A(n29022), .B(n29023), .Z(n29010) );
  AND U28774 ( .A(n29024), .B(n29025), .Z(n29023) );
  XOR U28775 ( .A(n29022), .B(n27211), .Z(n29025) );
  XOR U28776 ( .A(n29026), .B(n29027), .Z(n27211) );
  AND U28777 ( .A(n543), .B(n29028), .Z(n29027) );
  XOR U28778 ( .A(n29029), .B(n29026), .Z(n29028) );
  XNOR U28779 ( .A(n27208), .B(n29022), .Z(n29024) );
  XOR U28780 ( .A(n29030), .B(n29031), .Z(n27208) );
  AND U28781 ( .A(n540), .B(n29032), .Z(n29031) );
  XOR U28782 ( .A(n29033), .B(n29030), .Z(n29032) );
  XOR U28783 ( .A(n29034), .B(n29035), .Z(n29022) );
  AND U28784 ( .A(n29036), .B(n29037), .Z(n29035) );
  XOR U28785 ( .A(n29034), .B(n27223), .Z(n29037) );
  XOR U28786 ( .A(n29038), .B(n29039), .Z(n27223) );
  AND U28787 ( .A(n543), .B(n29040), .Z(n29039) );
  XOR U28788 ( .A(n29041), .B(n29038), .Z(n29040) );
  XNOR U28789 ( .A(n27220), .B(n29034), .Z(n29036) );
  XOR U28790 ( .A(n29042), .B(n29043), .Z(n27220) );
  AND U28791 ( .A(n540), .B(n29044), .Z(n29043) );
  XOR U28792 ( .A(n29045), .B(n29042), .Z(n29044) );
  XOR U28793 ( .A(n29046), .B(n29047), .Z(n29034) );
  AND U28794 ( .A(n29048), .B(n29049), .Z(n29047) );
  XOR U28795 ( .A(n29046), .B(n27235), .Z(n29049) );
  XOR U28796 ( .A(n29050), .B(n29051), .Z(n27235) );
  AND U28797 ( .A(n543), .B(n29052), .Z(n29051) );
  XOR U28798 ( .A(n29053), .B(n29050), .Z(n29052) );
  XNOR U28799 ( .A(n27232), .B(n29046), .Z(n29048) );
  XOR U28800 ( .A(n29054), .B(n29055), .Z(n27232) );
  AND U28801 ( .A(n540), .B(n29056), .Z(n29055) );
  XOR U28802 ( .A(n29057), .B(n29054), .Z(n29056) );
  XOR U28803 ( .A(n29058), .B(n29059), .Z(n29046) );
  AND U28804 ( .A(n29060), .B(n29061), .Z(n29059) );
  XOR U28805 ( .A(n29058), .B(n27247), .Z(n29061) );
  XOR U28806 ( .A(n29062), .B(n29063), .Z(n27247) );
  AND U28807 ( .A(n543), .B(n29064), .Z(n29063) );
  XOR U28808 ( .A(n29065), .B(n29062), .Z(n29064) );
  XNOR U28809 ( .A(n27244), .B(n29058), .Z(n29060) );
  XOR U28810 ( .A(n29066), .B(n29067), .Z(n27244) );
  AND U28811 ( .A(n540), .B(n29068), .Z(n29067) );
  XOR U28812 ( .A(n29069), .B(n29066), .Z(n29068) );
  XOR U28813 ( .A(n29070), .B(n29071), .Z(n29058) );
  AND U28814 ( .A(n29072), .B(n29073), .Z(n29071) );
  XOR U28815 ( .A(n29070), .B(n27259), .Z(n29073) );
  XOR U28816 ( .A(n29074), .B(n29075), .Z(n27259) );
  AND U28817 ( .A(n543), .B(n29076), .Z(n29075) );
  XOR U28818 ( .A(n29077), .B(n29074), .Z(n29076) );
  XNOR U28819 ( .A(n27256), .B(n29070), .Z(n29072) );
  XOR U28820 ( .A(n29078), .B(n29079), .Z(n27256) );
  AND U28821 ( .A(n540), .B(n29080), .Z(n29079) );
  XOR U28822 ( .A(n29081), .B(n29078), .Z(n29080) );
  XOR U28823 ( .A(n29082), .B(n29083), .Z(n29070) );
  AND U28824 ( .A(n29084), .B(n29085), .Z(n29083) );
  XOR U28825 ( .A(n29082), .B(n27271), .Z(n29085) );
  XOR U28826 ( .A(n29086), .B(n29087), .Z(n27271) );
  AND U28827 ( .A(n543), .B(n29088), .Z(n29087) );
  XOR U28828 ( .A(n29089), .B(n29086), .Z(n29088) );
  XNOR U28829 ( .A(n27268), .B(n29082), .Z(n29084) );
  XOR U28830 ( .A(n29090), .B(n29091), .Z(n27268) );
  AND U28831 ( .A(n540), .B(n29092), .Z(n29091) );
  XOR U28832 ( .A(n29093), .B(n29090), .Z(n29092) );
  XOR U28833 ( .A(n29094), .B(n29095), .Z(n29082) );
  AND U28834 ( .A(n29096), .B(n29097), .Z(n29095) );
  XOR U28835 ( .A(n29094), .B(n27283), .Z(n29097) );
  XOR U28836 ( .A(n29098), .B(n29099), .Z(n27283) );
  AND U28837 ( .A(n543), .B(n29100), .Z(n29099) );
  XOR U28838 ( .A(n29101), .B(n29098), .Z(n29100) );
  XNOR U28839 ( .A(n27280), .B(n29094), .Z(n29096) );
  XOR U28840 ( .A(n29102), .B(n29103), .Z(n27280) );
  AND U28841 ( .A(n540), .B(n29104), .Z(n29103) );
  XOR U28842 ( .A(n29105), .B(n29102), .Z(n29104) );
  XOR U28843 ( .A(n29106), .B(n29107), .Z(n29094) );
  AND U28844 ( .A(n29108), .B(n29109), .Z(n29107) );
  XOR U28845 ( .A(n29106), .B(n27295), .Z(n29109) );
  XOR U28846 ( .A(n29110), .B(n29111), .Z(n27295) );
  AND U28847 ( .A(n543), .B(n29112), .Z(n29111) );
  XOR U28848 ( .A(n29113), .B(n29110), .Z(n29112) );
  XNOR U28849 ( .A(n27292), .B(n29106), .Z(n29108) );
  XOR U28850 ( .A(n29114), .B(n29115), .Z(n27292) );
  AND U28851 ( .A(n540), .B(n29116), .Z(n29115) );
  XOR U28852 ( .A(n29117), .B(n29114), .Z(n29116) );
  XOR U28853 ( .A(n29118), .B(n29119), .Z(n29106) );
  AND U28854 ( .A(n29120), .B(n29121), .Z(n29119) );
  XOR U28855 ( .A(n29118), .B(n27307), .Z(n29121) );
  XOR U28856 ( .A(n29122), .B(n29123), .Z(n27307) );
  AND U28857 ( .A(n543), .B(n29124), .Z(n29123) );
  XOR U28858 ( .A(n29125), .B(n29122), .Z(n29124) );
  XNOR U28859 ( .A(n27304), .B(n29118), .Z(n29120) );
  XOR U28860 ( .A(n29126), .B(n29127), .Z(n27304) );
  AND U28861 ( .A(n540), .B(n29128), .Z(n29127) );
  XOR U28862 ( .A(n29129), .B(n29126), .Z(n29128) );
  XOR U28863 ( .A(n29130), .B(n29131), .Z(n29118) );
  AND U28864 ( .A(n29132), .B(n29133), .Z(n29131) );
  XOR U28865 ( .A(n29130), .B(n27319), .Z(n29133) );
  XOR U28866 ( .A(n29134), .B(n29135), .Z(n27319) );
  AND U28867 ( .A(n543), .B(n29136), .Z(n29135) );
  XOR U28868 ( .A(n29137), .B(n29134), .Z(n29136) );
  XNOR U28869 ( .A(n27316), .B(n29130), .Z(n29132) );
  XOR U28870 ( .A(n29138), .B(n29139), .Z(n27316) );
  AND U28871 ( .A(n540), .B(n29140), .Z(n29139) );
  XOR U28872 ( .A(n29141), .B(n29138), .Z(n29140) );
  XOR U28873 ( .A(n29142), .B(n29143), .Z(n29130) );
  AND U28874 ( .A(n29144), .B(n29145), .Z(n29143) );
  XOR U28875 ( .A(n29142), .B(n27331), .Z(n29145) );
  XOR U28876 ( .A(n29146), .B(n29147), .Z(n27331) );
  AND U28877 ( .A(n543), .B(n29148), .Z(n29147) );
  XOR U28878 ( .A(n29149), .B(n29146), .Z(n29148) );
  XNOR U28879 ( .A(n27328), .B(n29142), .Z(n29144) );
  XOR U28880 ( .A(n29150), .B(n29151), .Z(n27328) );
  AND U28881 ( .A(n540), .B(n29152), .Z(n29151) );
  XOR U28882 ( .A(n29153), .B(n29150), .Z(n29152) );
  XOR U28883 ( .A(n29154), .B(n29155), .Z(n29142) );
  AND U28884 ( .A(n29156), .B(n29157), .Z(n29155) );
  XOR U28885 ( .A(n29154), .B(n27343), .Z(n29157) );
  XOR U28886 ( .A(n29158), .B(n29159), .Z(n27343) );
  AND U28887 ( .A(n543), .B(n29160), .Z(n29159) );
  XOR U28888 ( .A(n29161), .B(n29158), .Z(n29160) );
  XNOR U28889 ( .A(n27340), .B(n29154), .Z(n29156) );
  XOR U28890 ( .A(n29162), .B(n29163), .Z(n27340) );
  AND U28891 ( .A(n540), .B(n29164), .Z(n29163) );
  XOR U28892 ( .A(n29165), .B(n29162), .Z(n29164) );
  XOR U28893 ( .A(n29166), .B(n29167), .Z(n29154) );
  AND U28894 ( .A(n29168), .B(n29169), .Z(n29167) );
  XOR U28895 ( .A(n29166), .B(n27355), .Z(n29169) );
  XOR U28896 ( .A(n29170), .B(n29171), .Z(n27355) );
  AND U28897 ( .A(n543), .B(n29172), .Z(n29171) );
  XOR U28898 ( .A(n29173), .B(n29170), .Z(n29172) );
  XNOR U28899 ( .A(n27352), .B(n29166), .Z(n29168) );
  XOR U28900 ( .A(n29174), .B(n29175), .Z(n27352) );
  AND U28901 ( .A(n540), .B(n29176), .Z(n29175) );
  XOR U28902 ( .A(n29177), .B(n29174), .Z(n29176) );
  XOR U28903 ( .A(n29178), .B(n29179), .Z(n29166) );
  AND U28904 ( .A(n29180), .B(n29181), .Z(n29179) );
  XOR U28905 ( .A(n29178), .B(n27367), .Z(n29181) );
  XOR U28906 ( .A(n29182), .B(n29183), .Z(n27367) );
  AND U28907 ( .A(n543), .B(n29184), .Z(n29183) );
  XOR U28908 ( .A(n29185), .B(n29182), .Z(n29184) );
  XNOR U28909 ( .A(n27364), .B(n29178), .Z(n29180) );
  XOR U28910 ( .A(n29186), .B(n29187), .Z(n27364) );
  AND U28911 ( .A(n540), .B(n29188), .Z(n29187) );
  XOR U28912 ( .A(n29189), .B(n29186), .Z(n29188) );
  XOR U28913 ( .A(n29190), .B(n29191), .Z(n29178) );
  AND U28914 ( .A(n29192), .B(n29193), .Z(n29191) );
  XOR U28915 ( .A(n29190), .B(n27379), .Z(n29193) );
  XOR U28916 ( .A(n29194), .B(n29195), .Z(n27379) );
  AND U28917 ( .A(n543), .B(n29196), .Z(n29195) );
  XOR U28918 ( .A(n29197), .B(n29194), .Z(n29196) );
  XNOR U28919 ( .A(n27376), .B(n29190), .Z(n29192) );
  XOR U28920 ( .A(n29198), .B(n29199), .Z(n27376) );
  AND U28921 ( .A(n540), .B(n29200), .Z(n29199) );
  XOR U28922 ( .A(n29201), .B(n29198), .Z(n29200) );
  XOR U28923 ( .A(n29202), .B(n29203), .Z(n29190) );
  AND U28924 ( .A(n29204), .B(n29205), .Z(n29203) );
  XOR U28925 ( .A(n29202), .B(n27391), .Z(n29205) );
  XOR U28926 ( .A(n29206), .B(n29207), .Z(n27391) );
  AND U28927 ( .A(n543), .B(n29208), .Z(n29207) );
  XOR U28928 ( .A(n29209), .B(n29206), .Z(n29208) );
  XNOR U28929 ( .A(n27388), .B(n29202), .Z(n29204) );
  XOR U28930 ( .A(n29210), .B(n29211), .Z(n27388) );
  AND U28931 ( .A(n540), .B(n29212), .Z(n29211) );
  XOR U28932 ( .A(n29213), .B(n29210), .Z(n29212) );
  XOR U28933 ( .A(n29214), .B(n29215), .Z(n29202) );
  AND U28934 ( .A(n29216), .B(n29217), .Z(n29215) );
  XNOR U28935 ( .A(n29218), .B(n27404), .Z(n29217) );
  XOR U28936 ( .A(n29219), .B(n29220), .Z(n27404) );
  AND U28937 ( .A(n543), .B(n29221), .Z(n29220) );
  XOR U28938 ( .A(n29219), .B(n29222), .Z(n29221) );
  XNOR U28939 ( .A(n27401), .B(n29214), .Z(n29216) );
  XOR U28940 ( .A(n29223), .B(n29224), .Z(n27401) );
  AND U28941 ( .A(n540), .B(n29225), .Z(n29224) );
  XOR U28942 ( .A(n29223), .B(n29226), .Z(n29225) );
  IV U28943 ( .A(n29218), .Z(n29214) );
  AND U28944 ( .A(n28850), .B(n28853), .Z(n29218) );
  XNOR U28945 ( .A(n29227), .B(n29228), .Z(n28853) );
  AND U28946 ( .A(n543), .B(n29229), .Z(n29228) );
  XNOR U28947 ( .A(n29230), .B(n29227), .Z(n29229) );
  XOR U28948 ( .A(n29231), .B(n29232), .Z(n543) );
  AND U28949 ( .A(n29233), .B(n29234), .Z(n29232) );
  XOR U28950 ( .A(n28861), .B(n29231), .Z(n29234) );
  IV U28951 ( .A(n29235), .Z(n28861) );
  AND U28952 ( .A(p_input[4351]), .B(p_input[4319]), .Z(n29235) );
  XOR U28953 ( .A(n29231), .B(n28858), .Z(n29233) );
  AND U28954 ( .A(p_input[4255]), .B(p_input[4287]), .Z(n28858) );
  XOR U28955 ( .A(n29236), .B(n29237), .Z(n29231) );
  AND U28956 ( .A(n29238), .B(n29239), .Z(n29237) );
  XOR U28957 ( .A(n29236), .B(n28873), .Z(n29239) );
  XNOR U28958 ( .A(p_input[4318]), .B(n29240), .Z(n28873) );
  AND U28959 ( .A(n411), .B(n29241), .Z(n29240) );
  XOR U28960 ( .A(p_input[4350]), .B(p_input[4318]), .Z(n29241) );
  XNOR U28961 ( .A(n28870), .B(n29236), .Z(n29238) );
  XOR U28962 ( .A(n29242), .B(n29243), .Z(n28870) );
  AND U28963 ( .A(n409), .B(n29244), .Z(n29243) );
  XOR U28964 ( .A(p_input[4286]), .B(p_input[4254]), .Z(n29244) );
  XOR U28965 ( .A(n29245), .B(n29246), .Z(n29236) );
  AND U28966 ( .A(n29247), .B(n29248), .Z(n29246) );
  XOR U28967 ( .A(n29245), .B(n28885), .Z(n29248) );
  XNOR U28968 ( .A(p_input[4317]), .B(n29249), .Z(n28885) );
  AND U28969 ( .A(n411), .B(n29250), .Z(n29249) );
  XOR U28970 ( .A(p_input[4349]), .B(p_input[4317]), .Z(n29250) );
  XNOR U28971 ( .A(n28882), .B(n29245), .Z(n29247) );
  XOR U28972 ( .A(n29251), .B(n29252), .Z(n28882) );
  AND U28973 ( .A(n409), .B(n29253), .Z(n29252) );
  XOR U28974 ( .A(p_input[4285]), .B(p_input[4253]), .Z(n29253) );
  XOR U28975 ( .A(n29254), .B(n29255), .Z(n29245) );
  AND U28976 ( .A(n29256), .B(n29257), .Z(n29255) );
  XOR U28977 ( .A(n29254), .B(n28897), .Z(n29257) );
  XNOR U28978 ( .A(p_input[4316]), .B(n29258), .Z(n28897) );
  AND U28979 ( .A(n411), .B(n29259), .Z(n29258) );
  XOR U28980 ( .A(p_input[4348]), .B(p_input[4316]), .Z(n29259) );
  XNOR U28981 ( .A(n28894), .B(n29254), .Z(n29256) );
  XOR U28982 ( .A(n29260), .B(n29261), .Z(n28894) );
  AND U28983 ( .A(n409), .B(n29262), .Z(n29261) );
  XOR U28984 ( .A(p_input[4284]), .B(p_input[4252]), .Z(n29262) );
  XOR U28985 ( .A(n29263), .B(n29264), .Z(n29254) );
  AND U28986 ( .A(n29265), .B(n29266), .Z(n29264) );
  XOR U28987 ( .A(n29263), .B(n28909), .Z(n29266) );
  XNOR U28988 ( .A(p_input[4315]), .B(n29267), .Z(n28909) );
  AND U28989 ( .A(n411), .B(n29268), .Z(n29267) );
  XOR U28990 ( .A(p_input[4347]), .B(p_input[4315]), .Z(n29268) );
  XNOR U28991 ( .A(n28906), .B(n29263), .Z(n29265) );
  XOR U28992 ( .A(n29269), .B(n29270), .Z(n28906) );
  AND U28993 ( .A(n409), .B(n29271), .Z(n29270) );
  XOR U28994 ( .A(p_input[4283]), .B(p_input[4251]), .Z(n29271) );
  XOR U28995 ( .A(n29272), .B(n29273), .Z(n29263) );
  AND U28996 ( .A(n29274), .B(n29275), .Z(n29273) );
  XOR U28997 ( .A(n29272), .B(n28921), .Z(n29275) );
  XNOR U28998 ( .A(p_input[4314]), .B(n29276), .Z(n28921) );
  AND U28999 ( .A(n411), .B(n29277), .Z(n29276) );
  XOR U29000 ( .A(p_input[4346]), .B(p_input[4314]), .Z(n29277) );
  XNOR U29001 ( .A(n28918), .B(n29272), .Z(n29274) );
  XOR U29002 ( .A(n29278), .B(n29279), .Z(n28918) );
  AND U29003 ( .A(n409), .B(n29280), .Z(n29279) );
  XOR U29004 ( .A(p_input[4282]), .B(p_input[4250]), .Z(n29280) );
  XOR U29005 ( .A(n29281), .B(n29282), .Z(n29272) );
  AND U29006 ( .A(n29283), .B(n29284), .Z(n29282) );
  XOR U29007 ( .A(n29281), .B(n28933), .Z(n29284) );
  XNOR U29008 ( .A(p_input[4313]), .B(n29285), .Z(n28933) );
  AND U29009 ( .A(n411), .B(n29286), .Z(n29285) );
  XOR U29010 ( .A(p_input[4345]), .B(p_input[4313]), .Z(n29286) );
  XNOR U29011 ( .A(n28930), .B(n29281), .Z(n29283) );
  XOR U29012 ( .A(n29287), .B(n29288), .Z(n28930) );
  AND U29013 ( .A(n409), .B(n29289), .Z(n29288) );
  XOR U29014 ( .A(p_input[4281]), .B(p_input[4249]), .Z(n29289) );
  XOR U29015 ( .A(n29290), .B(n29291), .Z(n29281) );
  AND U29016 ( .A(n29292), .B(n29293), .Z(n29291) );
  XOR U29017 ( .A(n29290), .B(n28945), .Z(n29293) );
  XNOR U29018 ( .A(p_input[4312]), .B(n29294), .Z(n28945) );
  AND U29019 ( .A(n411), .B(n29295), .Z(n29294) );
  XOR U29020 ( .A(p_input[4344]), .B(p_input[4312]), .Z(n29295) );
  XNOR U29021 ( .A(n28942), .B(n29290), .Z(n29292) );
  XOR U29022 ( .A(n29296), .B(n29297), .Z(n28942) );
  AND U29023 ( .A(n409), .B(n29298), .Z(n29297) );
  XOR U29024 ( .A(p_input[4280]), .B(p_input[4248]), .Z(n29298) );
  XOR U29025 ( .A(n29299), .B(n29300), .Z(n29290) );
  AND U29026 ( .A(n29301), .B(n29302), .Z(n29300) );
  XOR U29027 ( .A(n29299), .B(n28957), .Z(n29302) );
  XNOR U29028 ( .A(p_input[4311]), .B(n29303), .Z(n28957) );
  AND U29029 ( .A(n411), .B(n29304), .Z(n29303) );
  XOR U29030 ( .A(p_input[4343]), .B(p_input[4311]), .Z(n29304) );
  XNOR U29031 ( .A(n28954), .B(n29299), .Z(n29301) );
  XOR U29032 ( .A(n29305), .B(n29306), .Z(n28954) );
  AND U29033 ( .A(n409), .B(n29307), .Z(n29306) );
  XOR U29034 ( .A(p_input[4279]), .B(p_input[4247]), .Z(n29307) );
  XOR U29035 ( .A(n29308), .B(n29309), .Z(n29299) );
  AND U29036 ( .A(n29310), .B(n29311), .Z(n29309) );
  XOR U29037 ( .A(n29308), .B(n28969), .Z(n29311) );
  XNOR U29038 ( .A(p_input[4310]), .B(n29312), .Z(n28969) );
  AND U29039 ( .A(n411), .B(n29313), .Z(n29312) );
  XOR U29040 ( .A(p_input[4342]), .B(p_input[4310]), .Z(n29313) );
  XNOR U29041 ( .A(n28966), .B(n29308), .Z(n29310) );
  XOR U29042 ( .A(n29314), .B(n29315), .Z(n28966) );
  AND U29043 ( .A(n409), .B(n29316), .Z(n29315) );
  XOR U29044 ( .A(p_input[4278]), .B(p_input[4246]), .Z(n29316) );
  XOR U29045 ( .A(n29317), .B(n29318), .Z(n29308) );
  AND U29046 ( .A(n29319), .B(n29320), .Z(n29318) );
  XOR U29047 ( .A(n29317), .B(n28981), .Z(n29320) );
  XNOR U29048 ( .A(p_input[4309]), .B(n29321), .Z(n28981) );
  AND U29049 ( .A(n411), .B(n29322), .Z(n29321) );
  XOR U29050 ( .A(p_input[4341]), .B(p_input[4309]), .Z(n29322) );
  XNOR U29051 ( .A(n28978), .B(n29317), .Z(n29319) );
  XOR U29052 ( .A(n29323), .B(n29324), .Z(n28978) );
  AND U29053 ( .A(n409), .B(n29325), .Z(n29324) );
  XOR U29054 ( .A(p_input[4277]), .B(p_input[4245]), .Z(n29325) );
  XOR U29055 ( .A(n29326), .B(n29327), .Z(n29317) );
  AND U29056 ( .A(n29328), .B(n29329), .Z(n29327) );
  XOR U29057 ( .A(n29326), .B(n28993), .Z(n29329) );
  XNOR U29058 ( .A(p_input[4308]), .B(n29330), .Z(n28993) );
  AND U29059 ( .A(n411), .B(n29331), .Z(n29330) );
  XOR U29060 ( .A(p_input[4340]), .B(p_input[4308]), .Z(n29331) );
  XNOR U29061 ( .A(n28990), .B(n29326), .Z(n29328) );
  XOR U29062 ( .A(n29332), .B(n29333), .Z(n28990) );
  AND U29063 ( .A(n409), .B(n29334), .Z(n29333) );
  XOR U29064 ( .A(p_input[4276]), .B(p_input[4244]), .Z(n29334) );
  XOR U29065 ( .A(n29335), .B(n29336), .Z(n29326) );
  AND U29066 ( .A(n29337), .B(n29338), .Z(n29336) );
  XOR U29067 ( .A(n29335), .B(n29005), .Z(n29338) );
  XNOR U29068 ( .A(p_input[4307]), .B(n29339), .Z(n29005) );
  AND U29069 ( .A(n411), .B(n29340), .Z(n29339) );
  XOR U29070 ( .A(p_input[4339]), .B(p_input[4307]), .Z(n29340) );
  XNOR U29071 ( .A(n29002), .B(n29335), .Z(n29337) );
  XOR U29072 ( .A(n29341), .B(n29342), .Z(n29002) );
  AND U29073 ( .A(n409), .B(n29343), .Z(n29342) );
  XOR U29074 ( .A(p_input[4275]), .B(p_input[4243]), .Z(n29343) );
  XOR U29075 ( .A(n29344), .B(n29345), .Z(n29335) );
  AND U29076 ( .A(n29346), .B(n29347), .Z(n29345) );
  XOR U29077 ( .A(n29344), .B(n29017), .Z(n29347) );
  XNOR U29078 ( .A(p_input[4306]), .B(n29348), .Z(n29017) );
  AND U29079 ( .A(n411), .B(n29349), .Z(n29348) );
  XOR U29080 ( .A(p_input[4338]), .B(p_input[4306]), .Z(n29349) );
  XNOR U29081 ( .A(n29014), .B(n29344), .Z(n29346) );
  XOR U29082 ( .A(n29350), .B(n29351), .Z(n29014) );
  AND U29083 ( .A(n409), .B(n29352), .Z(n29351) );
  XOR U29084 ( .A(p_input[4274]), .B(p_input[4242]), .Z(n29352) );
  XOR U29085 ( .A(n29353), .B(n29354), .Z(n29344) );
  AND U29086 ( .A(n29355), .B(n29356), .Z(n29354) );
  XOR U29087 ( .A(n29353), .B(n29029), .Z(n29356) );
  XNOR U29088 ( .A(p_input[4305]), .B(n29357), .Z(n29029) );
  AND U29089 ( .A(n411), .B(n29358), .Z(n29357) );
  XOR U29090 ( .A(p_input[4337]), .B(p_input[4305]), .Z(n29358) );
  XNOR U29091 ( .A(n29026), .B(n29353), .Z(n29355) );
  XOR U29092 ( .A(n29359), .B(n29360), .Z(n29026) );
  AND U29093 ( .A(n409), .B(n29361), .Z(n29360) );
  XOR U29094 ( .A(p_input[4273]), .B(p_input[4241]), .Z(n29361) );
  XOR U29095 ( .A(n29362), .B(n29363), .Z(n29353) );
  AND U29096 ( .A(n29364), .B(n29365), .Z(n29363) );
  XOR U29097 ( .A(n29362), .B(n29041), .Z(n29365) );
  XNOR U29098 ( .A(p_input[4304]), .B(n29366), .Z(n29041) );
  AND U29099 ( .A(n411), .B(n29367), .Z(n29366) );
  XOR U29100 ( .A(p_input[4336]), .B(p_input[4304]), .Z(n29367) );
  XNOR U29101 ( .A(n29038), .B(n29362), .Z(n29364) );
  XOR U29102 ( .A(n29368), .B(n29369), .Z(n29038) );
  AND U29103 ( .A(n409), .B(n29370), .Z(n29369) );
  XOR U29104 ( .A(p_input[4272]), .B(p_input[4240]), .Z(n29370) );
  XOR U29105 ( .A(n29371), .B(n29372), .Z(n29362) );
  AND U29106 ( .A(n29373), .B(n29374), .Z(n29372) );
  XOR U29107 ( .A(n29371), .B(n29053), .Z(n29374) );
  XNOR U29108 ( .A(p_input[4303]), .B(n29375), .Z(n29053) );
  AND U29109 ( .A(n411), .B(n29376), .Z(n29375) );
  XOR U29110 ( .A(p_input[4335]), .B(p_input[4303]), .Z(n29376) );
  XNOR U29111 ( .A(n29050), .B(n29371), .Z(n29373) );
  XOR U29112 ( .A(n29377), .B(n29378), .Z(n29050) );
  AND U29113 ( .A(n409), .B(n29379), .Z(n29378) );
  XOR U29114 ( .A(p_input[4271]), .B(p_input[4239]), .Z(n29379) );
  XOR U29115 ( .A(n29380), .B(n29381), .Z(n29371) );
  AND U29116 ( .A(n29382), .B(n29383), .Z(n29381) );
  XOR U29117 ( .A(n29380), .B(n29065), .Z(n29383) );
  XNOR U29118 ( .A(p_input[4302]), .B(n29384), .Z(n29065) );
  AND U29119 ( .A(n411), .B(n29385), .Z(n29384) );
  XOR U29120 ( .A(p_input[4334]), .B(p_input[4302]), .Z(n29385) );
  XNOR U29121 ( .A(n29062), .B(n29380), .Z(n29382) );
  XOR U29122 ( .A(n29386), .B(n29387), .Z(n29062) );
  AND U29123 ( .A(n409), .B(n29388), .Z(n29387) );
  XOR U29124 ( .A(p_input[4270]), .B(p_input[4238]), .Z(n29388) );
  XOR U29125 ( .A(n29389), .B(n29390), .Z(n29380) );
  AND U29126 ( .A(n29391), .B(n29392), .Z(n29390) );
  XOR U29127 ( .A(n29389), .B(n29077), .Z(n29392) );
  XNOR U29128 ( .A(p_input[4301]), .B(n29393), .Z(n29077) );
  AND U29129 ( .A(n411), .B(n29394), .Z(n29393) );
  XOR U29130 ( .A(p_input[4333]), .B(p_input[4301]), .Z(n29394) );
  XNOR U29131 ( .A(n29074), .B(n29389), .Z(n29391) );
  XOR U29132 ( .A(n29395), .B(n29396), .Z(n29074) );
  AND U29133 ( .A(n409), .B(n29397), .Z(n29396) );
  XOR U29134 ( .A(p_input[4269]), .B(p_input[4237]), .Z(n29397) );
  XOR U29135 ( .A(n29398), .B(n29399), .Z(n29389) );
  AND U29136 ( .A(n29400), .B(n29401), .Z(n29399) );
  XOR U29137 ( .A(n29398), .B(n29089), .Z(n29401) );
  XNOR U29138 ( .A(p_input[4300]), .B(n29402), .Z(n29089) );
  AND U29139 ( .A(n411), .B(n29403), .Z(n29402) );
  XOR U29140 ( .A(p_input[4332]), .B(p_input[4300]), .Z(n29403) );
  XNOR U29141 ( .A(n29086), .B(n29398), .Z(n29400) );
  XOR U29142 ( .A(n29404), .B(n29405), .Z(n29086) );
  AND U29143 ( .A(n409), .B(n29406), .Z(n29405) );
  XOR U29144 ( .A(p_input[4268]), .B(p_input[4236]), .Z(n29406) );
  XOR U29145 ( .A(n29407), .B(n29408), .Z(n29398) );
  AND U29146 ( .A(n29409), .B(n29410), .Z(n29408) );
  XOR U29147 ( .A(n29407), .B(n29101), .Z(n29410) );
  XNOR U29148 ( .A(p_input[4299]), .B(n29411), .Z(n29101) );
  AND U29149 ( .A(n411), .B(n29412), .Z(n29411) );
  XOR U29150 ( .A(p_input[4331]), .B(p_input[4299]), .Z(n29412) );
  XNOR U29151 ( .A(n29098), .B(n29407), .Z(n29409) );
  XOR U29152 ( .A(n29413), .B(n29414), .Z(n29098) );
  AND U29153 ( .A(n409), .B(n29415), .Z(n29414) );
  XOR U29154 ( .A(p_input[4267]), .B(p_input[4235]), .Z(n29415) );
  XOR U29155 ( .A(n29416), .B(n29417), .Z(n29407) );
  AND U29156 ( .A(n29418), .B(n29419), .Z(n29417) );
  XOR U29157 ( .A(n29416), .B(n29113), .Z(n29419) );
  XNOR U29158 ( .A(p_input[4298]), .B(n29420), .Z(n29113) );
  AND U29159 ( .A(n411), .B(n29421), .Z(n29420) );
  XOR U29160 ( .A(p_input[4330]), .B(p_input[4298]), .Z(n29421) );
  XNOR U29161 ( .A(n29110), .B(n29416), .Z(n29418) );
  XOR U29162 ( .A(n29422), .B(n29423), .Z(n29110) );
  AND U29163 ( .A(n409), .B(n29424), .Z(n29423) );
  XOR U29164 ( .A(p_input[4266]), .B(p_input[4234]), .Z(n29424) );
  XOR U29165 ( .A(n29425), .B(n29426), .Z(n29416) );
  AND U29166 ( .A(n29427), .B(n29428), .Z(n29426) );
  XOR U29167 ( .A(n29425), .B(n29125), .Z(n29428) );
  XNOR U29168 ( .A(p_input[4297]), .B(n29429), .Z(n29125) );
  AND U29169 ( .A(n411), .B(n29430), .Z(n29429) );
  XOR U29170 ( .A(p_input[4329]), .B(p_input[4297]), .Z(n29430) );
  XNOR U29171 ( .A(n29122), .B(n29425), .Z(n29427) );
  XOR U29172 ( .A(n29431), .B(n29432), .Z(n29122) );
  AND U29173 ( .A(n409), .B(n29433), .Z(n29432) );
  XOR U29174 ( .A(p_input[4265]), .B(p_input[4233]), .Z(n29433) );
  XOR U29175 ( .A(n29434), .B(n29435), .Z(n29425) );
  AND U29176 ( .A(n29436), .B(n29437), .Z(n29435) );
  XOR U29177 ( .A(n29434), .B(n29137), .Z(n29437) );
  XNOR U29178 ( .A(p_input[4296]), .B(n29438), .Z(n29137) );
  AND U29179 ( .A(n411), .B(n29439), .Z(n29438) );
  XOR U29180 ( .A(p_input[4328]), .B(p_input[4296]), .Z(n29439) );
  XNOR U29181 ( .A(n29134), .B(n29434), .Z(n29436) );
  XOR U29182 ( .A(n29440), .B(n29441), .Z(n29134) );
  AND U29183 ( .A(n409), .B(n29442), .Z(n29441) );
  XOR U29184 ( .A(p_input[4264]), .B(p_input[4232]), .Z(n29442) );
  XOR U29185 ( .A(n29443), .B(n29444), .Z(n29434) );
  AND U29186 ( .A(n29445), .B(n29446), .Z(n29444) );
  XOR U29187 ( .A(n29443), .B(n29149), .Z(n29446) );
  XNOR U29188 ( .A(p_input[4295]), .B(n29447), .Z(n29149) );
  AND U29189 ( .A(n411), .B(n29448), .Z(n29447) );
  XOR U29190 ( .A(p_input[4327]), .B(p_input[4295]), .Z(n29448) );
  XNOR U29191 ( .A(n29146), .B(n29443), .Z(n29445) );
  XOR U29192 ( .A(n29449), .B(n29450), .Z(n29146) );
  AND U29193 ( .A(n409), .B(n29451), .Z(n29450) );
  XOR U29194 ( .A(p_input[4263]), .B(p_input[4231]), .Z(n29451) );
  XOR U29195 ( .A(n29452), .B(n29453), .Z(n29443) );
  AND U29196 ( .A(n29454), .B(n29455), .Z(n29453) );
  XOR U29197 ( .A(n29452), .B(n29161), .Z(n29455) );
  XNOR U29198 ( .A(p_input[4294]), .B(n29456), .Z(n29161) );
  AND U29199 ( .A(n411), .B(n29457), .Z(n29456) );
  XOR U29200 ( .A(p_input[4326]), .B(p_input[4294]), .Z(n29457) );
  XNOR U29201 ( .A(n29158), .B(n29452), .Z(n29454) );
  XOR U29202 ( .A(n29458), .B(n29459), .Z(n29158) );
  AND U29203 ( .A(n409), .B(n29460), .Z(n29459) );
  XOR U29204 ( .A(p_input[4262]), .B(p_input[4230]), .Z(n29460) );
  XOR U29205 ( .A(n29461), .B(n29462), .Z(n29452) );
  AND U29206 ( .A(n29463), .B(n29464), .Z(n29462) );
  XOR U29207 ( .A(n29461), .B(n29173), .Z(n29464) );
  XNOR U29208 ( .A(p_input[4293]), .B(n29465), .Z(n29173) );
  AND U29209 ( .A(n411), .B(n29466), .Z(n29465) );
  XOR U29210 ( .A(p_input[4325]), .B(p_input[4293]), .Z(n29466) );
  XNOR U29211 ( .A(n29170), .B(n29461), .Z(n29463) );
  XOR U29212 ( .A(n29467), .B(n29468), .Z(n29170) );
  AND U29213 ( .A(n409), .B(n29469), .Z(n29468) );
  XOR U29214 ( .A(p_input[4261]), .B(p_input[4229]), .Z(n29469) );
  XOR U29215 ( .A(n29470), .B(n29471), .Z(n29461) );
  AND U29216 ( .A(n29472), .B(n29473), .Z(n29471) );
  XOR U29217 ( .A(n29470), .B(n29185), .Z(n29473) );
  XNOR U29218 ( .A(p_input[4292]), .B(n29474), .Z(n29185) );
  AND U29219 ( .A(n411), .B(n29475), .Z(n29474) );
  XOR U29220 ( .A(p_input[4324]), .B(p_input[4292]), .Z(n29475) );
  XNOR U29221 ( .A(n29182), .B(n29470), .Z(n29472) );
  XOR U29222 ( .A(n29476), .B(n29477), .Z(n29182) );
  AND U29223 ( .A(n409), .B(n29478), .Z(n29477) );
  XOR U29224 ( .A(p_input[4260]), .B(p_input[4228]), .Z(n29478) );
  XOR U29225 ( .A(n29479), .B(n29480), .Z(n29470) );
  AND U29226 ( .A(n29481), .B(n29482), .Z(n29480) );
  XOR U29227 ( .A(n29479), .B(n29197), .Z(n29482) );
  XNOR U29228 ( .A(p_input[4291]), .B(n29483), .Z(n29197) );
  AND U29229 ( .A(n411), .B(n29484), .Z(n29483) );
  XOR U29230 ( .A(p_input[4323]), .B(p_input[4291]), .Z(n29484) );
  XNOR U29231 ( .A(n29194), .B(n29479), .Z(n29481) );
  XOR U29232 ( .A(n29485), .B(n29486), .Z(n29194) );
  AND U29233 ( .A(n409), .B(n29487), .Z(n29486) );
  XOR U29234 ( .A(p_input[4259]), .B(p_input[4227]), .Z(n29487) );
  XOR U29235 ( .A(n29488), .B(n29489), .Z(n29479) );
  AND U29236 ( .A(n29490), .B(n29491), .Z(n29489) );
  XOR U29237 ( .A(n29488), .B(n29209), .Z(n29491) );
  XNOR U29238 ( .A(p_input[4290]), .B(n29492), .Z(n29209) );
  AND U29239 ( .A(n411), .B(n29493), .Z(n29492) );
  XOR U29240 ( .A(p_input[4322]), .B(p_input[4290]), .Z(n29493) );
  XNOR U29241 ( .A(n29206), .B(n29488), .Z(n29490) );
  XOR U29242 ( .A(n29494), .B(n29495), .Z(n29206) );
  AND U29243 ( .A(n409), .B(n29496), .Z(n29495) );
  XOR U29244 ( .A(p_input[4258]), .B(p_input[4226]), .Z(n29496) );
  XOR U29245 ( .A(n29497), .B(n29498), .Z(n29488) );
  AND U29246 ( .A(n29499), .B(n29500), .Z(n29498) );
  XNOR U29247 ( .A(n29501), .B(n29222), .Z(n29500) );
  XNOR U29248 ( .A(p_input[4289]), .B(n29502), .Z(n29222) );
  AND U29249 ( .A(n411), .B(n29503), .Z(n29502) );
  XNOR U29250 ( .A(p_input[4321]), .B(n29504), .Z(n29503) );
  IV U29251 ( .A(p_input[4289]), .Z(n29504) );
  XNOR U29252 ( .A(n29219), .B(n29497), .Z(n29499) );
  XNOR U29253 ( .A(p_input[4225]), .B(n29505), .Z(n29219) );
  AND U29254 ( .A(n409), .B(n29506), .Z(n29505) );
  XOR U29255 ( .A(p_input[4257]), .B(p_input[4225]), .Z(n29506) );
  IV U29256 ( .A(n29501), .Z(n29497) );
  AND U29257 ( .A(n29227), .B(n29230), .Z(n29501) );
  XOR U29258 ( .A(p_input[4288]), .B(n29507), .Z(n29230) );
  AND U29259 ( .A(n411), .B(n29508), .Z(n29507) );
  XOR U29260 ( .A(p_input[4320]), .B(p_input[4288]), .Z(n29508) );
  XOR U29261 ( .A(n29509), .B(n29510), .Z(n411) );
  AND U29262 ( .A(n29511), .B(n29512), .Z(n29510) );
  XNOR U29263 ( .A(p_input[4351]), .B(n29509), .Z(n29512) );
  XOR U29264 ( .A(n29509), .B(p_input[4319]), .Z(n29511) );
  XOR U29265 ( .A(n29513), .B(n29514), .Z(n29509) );
  AND U29266 ( .A(n29515), .B(n29516), .Z(n29514) );
  XNOR U29267 ( .A(p_input[4350]), .B(n29513), .Z(n29516) );
  XOR U29268 ( .A(n29513), .B(p_input[4318]), .Z(n29515) );
  XOR U29269 ( .A(n29517), .B(n29518), .Z(n29513) );
  AND U29270 ( .A(n29519), .B(n29520), .Z(n29518) );
  XNOR U29271 ( .A(p_input[4349]), .B(n29517), .Z(n29520) );
  XOR U29272 ( .A(n29517), .B(p_input[4317]), .Z(n29519) );
  XOR U29273 ( .A(n29521), .B(n29522), .Z(n29517) );
  AND U29274 ( .A(n29523), .B(n29524), .Z(n29522) );
  XNOR U29275 ( .A(p_input[4348]), .B(n29521), .Z(n29524) );
  XOR U29276 ( .A(n29521), .B(p_input[4316]), .Z(n29523) );
  XOR U29277 ( .A(n29525), .B(n29526), .Z(n29521) );
  AND U29278 ( .A(n29527), .B(n29528), .Z(n29526) );
  XNOR U29279 ( .A(p_input[4347]), .B(n29525), .Z(n29528) );
  XOR U29280 ( .A(n29525), .B(p_input[4315]), .Z(n29527) );
  XOR U29281 ( .A(n29529), .B(n29530), .Z(n29525) );
  AND U29282 ( .A(n29531), .B(n29532), .Z(n29530) );
  XNOR U29283 ( .A(p_input[4346]), .B(n29529), .Z(n29532) );
  XOR U29284 ( .A(n29529), .B(p_input[4314]), .Z(n29531) );
  XOR U29285 ( .A(n29533), .B(n29534), .Z(n29529) );
  AND U29286 ( .A(n29535), .B(n29536), .Z(n29534) );
  XNOR U29287 ( .A(p_input[4345]), .B(n29533), .Z(n29536) );
  XOR U29288 ( .A(n29533), .B(p_input[4313]), .Z(n29535) );
  XOR U29289 ( .A(n29537), .B(n29538), .Z(n29533) );
  AND U29290 ( .A(n29539), .B(n29540), .Z(n29538) );
  XNOR U29291 ( .A(p_input[4344]), .B(n29537), .Z(n29540) );
  XOR U29292 ( .A(n29537), .B(p_input[4312]), .Z(n29539) );
  XOR U29293 ( .A(n29541), .B(n29542), .Z(n29537) );
  AND U29294 ( .A(n29543), .B(n29544), .Z(n29542) );
  XNOR U29295 ( .A(p_input[4343]), .B(n29541), .Z(n29544) );
  XOR U29296 ( .A(n29541), .B(p_input[4311]), .Z(n29543) );
  XOR U29297 ( .A(n29545), .B(n29546), .Z(n29541) );
  AND U29298 ( .A(n29547), .B(n29548), .Z(n29546) );
  XNOR U29299 ( .A(p_input[4342]), .B(n29545), .Z(n29548) );
  XOR U29300 ( .A(n29545), .B(p_input[4310]), .Z(n29547) );
  XOR U29301 ( .A(n29549), .B(n29550), .Z(n29545) );
  AND U29302 ( .A(n29551), .B(n29552), .Z(n29550) );
  XNOR U29303 ( .A(p_input[4341]), .B(n29549), .Z(n29552) );
  XOR U29304 ( .A(n29549), .B(p_input[4309]), .Z(n29551) );
  XOR U29305 ( .A(n29553), .B(n29554), .Z(n29549) );
  AND U29306 ( .A(n29555), .B(n29556), .Z(n29554) );
  XNOR U29307 ( .A(p_input[4340]), .B(n29553), .Z(n29556) );
  XOR U29308 ( .A(n29553), .B(p_input[4308]), .Z(n29555) );
  XOR U29309 ( .A(n29557), .B(n29558), .Z(n29553) );
  AND U29310 ( .A(n29559), .B(n29560), .Z(n29558) );
  XNOR U29311 ( .A(p_input[4339]), .B(n29557), .Z(n29560) );
  XOR U29312 ( .A(n29557), .B(p_input[4307]), .Z(n29559) );
  XOR U29313 ( .A(n29561), .B(n29562), .Z(n29557) );
  AND U29314 ( .A(n29563), .B(n29564), .Z(n29562) );
  XNOR U29315 ( .A(p_input[4338]), .B(n29561), .Z(n29564) );
  XOR U29316 ( .A(n29561), .B(p_input[4306]), .Z(n29563) );
  XOR U29317 ( .A(n29565), .B(n29566), .Z(n29561) );
  AND U29318 ( .A(n29567), .B(n29568), .Z(n29566) );
  XNOR U29319 ( .A(p_input[4337]), .B(n29565), .Z(n29568) );
  XOR U29320 ( .A(n29565), .B(p_input[4305]), .Z(n29567) );
  XOR U29321 ( .A(n29569), .B(n29570), .Z(n29565) );
  AND U29322 ( .A(n29571), .B(n29572), .Z(n29570) );
  XNOR U29323 ( .A(p_input[4336]), .B(n29569), .Z(n29572) );
  XOR U29324 ( .A(n29569), .B(p_input[4304]), .Z(n29571) );
  XOR U29325 ( .A(n29573), .B(n29574), .Z(n29569) );
  AND U29326 ( .A(n29575), .B(n29576), .Z(n29574) );
  XNOR U29327 ( .A(p_input[4335]), .B(n29573), .Z(n29576) );
  XOR U29328 ( .A(n29573), .B(p_input[4303]), .Z(n29575) );
  XOR U29329 ( .A(n29577), .B(n29578), .Z(n29573) );
  AND U29330 ( .A(n29579), .B(n29580), .Z(n29578) );
  XNOR U29331 ( .A(p_input[4334]), .B(n29577), .Z(n29580) );
  XOR U29332 ( .A(n29577), .B(p_input[4302]), .Z(n29579) );
  XOR U29333 ( .A(n29581), .B(n29582), .Z(n29577) );
  AND U29334 ( .A(n29583), .B(n29584), .Z(n29582) );
  XNOR U29335 ( .A(p_input[4333]), .B(n29581), .Z(n29584) );
  XOR U29336 ( .A(n29581), .B(p_input[4301]), .Z(n29583) );
  XOR U29337 ( .A(n29585), .B(n29586), .Z(n29581) );
  AND U29338 ( .A(n29587), .B(n29588), .Z(n29586) );
  XNOR U29339 ( .A(p_input[4332]), .B(n29585), .Z(n29588) );
  XOR U29340 ( .A(n29585), .B(p_input[4300]), .Z(n29587) );
  XOR U29341 ( .A(n29589), .B(n29590), .Z(n29585) );
  AND U29342 ( .A(n29591), .B(n29592), .Z(n29590) );
  XNOR U29343 ( .A(p_input[4331]), .B(n29589), .Z(n29592) );
  XOR U29344 ( .A(n29589), .B(p_input[4299]), .Z(n29591) );
  XOR U29345 ( .A(n29593), .B(n29594), .Z(n29589) );
  AND U29346 ( .A(n29595), .B(n29596), .Z(n29594) );
  XNOR U29347 ( .A(p_input[4330]), .B(n29593), .Z(n29596) );
  XOR U29348 ( .A(n29593), .B(p_input[4298]), .Z(n29595) );
  XOR U29349 ( .A(n29597), .B(n29598), .Z(n29593) );
  AND U29350 ( .A(n29599), .B(n29600), .Z(n29598) );
  XNOR U29351 ( .A(p_input[4329]), .B(n29597), .Z(n29600) );
  XOR U29352 ( .A(n29597), .B(p_input[4297]), .Z(n29599) );
  XOR U29353 ( .A(n29601), .B(n29602), .Z(n29597) );
  AND U29354 ( .A(n29603), .B(n29604), .Z(n29602) );
  XNOR U29355 ( .A(p_input[4328]), .B(n29601), .Z(n29604) );
  XOR U29356 ( .A(n29601), .B(p_input[4296]), .Z(n29603) );
  XOR U29357 ( .A(n29605), .B(n29606), .Z(n29601) );
  AND U29358 ( .A(n29607), .B(n29608), .Z(n29606) );
  XNOR U29359 ( .A(p_input[4327]), .B(n29605), .Z(n29608) );
  XOR U29360 ( .A(n29605), .B(p_input[4295]), .Z(n29607) );
  XOR U29361 ( .A(n29609), .B(n29610), .Z(n29605) );
  AND U29362 ( .A(n29611), .B(n29612), .Z(n29610) );
  XNOR U29363 ( .A(p_input[4326]), .B(n29609), .Z(n29612) );
  XOR U29364 ( .A(n29609), .B(p_input[4294]), .Z(n29611) );
  XOR U29365 ( .A(n29613), .B(n29614), .Z(n29609) );
  AND U29366 ( .A(n29615), .B(n29616), .Z(n29614) );
  XNOR U29367 ( .A(p_input[4325]), .B(n29613), .Z(n29616) );
  XOR U29368 ( .A(n29613), .B(p_input[4293]), .Z(n29615) );
  XOR U29369 ( .A(n29617), .B(n29618), .Z(n29613) );
  AND U29370 ( .A(n29619), .B(n29620), .Z(n29618) );
  XNOR U29371 ( .A(p_input[4324]), .B(n29617), .Z(n29620) );
  XOR U29372 ( .A(n29617), .B(p_input[4292]), .Z(n29619) );
  XOR U29373 ( .A(n29621), .B(n29622), .Z(n29617) );
  AND U29374 ( .A(n29623), .B(n29624), .Z(n29622) );
  XNOR U29375 ( .A(p_input[4323]), .B(n29621), .Z(n29624) );
  XOR U29376 ( .A(n29621), .B(p_input[4291]), .Z(n29623) );
  XOR U29377 ( .A(n29625), .B(n29626), .Z(n29621) );
  AND U29378 ( .A(n29627), .B(n29628), .Z(n29626) );
  XNOR U29379 ( .A(p_input[4322]), .B(n29625), .Z(n29628) );
  XOR U29380 ( .A(n29625), .B(p_input[4290]), .Z(n29627) );
  XNOR U29381 ( .A(n29629), .B(n29630), .Z(n29625) );
  AND U29382 ( .A(n29631), .B(n29632), .Z(n29630) );
  XOR U29383 ( .A(p_input[4321]), .B(n29629), .Z(n29632) );
  XNOR U29384 ( .A(p_input[4289]), .B(n29629), .Z(n29631) );
  AND U29385 ( .A(p_input[4320]), .B(n29633), .Z(n29629) );
  IV U29386 ( .A(p_input[4288]), .Z(n29633) );
  XNOR U29387 ( .A(p_input[4224]), .B(n29634), .Z(n29227) );
  AND U29388 ( .A(n409), .B(n29635), .Z(n29634) );
  XOR U29389 ( .A(p_input[4256]), .B(p_input[4224]), .Z(n29635) );
  XOR U29390 ( .A(n29636), .B(n29637), .Z(n409) );
  AND U29391 ( .A(n29638), .B(n29639), .Z(n29637) );
  XNOR U29392 ( .A(p_input[4287]), .B(n29636), .Z(n29639) );
  XOR U29393 ( .A(n29636), .B(p_input[4255]), .Z(n29638) );
  XOR U29394 ( .A(n29640), .B(n29641), .Z(n29636) );
  AND U29395 ( .A(n29642), .B(n29643), .Z(n29641) );
  XNOR U29396 ( .A(p_input[4286]), .B(n29640), .Z(n29643) );
  XNOR U29397 ( .A(n29640), .B(n29242), .Z(n29642) );
  IV U29398 ( .A(p_input[4254]), .Z(n29242) );
  XOR U29399 ( .A(n29644), .B(n29645), .Z(n29640) );
  AND U29400 ( .A(n29646), .B(n29647), .Z(n29645) );
  XNOR U29401 ( .A(p_input[4285]), .B(n29644), .Z(n29647) );
  XNOR U29402 ( .A(n29644), .B(n29251), .Z(n29646) );
  IV U29403 ( .A(p_input[4253]), .Z(n29251) );
  XOR U29404 ( .A(n29648), .B(n29649), .Z(n29644) );
  AND U29405 ( .A(n29650), .B(n29651), .Z(n29649) );
  XNOR U29406 ( .A(p_input[4284]), .B(n29648), .Z(n29651) );
  XNOR U29407 ( .A(n29648), .B(n29260), .Z(n29650) );
  IV U29408 ( .A(p_input[4252]), .Z(n29260) );
  XOR U29409 ( .A(n29652), .B(n29653), .Z(n29648) );
  AND U29410 ( .A(n29654), .B(n29655), .Z(n29653) );
  XNOR U29411 ( .A(p_input[4283]), .B(n29652), .Z(n29655) );
  XNOR U29412 ( .A(n29652), .B(n29269), .Z(n29654) );
  IV U29413 ( .A(p_input[4251]), .Z(n29269) );
  XOR U29414 ( .A(n29656), .B(n29657), .Z(n29652) );
  AND U29415 ( .A(n29658), .B(n29659), .Z(n29657) );
  XNOR U29416 ( .A(p_input[4282]), .B(n29656), .Z(n29659) );
  XNOR U29417 ( .A(n29656), .B(n29278), .Z(n29658) );
  IV U29418 ( .A(p_input[4250]), .Z(n29278) );
  XOR U29419 ( .A(n29660), .B(n29661), .Z(n29656) );
  AND U29420 ( .A(n29662), .B(n29663), .Z(n29661) );
  XNOR U29421 ( .A(p_input[4281]), .B(n29660), .Z(n29663) );
  XNOR U29422 ( .A(n29660), .B(n29287), .Z(n29662) );
  IV U29423 ( .A(p_input[4249]), .Z(n29287) );
  XOR U29424 ( .A(n29664), .B(n29665), .Z(n29660) );
  AND U29425 ( .A(n29666), .B(n29667), .Z(n29665) );
  XNOR U29426 ( .A(p_input[4280]), .B(n29664), .Z(n29667) );
  XNOR U29427 ( .A(n29664), .B(n29296), .Z(n29666) );
  IV U29428 ( .A(p_input[4248]), .Z(n29296) );
  XOR U29429 ( .A(n29668), .B(n29669), .Z(n29664) );
  AND U29430 ( .A(n29670), .B(n29671), .Z(n29669) );
  XNOR U29431 ( .A(p_input[4279]), .B(n29668), .Z(n29671) );
  XNOR U29432 ( .A(n29668), .B(n29305), .Z(n29670) );
  IV U29433 ( .A(p_input[4247]), .Z(n29305) );
  XOR U29434 ( .A(n29672), .B(n29673), .Z(n29668) );
  AND U29435 ( .A(n29674), .B(n29675), .Z(n29673) );
  XNOR U29436 ( .A(p_input[4278]), .B(n29672), .Z(n29675) );
  XNOR U29437 ( .A(n29672), .B(n29314), .Z(n29674) );
  IV U29438 ( .A(p_input[4246]), .Z(n29314) );
  XOR U29439 ( .A(n29676), .B(n29677), .Z(n29672) );
  AND U29440 ( .A(n29678), .B(n29679), .Z(n29677) );
  XNOR U29441 ( .A(p_input[4277]), .B(n29676), .Z(n29679) );
  XNOR U29442 ( .A(n29676), .B(n29323), .Z(n29678) );
  IV U29443 ( .A(p_input[4245]), .Z(n29323) );
  XOR U29444 ( .A(n29680), .B(n29681), .Z(n29676) );
  AND U29445 ( .A(n29682), .B(n29683), .Z(n29681) );
  XNOR U29446 ( .A(p_input[4276]), .B(n29680), .Z(n29683) );
  XNOR U29447 ( .A(n29680), .B(n29332), .Z(n29682) );
  IV U29448 ( .A(p_input[4244]), .Z(n29332) );
  XOR U29449 ( .A(n29684), .B(n29685), .Z(n29680) );
  AND U29450 ( .A(n29686), .B(n29687), .Z(n29685) );
  XNOR U29451 ( .A(p_input[4275]), .B(n29684), .Z(n29687) );
  XNOR U29452 ( .A(n29684), .B(n29341), .Z(n29686) );
  IV U29453 ( .A(p_input[4243]), .Z(n29341) );
  XOR U29454 ( .A(n29688), .B(n29689), .Z(n29684) );
  AND U29455 ( .A(n29690), .B(n29691), .Z(n29689) );
  XNOR U29456 ( .A(p_input[4274]), .B(n29688), .Z(n29691) );
  XNOR U29457 ( .A(n29688), .B(n29350), .Z(n29690) );
  IV U29458 ( .A(p_input[4242]), .Z(n29350) );
  XOR U29459 ( .A(n29692), .B(n29693), .Z(n29688) );
  AND U29460 ( .A(n29694), .B(n29695), .Z(n29693) );
  XNOR U29461 ( .A(p_input[4273]), .B(n29692), .Z(n29695) );
  XNOR U29462 ( .A(n29692), .B(n29359), .Z(n29694) );
  IV U29463 ( .A(p_input[4241]), .Z(n29359) );
  XOR U29464 ( .A(n29696), .B(n29697), .Z(n29692) );
  AND U29465 ( .A(n29698), .B(n29699), .Z(n29697) );
  XNOR U29466 ( .A(p_input[4272]), .B(n29696), .Z(n29699) );
  XNOR U29467 ( .A(n29696), .B(n29368), .Z(n29698) );
  IV U29468 ( .A(p_input[4240]), .Z(n29368) );
  XOR U29469 ( .A(n29700), .B(n29701), .Z(n29696) );
  AND U29470 ( .A(n29702), .B(n29703), .Z(n29701) );
  XNOR U29471 ( .A(p_input[4271]), .B(n29700), .Z(n29703) );
  XNOR U29472 ( .A(n29700), .B(n29377), .Z(n29702) );
  IV U29473 ( .A(p_input[4239]), .Z(n29377) );
  XOR U29474 ( .A(n29704), .B(n29705), .Z(n29700) );
  AND U29475 ( .A(n29706), .B(n29707), .Z(n29705) );
  XNOR U29476 ( .A(p_input[4270]), .B(n29704), .Z(n29707) );
  XNOR U29477 ( .A(n29704), .B(n29386), .Z(n29706) );
  IV U29478 ( .A(p_input[4238]), .Z(n29386) );
  XOR U29479 ( .A(n29708), .B(n29709), .Z(n29704) );
  AND U29480 ( .A(n29710), .B(n29711), .Z(n29709) );
  XNOR U29481 ( .A(p_input[4269]), .B(n29708), .Z(n29711) );
  XNOR U29482 ( .A(n29708), .B(n29395), .Z(n29710) );
  IV U29483 ( .A(p_input[4237]), .Z(n29395) );
  XOR U29484 ( .A(n29712), .B(n29713), .Z(n29708) );
  AND U29485 ( .A(n29714), .B(n29715), .Z(n29713) );
  XNOR U29486 ( .A(p_input[4268]), .B(n29712), .Z(n29715) );
  XNOR U29487 ( .A(n29712), .B(n29404), .Z(n29714) );
  IV U29488 ( .A(p_input[4236]), .Z(n29404) );
  XOR U29489 ( .A(n29716), .B(n29717), .Z(n29712) );
  AND U29490 ( .A(n29718), .B(n29719), .Z(n29717) );
  XNOR U29491 ( .A(p_input[4267]), .B(n29716), .Z(n29719) );
  XNOR U29492 ( .A(n29716), .B(n29413), .Z(n29718) );
  IV U29493 ( .A(p_input[4235]), .Z(n29413) );
  XOR U29494 ( .A(n29720), .B(n29721), .Z(n29716) );
  AND U29495 ( .A(n29722), .B(n29723), .Z(n29721) );
  XNOR U29496 ( .A(p_input[4266]), .B(n29720), .Z(n29723) );
  XNOR U29497 ( .A(n29720), .B(n29422), .Z(n29722) );
  IV U29498 ( .A(p_input[4234]), .Z(n29422) );
  XOR U29499 ( .A(n29724), .B(n29725), .Z(n29720) );
  AND U29500 ( .A(n29726), .B(n29727), .Z(n29725) );
  XNOR U29501 ( .A(p_input[4265]), .B(n29724), .Z(n29727) );
  XNOR U29502 ( .A(n29724), .B(n29431), .Z(n29726) );
  IV U29503 ( .A(p_input[4233]), .Z(n29431) );
  XOR U29504 ( .A(n29728), .B(n29729), .Z(n29724) );
  AND U29505 ( .A(n29730), .B(n29731), .Z(n29729) );
  XNOR U29506 ( .A(p_input[4264]), .B(n29728), .Z(n29731) );
  XNOR U29507 ( .A(n29728), .B(n29440), .Z(n29730) );
  IV U29508 ( .A(p_input[4232]), .Z(n29440) );
  XOR U29509 ( .A(n29732), .B(n29733), .Z(n29728) );
  AND U29510 ( .A(n29734), .B(n29735), .Z(n29733) );
  XNOR U29511 ( .A(p_input[4263]), .B(n29732), .Z(n29735) );
  XNOR U29512 ( .A(n29732), .B(n29449), .Z(n29734) );
  IV U29513 ( .A(p_input[4231]), .Z(n29449) );
  XOR U29514 ( .A(n29736), .B(n29737), .Z(n29732) );
  AND U29515 ( .A(n29738), .B(n29739), .Z(n29737) );
  XNOR U29516 ( .A(p_input[4262]), .B(n29736), .Z(n29739) );
  XNOR U29517 ( .A(n29736), .B(n29458), .Z(n29738) );
  IV U29518 ( .A(p_input[4230]), .Z(n29458) );
  XOR U29519 ( .A(n29740), .B(n29741), .Z(n29736) );
  AND U29520 ( .A(n29742), .B(n29743), .Z(n29741) );
  XNOR U29521 ( .A(p_input[4261]), .B(n29740), .Z(n29743) );
  XNOR U29522 ( .A(n29740), .B(n29467), .Z(n29742) );
  IV U29523 ( .A(p_input[4229]), .Z(n29467) );
  XOR U29524 ( .A(n29744), .B(n29745), .Z(n29740) );
  AND U29525 ( .A(n29746), .B(n29747), .Z(n29745) );
  XNOR U29526 ( .A(p_input[4260]), .B(n29744), .Z(n29747) );
  XNOR U29527 ( .A(n29744), .B(n29476), .Z(n29746) );
  IV U29528 ( .A(p_input[4228]), .Z(n29476) );
  XOR U29529 ( .A(n29748), .B(n29749), .Z(n29744) );
  AND U29530 ( .A(n29750), .B(n29751), .Z(n29749) );
  XNOR U29531 ( .A(p_input[4259]), .B(n29748), .Z(n29751) );
  XNOR U29532 ( .A(n29748), .B(n29485), .Z(n29750) );
  IV U29533 ( .A(p_input[4227]), .Z(n29485) );
  XOR U29534 ( .A(n29752), .B(n29753), .Z(n29748) );
  AND U29535 ( .A(n29754), .B(n29755), .Z(n29753) );
  XNOR U29536 ( .A(p_input[4258]), .B(n29752), .Z(n29755) );
  XNOR U29537 ( .A(n29752), .B(n29494), .Z(n29754) );
  IV U29538 ( .A(p_input[4226]), .Z(n29494) );
  XNOR U29539 ( .A(n29756), .B(n29757), .Z(n29752) );
  AND U29540 ( .A(n29758), .B(n29759), .Z(n29757) );
  XOR U29541 ( .A(p_input[4257]), .B(n29756), .Z(n29759) );
  XNOR U29542 ( .A(p_input[4225]), .B(n29756), .Z(n29758) );
  AND U29543 ( .A(p_input[4256]), .B(n29760), .Z(n29756) );
  IV U29544 ( .A(p_input[4224]), .Z(n29760) );
  XOR U29545 ( .A(n29761), .B(n29762), .Z(n28850) );
  AND U29546 ( .A(n540), .B(n29763), .Z(n29762) );
  XNOR U29547 ( .A(n29764), .B(n29761), .Z(n29763) );
  XOR U29548 ( .A(n29765), .B(n29766), .Z(n540) );
  AND U29549 ( .A(n29767), .B(n29768), .Z(n29766) );
  XNOR U29550 ( .A(n28865), .B(n29765), .Z(n29768) );
  AND U29551 ( .A(p_input[4223]), .B(p_input[4191]), .Z(n28865) );
  XNOR U29552 ( .A(n29765), .B(n28862), .Z(n29767) );
  IV U29553 ( .A(n29769), .Z(n28862) );
  AND U29554 ( .A(p_input[4127]), .B(p_input[4159]), .Z(n29769) );
  XOR U29555 ( .A(n29770), .B(n29771), .Z(n29765) );
  AND U29556 ( .A(n29772), .B(n29773), .Z(n29771) );
  XOR U29557 ( .A(n29770), .B(n28877), .Z(n29773) );
  XNOR U29558 ( .A(p_input[4190]), .B(n29774), .Z(n28877) );
  AND U29559 ( .A(n415), .B(n29775), .Z(n29774) );
  XOR U29560 ( .A(p_input[4222]), .B(p_input[4190]), .Z(n29775) );
  XNOR U29561 ( .A(n28874), .B(n29770), .Z(n29772) );
  XOR U29562 ( .A(n29776), .B(n29777), .Z(n28874) );
  AND U29563 ( .A(n412), .B(n29778), .Z(n29777) );
  XOR U29564 ( .A(p_input[4158]), .B(p_input[4126]), .Z(n29778) );
  XOR U29565 ( .A(n29779), .B(n29780), .Z(n29770) );
  AND U29566 ( .A(n29781), .B(n29782), .Z(n29780) );
  XOR U29567 ( .A(n29779), .B(n28889), .Z(n29782) );
  XNOR U29568 ( .A(p_input[4189]), .B(n29783), .Z(n28889) );
  AND U29569 ( .A(n415), .B(n29784), .Z(n29783) );
  XOR U29570 ( .A(p_input[4221]), .B(p_input[4189]), .Z(n29784) );
  XNOR U29571 ( .A(n28886), .B(n29779), .Z(n29781) );
  XOR U29572 ( .A(n29785), .B(n29786), .Z(n28886) );
  AND U29573 ( .A(n412), .B(n29787), .Z(n29786) );
  XOR U29574 ( .A(p_input[4157]), .B(p_input[4125]), .Z(n29787) );
  XOR U29575 ( .A(n29788), .B(n29789), .Z(n29779) );
  AND U29576 ( .A(n29790), .B(n29791), .Z(n29789) );
  XOR U29577 ( .A(n29788), .B(n28901), .Z(n29791) );
  XNOR U29578 ( .A(p_input[4188]), .B(n29792), .Z(n28901) );
  AND U29579 ( .A(n415), .B(n29793), .Z(n29792) );
  XOR U29580 ( .A(p_input[4220]), .B(p_input[4188]), .Z(n29793) );
  XNOR U29581 ( .A(n28898), .B(n29788), .Z(n29790) );
  XOR U29582 ( .A(n29794), .B(n29795), .Z(n28898) );
  AND U29583 ( .A(n412), .B(n29796), .Z(n29795) );
  XOR U29584 ( .A(p_input[4156]), .B(p_input[4124]), .Z(n29796) );
  XOR U29585 ( .A(n29797), .B(n29798), .Z(n29788) );
  AND U29586 ( .A(n29799), .B(n29800), .Z(n29798) );
  XOR U29587 ( .A(n29797), .B(n28913), .Z(n29800) );
  XNOR U29588 ( .A(p_input[4187]), .B(n29801), .Z(n28913) );
  AND U29589 ( .A(n415), .B(n29802), .Z(n29801) );
  XOR U29590 ( .A(p_input[4219]), .B(p_input[4187]), .Z(n29802) );
  XNOR U29591 ( .A(n28910), .B(n29797), .Z(n29799) );
  XOR U29592 ( .A(n29803), .B(n29804), .Z(n28910) );
  AND U29593 ( .A(n412), .B(n29805), .Z(n29804) );
  XOR U29594 ( .A(p_input[4155]), .B(p_input[4123]), .Z(n29805) );
  XOR U29595 ( .A(n29806), .B(n29807), .Z(n29797) );
  AND U29596 ( .A(n29808), .B(n29809), .Z(n29807) );
  XOR U29597 ( .A(n29806), .B(n28925), .Z(n29809) );
  XNOR U29598 ( .A(p_input[4186]), .B(n29810), .Z(n28925) );
  AND U29599 ( .A(n415), .B(n29811), .Z(n29810) );
  XOR U29600 ( .A(p_input[4218]), .B(p_input[4186]), .Z(n29811) );
  XNOR U29601 ( .A(n28922), .B(n29806), .Z(n29808) );
  XOR U29602 ( .A(n29812), .B(n29813), .Z(n28922) );
  AND U29603 ( .A(n412), .B(n29814), .Z(n29813) );
  XOR U29604 ( .A(p_input[4154]), .B(p_input[4122]), .Z(n29814) );
  XOR U29605 ( .A(n29815), .B(n29816), .Z(n29806) );
  AND U29606 ( .A(n29817), .B(n29818), .Z(n29816) );
  XOR U29607 ( .A(n29815), .B(n28937), .Z(n29818) );
  XNOR U29608 ( .A(p_input[4185]), .B(n29819), .Z(n28937) );
  AND U29609 ( .A(n415), .B(n29820), .Z(n29819) );
  XOR U29610 ( .A(p_input[4217]), .B(p_input[4185]), .Z(n29820) );
  XNOR U29611 ( .A(n28934), .B(n29815), .Z(n29817) );
  XOR U29612 ( .A(n29821), .B(n29822), .Z(n28934) );
  AND U29613 ( .A(n412), .B(n29823), .Z(n29822) );
  XOR U29614 ( .A(p_input[4153]), .B(p_input[4121]), .Z(n29823) );
  XOR U29615 ( .A(n29824), .B(n29825), .Z(n29815) );
  AND U29616 ( .A(n29826), .B(n29827), .Z(n29825) );
  XOR U29617 ( .A(n29824), .B(n28949), .Z(n29827) );
  XNOR U29618 ( .A(p_input[4184]), .B(n29828), .Z(n28949) );
  AND U29619 ( .A(n415), .B(n29829), .Z(n29828) );
  XOR U29620 ( .A(p_input[4216]), .B(p_input[4184]), .Z(n29829) );
  XNOR U29621 ( .A(n28946), .B(n29824), .Z(n29826) );
  XOR U29622 ( .A(n29830), .B(n29831), .Z(n28946) );
  AND U29623 ( .A(n412), .B(n29832), .Z(n29831) );
  XOR U29624 ( .A(p_input[4152]), .B(p_input[4120]), .Z(n29832) );
  XOR U29625 ( .A(n29833), .B(n29834), .Z(n29824) );
  AND U29626 ( .A(n29835), .B(n29836), .Z(n29834) );
  XOR U29627 ( .A(n29833), .B(n28961), .Z(n29836) );
  XNOR U29628 ( .A(p_input[4183]), .B(n29837), .Z(n28961) );
  AND U29629 ( .A(n415), .B(n29838), .Z(n29837) );
  XOR U29630 ( .A(p_input[4215]), .B(p_input[4183]), .Z(n29838) );
  XNOR U29631 ( .A(n28958), .B(n29833), .Z(n29835) );
  XOR U29632 ( .A(n29839), .B(n29840), .Z(n28958) );
  AND U29633 ( .A(n412), .B(n29841), .Z(n29840) );
  XOR U29634 ( .A(p_input[4151]), .B(p_input[4119]), .Z(n29841) );
  XOR U29635 ( .A(n29842), .B(n29843), .Z(n29833) );
  AND U29636 ( .A(n29844), .B(n29845), .Z(n29843) );
  XOR U29637 ( .A(n29842), .B(n28973), .Z(n29845) );
  XNOR U29638 ( .A(p_input[4182]), .B(n29846), .Z(n28973) );
  AND U29639 ( .A(n415), .B(n29847), .Z(n29846) );
  XOR U29640 ( .A(p_input[4214]), .B(p_input[4182]), .Z(n29847) );
  XNOR U29641 ( .A(n28970), .B(n29842), .Z(n29844) );
  XOR U29642 ( .A(n29848), .B(n29849), .Z(n28970) );
  AND U29643 ( .A(n412), .B(n29850), .Z(n29849) );
  XOR U29644 ( .A(p_input[4150]), .B(p_input[4118]), .Z(n29850) );
  XOR U29645 ( .A(n29851), .B(n29852), .Z(n29842) );
  AND U29646 ( .A(n29853), .B(n29854), .Z(n29852) );
  XOR U29647 ( .A(n29851), .B(n28985), .Z(n29854) );
  XNOR U29648 ( .A(p_input[4181]), .B(n29855), .Z(n28985) );
  AND U29649 ( .A(n415), .B(n29856), .Z(n29855) );
  XOR U29650 ( .A(p_input[4213]), .B(p_input[4181]), .Z(n29856) );
  XNOR U29651 ( .A(n28982), .B(n29851), .Z(n29853) );
  XOR U29652 ( .A(n29857), .B(n29858), .Z(n28982) );
  AND U29653 ( .A(n412), .B(n29859), .Z(n29858) );
  XOR U29654 ( .A(p_input[4149]), .B(p_input[4117]), .Z(n29859) );
  XOR U29655 ( .A(n29860), .B(n29861), .Z(n29851) );
  AND U29656 ( .A(n29862), .B(n29863), .Z(n29861) );
  XOR U29657 ( .A(n29860), .B(n28997), .Z(n29863) );
  XNOR U29658 ( .A(p_input[4180]), .B(n29864), .Z(n28997) );
  AND U29659 ( .A(n415), .B(n29865), .Z(n29864) );
  XOR U29660 ( .A(p_input[4212]), .B(p_input[4180]), .Z(n29865) );
  XNOR U29661 ( .A(n28994), .B(n29860), .Z(n29862) );
  XOR U29662 ( .A(n29866), .B(n29867), .Z(n28994) );
  AND U29663 ( .A(n412), .B(n29868), .Z(n29867) );
  XOR U29664 ( .A(p_input[4148]), .B(p_input[4116]), .Z(n29868) );
  XOR U29665 ( .A(n29869), .B(n29870), .Z(n29860) );
  AND U29666 ( .A(n29871), .B(n29872), .Z(n29870) );
  XOR U29667 ( .A(n29869), .B(n29009), .Z(n29872) );
  XNOR U29668 ( .A(p_input[4179]), .B(n29873), .Z(n29009) );
  AND U29669 ( .A(n415), .B(n29874), .Z(n29873) );
  XOR U29670 ( .A(p_input[4211]), .B(p_input[4179]), .Z(n29874) );
  XNOR U29671 ( .A(n29006), .B(n29869), .Z(n29871) );
  XOR U29672 ( .A(n29875), .B(n29876), .Z(n29006) );
  AND U29673 ( .A(n412), .B(n29877), .Z(n29876) );
  XOR U29674 ( .A(p_input[4147]), .B(p_input[4115]), .Z(n29877) );
  XOR U29675 ( .A(n29878), .B(n29879), .Z(n29869) );
  AND U29676 ( .A(n29880), .B(n29881), .Z(n29879) );
  XOR U29677 ( .A(n29878), .B(n29021), .Z(n29881) );
  XNOR U29678 ( .A(p_input[4178]), .B(n29882), .Z(n29021) );
  AND U29679 ( .A(n415), .B(n29883), .Z(n29882) );
  XOR U29680 ( .A(p_input[4210]), .B(p_input[4178]), .Z(n29883) );
  XNOR U29681 ( .A(n29018), .B(n29878), .Z(n29880) );
  XOR U29682 ( .A(n29884), .B(n29885), .Z(n29018) );
  AND U29683 ( .A(n412), .B(n29886), .Z(n29885) );
  XOR U29684 ( .A(p_input[4146]), .B(p_input[4114]), .Z(n29886) );
  XOR U29685 ( .A(n29887), .B(n29888), .Z(n29878) );
  AND U29686 ( .A(n29889), .B(n29890), .Z(n29888) );
  XOR U29687 ( .A(n29887), .B(n29033), .Z(n29890) );
  XNOR U29688 ( .A(p_input[4177]), .B(n29891), .Z(n29033) );
  AND U29689 ( .A(n415), .B(n29892), .Z(n29891) );
  XOR U29690 ( .A(p_input[4209]), .B(p_input[4177]), .Z(n29892) );
  XNOR U29691 ( .A(n29030), .B(n29887), .Z(n29889) );
  XOR U29692 ( .A(n29893), .B(n29894), .Z(n29030) );
  AND U29693 ( .A(n412), .B(n29895), .Z(n29894) );
  XOR U29694 ( .A(p_input[4145]), .B(p_input[4113]), .Z(n29895) );
  XOR U29695 ( .A(n29896), .B(n29897), .Z(n29887) );
  AND U29696 ( .A(n29898), .B(n29899), .Z(n29897) );
  XOR U29697 ( .A(n29896), .B(n29045), .Z(n29899) );
  XNOR U29698 ( .A(p_input[4176]), .B(n29900), .Z(n29045) );
  AND U29699 ( .A(n415), .B(n29901), .Z(n29900) );
  XOR U29700 ( .A(p_input[4208]), .B(p_input[4176]), .Z(n29901) );
  XNOR U29701 ( .A(n29042), .B(n29896), .Z(n29898) );
  XOR U29702 ( .A(n29902), .B(n29903), .Z(n29042) );
  AND U29703 ( .A(n412), .B(n29904), .Z(n29903) );
  XOR U29704 ( .A(p_input[4144]), .B(p_input[4112]), .Z(n29904) );
  XOR U29705 ( .A(n29905), .B(n29906), .Z(n29896) );
  AND U29706 ( .A(n29907), .B(n29908), .Z(n29906) );
  XOR U29707 ( .A(n29905), .B(n29057), .Z(n29908) );
  XNOR U29708 ( .A(p_input[4175]), .B(n29909), .Z(n29057) );
  AND U29709 ( .A(n415), .B(n29910), .Z(n29909) );
  XOR U29710 ( .A(p_input[4207]), .B(p_input[4175]), .Z(n29910) );
  XNOR U29711 ( .A(n29054), .B(n29905), .Z(n29907) );
  XOR U29712 ( .A(n29911), .B(n29912), .Z(n29054) );
  AND U29713 ( .A(n412), .B(n29913), .Z(n29912) );
  XOR U29714 ( .A(p_input[4143]), .B(p_input[4111]), .Z(n29913) );
  XOR U29715 ( .A(n29914), .B(n29915), .Z(n29905) );
  AND U29716 ( .A(n29916), .B(n29917), .Z(n29915) );
  XOR U29717 ( .A(n29914), .B(n29069), .Z(n29917) );
  XNOR U29718 ( .A(p_input[4174]), .B(n29918), .Z(n29069) );
  AND U29719 ( .A(n415), .B(n29919), .Z(n29918) );
  XOR U29720 ( .A(p_input[4206]), .B(p_input[4174]), .Z(n29919) );
  XNOR U29721 ( .A(n29066), .B(n29914), .Z(n29916) );
  XOR U29722 ( .A(n29920), .B(n29921), .Z(n29066) );
  AND U29723 ( .A(n412), .B(n29922), .Z(n29921) );
  XOR U29724 ( .A(p_input[4142]), .B(p_input[4110]), .Z(n29922) );
  XOR U29725 ( .A(n29923), .B(n29924), .Z(n29914) );
  AND U29726 ( .A(n29925), .B(n29926), .Z(n29924) );
  XOR U29727 ( .A(n29923), .B(n29081), .Z(n29926) );
  XNOR U29728 ( .A(p_input[4173]), .B(n29927), .Z(n29081) );
  AND U29729 ( .A(n415), .B(n29928), .Z(n29927) );
  XOR U29730 ( .A(p_input[4205]), .B(p_input[4173]), .Z(n29928) );
  XNOR U29731 ( .A(n29078), .B(n29923), .Z(n29925) );
  XOR U29732 ( .A(n29929), .B(n29930), .Z(n29078) );
  AND U29733 ( .A(n412), .B(n29931), .Z(n29930) );
  XOR U29734 ( .A(p_input[4141]), .B(p_input[4109]), .Z(n29931) );
  XOR U29735 ( .A(n29932), .B(n29933), .Z(n29923) );
  AND U29736 ( .A(n29934), .B(n29935), .Z(n29933) );
  XOR U29737 ( .A(n29932), .B(n29093), .Z(n29935) );
  XNOR U29738 ( .A(p_input[4172]), .B(n29936), .Z(n29093) );
  AND U29739 ( .A(n415), .B(n29937), .Z(n29936) );
  XOR U29740 ( .A(p_input[4204]), .B(p_input[4172]), .Z(n29937) );
  XNOR U29741 ( .A(n29090), .B(n29932), .Z(n29934) );
  XOR U29742 ( .A(n29938), .B(n29939), .Z(n29090) );
  AND U29743 ( .A(n412), .B(n29940), .Z(n29939) );
  XOR U29744 ( .A(p_input[4140]), .B(p_input[4108]), .Z(n29940) );
  XOR U29745 ( .A(n29941), .B(n29942), .Z(n29932) );
  AND U29746 ( .A(n29943), .B(n29944), .Z(n29942) );
  XOR U29747 ( .A(n29941), .B(n29105), .Z(n29944) );
  XNOR U29748 ( .A(p_input[4171]), .B(n29945), .Z(n29105) );
  AND U29749 ( .A(n415), .B(n29946), .Z(n29945) );
  XOR U29750 ( .A(p_input[4203]), .B(p_input[4171]), .Z(n29946) );
  XNOR U29751 ( .A(n29102), .B(n29941), .Z(n29943) );
  XOR U29752 ( .A(n29947), .B(n29948), .Z(n29102) );
  AND U29753 ( .A(n412), .B(n29949), .Z(n29948) );
  XOR U29754 ( .A(p_input[4139]), .B(p_input[4107]), .Z(n29949) );
  XOR U29755 ( .A(n29950), .B(n29951), .Z(n29941) );
  AND U29756 ( .A(n29952), .B(n29953), .Z(n29951) );
  XOR U29757 ( .A(n29950), .B(n29117), .Z(n29953) );
  XNOR U29758 ( .A(p_input[4170]), .B(n29954), .Z(n29117) );
  AND U29759 ( .A(n415), .B(n29955), .Z(n29954) );
  XOR U29760 ( .A(p_input[4202]), .B(p_input[4170]), .Z(n29955) );
  XNOR U29761 ( .A(n29114), .B(n29950), .Z(n29952) );
  XOR U29762 ( .A(n29956), .B(n29957), .Z(n29114) );
  AND U29763 ( .A(n412), .B(n29958), .Z(n29957) );
  XOR U29764 ( .A(p_input[4138]), .B(p_input[4106]), .Z(n29958) );
  XOR U29765 ( .A(n29959), .B(n29960), .Z(n29950) );
  AND U29766 ( .A(n29961), .B(n29962), .Z(n29960) );
  XOR U29767 ( .A(n29959), .B(n29129), .Z(n29962) );
  XNOR U29768 ( .A(p_input[4169]), .B(n29963), .Z(n29129) );
  AND U29769 ( .A(n415), .B(n29964), .Z(n29963) );
  XOR U29770 ( .A(p_input[4201]), .B(p_input[4169]), .Z(n29964) );
  XNOR U29771 ( .A(n29126), .B(n29959), .Z(n29961) );
  XOR U29772 ( .A(n29965), .B(n29966), .Z(n29126) );
  AND U29773 ( .A(n412), .B(n29967), .Z(n29966) );
  XOR U29774 ( .A(p_input[4137]), .B(p_input[4105]), .Z(n29967) );
  XOR U29775 ( .A(n29968), .B(n29969), .Z(n29959) );
  AND U29776 ( .A(n29970), .B(n29971), .Z(n29969) );
  XOR U29777 ( .A(n29968), .B(n29141), .Z(n29971) );
  XNOR U29778 ( .A(p_input[4168]), .B(n29972), .Z(n29141) );
  AND U29779 ( .A(n415), .B(n29973), .Z(n29972) );
  XOR U29780 ( .A(p_input[4200]), .B(p_input[4168]), .Z(n29973) );
  XNOR U29781 ( .A(n29138), .B(n29968), .Z(n29970) );
  XOR U29782 ( .A(n29974), .B(n29975), .Z(n29138) );
  AND U29783 ( .A(n412), .B(n29976), .Z(n29975) );
  XOR U29784 ( .A(p_input[4136]), .B(p_input[4104]), .Z(n29976) );
  XOR U29785 ( .A(n29977), .B(n29978), .Z(n29968) );
  AND U29786 ( .A(n29979), .B(n29980), .Z(n29978) );
  XOR U29787 ( .A(n29977), .B(n29153), .Z(n29980) );
  XNOR U29788 ( .A(p_input[4167]), .B(n29981), .Z(n29153) );
  AND U29789 ( .A(n415), .B(n29982), .Z(n29981) );
  XOR U29790 ( .A(p_input[4199]), .B(p_input[4167]), .Z(n29982) );
  XNOR U29791 ( .A(n29150), .B(n29977), .Z(n29979) );
  XOR U29792 ( .A(n29983), .B(n29984), .Z(n29150) );
  AND U29793 ( .A(n412), .B(n29985), .Z(n29984) );
  XOR U29794 ( .A(p_input[4135]), .B(p_input[4103]), .Z(n29985) );
  XOR U29795 ( .A(n29986), .B(n29987), .Z(n29977) );
  AND U29796 ( .A(n29988), .B(n29989), .Z(n29987) );
  XOR U29797 ( .A(n29986), .B(n29165), .Z(n29989) );
  XNOR U29798 ( .A(p_input[4166]), .B(n29990), .Z(n29165) );
  AND U29799 ( .A(n415), .B(n29991), .Z(n29990) );
  XOR U29800 ( .A(p_input[4198]), .B(p_input[4166]), .Z(n29991) );
  XNOR U29801 ( .A(n29162), .B(n29986), .Z(n29988) );
  XOR U29802 ( .A(n29992), .B(n29993), .Z(n29162) );
  AND U29803 ( .A(n412), .B(n29994), .Z(n29993) );
  XOR U29804 ( .A(p_input[4134]), .B(p_input[4102]), .Z(n29994) );
  XOR U29805 ( .A(n29995), .B(n29996), .Z(n29986) );
  AND U29806 ( .A(n29997), .B(n29998), .Z(n29996) );
  XOR U29807 ( .A(n29995), .B(n29177), .Z(n29998) );
  XNOR U29808 ( .A(p_input[4165]), .B(n29999), .Z(n29177) );
  AND U29809 ( .A(n415), .B(n30000), .Z(n29999) );
  XOR U29810 ( .A(p_input[4197]), .B(p_input[4165]), .Z(n30000) );
  XNOR U29811 ( .A(n29174), .B(n29995), .Z(n29997) );
  XOR U29812 ( .A(n30001), .B(n30002), .Z(n29174) );
  AND U29813 ( .A(n412), .B(n30003), .Z(n30002) );
  XOR U29814 ( .A(p_input[4133]), .B(p_input[4101]), .Z(n30003) );
  XOR U29815 ( .A(n30004), .B(n30005), .Z(n29995) );
  AND U29816 ( .A(n30006), .B(n30007), .Z(n30005) );
  XOR U29817 ( .A(n30004), .B(n29189), .Z(n30007) );
  XNOR U29818 ( .A(p_input[4164]), .B(n30008), .Z(n29189) );
  AND U29819 ( .A(n415), .B(n30009), .Z(n30008) );
  XOR U29820 ( .A(p_input[4196]), .B(p_input[4164]), .Z(n30009) );
  XNOR U29821 ( .A(n29186), .B(n30004), .Z(n30006) );
  XOR U29822 ( .A(n30010), .B(n30011), .Z(n29186) );
  AND U29823 ( .A(n412), .B(n30012), .Z(n30011) );
  XOR U29824 ( .A(p_input[4132]), .B(p_input[4100]), .Z(n30012) );
  XOR U29825 ( .A(n30013), .B(n30014), .Z(n30004) );
  AND U29826 ( .A(n30015), .B(n30016), .Z(n30014) );
  XOR U29827 ( .A(n30013), .B(n29201), .Z(n30016) );
  XNOR U29828 ( .A(p_input[4163]), .B(n30017), .Z(n29201) );
  AND U29829 ( .A(n415), .B(n30018), .Z(n30017) );
  XOR U29830 ( .A(p_input[4195]), .B(p_input[4163]), .Z(n30018) );
  XNOR U29831 ( .A(n29198), .B(n30013), .Z(n30015) );
  XOR U29832 ( .A(n30019), .B(n30020), .Z(n29198) );
  AND U29833 ( .A(n412), .B(n30021), .Z(n30020) );
  XOR U29834 ( .A(p_input[4131]), .B(p_input[4099]), .Z(n30021) );
  XOR U29835 ( .A(n30022), .B(n30023), .Z(n30013) );
  AND U29836 ( .A(n30024), .B(n30025), .Z(n30023) );
  XOR U29837 ( .A(n30022), .B(n29213), .Z(n30025) );
  XNOR U29838 ( .A(p_input[4162]), .B(n30026), .Z(n29213) );
  AND U29839 ( .A(n415), .B(n30027), .Z(n30026) );
  XOR U29840 ( .A(p_input[4194]), .B(p_input[4162]), .Z(n30027) );
  XNOR U29841 ( .A(n29210), .B(n30022), .Z(n30024) );
  XOR U29842 ( .A(n30028), .B(n30029), .Z(n29210) );
  AND U29843 ( .A(n412), .B(n30030), .Z(n30029) );
  XOR U29844 ( .A(p_input[4130]), .B(p_input[4098]), .Z(n30030) );
  XOR U29845 ( .A(n30031), .B(n30032), .Z(n30022) );
  AND U29846 ( .A(n30033), .B(n30034), .Z(n30032) );
  XNOR U29847 ( .A(n30035), .B(n29226), .Z(n30034) );
  XNOR U29848 ( .A(p_input[4161]), .B(n30036), .Z(n29226) );
  AND U29849 ( .A(n415), .B(n30037), .Z(n30036) );
  XNOR U29850 ( .A(p_input[4193]), .B(n30038), .Z(n30037) );
  IV U29851 ( .A(p_input[4161]), .Z(n30038) );
  XNOR U29852 ( .A(n29223), .B(n30031), .Z(n30033) );
  XNOR U29853 ( .A(p_input[4097]), .B(n30039), .Z(n29223) );
  AND U29854 ( .A(n412), .B(n30040), .Z(n30039) );
  XOR U29855 ( .A(p_input[4129]), .B(p_input[4097]), .Z(n30040) );
  IV U29856 ( .A(n30035), .Z(n30031) );
  AND U29857 ( .A(n29761), .B(n29764), .Z(n30035) );
  XOR U29858 ( .A(p_input[4160]), .B(n30041), .Z(n29764) );
  AND U29859 ( .A(n415), .B(n30042), .Z(n30041) );
  XOR U29860 ( .A(p_input[4192]), .B(p_input[4160]), .Z(n30042) );
  XOR U29861 ( .A(n30043), .B(n30044), .Z(n415) );
  AND U29862 ( .A(n30045), .B(n30046), .Z(n30044) );
  XNOR U29863 ( .A(p_input[4223]), .B(n30043), .Z(n30046) );
  XOR U29864 ( .A(n30043), .B(p_input[4191]), .Z(n30045) );
  XOR U29865 ( .A(n30047), .B(n30048), .Z(n30043) );
  AND U29866 ( .A(n30049), .B(n30050), .Z(n30048) );
  XNOR U29867 ( .A(p_input[4222]), .B(n30047), .Z(n30050) );
  XOR U29868 ( .A(n30047), .B(p_input[4190]), .Z(n30049) );
  XOR U29869 ( .A(n30051), .B(n30052), .Z(n30047) );
  AND U29870 ( .A(n30053), .B(n30054), .Z(n30052) );
  XNOR U29871 ( .A(p_input[4221]), .B(n30051), .Z(n30054) );
  XOR U29872 ( .A(n30051), .B(p_input[4189]), .Z(n30053) );
  XOR U29873 ( .A(n30055), .B(n30056), .Z(n30051) );
  AND U29874 ( .A(n30057), .B(n30058), .Z(n30056) );
  XNOR U29875 ( .A(p_input[4220]), .B(n30055), .Z(n30058) );
  XOR U29876 ( .A(n30055), .B(p_input[4188]), .Z(n30057) );
  XOR U29877 ( .A(n30059), .B(n30060), .Z(n30055) );
  AND U29878 ( .A(n30061), .B(n30062), .Z(n30060) );
  XNOR U29879 ( .A(p_input[4219]), .B(n30059), .Z(n30062) );
  XOR U29880 ( .A(n30059), .B(p_input[4187]), .Z(n30061) );
  XOR U29881 ( .A(n30063), .B(n30064), .Z(n30059) );
  AND U29882 ( .A(n30065), .B(n30066), .Z(n30064) );
  XNOR U29883 ( .A(p_input[4218]), .B(n30063), .Z(n30066) );
  XOR U29884 ( .A(n30063), .B(p_input[4186]), .Z(n30065) );
  XOR U29885 ( .A(n30067), .B(n30068), .Z(n30063) );
  AND U29886 ( .A(n30069), .B(n30070), .Z(n30068) );
  XNOR U29887 ( .A(p_input[4217]), .B(n30067), .Z(n30070) );
  XOR U29888 ( .A(n30067), .B(p_input[4185]), .Z(n30069) );
  XOR U29889 ( .A(n30071), .B(n30072), .Z(n30067) );
  AND U29890 ( .A(n30073), .B(n30074), .Z(n30072) );
  XNOR U29891 ( .A(p_input[4216]), .B(n30071), .Z(n30074) );
  XOR U29892 ( .A(n30071), .B(p_input[4184]), .Z(n30073) );
  XOR U29893 ( .A(n30075), .B(n30076), .Z(n30071) );
  AND U29894 ( .A(n30077), .B(n30078), .Z(n30076) );
  XNOR U29895 ( .A(p_input[4215]), .B(n30075), .Z(n30078) );
  XOR U29896 ( .A(n30075), .B(p_input[4183]), .Z(n30077) );
  XOR U29897 ( .A(n30079), .B(n30080), .Z(n30075) );
  AND U29898 ( .A(n30081), .B(n30082), .Z(n30080) );
  XNOR U29899 ( .A(p_input[4214]), .B(n30079), .Z(n30082) );
  XOR U29900 ( .A(n30079), .B(p_input[4182]), .Z(n30081) );
  XOR U29901 ( .A(n30083), .B(n30084), .Z(n30079) );
  AND U29902 ( .A(n30085), .B(n30086), .Z(n30084) );
  XNOR U29903 ( .A(p_input[4213]), .B(n30083), .Z(n30086) );
  XOR U29904 ( .A(n30083), .B(p_input[4181]), .Z(n30085) );
  XOR U29905 ( .A(n30087), .B(n30088), .Z(n30083) );
  AND U29906 ( .A(n30089), .B(n30090), .Z(n30088) );
  XNOR U29907 ( .A(p_input[4212]), .B(n30087), .Z(n30090) );
  XOR U29908 ( .A(n30087), .B(p_input[4180]), .Z(n30089) );
  XOR U29909 ( .A(n30091), .B(n30092), .Z(n30087) );
  AND U29910 ( .A(n30093), .B(n30094), .Z(n30092) );
  XNOR U29911 ( .A(p_input[4211]), .B(n30091), .Z(n30094) );
  XOR U29912 ( .A(n30091), .B(p_input[4179]), .Z(n30093) );
  XOR U29913 ( .A(n30095), .B(n30096), .Z(n30091) );
  AND U29914 ( .A(n30097), .B(n30098), .Z(n30096) );
  XNOR U29915 ( .A(p_input[4210]), .B(n30095), .Z(n30098) );
  XOR U29916 ( .A(n30095), .B(p_input[4178]), .Z(n30097) );
  XOR U29917 ( .A(n30099), .B(n30100), .Z(n30095) );
  AND U29918 ( .A(n30101), .B(n30102), .Z(n30100) );
  XNOR U29919 ( .A(p_input[4209]), .B(n30099), .Z(n30102) );
  XOR U29920 ( .A(n30099), .B(p_input[4177]), .Z(n30101) );
  XOR U29921 ( .A(n30103), .B(n30104), .Z(n30099) );
  AND U29922 ( .A(n30105), .B(n30106), .Z(n30104) );
  XNOR U29923 ( .A(p_input[4208]), .B(n30103), .Z(n30106) );
  XOR U29924 ( .A(n30103), .B(p_input[4176]), .Z(n30105) );
  XOR U29925 ( .A(n30107), .B(n30108), .Z(n30103) );
  AND U29926 ( .A(n30109), .B(n30110), .Z(n30108) );
  XNOR U29927 ( .A(p_input[4207]), .B(n30107), .Z(n30110) );
  XOR U29928 ( .A(n30107), .B(p_input[4175]), .Z(n30109) );
  XOR U29929 ( .A(n30111), .B(n30112), .Z(n30107) );
  AND U29930 ( .A(n30113), .B(n30114), .Z(n30112) );
  XNOR U29931 ( .A(p_input[4206]), .B(n30111), .Z(n30114) );
  XOR U29932 ( .A(n30111), .B(p_input[4174]), .Z(n30113) );
  XOR U29933 ( .A(n30115), .B(n30116), .Z(n30111) );
  AND U29934 ( .A(n30117), .B(n30118), .Z(n30116) );
  XNOR U29935 ( .A(p_input[4205]), .B(n30115), .Z(n30118) );
  XOR U29936 ( .A(n30115), .B(p_input[4173]), .Z(n30117) );
  XOR U29937 ( .A(n30119), .B(n30120), .Z(n30115) );
  AND U29938 ( .A(n30121), .B(n30122), .Z(n30120) );
  XNOR U29939 ( .A(p_input[4204]), .B(n30119), .Z(n30122) );
  XOR U29940 ( .A(n30119), .B(p_input[4172]), .Z(n30121) );
  XOR U29941 ( .A(n30123), .B(n30124), .Z(n30119) );
  AND U29942 ( .A(n30125), .B(n30126), .Z(n30124) );
  XNOR U29943 ( .A(p_input[4203]), .B(n30123), .Z(n30126) );
  XOR U29944 ( .A(n30123), .B(p_input[4171]), .Z(n30125) );
  XOR U29945 ( .A(n30127), .B(n30128), .Z(n30123) );
  AND U29946 ( .A(n30129), .B(n30130), .Z(n30128) );
  XNOR U29947 ( .A(p_input[4202]), .B(n30127), .Z(n30130) );
  XOR U29948 ( .A(n30127), .B(p_input[4170]), .Z(n30129) );
  XOR U29949 ( .A(n30131), .B(n30132), .Z(n30127) );
  AND U29950 ( .A(n30133), .B(n30134), .Z(n30132) );
  XNOR U29951 ( .A(p_input[4201]), .B(n30131), .Z(n30134) );
  XOR U29952 ( .A(n30131), .B(p_input[4169]), .Z(n30133) );
  XOR U29953 ( .A(n30135), .B(n30136), .Z(n30131) );
  AND U29954 ( .A(n30137), .B(n30138), .Z(n30136) );
  XNOR U29955 ( .A(p_input[4200]), .B(n30135), .Z(n30138) );
  XOR U29956 ( .A(n30135), .B(p_input[4168]), .Z(n30137) );
  XOR U29957 ( .A(n30139), .B(n30140), .Z(n30135) );
  AND U29958 ( .A(n30141), .B(n30142), .Z(n30140) );
  XNOR U29959 ( .A(p_input[4199]), .B(n30139), .Z(n30142) );
  XOR U29960 ( .A(n30139), .B(p_input[4167]), .Z(n30141) );
  XOR U29961 ( .A(n30143), .B(n30144), .Z(n30139) );
  AND U29962 ( .A(n30145), .B(n30146), .Z(n30144) );
  XNOR U29963 ( .A(p_input[4198]), .B(n30143), .Z(n30146) );
  XOR U29964 ( .A(n30143), .B(p_input[4166]), .Z(n30145) );
  XOR U29965 ( .A(n30147), .B(n30148), .Z(n30143) );
  AND U29966 ( .A(n30149), .B(n30150), .Z(n30148) );
  XNOR U29967 ( .A(p_input[4197]), .B(n30147), .Z(n30150) );
  XOR U29968 ( .A(n30147), .B(p_input[4165]), .Z(n30149) );
  XOR U29969 ( .A(n30151), .B(n30152), .Z(n30147) );
  AND U29970 ( .A(n30153), .B(n30154), .Z(n30152) );
  XNOR U29971 ( .A(p_input[4196]), .B(n30151), .Z(n30154) );
  XOR U29972 ( .A(n30151), .B(p_input[4164]), .Z(n30153) );
  XOR U29973 ( .A(n30155), .B(n30156), .Z(n30151) );
  AND U29974 ( .A(n30157), .B(n30158), .Z(n30156) );
  XNOR U29975 ( .A(p_input[4195]), .B(n30155), .Z(n30158) );
  XOR U29976 ( .A(n30155), .B(p_input[4163]), .Z(n30157) );
  XOR U29977 ( .A(n30159), .B(n30160), .Z(n30155) );
  AND U29978 ( .A(n30161), .B(n30162), .Z(n30160) );
  XNOR U29979 ( .A(p_input[4194]), .B(n30159), .Z(n30162) );
  XOR U29980 ( .A(n30159), .B(p_input[4162]), .Z(n30161) );
  XNOR U29981 ( .A(n30163), .B(n30164), .Z(n30159) );
  AND U29982 ( .A(n30165), .B(n30166), .Z(n30164) );
  XOR U29983 ( .A(p_input[4193]), .B(n30163), .Z(n30166) );
  XNOR U29984 ( .A(p_input[4161]), .B(n30163), .Z(n30165) );
  AND U29985 ( .A(p_input[4192]), .B(n30167), .Z(n30163) );
  IV U29986 ( .A(p_input[4160]), .Z(n30167) );
  XNOR U29987 ( .A(p_input[4096]), .B(n30168), .Z(n29761) );
  AND U29988 ( .A(n412), .B(n30169), .Z(n30168) );
  XOR U29989 ( .A(p_input[4128]), .B(p_input[4096]), .Z(n30169) );
  XOR U29990 ( .A(n30170), .B(n30171), .Z(n412) );
  AND U29991 ( .A(n30172), .B(n30173), .Z(n30171) );
  XNOR U29992 ( .A(p_input[4159]), .B(n30170), .Z(n30173) );
  XOR U29993 ( .A(n30170), .B(p_input[4127]), .Z(n30172) );
  XOR U29994 ( .A(n30174), .B(n30175), .Z(n30170) );
  AND U29995 ( .A(n30176), .B(n30177), .Z(n30175) );
  XNOR U29996 ( .A(p_input[4158]), .B(n30174), .Z(n30177) );
  XNOR U29997 ( .A(n30174), .B(n29776), .Z(n30176) );
  IV U29998 ( .A(p_input[4126]), .Z(n29776) );
  XOR U29999 ( .A(n30178), .B(n30179), .Z(n30174) );
  AND U30000 ( .A(n30180), .B(n30181), .Z(n30179) );
  XNOR U30001 ( .A(p_input[4157]), .B(n30178), .Z(n30181) );
  XNOR U30002 ( .A(n30178), .B(n29785), .Z(n30180) );
  IV U30003 ( .A(p_input[4125]), .Z(n29785) );
  XOR U30004 ( .A(n30182), .B(n30183), .Z(n30178) );
  AND U30005 ( .A(n30184), .B(n30185), .Z(n30183) );
  XNOR U30006 ( .A(p_input[4156]), .B(n30182), .Z(n30185) );
  XNOR U30007 ( .A(n30182), .B(n29794), .Z(n30184) );
  IV U30008 ( .A(p_input[4124]), .Z(n29794) );
  XOR U30009 ( .A(n30186), .B(n30187), .Z(n30182) );
  AND U30010 ( .A(n30188), .B(n30189), .Z(n30187) );
  XNOR U30011 ( .A(p_input[4155]), .B(n30186), .Z(n30189) );
  XNOR U30012 ( .A(n30186), .B(n29803), .Z(n30188) );
  IV U30013 ( .A(p_input[4123]), .Z(n29803) );
  XOR U30014 ( .A(n30190), .B(n30191), .Z(n30186) );
  AND U30015 ( .A(n30192), .B(n30193), .Z(n30191) );
  XNOR U30016 ( .A(p_input[4154]), .B(n30190), .Z(n30193) );
  XNOR U30017 ( .A(n30190), .B(n29812), .Z(n30192) );
  IV U30018 ( .A(p_input[4122]), .Z(n29812) );
  XOR U30019 ( .A(n30194), .B(n30195), .Z(n30190) );
  AND U30020 ( .A(n30196), .B(n30197), .Z(n30195) );
  XNOR U30021 ( .A(p_input[4153]), .B(n30194), .Z(n30197) );
  XNOR U30022 ( .A(n30194), .B(n29821), .Z(n30196) );
  IV U30023 ( .A(p_input[4121]), .Z(n29821) );
  XOR U30024 ( .A(n30198), .B(n30199), .Z(n30194) );
  AND U30025 ( .A(n30200), .B(n30201), .Z(n30199) );
  XNOR U30026 ( .A(p_input[4152]), .B(n30198), .Z(n30201) );
  XNOR U30027 ( .A(n30198), .B(n29830), .Z(n30200) );
  IV U30028 ( .A(p_input[4120]), .Z(n29830) );
  XOR U30029 ( .A(n30202), .B(n30203), .Z(n30198) );
  AND U30030 ( .A(n30204), .B(n30205), .Z(n30203) );
  XNOR U30031 ( .A(p_input[4151]), .B(n30202), .Z(n30205) );
  XNOR U30032 ( .A(n30202), .B(n29839), .Z(n30204) );
  IV U30033 ( .A(p_input[4119]), .Z(n29839) );
  XOR U30034 ( .A(n30206), .B(n30207), .Z(n30202) );
  AND U30035 ( .A(n30208), .B(n30209), .Z(n30207) );
  XNOR U30036 ( .A(p_input[4150]), .B(n30206), .Z(n30209) );
  XNOR U30037 ( .A(n30206), .B(n29848), .Z(n30208) );
  IV U30038 ( .A(p_input[4118]), .Z(n29848) );
  XOR U30039 ( .A(n30210), .B(n30211), .Z(n30206) );
  AND U30040 ( .A(n30212), .B(n30213), .Z(n30211) );
  XNOR U30041 ( .A(p_input[4149]), .B(n30210), .Z(n30213) );
  XNOR U30042 ( .A(n30210), .B(n29857), .Z(n30212) );
  IV U30043 ( .A(p_input[4117]), .Z(n29857) );
  XOR U30044 ( .A(n30214), .B(n30215), .Z(n30210) );
  AND U30045 ( .A(n30216), .B(n30217), .Z(n30215) );
  XNOR U30046 ( .A(p_input[4148]), .B(n30214), .Z(n30217) );
  XNOR U30047 ( .A(n30214), .B(n29866), .Z(n30216) );
  IV U30048 ( .A(p_input[4116]), .Z(n29866) );
  XOR U30049 ( .A(n30218), .B(n30219), .Z(n30214) );
  AND U30050 ( .A(n30220), .B(n30221), .Z(n30219) );
  XNOR U30051 ( .A(p_input[4147]), .B(n30218), .Z(n30221) );
  XNOR U30052 ( .A(n30218), .B(n29875), .Z(n30220) );
  IV U30053 ( .A(p_input[4115]), .Z(n29875) );
  XOR U30054 ( .A(n30222), .B(n30223), .Z(n30218) );
  AND U30055 ( .A(n30224), .B(n30225), .Z(n30223) );
  XNOR U30056 ( .A(p_input[4146]), .B(n30222), .Z(n30225) );
  XNOR U30057 ( .A(n30222), .B(n29884), .Z(n30224) );
  IV U30058 ( .A(p_input[4114]), .Z(n29884) );
  XOR U30059 ( .A(n30226), .B(n30227), .Z(n30222) );
  AND U30060 ( .A(n30228), .B(n30229), .Z(n30227) );
  XNOR U30061 ( .A(p_input[4145]), .B(n30226), .Z(n30229) );
  XNOR U30062 ( .A(n30226), .B(n29893), .Z(n30228) );
  IV U30063 ( .A(p_input[4113]), .Z(n29893) );
  XOR U30064 ( .A(n30230), .B(n30231), .Z(n30226) );
  AND U30065 ( .A(n30232), .B(n30233), .Z(n30231) );
  XNOR U30066 ( .A(p_input[4144]), .B(n30230), .Z(n30233) );
  XNOR U30067 ( .A(n30230), .B(n29902), .Z(n30232) );
  IV U30068 ( .A(p_input[4112]), .Z(n29902) );
  XOR U30069 ( .A(n30234), .B(n30235), .Z(n30230) );
  AND U30070 ( .A(n30236), .B(n30237), .Z(n30235) );
  XNOR U30071 ( .A(p_input[4143]), .B(n30234), .Z(n30237) );
  XNOR U30072 ( .A(n30234), .B(n29911), .Z(n30236) );
  IV U30073 ( .A(p_input[4111]), .Z(n29911) );
  XOR U30074 ( .A(n30238), .B(n30239), .Z(n30234) );
  AND U30075 ( .A(n30240), .B(n30241), .Z(n30239) );
  XNOR U30076 ( .A(p_input[4142]), .B(n30238), .Z(n30241) );
  XNOR U30077 ( .A(n30238), .B(n29920), .Z(n30240) );
  IV U30078 ( .A(p_input[4110]), .Z(n29920) );
  XOR U30079 ( .A(n30242), .B(n30243), .Z(n30238) );
  AND U30080 ( .A(n30244), .B(n30245), .Z(n30243) );
  XNOR U30081 ( .A(p_input[4141]), .B(n30242), .Z(n30245) );
  XNOR U30082 ( .A(n30242), .B(n29929), .Z(n30244) );
  IV U30083 ( .A(p_input[4109]), .Z(n29929) );
  XOR U30084 ( .A(n30246), .B(n30247), .Z(n30242) );
  AND U30085 ( .A(n30248), .B(n30249), .Z(n30247) );
  XNOR U30086 ( .A(p_input[4140]), .B(n30246), .Z(n30249) );
  XNOR U30087 ( .A(n30246), .B(n29938), .Z(n30248) );
  IV U30088 ( .A(p_input[4108]), .Z(n29938) );
  XOR U30089 ( .A(n30250), .B(n30251), .Z(n30246) );
  AND U30090 ( .A(n30252), .B(n30253), .Z(n30251) );
  XNOR U30091 ( .A(p_input[4139]), .B(n30250), .Z(n30253) );
  XNOR U30092 ( .A(n30250), .B(n29947), .Z(n30252) );
  IV U30093 ( .A(p_input[4107]), .Z(n29947) );
  XOR U30094 ( .A(n30254), .B(n30255), .Z(n30250) );
  AND U30095 ( .A(n30256), .B(n30257), .Z(n30255) );
  XNOR U30096 ( .A(p_input[4138]), .B(n30254), .Z(n30257) );
  XNOR U30097 ( .A(n30254), .B(n29956), .Z(n30256) );
  IV U30098 ( .A(p_input[4106]), .Z(n29956) );
  XOR U30099 ( .A(n30258), .B(n30259), .Z(n30254) );
  AND U30100 ( .A(n30260), .B(n30261), .Z(n30259) );
  XNOR U30101 ( .A(p_input[4137]), .B(n30258), .Z(n30261) );
  XNOR U30102 ( .A(n30258), .B(n29965), .Z(n30260) );
  IV U30103 ( .A(p_input[4105]), .Z(n29965) );
  XOR U30104 ( .A(n30262), .B(n30263), .Z(n30258) );
  AND U30105 ( .A(n30264), .B(n30265), .Z(n30263) );
  XNOR U30106 ( .A(p_input[4136]), .B(n30262), .Z(n30265) );
  XNOR U30107 ( .A(n30262), .B(n29974), .Z(n30264) );
  IV U30108 ( .A(p_input[4104]), .Z(n29974) );
  XOR U30109 ( .A(n30266), .B(n30267), .Z(n30262) );
  AND U30110 ( .A(n30268), .B(n30269), .Z(n30267) );
  XNOR U30111 ( .A(p_input[4135]), .B(n30266), .Z(n30269) );
  XNOR U30112 ( .A(n30266), .B(n29983), .Z(n30268) );
  IV U30113 ( .A(p_input[4103]), .Z(n29983) );
  XOR U30114 ( .A(n30270), .B(n30271), .Z(n30266) );
  AND U30115 ( .A(n30272), .B(n30273), .Z(n30271) );
  XNOR U30116 ( .A(p_input[4134]), .B(n30270), .Z(n30273) );
  XNOR U30117 ( .A(n30270), .B(n29992), .Z(n30272) );
  IV U30118 ( .A(p_input[4102]), .Z(n29992) );
  XOR U30119 ( .A(n30274), .B(n30275), .Z(n30270) );
  AND U30120 ( .A(n30276), .B(n30277), .Z(n30275) );
  XNOR U30121 ( .A(p_input[4133]), .B(n30274), .Z(n30277) );
  XNOR U30122 ( .A(n30274), .B(n30001), .Z(n30276) );
  IV U30123 ( .A(p_input[4101]), .Z(n30001) );
  XOR U30124 ( .A(n30278), .B(n30279), .Z(n30274) );
  AND U30125 ( .A(n30280), .B(n30281), .Z(n30279) );
  XNOR U30126 ( .A(p_input[4132]), .B(n30278), .Z(n30281) );
  XNOR U30127 ( .A(n30278), .B(n30010), .Z(n30280) );
  IV U30128 ( .A(p_input[4100]), .Z(n30010) );
  XOR U30129 ( .A(n30282), .B(n30283), .Z(n30278) );
  AND U30130 ( .A(n30284), .B(n30285), .Z(n30283) );
  XNOR U30131 ( .A(p_input[4131]), .B(n30282), .Z(n30285) );
  XNOR U30132 ( .A(n30282), .B(n30019), .Z(n30284) );
  IV U30133 ( .A(p_input[4099]), .Z(n30019) );
  XOR U30134 ( .A(n30286), .B(n30287), .Z(n30282) );
  AND U30135 ( .A(n30288), .B(n30289), .Z(n30287) );
  XNOR U30136 ( .A(p_input[4130]), .B(n30286), .Z(n30289) );
  XNOR U30137 ( .A(n30286), .B(n30028), .Z(n30288) );
  IV U30138 ( .A(p_input[4098]), .Z(n30028) );
  XNOR U30139 ( .A(n30290), .B(n30291), .Z(n30286) );
  AND U30140 ( .A(n30292), .B(n30293), .Z(n30291) );
  XOR U30141 ( .A(p_input[4129]), .B(n30290), .Z(n30293) );
  XNOR U30142 ( .A(p_input[4097]), .B(n30290), .Z(n30292) );
  AND U30143 ( .A(p_input[4128]), .B(n30294), .Z(n30290) );
  IV U30144 ( .A(p_input[4096]), .Z(n30294) );
  XOR U30145 ( .A(n30295), .B(n30296), .Z(n7) );
  AND U30146 ( .A(n1140), .B(n30297), .Z(n30296) );
  XNOR U30147 ( .A(n30298), .B(n30295), .Z(n30297) );
  XOR U30148 ( .A(n30299), .B(n30300), .Z(n1140) );
  AND U30149 ( .A(n30301), .B(n30302), .Z(n30300) );
  XOR U30150 ( .A(n30299), .B(n1159), .Z(n30302) );
  XOR U30151 ( .A(n30303), .B(n30304), .Z(n1159) );
  AND U30152 ( .A(n1131), .B(n30305), .Z(n30304) );
  XOR U30153 ( .A(n30306), .B(n30303), .Z(n30305) );
  XNOR U30154 ( .A(n1156), .B(n30299), .Z(n30301) );
  XOR U30155 ( .A(n30307), .B(n30308), .Z(n1156) );
  AND U30156 ( .A(n1128), .B(n30309), .Z(n30308) );
  XOR U30157 ( .A(n30310), .B(n30307), .Z(n30309) );
  XOR U30158 ( .A(n30311), .B(n30312), .Z(n30299) );
  AND U30159 ( .A(n30313), .B(n30314), .Z(n30312) );
  XOR U30160 ( .A(n30311), .B(n1171), .Z(n30314) );
  XOR U30161 ( .A(n30315), .B(n30316), .Z(n1171) );
  AND U30162 ( .A(n1131), .B(n30317), .Z(n30316) );
  XOR U30163 ( .A(n30318), .B(n30315), .Z(n30317) );
  XNOR U30164 ( .A(n1168), .B(n30311), .Z(n30313) );
  XOR U30165 ( .A(n30319), .B(n30320), .Z(n1168) );
  AND U30166 ( .A(n1128), .B(n30321), .Z(n30320) );
  XOR U30167 ( .A(n30322), .B(n30319), .Z(n30321) );
  XOR U30168 ( .A(n30323), .B(n30324), .Z(n30311) );
  AND U30169 ( .A(n30325), .B(n30326), .Z(n30324) );
  XOR U30170 ( .A(n30323), .B(n1183), .Z(n30326) );
  XOR U30171 ( .A(n30327), .B(n30328), .Z(n1183) );
  AND U30172 ( .A(n1131), .B(n30329), .Z(n30328) );
  XOR U30173 ( .A(n30330), .B(n30327), .Z(n30329) );
  XNOR U30174 ( .A(n1180), .B(n30323), .Z(n30325) );
  XOR U30175 ( .A(n30331), .B(n30332), .Z(n1180) );
  AND U30176 ( .A(n1128), .B(n30333), .Z(n30332) );
  XOR U30177 ( .A(n30334), .B(n30331), .Z(n30333) );
  XOR U30178 ( .A(n30335), .B(n30336), .Z(n30323) );
  AND U30179 ( .A(n30337), .B(n30338), .Z(n30336) );
  XOR U30180 ( .A(n30335), .B(n1195), .Z(n30338) );
  XOR U30181 ( .A(n30339), .B(n30340), .Z(n1195) );
  AND U30182 ( .A(n1131), .B(n30341), .Z(n30340) );
  XOR U30183 ( .A(n30342), .B(n30339), .Z(n30341) );
  XNOR U30184 ( .A(n1192), .B(n30335), .Z(n30337) );
  XOR U30185 ( .A(n30343), .B(n30344), .Z(n1192) );
  AND U30186 ( .A(n1128), .B(n30345), .Z(n30344) );
  XOR U30187 ( .A(n30346), .B(n30343), .Z(n30345) );
  XOR U30188 ( .A(n30347), .B(n30348), .Z(n30335) );
  AND U30189 ( .A(n30349), .B(n30350), .Z(n30348) );
  XOR U30190 ( .A(n30347), .B(n1207), .Z(n30350) );
  XOR U30191 ( .A(n30351), .B(n30352), .Z(n1207) );
  AND U30192 ( .A(n1131), .B(n30353), .Z(n30352) );
  XOR U30193 ( .A(n30354), .B(n30351), .Z(n30353) );
  XNOR U30194 ( .A(n1204), .B(n30347), .Z(n30349) );
  XOR U30195 ( .A(n30355), .B(n30356), .Z(n1204) );
  AND U30196 ( .A(n1128), .B(n30357), .Z(n30356) );
  XOR U30197 ( .A(n30358), .B(n30355), .Z(n30357) );
  XOR U30198 ( .A(n30359), .B(n30360), .Z(n30347) );
  AND U30199 ( .A(n30361), .B(n30362), .Z(n30360) );
  XOR U30200 ( .A(n30359), .B(n1219), .Z(n30362) );
  XOR U30201 ( .A(n30363), .B(n30364), .Z(n1219) );
  AND U30202 ( .A(n1131), .B(n30365), .Z(n30364) );
  XOR U30203 ( .A(n30366), .B(n30363), .Z(n30365) );
  XNOR U30204 ( .A(n1216), .B(n30359), .Z(n30361) );
  XOR U30205 ( .A(n30367), .B(n30368), .Z(n1216) );
  AND U30206 ( .A(n1128), .B(n30369), .Z(n30368) );
  XOR U30207 ( .A(n30370), .B(n30367), .Z(n30369) );
  XOR U30208 ( .A(n30371), .B(n30372), .Z(n30359) );
  AND U30209 ( .A(n30373), .B(n30374), .Z(n30372) );
  XOR U30210 ( .A(n30371), .B(n1231), .Z(n30374) );
  XOR U30211 ( .A(n30375), .B(n30376), .Z(n1231) );
  AND U30212 ( .A(n1131), .B(n30377), .Z(n30376) );
  XOR U30213 ( .A(n30378), .B(n30375), .Z(n30377) );
  XNOR U30214 ( .A(n1228), .B(n30371), .Z(n30373) );
  XOR U30215 ( .A(n30379), .B(n30380), .Z(n1228) );
  AND U30216 ( .A(n1128), .B(n30381), .Z(n30380) );
  XOR U30217 ( .A(n30382), .B(n30379), .Z(n30381) );
  XOR U30218 ( .A(n30383), .B(n30384), .Z(n30371) );
  AND U30219 ( .A(n30385), .B(n30386), .Z(n30384) );
  XOR U30220 ( .A(n30383), .B(n1243), .Z(n30386) );
  XOR U30221 ( .A(n30387), .B(n30388), .Z(n1243) );
  AND U30222 ( .A(n1131), .B(n30389), .Z(n30388) );
  XOR U30223 ( .A(n30390), .B(n30387), .Z(n30389) );
  XNOR U30224 ( .A(n1240), .B(n30383), .Z(n30385) );
  XOR U30225 ( .A(n30391), .B(n30392), .Z(n1240) );
  AND U30226 ( .A(n1128), .B(n30393), .Z(n30392) );
  XOR U30227 ( .A(n30394), .B(n30391), .Z(n30393) );
  XOR U30228 ( .A(n30395), .B(n30396), .Z(n30383) );
  AND U30229 ( .A(n30397), .B(n30398), .Z(n30396) );
  XOR U30230 ( .A(n30395), .B(n1255), .Z(n30398) );
  XOR U30231 ( .A(n30399), .B(n30400), .Z(n1255) );
  AND U30232 ( .A(n1131), .B(n30401), .Z(n30400) );
  XOR U30233 ( .A(n30402), .B(n30399), .Z(n30401) );
  XNOR U30234 ( .A(n1252), .B(n30395), .Z(n30397) );
  XOR U30235 ( .A(n30403), .B(n30404), .Z(n1252) );
  AND U30236 ( .A(n1128), .B(n30405), .Z(n30404) );
  XOR U30237 ( .A(n30406), .B(n30403), .Z(n30405) );
  XOR U30238 ( .A(n30407), .B(n30408), .Z(n30395) );
  AND U30239 ( .A(n30409), .B(n30410), .Z(n30408) );
  XOR U30240 ( .A(n30407), .B(n1267), .Z(n30410) );
  XOR U30241 ( .A(n30411), .B(n30412), .Z(n1267) );
  AND U30242 ( .A(n1131), .B(n30413), .Z(n30412) );
  XOR U30243 ( .A(n30414), .B(n30411), .Z(n30413) );
  XNOR U30244 ( .A(n1264), .B(n30407), .Z(n30409) );
  XOR U30245 ( .A(n30415), .B(n30416), .Z(n1264) );
  AND U30246 ( .A(n1128), .B(n30417), .Z(n30416) );
  XOR U30247 ( .A(n30418), .B(n30415), .Z(n30417) );
  XOR U30248 ( .A(n30419), .B(n30420), .Z(n30407) );
  AND U30249 ( .A(n30421), .B(n30422), .Z(n30420) );
  XOR U30250 ( .A(n30419), .B(n1279), .Z(n30422) );
  XOR U30251 ( .A(n30423), .B(n30424), .Z(n1279) );
  AND U30252 ( .A(n1131), .B(n30425), .Z(n30424) );
  XOR U30253 ( .A(n30426), .B(n30423), .Z(n30425) );
  XNOR U30254 ( .A(n1276), .B(n30419), .Z(n30421) );
  XOR U30255 ( .A(n30427), .B(n30428), .Z(n1276) );
  AND U30256 ( .A(n1128), .B(n30429), .Z(n30428) );
  XOR U30257 ( .A(n30430), .B(n30427), .Z(n30429) );
  XOR U30258 ( .A(n30431), .B(n30432), .Z(n30419) );
  AND U30259 ( .A(n30433), .B(n30434), .Z(n30432) );
  XOR U30260 ( .A(n30431), .B(n1291), .Z(n30434) );
  XOR U30261 ( .A(n30435), .B(n30436), .Z(n1291) );
  AND U30262 ( .A(n1131), .B(n30437), .Z(n30436) );
  XOR U30263 ( .A(n30438), .B(n30435), .Z(n30437) );
  XNOR U30264 ( .A(n1288), .B(n30431), .Z(n30433) );
  XOR U30265 ( .A(n30439), .B(n30440), .Z(n1288) );
  AND U30266 ( .A(n1128), .B(n30441), .Z(n30440) );
  XOR U30267 ( .A(n30442), .B(n30439), .Z(n30441) );
  XOR U30268 ( .A(n30443), .B(n30444), .Z(n30431) );
  AND U30269 ( .A(n30445), .B(n30446), .Z(n30444) );
  XOR U30270 ( .A(n30443), .B(n1303), .Z(n30446) );
  XOR U30271 ( .A(n30447), .B(n30448), .Z(n1303) );
  AND U30272 ( .A(n1131), .B(n30449), .Z(n30448) );
  XOR U30273 ( .A(n30450), .B(n30447), .Z(n30449) );
  XNOR U30274 ( .A(n1300), .B(n30443), .Z(n30445) );
  XOR U30275 ( .A(n30451), .B(n30452), .Z(n1300) );
  AND U30276 ( .A(n1128), .B(n30453), .Z(n30452) );
  XOR U30277 ( .A(n30454), .B(n30451), .Z(n30453) );
  XOR U30278 ( .A(n30455), .B(n30456), .Z(n30443) );
  AND U30279 ( .A(n30457), .B(n30458), .Z(n30456) );
  XOR U30280 ( .A(n30455), .B(n1315), .Z(n30458) );
  XOR U30281 ( .A(n30459), .B(n30460), .Z(n1315) );
  AND U30282 ( .A(n1131), .B(n30461), .Z(n30460) );
  XOR U30283 ( .A(n30462), .B(n30459), .Z(n30461) );
  XNOR U30284 ( .A(n1312), .B(n30455), .Z(n30457) );
  XOR U30285 ( .A(n30463), .B(n30464), .Z(n1312) );
  AND U30286 ( .A(n1128), .B(n30465), .Z(n30464) );
  XOR U30287 ( .A(n30466), .B(n30463), .Z(n30465) );
  XOR U30288 ( .A(n30467), .B(n30468), .Z(n30455) );
  AND U30289 ( .A(n30469), .B(n30470), .Z(n30468) );
  XOR U30290 ( .A(n30467), .B(n1327), .Z(n30470) );
  XOR U30291 ( .A(n30471), .B(n30472), .Z(n1327) );
  AND U30292 ( .A(n1131), .B(n30473), .Z(n30472) );
  XOR U30293 ( .A(n30474), .B(n30471), .Z(n30473) );
  XNOR U30294 ( .A(n1324), .B(n30467), .Z(n30469) );
  XOR U30295 ( .A(n30475), .B(n30476), .Z(n1324) );
  AND U30296 ( .A(n1128), .B(n30477), .Z(n30476) );
  XOR U30297 ( .A(n30478), .B(n30475), .Z(n30477) );
  XOR U30298 ( .A(n30479), .B(n30480), .Z(n30467) );
  AND U30299 ( .A(n30481), .B(n30482), .Z(n30480) );
  XOR U30300 ( .A(n30479), .B(n1339), .Z(n30482) );
  XOR U30301 ( .A(n30483), .B(n30484), .Z(n1339) );
  AND U30302 ( .A(n1131), .B(n30485), .Z(n30484) );
  XOR U30303 ( .A(n30486), .B(n30483), .Z(n30485) );
  XNOR U30304 ( .A(n1336), .B(n30479), .Z(n30481) );
  XOR U30305 ( .A(n30487), .B(n30488), .Z(n1336) );
  AND U30306 ( .A(n1128), .B(n30489), .Z(n30488) );
  XOR U30307 ( .A(n30490), .B(n30487), .Z(n30489) );
  XOR U30308 ( .A(n30491), .B(n30492), .Z(n30479) );
  AND U30309 ( .A(n30493), .B(n30494), .Z(n30492) );
  XOR U30310 ( .A(n30491), .B(n1351), .Z(n30494) );
  XOR U30311 ( .A(n30495), .B(n30496), .Z(n1351) );
  AND U30312 ( .A(n1131), .B(n30497), .Z(n30496) );
  XOR U30313 ( .A(n30498), .B(n30495), .Z(n30497) );
  XNOR U30314 ( .A(n1348), .B(n30491), .Z(n30493) );
  XOR U30315 ( .A(n30499), .B(n30500), .Z(n1348) );
  AND U30316 ( .A(n1128), .B(n30501), .Z(n30500) );
  XOR U30317 ( .A(n30502), .B(n30499), .Z(n30501) );
  XOR U30318 ( .A(n30503), .B(n30504), .Z(n30491) );
  AND U30319 ( .A(n30505), .B(n30506), .Z(n30504) );
  XOR U30320 ( .A(n30503), .B(n1363), .Z(n30506) );
  XOR U30321 ( .A(n30507), .B(n30508), .Z(n1363) );
  AND U30322 ( .A(n1131), .B(n30509), .Z(n30508) );
  XOR U30323 ( .A(n30510), .B(n30507), .Z(n30509) );
  XNOR U30324 ( .A(n1360), .B(n30503), .Z(n30505) );
  XOR U30325 ( .A(n30511), .B(n30512), .Z(n1360) );
  AND U30326 ( .A(n1128), .B(n30513), .Z(n30512) );
  XOR U30327 ( .A(n30514), .B(n30511), .Z(n30513) );
  XOR U30328 ( .A(n30515), .B(n30516), .Z(n30503) );
  AND U30329 ( .A(n30517), .B(n30518), .Z(n30516) );
  XOR U30330 ( .A(n30515), .B(n1375), .Z(n30518) );
  XOR U30331 ( .A(n30519), .B(n30520), .Z(n1375) );
  AND U30332 ( .A(n1131), .B(n30521), .Z(n30520) );
  XOR U30333 ( .A(n30522), .B(n30519), .Z(n30521) );
  XNOR U30334 ( .A(n1372), .B(n30515), .Z(n30517) );
  XOR U30335 ( .A(n30523), .B(n30524), .Z(n1372) );
  AND U30336 ( .A(n1128), .B(n30525), .Z(n30524) );
  XOR U30337 ( .A(n30526), .B(n30523), .Z(n30525) );
  XOR U30338 ( .A(n30527), .B(n30528), .Z(n30515) );
  AND U30339 ( .A(n30529), .B(n30530), .Z(n30528) );
  XOR U30340 ( .A(n30527), .B(n1387), .Z(n30530) );
  XOR U30341 ( .A(n30531), .B(n30532), .Z(n1387) );
  AND U30342 ( .A(n1131), .B(n30533), .Z(n30532) );
  XOR U30343 ( .A(n30534), .B(n30531), .Z(n30533) );
  XNOR U30344 ( .A(n1384), .B(n30527), .Z(n30529) );
  XOR U30345 ( .A(n30535), .B(n30536), .Z(n1384) );
  AND U30346 ( .A(n1128), .B(n30537), .Z(n30536) );
  XOR U30347 ( .A(n30538), .B(n30535), .Z(n30537) );
  XOR U30348 ( .A(n30539), .B(n30540), .Z(n30527) );
  AND U30349 ( .A(n30541), .B(n30542), .Z(n30540) );
  XOR U30350 ( .A(n30539), .B(n1399), .Z(n30542) );
  XOR U30351 ( .A(n30543), .B(n30544), .Z(n1399) );
  AND U30352 ( .A(n1131), .B(n30545), .Z(n30544) );
  XOR U30353 ( .A(n30546), .B(n30543), .Z(n30545) );
  XNOR U30354 ( .A(n1396), .B(n30539), .Z(n30541) );
  XOR U30355 ( .A(n30547), .B(n30548), .Z(n1396) );
  AND U30356 ( .A(n1128), .B(n30549), .Z(n30548) );
  XOR U30357 ( .A(n30550), .B(n30547), .Z(n30549) );
  XOR U30358 ( .A(n30551), .B(n30552), .Z(n30539) );
  AND U30359 ( .A(n30553), .B(n30554), .Z(n30552) );
  XOR U30360 ( .A(n30551), .B(n1411), .Z(n30554) );
  XOR U30361 ( .A(n30555), .B(n30556), .Z(n1411) );
  AND U30362 ( .A(n1131), .B(n30557), .Z(n30556) );
  XOR U30363 ( .A(n30558), .B(n30555), .Z(n30557) );
  XNOR U30364 ( .A(n1408), .B(n30551), .Z(n30553) );
  XOR U30365 ( .A(n30559), .B(n30560), .Z(n1408) );
  AND U30366 ( .A(n1128), .B(n30561), .Z(n30560) );
  XOR U30367 ( .A(n30562), .B(n30559), .Z(n30561) );
  XOR U30368 ( .A(n30563), .B(n30564), .Z(n30551) );
  AND U30369 ( .A(n30565), .B(n30566), .Z(n30564) );
  XOR U30370 ( .A(n30563), .B(n1423), .Z(n30566) );
  XOR U30371 ( .A(n30567), .B(n30568), .Z(n1423) );
  AND U30372 ( .A(n1131), .B(n30569), .Z(n30568) );
  XOR U30373 ( .A(n30570), .B(n30567), .Z(n30569) );
  XNOR U30374 ( .A(n1420), .B(n30563), .Z(n30565) );
  XOR U30375 ( .A(n30571), .B(n30572), .Z(n1420) );
  AND U30376 ( .A(n1128), .B(n30573), .Z(n30572) );
  XOR U30377 ( .A(n30574), .B(n30571), .Z(n30573) );
  XOR U30378 ( .A(n30575), .B(n30576), .Z(n30563) );
  AND U30379 ( .A(n30577), .B(n30578), .Z(n30576) );
  XOR U30380 ( .A(n30575), .B(n1435), .Z(n30578) );
  XOR U30381 ( .A(n30579), .B(n30580), .Z(n1435) );
  AND U30382 ( .A(n1131), .B(n30581), .Z(n30580) );
  XOR U30383 ( .A(n30582), .B(n30579), .Z(n30581) );
  XNOR U30384 ( .A(n1432), .B(n30575), .Z(n30577) );
  XOR U30385 ( .A(n30583), .B(n30584), .Z(n1432) );
  AND U30386 ( .A(n1128), .B(n30585), .Z(n30584) );
  XOR U30387 ( .A(n30586), .B(n30583), .Z(n30585) );
  XOR U30388 ( .A(n30587), .B(n30588), .Z(n30575) );
  AND U30389 ( .A(n30589), .B(n30590), .Z(n30588) );
  XOR U30390 ( .A(n30587), .B(n1447), .Z(n30590) );
  XOR U30391 ( .A(n30591), .B(n30592), .Z(n1447) );
  AND U30392 ( .A(n1131), .B(n30593), .Z(n30592) );
  XOR U30393 ( .A(n30594), .B(n30591), .Z(n30593) );
  XNOR U30394 ( .A(n1444), .B(n30587), .Z(n30589) );
  XOR U30395 ( .A(n30595), .B(n30596), .Z(n1444) );
  AND U30396 ( .A(n1128), .B(n30597), .Z(n30596) );
  XOR U30397 ( .A(n30598), .B(n30595), .Z(n30597) );
  XOR U30398 ( .A(n30599), .B(n30600), .Z(n30587) );
  AND U30399 ( .A(n30601), .B(n30602), .Z(n30600) );
  XOR U30400 ( .A(n30599), .B(n1459), .Z(n30602) );
  XOR U30401 ( .A(n30603), .B(n30604), .Z(n1459) );
  AND U30402 ( .A(n1131), .B(n30605), .Z(n30604) );
  XOR U30403 ( .A(n30606), .B(n30603), .Z(n30605) );
  XNOR U30404 ( .A(n1456), .B(n30599), .Z(n30601) );
  XOR U30405 ( .A(n30607), .B(n30608), .Z(n1456) );
  AND U30406 ( .A(n1128), .B(n30609), .Z(n30608) );
  XOR U30407 ( .A(n30610), .B(n30607), .Z(n30609) );
  XOR U30408 ( .A(n30611), .B(n30612), .Z(n30599) );
  AND U30409 ( .A(n30613), .B(n30614), .Z(n30612) );
  XOR U30410 ( .A(n30611), .B(n1471), .Z(n30614) );
  XOR U30411 ( .A(n30615), .B(n30616), .Z(n1471) );
  AND U30412 ( .A(n1131), .B(n30617), .Z(n30616) );
  XOR U30413 ( .A(n30618), .B(n30615), .Z(n30617) );
  XNOR U30414 ( .A(n1468), .B(n30611), .Z(n30613) );
  XOR U30415 ( .A(n30619), .B(n30620), .Z(n1468) );
  AND U30416 ( .A(n1128), .B(n30621), .Z(n30620) );
  XOR U30417 ( .A(n30622), .B(n30619), .Z(n30621) );
  XOR U30418 ( .A(n30623), .B(n30624), .Z(n30611) );
  AND U30419 ( .A(n30625), .B(n30626), .Z(n30624) );
  XOR U30420 ( .A(n30623), .B(n1483), .Z(n30626) );
  XOR U30421 ( .A(n30627), .B(n30628), .Z(n1483) );
  AND U30422 ( .A(n1131), .B(n30629), .Z(n30628) );
  XOR U30423 ( .A(n30630), .B(n30627), .Z(n30629) );
  XNOR U30424 ( .A(n1480), .B(n30623), .Z(n30625) );
  XOR U30425 ( .A(n30631), .B(n30632), .Z(n1480) );
  AND U30426 ( .A(n1128), .B(n30633), .Z(n30632) );
  XOR U30427 ( .A(n30634), .B(n30631), .Z(n30633) );
  XOR U30428 ( .A(n30635), .B(n30636), .Z(n30623) );
  AND U30429 ( .A(n30637), .B(n30638), .Z(n30636) );
  XOR U30430 ( .A(n30635), .B(n1495), .Z(n30638) );
  XOR U30431 ( .A(n30639), .B(n30640), .Z(n1495) );
  AND U30432 ( .A(n1131), .B(n30641), .Z(n30640) );
  XOR U30433 ( .A(n30642), .B(n30639), .Z(n30641) );
  XNOR U30434 ( .A(n1492), .B(n30635), .Z(n30637) );
  XOR U30435 ( .A(n30643), .B(n30644), .Z(n1492) );
  AND U30436 ( .A(n1128), .B(n30645), .Z(n30644) );
  XOR U30437 ( .A(n30646), .B(n30643), .Z(n30645) );
  XOR U30438 ( .A(n30647), .B(n30648), .Z(n30635) );
  AND U30439 ( .A(n30649), .B(n30650), .Z(n30648) );
  XOR U30440 ( .A(n30647), .B(n1507), .Z(n30650) );
  XOR U30441 ( .A(n30651), .B(n30652), .Z(n1507) );
  AND U30442 ( .A(n1131), .B(n30653), .Z(n30652) );
  XOR U30443 ( .A(n30654), .B(n30651), .Z(n30653) );
  XNOR U30444 ( .A(n1504), .B(n30647), .Z(n30649) );
  XOR U30445 ( .A(n30655), .B(n30656), .Z(n1504) );
  AND U30446 ( .A(n1128), .B(n30657), .Z(n30656) );
  XOR U30447 ( .A(n30658), .B(n30655), .Z(n30657) );
  XOR U30448 ( .A(n30659), .B(n30660), .Z(n30647) );
  AND U30449 ( .A(n30661), .B(n30662), .Z(n30660) );
  XNOR U30450 ( .A(n30663), .B(n1519), .Z(n30662) );
  XOR U30451 ( .A(n30664), .B(n30665), .Z(n1519) );
  AND U30452 ( .A(n1131), .B(n30666), .Z(n30665) );
  XOR U30453 ( .A(n30664), .B(n30667), .Z(n30666) );
  XNOR U30454 ( .A(n1516), .B(n30659), .Z(n30661) );
  XOR U30455 ( .A(n30668), .B(n30669), .Z(n1516) );
  AND U30456 ( .A(n1128), .B(n30670), .Z(n30669) );
  XOR U30457 ( .A(n30668), .B(n30671), .Z(n30670) );
  IV U30458 ( .A(n30663), .Z(n30659) );
  AND U30459 ( .A(n30295), .B(n30298), .Z(n30663) );
  XNOR U30460 ( .A(n30672), .B(n30673), .Z(n30298) );
  AND U30461 ( .A(n1131), .B(n30674), .Z(n30673) );
  XNOR U30462 ( .A(n30675), .B(n30672), .Z(n30674) );
  XOR U30463 ( .A(n30676), .B(n30677), .Z(n1131) );
  AND U30464 ( .A(n30678), .B(n30679), .Z(n30677) );
  XOR U30465 ( .A(n30676), .B(n30306), .Z(n30679) );
  XOR U30466 ( .A(n30680), .B(n30681), .Z(n30306) );
  AND U30467 ( .A(n1099), .B(n30682), .Z(n30681) );
  XOR U30468 ( .A(n30683), .B(n30680), .Z(n30682) );
  XNOR U30469 ( .A(n30303), .B(n30676), .Z(n30678) );
  XOR U30470 ( .A(n30684), .B(n30685), .Z(n30303) );
  AND U30471 ( .A(n1097), .B(n30686), .Z(n30685) );
  XOR U30472 ( .A(n30687), .B(n30684), .Z(n30686) );
  XOR U30473 ( .A(n30688), .B(n30689), .Z(n30676) );
  AND U30474 ( .A(n30690), .B(n30691), .Z(n30689) );
  XOR U30475 ( .A(n30688), .B(n30318), .Z(n30691) );
  XOR U30476 ( .A(n30692), .B(n30693), .Z(n30318) );
  AND U30477 ( .A(n1099), .B(n30694), .Z(n30693) );
  XOR U30478 ( .A(n30695), .B(n30692), .Z(n30694) );
  XNOR U30479 ( .A(n30315), .B(n30688), .Z(n30690) );
  XOR U30480 ( .A(n30696), .B(n30697), .Z(n30315) );
  AND U30481 ( .A(n1097), .B(n30698), .Z(n30697) );
  XOR U30482 ( .A(n30699), .B(n30696), .Z(n30698) );
  XOR U30483 ( .A(n30700), .B(n30701), .Z(n30688) );
  AND U30484 ( .A(n30702), .B(n30703), .Z(n30701) );
  XOR U30485 ( .A(n30700), .B(n30330), .Z(n30703) );
  XOR U30486 ( .A(n30704), .B(n30705), .Z(n30330) );
  AND U30487 ( .A(n1099), .B(n30706), .Z(n30705) );
  XOR U30488 ( .A(n30707), .B(n30704), .Z(n30706) );
  XNOR U30489 ( .A(n30327), .B(n30700), .Z(n30702) );
  XOR U30490 ( .A(n30708), .B(n30709), .Z(n30327) );
  AND U30491 ( .A(n1097), .B(n30710), .Z(n30709) );
  XOR U30492 ( .A(n30711), .B(n30708), .Z(n30710) );
  XOR U30493 ( .A(n30712), .B(n30713), .Z(n30700) );
  AND U30494 ( .A(n30714), .B(n30715), .Z(n30713) );
  XOR U30495 ( .A(n30712), .B(n30342), .Z(n30715) );
  XOR U30496 ( .A(n30716), .B(n30717), .Z(n30342) );
  AND U30497 ( .A(n1099), .B(n30718), .Z(n30717) );
  XOR U30498 ( .A(n30719), .B(n30716), .Z(n30718) );
  XNOR U30499 ( .A(n30339), .B(n30712), .Z(n30714) );
  XOR U30500 ( .A(n30720), .B(n30721), .Z(n30339) );
  AND U30501 ( .A(n1097), .B(n30722), .Z(n30721) );
  XOR U30502 ( .A(n30723), .B(n30720), .Z(n30722) );
  XOR U30503 ( .A(n30724), .B(n30725), .Z(n30712) );
  AND U30504 ( .A(n30726), .B(n30727), .Z(n30725) );
  XOR U30505 ( .A(n30724), .B(n30354), .Z(n30727) );
  XOR U30506 ( .A(n30728), .B(n30729), .Z(n30354) );
  AND U30507 ( .A(n1099), .B(n30730), .Z(n30729) );
  XOR U30508 ( .A(n30731), .B(n30728), .Z(n30730) );
  XNOR U30509 ( .A(n30351), .B(n30724), .Z(n30726) );
  XOR U30510 ( .A(n30732), .B(n30733), .Z(n30351) );
  AND U30511 ( .A(n1097), .B(n30734), .Z(n30733) );
  XOR U30512 ( .A(n30735), .B(n30732), .Z(n30734) );
  XOR U30513 ( .A(n30736), .B(n30737), .Z(n30724) );
  AND U30514 ( .A(n30738), .B(n30739), .Z(n30737) );
  XOR U30515 ( .A(n30736), .B(n30366), .Z(n30739) );
  XOR U30516 ( .A(n30740), .B(n30741), .Z(n30366) );
  AND U30517 ( .A(n1099), .B(n30742), .Z(n30741) );
  XOR U30518 ( .A(n30743), .B(n30740), .Z(n30742) );
  XNOR U30519 ( .A(n30363), .B(n30736), .Z(n30738) );
  XOR U30520 ( .A(n30744), .B(n30745), .Z(n30363) );
  AND U30521 ( .A(n1097), .B(n30746), .Z(n30745) );
  XOR U30522 ( .A(n30747), .B(n30744), .Z(n30746) );
  XOR U30523 ( .A(n30748), .B(n30749), .Z(n30736) );
  AND U30524 ( .A(n30750), .B(n30751), .Z(n30749) );
  XOR U30525 ( .A(n30748), .B(n30378), .Z(n30751) );
  XOR U30526 ( .A(n30752), .B(n30753), .Z(n30378) );
  AND U30527 ( .A(n1099), .B(n30754), .Z(n30753) );
  XOR U30528 ( .A(n30755), .B(n30752), .Z(n30754) );
  XNOR U30529 ( .A(n30375), .B(n30748), .Z(n30750) );
  XOR U30530 ( .A(n30756), .B(n30757), .Z(n30375) );
  AND U30531 ( .A(n1097), .B(n30758), .Z(n30757) );
  XOR U30532 ( .A(n30759), .B(n30756), .Z(n30758) );
  XOR U30533 ( .A(n30760), .B(n30761), .Z(n30748) );
  AND U30534 ( .A(n30762), .B(n30763), .Z(n30761) );
  XOR U30535 ( .A(n30760), .B(n30390), .Z(n30763) );
  XOR U30536 ( .A(n30764), .B(n30765), .Z(n30390) );
  AND U30537 ( .A(n1099), .B(n30766), .Z(n30765) );
  XOR U30538 ( .A(n30767), .B(n30764), .Z(n30766) );
  XNOR U30539 ( .A(n30387), .B(n30760), .Z(n30762) );
  XOR U30540 ( .A(n30768), .B(n30769), .Z(n30387) );
  AND U30541 ( .A(n1097), .B(n30770), .Z(n30769) );
  XOR U30542 ( .A(n30771), .B(n30768), .Z(n30770) );
  XOR U30543 ( .A(n30772), .B(n30773), .Z(n30760) );
  AND U30544 ( .A(n30774), .B(n30775), .Z(n30773) );
  XOR U30545 ( .A(n30772), .B(n30402), .Z(n30775) );
  XOR U30546 ( .A(n30776), .B(n30777), .Z(n30402) );
  AND U30547 ( .A(n1099), .B(n30778), .Z(n30777) );
  XOR U30548 ( .A(n30779), .B(n30776), .Z(n30778) );
  XNOR U30549 ( .A(n30399), .B(n30772), .Z(n30774) );
  XOR U30550 ( .A(n30780), .B(n30781), .Z(n30399) );
  AND U30551 ( .A(n1097), .B(n30782), .Z(n30781) );
  XOR U30552 ( .A(n30783), .B(n30780), .Z(n30782) );
  XOR U30553 ( .A(n30784), .B(n30785), .Z(n30772) );
  AND U30554 ( .A(n30786), .B(n30787), .Z(n30785) );
  XOR U30555 ( .A(n30784), .B(n30414), .Z(n30787) );
  XOR U30556 ( .A(n30788), .B(n30789), .Z(n30414) );
  AND U30557 ( .A(n1099), .B(n30790), .Z(n30789) );
  XOR U30558 ( .A(n30791), .B(n30788), .Z(n30790) );
  XNOR U30559 ( .A(n30411), .B(n30784), .Z(n30786) );
  XOR U30560 ( .A(n30792), .B(n30793), .Z(n30411) );
  AND U30561 ( .A(n1097), .B(n30794), .Z(n30793) );
  XOR U30562 ( .A(n30795), .B(n30792), .Z(n30794) );
  XOR U30563 ( .A(n30796), .B(n30797), .Z(n30784) );
  AND U30564 ( .A(n30798), .B(n30799), .Z(n30797) );
  XOR U30565 ( .A(n30796), .B(n30426), .Z(n30799) );
  XOR U30566 ( .A(n30800), .B(n30801), .Z(n30426) );
  AND U30567 ( .A(n1099), .B(n30802), .Z(n30801) );
  XOR U30568 ( .A(n30803), .B(n30800), .Z(n30802) );
  XNOR U30569 ( .A(n30423), .B(n30796), .Z(n30798) );
  XOR U30570 ( .A(n30804), .B(n30805), .Z(n30423) );
  AND U30571 ( .A(n1097), .B(n30806), .Z(n30805) );
  XOR U30572 ( .A(n30807), .B(n30804), .Z(n30806) );
  XOR U30573 ( .A(n30808), .B(n30809), .Z(n30796) );
  AND U30574 ( .A(n30810), .B(n30811), .Z(n30809) );
  XOR U30575 ( .A(n30808), .B(n30438), .Z(n30811) );
  XOR U30576 ( .A(n30812), .B(n30813), .Z(n30438) );
  AND U30577 ( .A(n1099), .B(n30814), .Z(n30813) );
  XOR U30578 ( .A(n30815), .B(n30812), .Z(n30814) );
  XNOR U30579 ( .A(n30435), .B(n30808), .Z(n30810) );
  XOR U30580 ( .A(n30816), .B(n30817), .Z(n30435) );
  AND U30581 ( .A(n1097), .B(n30818), .Z(n30817) );
  XOR U30582 ( .A(n30819), .B(n30816), .Z(n30818) );
  XOR U30583 ( .A(n30820), .B(n30821), .Z(n30808) );
  AND U30584 ( .A(n30822), .B(n30823), .Z(n30821) );
  XOR U30585 ( .A(n30820), .B(n30450), .Z(n30823) );
  XOR U30586 ( .A(n30824), .B(n30825), .Z(n30450) );
  AND U30587 ( .A(n1099), .B(n30826), .Z(n30825) );
  XOR U30588 ( .A(n30827), .B(n30824), .Z(n30826) );
  XNOR U30589 ( .A(n30447), .B(n30820), .Z(n30822) );
  XOR U30590 ( .A(n30828), .B(n30829), .Z(n30447) );
  AND U30591 ( .A(n1097), .B(n30830), .Z(n30829) );
  XOR U30592 ( .A(n30831), .B(n30828), .Z(n30830) );
  XOR U30593 ( .A(n30832), .B(n30833), .Z(n30820) );
  AND U30594 ( .A(n30834), .B(n30835), .Z(n30833) );
  XOR U30595 ( .A(n30832), .B(n30462), .Z(n30835) );
  XOR U30596 ( .A(n30836), .B(n30837), .Z(n30462) );
  AND U30597 ( .A(n1099), .B(n30838), .Z(n30837) );
  XOR U30598 ( .A(n30839), .B(n30836), .Z(n30838) );
  XNOR U30599 ( .A(n30459), .B(n30832), .Z(n30834) );
  XOR U30600 ( .A(n30840), .B(n30841), .Z(n30459) );
  AND U30601 ( .A(n1097), .B(n30842), .Z(n30841) );
  XOR U30602 ( .A(n30843), .B(n30840), .Z(n30842) );
  XOR U30603 ( .A(n30844), .B(n30845), .Z(n30832) );
  AND U30604 ( .A(n30846), .B(n30847), .Z(n30845) );
  XOR U30605 ( .A(n30844), .B(n30474), .Z(n30847) );
  XOR U30606 ( .A(n30848), .B(n30849), .Z(n30474) );
  AND U30607 ( .A(n1099), .B(n30850), .Z(n30849) );
  XOR U30608 ( .A(n30851), .B(n30848), .Z(n30850) );
  XNOR U30609 ( .A(n30471), .B(n30844), .Z(n30846) );
  XOR U30610 ( .A(n30852), .B(n30853), .Z(n30471) );
  AND U30611 ( .A(n1097), .B(n30854), .Z(n30853) );
  XOR U30612 ( .A(n30855), .B(n30852), .Z(n30854) );
  XOR U30613 ( .A(n30856), .B(n30857), .Z(n30844) );
  AND U30614 ( .A(n30858), .B(n30859), .Z(n30857) );
  XOR U30615 ( .A(n30856), .B(n30486), .Z(n30859) );
  XOR U30616 ( .A(n30860), .B(n30861), .Z(n30486) );
  AND U30617 ( .A(n1099), .B(n30862), .Z(n30861) );
  XOR U30618 ( .A(n30863), .B(n30860), .Z(n30862) );
  XNOR U30619 ( .A(n30483), .B(n30856), .Z(n30858) );
  XOR U30620 ( .A(n30864), .B(n30865), .Z(n30483) );
  AND U30621 ( .A(n1097), .B(n30866), .Z(n30865) );
  XOR U30622 ( .A(n30867), .B(n30864), .Z(n30866) );
  XOR U30623 ( .A(n30868), .B(n30869), .Z(n30856) );
  AND U30624 ( .A(n30870), .B(n30871), .Z(n30869) );
  XOR U30625 ( .A(n30868), .B(n30498), .Z(n30871) );
  XOR U30626 ( .A(n30872), .B(n30873), .Z(n30498) );
  AND U30627 ( .A(n1099), .B(n30874), .Z(n30873) );
  XOR U30628 ( .A(n30875), .B(n30872), .Z(n30874) );
  XNOR U30629 ( .A(n30495), .B(n30868), .Z(n30870) );
  XOR U30630 ( .A(n30876), .B(n30877), .Z(n30495) );
  AND U30631 ( .A(n1097), .B(n30878), .Z(n30877) );
  XOR U30632 ( .A(n30879), .B(n30876), .Z(n30878) );
  XOR U30633 ( .A(n30880), .B(n30881), .Z(n30868) );
  AND U30634 ( .A(n30882), .B(n30883), .Z(n30881) );
  XOR U30635 ( .A(n30880), .B(n30510), .Z(n30883) );
  XOR U30636 ( .A(n30884), .B(n30885), .Z(n30510) );
  AND U30637 ( .A(n1099), .B(n30886), .Z(n30885) );
  XOR U30638 ( .A(n30887), .B(n30884), .Z(n30886) );
  XNOR U30639 ( .A(n30507), .B(n30880), .Z(n30882) );
  XOR U30640 ( .A(n30888), .B(n30889), .Z(n30507) );
  AND U30641 ( .A(n1097), .B(n30890), .Z(n30889) );
  XOR U30642 ( .A(n30891), .B(n30888), .Z(n30890) );
  XOR U30643 ( .A(n30892), .B(n30893), .Z(n30880) );
  AND U30644 ( .A(n30894), .B(n30895), .Z(n30893) );
  XOR U30645 ( .A(n30892), .B(n30522), .Z(n30895) );
  XOR U30646 ( .A(n30896), .B(n30897), .Z(n30522) );
  AND U30647 ( .A(n1099), .B(n30898), .Z(n30897) );
  XOR U30648 ( .A(n30899), .B(n30896), .Z(n30898) );
  XNOR U30649 ( .A(n30519), .B(n30892), .Z(n30894) );
  XOR U30650 ( .A(n30900), .B(n30901), .Z(n30519) );
  AND U30651 ( .A(n1097), .B(n30902), .Z(n30901) );
  XOR U30652 ( .A(n30903), .B(n30900), .Z(n30902) );
  XOR U30653 ( .A(n30904), .B(n30905), .Z(n30892) );
  AND U30654 ( .A(n30906), .B(n30907), .Z(n30905) );
  XOR U30655 ( .A(n30904), .B(n30534), .Z(n30907) );
  XOR U30656 ( .A(n30908), .B(n30909), .Z(n30534) );
  AND U30657 ( .A(n1099), .B(n30910), .Z(n30909) );
  XOR U30658 ( .A(n30911), .B(n30908), .Z(n30910) );
  XNOR U30659 ( .A(n30531), .B(n30904), .Z(n30906) );
  XOR U30660 ( .A(n30912), .B(n30913), .Z(n30531) );
  AND U30661 ( .A(n1097), .B(n30914), .Z(n30913) );
  XOR U30662 ( .A(n30915), .B(n30912), .Z(n30914) );
  XOR U30663 ( .A(n30916), .B(n30917), .Z(n30904) );
  AND U30664 ( .A(n30918), .B(n30919), .Z(n30917) );
  XOR U30665 ( .A(n30916), .B(n30546), .Z(n30919) );
  XOR U30666 ( .A(n30920), .B(n30921), .Z(n30546) );
  AND U30667 ( .A(n1099), .B(n30922), .Z(n30921) );
  XOR U30668 ( .A(n30923), .B(n30920), .Z(n30922) );
  XNOR U30669 ( .A(n30543), .B(n30916), .Z(n30918) );
  XOR U30670 ( .A(n30924), .B(n30925), .Z(n30543) );
  AND U30671 ( .A(n1097), .B(n30926), .Z(n30925) );
  XOR U30672 ( .A(n30927), .B(n30924), .Z(n30926) );
  XOR U30673 ( .A(n30928), .B(n30929), .Z(n30916) );
  AND U30674 ( .A(n30930), .B(n30931), .Z(n30929) );
  XOR U30675 ( .A(n30928), .B(n30558), .Z(n30931) );
  XOR U30676 ( .A(n30932), .B(n30933), .Z(n30558) );
  AND U30677 ( .A(n1099), .B(n30934), .Z(n30933) );
  XOR U30678 ( .A(n30935), .B(n30932), .Z(n30934) );
  XNOR U30679 ( .A(n30555), .B(n30928), .Z(n30930) );
  XOR U30680 ( .A(n30936), .B(n30937), .Z(n30555) );
  AND U30681 ( .A(n1097), .B(n30938), .Z(n30937) );
  XOR U30682 ( .A(n30939), .B(n30936), .Z(n30938) );
  XOR U30683 ( .A(n30940), .B(n30941), .Z(n30928) );
  AND U30684 ( .A(n30942), .B(n30943), .Z(n30941) );
  XOR U30685 ( .A(n30940), .B(n30570), .Z(n30943) );
  XOR U30686 ( .A(n30944), .B(n30945), .Z(n30570) );
  AND U30687 ( .A(n1099), .B(n30946), .Z(n30945) );
  XOR U30688 ( .A(n30947), .B(n30944), .Z(n30946) );
  XNOR U30689 ( .A(n30567), .B(n30940), .Z(n30942) );
  XOR U30690 ( .A(n30948), .B(n30949), .Z(n30567) );
  AND U30691 ( .A(n1097), .B(n30950), .Z(n30949) );
  XOR U30692 ( .A(n30951), .B(n30948), .Z(n30950) );
  XOR U30693 ( .A(n30952), .B(n30953), .Z(n30940) );
  AND U30694 ( .A(n30954), .B(n30955), .Z(n30953) );
  XOR U30695 ( .A(n30952), .B(n30582), .Z(n30955) );
  XOR U30696 ( .A(n30956), .B(n30957), .Z(n30582) );
  AND U30697 ( .A(n1099), .B(n30958), .Z(n30957) );
  XOR U30698 ( .A(n30959), .B(n30956), .Z(n30958) );
  XNOR U30699 ( .A(n30579), .B(n30952), .Z(n30954) );
  XOR U30700 ( .A(n30960), .B(n30961), .Z(n30579) );
  AND U30701 ( .A(n1097), .B(n30962), .Z(n30961) );
  XOR U30702 ( .A(n30963), .B(n30960), .Z(n30962) );
  XOR U30703 ( .A(n30964), .B(n30965), .Z(n30952) );
  AND U30704 ( .A(n30966), .B(n30967), .Z(n30965) );
  XOR U30705 ( .A(n30964), .B(n30594), .Z(n30967) );
  XOR U30706 ( .A(n30968), .B(n30969), .Z(n30594) );
  AND U30707 ( .A(n1099), .B(n30970), .Z(n30969) );
  XOR U30708 ( .A(n30971), .B(n30968), .Z(n30970) );
  XNOR U30709 ( .A(n30591), .B(n30964), .Z(n30966) );
  XOR U30710 ( .A(n30972), .B(n30973), .Z(n30591) );
  AND U30711 ( .A(n1097), .B(n30974), .Z(n30973) );
  XOR U30712 ( .A(n30975), .B(n30972), .Z(n30974) );
  XOR U30713 ( .A(n30976), .B(n30977), .Z(n30964) );
  AND U30714 ( .A(n30978), .B(n30979), .Z(n30977) );
  XOR U30715 ( .A(n30976), .B(n30606), .Z(n30979) );
  XOR U30716 ( .A(n30980), .B(n30981), .Z(n30606) );
  AND U30717 ( .A(n1099), .B(n30982), .Z(n30981) );
  XOR U30718 ( .A(n30983), .B(n30980), .Z(n30982) );
  XNOR U30719 ( .A(n30603), .B(n30976), .Z(n30978) );
  XOR U30720 ( .A(n30984), .B(n30985), .Z(n30603) );
  AND U30721 ( .A(n1097), .B(n30986), .Z(n30985) );
  XOR U30722 ( .A(n30987), .B(n30984), .Z(n30986) );
  XOR U30723 ( .A(n30988), .B(n30989), .Z(n30976) );
  AND U30724 ( .A(n30990), .B(n30991), .Z(n30989) );
  XOR U30725 ( .A(n30988), .B(n30618), .Z(n30991) );
  XOR U30726 ( .A(n30992), .B(n30993), .Z(n30618) );
  AND U30727 ( .A(n1099), .B(n30994), .Z(n30993) );
  XOR U30728 ( .A(n30995), .B(n30992), .Z(n30994) );
  XNOR U30729 ( .A(n30615), .B(n30988), .Z(n30990) );
  XOR U30730 ( .A(n30996), .B(n30997), .Z(n30615) );
  AND U30731 ( .A(n1097), .B(n30998), .Z(n30997) );
  XOR U30732 ( .A(n30999), .B(n30996), .Z(n30998) );
  XOR U30733 ( .A(n31000), .B(n31001), .Z(n30988) );
  AND U30734 ( .A(n31002), .B(n31003), .Z(n31001) );
  XOR U30735 ( .A(n31000), .B(n30630), .Z(n31003) );
  XOR U30736 ( .A(n31004), .B(n31005), .Z(n30630) );
  AND U30737 ( .A(n1099), .B(n31006), .Z(n31005) );
  XOR U30738 ( .A(n31007), .B(n31004), .Z(n31006) );
  XNOR U30739 ( .A(n30627), .B(n31000), .Z(n31002) );
  XOR U30740 ( .A(n31008), .B(n31009), .Z(n30627) );
  AND U30741 ( .A(n1097), .B(n31010), .Z(n31009) );
  XOR U30742 ( .A(n31011), .B(n31008), .Z(n31010) );
  XOR U30743 ( .A(n31012), .B(n31013), .Z(n31000) );
  AND U30744 ( .A(n31014), .B(n31015), .Z(n31013) );
  XOR U30745 ( .A(n31012), .B(n30642), .Z(n31015) );
  XOR U30746 ( .A(n31016), .B(n31017), .Z(n30642) );
  AND U30747 ( .A(n1099), .B(n31018), .Z(n31017) );
  XOR U30748 ( .A(n31019), .B(n31016), .Z(n31018) );
  XNOR U30749 ( .A(n30639), .B(n31012), .Z(n31014) );
  XOR U30750 ( .A(n31020), .B(n31021), .Z(n30639) );
  AND U30751 ( .A(n1097), .B(n31022), .Z(n31021) );
  XOR U30752 ( .A(n31023), .B(n31020), .Z(n31022) );
  XOR U30753 ( .A(n31024), .B(n31025), .Z(n31012) );
  AND U30754 ( .A(n31026), .B(n31027), .Z(n31025) );
  XOR U30755 ( .A(n31024), .B(n30654), .Z(n31027) );
  XOR U30756 ( .A(n31028), .B(n31029), .Z(n30654) );
  AND U30757 ( .A(n1099), .B(n31030), .Z(n31029) );
  XOR U30758 ( .A(n31031), .B(n31028), .Z(n31030) );
  XNOR U30759 ( .A(n30651), .B(n31024), .Z(n31026) );
  XOR U30760 ( .A(n31032), .B(n31033), .Z(n30651) );
  AND U30761 ( .A(n1097), .B(n31034), .Z(n31033) );
  XOR U30762 ( .A(n31035), .B(n31032), .Z(n31034) );
  XOR U30763 ( .A(n31036), .B(n31037), .Z(n31024) );
  AND U30764 ( .A(n31038), .B(n31039), .Z(n31037) );
  XNOR U30765 ( .A(n31040), .B(n30667), .Z(n31039) );
  XOR U30766 ( .A(n31041), .B(n31042), .Z(n30667) );
  AND U30767 ( .A(n1099), .B(n31043), .Z(n31042) );
  XOR U30768 ( .A(n31041), .B(n31044), .Z(n31043) );
  XNOR U30769 ( .A(n30664), .B(n31036), .Z(n31038) );
  XOR U30770 ( .A(n31045), .B(n31046), .Z(n30664) );
  AND U30771 ( .A(n1097), .B(n31047), .Z(n31046) );
  XOR U30772 ( .A(n31045), .B(n31048), .Z(n31047) );
  IV U30773 ( .A(n31040), .Z(n31036) );
  AND U30774 ( .A(n30672), .B(n30675), .Z(n31040) );
  XNOR U30775 ( .A(n31049), .B(n31050), .Z(n30675) );
  AND U30776 ( .A(n1099), .B(n31051), .Z(n31050) );
  XNOR U30777 ( .A(n31052), .B(n31049), .Z(n31051) );
  XOR U30778 ( .A(n31053), .B(n31054), .Z(n1099) );
  AND U30779 ( .A(n31055), .B(n31056), .Z(n31054) );
  XOR U30780 ( .A(n31053), .B(n30683), .Z(n31056) );
  XOR U30781 ( .A(n31057), .B(n31058), .Z(n30683) );
  AND U30782 ( .A(n1027), .B(n31059), .Z(n31058) );
  XOR U30783 ( .A(n31060), .B(n31057), .Z(n31059) );
  XNOR U30784 ( .A(n30680), .B(n31053), .Z(n31055) );
  XOR U30785 ( .A(n31061), .B(n31062), .Z(n30680) );
  AND U30786 ( .A(n1025), .B(n31063), .Z(n31062) );
  XOR U30787 ( .A(n31064), .B(n31061), .Z(n31063) );
  XOR U30788 ( .A(n31065), .B(n31066), .Z(n31053) );
  AND U30789 ( .A(n31067), .B(n31068), .Z(n31066) );
  XOR U30790 ( .A(n31065), .B(n30695), .Z(n31068) );
  XOR U30791 ( .A(n31069), .B(n31070), .Z(n30695) );
  AND U30792 ( .A(n1027), .B(n31071), .Z(n31070) );
  XOR U30793 ( .A(n31072), .B(n31069), .Z(n31071) );
  XNOR U30794 ( .A(n30692), .B(n31065), .Z(n31067) );
  XOR U30795 ( .A(n31073), .B(n31074), .Z(n30692) );
  AND U30796 ( .A(n1025), .B(n31075), .Z(n31074) );
  XOR U30797 ( .A(n31076), .B(n31073), .Z(n31075) );
  XOR U30798 ( .A(n31077), .B(n31078), .Z(n31065) );
  AND U30799 ( .A(n31079), .B(n31080), .Z(n31078) );
  XOR U30800 ( .A(n31077), .B(n30707), .Z(n31080) );
  XOR U30801 ( .A(n31081), .B(n31082), .Z(n30707) );
  AND U30802 ( .A(n1027), .B(n31083), .Z(n31082) );
  XOR U30803 ( .A(n31084), .B(n31081), .Z(n31083) );
  XNOR U30804 ( .A(n30704), .B(n31077), .Z(n31079) );
  XOR U30805 ( .A(n31085), .B(n31086), .Z(n30704) );
  AND U30806 ( .A(n1025), .B(n31087), .Z(n31086) );
  XOR U30807 ( .A(n31088), .B(n31085), .Z(n31087) );
  XOR U30808 ( .A(n31089), .B(n31090), .Z(n31077) );
  AND U30809 ( .A(n31091), .B(n31092), .Z(n31090) );
  XOR U30810 ( .A(n31089), .B(n30719), .Z(n31092) );
  XOR U30811 ( .A(n31093), .B(n31094), .Z(n30719) );
  AND U30812 ( .A(n1027), .B(n31095), .Z(n31094) );
  XOR U30813 ( .A(n31096), .B(n31093), .Z(n31095) );
  XNOR U30814 ( .A(n30716), .B(n31089), .Z(n31091) );
  XOR U30815 ( .A(n31097), .B(n31098), .Z(n30716) );
  AND U30816 ( .A(n1025), .B(n31099), .Z(n31098) );
  XOR U30817 ( .A(n31100), .B(n31097), .Z(n31099) );
  XOR U30818 ( .A(n31101), .B(n31102), .Z(n31089) );
  AND U30819 ( .A(n31103), .B(n31104), .Z(n31102) );
  XOR U30820 ( .A(n31101), .B(n30731), .Z(n31104) );
  XOR U30821 ( .A(n31105), .B(n31106), .Z(n30731) );
  AND U30822 ( .A(n1027), .B(n31107), .Z(n31106) );
  XOR U30823 ( .A(n31108), .B(n31105), .Z(n31107) );
  XNOR U30824 ( .A(n30728), .B(n31101), .Z(n31103) );
  XOR U30825 ( .A(n31109), .B(n31110), .Z(n30728) );
  AND U30826 ( .A(n1025), .B(n31111), .Z(n31110) );
  XOR U30827 ( .A(n31112), .B(n31109), .Z(n31111) );
  XOR U30828 ( .A(n31113), .B(n31114), .Z(n31101) );
  AND U30829 ( .A(n31115), .B(n31116), .Z(n31114) );
  XOR U30830 ( .A(n31113), .B(n30743), .Z(n31116) );
  XOR U30831 ( .A(n31117), .B(n31118), .Z(n30743) );
  AND U30832 ( .A(n1027), .B(n31119), .Z(n31118) );
  XOR U30833 ( .A(n31120), .B(n31117), .Z(n31119) );
  XNOR U30834 ( .A(n30740), .B(n31113), .Z(n31115) );
  XOR U30835 ( .A(n31121), .B(n31122), .Z(n30740) );
  AND U30836 ( .A(n1025), .B(n31123), .Z(n31122) );
  XOR U30837 ( .A(n31124), .B(n31121), .Z(n31123) );
  XOR U30838 ( .A(n31125), .B(n31126), .Z(n31113) );
  AND U30839 ( .A(n31127), .B(n31128), .Z(n31126) );
  XOR U30840 ( .A(n31125), .B(n30755), .Z(n31128) );
  XOR U30841 ( .A(n31129), .B(n31130), .Z(n30755) );
  AND U30842 ( .A(n1027), .B(n31131), .Z(n31130) );
  XOR U30843 ( .A(n31132), .B(n31129), .Z(n31131) );
  XNOR U30844 ( .A(n30752), .B(n31125), .Z(n31127) );
  XOR U30845 ( .A(n31133), .B(n31134), .Z(n30752) );
  AND U30846 ( .A(n1025), .B(n31135), .Z(n31134) );
  XOR U30847 ( .A(n31136), .B(n31133), .Z(n31135) );
  XOR U30848 ( .A(n31137), .B(n31138), .Z(n31125) );
  AND U30849 ( .A(n31139), .B(n31140), .Z(n31138) );
  XOR U30850 ( .A(n31137), .B(n30767), .Z(n31140) );
  XOR U30851 ( .A(n31141), .B(n31142), .Z(n30767) );
  AND U30852 ( .A(n1027), .B(n31143), .Z(n31142) );
  XOR U30853 ( .A(n31144), .B(n31141), .Z(n31143) );
  XNOR U30854 ( .A(n30764), .B(n31137), .Z(n31139) );
  XOR U30855 ( .A(n31145), .B(n31146), .Z(n30764) );
  AND U30856 ( .A(n1025), .B(n31147), .Z(n31146) );
  XOR U30857 ( .A(n31148), .B(n31145), .Z(n31147) );
  XOR U30858 ( .A(n31149), .B(n31150), .Z(n31137) );
  AND U30859 ( .A(n31151), .B(n31152), .Z(n31150) );
  XOR U30860 ( .A(n31149), .B(n30779), .Z(n31152) );
  XOR U30861 ( .A(n31153), .B(n31154), .Z(n30779) );
  AND U30862 ( .A(n1027), .B(n31155), .Z(n31154) );
  XOR U30863 ( .A(n31156), .B(n31153), .Z(n31155) );
  XNOR U30864 ( .A(n30776), .B(n31149), .Z(n31151) );
  XOR U30865 ( .A(n31157), .B(n31158), .Z(n30776) );
  AND U30866 ( .A(n1025), .B(n31159), .Z(n31158) );
  XOR U30867 ( .A(n31160), .B(n31157), .Z(n31159) );
  XOR U30868 ( .A(n31161), .B(n31162), .Z(n31149) );
  AND U30869 ( .A(n31163), .B(n31164), .Z(n31162) );
  XOR U30870 ( .A(n31161), .B(n30791), .Z(n31164) );
  XOR U30871 ( .A(n31165), .B(n31166), .Z(n30791) );
  AND U30872 ( .A(n1027), .B(n31167), .Z(n31166) );
  XOR U30873 ( .A(n31168), .B(n31165), .Z(n31167) );
  XNOR U30874 ( .A(n30788), .B(n31161), .Z(n31163) );
  XOR U30875 ( .A(n31169), .B(n31170), .Z(n30788) );
  AND U30876 ( .A(n1025), .B(n31171), .Z(n31170) );
  XOR U30877 ( .A(n31172), .B(n31169), .Z(n31171) );
  XOR U30878 ( .A(n31173), .B(n31174), .Z(n31161) );
  AND U30879 ( .A(n31175), .B(n31176), .Z(n31174) );
  XOR U30880 ( .A(n31173), .B(n30803), .Z(n31176) );
  XOR U30881 ( .A(n31177), .B(n31178), .Z(n30803) );
  AND U30882 ( .A(n1027), .B(n31179), .Z(n31178) );
  XOR U30883 ( .A(n31180), .B(n31177), .Z(n31179) );
  XNOR U30884 ( .A(n30800), .B(n31173), .Z(n31175) );
  XOR U30885 ( .A(n31181), .B(n31182), .Z(n30800) );
  AND U30886 ( .A(n1025), .B(n31183), .Z(n31182) );
  XOR U30887 ( .A(n31184), .B(n31181), .Z(n31183) );
  XOR U30888 ( .A(n31185), .B(n31186), .Z(n31173) );
  AND U30889 ( .A(n31187), .B(n31188), .Z(n31186) );
  XOR U30890 ( .A(n31185), .B(n30815), .Z(n31188) );
  XOR U30891 ( .A(n31189), .B(n31190), .Z(n30815) );
  AND U30892 ( .A(n1027), .B(n31191), .Z(n31190) );
  XOR U30893 ( .A(n31192), .B(n31189), .Z(n31191) );
  XNOR U30894 ( .A(n30812), .B(n31185), .Z(n31187) );
  XOR U30895 ( .A(n31193), .B(n31194), .Z(n30812) );
  AND U30896 ( .A(n1025), .B(n31195), .Z(n31194) );
  XOR U30897 ( .A(n31196), .B(n31193), .Z(n31195) );
  XOR U30898 ( .A(n31197), .B(n31198), .Z(n31185) );
  AND U30899 ( .A(n31199), .B(n31200), .Z(n31198) );
  XOR U30900 ( .A(n31197), .B(n30827), .Z(n31200) );
  XOR U30901 ( .A(n31201), .B(n31202), .Z(n30827) );
  AND U30902 ( .A(n1027), .B(n31203), .Z(n31202) );
  XOR U30903 ( .A(n31204), .B(n31201), .Z(n31203) );
  XNOR U30904 ( .A(n30824), .B(n31197), .Z(n31199) );
  XOR U30905 ( .A(n31205), .B(n31206), .Z(n30824) );
  AND U30906 ( .A(n1025), .B(n31207), .Z(n31206) );
  XOR U30907 ( .A(n31208), .B(n31205), .Z(n31207) );
  XOR U30908 ( .A(n31209), .B(n31210), .Z(n31197) );
  AND U30909 ( .A(n31211), .B(n31212), .Z(n31210) );
  XOR U30910 ( .A(n31209), .B(n30839), .Z(n31212) );
  XOR U30911 ( .A(n31213), .B(n31214), .Z(n30839) );
  AND U30912 ( .A(n1027), .B(n31215), .Z(n31214) );
  XOR U30913 ( .A(n31216), .B(n31213), .Z(n31215) );
  XNOR U30914 ( .A(n30836), .B(n31209), .Z(n31211) );
  XOR U30915 ( .A(n31217), .B(n31218), .Z(n30836) );
  AND U30916 ( .A(n1025), .B(n31219), .Z(n31218) );
  XOR U30917 ( .A(n31220), .B(n31217), .Z(n31219) );
  XOR U30918 ( .A(n31221), .B(n31222), .Z(n31209) );
  AND U30919 ( .A(n31223), .B(n31224), .Z(n31222) );
  XOR U30920 ( .A(n31221), .B(n30851), .Z(n31224) );
  XOR U30921 ( .A(n31225), .B(n31226), .Z(n30851) );
  AND U30922 ( .A(n1027), .B(n31227), .Z(n31226) );
  XOR U30923 ( .A(n31228), .B(n31225), .Z(n31227) );
  XNOR U30924 ( .A(n30848), .B(n31221), .Z(n31223) );
  XOR U30925 ( .A(n31229), .B(n31230), .Z(n30848) );
  AND U30926 ( .A(n1025), .B(n31231), .Z(n31230) );
  XOR U30927 ( .A(n31232), .B(n31229), .Z(n31231) );
  XOR U30928 ( .A(n31233), .B(n31234), .Z(n31221) );
  AND U30929 ( .A(n31235), .B(n31236), .Z(n31234) );
  XOR U30930 ( .A(n31233), .B(n30863), .Z(n31236) );
  XOR U30931 ( .A(n31237), .B(n31238), .Z(n30863) );
  AND U30932 ( .A(n1027), .B(n31239), .Z(n31238) );
  XOR U30933 ( .A(n31240), .B(n31237), .Z(n31239) );
  XNOR U30934 ( .A(n30860), .B(n31233), .Z(n31235) );
  XOR U30935 ( .A(n31241), .B(n31242), .Z(n30860) );
  AND U30936 ( .A(n1025), .B(n31243), .Z(n31242) );
  XOR U30937 ( .A(n31244), .B(n31241), .Z(n31243) );
  XOR U30938 ( .A(n31245), .B(n31246), .Z(n31233) );
  AND U30939 ( .A(n31247), .B(n31248), .Z(n31246) );
  XOR U30940 ( .A(n31245), .B(n30875), .Z(n31248) );
  XOR U30941 ( .A(n31249), .B(n31250), .Z(n30875) );
  AND U30942 ( .A(n1027), .B(n31251), .Z(n31250) );
  XOR U30943 ( .A(n31252), .B(n31249), .Z(n31251) );
  XNOR U30944 ( .A(n30872), .B(n31245), .Z(n31247) );
  XOR U30945 ( .A(n31253), .B(n31254), .Z(n30872) );
  AND U30946 ( .A(n1025), .B(n31255), .Z(n31254) );
  XOR U30947 ( .A(n31256), .B(n31253), .Z(n31255) );
  XOR U30948 ( .A(n31257), .B(n31258), .Z(n31245) );
  AND U30949 ( .A(n31259), .B(n31260), .Z(n31258) );
  XOR U30950 ( .A(n31257), .B(n30887), .Z(n31260) );
  XOR U30951 ( .A(n31261), .B(n31262), .Z(n30887) );
  AND U30952 ( .A(n1027), .B(n31263), .Z(n31262) );
  XOR U30953 ( .A(n31264), .B(n31261), .Z(n31263) );
  XNOR U30954 ( .A(n30884), .B(n31257), .Z(n31259) );
  XOR U30955 ( .A(n31265), .B(n31266), .Z(n30884) );
  AND U30956 ( .A(n1025), .B(n31267), .Z(n31266) );
  XOR U30957 ( .A(n31268), .B(n31265), .Z(n31267) );
  XOR U30958 ( .A(n31269), .B(n31270), .Z(n31257) );
  AND U30959 ( .A(n31271), .B(n31272), .Z(n31270) );
  XOR U30960 ( .A(n31269), .B(n30899), .Z(n31272) );
  XOR U30961 ( .A(n31273), .B(n31274), .Z(n30899) );
  AND U30962 ( .A(n1027), .B(n31275), .Z(n31274) );
  XOR U30963 ( .A(n31276), .B(n31273), .Z(n31275) );
  XNOR U30964 ( .A(n30896), .B(n31269), .Z(n31271) );
  XOR U30965 ( .A(n31277), .B(n31278), .Z(n30896) );
  AND U30966 ( .A(n1025), .B(n31279), .Z(n31278) );
  XOR U30967 ( .A(n31280), .B(n31277), .Z(n31279) );
  XOR U30968 ( .A(n31281), .B(n31282), .Z(n31269) );
  AND U30969 ( .A(n31283), .B(n31284), .Z(n31282) );
  XOR U30970 ( .A(n31281), .B(n30911), .Z(n31284) );
  XOR U30971 ( .A(n31285), .B(n31286), .Z(n30911) );
  AND U30972 ( .A(n1027), .B(n31287), .Z(n31286) );
  XOR U30973 ( .A(n31288), .B(n31285), .Z(n31287) );
  XNOR U30974 ( .A(n30908), .B(n31281), .Z(n31283) );
  XOR U30975 ( .A(n31289), .B(n31290), .Z(n30908) );
  AND U30976 ( .A(n1025), .B(n31291), .Z(n31290) );
  XOR U30977 ( .A(n31292), .B(n31289), .Z(n31291) );
  XOR U30978 ( .A(n31293), .B(n31294), .Z(n31281) );
  AND U30979 ( .A(n31295), .B(n31296), .Z(n31294) );
  XOR U30980 ( .A(n31293), .B(n30923), .Z(n31296) );
  XOR U30981 ( .A(n31297), .B(n31298), .Z(n30923) );
  AND U30982 ( .A(n1027), .B(n31299), .Z(n31298) );
  XOR U30983 ( .A(n31300), .B(n31297), .Z(n31299) );
  XNOR U30984 ( .A(n30920), .B(n31293), .Z(n31295) );
  XOR U30985 ( .A(n31301), .B(n31302), .Z(n30920) );
  AND U30986 ( .A(n1025), .B(n31303), .Z(n31302) );
  XOR U30987 ( .A(n31304), .B(n31301), .Z(n31303) );
  XOR U30988 ( .A(n31305), .B(n31306), .Z(n31293) );
  AND U30989 ( .A(n31307), .B(n31308), .Z(n31306) );
  XOR U30990 ( .A(n31305), .B(n30935), .Z(n31308) );
  XOR U30991 ( .A(n31309), .B(n31310), .Z(n30935) );
  AND U30992 ( .A(n1027), .B(n31311), .Z(n31310) );
  XOR U30993 ( .A(n31312), .B(n31309), .Z(n31311) );
  XNOR U30994 ( .A(n30932), .B(n31305), .Z(n31307) );
  XOR U30995 ( .A(n31313), .B(n31314), .Z(n30932) );
  AND U30996 ( .A(n1025), .B(n31315), .Z(n31314) );
  XOR U30997 ( .A(n31316), .B(n31313), .Z(n31315) );
  XOR U30998 ( .A(n31317), .B(n31318), .Z(n31305) );
  AND U30999 ( .A(n31319), .B(n31320), .Z(n31318) );
  XOR U31000 ( .A(n31317), .B(n30947), .Z(n31320) );
  XOR U31001 ( .A(n31321), .B(n31322), .Z(n30947) );
  AND U31002 ( .A(n1027), .B(n31323), .Z(n31322) );
  XOR U31003 ( .A(n31324), .B(n31321), .Z(n31323) );
  XNOR U31004 ( .A(n30944), .B(n31317), .Z(n31319) );
  XOR U31005 ( .A(n31325), .B(n31326), .Z(n30944) );
  AND U31006 ( .A(n1025), .B(n31327), .Z(n31326) );
  XOR U31007 ( .A(n31328), .B(n31325), .Z(n31327) );
  XOR U31008 ( .A(n31329), .B(n31330), .Z(n31317) );
  AND U31009 ( .A(n31331), .B(n31332), .Z(n31330) );
  XOR U31010 ( .A(n31329), .B(n30959), .Z(n31332) );
  XOR U31011 ( .A(n31333), .B(n31334), .Z(n30959) );
  AND U31012 ( .A(n1027), .B(n31335), .Z(n31334) );
  XOR U31013 ( .A(n31336), .B(n31333), .Z(n31335) );
  XNOR U31014 ( .A(n30956), .B(n31329), .Z(n31331) );
  XOR U31015 ( .A(n31337), .B(n31338), .Z(n30956) );
  AND U31016 ( .A(n1025), .B(n31339), .Z(n31338) );
  XOR U31017 ( .A(n31340), .B(n31337), .Z(n31339) );
  XOR U31018 ( .A(n31341), .B(n31342), .Z(n31329) );
  AND U31019 ( .A(n31343), .B(n31344), .Z(n31342) );
  XOR U31020 ( .A(n31341), .B(n30971), .Z(n31344) );
  XOR U31021 ( .A(n31345), .B(n31346), .Z(n30971) );
  AND U31022 ( .A(n1027), .B(n31347), .Z(n31346) );
  XOR U31023 ( .A(n31348), .B(n31345), .Z(n31347) );
  XNOR U31024 ( .A(n30968), .B(n31341), .Z(n31343) );
  XOR U31025 ( .A(n31349), .B(n31350), .Z(n30968) );
  AND U31026 ( .A(n1025), .B(n31351), .Z(n31350) );
  XOR U31027 ( .A(n31352), .B(n31349), .Z(n31351) );
  XOR U31028 ( .A(n31353), .B(n31354), .Z(n31341) );
  AND U31029 ( .A(n31355), .B(n31356), .Z(n31354) );
  XOR U31030 ( .A(n31353), .B(n30983), .Z(n31356) );
  XOR U31031 ( .A(n31357), .B(n31358), .Z(n30983) );
  AND U31032 ( .A(n1027), .B(n31359), .Z(n31358) );
  XOR U31033 ( .A(n31360), .B(n31357), .Z(n31359) );
  XNOR U31034 ( .A(n30980), .B(n31353), .Z(n31355) );
  XOR U31035 ( .A(n31361), .B(n31362), .Z(n30980) );
  AND U31036 ( .A(n1025), .B(n31363), .Z(n31362) );
  XOR U31037 ( .A(n31364), .B(n31361), .Z(n31363) );
  XOR U31038 ( .A(n31365), .B(n31366), .Z(n31353) );
  AND U31039 ( .A(n31367), .B(n31368), .Z(n31366) );
  XOR U31040 ( .A(n31365), .B(n30995), .Z(n31368) );
  XOR U31041 ( .A(n31369), .B(n31370), .Z(n30995) );
  AND U31042 ( .A(n1027), .B(n31371), .Z(n31370) );
  XOR U31043 ( .A(n31372), .B(n31369), .Z(n31371) );
  XNOR U31044 ( .A(n30992), .B(n31365), .Z(n31367) );
  XOR U31045 ( .A(n31373), .B(n31374), .Z(n30992) );
  AND U31046 ( .A(n1025), .B(n31375), .Z(n31374) );
  XOR U31047 ( .A(n31376), .B(n31373), .Z(n31375) );
  XOR U31048 ( .A(n31377), .B(n31378), .Z(n31365) );
  AND U31049 ( .A(n31379), .B(n31380), .Z(n31378) );
  XOR U31050 ( .A(n31377), .B(n31007), .Z(n31380) );
  XOR U31051 ( .A(n31381), .B(n31382), .Z(n31007) );
  AND U31052 ( .A(n1027), .B(n31383), .Z(n31382) );
  XOR U31053 ( .A(n31384), .B(n31381), .Z(n31383) );
  XNOR U31054 ( .A(n31004), .B(n31377), .Z(n31379) );
  XOR U31055 ( .A(n31385), .B(n31386), .Z(n31004) );
  AND U31056 ( .A(n1025), .B(n31387), .Z(n31386) );
  XOR U31057 ( .A(n31388), .B(n31385), .Z(n31387) );
  XOR U31058 ( .A(n31389), .B(n31390), .Z(n31377) );
  AND U31059 ( .A(n31391), .B(n31392), .Z(n31390) );
  XOR U31060 ( .A(n31389), .B(n31019), .Z(n31392) );
  XOR U31061 ( .A(n31393), .B(n31394), .Z(n31019) );
  AND U31062 ( .A(n1027), .B(n31395), .Z(n31394) );
  XOR U31063 ( .A(n31396), .B(n31393), .Z(n31395) );
  XNOR U31064 ( .A(n31016), .B(n31389), .Z(n31391) );
  XOR U31065 ( .A(n31397), .B(n31398), .Z(n31016) );
  AND U31066 ( .A(n1025), .B(n31399), .Z(n31398) );
  XOR U31067 ( .A(n31400), .B(n31397), .Z(n31399) );
  XOR U31068 ( .A(n31401), .B(n31402), .Z(n31389) );
  AND U31069 ( .A(n31403), .B(n31404), .Z(n31402) );
  XOR U31070 ( .A(n31401), .B(n31031), .Z(n31404) );
  XOR U31071 ( .A(n31405), .B(n31406), .Z(n31031) );
  AND U31072 ( .A(n1027), .B(n31407), .Z(n31406) );
  XOR U31073 ( .A(n31408), .B(n31405), .Z(n31407) );
  XNOR U31074 ( .A(n31028), .B(n31401), .Z(n31403) );
  XOR U31075 ( .A(n31409), .B(n31410), .Z(n31028) );
  AND U31076 ( .A(n1025), .B(n31411), .Z(n31410) );
  XOR U31077 ( .A(n31412), .B(n31409), .Z(n31411) );
  XOR U31078 ( .A(n31413), .B(n31414), .Z(n31401) );
  AND U31079 ( .A(n31415), .B(n31416), .Z(n31414) );
  XNOR U31080 ( .A(n31417), .B(n31044), .Z(n31416) );
  XOR U31081 ( .A(n31418), .B(n31419), .Z(n31044) );
  AND U31082 ( .A(n1027), .B(n31420), .Z(n31419) );
  XOR U31083 ( .A(n31418), .B(n31421), .Z(n31420) );
  XNOR U31084 ( .A(n31041), .B(n31413), .Z(n31415) );
  XOR U31085 ( .A(n31422), .B(n31423), .Z(n31041) );
  AND U31086 ( .A(n1025), .B(n31424), .Z(n31423) );
  XOR U31087 ( .A(n31422), .B(n31425), .Z(n31424) );
  IV U31088 ( .A(n31417), .Z(n31413) );
  AND U31089 ( .A(n31049), .B(n31052), .Z(n31417) );
  XNOR U31090 ( .A(n31426), .B(n31427), .Z(n31052) );
  AND U31091 ( .A(n1027), .B(n31428), .Z(n31427) );
  XNOR U31092 ( .A(n31429), .B(n31426), .Z(n31428) );
  XOR U31093 ( .A(n31430), .B(n31431), .Z(n1027) );
  AND U31094 ( .A(n31432), .B(n31433), .Z(n31431) );
  XOR U31095 ( .A(n31430), .B(n31060), .Z(n31433) );
  XOR U31096 ( .A(n31434), .B(n31435), .Z(n31060) );
  AND U31097 ( .A(n875), .B(n31436), .Z(n31435) );
  XOR U31098 ( .A(n31437), .B(n31434), .Z(n31436) );
  XNOR U31099 ( .A(n31057), .B(n31430), .Z(n31432) );
  XOR U31100 ( .A(n31438), .B(n31439), .Z(n31057) );
  AND U31101 ( .A(n873), .B(n31440), .Z(n31439) );
  XOR U31102 ( .A(n31441), .B(n31438), .Z(n31440) );
  XOR U31103 ( .A(n31442), .B(n31443), .Z(n31430) );
  AND U31104 ( .A(n31444), .B(n31445), .Z(n31443) );
  XOR U31105 ( .A(n31442), .B(n31072), .Z(n31445) );
  XOR U31106 ( .A(n31446), .B(n31447), .Z(n31072) );
  AND U31107 ( .A(n875), .B(n31448), .Z(n31447) );
  XOR U31108 ( .A(n31449), .B(n31446), .Z(n31448) );
  XNOR U31109 ( .A(n31069), .B(n31442), .Z(n31444) );
  XOR U31110 ( .A(n31450), .B(n31451), .Z(n31069) );
  AND U31111 ( .A(n873), .B(n31452), .Z(n31451) );
  XOR U31112 ( .A(n31453), .B(n31450), .Z(n31452) );
  XOR U31113 ( .A(n31454), .B(n31455), .Z(n31442) );
  AND U31114 ( .A(n31456), .B(n31457), .Z(n31455) );
  XOR U31115 ( .A(n31454), .B(n31084), .Z(n31457) );
  XOR U31116 ( .A(n31458), .B(n31459), .Z(n31084) );
  AND U31117 ( .A(n875), .B(n31460), .Z(n31459) );
  XOR U31118 ( .A(n31461), .B(n31458), .Z(n31460) );
  XNOR U31119 ( .A(n31081), .B(n31454), .Z(n31456) );
  XOR U31120 ( .A(n31462), .B(n31463), .Z(n31081) );
  AND U31121 ( .A(n873), .B(n31464), .Z(n31463) );
  XOR U31122 ( .A(n31465), .B(n31462), .Z(n31464) );
  XOR U31123 ( .A(n31466), .B(n31467), .Z(n31454) );
  AND U31124 ( .A(n31468), .B(n31469), .Z(n31467) );
  XOR U31125 ( .A(n31466), .B(n31096), .Z(n31469) );
  XOR U31126 ( .A(n31470), .B(n31471), .Z(n31096) );
  AND U31127 ( .A(n875), .B(n31472), .Z(n31471) );
  XOR U31128 ( .A(n31473), .B(n31470), .Z(n31472) );
  XNOR U31129 ( .A(n31093), .B(n31466), .Z(n31468) );
  XOR U31130 ( .A(n31474), .B(n31475), .Z(n31093) );
  AND U31131 ( .A(n873), .B(n31476), .Z(n31475) );
  XOR U31132 ( .A(n31477), .B(n31474), .Z(n31476) );
  XOR U31133 ( .A(n31478), .B(n31479), .Z(n31466) );
  AND U31134 ( .A(n31480), .B(n31481), .Z(n31479) );
  XOR U31135 ( .A(n31478), .B(n31108), .Z(n31481) );
  XOR U31136 ( .A(n31482), .B(n31483), .Z(n31108) );
  AND U31137 ( .A(n875), .B(n31484), .Z(n31483) );
  XOR U31138 ( .A(n31485), .B(n31482), .Z(n31484) );
  XNOR U31139 ( .A(n31105), .B(n31478), .Z(n31480) );
  XOR U31140 ( .A(n31486), .B(n31487), .Z(n31105) );
  AND U31141 ( .A(n873), .B(n31488), .Z(n31487) );
  XOR U31142 ( .A(n31489), .B(n31486), .Z(n31488) );
  XOR U31143 ( .A(n31490), .B(n31491), .Z(n31478) );
  AND U31144 ( .A(n31492), .B(n31493), .Z(n31491) );
  XOR U31145 ( .A(n31490), .B(n31120), .Z(n31493) );
  XOR U31146 ( .A(n31494), .B(n31495), .Z(n31120) );
  AND U31147 ( .A(n875), .B(n31496), .Z(n31495) );
  XOR U31148 ( .A(n31497), .B(n31494), .Z(n31496) );
  XNOR U31149 ( .A(n31117), .B(n31490), .Z(n31492) );
  XOR U31150 ( .A(n31498), .B(n31499), .Z(n31117) );
  AND U31151 ( .A(n873), .B(n31500), .Z(n31499) );
  XOR U31152 ( .A(n31501), .B(n31498), .Z(n31500) );
  XOR U31153 ( .A(n31502), .B(n31503), .Z(n31490) );
  AND U31154 ( .A(n31504), .B(n31505), .Z(n31503) );
  XOR U31155 ( .A(n31502), .B(n31132), .Z(n31505) );
  XOR U31156 ( .A(n31506), .B(n31507), .Z(n31132) );
  AND U31157 ( .A(n875), .B(n31508), .Z(n31507) );
  XOR U31158 ( .A(n31509), .B(n31506), .Z(n31508) );
  XNOR U31159 ( .A(n31129), .B(n31502), .Z(n31504) );
  XOR U31160 ( .A(n31510), .B(n31511), .Z(n31129) );
  AND U31161 ( .A(n873), .B(n31512), .Z(n31511) );
  XOR U31162 ( .A(n31513), .B(n31510), .Z(n31512) );
  XOR U31163 ( .A(n31514), .B(n31515), .Z(n31502) );
  AND U31164 ( .A(n31516), .B(n31517), .Z(n31515) );
  XOR U31165 ( .A(n31514), .B(n31144), .Z(n31517) );
  XOR U31166 ( .A(n31518), .B(n31519), .Z(n31144) );
  AND U31167 ( .A(n875), .B(n31520), .Z(n31519) );
  XOR U31168 ( .A(n31521), .B(n31518), .Z(n31520) );
  XNOR U31169 ( .A(n31141), .B(n31514), .Z(n31516) );
  XOR U31170 ( .A(n31522), .B(n31523), .Z(n31141) );
  AND U31171 ( .A(n873), .B(n31524), .Z(n31523) );
  XOR U31172 ( .A(n31525), .B(n31522), .Z(n31524) );
  XOR U31173 ( .A(n31526), .B(n31527), .Z(n31514) );
  AND U31174 ( .A(n31528), .B(n31529), .Z(n31527) );
  XOR U31175 ( .A(n31526), .B(n31156), .Z(n31529) );
  XOR U31176 ( .A(n31530), .B(n31531), .Z(n31156) );
  AND U31177 ( .A(n875), .B(n31532), .Z(n31531) );
  XOR U31178 ( .A(n31533), .B(n31530), .Z(n31532) );
  XNOR U31179 ( .A(n31153), .B(n31526), .Z(n31528) );
  XOR U31180 ( .A(n31534), .B(n31535), .Z(n31153) );
  AND U31181 ( .A(n873), .B(n31536), .Z(n31535) );
  XOR U31182 ( .A(n31537), .B(n31534), .Z(n31536) );
  XOR U31183 ( .A(n31538), .B(n31539), .Z(n31526) );
  AND U31184 ( .A(n31540), .B(n31541), .Z(n31539) );
  XOR U31185 ( .A(n31538), .B(n31168), .Z(n31541) );
  XOR U31186 ( .A(n31542), .B(n31543), .Z(n31168) );
  AND U31187 ( .A(n875), .B(n31544), .Z(n31543) );
  XOR U31188 ( .A(n31545), .B(n31542), .Z(n31544) );
  XNOR U31189 ( .A(n31165), .B(n31538), .Z(n31540) );
  XOR U31190 ( .A(n31546), .B(n31547), .Z(n31165) );
  AND U31191 ( .A(n873), .B(n31548), .Z(n31547) );
  XOR U31192 ( .A(n31549), .B(n31546), .Z(n31548) );
  XOR U31193 ( .A(n31550), .B(n31551), .Z(n31538) );
  AND U31194 ( .A(n31552), .B(n31553), .Z(n31551) );
  XOR U31195 ( .A(n31550), .B(n31180), .Z(n31553) );
  XOR U31196 ( .A(n31554), .B(n31555), .Z(n31180) );
  AND U31197 ( .A(n875), .B(n31556), .Z(n31555) );
  XOR U31198 ( .A(n31557), .B(n31554), .Z(n31556) );
  XNOR U31199 ( .A(n31177), .B(n31550), .Z(n31552) );
  XOR U31200 ( .A(n31558), .B(n31559), .Z(n31177) );
  AND U31201 ( .A(n873), .B(n31560), .Z(n31559) );
  XOR U31202 ( .A(n31561), .B(n31558), .Z(n31560) );
  XOR U31203 ( .A(n31562), .B(n31563), .Z(n31550) );
  AND U31204 ( .A(n31564), .B(n31565), .Z(n31563) );
  XOR U31205 ( .A(n31562), .B(n31192), .Z(n31565) );
  XOR U31206 ( .A(n31566), .B(n31567), .Z(n31192) );
  AND U31207 ( .A(n875), .B(n31568), .Z(n31567) );
  XOR U31208 ( .A(n31569), .B(n31566), .Z(n31568) );
  XNOR U31209 ( .A(n31189), .B(n31562), .Z(n31564) );
  XOR U31210 ( .A(n31570), .B(n31571), .Z(n31189) );
  AND U31211 ( .A(n873), .B(n31572), .Z(n31571) );
  XOR U31212 ( .A(n31573), .B(n31570), .Z(n31572) );
  XOR U31213 ( .A(n31574), .B(n31575), .Z(n31562) );
  AND U31214 ( .A(n31576), .B(n31577), .Z(n31575) );
  XOR U31215 ( .A(n31574), .B(n31204), .Z(n31577) );
  XOR U31216 ( .A(n31578), .B(n31579), .Z(n31204) );
  AND U31217 ( .A(n875), .B(n31580), .Z(n31579) );
  XOR U31218 ( .A(n31581), .B(n31578), .Z(n31580) );
  XNOR U31219 ( .A(n31201), .B(n31574), .Z(n31576) );
  XOR U31220 ( .A(n31582), .B(n31583), .Z(n31201) );
  AND U31221 ( .A(n873), .B(n31584), .Z(n31583) );
  XOR U31222 ( .A(n31585), .B(n31582), .Z(n31584) );
  XOR U31223 ( .A(n31586), .B(n31587), .Z(n31574) );
  AND U31224 ( .A(n31588), .B(n31589), .Z(n31587) );
  XOR U31225 ( .A(n31586), .B(n31216), .Z(n31589) );
  XOR U31226 ( .A(n31590), .B(n31591), .Z(n31216) );
  AND U31227 ( .A(n875), .B(n31592), .Z(n31591) );
  XOR U31228 ( .A(n31593), .B(n31590), .Z(n31592) );
  XNOR U31229 ( .A(n31213), .B(n31586), .Z(n31588) );
  XOR U31230 ( .A(n31594), .B(n31595), .Z(n31213) );
  AND U31231 ( .A(n873), .B(n31596), .Z(n31595) );
  XOR U31232 ( .A(n31597), .B(n31594), .Z(n31596) );
  XOR U31233 ( .A(n31598), .B(n31599), .Z(n31586) );
  AND U31234 ( .A(n31600), .B(n31601), .Z(n31599) );
  XOR U31235 ( .A(n31598), .B(n31228), .Z(n31601) );
  XOR U31236 ( .A(n31602), .B(n31603), .Z(n31228) );
  AND U31237 ( .A(n875), .B(n31604), .Z(n31603) );
  XOR U31238 ( .A(n31605), .B(n31602), .Z(n31604) );
  XNOR U31239 ( .A(n31225), .B(n31598), .Z(n31600) );
  XOR U31240 ( .A(n31606), .B(n31607), .Z(n31225) );
  AND U31241 ( .A(n873), .B(n31608), .Z(n31607) );
  XOR U31242 ( .A(n31609), .B(n31606), .Z(n31608) );
  XOR U31243 ( .A(n31610), .B(n31611), .Z(n31598) );
  AND U31244 ( .A(n31612), .B(n31613), .Z(n31611) );
  XOR U31245 ( .A(n31610), .B(n31240), .Z(n31613) );
  XOR U31246 ( .A(n31614), .B(n31615), .Z(n31240) );
  AND U31247 ( .A(n875), .B(n31616), .Z(n31615) );
  XOR U31248 ( .A(n31617), .B(n31614), .Z(n31616) );
  XNOR U31249 ( .A(n31237), .B(n31610), .Z(n31612) );
  XOR U31250 ( .A(n31618), .B(n31619), .Z(n31237) );
  AND U31251 ( .A(n873), .B(n31620), .Z(n31619) );
  XOR U31252 ( .A(n31621), .B(n31618), .Z(n31620) );
  XOR U31253 ( .A(n31622), .B(n31623), .Z(n31610) );
  AND U31254 ( .A(n31624), .B(n31625), .Z(n31623) );
  XOR U31255 ( .A(n31622), .B(n31252), .Z(n31625) );
  XOR U31256 ( .A(n31626), .B(n31627), .Z(n31252) );
  AND U31257 ( .A(n875), .B(n31628), .Z(n31627) );
  XOR U31258 ( .A(n31629), .B(n31626), .Z(n31628) );
  XNOR U31259 ( .A(n31249), .B(n31622), .Z(n31624) );
  XOR U31260 ( .A(n31630), .B(n31631), .Z(n31249) );
  AND U31261 ( .A(n873), .B(n31632), .Z(n31631) );
  XOR U31262 ( .A(n31633), .B(n31630), .Z(n31632) );
  XOR U31263 ( .A(n31634), .B(n31635), .Z(n31622) );
  AND U31264 ( .A(n31636), .B(n31637), .Z(n31635) );
  XOR U31265 ( .A(n31634), .B(n31264), .Z(n31637) );
  XOR U31266 ( .A(n31638), .B(n31639), .Z(n31264) );
  AND U31267 ( .A(n875), .B(n31640), .Z(n31639) );
  XOR U31268 ( .A(n31641), .B(n31638), .Z(n31640) );
  XNOR U31269 ( .A(n31261), .B(n31634), .Z(n31636) );
  XOR U31270 ( .A(n31642), .B(n31643), .Z(n31261) );
  AND U31271 ( .A(n873), .B(n31644), .Z(n31643) );
  XOR U31272 ( .A(n31645), .B(n31642), .Z(n31644) );
  XOR U31273 ( .A(n31646), .B(n31647), .Z(n31634) );
  AND U31274 ( .A(n31648), .B(n31649), .Z(n31647) );
  XOR U31275 ( .A(n31646), .B(n31276), .Z(n31649) );
  XOR U31276 ( .A(n31650), .B(n31651), .Z(n31276) );
  AND U31277 ( .A(n875), .B(n31652), .Z(n31651) );
  XOR U31278 ( .A(n31653), .B(n31650), .Z(n31652) );
  XNOR U31279 ( .A(n31273), .B(n31646), .Z(n31648) );
  XOR U31280 ( .A(n31654), .B(n31655), .Z(n31273) );
  AND U31281 ( .A(n873), .B(n31656), .Z(n31655) );
  XOR U31282 ( .A(n31657), .B(n31654), .Z(n31656) );
  XOR U31283 ( .A(n31658), .B(n31659), .Z(n31646) );
  AND U31284 ( .A(n31660), .B(n31661), .Z(n31659) );
  XOR U31285 ( .A(n31658), .B(n31288), .Z(n31661) );
  XOR U31286 ( .A(n31662), .B(n31663), .Z(n31288) );
  AND U31287 ( .A(n875), .B(n31664), .Z(n31663) );
  XOR U31288 ( .A(n31665), .B(n31662), .Z(n31664) );
  XNOR U31289 ( .A(n31285), .B(n31658), .Z(n31660) );
  XOR U31290 ( .A(n31666), .B(n31667), .Z(n31285) );
  AND U31291 ( .A(n873), .B(n31668), .Z(n31667) );
  XOR U31292 ( .A(n31669), .B(n31666), .Z(n31668) );
  XOR U31293 ( .A(n31670), .B(n31671), .Z(n31658) );
  AND U31294 ( .A(n31672), .B(n31673), .Z(n31671) );
  XOR U31295 ( .A(n31670), .B(n31300), .Z(n31673) );
  XOR U31296 ( .A(n31674), .B(n31675), .Z(n31300) );
  AND U31297 ( .A(n875), .B(n31676), .Z(n31675) );
  XOR U31298 ( .A(n31677), .B(n31674), .Z(n31676) );
  XNOR U31299 ( .A(n31297), .B(n31670), .Z(n31672) );
  XOR U31300 ( .A(n31678), .B(n31679), .Z(n31297) );
  AND U31301 ( .A(n873), .B(n31680), .Z(n31679) );
  XOR U31302 ( .A(n31681), .B(n31678), .Z(n31680) );
  XOR U31303 ( .A(n31682), .B(n31683), .Z(n31670) );
  AND U31304 ( .A(n31684), .B(n31685), .Z(n31683) );
  XOR U31305 ( .A(n31682), .B(n31312), .Z(n31685) );
  XOR U31306 ( .A(n31686), .B(n31687), .Z(n31312) );
  AND U31307 ( .A(n875), .B(n31688), .Z(n31687) );
  XOR U31308 ( .A(n31689), .B(n31686), .Z(n31688) );
  XNOR U31309 ( .A(n31309), .B(n31682), .Z(n31684) );
  XOR U31310 ( .A(n31690), .B(n31691), .Z(n31309) );
  AND U31311 ( .A(n873), .B(n31692), .Z(n31691) );
  XOR U31312 ( .A(n31693), .B(n31690), .Z(n31692) );
  XOR U31313 ( .A(n31694), .B(n31695), .Z(n31682) );
  AND U31314 ( .A(n31696), .B(n31697), .Z(n31695) );
  XOR U31315 ( .A(n31694), .B(n31324), .Z(n31697) );
  XOR U31316 ( .A(n31698), .B(n31699), .Z(n31324) );
  AND U31317 ( .A(n875), .B(n31700), .Z(n31699) );
  XOR U31318 ( .A(n31701), .B(n31698), .Z(n31700) );
  XNOR U31319 ( .A(n31321), .B(n31694), .Z(n31696) );
  XOR U31320 ( .A(n31702), .B(n31703), .Z(n31321) );
  AND U31321 ( .A(n873), .B(n31704), .Z(n31703) );
  XOR U31322 ( .A(n31705), .B(n31702), .Z(n31704) );
  XOR U31323 ( .A(n31706), .B(n31707), .Z(n31694) );
  AND U31324 ( .A(n31708), .B(n31709), .Z(n31707) );
  XOR U31325 ( .A(n31706), .B(n31336), .Z(n31709) );
  XOR U31326 ( .A(n31710), .B(n31711), .Z(n31336) );
  AND U31327 ( .A(n875), .B(n31712), .Z(n31711) );
  XOR U31328 ( .A(n31713), .B(n31710), .Z(n31712) );
  XNOR U31329 ( .A(n31333), .B(n31706), .Z(n31708) );
  XOR U31330 ( .A(n31714), .B(n31715), .Z(n31333) );
  AND U31331 ( .A(n873), .B(n31716), .Z(n31715) );
  XOR U31332 ( .A(n31717), .B(n31714), .Z(n31716) );
  XOR U31333 ( .A(n31718), .B(n31719), .Z(n31706) );
  AND U31334 ( .A(n31720), .B(n31721), .Z(n31719) );
  XOR U31335 ( .A(n31718), .B(n31348), .Z(n31721) );
  XOR U31336 ( .A(n31722), .B(n31723), .Z(n31348) );
  AND U31337 ( .A(n875), .B(n31724), .Z(n31723) );
  XOR U31338 ( .A(n31725), .B(n31722), .Z(n31724) );
  XNOR U31339 ( .A(n31345), .B(n31718), .Z(n31720) );
  XOR U31340 ( .A(n31726), .B(n31727), .Z(n31345) );
  AND U31341 ( .A(n873), .B(n31728), .Z(n31727) );
  XOR U31342 ( .A(n31729), .B(n31726), .Z(n31728) );
  XOR U31343 ( .A(n31730), .B(n31731), .Z(n31718) );
  AND U31344 ( .A(n31732), .B(n31733), .Z(n31731) );
  XOR U31345 ( .A(n31730), .B(n31360), .Z(n31733) );
  XOR U31346 ( .A(n31734), .B(n31735), .Z(n31360) );
  AND U31347 ( .A(n875), .B(n31736), .Z(n31735) );
  XOR U31348 ( .A(n31737), .B(n31734), .Z(n31736) );
  XNOR U31349 ( .A(n31357), .B(n31730), .Z(n31732) );
  XOR U31350 ( .A(n31738), .B(n31739), .Z(n31357) );
  AND U31351 ( .A(n873), .B(n31740), .Z(n31739) );
  XOR U31352 ( .A(n31741), .B(n31738), .Z(n31740) );
  XOR U31353 ( .A(n31742), .B(n31743), .Z(n31730) );
  AND U31354 ( .A(n31744), .B(n31745), .Z(n31743) );
  XOR U31355 ( .A(n31742), .B(n31372), .Z(n31745) );
  XOR U31356 ( .A(n31746), .B(n31747), .Z(n31372) );
  AND U31357 ( .A(n875), .B(n31748), .Z(n31747) );
  XOR U31358 ( .A(n31749), .B(n31746), .Z(n31748) );
  XNOR U31359 ( .A(n31369), .B(n31742), .Z(n31744) );
  XOR U31360 ( .A(n31750), .B(n31751), .Z(n31369) );
  AND U31361 ( .A(n873), .B(n31752), .Z(n31751) );
  XOR U31362 ( .A(n31753), .B(n31750), .Z(n31752) );
  XOR U31363 ( .A(n31754), .B(n31755), .Z(n31742) );
  AND U31364 ( .A(n31756), .B(n31757), .Z(n31755) );
  XOR U31365 ( .A(n31754), .B(n31384), .Z(n31757) );
  XOR U31366 ( .A(n31758), .B(n31759), .Z(n31384) );
  AND U31367 ( .A(n875), .B(n31760), .Z(n31759) );
  XOR U31368 ( .A(n31761), .B(n31758), .Z(n31760) );
  XNOR U31369 ( .A(n31381), .B(n31754), .Z(n31756) );
  XOR U31370 ( .A(n31762), .B(n31763), .Z(n31381) );
  AND U31371 ( .A(n873), .B(n31764), .Z(n31763) );
  XOR U31372 ( .A(n31765), .B(n31762), .Z(n31764) );
  XOR U31373 ( .A(n31766), .B(n31767), .Z(n31754) );
  AND U31374 ( .A(n31768), .B(n31769), .Z(n31767) );
  XOR U31375 ( .A(n31766), .B(n31396), .Z(n31769) );
  XOR U31376 ( .A(n31770), .B(n31771), .Z(n31396) );
  AND U31377 ( .A(n875), .B(n31772), .Z(n31771) );
  XOR U31378 ( .A(n31773), .B(n31770), .Z(n31772) );
  XNOR U31379 ( .A(n31393), .B(n31766), .Z(n31768) );
  XOR U31380 ( .A(n31774), .B(n31775), .Z(n31393) );
  AND U31381 ( .A(n873), .B(n31776), .Z(n31775) );
  XOR U31382 ( .A(n31777), .B(n31774), .Z(n31776) );
  XOR U31383 ( .A(n31778), .B(n31779), .Z(n31766) );
  AND U31384 ( .A(n31780), .B(n31781), .Z(n31779) );
  XOR U31385 ( .A(n31778), .B(n31408), .Z(n31781) );
  XOR U31386 ( .A(n31782), .B(n31783), .Z(n31408) );
  AND U31387 ( .A(n875), .B(n31784), .Z(n31783) );
  XOR U31388 ( .A(n31785), .B(n31782), .Z(n31784) );
  XNOR U31389 ( .A(n31405), .B(n31778), .Z(n31780) );
  XOR U31390 ( .A(n31786), .B(n31787), .Z(n31405) );
  AND U31391 ( .A(n873), .B(n31788), .Z(n31787) );
  XOR U31392 ( .A(n31789), .B(n31786), .Z(n31788) );
  XOR U31393 ( .A(n31790), .B(n31791), .Z(n31778) );
  AND U31394 ( .A(n31792), .B(n31793), .Z(n31791) );
  XNOR U31395 ( .A(n31794), .B(n31421), .Z(n31793) );
  XOR U31396 ( .A(n31795), .B(n31796), .Z(n31421) );
  AND U31397 ( .A(n875), .B(n31797), .Z(n31796) );
  XOR U31398 ( .A(n31795), .B(n31798), .Z(n31797) );
  XNOR U31399 ( .A(n31418), .B(n31790), .Z(n31792) );
  XOR U31400 ( .A(n31799), .B(n31800), .Z(n31418) );
  AND U31401 ( .A(n873), .B(n31801), .Z(n31800) );
  XOR U31402 ( .A(n31799), .B(n31802), .Z(n31801) );
  IV U31403 ( .A(n31794), .Z(n31790) );
  AND U31404 ( .A(n31426), .B(n31429), .Z(n31794) );
  XNOR U31405 ( .A(n31803), .B(n31804), .Z(n31429) );
  AND U31406 ( .A(n875), .B(n31805), .Z(n31804) );
  XNOR U31407 ( .A(n31806), .B(n31803), .Z(n31805) );
  XOR U31408 ( .A(n31807), .B(n31808), .Z(n875) );
  AND U31409 ( .A(n31809), .B(n31810), .Z(n31808) );
  XOR U31410 ( .A(n31807), .B(n31437), .Z(n31810) );
  XNOR U31411 ( .A(n31811), .B(n31812), .Z(n31437) );
  AND U31412 ( .A(n31813), .B(n563), .Z(n31812) );
  AND U31413 ( .A(n31811), .B(n31814), .Z(n31813) );
  XNOR U31414 ( .A(n31434), .B(n31807), .Z(n31809) );
  XOR U31415 ( .A(n31815), .B(n31816), .Z(n31434) );
  AND U31416 ( .A(n31817), .B(n561), .Z(n31816) );
  NOR U31417 ( .A(n31815), .B(n31818), .Z(n31817) );
  XOR U31418 ( .A(n31819), .B(n31820), .Z(n31807) );
  AND U31419 ( .A(n31821), .B(n31822), .Z(n31820) );
  XOR U31420 ( .A(n31819), .B(n31449), .Z(n31822) );
  XOR U31421 ( .A(n31823), .B(n31824), .Z(n31449) );
  AND U31422 ( .A(n563), .B(n31825), .Z(n31824) );
  XOR U31423 ( .A(n31826), .B(n31823), .Z(n31825) );
  XNOR U31424 ( .A(n31446), .B(n31819), .Z(n31821) );
  XOR U31425 ( .A(n31827), .B(n31828), .Z(n31446) );
  AND U31426 ( .A(n561), .B(n31829), .Z(n31828) );
  XOR U31427 ( .A(n31830), .B(n31827), .Z(n31829) );
  XOR U31428 ( .A(n31831), .B(n31832), .Z(n31819) );
  AND U31429 ( .A(n31833), .B(n31834), .Z(n31832) );
  XOR U31430 ( .A(n31831), .B(n31461), .Z(n31834) );
  XOR U31431 ( .A(n31835), .B(n31836), .Z(n31461) );
  AND U31432 ( .A(n563), .B(n31837), .Z(n31836) );
  XOR U31433 ( .A(n31838), .B(n31835), .Z(n31837) );
  XNOR U31434 ( .A(n31458), .B(n31831), .Z(n31833) );
  XOR U31435 ( .A(n31839), .B(n31840), .Z(n31458) );
  AND U31436 ( .A(n561), .B(n31841), .Z(n31840) );
  XOR U31437 ( .A(n31842), .B(n31839), .Z(n31841) );
  XOR U31438 ( .A(n31843), .B(n31844), .Z(n31831) );
  AND U31439 ( .A(n31845), .B(n31846), .Z(n31844) );
  XOR U31440 ( .A(n31843), .B(n31473), .Z(n31846) );
  XOR U31441 ( .A(n31847), .B(n31848), .Z(n31473) );
  AND U31442 ( .A(n563), .B(n31849), .Z(n31848) );
  XOR U31443 ( .A(n31850), .B(n31847), .Z(n31849) );
  XNOR U31444 ( .A(n31470), .B(n31843), .Z(n31845) );
  XOR U31445 ( .A(n31851), .B(n31852), .Z(n31470) );
  AND U31446 ( .A(n561), .B(n31853), .Z(n31852) );
  XOR U31447 ( .A(n31854), .B(n31851), .Z(n31853) );
  XOR U31448 ( .A(n31855), .B(n31856), .Z(n31843) );
  AND U31449 ( .A(n31857), .B(n31858), .Z(n31856) );
  XOR U31450 ( .A(n31855), .B(n31485), .Z(n31858) );
  XOR U31451 ( .A(n31859), .B(n31860), .Z(n31485) );
  AND U31452 ( .A(n563), .B(n31861), .Z(n31860) );
  XOR U31453 ( .A(n31862), .B(n31859), .Z(n31861) );
  XNOR U31454 ( .A(n31482), .B(n31855), .Z(n31857) );
  XOR U31455 ( .A(n31863), .B(n31864), .Z(n31482) );
  AND U31456 ( .A(n561), .B(n31865), .Z(n31864) );
  XOR U31457 ( .A(n31866), .B(n31863), .Z(n31865) );
  XOR U31458 ( .A(n31867), .B(n31868), .Z(n31855) );
  AND U31459 ( .A(n31869), .B(n31870), .Z(n31868) );
  XOR U31460 ( .A(n31867), .B(n31497), .Z(n31870) );
  XOR U31461 ( .A(n31871), .B(n31872), .Z(n31497) );
  AND U31462 ( .A(n563), .B(n31873), .Z(n31872) );
  XOR U31463 ( .A(n31874), .B(n31871), .Z(n31873) );
  XNOR U31464 ( .A(n31494), .B(n31867), .Z(n31869) );
  XOR U31465 ( .A(n31875), .B(n31876), .Z(n31494) );
  AND U31466 ( .A(n561), .B(n31877), .Z(n31876) );
  XOR U31467 ( .A(n31878), .B(n31875), .Z(n31877) );
  XOR U31468 ( .A(n31879), .B(n31880), .Z(n31867) );
  AND U31469 ( .A(n31881), .B(n31882), .Z(n31880) );
  XOR U31470 ( .A(n31879), .B(n31509), .Z(n31882) );
  XOR U31471 ( .A(n31883), .B(n31884), .Z(n31509) );
  AND U31472 ( .A(n563), .B(n31885), .Z(n31884) );
  XOR U31473 ( .A(n31886), .B(n31883), .Z(n31885) );
  XNOR U31474 ( .A(n31506), .B(n31879), .Z(n31881) );
  XOR U31475 ( .A(n31887), .B(n31888), .Z(n31506) );
  AND U31476 ( .A(n561), .B(n31889), .Z(n31888) );
  XOR U31477 ( .A(n31890), .B(n31887), .Z(n31889) );
  XOR U31478 ( .A(n31891), .B(n31892), .Z(n31879) );
  AND U31479 ( .A(n31893), .B(n31894), .Z(n31892) );
  XOR U31480 ( .A(n31891), .B(n31521), .Z(n31894) );
  XOR U31481 ( .A(n31895), .B(n31896), .Z(n31521) );
  AND U31482 ( .A(n563), .B(n31897), .Z(n31896) );
  XOR U31483 ( .A(n31898), .B(n31895), .Z(n31897) );
  XNOR U31484 ( .A(n31518), .B(n31891), .Z(n31893) );
  XOR U31485 ( .A(n31899), .B(n31900), .Z(n31518) );
  AND U31486 ( .A(n561), .B(n31901), .Z(n31900) );
  XOR U31487 ( .A(n31902), .B(n31899), .Z(n31901) );
  XOR U31488 ( .A(n31903), .B(n31904), .Z(n31891) );
  AND U31489 ( .A(n31905), .B(n31906), .Z(n31904) );
  XOR U31490 ( .A(n31903), .B(n31533), .Z(n31906) );
  XOR U31491 ( .A(n31907), .B(n31908), .Z(n31533) );
  AND U31492 ( .A(n563), .B(n31909), .Z(n31908) );
  XOR U31493 ( .A(n31910), .B(n31907), .Z(n31909) );
  XNOR U31494 ( .A(n31530), .B(n31903), .Z(n31905) );
  XOR U31495 ( .A(n31911), .B(n31912), .Z(n31530) );
  AND U31496 ( .A(n561), .B(n31913), .Z(n31912) );
  XOR U31497 ( .A(n31914), .B(n31911), .Z(n31913) );
  XOR U31498 ( .A(n31915), .B(n31916), .Z(n31903) );
  AND U31499 ( .A(n31917), .B(n31918), .Z(n31916) );
  XOR U31500 ( .A(n31915), .B(n31545), .Z(n31918) );
  XOR U31501 ( .A(n31919), .B(n31920), .Z(n31545) );
  AND U31502 ( .A(n563), .B(n31921), .Z(n31920) );
  XOR U31503 ( .A(n31922), .B(n31919), .Z(n31921) );
  XNOR U31504 ( .A(n31542), .B(n31915), .Z(n31917) );
  XOR U31505 ( .A(n31923), .B(n31924), .Z(n31542) );
  AND U31506 ( .A(n561), .B(n31925), .Z(n31924) );
  XOR U31507 ( .A(n31926), .B(n31923), .Z(n31925) );
  XOR U31508 ( .A(n31927), .B(n31928), .Z(n31915) );
  AND U31509 ( .A(n31929), .B(n31930), .Z(n31928) );
  XOR U31510 ( .A(n31927), .B(n31557), .Z(n31930) );
  XOR U31511 ( .A(n31931), .B(n31932), .Z(n31557) );
  AND U31512 ( .A(n563), .B(n31933), .Z(n31932) );
  XOR U31513 ( .A(n31934), .B(n31931), .Z(n31933) );
  XNOR U31514 ( .A(n31554), .B(n31927), .Z(n31929) );
  XOR U31515 ( .A(n31935), .B(n31936), .Z(n31554) );
  AND U31516 ( .A(n561), .B(n31937), .Z(n31936) );
  XOR U31517 ( .A(n31938), .B(n31935), .Z(n31937) );
  XOR U31518 ( .A(n31939), .B(n31940), .Z(n31927) );
  AND U31519 ( .A(n31941), .B(n31942), .Z(n31940) );
  XOR U31520 ( .A(n31939), .B(n31569), .Z(n31942) );
  XOR U31521 ( .A(n31943), .B(n31944), .Z(n31569) );
  AND U31522 ( .A(n563), .B(n31945), .Z(n31944) );
  XOR U31523 ( .A(n31946), .B(n31943), .Z(n31945) );
  XNOR U31524 ( .A(n31566), .B(n31939), .Z(n31941) );
  XOR U31525 ( .A(n31947), .B(n31948), .Z(n31566) );
  AND U31526 ( .A(n561), .B(n31949), .Z(n31948) );
  XOR U31527 ( .A(n31950), .B(n31947), .Z(n31949) );
  XOR U31528 ( .A(n31951), .B(n31952), .Z(n31939) );
  AND U31529 ( .A(n31953), .B(n31954), .Z(n31952) );
  XOR U31530 ( .A(n31951), .B(n31581), .Z(n31954) );
  XOR U31531 ( .A(n31955), .B(n31956), .Z(n31581) );
  AND U31532 ( .A(n563), .B(n31957), .Z(n31956) );
  XOR U31533 ( .A(n31958), .B(n31955), .Z(n31957) );
  XNOR U31534 ( .A(n31578), .B(n31951), .Z(n31953) );
  XOR U31535 ( .A(n31959), .B(n31960), .Z(n31578) );
  AND U31536 ( .A(n561), .B(n31961), .Z(n31960) );
  XOR U31537 ( .A(n31962), .B(n31959), .Z(n31961) );
  XOR U31538 ( .A(n31963), .B(n31964), .Z(n31951) );
  AND U31539 ( .A(n31965), .B(n31966), .Z(n31964) );
  XOR U31540 ( .A(n31963), .B(n31593), .Z(n31966) );
  XOR U31541 ( .A(n31967), .B(n31968), .Z(n31593) );
  AND U31542 ( .A(n563), .B(n31969), .Z(n31968) );
  XOR U31543 ( .A(n31970), .B(n31967), .Z(n31969) );
  XNOR U31544 ( .A(n31590), .B(n31963), .Z(n31965) );
  XOR U31545 ( .A(n31971), .B(n31972), .Z(n31590) );
  AND U31546 ( .A(n561), .B(n31973), .Z(n31972) );
  XOR U31547 ( .A(n31974), .B(n31971), .Z(n31973) );
  XOR U31548 ( .A(n31975), .B(n31976), .Z(n31963) );
  AND U31549 ( .A(n31977), .B(n31978), .Z(n31976) );
  XOR U31550 ( .A(n31975), .B(n31605), .Z(n31978) );
  XOR U31551 ( .A(n31979), .B(n31980), .Z(n31605) );
  AND U31552 ( .A(n563), .B(n31981), .Z(n31980) );
  XOR U31553 ( .A(n31982), .B(n31979), .Z(n31981) );
  XNOR U31554 ( .A(n31602), .B(n31975), .Z(n31977) );
  XOR U31555 ( .A(n31983), .B(n31984), .Z(n31602) );
  AND U31556 ( .A(n561), .B(n31985), .Z(n31984) );
  XOR U31557 ( .A(n31986), .B(n31983), .Z(n31985) );
  XOR U31558 ( .A(n31987), .B(n31988), .Z(n31975) );
  AND U31559 ( .A(n31989), .B(n31990), .Z(n31988) );
  XOR U31560 ( .A(n31987), .B(n31617), .Z(n31990) );
  XOR U31561 ( .A(n31991), .B(n31992), .Z(n31617) );
  AND U31562 ( .A(n563), .B(n31993), .Z(n31992) );
  XOR U31563 ( .A(n31994), .B(n31991), .Z(n31993) );
  XNOR U31564 ( .A(n31614), .B(n31987), .Z(n31989) );
  XOR U31565 ( .A(n31995), .B(n31996), .Z(n31614) );
  AND U31566 ( .A(n561), .B(n31997), .Z(n31996) );
  XOR U31567 ( .A(n31998), .B(n31995), .Z(n31997) );
  XOR U31568 ( .A(n31999), .B(n32000), .Z(n31987) );
  AND U31569 ( .A(n32001), .B(n32002), .Z(n32000) );
  XOR U31570 ( .A(n31999), .B(n31629), .Z(n32002) );
  XOR U31571 ( .A(n32003), .B(n32004), .Z(n31629) );
  AND U31572 ( .A(n563), .B(n32005), .Z(n32004) );
  XOR U31573 ( .A(n32006), .B(n32003), .Z(n32005) );
  XNOR U31574 ( .A(n31626), .B(n31999), .Z(n32001) );
  XOR U31575 ( .A(n32007), .B(n32008), .Z(n31626) );
  AND U31576 ( .A(n561), .B(n32009), .Z(n32008) );
  XOR U31577 ( .A(n32010), .B(n32007), .Z(n32009) );
  XOR U31578 ( .A(n32011), .B(n32012), .Z(n31999) );
  AND U31579 ( .A(n32013), .B(n32014), .Z(n32012) );
  XOR U31580 ( .A(n32011), .B(n31641), .Z(n32014) );
  XOR U31581 ( .A(n32015), .B(n32016), .Z(n31641) );
  AND U31582 ( .A(n563), .B(n32017), .Z(n32016) );
  XOR U31583 ( .A(n32018), .B(n32015), .Z(n32017) );
  XNOR U31584 ( .A(n31638), .B(n32011), .Z(n32013) );
  XOR U31585 ( .A(n32019), .B(n32020), .Z(n31638) );
  AND U31586 ( .A(n561), .B(n32021), .Z(n32020) );
  XOR U31587 ( .A(n32022), .B(n32019), .Z(n32021) );
  XOR U31588 ( .A(n32023), .B(n32024), .Z(n32011) );
  AND U31589 ( .A(n32025), .B(n32026), .Z(n32024) );
  XOR U31590 ( .A(n32023), .B(n31653), .Z(n32026) );
  XOR U31591 ( .A(n32027), .B(n32028), .Z(n31653) );
  AND U31592 ( .A(n563), .B(n32029), .Z(n32028) );
  XOR U31593 ( .A(n32030), .B(n32027), .Z(n32029) );
  XNOR U31594 ( .A(n31650), .B(n32023), .Z(n32025) );
  XOR U31595 ( .A(n32031), .B(n32032), .Z(n31650) );
  AND U31596 ( .A(n561), .B(n32033), .Z(n32032) );
  XOR U31597 ( .A(n32034), .B(n32031), .Z(n32033) );
  XOR U31598 ( .A(n32035), .B(n32036), .Z(n32023) );
  AND U31599 ( .A(n32037), .B(n32038), .Z(n32036) );
  XOR U31600 ( .A(n32035), .B(n31665), .Z(n32038) );
  XOR U31601 ( .A(n32039), .B(n32040), .Z(n31665) );
  AND U31602 ( .A(n563), .B(n32041), .Z(n32040) );
  XOR U31603 ( .A(n32042), .B(n32039), .Z(n32041) );
  XNOR U31604 ( .A(n31662), .B(n32035), .Z(n32037) );
  XOR U31605 ( .A(n32043), .B(n32044), .Z(n31662) );
  AND U31606 ( .A(n561), .B(n32045), .Z(n32044) );
  XOR U31607 ( .A(n32046), .B(n32043), .Z(n32045) );
  XOR U31608 ( .A(n32047), .B(n32048), .Z(n32035) );
  AND U31609 ( .A(n32049), .B(n32050), .Z(n32048) );
  XOR U31610 ( .A(n32047), .B(n31677), .Z(n32050) );
  XOR U31611 ( .A(n32051), .B(n32052), .Z(n31677) );
  AND U31612 ( .A(n563), .B(n32053), .Z(n32052) );
  XOR U31613 ( .A(n32054), .B(n32051), .Z(n32053) );
  XNOR U31614 ( .A(n31674), .B(n32047), .Z(n32049) );
  XOR U31615 ( .A(n32055), .B(n32056), .Z(n31674) );
  AND U31616 ( .A(n561), .B(n32057), .Z(n32056) );
  XOR U31617 ( .A(n32058), .B(n32055), .Z(n32057) );
  XOR U31618 ( .A(n32059), .B(n32060), .Z(n32047) );
  AND U31619 ( .A(n32061), .B(n32062), .Z(n32060) );
  XOR U31620 ( .A(n32059), .B(n31689), .Z(n32062) );
  XOR U31621 ( .A(n32063), .B(n32064), .Z(n31689) );
  AND U31622 ( .A(n563), .B(n32065), .Z(n32064) );
  XOR U31623 ( .A(n32066), .B(n32063), .Z(n32065) );
  XNOR U31624 ( .A(n31686), .B(n32059), .Z(n32061) );
  XOR U31625 ( .A(n32067), .B(n32068), .Z(n31686) );
  AND U31626 ( .A(n561), .B(n32069), .Z(n32068) );
  XOR U31627 ( .A(n32070), .B(n32067), .Z(n32069) );
  XOR U31628 ( .A(n32071), .B(n32072), .Z(n32059) );
  AND U31629 ( .A(n32073), .B(n32074), .Z(n32072) );
  XOR U31630 ( .A(n32071), .B(n31701), .Z(n32074) );
  XOR U31631 ( .A(n32075), .B(n32076), .Z(n31701) );
  AND U31632 ( .A(n563), .B(n32077), .Z(n32076) );
  XOR U31633 ( .A(n32078), .B(n32075), .Z(n32077) );
  XNOR U31634 ( .A(n31698), .B(n32071), .Z(n32073) );
  XOR U31635 ( .A(n32079), .B(n32080), .Z(n31698) );
  AND U31636 ( .A(n561), .B(n32081), .Z(n32080) );
  XOR U31637 ( .A(n32082), .B(n32079), .Z(n32081) );
  XOR U31638 ( .A(n32083), .B(n32084), .Z(n32071) );
  AND U31639 ( .A(n32085), .B(n32086), .Z(n32084) );
  XOR U31640 ( .A(n32083), .B(n31713), .Z(n32086) );
  XOR U31641 ( .A(n32087), .B(n32088), .Z(n31713) );
  AND U31642 ( .A(n563), .B(n32089), .Z(n32088) );
  XOR U31643 ( .A(n32090), .B(n32087), .Z(n32089) );
  XNOR U31644 ( .A(n31710), .B(n32083), .Z(n32085) );
  XOR U31645 ( .A(n32091), .B(n32092), .Z(n31710) );
  AND U31646 ( .A(n561), .B(n32093), .Z(n32092) );
  XOR U31647 ( .A(n32094), .B(n32091), .Z(n32093) );
  XOR U31648 ( .A(n32095), .B(n32096), .Z(n32083) );
  AND U31649 ( .A(n32097), .B(n32098), .Z(n32096) );
  XOR U31650 ( .A(n32095), .B(n31725), .Z(n32098) );
  XOR U31651 ( .A(n32099), .B(n32100), .Z(n31725) );
  AND U31652 ( .A(n563), .B(n32101), .Z(n32100) );
  XOR U31653 ( .A(n32102), .B(n32099), .Z(n32101) );
  XNOR U31654 ( .A(n31722), .B(n32095), .Z(n32097) );
  XOR U31655 ( .A(n32103), .B(n32104), .Z(n31722) );
  AND U31656 ( .A(n561), .B(n32105), .Z(n32104) );
  XOR U31657 ( .A(n32106), .B(n32103), .Z(n32105) );
  XOR U31658 ( .A(n32107), .B(n32108), .Z(n32095) );
  AND U31659 ( .A(n32109), .B(n32110), .Z(n32108) );
  XOR U31660 ( .A(n32107), .B(n31737), .Z(n32110) );
  XOR U31661 ( .A(n32111), .B(n32112), .Z(n31737) );
  AND U31662 ( .A(n563), .B(n32113), .Z(n32112) );
  XOR U31663 ( .A(n32114), .B(n32111), .Z(n32113) );
  XNOR U31664 ( .A(n31734), .B(n32107), .Z(n32109) );
  XOR U31665 ( .A(n32115), .B(n32116), .Z(n31734) );
  AND U31666 ( .A(n561), .B(n32117), .Z(n32116) );
  XOR U31667 ( .A(n32118), .B(n32115), .Z(n32117) );
  XOR U31668 ( .A(n32119), .B(n32120), .Z(n32107) );
  AND U31669 ( .A(n32121), .B(n32122), .Z(n32120) );
  XOR U31670 ( .A(n32119), .B(n31749), .Z(n32122) );
  XOR U31671 ( .A(n32123), .B(n32124), .Z(n31749) );
  AND U31672 ( .A(n563), .B(n32125), .Z(n32124) );
  XOR U31673 ( .A(n32126), .B(n32123), .Z(n32125) );
  XNOR U31674 ( .A(n31746), .B(n32119), .Z(n32121) );
  XOR U31675 ( .A(n32127), .B(n32128), .Z(n31746) );
  AND U31676 ( .A(n561), .B(n32129), .Z(n32128) );
  XOR U31677 ( .A(n32130), .B(n32127), .Z(n32129) );
  XOR U31678 ( .A(n32131), .B(n32132), .Z(n32119) );
  AND U31679 ( .A(n32133), .B(n32134), .Z(n32132) );
  XOR U31680 ( .A(n32131), .B(n31761), .Z(n32134) );
  XOR U31681 ( .A(n32135), .B(n32136), .Z(n31761) );
  AND U31682 ( .A(n563), .B(n32137), .Z(n32136) );
  XOR U31683 ( .A(n32138), .B(n32135), .Z(n32137) );
  XNOR U31684 ( .A(n31758), .B(n32131), .Z(n32133) );
  XOR U31685 ( .A(n32139), .B(n32140), .Z(n31758) );
  AND U31686 ( .A(n561), .B(n32141), .Z(n32140) );
  XOR U31687 ( .A(n32142), .B(n32139), .Z(n32141) );
  XOR U31688 ( .A(n32143), .B(n32144), .Z(n32131) );
  AND U31689 ( .A(n32145), .B(n32146), .Z(n32144) );
  XOR U31690 ( .A(n32143), .B(n31773), .Z(n32146) );
  XOR U31691 ( .A(n32147), .B(n32148), .Z(n31773) );
  AND U31692 ( .A(n563), .B(n32149), .Z(n32148) );
  XOR U31693 ( .A(n32150), .B(n32147), .Z(n32149) );
  XNOR U31694 ( .A(n31770), .B(n32143), .Z(n32145) );
  XOR U31695 ( .A(n32151), .B(n32152), .Z(n31770) );
  AND U31696 ( .A(n561), .B(n32153), .Z(n32152) );
  XOR U31697 ( .A(n32154), .B(n32151), .Z(n32153) );
  XOR U31698 ( .A(n32155), .B(n32156), .Z(n32143) );
  AND U31699 ( .A(n32157), .B(n32158), .Z(n32156) );
  XOR U31700 ( .A(n32155), .B(n31785), .Z(n32158) );
  XOR U31701 ( .A(n32159), .B(n32160), .Z(n31785) );
  AND U31702 ( .A(n563), .B(n32161), .Z(n32160) );
  XOR U31703 ( .A(n32162), .B(n32159), .Z(n32161) );
  XNOR U31704 ( .A(n31782), .B(n32155), .Z(n32157) );
  XOR U31705 ( .A(n32163), .B(n32164), .Z(n31782) );
  AND U31706 ( .A(n561), .B(n32165), .Z(n32164) );
  XOR U31707 ( .A(n32166), .B(n32163), .Z(n32165) );
  XOR U31708 ( .A(n32167), .B(n32168), .Z(n32155) );
  AND U31709 ( .A(n32169), .B(n32170), .Z(n32168) );
  XNOR U31710 ( .A(n32171), .B(n31798), .Z(n32170) );
  XOR U31711 ( .A(n32172), .B(n32173), .Z(n31798) );
  AND U31712 ( .A(n563), .B(n32174), .Z(n32173) );
  XOR U31713 ( .A(n32172), .B(n32175), .Z(n32174) );
  XNOR U31714 ( .A(n31795), .B(n32167), .Z(n32169) );
  XOR U31715 ( .A(n32176), .B(n32177), .Z(n31795) );
  AND U31716 ( .A(n561), .B(n32178), .Z(n32177) );
  XOR U31717 ( .A(n32176), .B(n32179), .Z(n32178) );
  IV U31718 ( .A(n32171), .Z(n32167) );
  AND U31719 ( .A(n31803), .B(n31806), .Z(n32171) );
  XNOR U31720 ( .A(n32180), .B(n32181), .Z(n31806) );
  AND U31721 ( .A(n563), .B(n32182), .Z(n32181) );
  XNOR U31722 ( .A(n32183), .B(n32180), .Z(n32182) );
  XOR U31723 ( .A(n32184), .B(n32185), .Z(n563) );
  AND U31724 ( .A(n32186), .B(n32187), .Z(n32185) );
  XOR U31725 ( .A(n31814), .B(n32184), .Z(n32187) );
  IV U31726 ( .A(n32188), .Z(n31814) );
  AND U31727 ( .A(p_input[4095]), .B(p_input[4063]), .Z(n32188) );
  XOR U31728 ( .A(n32184), .B(n31811), .Z(n32186) );
  AND U31729 ( .A(p_input[3999]), .B(p_input[4031]), .Z(n31811) );
  XOR U31730 ( .A(n32189), .B(n32190), .Z(n32184) );
  AND U31731 ( .A(n32191), .B(n32192), .Z(n32190) );
  XOR U31732 ( .A(n32189), .B(n31826), .Z(n32192) );
  XNOR U31733 ( .A(p_input[4062]), .B(n32193), .Z(n31826) );
  AND U31734 ( .A(n691), .B(n32194), .Z(n32193) );
  XOR U31735 ( .A(p_input[4094]), .B(p_input[4062]), .Z(n32194) );
  XNOR U31736 ( .A(n31823), .B(n32189), .Z(n32191) );
  XOR U31737 ( .A(n32195), .B(n32196), .Z(n31823) );
  AND U31738 ( .A(n689), .B(n32197), .Z(n32196) );
  XOR U31739 ( .A(p_input[4030]), .B(p_input[3998]), .Z(n32197) );
  XOR U31740 ( .A(n32198), .B(n32199), .Z(n32189) );
  AND U31741 ( .A(n32200), .B(n32201), .Z(n32199) );
  XOR U31742 ( .A(n32198), .B(n31838), .Z(n32201) );
  XNOR U31743 ( .A(p_input[4061]), .B(n32202), .Z(n31838) );
  AND U31744 ( .A(n691), .B(n32203), .Z(n32202) );
  XOR U31745 ( .A(p_input[4093]), .B(p_input[4061]), .Z(n32203) );
  XNOR U31746 ( .A(n31835), .B(n32198), .Z(n32200) );
  XOR U31747 ( .A(n32204), .B(n32205), .Z(n31835) );
  AND U31748 ( .A(n689), .B(n32206), .Z(n32205) );
  XOR U31749 ( .A(p_input[4029]), .B(p_input[3997]), .Z(n32206) );
  XOR U31750 ( .A(n32207), .B(n32208), .Z(n32198) );
  AND U31751 ( .A(n32209), .B(n32210), .Z(n32208) );
  XOR U31752 ( .A(n32207), .B(n31850), .Z(n32210) );
  XNOR U31753 ( .A(p_input[4060]), .B(n32211), .Z(n31850) );
  AND U31754 ( .A(n691), .B(n32212), .Z(n32211) );
  XOR U31755 ( .A(p_input[4092]), .B(p_input[4060]), .Z(n32212) );
  XNOR U31756 ( .A(n31847), .B(n32207), .Z(n32209) );
  XOR U31757 ( .A(n32213), .B(n32214), .Z(n31847) );
  AND U31758 ( .A(n689), .B(n32215), .Z(n32214) );
  XOR U31759 ( .A(p_input[4028]), .B(p_input[3996]), .Z(n32215) );
  XOR U31760 ( .A(n32216), .B(n32217), .Z(n32207) );
  AND U31761 ( .A(n32218), .B(n32219), .Z(n32217) );
  XOR U31762 ( .A(n32216), .B(n31862), .Z(n32219) );
  XNOR U31763 ( .A(p_input[4059]), .B(n32220), .Z(n31862) );
  AND U31764 ( .A(n691), .B(n32221), .Z(n32220) );
  XOR U31765 ( .A(p_input[4091]), .B(p_input[4059]), .Z(n32221) );
  XNOR U31766 ( .A(n31859), .B(n32216), .Z(n32218) );
  XOR U31767 ( .A(n32222), .B(n32223), .Z(n31859) );
  AND U31768 ( .A(n689), .B(n32224), .Z(n32223) );
  XOR U31769 ( .A(p_input[4027]), .B(p_input[3995]), .Z(n32224) );
  XOR U31770 ( .A(n32225), .B(n32226), .Z(n32216) );
  AND U31771 ( .A(n32227), .B(n32228), .Z(n32226) );
  XOR U31772 ( .A(n32225), .B(n31874), .Z(n32228) );
  XNOR U31773 ( .A(p_input[4058]), .B(n32229), .Z(n31874) );
  AND U31774 ( .A(n691), .B(n32230), .Z(n32229) );
  XOR U31775 ( .A(p_input[4090]), .B(p_input[4058]), .Z(n32230) );
  XNOR U31776 ( .A(n31871), .B(n32225), .Z(n32227) );
  XOR U31777 ( .A(n32231), .B(n32232), .Z(n31871) );
  AND U31778 ( .A(n689), .B(n32233), .Z(n32232) );
  XOR U31779 ( .A(p_input[4026]), .B(p_input[3994]), .Z(n32233) );
  XOR U31780 ( .A(n32234), .B(n32235), .Z(n32225) );
  AND U31781 ( .A(n32236), .B(n32237), .Z(n32235) );
  XOR U31782 ( .A(n32234), .B(n31886), .Z(n32237) );
  XNOR U31783 ( .A(p_input[4057]), .B(n32238), .Z(n31886) );
  AND U31784 ( .A(n691), .B(n32239), .Z(n32238) );
  XOR U31785 ( .A(p_input[4089]), .B(p_input[4057]), .Z(n32239) );
  XNOR U31786 ( .A(n31883), .B(n32234), .Z(n32236) );
  XOR U31787 ( .A(n32240), .B(n32241), .Z(n31883) );
  AND U31788 ( .A(n689), .B(n32242), .Z(n32241) );
  XOR U31789 ( .A(p_input[4025]), .B(p_input[3993]), .Z(n32242) );
  XOR U31790 ( .A(n32243), .B(n32244), .Z(n32234) );
  AND U31791 ( .A(n32245), .B(n32246), .Z(n32244) );
  XOR U31792 ( .A(n32243), .B(n31898), .Z(n32246) );
  XNOR U31793 ( .A(p_input[4056]), .B(n32247), .Z(n31898) );
  AND U31794 ( .A(n691), .B(n32248), .Z(n32247) );
  XOR U31795 ( .A(p_input[4088]), .B(p_input[4056]), .Z(n32248) );
  XNOR U31796 ( .A(n31895), .B(n32243), .Z(n32245) );
  XOR U31797 ( .A(n32249), .B(n32250), .Z(n31895) );
  AND U31798 ( .A(n689), .B(n32251), .Z(n32250) );
  XOR U31799 ( .A(p_input[4024]), .B(p_input[3992]), .Z(n32251) );
  XOR U31800 ( .A(n32252), .B(n32253), .Z(n32243) );
  AND U31801 ( .A(n32254), .B(n32255), .Z(n32253) );
  XOR U31802 ( .A(n32252), .B(n31910), .Z(n32255) );
  XNOR U31803 ( .A(p_input[4055]), .B(n32256), .Z(n31910) );
  AND U31804 ( .A(n691), .B(n32257), .Z(n32256) );
  XOR U31805 ( .A(p_input[4087]), .B(p_input[4055]), .Z(n32257) );
  XNOR U31806 ( .A(n31907), .B(n32252), .Z(n32254) );
  XOR U31807 ( .A(n32258), .B(n32259), .Z(n31907) );
  AND U31808 ( .A(n689), .B(n32260), .Z(n32259) );
  XOR U31809 ( .A(p_input[4023]), .B(p_input[3991]), .Z(n32260) );
  XOR U31810 ( .A(n32261), .B(n32262), .Z(n32252) );
  AND U31811 ( .A(n32263), .B(n32264), .Z(n32262) );
  XOR U31812 ( .A(n32261), .B(n31922), .Z(n32264) );
  XNOR U31813 ( .A(p_input[4054]), .B(n32265), .Z(n31922) );
  AND U31814 ( .A(n691), .B(n32266), .Z(n32265) );
  XOR U31815 ( .A(p_input[4086]), .B(p_input[4054]), .Z(n32266) );
  XNOR U31816 ( .A(n31919), .B(n32261), .Z(n32263) );
  XOR U31817 ( .A(n32267), .B(n32268), .Z(n31919) );
  AND U31818 ( .A(n689), .B(n32269), .Z(n32268) );
  XOR U31819 ( .A(p_input[4022]), .B(p_input[3990]), .Z(n32269) );
  XOR U31820 ( .A(n32270), .B(n32271), .Z(n32261) );
  AND U31821 ( .A(n32272), .B(n32273), .Z(n32271) );
  XOR U31822 ( .A(n32270), .B(n31934), .Z(n32273) );
  XNOR U31823 ( .A(p_input[4053]), .B(n32274), .Z(n31934) );
  AND U31824 ( .A(n691), .B(n32275), .Z(n32274) );
  XOR U31825 ( .A(p_input[4085]), .B(p_input[4053]), .Z(n32275) );
  XNOR U31826 ( .A(n31931), .B(n32270), .Z(n32272) );
  XOR U31827 ( .A(n32276), .B(n32277), .Z(n31931) );
  AND U31828 ( .A(n689), .B(n32278), .Z(n32277) );
  XOR U31829 ( .A(p_input[4021]), .B(p_input[3989]), .Z(n32278) );
  XOR U31830 ( .A(n32279), .B(n32280), .Z(n32270) );
  AND U31831 ( .A(n32281), .B(n32282), .Z(n32280) );
  XOR U31832 ( .A(n32279), .B(n31946), .Z(n32282) );
  XNOR U31833 ( .A(p_input[4052]), .B(n32283), .Z(n31946) );
  AND U31834 ( .A(n691), .B(n32284), .Z(n32283) );
  XOR U31835 ( .A(p_input[4084]), .B(p_input[4052]), .Z(n32284) );
  XNOR U31836 ( .A(n31943), .B(n32279), .Z(n32281) );
  XOR U31837 ( .A(n32285), .B(n32286), .Z(n31943) );
  AND U31838 ( .A(n689), .B(n32287), .Z(n32286) );
  XOR U31839 ( .A(p_input[4020]), .B(p_input[3988]), .Z(n32287) );
  XOR U31840 ( .A(n32288), .B(n32289), .Z(n32279) );
  AND U31841 ( .A(n32290), .B(n32291), .Z(n32289) );
  XOR U31842 ( .A(n32288), .B(n31958), .Z(n32291) );
  XNOR U31843 ( .A(p_input[4051]), .B(n32292), .Z(n31958) );
  AND U31844 ( .A(n691), .B(n32293), .Z(n32292) );
  XOR U31845 ( .A(p_input[4083]), .B(p_input[4051]), .Z(n32293) );
  XNOR U31846 ( .A(n31955), .B(n32288), .Z(n32290) );
  XOR U31847 ( .A(n32294), .B(n32295), .Z(n31955) );
  AND U31848 ( .A(n689), .B(n32296), .Z(n32295) );
  XOR U31849 ( .A(p_input[4019]), .B(p_input[3987]), .Z(n32296) );
  XOR U31850 ( .A(n32297), .B(n32298), .Z(n32288) );
  AND U31851 ( .A(n32299), .B(n32300), .Z(n32298) );
  XOR U31852 ( .A(n32297), .B(n31970), .Z(n32300) );
  XNOR U31853 ( .A(p_input[4050]), .B(n32301), .Z(n31970) );
  AND U31854 ( .A(n691), .B(n32302), .Z(n32301) );
  XOR U31855 ( .A(p_input[4082]), .B(p_input[4050]), .Z(n32302) );
  XNOR U31856 ( .A(n31967), .B(n32297), .Z(n32299) );
  XOR U31857 ( .A(n32303), .B(n32304), .Z(n31967) );
  AND U31858 ( .A(n689), .B(n32305), .Z(n32304) );
  XOR U31859 ( .A(p_input[4018]), .B(p_input[3986]), .Z(n32305) );
  XOR U31860 ( .A(n32306), .B(n32307), .Z(n32297) );
  AND U31861 ( .A(n32308), .B(n32309), .Z(n32307) );
  XOR U31862 ( .A(n32306), .B(n31982), .Z(n32309) );
  XNOR U31863 ( .A(p_input[4049]), .B(n32310), .Z(n31982) );
  AND U31864 ( .A(n691), .B(n32311), .Z(n32310) );
  XOR U31865 ( .A(p_input[4081]), .B(p_input[4049]), .Z(n32311) );
  XNOR U31866 ( .A(n31979), .B(n32306), .Z(n32308) );
  XOR U31867 ( .A(n32312), .B(n32313), .Z(n31979) );
  AND U31868 ( .A(n689), .B(n32314), .Z(n32313) );
  XOR U31869 ( .A(p_input[4017]), .B(p_input[3985]), .Z(n32314) );
  XOR U31870 ( .A(n32315), .B(n32316), .Z(n32306) );
  AND U31871 ( .A(n32317), .B(n32318), .Z(n32316) );
  XOR U31872 ( .A(n32315), .B(n31994), .Z(n32318) );
  XNOR U31873 ( .A(p_input[4048]), .B(n32319), .Z(n31994) );
  AND U31874 ( .A(n691), .B(n32320), .Z(n32319) );
  XOR U31875 ( .A(p_input[4080]), .B(p_input[4048]), .Z(n32320) );
  XNOR U31876 ( .A(n31991), .B(n32315), .Z(n32317) );
  XOR U31877 ( .A(n32321), .B(n32322), .Z(n31991) );
  AND U31878 ( .A(n689), .B(n32323), .Z(n32322) );
  XOR U31879 ( .A(p_input[4016]), .B(p_input[3984]), .Z(n32323) );
  XOR U31880 ( .A(n32324), .B(n32325), .Z(n32315) );
  AND U31881 ( .A(n32326), .B(n32327), .Z(n32325) );
  XOR U31882 ( .A(n32324), .B(n32006), .Z(n32327) );
  XNOR U31883 ( .A(p_input[4047]), .B(n32328), .Z(n32006) );
  AND U31884 ( .A(n691), .B(n32329), .Z(n32328) );
  XOR U31885 ( .A(p_input[4079]), .B(p_input[4047]), .Z(n32329) );
  XNOR U31886 ( .A(n32003), .B(n32324), .Z(n32326) );
  XOR U31887 ( .A(n32330), .B(n32331), .Z(n32003) );
  AND U31888 ( .A(n689), .B(n32332), .Z(n32331) );
  XOR U31889 ( .A(p_input[4015]), .B(p_input[3983]), .Z(n32332) );
  XOR U31890 ( .A(n32333), .B(n32334), .Z(n32324) );
  AND U31891 ( .A(n32335), .B(n32336), .Z(n32334) );
  XOR U31892 ( .A(n32333), .B(n32018), .Z(n32336) );
  XNOR U31893 ( .A(p_input[4046]), .B(n32337), .Z(n32018) );
  AND U31894 ( .A(n691), .B(n32338), .Z(n32337) );
  XOR U31895 ( .A(p_input[4078]), .B(p_input[4046]), .Z(n32338) );
  XNOR U31896 ( .A(n32015), .B(n32333), .Z(n32335) );
  XOR U31897 ( .A(n32339), .B(n32340), .Z(n32015) );
  AND U31898 ( .A(n689), .B(n32341), .Z(n32340) );
  XOR U31899 ( .A(p_input[4014]), .B(p_input[3982]), .Z(n32341) );
  XOR U31900 ( .A(n32342), .B(n32343), .Z(n32333) );
  AND U31901 ( .A(n32344), .B(n32345), .Z(n32343) );
  XOR U31902 ( .A(n32342), .B(n32030), .Z(n32345) );
  XNOR U31903 ( .A(p_input[4045]), .B(n32346), .Z(n32030) );
  AND U31904 ( .A(n691), .B(n32347), .Z(n32346) );
  XOR U31905 ( .A(p_input[4077]), .B(p_input[4045]), .Z(n32347) );
  XNOR U31906 ( .A(n32027), .B(n32342), .Z(n32344) );
  XOR U31907 ( .A(n32348), .B(n32349), .Z(n32027) );
  AND U31908 ( .A(n689), .B(n32350), .Z(n32349) );
  XOR U31909 ( .A(p_input[4013]), .B(p_input[3981]), .Z(n32350) );
  XOR U31910 ( .A(n32351), .B(n32352), .Z(n32342) );
  AND U31911 ( .A(n32353), .B(n32354), .Z(n32352) );
  XOR U31912 ( .A(n32351), .B(n32042), .Z(n32354) );
  XNOR U31913 ( .A(p_input[4044]), .B(n32355), .Z(n32042) );
  AND U31914 ( .A(n691), .B(n32356), .Z(n32355) );
  XOR U31915 ( .A(p_input[4076]), .B(p_input[4044]), .Z(n32356) );
  XNOR U31916 ( .A(n32039), .B(n32351), .Z(n32353) );
  XOR U31917 ( .A(n32357), .B(n32358), .Z(n32039) );
  AND U31918 ( .A(n689), .B(n32359), .Z(n32358) );
  XOR U31919 ( .A(p_input[4012]), .B(p_input[3980]), .Z(n32359) );
  XOR U31920 ( .A(n32360), .B(n32361), .Z(n32351) );
  AND U31921 ( .A(n32362), .B(n32363), .Z(n32361) );
  XOR U31922 ( .A(n32360), .B(n32054), .Z(n32363) );
  XNOR U31923 ( .A(p_input[4043]), .B(n32364), .Z(n32054) );
  AND U31924 ( .A(n691), .B(n32365), .Z(n32364) );
  XOR U31925 ( .A(p_input[4075]), .B(p_input[4043]), .Z(n32365) );
  XNOR U31926 ( .A(n32051), .B(n32360), .Z(n32362) );
  XOR U31927 ( .A(n32366), .B(n32367), .Z(n32051) );
  AND U31928 ( .A(n689), .B(n32368), .Z(n32367) );
  XOR U31929 ( .A(p_input[4011]), .B(p_input[3979]), .Z(n32368) );
  XOR U31930 ( .A(n32369), .B(n32370), .Z(n32360) );
  AND U31931 ( .A(n32371), .B(n32372), .Z(n32370) );
  XOR U31932 ( .A(n32369), .B(n32066), .Z(n32372) );
  XNOR U31933 ( .A(p_input[4042]), .B(n32373), .Z(n32066) );
  AND U31934 ( .A(n691), .B(n32374), .Z(n32373) );
  XOR U31935 ( .A(p_input[4074]), .B(p_input[4042]), .Z(n32374) );
  XNOR U31936 ( .A(n32063), .B(n32369), .Z(n32371) );
  XOR U31937 ( .A(n32375), .B(n32376), .Z(n32063) );
  AND U31938 ( .A(n689), .B(n32377), .Z(n32376) );
  XOR U31939 ( .A(p_input[4010]), .B(p_input[3978]), .Z(n32377) );
  XOR U31940 ( .A(n32378), .B(n32379), .Z(n32369) );
  AND U31941 ( .A(n32380), .B(n32381), .Z(n32379) );
  XOR U31942 ( .A(n32378), .B(n32078), .Z(n32381) );
  XNOR U31943 ( .A(p_input[4041]), .B(n32382), .Z(n32078) );
  AND U31944 ( .A(n691), .B(n32383), .Z(n32382) );
  XOR U31945 ( .A(p_input[4073]), .B(p_input[4041]), .Z(n32383) );
  XNOR U31946 ( .A(n32075), .B(n32378), .Z(n32380) );
  XOR U31947 ( .A(n32384), .B(n32385), .Z(n32075) );
  AND U31948 ( .A(n689), .B(n32386), .Z(n32385) );
  XOR U31949 ( .A(p_input[4009]), .B(p_input[3977]), .Z(n32386) );
  XOR U31950 ( .A(n32387), .B(n32388), .Z(n32378) );
  AND U31951 ( .A(n32389), .B(n32390), .Z(n32388) );
  XOR U31952 ( .A(n32387), .B(n32090), .Z(n32390) );
  XNOR U31953 ( .A(p_input[4040]), .B(n32391), .Z(n32090) );
  AND U31954 ( .A(n691), .B(n32392), .Z(n32391) );
  XOR U31955 ( .A(p_input[4072]), .B(p_input[4040]), .Z(n32392) );
  XNOR U31956 ( .A(n32087), .B(n32387), .Z(n32389) );
  XOR U31957 ( .A(n32393), .B(n32394), .Z(n32087) );
  AND U31958 ( .A(n689), .B(n32395), .Z(n32394) );
  XOR U31959 ( .A(p_input[4008]), .B(p_input[3976]), .Z(n32395) );
  XOR U31960 ( .A(n32396), .B(n32397), .Z(n32387) );
  AND U31961 ( .A(n32398), .B(n32399), .Z(n32397) );
  XOR U31962 ( .A(n32396), .B(n32102), .Z(n32399) );
  XNOR U31963 ( .A(p_input[4039]), .B(n32400), .Z(n32102) );
  AND U31964 ( .A(n691), .B(n32401), .Z(n32400) );
  XOR U31965 ( .A(p_input[4071]), .B(p_input[4039]), .Z(n32401) );
  XNOR U31966 ( .A(n32099), .B(n32396), .Z(n32398) );
  XOR U31967 ( .A(n32402), .B(n32403), .Z(n32099) );
  AND U31968 ( .A(n689), .B(n32404), .Z(n32403) );
  XOR U31969 ( .A(p_input[4007]), .B(p_input[3975]), .Z(n32404) );
  XOR U31970 ( .A(n32405), .B(n32406), .Z(n32396) );
  AND U31971 ( .A(n32407), .B(n32408), .Z(n32406) );
  XOR U31972 ( .A(n32405), .B(n32114), .Z(n32408) );
  XNOR U31973 ( .A(p_input[4038]), .B(n32409), .Z(n32114) );
  AND U31974 ( .A(n691), .B(n32410), .Z(n32409) );
  XOR U31975 ( .A(p_input[4070]), .B(p_input[4038]), .Z(n32410) );
  XNOR U31976 ( .A(n32111), .B(n32405), .Z(n32407) );
  XOR U31977 ( .A(n32411), .B(n32412), .Z(n32111) );
  AND U31978 ( .A(n689), .B(n32413), .Z(n32412) );
  XOR U31979 ( .A(p_input[4006]), .B(p_input[3974]), .Z(n32413) );
  XOR U31980 ( .A(n32414), .B(n32415), .Z(n32405) );
  AND U31981 ( .A(n32416), .B(n32417), .Z(n32415) );
  XOR U31982 ( .A(n32414), .B(n32126), .Z(n32417) );
  XNOR U31983 ( .A(p_input[4037]), .B(n32418), .Z(n32126) );
  AND U31984 ( .A(n691), .B(n32419), .Z(n32418) );
  XOR U31985 ( .A(p_input[4069]), .B(p_input[4037]), .Z(n32419) );
  XNOR U31986 ( .A(n32123), .B(n32414), .Z(n32416) );
  XOR U31987 ( .A(n32420), .B(n32421), .Z(n32123) );
  AND U31988 ( .A(n689), .B(n32422), .Z(n32421) );
  XOR U31989 ( .A(p_input[4005]), .B(p_input[3973]), .Z(n32422) );
  XOR U31990 ( .A(n32423), .B(n32424), .Z(n32414) );
  AND U31991 ( .A(n32425), .B(n32426), .Z(n32424) );
  XOR U31992 ( .A(n32423), .B(n32138), .Z(n32426) );
  XNOR U31993 ( .A(p_input[4036]), .B(n32427), .Z(n32138) );
  AND U31994 ( .A(n691), .B(n32428), .Z(n32427) );
  XOR U31995 ( .A(p_input[4068]), .B(p_input[4036]), .Z(n32428) );
  XNOR U31996 ( .A(n32135), .B(n32423), .Z(n32425) );
  XOR U31997 ( .A(n32429), .B(n32430), .Z(n32135) );
  AND U31998 ( .A(n689), .B(n32431), .Z(n32430) );
  XOR U31999 ( .A(p_input[4004]), .B(p_input[3972]), .Z(n32431) );
  XOR U32000 ( .A(n32432), .B(n32433), .Z(n32423) );
  AND U32001 ( .A(n32434), .B(n32435), .Z(n32433) );
  XOR U32002 ( .A(n32432), .B(n32150), .Z(n32435) );
  XNOR U32003 ( .A(p_input[4035]), .B(n32436), .Z(n32150) );
  AND U32004 ( .A(n691), .B(n32437), .Z(n32436) );
  XOR U32005 ( .A(p_input[4067]), .B(p_input[4035]), .Z(n32437) );
  XNOR U32006 ( .A(n32147), .B(n32432), .Z(n32434) );
  XOR U32007 ( .A(n32438), .B(n32439), .Z(n32147) );
  AND U32008 ( .A(n689), .B(n32440), .Z(n32439) );
  XOR U32009 ( .A(p_input[4003]), .B(p_input[3971]), .Z(n32440) );
  XOR U32010 ( .A(n32441), .B(n32442), .Z(n32432) );
  AND U32011 ( .A(n32443), .B(n32444), .Z(n32442) );
  XOR U32012 ( .A(n32441), .B(n32162), .Z(n32444) );
  XNOR U32013 ( .A(p_input[4034]), .B(n32445), .Z(n32162) );
  AND U32014 ( .A(n691), .B(n32446), .Z(n32445) );
  XOR U32015 ( .A(p_input[4066]), .B(p_input[4034]), .Z(n32446) );
  XNOR U32016 ( .A(n32159), .B(n32441), .Z(n32443) );
  XOR U32017 ( .A(n32447), .B(n32448), .Z(n32159) );
  AND U32018 ( .A(n689), .B(n32449), .Z(n32448) );
  XOR U32019 ( .A(p_input[4002]), .B(p_input[3970]), .Z(n32449) );
  XOR U32020 ( .A(n32450), .B(n32451), .Z(n32441) );
  AND U32021 ( .A(n32452), .B(n32453), .Z(n32451) );
  XNOR U32022 ( .A(n32454), .B(n32175), .Z(n32453) );
  XNOR U32023 ( .A(p_input[4033]), .B(n32455), .Z(n32175) );
  AND U32024 ( .A(n691), .B(n32456), .Z(n32455) );
  XNOR U32025 ( .A(p_input[4065]), .B(n32457), .Z(n32456) );
  IV U32026 ( .A(p_input[4033]), .Z(n32457) );
  XNOR U32027 ( .A(n32172), .B(n32450), .Z(n32452) );
  XNOR U32028 ( .A(p_input[3969]), .B(n32458), .Z(n32172) );
  AND U32029 ( .A(n689), .B(n32459), .Z(n32458) );
  XOR U32030 ( .A(p_input[4001]), .B(p_input[3969]), .Z(n32459) );
  IV U32031 ( .A(n32454), .Z(n32450) );
  AND U32032 ( .A(n32180), .B(n32183), .Z(n32454) );
  XOR U32033 ( .A(p_input[4032]), .B(n32460), .Z(n32183) );
  AND U32034 ( .A(n691), .B(n32461), .Z(n32460) );
  XOR U32035 ( .A(p_input[4064]), .B(p_input[4032]), .Z(n32461) );
  XOR U32036 ( .A(n32462), .B(n32463), .Z(n691) );
  AND U32037 ( .A(n32464), .B(n32465), .Z(n32463) );
  XNOR U32038 ( .A(p_input[4095]), .B(n32462), .Z(n32465) );
  XOR U32039 ( .A(n32462), .B(p_input[4063]), .Z(n32464) );
  XOR U32040 ( .A(n32466), .B(n32467), .Z(n32462) );
  AND U32041 ( .A(n32468), .B(n32469), .Z(n32467) );
  XNOR U32042 ( .A(p_input[4094]), .B(n32466), .Z(n32469) );
  XOR U32043 ( .A(n32466), .B(p_input[4062]), .Z(n32468) );
  XOR U32044 ( .A(n32470), .B(n32471), .Z(n32466) );
  AND U32045 ( .A(n32472), .B(n32473), .Z(n32471) );
  XNOR U32046 ( .A(p_input[4093]), .B(n32470), .Z(n32473) );
  XOR U32047 ( .A(n32470), .B(p_input[4061]), .Z(n32472) );
  XOR U32048 ( .A(n32474), .B(n32475), .Z(n32470) );
  AND U32049 ( .A(n32476), .B(n32477), .Z(n32475) );
  XNOR U32050 ( .A(p_input[4092]), .B(n32474), .Z(n32477) );
  XOR U32051 ( .A(n32474), .B(p_input[4060]), .Z(n32476) );
  XOR U32052 ( .A(n32478), .B(n32479), .Z(n32474) );
  AND U32053 ( .A(n32480), .B(n32481), .Z(n32479) );
  XNOR U32054 ( .A(p_input[4091]), .B(n32478), .Z(n32481) );
  XOR U32055 ( .A(n32478), .B(p_input[4059]), .Z(n32480) );
  XOR U32056 ( .A(n32482), .B(n32483), .Z(n32478) );
  AND U32057 ( .A(n32484), .B(n32485), .Z(n32483) );
  XNOR U32058 ( .A(p_input[4090]), .B(n32482), .Z(n32485) );
  XOR U32059 ( .A(n32482), .B(p_input[4058]), .Z(n32484) );
  XOR U32060 ( .A(n32486), .B(n32487), .Z(n32482) );
  AND U32061 ( .A(n32488), .B(n32489), .Z(n32487) );
  XNOR U32062 ( .A(p_input[4089]), .B(n32486), .Z(n32489) );
  XOR U32063 ( .A(n32486), .B(p_input[4057]), .Z(n32488) );
  XOR U32064 ( .A(n32490), .B(n32491), .Z(n32486) );
  AND U32065 ( .A(n32492), .B(n32493), .Z(n32491) );
  XNOR U32066 ( .A(p_input[4088]), .B(n32490), .Z(n32493) );
  XOR U32067 ( .A(n32490), .B(p_input[4056]), .Z(n32492) );
  XOR U32068 ( .A(n32494), .B(n32495), .Z(n32490) );
  AND U32069 ( .A(n32496), .B(n32497), .Z(n32495) );
  XNOR U32070 ( .A(p_input[4087]), .B(n32494), .Z(n32497) );
  XOR U32071 ( .A(n32494), .B(p_input[4055]), .Z(n32496) );
  XOR U32072 ( .A(n32498), .B(n32499), .Z(n32494) );
  AND U32073 ( .A(n32500), .B(n32501), .Z(n32499) );
  XNOR U32074 ( .A(p_input[4086]), .B(n32498), .Z(n32501) );
  XOR U32075 ( .A(n32498), .B(p_input[4054]), .Z(n32500) );
  XOR U32076 ( .A(n32502), .B(n32503), .Z(n32498) );
  AND U32077 ( .A(n32504), .B(n32505), .Z(n32503) );
  XNOR U32078 ( .A(p_input[4085]), .B(n32502), .Z(n32505) );
  XOR U32079 ( .A(n32502), .B(p_input[4053]), .Z(n32504) );
  XOR U32080 ( .A(n32506), .B(n32507), .Z(n32502) );
  AND U32081 ( .A(n32508), .B(n32509), .Z(n32507) );
  XNOR U32082 ( .A(p_input[4084]), .B(n32506), .Z(n32509) );
  XOR U32083 ( .A(n32506), .B(p_input[4052]), .Z(n32508) );
  XOR U32084 ( .A(n32510), .B(n32511), .Z(n32506) );
  AND U32085 ( .A(n32512), .B(n32513), .Z(n32511) );
  XNOR U32086 ( .A(p_input[4083]), .B(n32510), .Z(n32513) );
  XOR U32087 ( .A(n32510), .B(p_input[4051]), .Z(n32512) );
  XOR U32088 ( .A(n32514), .B(n32515), .Z(n32510) );
  AND U32089 ( .A(n32516), .B(n32517), .Z(n32515) );
  XNOR U32090 ( .A(p_input[4082]), .B(n32514), .Z(n32517) );
  XOR U32091 ( .A(n32514), .B(p_input[4050]), .Z(n32516) );
  XOR U32092 ( .A(n32518), .B(n32519), .Z(n32514) );
  AND U32093 ( .A(n32520), .B(n32521), .Z(n32519) );
  XNOR U32094 ( .A(p_input[4081]), .B(n32518), .Z(n32521) );
  XOR U32095 ( .A(n32518), .B(p_input[4049]), .Z(n32520) );
  XOR U32096 ( .A(n32522), .B(n32523), .Z(n32518) );
  AND U32097 ( .A(n32524), .B(n32525), .Z(n32523) );
  XNOR U32098 ( .A(p_input[4080]), .B(n32522), .Z(n32525) );
  XOR U32099 ( .A(n32522), .B(p_input[4048]), .Z(n32524) );
  XOR U32100 ( .A(n32526), .B(n32527), .Z(n32522) );
  AND U32101 ( .A(n32528), .B(n32529), .Z(n32527) );
  XNOR U32102 ( .A(p_input[4079]), .B(n32526), .Z(n32529) );
  XOR U32103 ( .A(n32526), .B(p_input[4047]), .Z(n32528) );
  XOR U32104 ( .A(n32530), .B(n32531), .Z(n32526) );
  AND U32105 ( .A(n32532), .B(n32533), .Z(n32531) );
  XNOR U32106 ( .A(p_input[4078]), .B(n32530), .Z(n32533) );
  XOR U32107 ( .A(n32530), .B(p_input[4046]), .Z(n32532) );
  XOR U32108 ( .A(n32534), .B(n32535), .Z(n32530) );
  AND U32109 ( .A(n32536), .B(n32537), .Z(n32535) );
  XNOR U32110 ( .A(p_input[4077]), .B(n32534), .Z(n32537) );
  XOR U32111 ( .A(n32534), .B(p_input[4045]), .Z(n32536) );
  XOR U32112 ( .A(n32538), .B(n32539), .Z(n32534) );
  AND U32113 ( .A(n32540), .B(n32541), .Z(n32539) );
  XNOR U32114 ( .A(p_input[4076]), .B(n32538), .Z(n32541) );
  XOR U32115 ( .A(n32538), .B(p_input[4044]), .Z(n32540) );
  XOR U32116 ( .A(n32542), .B(n32543), .Z(n32538) );
  AND U32117 ( .A(n32544), .B(n32545), .Z(n32543) );
  XNOR U32118 ( .A(p_input[4075]), .B(n32542), .Z(n32545) );
  XOR U32119 ( .A(n32542), .B(p_input[4043]), .Z(n32544) );
  XOR U32120 ( .A(n32546), .B(n32547), .Z(n32542) );
  AND U32121 ( .A(n32548), .B(n32549), .Z(n32547) );
  XNOR U32122 ( .A(p_input[4074]), .B(n32546), .Z(n32549) );
  XOR U32123 ( .A(n32546), .B(p_input[4042]), .Z(n32548) );
  XOR U32124 ( .A(n32550), .B(n32551), .Z(n32546) );
  AND U32125 ( .A(n32552), .B(n32553), .Z(n32551) );
  XNOR U32126 ( .A(p_input[4073]), .B(n32550), .Z(n32553) );
  XOR U32127 ( .A(n32550), .B(p_input[4041]), .Z(n32552) );
  XOR U32128 ( .A(n32554), .B(n32555), .Z(n32550) );
  AND U32129 ( .A(n32556), .B(n32557), .Z(n32555) );
  XNOR U32130 ( .A(p_input[4072]), .B(n32554), .Z(n32557) );
  XOR U32131 ( .A(n32554), .B(p_input[4040]), .Z(n32556) );
  XOR U32132 ( .A(n32558), .B(n32559), .Z(n32554) );
  AND U32133 ( .A(n32560), .B(n32561), .Z(n32559) );
  XNOR U32134 ( .A(p_input[4071]), .B(n32558), .Z(n32561) );
  XOR U32135 ( .A(n32558), .B(p_input[4039]), .Z(n32560) );
  XOR U32136 ( .A(n32562), .B(n32563), .Z(n32558) );
  AND U32137 ( .A(n32564), .B(n32565), .Z(n32563) );
  XNOR U32138 ( .A(p_input[4070]), .B(n32562), .Z(n32565) );
  XOR U32139 ( .A(n32562), .B(p_input[4038]), .Z(n32564) );
  XOR U32140 ( .A(n32566), .B(n32567), .Z(n32562) );
  AND U32141 ( .A(n32568), .B(n32569), .Z(n32567) );
  XNOR U32142 ( .A(p_input[4069]), .B(n32566), .Z(n32569) );
  XOR U32143 ( .A(n32566), .B(p_input[4037]), .Z(n32568) );
  XOR U32144 ( .A(n32570), .B(n32571), .Z(n32566) );
  AND U32145 ( .A(n32572), .B(n32573), .Z(n32571) );
  XNOR U32146 ( .A(p_input[4068]), .B(n32570), .Z(n32573) );
  XOR U32147 ( .A(n32570), .B(p_input[4036]), .Z(n32572) );
  XOR U32148 ( .A(n32574), .B(n32575), .Z(n32570) );
  AND U32149 ( .A(n32576), .B(n32577), .Z(n32575) );
  XNOR U32150 ( .A(p_input[4067]), .B(n32574), .Z(n32577) );
  XOR U32151 ( .A(n32574), .B(p_input[4035]), .Z(n32576) );
  XOR U32152 ( .A(n32578), .B(n32579), .Z(n32574) );
  AND U32153 ( .A(n32580), .B(n32581), .Z(n32579) );
  XNOR U32154 ( .A(p_input[4066]), .B(n32578), .Z(n32581) );
  XOR U32155 ( .A(n32578), .B(p_input[4034]), .Z(n32580) );
  XNOR U32156 ( .A(n32582), .B(n32583), .Z(n32578) );
  AND U32157 ( .A(n32584), .B(n32585), .Z(n32583) );
  XOR U32158 ( .A(p_input[4065]), .B(n32582), .Z(n32585) );
  XNOR U32159 ( .A(p_input[4033]), .B(n32582), .Z(n32584) );
  AND U32160 ( .A(p_input[4064]), .B(n32586), .Z(n32582) );
  IV U32161 ( .A(p_input[4032]), .Z(n32586) );
  XNOR U32162 ( .A(p_input[3968]), .B(n32587), .Z(n32180) );
  AND U32163 ( .A(n689), .B(n32588), .Z(n32587) );
  XOR U32164 ( .A(p_input[4000]), .B(p_input[3968]), .Z(n32588) );
  XOR U32165 ( .A(n32589), .B(n32590), .Z(n689) );
  AND U32166 ( .A(n32591), .B(n32592), .Z(n32590) );
  XNOR U32167 ( .A(p_input[4031]), .B(n32589), .Z(n32592) );
  XOR U32168 ( .A(n32589), .B(p_input[3999]), .Z(n32591) );
  XOR U32169 ( .A(n32593), .B(n32594), .Z(n32589) );
  AND U32170 ( .A(n32595), .B(n32596), .Z(n32594) );
  XNOR U32171 ( .A(p_input[4030]), .B(n32593), .Z(n32596) );
  XNOR U32172 ( .A(n32593), .B(n32195), .Z(n32595) );
  IV U32173 ( .A(p_input[3998]), .Z(n32195) );
  XOR U32174 ( .A(n32597), .B(n32598), .Z(n32593) );
  AND U32175 ( .A(n32599), .B(n32600), .Z(n32598) );
  XNOR U32176 ( .A(p_input[4029]), .B(n32597), .Z(n32600) );
  XNOR U32177 ( .A(n32597), .B(n32204), .Z(n32599) );
  IV U32178 ( .A(p_input[3997]), .Z(n32204) );
  XOR U32179 ( .A(n32601), .B(n32602), .Z(n32597) );
  AND U32180 ( .A(n32603), .B(n32604), .Z(n32602) );
  XNOR U32181 ( .A(p_input[4028]), .B(n32601), .Z(n32604) );
  XNOR U32182 ( .A(n32601), .B(n32213), .Z(n32603) );
  IV U32183 ( .A(p_input[3996]), .Z(n32213) );
  XOR U32184 ( .A(n32605), .B(n32606), .Z(n32601) );
  AND U32185 ( .A(n32607), .B(n32608), .Z(n32606) );
  XNOR U32186 ( .A(p_input[4027]), .B(n32605), .Z(n32608) );
  XNOR U32187 ( .A(n32605), .B(n32222), .Z(n32607) );
  IV U32188 ( .A(p_input[3995]), .Z(n32222) );
  XOR U32189 ( .A(n32609), .B(n32610), .Z(n32605) );
  AND U32190 ( .A(n32611), .B(n32612), .Z(n32610) );
  XNOR U32191 ( .A(p_input[4026]), .B(n32609), .Z(n32612) );
  XNOR U32192 ( .A(n32609), .B(n32231), .Z(n32611) );
  IV U32193 ( .A(p_input[3994]), .Z(n32231) );
  XOR U32194 ( .A(n32613), .B(n32614), .Z(n32609) );
  AND U32195 ( .A(n32615), .B(n32616), .Z(n32614) );
  XNOR U32196 ( .A(p_input[4025]), .B(n32613), .Z(n32616) );
  XNOR U32197 ( .A(n32613), .B(n32240), .Z(n32615) );
  IV U32198 ( .A(p_input[3993]), .Z(n32240) );
  XOR U32199 ( .A(n32617), .B(n32618), .Z(n32613) );
  AND U32200 ( .A(n32619), .B(n32620), .Z(n32618) );
  XNOR U32201 ( .A(p_input[4024]), .B(n32617), .Z(n32620) );
  XNOR U32202 ( .A(n32617), .B(n32249), .Z(n32619) );
  IV U32203 ( .A(p_input[3992]), .Z(n32249) );
  XOR U32204 ( .A(n32621), .B(n32622), .Z(n32617) );
  AND U32205 ( .A(n32623), .B(n32624), .Z(n32622) );
  XNOR U32206 ( .A(p_input[4023]), .B(n32621), .Z(n32624) );
  XNOR U32207 ( .A(n32621), .B(n32258), .Z(n32623) );
  IV U32208 ( .A(p_input[3991]), .Z(n32258) );
  XOR U32209 ( .A(n32625), .B(n32626), .Z(n32621) );
  AND U32210 ( .A(n32627), .B(n32628), .Z(n32626) );
  XNOR U32211 ( .A(p_input[4022]), .B(n32625), .Z(n32628) );
  XNOR U32212 ( .A(n32625), .B(n32267), .Z(n32627) );
  IV U32213 ( .A(p_input[3990]), .Z(n32267) );
  XOR U32214 ( .A(n32629), .B(n32630), .Z(n32625) );
  AND U32215 ( .A(n32631), .B(n32632), .Z(n32630) );
  XNOR U32216 ( .A(p_input[4021]), .B(n32629), .Z(n32632) );
  XNOR U32217 ( .A(n32629), .B(n32276), .Z(n32631) );
  IV U32218 ( .A(p_input[3989]), .Z(n32276) );
  XOR U32219 ( .A(n32633), .B(n32634), .Z(n32629) );
  AND U32220 ( .A(n32635), .B(n32636), .Z(n32634) );
  XNOR U32221 ( .A(p_input[4020]), .B(n32633), .Z(n32636) );
  XNOR U32222 ( .A(n32633), .B(n32285), .Z(n32635) );
  IV U32223 ( .A(p_input[3988]), .Z(n32285) );
  XOR U32224 ( .A(n32637), .B(n32638), .Z(n32633) );
  AND U32225 ( .A(n32639), .B(n32640), .Z(n32638) );
  XNOR U32226 ( .A(p_input[4019]), .B(n32637), .Z(n32640) );
  XNOR U32227 ( .A(n32637), .B(n32294), .Z(n32639) );
  IV U32228 ( .A(p_input[3987]), .Z(n32294) );
  XOR U32229 ( .A(n32641), .B(n32642), .Z(n32637) );
  AND U32230 ( .A(n32643), .B(n32644), .Z(n32642) );
  XNOR U32231 ( .A(p_input[4018]), .B(n32641), .Z(n32644) );
  XNOR U32232 ( .A(n32641), .B(n32303), .Z(n32643) );
  IV U32233 ( .A(p_input[3986]), .Z(n32303) );
  XOR U32234 ( .A(n32645), .B(n32646), .Z(n32641) );
  AND U32235 ( .A(n32647), .B(n32648), .Z(n32646) );
  XNOR U32236 ( .A(p_input[4017]), .B(n32645), .Z(n32648) );
  XNOR U32237 ( .A(n32645), .B(n32312), .Z(n32647) );
  IV U32238 ( .A(p_input[3985]), .Z(n32312) );
  XOR U32239 ( .A(n32649), .B(n32650), .Z(n32645) );
  AND U32240 ( .A(n32651), .B(n32652), .Z(n32650) );
  XNOR U32241 ( .A(p_input[4016]), .B(n32649), .Z(n32652) );
  XNOR U32242 ( .A(n32649), .B(n32321), .Z(n32651) );
  IV U32243 ( .A(p_input[3984]), .Z(n32321) );
  XOR U32244 ( .A(n32653), .B(n32654), .Z(n32649) );
  AND U32245 ( .A(n32655), .B(n32656), .Z(n32654) );
  XNOR U32246 ( .A(p_input[4015]), .B(n32653), .Z(n32656) );
  XNOR U32247 ( .A(n32653), .B(n32330), .Z(n32655) );
  IV U32248 ( .A(p_input[3983]), .Z(n32330) );
  XOR U32249 ( .A(n32657), .B(n32658), .Z(n32653) );
  AND U32250 ( .A(n32659), .B(n32660), .Z(n32658) );
  XNOR U32251 ( .A(p_input[4014]), .B(n32657), .Z(n32660) );
  XNOR U32252 ( .A(n32657), .B(n32339), .Z(n32659) );
  IV U32253 ( .A(p_input[3982]), .Z(n32339) );
  XOR U32254 ( .A(n32661), .B(n32662), .Z(n32657) );
  AND U32255 ( .A(n32663), .B(n32664), .Z(n32662) );
  XNOR U32256 ( .A(p_input[4013]), .B(n32661), .Z(n32664) );
  XNOR U32257 ( .A(n32661), .B(n32348), .Z(n32663) );
  IV U32258 ( .A(p_input[3981]), .Z(n32348) );
  XOR U32259 ( .A(n32665), .B(n32666), .Z(n32661) );
  AND U32260 ( .A(n32667), .B(n32668), .Z(n32666) );
  XNOR U32261 ( .A(p_input[4012]), .B(n32665), .Z(n32668) );
  XNOR U32262 ( .A(n32665), .B(n32357), .Z(n32667) );
  IV U32263 ( .A(p_input[3980]), .Z(n32357) );
  XOR U32264 ( .A(n32669), .B(n32670), .Z(n32665) );
  AND U32265 ( .A(n32671), .B(n32672), .Z(n32670) );
  XNOR U32266 ( .A(p_input[4011]), .B(n32669), .Z(n32672) );
  XNOR U32267 ( .A(n32669), .B(n32366), .Z(n32671) );
  IV U32268 ( .A(p_input[3979]), .Z(n32366) );
  XOR U32269 ( .A(n32673), .B(n32674), .Z(n32669) );
  AND U32270 ( .A(n32675), .B(n32676), .Z(n32674) );
  XNOR U32271 ( .A(p_input[4010]), .B(n32673), .Z(n32676) );
  XNOR U32272 ( .A(n32673), .B(n32375), .Z(n32675) );
  IV U32273 ( .A(p_input[3978]), .Z(n32375) );
  XOR U32274 ( .A(n32677), .B(n32678), .Z(n32673) );
  AND U32275 ( .A(n32679), .B(n32680), .Z(n32678) );
  XNOR U32276 ( .A(p_input[4009]), .B(n32677), .Z(n32680) );
  XNOR U32277 ( .A(n32677), .B(n32384), .Z(n32679) );
  IV U32278 ( .A(p_input[3977]), .Z(n32384) );
  XOR U32279 ( .A(n32681), .B(n32682), .Z(n32677) );
  AND U32280 ( .A(n32683), .B(n32684), .Z(n32682) );
  XNOR U32281 ( .A(p_input[4008]), .B(n32681), .Z(n32684) );
  XNOR U32282 ( .A(n32681), .B(n32393), .Z(n32683) );
  IV U32283 ( .A(p_input[3976]), .Z(n32393) );
  XOR U32284 ( .A(n32685), .B(n32686), .Z(n32681) );
  AND U32285 ( .A(n32687), .B(n32688), .Z(n32686) );
  XNOR U32286 ( .A(p_input[4007]), .B(n32685), .Z(n32688) );
  XNOR U32287 ( .A(n32685), .B(n32402), .Z(n32687) );
  IV U32288 ( .A(p_input[3975]), .Z(n32402) );
  XOR U32289 ( .A(n32689), .B(n32690), .Z(n32685) );
  AND U32290 ( .A(n32691), .B(n32692), .Z(n32690) );
  XNOR U32291 ( .A(p_input[4006]), .B(n32689), .Z(n32692) );
  XNOR U32292 ( .A(n32689), .B(n32411), .Z(n32691) );
  IV U32293 ( .A(p_input[3974]), .Z(n32411) );
  XOR U32294 ( .A(n32693), .B(n32694), .Z(n32689) );
  AND U32295 ( .A(n32695), .B(n32696), .Z(n32694) );
  XNOR U32296 ( .A(p_input[4005]), .B(n32693), .Z(n32696) );
  XNOR U32297 ( .A(n32693), .B(n32420), .Z(n32695) );
  IV U32298 ( .A(p_input[3973]), .Z(n32420) );
  XOR U32299 ( .A(n32697), .B(n32698), .Z(n32693) );
  AND U32300 ( .A(n32699), .B(n32700), .Z(n32698) );
  XNOR U32301 ( .A(p_input[4004]), .B(n32697), .Z(n32700) );
  XNOR U32302 ( .A(n32697), .B(n32429), .Z(n32699) );
  IV U32303 ( .A(p_input[3972]), .Z(n32429) );
  XOR U32304 ( .A(n32701), .B(n32702), .Z(n32697) );
  AND U32305 ( .A(n32703), .B(n32704), .Z(n32702) );
  XNOR U32306 ( .A(p_input[4003]), .B(n32701), .Z(n32704) );
  XNOR U32307 ( .A(n32701), .B(n32438), .Z(n32703) );
  IV U32308 ( .A(p_input[3971]), .Z(n32438) );
  XOR U32309 ( .A(n32705), .B(n32706), .Z(n32701) );
  AND U32310 ( .A(n32707), .B(n32708), .Z(n32706) );
  XNOR U32311 ( .A(p_input[4002]), .B(n32705), .Z(n32708) );
  XNOR U32312 ( .A(n32705), .B(n32447), .Z(n32707) );
  IV U32313 ( .A(p_input[3970]), .Z(n32447) );
  XNOR U32314 ( .A(n32709), .B(n32710), .Z(n32705) );
  AND U32315 ( .A(n32711), .B(n32712), .Z(n32710) );
  XOR U32316 ( .A(p_input[4001]), .B(n32709), .Z(n32712) );
  XNOR U32317 ( .A(p_input[3969]), .B(n32709), .Z(n32711) );
  AND U32318 ( .A(p_input[4000]), .B(n32713), .Z(n32709) );
  IV U32319 ( .A(p_input[3968]), .Z(n32713) );
  XOR U32320 ( .A(n32714), .B(n32715), .Z(n31803) );
  AND U32321 ( .A(n561), .B(n32716), .Z(n32715) );
  XNOR U32322 ( .A(n32717), .B(n32714), .Z(n32716) );
  XOR U32323 ( .A(n32718), .B(n32719), .Z(n561) );
  AND U32324 ( .A(n32720), .B(n32721), .Z(n32719) );
  XNOR U32325 ( .A(n31818), .B(n32718), .Z(n32721) );
  AND U32326 ( .A(p_input[3967]), .B(p_input[3935]), .Z(n31818) );
  XNOR U32327 ( .A(n32718), .B(n31815), .Z(n32720) );
  IV U32328 ( .A(n32722), .Z(n31815) );
  AND U32329 ( .A(p_input[3871]), .B(p_input[3903]), .Z(n32722) );
  XOR U32330 ( .A(n32723), .B(n32724), .Z(n32718) );
  AND U32331 ( .A(n32725), .B(n32726), .Z(n32724) );
  XOR U32332 ( .A(n32723), .B(n31830), .Z(n32726) );
  XNOR U32333 ( .A(p_input[3934]), .B(n32727), .Z(n31830) );
  AND U32334 ( .A(n695), .B(n32728), .Z(n32727) );
  XOR U32335 ( .A(p_input[3966]), .B(p_input[3934]), .Z(n32728) );
  XNOR U32336 ( .A(n31827), .B(n32723), .Z(n32725) );
  XOR U32337 ( .A(n32729), .B(n32730), .Z(n31827) );
  AND U32338 ( .A(n692), .B(n32731), .Z(n32730) );
  XOR U32339 ( .A(p_input[3902]), .B(p_input[3870]), .Z(n32731) );
  XOR U32340 ( .A(n32732), .B(n32733), .Z(n32723) );
  AND U32341 ( .A(n32734), .B(n32735), .Z(n32733) );
  XOR U32342 ( .A(n32732), .B(n31842), .Z(n32735) );
  XNOR U32343 ( .A(p_input[3933]), .B(n32736), .Z(n31842) );
  AND U32344 ( .A(n695), .B(n32737), .Z(n32736) );
  XOR U32345 ( .A(p_input[3965]), .B(p_input[3933]), .Z(n32737) );
  XNOR U32346 ( .A(n31839), .B(n32732), .Z(n32734) );
  XOR U32347 ( .A(n32738), .B(n32739), .Z(n31839) );
  AND U32348 ( .A(n692), .B(n32740), .Z(n32739) );
  XOR U32349 ( .A(p_input[3901]), .B(p_input[3869]), .Z(n32740) );
  XOR U32350 ( .A(n32741), .B(n32742), .Z(n32732) );
  AND U32351 ( .A(n32743), .B(n32744), .Z(n32742) );
  XOR U32352 ( .A(n32741), .B(n31854), .Z(n32744) );
  XNOR U32353 ( .A(p_input[3932]), .B(n32745), .Z(n31854) );
  AND U32354 ( .A(n695), .B(n32746), .Z(n32745) );
  XOR U32355 ( .A(p_input[3964]), .B(p_input[3932]), .Z(n32746) );
  XNOR U32356 ( .A(n31851), .B(n32741), .Z(n32743) );
  XOR U32357 ( .A(n32747), .B(n32748), .Z(n31851) );
  AND U32358 ( .A(n692), .B(n32749), .Z(n32748) );
  XOR U32359 ( .A(p_input[3900]), .B(p_input[3868]), .Z(n32749) );
  XOR U32360 ( .A(n32750), .B(n32751), .Z(n32741) );
  AND U32361 ( .A(n32752), .B(n32753), .Z(n32751) );
  XOR U32362 ( .A(n32750), .B(n31866), .Z(n32753) );
  XNOR U32363 ( .A(p_input[3931]), .B(n32754), .Z(n31866) );
  AND U32364 ( .A(n695), .B(n32755), .Z(n32754) );
  XOR U32365 ( .A(p_input[3963]), .B(p_input[3931]), .Z(n32755) );
  XNOR U32366 ( .A(n31863), .B(n32750), .Z(n32752) );
  XOR U32367 ( .A(n32756), .B(n32757), .Z(n31863) );
  AND U32368 ( .A(n692), .B(n32758), .Z(n32757) );
  XOR U32369 ( .A(p_input[3899]), .B(p_input[3867]), .Z(n32758) );
  XOR U32370 ( .A(n32759), .B(n32760), .Z(n32750) );
  AND U32371 ( .A(n32761), .B(n32762), .Z(n32760) );
  XOR U32372 ( .A(n32759), .B(n31878), .Z(n32762) );
  XNOR U32373 ( .A(p_input[3930]), .B(n32763), .Z(n31878) );
  AND U32374 ( .A(n695), .B(n32764), .Z(n32763) );
  XOR U32375 ( .A(p_input[3962]), .B(p_input[3930]), .Z(n32764) );
  XNOR U32376 ( .A(n31875), .B(n32759), .Z(n32761) );
  XOR U32377 ( .A(n32765), .B(n32766), .Z(n31875) );
  AND U32378 ( .A(n692), .B(n32767), .Z(n32766) );
  XOR U32379 ( .A(p_input[3898]), .B(p_input[3866]), .Z(n32767) );
  XOR U32380 ( .A(n32768), .B(n32769), .Z(n32759) );
  AND U32381 ( .A(n32770), .B(n32771), .Z(n32769) );
  XOR U32382 ( .A(n32768), .B(n31890), .Z(n32771) );
  XNOR U32383 ( .A(p_input[3929]), .B(n32772), .Z(n31890) );
  AND U32384 ( .A(n695), .B(n32773), .Z(n32772) );
  XOR U32385 ( .A(p_input[3961]), .B(p_input[3929]), .Z(n32773) );
  XNOR U32386 ( .A(n31887), .B(n32768), .Z(n32770) );
  XOR U32387 ( .A(n32774), .B(n32775), .Z(n31887) );
  AND U32388 ( .A(n692), .B(n32776), .Z(n32775) );
  XOR U32389 ( .A(p_input[3897]), .B(p_input[3865]), .Z(n32776) );
  XOR U32390 ( .A(n32777), .B(n32778), .Z(n32768) );
  AND U32391 ( .A(n32779), .B(n32780), .Z(n32778) );
  XOR U32392 ( .A(n32777), .B(n31902), .Z(n32780) );
  XNOR U32393 ( .A(p_input[3928]), .B(n32781), .Z(n31902) );
  AND U32394 ( .A(n695), .B(n32782), .Z(n32781) );
  XOR U32395 ( .A(p_input[3960]), .B(p_input[3928]), .Z(n32782) );
  XNOR U32396 ( .A(n31899), .B(n32777), .Z(n32779) );
  XOR U32397 ( .A(n32783), .B(n32784), .Z(n31899) );
  AND U32398 ( .A(n692), .B(n32785), .Z(n32784) );
  XOR U32399 ( .A(p_input[3896]), .B(p_input[3864]), .Z(n32785) );
  XOR U32400 ( .A(n32786), .B(n32787), .Z(n32777) );
  AND U32401 ( .A(n32788), .B(n32789), .Z(n32787) );
  XOR U32402 ( .A(n32786), .B(n31914), .Z(n32789) );
  XNOR U32403 ( .A(p_input[3927]), .B(n32790), .Z(n31914) );
  AND U32404 ( .A(n695), .B(n32791), .Z(n32790) );
  XOR U32405 ( .A(p_input[3959]), .B(p_input[3927]), .Z(n32791) );
  XNOR U32406 ( .A(n31911), .B(n32786), .Z(n32788) );
  XOR U32407 ( .A(n32792), .B(n32793), .Z(n31911) );
  AND U32408 ( .A(n692), .B(n32794), .Z(n32793) );
  XOR U32409 ( .A(p_input[3895]), .B(p_input[3863]), .Z(n32794) );
  XOR U32410 ( .A(n32795), .B(n32796), .Z(n32786) );
  AND U32411 ( .A(n32797), .B(n32798), .Z(n32796) );
  XOR U32412 ( .A(n32795), .B(n31926), .Z(n32798) );
  XNOR U32413 ( .A(p_input[3926]), .B(n32799), .Z(n31926) );
  AND U32414 ( .A(n695), .B(n32800), .Z(n32799) );
  XOR U32415 ( .A(p_input[3958]), .B(p_input[3926]), .Z(n32800) );
  XNOR U32416 ( .A(n31923), .B(n32795), .Z(n32797) );
  XOR U32417 ( .A(n32801), .B(n32802), .Z(n31923) );
  AND U32418 ( .A(n692), .B(n32803), .Z(n32802) );
  XOR U32419 ( .A(p_input[3894]), .B(p_input[3862]), .Z(n32803) );
  XOR U32420 ( .A(n32804), .B(n32805), .Z(n32795) );
  AND U32421 ( .A(n32806), .B(n32807), .Z(n32805) );
  XOR U32422 ( .A(n32804), .B(n31938), .Z(n32807) );
  XNOR U32423 ( .A(p_input[3925]), .B(n32808), .Z(n31938) );
  AND U32424 ( .A(n695), .B(n32809), .Z(n32808) );
  XOR U32425 ( .A(p_input[3957]), .B(p_input[3925]), .Z(n32809) );
  XNOR U32426 ( .A(n31935), .B(n32804), .Z(n32806) );
  XOR U32427 ( .A(n32810), .B(n32811), .Z(n31935) );
  AND U32428 ( .A(n692), .B(n32812), .Z(n32811) );
  XOR U32429 ( .A(p_input[3893]), .B(p_input[3861]), .Z(n32812) );
  XOR U32430 ( .A(n32813), .B(n32814), .Z(n32804) );
  AND U32431 ( .A(n32815), .B(n32816), .Z(n32814) );
  XOR U32432 ( .A(n32813), .B(n31950), .Z(n32816) );
  XNOR U32433 ( .A(p_input[3924]), .B(n32817), .Z(n31950) );
  AND U32434 ( .A(n695), .B(n32818), .Z(n32817) );
  XOR U32435 ( .A(p_input[3956]), .B(p_input[3924]), .Z(n32818) );
  XNOR U32436 ( .A(n31947), .B(n32813), .Z(n32815) );
  XOR U32437 ( .A(n32819), .B(n32820), .Z(n31947) );
  AND U32438 ( .A(n692), .B(n32821), .Z(n32820) );
  XOR U32439 ( .A(p_input[3892]), .B(p_input[3860]), .Z(n32821) );
  XOR U32440 ( .A(n32822), .B(n32823), .Z(n32813) );
  AND U32441 ( .A(n32824), .B(n32825), .Z(n32823) );
  XOR U32442 ( .A(n32822), .B(n31962), .Z(n32825) );
  XNOR U32443 ( .A(p_input[3923]), .B(n32826), .Z(n31962) );
  AND U32444 ( .A(n695), .B(n32827), .Z(n32826) );
  XOR U32445 ( .A(p_input[3955]), .B(p_input[3923]), .Z(n32827) );
  XNOR U32446 ( .A(n31959), .B(n32822), .Z(n32824) );
  XOR U32447 ( .A(n32828), .B(n32829), .Z(n31959) );
  AND U32448 ( .A(n692), .B(n32830), .Z(n32829) );
  XOR U32449 ( .A(p_input[3891]), .B(p_input[3859]), .Z(n32830) );
  XOR U32450 ( .A(n32831), .B(n32832), .Z(n32822) );
  AND U32451 ( .A(n32833), .B(n32834), .Z(n32832) );
  XOR U32452 ( .A(n32831), .B(n31974), .Z(n32834) );
  XNOR U32453 ( .A(p_input[3922]), .B(n32835), .Z(n31974) );
  AND U32454 ( .A(n695), .B(n32836), .Z(n32835) );
  XOR U32455 ( .A(p_input[3954]), .B(p_input[3922]), .Z(n32836) );
  XNOR U32456 ( .A(n31971), .B(n32831), .Z(n32833) );
  XOR U32457 ( .A(n32837), .B(n32838), .Z(n31971) );
  AND U32458 ( .A(n692), .B(n32839), .Z(n32838) );
  XOR U32459 ( .A(p_input[3890]), .B(p_input[3858]), .Z(n32839) );
  XOR U32460 ( .A(n32840), .B(n32841), .Z(n32831) );
  AND U32461 ( .A(n32842), .B(n32843), .Z(n32841) );
  XOR U32462 ( .A(n32840), .B(n31986), .Z(n32843) );
  XNOR U32463 ( .A(p_input[3921]), .B(n32844), .Z(n31986) );
  AND U32464 ( .A(n695), .B(n32845), .Z(n32844) );
  XOR U32465 ( .A(p_input[3953]), .B(p_input[3921]), .Z(n32845) );
  XNOR U32466 ( .A(n31983), .B(n32840), .Z(n32842) );
  XOR U32467 ( .A(n32846), .B(n32847), .Z(n31983) );
  AND U32468 ( .A(n692), .B(n32848), .Z(n32847) );
  XOR U32469 ( .A(p_input[3889]), .B(p_input[3857]), .Z(n32848) );
  XOR U32470 ( .A(n32849), .B(n32850), .Z(n32840) );
  AND U32471 ( .A(n32851), .B(n32852), .Z(n32850) );
  XOR U32472 ( .A(n32849), .B(n31998), .Z(n32852) );
  XNOR U32473 ( .A(p_input[3920]), .B(n32853), .Z(n31998) );
  AND U32474 ( .A(n695), .B(n32854), .Z(n32853) );
  XOR U32475 ( .A(p_input[3952]), .B(p_input[3920]), .Z(n32854) );
  XNOR U32476 ( .A(n31995), .B(n32849), .Z(n32851) );
  XOR U32477 ( .A(n32855), .B(n32856), .Z(n31995) );
  AND U32478 ( .A(n692), .B(n32857), .Z(n32856) );
  XOR U32479 ( .A(p_input[3888]), .B(p_input[3856]), .Z(n32857) );
  XOR U32480 ( .A(n32858), .B(n32859), .Z(n32849) );
  AND U32481 ( .A(n32860), .B(n32861), .Z(n32859) );
  XOR U32482 ( .A(n32858), .B(n32010), .Z(n32861) );
  XNOR U32483 ( .A(p_input[3919]), .B(n32862), .Z(n32010) );
  AND U32484 ( .A(n695), .B(n32863), .Z(n32862) );
  XOR U32485 ( .A(p_input[3951]), .B(p_input[3919]), .Z(n32863) );
  XNOR U32486 ( .A(n32007), .B(n32858), .Z(n32860) );
  XOR U32487 ( .A(n32864), .B(n32865), .Z(n32007) );
  AND U32488 ( .A(n692), .B(n32866), .Z(n32865) );
  XOR U32489 ( .A(p_input[3887]), .B(p_input[3855]), .Z(n32866) );
  XOR U32490 ( .A(n32867), .B(n32868), .Z(n32858) );
  AND U32491 ( .A(n32869), .B(n32870), .Z(n32868) );
  XOR U32492 ( .A(n32867), .B(n32022), .Z(n32870) );
  XNOR U32493 ( .A(p_input[3918]), .B(n32871), .Z(n32022) );
  AND U32494 ( .A(n695), .B(n32872), .Z(n32871) );
  XOR U32495 ( .A(p_input[3950]), .B(p_input[3918]), .Z(n32872) );
  XNOR U32496 ( .A(n32019), .B(n32867), .Z(n32869) );
  XOR U32497 ( .A(n32873), .B(n32874), .Z(n32019) );
  AND U32498 ( .A(n692), .B(n32875), .Z(n32874) );
  XOR U32499 ( .A(p_input[3886]), .B(p_input[3854]), .Z(n32875) );
  XOR U32500 ( .A(n32876), .B(n32877), .Z(n32867) );
  AND U32501 ( .A(n32878), .B(n32879), .Z(n32877) );
  XOR U32502 ( .A(n32876), .B(n32034), .Z(n32879) );
  XNOR U32503 ( .A(p_input[3917]), .B(n32880), .Z(n32034) );
  AND U32504 ( .A(n695), .B(n32881), .Z(n32880) );
  XOR U32505 ( .A(p_input[3949]), .B(p_input[3917]), .Z(n32881) );
  XNOR U32506 ( .A(n32031), .B(n32876), .Z(n32878) );
  XOR U32507 ( .A(n32882), .B(n32883), .Z(n32031) );
  AND U32508 ( .A(n692), .B(n32884), .Z(n32883) );
  XOR U32509 ( .A(p_input[3885]), .B(p_input[3853]), .Z(n32884) );
  XOR U32510 ( .A(n32885), .B(n32886), .Z(n32876) );
  AND U32511 ( .A(n32887), .B(n32888), .Z(n32886) );
  XOR U32512 ( .A(n32885), .B(n32046), .Z(n32888) );
  XNOR U32513 ( .A(p_input[3916]), .B(n32889), .Z(n32046) );
  AND U32514 ( .A(n695), .B(n32890), .Z(n32889) );
  XOR U32515 ( .A(p_input[3948]), .B(p_input[3916]), .Z(n32890) );
  XNOR U32516 ( .A(n32043), .B(n32885), .Z(n32887) );
  XOR U32517 ( .A(n32891), .B(n32892), .Z(n32043) );
  AND U32518 ( .A(n692), .B(n32893), .Z(n32892) );
  XOR U32519 ( .A(p_input[3884]), .B(p_input[3852]), .Z(n32893) );
  XOR U32520 ( .A(n32894), .B(n32895), .Z(n32885) );
  AND U32521 ( .A(n32896), .B(n32897), .Z(n32895) );
  XOR U32522 ( .A(n32894), .B(n32058), .Z(n32897) );
  XNOR U32523 ( .A(p_input[3915]), .B(n32898), .Z(n32058) );
  AND U32524 ( .A(n695), .B(n32899), .Z(n32898) );
  XOR U32525 ( .A(p_input[3947]), .B(p_input[3915]), .Z(n32899) );
  XNOR U32526 ( .A(n32055), .B(n32894), .Z(n32896) );
  XOR U32527 ( .A(n32900), .B(n32901), .Z(n32055) );
  AND U32528 ( .A(n692), .B(n32902), .Z(n32901) );
  XOR U32529 ( .A(p_input[3883]), .B(p_input[3851]), .Z(n32902) );
  XOR U32530 ( .A(n32903), .B(n32904), .Z(n32894) );
  AND U32531 ( .A(n32905), .B(n32906), .Z(n32904) );
  XOR U32532 ( .A(n32903), .B(n32070), .Z(n32906) );
  XNOR U32533 ( .A(p_input[3914]), .B(n32907), .Z(n32070) );
  AND U32534 ( .A(n695), .B(n32908), .Z(n32907) );
  XOR U32535 ( .A(p_input[3946]), .B(p_input[3914]), .Z(n32908) );
  XNOR U32536 ( .A(n32067), .B(n32903), .Z(n32905) );
  XOR U32537 ( .A(n32909), .B(n32910), .Z(n32067) );
  AND U32538 ( .A(n692), .B(n32911), .Z(n32910) );
  XOR U32539 ( .A(p_input[3882]), .B(p_input[3850]), .Z(n32911) );
  XOR U32540 ( .A(n32912), .B(n32913), .Z(n32903) );
  AND U32541 ( .A(n32914), .B(n32915), .Z(n32913) );
  XOR U32542 ( .A(n32912), .B(n32082), .Z(n32915) );
  XNOR U32543 ( .A(p_input[3913]), .B(n32916), .Z(n32082) );
  AND U32544 ( .A(n695), .B(n32917), .Z(n32916) );
  XOR U32545 ( .A(p_input[3945]), .B(p_input[3913]), .Z(n32917) );
  XNOR U32546 ( .A(n32079), .B(n32912), .Z(n32914) );
  XOR U32547 ( .A(n32918), .B(n32919), .Z(n32079) );
  AND U32548 ( .A(n692), .B(n32920), .Z(n32919) );
  XOR U32549 ( .A(p_input[3881]), .B(p_input[3849]), .Z(n32920) );
  XOR U32550 ( .A(n32921), .B(n32922), .Z(n32912) );
  AND U32551 ( .A(n32923), .B(n32924), .Z(n32922) );
  XOR U32552 ( .A(n32921), .B(n32094), .Z(n32924) );
  XNOR U32553 ( .A(p_input[3912]), .B(n32925), .Z(n32094) );
  AND U32554 ( .A(n695), .B(n32926), .Z(n32925) );
  XOR U32555 ( .A(p_input[3944]), .B(p_input[3912]), .Z(n32926) );
  XNOR U32556 ( .A(n32091), .B(n32921), .Z(n32923) );
  XOR U32557 ( .A(n32927), .B(n32928), .Z(n32091) );
  AND U32558 ( .A(n692), .B(n32929), .Z(n32928) );
  XOR U32559 ( .A(p_input[3880]), .B(p_input[3848]), .Z(n32929) );
  XOR U32560 ( .A(n32930), .B(n32931), .Z(n32921) );
  AND U32561 ( .A(n32932), .B(n32933), .Z(n32931) );
  XOR U32562 ( .A(n32930), .B(n32106), .Z(n32933) );
  XNOR U32563 ( .A(p_input[3911]), .B(n32934), .Z(n32106) );
  AND U32564 ( .A(n695), .B(n32935), .Z(n32934) );
  XOR U32565 ( .A(p_input[3943]), .B(p_input[3911]), .Z(n32935) );
  XNOR U32566 ( .A(n32103), .B(n32930), .Z(n32932) );
  XOR U32567 ( .A(n32936), .B(n32937), .Z(n32103) );
  AND U32568 ( .A(n692), .B(n32938), .Z(n32937) );
  XOR U32569 ( .A(p_input[3879]), .B(p_input[3847]), .Z(n32938) );
  XOR U32570 ( .A(n32939), .B(n32940), .Z(n32930) );
  AND U32571 ( .A(n32941), .B(n32942), .Z(n32940) );
  XOR U32572 ( .A(n32939), .B(n32118), .Z(n32942) );
  XNOR U32573 ( .A(p_input[3910]), .B(n32943), .Z(n32118) );
  AND U32574 ( .A(n695), .B(n32944), .Z(n32943) );
  XOR U32575 ( .A(p_input[3942]), .B(p_input[3910]), .Z(n32944) );
  XNOR U32576 ( .A(n32115), .B(n32939), .Z(n32941) );
  XOR U32577 ( .A(n32945), .B(n32946), .Z(n32115) );
  AND U32578 ( .A(n692), .B(n32947), .Z(n32946) );
  XOR U32579 ( .A(p_input[3878]), .B(p_input[3846]), .Z(n32947) );
  XOR U32580 ( .A(n32948), .B(n32949), .Z(n32939) );
  AND U32581 ( .A(n32950), .B(n32951), .Z(n32949) );
  XOR U32582 ( .A(n32948), .B(n32130), .Z(n32951) );
  XNOR U32583 ( .A(p_input[3909]), .B(n32952), .Z(n32130) );
  AND U32584 ( .A(n695), .B(n32953), .Z(n32952) );
  XOR U32585 ( .A(p_input[3941]), .B(p_input[3909]), .Z(n32953) );
  XNOR U32586 ( .A(n32127), .B(n32948), .Z(n32950) );
  XOR U32587 ( .A(n32954), .B(n32955), .Z(n32127) );
  AND U32588 ( .A(n692), .B(n32956), .Z(n32955) );
  XOR U32589 ( .A(p_input[3877]), .B(p_input[3845]), .Z(n32956) );
  XOR U32590 ( .A(n32957), .B(n32958), .Z(n32948) );
  AND U32591 ( .A(n32959), .B(n32960), .Z(n32958) );
  XOR U32592 ( .A(n32957), .B(n32142), .Z(n32960) );
  XNOR U32593 ( .A(p_input[3908]), .B(n32961), .Z(n32142) );
  AND U32594 ( .A(n695), .B(n32962), .Z(n32961) );
  XOR U32595 ( .A(p_input[3940]), .B(p_input[3908]), .Z(n32962) );
  XNOR U32596 ( .A(n32139), .B(n32957), .Z(n32959) );
  XOR U32597 ( .A(n32963), .B(n32964), .Z(n32139) );
  AND U32598 ( .A(n692), .B(n32965), .Z(n32964) );
  XOR U32599 ( .A(p_input[3876]), .B(p_input[3844]), .Z(n32965) );
  XOR U32600 ( .A(n32966), .B(n32967), .Z(n32957) );
  AND U32601 ( .A(n32968), .B(n32969), .Z(n32967) );
  XOR U32602 ( .A(n32966), .B(n32154), .Z(n32969) );
  XNOR U32603 ( .A(p_input[3907]), .B(n32970), .Z(n32154) );
  AND U32604 ( .A(n695), .B(n32971), .Z(n32970) );
  XOR U32605 ( .A(p_input[3939]), .B(p_input[3907]), .Z(n32971) );
  XNOR U32606 ( .A(n32151), .B(n32966), .Z(n32968) );
  XOR U32607 ( .A(n32972), .B(n32973), .Z(n32151) );
  AND U32608 ( .A(n692), .B(n32974), .Z(n32973) );
  XOR U32609 ( .A(p_input[3875]), .B(p_input[3843]), .Z(n32974) );
  XOR U32610 ( .A(n32975), .B(n32976), .Z(n32966) );
  AND U32611 ( .A(n32977), .B(n32978), .Z(n32976) );
  XOR U32612 ( .A(n32975), .B(n32166), .Z(n32978) );
  XNOR U32613 ( .A(p_input[3906]), .B(n32979), .Z(n32166) );
  AND U32614 ( .A(n695), .B(n32980), .Z(n32979) );
  XOR U32615 ( .A(p_input[3938]), .B(p_input[3906]), .Z(n32980) );
  XNOR U32616 ( .A(n32163), .B(n32975), .Z(n32977) );
  XOR U32617 ( .A(n32981), .B(n32982), .Z(n32163) );
  AND U32618 ( .A(n692), .B(n32983), .Z(n32982) );
  XOR U32619 ( .A(p_input[3874]), .B(p_input[3842]), .Z(n32983) );
  XOR U32620 ( .A(n32984), .B(n32985), .Z(n32975) );
  AND U32621 ( .A(n32986), .B(n32987), .Z(n32985) );
  XNOR U32622 ( .A(n32988), .B(n32179), .Z(n32987) );
  XNOR U32623 ( .A(p_input[3905]), .B(n32989), .Z(n32179) );
  AND U32624 ( .A(n695), .B(n32990), .Z(n32989) );
  XNOR U32625 ( .A(p_input[3937]), .B(n32991), .Z(n32990) );
  IV U32626 ( .A(p_input[3905]), .Z(n32991) );
  XNOR U32627 ( .A(n32176), .B(n32984), .Z(n32986) );
  XNOR U32628 ( .A(p_input[3841]), .B(n32992), .Z(n32176) );
  AND U32629 ( .A(n692), .B(n32993), .Z(n32992) );
  XOR U32630 ( .A(p_input[3873]), .B(p_input[3841]), .Z(n32993) );
  IV U32631 ( .A(n32988), .Z(n32984) );
  AND U32632 ( .A(n32714), .B(n32717), .Z(n32988) );
  XOR U32633 ( .A(p_input[3904]), .B(n32994), .Z(n32717) );
  AND U32634 ( .A(n695), .B(n32995), .Z(n32994) );
  XOR U32635 ( .A(p_input[3936]), .B(p_input[3904]), .Z(n32995) );
  XOR U32636 ( .A(n32996), .B(n32997), .Z(n695) );
  AND U32637 ( .A(n32998), .B(n32999), .Z(n32997) );
  XNOR U32638 ( .A(p_input[3967]), .B(n32996), .Z(n32999) );
  XOR U32639 ( .A(n32996), .B(p_input[3935]), .Z(n32998) );
  XOR U32640 ( .A(n33000), .B(n33001), .Z(n32996) );
  AND U32641 ( .A(n33002), .B(n33003), .Z(n33001) );
  XNOR U32642 ( .A(p_input[3966]), .B(n33000), .Z(n33003) );
  XOR U32643 ( .A(n33000), .B(p_input[3934]), .Z(n33002) );
  XOR U32644 ( .A(n33004), .B(n33005), .Z(n33000) );
  AND U32645 ( .A(n33006), .B(n33007), .Z(n33005) );
  XNOR U32646 ( .A(p_input[3965]), .B(n33004), .Z(n33007) );
  XOR U32647 ( .A(n33004), .B(p_input[3933]), .Z(n33006) );
  XOR U32648 ( .A(n33008), .B(n33009), .Z(n33004) );
  AND U32649 ( .A(n33010), .B(n33011), .Z(n33009) );
  XNOR U32650 ( .A(p_input[3964]), .B(n33008), .Z(n33011) );
  XOR U32651 ( .A(n33008), .B(p_input[3932]), .Z(n33010) );
  XOR U32652 ( .A(n33012), .B(n33013), .Z(n33008) );
  AND U32653 ( .A(n33014), .B(n33015), .Z(n33013) );
  XNOR U32654 ( .A(p_input[3963]), .B(n33012), .Z(n33015) );
  XOR U32655 ( .A(n33012), .B(p_input[3931]), .Z(n33014) );
  XOR U32656 ( .A(n33016), .B(n33017), .Z(n33012) );
  AND U32657 ( .A(n33018), .B(n33019), .Z(n33017) );
  XNOR U32658 ( .A(p_input[3962]), .B(n33016), .Z(n33019) );
  XOR U32659 ( .A(n33016), .B(p_input[3930]), .Z(n33018) );
  XOR U32660 ( .A(n33020), .B(n33021), .Z(n33016) );
  AND U32661 ( .A(n33022), .B(n33023), .Z(n33021) );
  XNOR U32662 ( .A(p_input[3961]), .B(n33020), .Z(n33023) );
  XOR U32663 ( .A(n33020), .B(p_input[3929]), .Z(n33022) );
  XOR U32664 ( .A(n33024), .B(n33025), .Z(n33020) );
  AND U32665 ( .A(n33026), .B(n33027), .Z(n33025) );
  XNOR U32666 ( .A(p_input[3960]), .B(n33024), .Z(n33027) );
  XOR U32667 ( .A(n33024), .B(p_input[3928]), .Z(n33026) );
  XOR U32668 ( .A(n33028), .B(n33029), .Z(n33024) );
  AND U32669 ( .A(n33030), .B(n33031), .Z(n33029) );
  XNOR U32670 ( .A(p_input[3959]), .B(n33028), .Z(n33031) );
  XOR U32671 ( .A(n33028), .B(p_input[3927]), .Z(n33030) );
  XOR U32672 ( .A(n33032), .B(n33033), .Z(n33028) );
  AND U32673 ( .A(n33034), .B(n33035), .Z(n33033) );
  XNOR U32674 ( .A(p_input[3958]), .B(n33032), .Z(n33035) );
  XOR U32675 ( .A(n33032), .B(p_input[3926]), .Z(n33034) );
  XOR U32676 ( .A(n33036), .B(n33037), .Z(n33032) );
  AND U32677 ( .A(n33038), .B(n33039), .Z(n33037) );
  XNOR U32678 ( .A(p_input[3957]), .B(n33036), .Z(n33039) );
  XOR U32679 ( .A(n33036), .B(p_input[3925]), .Z(n33038) );
  XOR U32680 ( .A(n33040), .B(n33041), .Z(n33036) );
  AND U32681 ( .A(n33042), .B(n33043), .Z(n33041) );
  XNOR U32682 ( .A(p_input[3956]), .B(n33040), .Z(n33043) );
  XOR U32683 ( .A(n33040), .B(p_input[3924]), .Z(n33042) );
  XOR U32684 ( .A(n33044), .B(n33045), .Z(n33040) );
  AND U32685 ( .A(n33046), .B(n33047), .Z(n33045) );
  XNOR U32686 ( .A(p_input[3955]), .B(n33044), .Z(n33047) );
  XOR U32687 ( .A(n33044), .B(p_input[3923]), .Z(n33046) );
  XOR U32688 ( .A(n33048), .B(n33049), .Z(n33044) );
  AND U32689 ( .A(n33050), .B(n33051), .Z(n33049) );
  XNOR U32690 ( .A(p_input[3954]), .B(n33048), .Z(n33051) );
  XOR U32691 ( .A(n33048), .B(p_input[3922]), .Z(n33050) );
  XOR U32692 ( .A(n33052), .B(n33053), .Z(n33048) );
  AND U32693 ( .A(n33054), .B(n33055), .Z(n33053) );
  XNOR U32694 ( .A(p_input[3953]), .B(n33052), .Z(n33055) );
  XOR U32695 ( .A(n33052), .B(p_input[3921]), .Z(n33054) );
  XOR U32696 ( .A(n33056), .B(n33057), .Z(n33052) );
  AND U32697 ( .A(n33058), .B(n33059), .Z(n33057) );
  XNOR U32698 ( .A(p_input[3952]), .B(n33056), .Z(n33059) );
  XOR U32699 ( .A(n33056), .B(p_input[3920]), .Z(n33058) );
  XOR U32700 ( .A(n33060), .B(n33061), .Z(n33056) );
  AND U32701 ( .A(n33062), .B(n33063), .Z(n33061) );
  XNOR U32702 ( .A(p_input[3951]), .B(n33060), .Z(n33063) );
  XOR U32703 ( .A(n33060), .B(p_input[3919]), .Z(n33062) );
  XOR U32704 ( .A(n33064), .B(n33065), .Z(n33060) );
  AND U32705 ( .A(n33066), .B(n33067), .Z(n33065) );
  XNOR U32706 ( .A(p_input[3950]), .B(n33064), .Z(n33067) );
  XOR U32707 ( .A(n33064), .B(p_input[3918]), .Z(n33066) );
  XOR U32708 ( .A(n33068), .B(n33069), .Z(n33064) );
  AND U32709 ( .A(n33070), .B(n33071), .Z(n33069) );
  XNOR U32710 ( .A(p_input[3949]), .B(n33068), .Z(n33071) );
  XOR U32711 ( .A(n33068), .B(p_input[3917]), .Z(n33070) );
  XOR U32712 ( .A(n33072), .B(n33073), .Z(n33068) );
  AND U32713 ( .A(n33074), .B(n33075), .Z(n33073) );
  XNOR U32714 ( .A(p_input[3948]), .B(n33072), .Z(n33075) );
  XOR U32715 ( .A(n33072), .B(p_input[3916]), .Z(n33074) );
  XOR U32716 ( .A(n33076), .B(n33077), .Z(n33072) );
  AND U32717 ( .A(n33078), .B(n33079), .Z(n33077) );
  XNOR U32718 ( .A(p_input[3947]), .B(n33076), .Z(n33079) );
  XOR U32719 ( .A(n33076), .B(p_input[3915]), .Z(n33078) );
  XOR U32720 ( .A(n33080), .B(n33081), .Z(n33076) );
  AND U32721 ( .A(n33082), .B(n33083), .Z(n33081) );
  XNOR U32722 ( .A(p_input[3946]), .B(n33080), .Z(n33083) );
  XOR U32723 ( .A(n33080), .B(p_input[3914]), .Z(n33082) );
  XOR U32724 ( .A(n33084), .B(n33085), .Z(n33080) );
  AND U32725 ( .A(n33086), .B(n33087), .Z(n33085) );
  XNOR U32726 ( .A(p_input[3945]), .B(n33084), .Z(n33087) );
  XOR U32727 ( .A(n33084), .B(p_input[3913]), .Z(n33086) );
  XOR U32728 ( .A(n33088), .B(n33089), .Z(n33084) );
  AND U32729 ( .A(n33090), .B(n33091), .Z(n33089) );
  XNOR U32730 ( .A(p_input[3944]), .B(n33088), .Z(n33091) );
  XOR U32731 ( .A(n33088), .B(p_input[3912]), .Z(n33090) );
  XOR U32732 ( .A(n33092), .B(n33093), .Z(n33088) );
  AND U32733 ( .A(n33094), .B(n33095), .Z(n33093) );
  XNOR U32734 ( .A(p_input[3943]), .B(n33092), .Z(n33095) );
  XOR U32735 ( .A(n33092), .B(p_input[3911]), .Z(n33094) );
  XOR U32736 ( .A(n33096), .B(n33097), .Z(n33092) );
  AND U32737 ( .A(n33098), .B(n33099), .Z(n33097) );
  XNOR U32738 ( .A(p_input[3942]), .B(n33096), .Z(n33099) );
  XOR U32739 ( .A(n33096), .B(p_input[3910]), .Z(n33098) );
  XOR U32740 ( .A(n33100), .B(n33101), .Z(n33096) );
  AND U32741 ( .A(n33102), .B(n33103), .Z(n33101) );
  XNOR U32742 ( .A(p_input[3941]), .B(n33100), .Z(n33103) );
  XOR U32743 ( .A(n33100), .B(p_input[3909]), .Z(n33102) );
  XOR U32744 ( .A(n33104), .B(n33105), .Z(n33100) );
  AND U32745 ( .A(n33106), .B(n33107), .Z(n33105) );
  XNOR U32746 ( .A(p_input[3940]), .B(n33104), .Z(n33107) );
  XOR U32747 ( .A(n33104), .B(p_input[3908]), .Z(n33106) );
  XOR U32748 ( .A(n33108), .B(n33109), .Z(n33104) );
  AND U32749 ( .A(n33110), .B(n33111), .Z(n33109) );
  XNOR U32750 ( .A(p_input[3939]), .B(n33108), .Z(n33111) );
  XOR U32751 ( .A(n33108), .B(p_input[3907]), .Z(n33110) );
  XOR U32752 ( .A(n33112), .B(n33113), .Z(n33108) );
  AND U32753 ( .A(n33114), .B(n33115), .Z(n33113) );
  XNOR U32754 ( .A(p_input[3938]), .B(n33112), .Z(n33115) );
  XOR U32755 ( .A(n33112), .B(p_input[3906]), .Z(n33114) );
  XNOR U32756 ( .A(n33116), .B(n33117), .Z(n33112) );
  AND U32757 ( .A(n33118), .B(n33119), .Z(n33117) );
  XOR U32758 ( .A(p_input[3937]), .B(n33116), .Z(n33119) );
  XNOR U32759 ( .A(p_input[3905]), .B(n33116), .Z(n33118) );
  AND U32760 ( .A(p_input[3936]), .B(n33120), .Z(n33116) );
  IV U32761 ( .A(p_input[3904]), .Z(n33120) );
  XNOR U32762 ( .A(p_input[3840]), .B(n33121), .Z(n32714) );
  AND U32763 ( .A(n692), .B(n33122), .Z(n33121) );
  XOR U32764 ( .A(p_input[3872]), .B(p_input[3840]), .Z(n33122) );
  XOR U32765 ( .A(n33123), .B(n33124), .Z(n692) );
  AND U32766 ( .A(n33125), .B(n33126), .Z(n33124) );
  XNOR U32767 ( .A(p_input[3903]), .B(n33123), .Z(n33126) );
  XOR U32768 ( .A(n33123), .B(p_input[3871]), .Z(n33125) );
  XOR U32769 ( .A(n33127), .B(n33128), .Z(n33123) );
  AND U32770 ( .A(n33129), .B(n33130), .Z(n33128) );
  XNOR U32771 ( .A(p_input[3902]), .B(n33127), .Z(n33130) );
  XNOR U32772 ( .A(n33127), .B(n32729), .Z(n33129) );
  IV U32773 ( .A(p_input[3870]), .Z(n32729) );
  XOR U32774 ( .A(n33131), .B(n33132), .Z(n33127) );
  AND U32775 ( .A(n33133), .B(n33134), .Z(n33132) );
  XNOR U32776 ( .A(p_input[3901]), .B(n33131), .Z(n33134) );
  XNOR U32777 ( .A(n33131), .B(n32738), .Z(n33133) );
  IV U32778 ( .A(p_input[3869]), .Z(n32738) );
  XOR U32779 ( .A(n33135), .B(n33136), .Z(n33131) );
  AND U32780 ( .A(n33137), .B(n33138), .Z(n33136) );
  XNOR U32781 ( .A(p_input[3900]), .B(n33135), .Z(n33138) );
  XNOR U32782 ( .A(n33135), .B(n32747), .Z(n33137) );
  IV U32783 ( .A(p_input[3868]), .Z(n32747) );
  XOR U32784 ( .A(n33139), .B(n33140), .Z(n33135) );
  AND U32785 ( .A(n33141), .B(n33142), .Z(n33140) );
  XNOR U32786 ( .A(p_input[3899]), .B(n33139), .Z(n33142) );
  XNOR U32787 ( .A(n33139), .B(n32756), .Z(n33141) );
  IV U32788 ( .A(p_input[3867]), .Z(n32756) );
  XOR U32789 ( .A(n33143), .B(n33144), .Z(n33139) );
  AND U32790 ( .A(n33145), .B(n33146), .Z(n33144) );
  XNOR U32791 ( .A(p_input[3898]), .B(n33143), .Z(n33146) );
  XNOR U32792 ( .A(n33143), .B(n32765), .Z(n33145) );
  IV U32793 ( .A(p_input[3866]), .Z(n32765) );
  XOR U32794 ( .A(n33147), .B(n33148), .Z(n33143) );
  AND U32795 ( .A(n33149), .B(n33150), .Z(n33148) );
  XNOR U32796 ( .A(p_input[3897]), .B(n33147), .Z(n33150) );
  XNOR U32797 ( .A(n33147), .B(n32774), .Z(n33149) );
  IV U32798 ( .A(p_input[3865]), .Z(n32774) );
  XOR U32799 ( .A(n33151), .B(n33152), .Z(n33147) );
  AND U32800 ( .A(n33153), .B(n33154), .Z(n33152) );
  XNOR U32801 ( .A(p_input[3896]), .B(n33151), .Z(n33154) );
  XNOR U32802 ( .A(n33151), .B(n32783), .Z(n33153) );
  IV U32803 ( .A(p_input[3864]), .Z(n32783) );
  XOR U32804 ( .A(n33155), .B(n33156), .Z(n33151) );
  AND U32805 ( .A(n33157), .B(n33158), .Z(n33156) );
  XNOR U32806 ( .A(p_input[3895]), .B(n33155), .Z(n33158) );
  XNOR U32807 ( .A(n33155), .B(n32792), .Z(n33157) );
  IV U32808 ( .A(p_input[3863]), .Z(n32792) );
  XOR U32809 ( .A(n33159), .B(n33160), .Z(n33155) );
  AND U32810 ( .A(n33161), .B(n33162), .Z(n33160) );
  XNOR U32811 ( .A(p_input[3894]), .B(n33159), .Z(n33162) );
  XNOR U32812 ( .A(n33159), .B(n32801), .Z(n33161) );
  IV U32813 ( .A(p_input[3862]), .Z(n32801) );
  XOR U32814 ( .A(n33163), .B(n33164), .Z(n33159) );
  AND U32815 ( .A(n33165), .B(n33166), .Z(n33164) );
  XNOR U32816 ( .A(p_input[3893]), .B(n33163), .Z(n33166) );
  XNOR U32817 ( .A(n33163), .B(n32810), .Z(n33165) );
  IV U32818 ( .A(p_input[3861]), .Z(n32810) );
  XOR U32819 ( .A(n33167), .B(n33168), .Z(n33163) );
  AND U32820 ( .A(n33169), .B(n33170), .Z(n33168) );
  XNOR U32821 ( .A(p_input[3892]), .B(n33167), .Z(n33170) );
  XNOR U32822 ( .A(n33167), .B(n32819), .Z(n33169) );
  IV U32823 ( .A(p_input[3860]), .Z(n32819) );
  XOR U32824 ( .A(n33171), .B(n33172), .Z(n33167) );
  AND U32825 ( .A(n33173), .B(n33174), .Z(n33172) );
  XNOR U32826 ( .A(p_input[3891]), .B(n33171), .Z(n33174) );
  XNOR U32827 ( .A(n33171), .B(n32828), .Z(n33173) );
  IV U32828 ( .A(p_input[3859]), .Z(n32828) );
  XOR U32829 ( .A(n33175), .B(n33176), .Z(n33171) );
  AND U32830 ( .A(n33177), .B(n33178), .Z(n33176) );
  XNOR U32831 ( .A(p_input[3890]), .B(n33175), .Z(n33178) );
  XNOR U32832 ( .A(n33175), .B(n32837), .Z(n33177) );
  IV U32833 ( .A(p_input[3858]), .Z(n32837) );
  XOR U32834 ( .A(n33179), .B(n33180), .Z(n33175) );
  AND U32835 ( .A(n33181), .B(n33182), .Z(n33180) );
  XNOR U32836 ( .A(p_input[3889]), .B(n33179), .Z(n33182) );
  XNOR U32837 ( .A(n33179), .B(n32846), .Z(n33181) );
  IV U32838 ( .A(p_input[3857]), .Z(n32846) );
  XOR U32839 ( .A(n33183), .B(n33184), .Z(n33179) );
  AND U32840 ( .A(n33185), .B(n33186), .Z(n33184) );
  XNOR U32841 ( .A(p_input[3888]), .B(n33183), .Z(n33186) );
  XNOR U32842 ( .A(n33183), .B(n32855), .Z(n33185) );
  IV U32843 ( .A(p_input[3856]), .Z(n32855) );
  XOR U32844 ( .A(n33187), .B(n33188), .Z(n33183) );
  AND U32845 ( .A(n33189), .B(n33190), .Z(n33188) );
  XNOR U32846 ( .A(p_input[3887]), .B(n33187), .Z(n33190) );
  XNOR U32847 ( .A(n33187), .B(n32864), .Z(n33189) );
  IV U32848 ( .A(p_input[3855]), .Z(n32864) );
  XOR U32849 ( .A(n33191), .B(n33192), .Z(n33187) );
  AND U32850 ( .A(n33193), .B(n33194), .Z(n33192) );
  XNOR U32851 ( .A(p_input[3886]), .B(n33191), .Z(n33194) );
  XNOR U32852 ( .A(n33191), .B(n32873), .Z(n33193) );
  IV U32853 ( .A(p_input[3854]), .Z(n32873) );
  XOR U32854 ( .A(n33195), .B(n33196), .Z(n33191) );
  AND U32855 ( .A(n33197), .B(n33198), .Z(n33196) );
  XNOR U32856 ( .A(p_input[3885]), .B(n33195), .Z(n33198) );
  XNOR U32857 ( .A(n33195), .B(n32882), .Z(n33197) );
  IV U32858 ( .A(p_input[3853]), .Z(n32882) );
  XOR U32859 ( .A(n33199), .B(n33200), .Z(n33195) );
  AND U32860 ( .A(n33201), .B(n33202), .Z(n33200) );
  XNOR U32861 ( .A(p_input[3884]), .B(n33199), .Z(n33202) );
  XNOR U32862 ( .A(n33199), .B(n32891), .Z(n33201) );
  IV U32863 ( .A(p_input[3852]), .Z(n32891) );
  XOR U32864 ( .A(n33203), .B(n33204), .Z(n33199) );
  AND U32865 ( .A(n33205), .B(n33206), .Z(n33204) );
  XNOR U32866 ( .A(p_input[3883]), .B(n33203), .Z(n33206) );
  XNOR U32867 ( .A(n33203), .B(n32900), .Z(n33205) );
  IV U32868 ( .A(p_input[3851]), .Z(n32900) );
  XOR U32869 ( .A(n33207), .B(n33208), .Z(n33203) );
  AND U32870 ( .A(n33209), .B(n33210), .Z(n33208) );
  XNOR U32871 ( .A(p_input[3882]), .B(n33207), .Z(n33210) );
  XNOR U32872 ( .A(n33207), .B(n32909), .Z(n33209) );
  IV U32873 ( .A(p_input[3850]), .Z(n32909) );
  XOR U32874 ( .A(n33211), .B(n33212), .Z(n33207) );
  AND U32875 ( .A(n33213), .B(n33214), .Z(n33212) );
  XNOR U32876 ( .A(p_input[3881]), .B(n33211), .Z(n33214) );
  XNOR U32877 ( .A(n33211), .B(n32918), .Z(n33213) );
  IV U32878 ( .A(p_input[3849]), .Z(n32918) );
  XOR U32879 ( .A(n33215), .B(n33216), .Z(n33211) );
  AND U32880 ( .A(n33217), .B(n33218), .Z(n33216) );
  XNOR U32881 ( .A(p_input[3880]), .B(n33215), .Z(n33218) );
  XNOR U32882 ( .A(n33215), .B(n32927), .Z(n33217) );
  IV U32883 ( .A(p_input[3848]), .Z(n32927) );
  XOR U32884 ( .A(n33219), .B(n33220), .Z(n33215) );
  AND U32885 ( .A(n33221), .B(n33222), .Z(n33220) );
  XNOR U32886 ( .A(p_input[3879]), .B(n33219), .Z(n33222) );
  XNOR U32887 ( .A(n33219), .B(n32936), .Z(n33221) );
  IV U32888 ( .A(p_input[3847]), .Z(n32936) );
  XOR U32889 ( .A(n33223), .B(n33224), .Z(n33219) );
  AND U32890 ( .A(n33225), .B(n33226), .Z(n33224) );
  XNOR U32891 ( .A(p_input[3878]), .B(n33223), .Z(n33226) );
  XNOR U32892 ( .A(n33223), .B(n32945), .Z(n33225) );
  IV U32893 ( .A(p_input[3846]), .Z(n32945) );
  XOR U32894 ( .A(n33227), .B(n33228), .Z(n33223) );
  AND U32895 ( .A(n33229), .B(n33230), .Z(n33228) );
  XNOR U32896 ( .A(p_input[3877]), .B(n33227), .Z(n33230) );
  XNOR U32897 ( .A(n33227), .B(n32954), .Z(n33229) );
  IV U32898 ( .A(p_input[3845]), .Z(n32954) );
  XOR U32899 ( .A(n33231), .B(n33232), .Z(n33227) );
  AND U32900 ( .A(n33233), .B(n33234), .Z(n33232) );
  XNOR U32901 ( .A(p_input[3876]), .B(n33231), .Z(n33234) );
  XNOR U32902 ( .A(n33231), .B(n32963), .Z(n33233) );
  IV U32903 ( .A(p_input[3844]), .Z(n32963) );
  XOR U32904 ( .A(n33235), .B(n33236), .Z(n33231) );
  AND U32905 ( .A(n33237), .B(n33238), .Z(n33236) );
  XNOR U32906 ( .A(p_input[3875]), .B(n33235), .Z(n33238) );
  XNOR U32907 ( .A(n33235), .B(n32972), .Z(n33237) );
  IV U32908 ( .A(p_input[3843]), .Z(n32972) );
  XOR U32909 ( .A(n33239), .B(n33240), .Z(n33235) );
  AND U32910 ( .A(n33241), .B(n33242), .Z(n33240) );
  XNOR U32911 ( .A(p_input[3874]), .B(n33239), .Z(n33242) );
  XNOR U32912 ( .A(n33239), .B(n32981), .Z(n33241) );
  IV U32913 ( .A(p_input[3842]), .Z(n32981) );
  XNOR U32914 ( .A(n33243), .B(n33244), .Z(n33239) );
  AND U32915 ( .A(n33245), .B(n33246), .Z(n33244) );
  XOR U32916 ( .A(p_input[3873]), .B(n33243), .Z(n33246) );
  XNOR U32917 ( .A(p_input[3841]), .B(n33243), .Z(n33245) );
  AND U32918 ( .A(p_input[3872]), .B(n33247), .Z(n33243) );
  IV U32919 ( .A(p_input[3840]), .Z(n33247) );
  XOR U32920 ( .A(n33248), .B(n33249), .Z(n31426) );
  AND U32921 ( .A(n873), .B(n33250), .Z(n33249) );
  XNOR U32922 ( .A(n33251), .B(n33248), .Z(n33250) );
  XOR U32923 ( .A(n33252), .B(n33253), .Z(n873) );
  AND U32924 ( .A(n33254), .B(n33255), .Z(n33253) );
  XOR U32925 ( .A(n33252), .B(n31441), .Z(n33255) );
  XNOR U32926 ( .A(n33256), .B(n33257), .Z(n31441) );
  AND U32927 ( .A(n33258), .B(n567), .Z(n33257) );
  AND U32928 ( .A(n33256), .B(n33259), .Z(n33258) );
  XNOR U32929 ( .A(n31438), .B(n33252), .Z(n33254) );
  XOR U32930 ( .A(n33260), .B(n33261), .Z(n31438) );
  AND U32931 ( .A(n33262), .B(n564), .Z(n33261) );
  NOR U32932 ( .A(n33260), .B(n33263), .Z(n33262) );
  XOR U32933 ( .A(n33264), .B(n33265), .Z(n33252) );
  AND U32934 ( .A(n33266), .B(n33267), .Z(n33265) );
  XOR U32935 ( .A(n33264), .B(n31453), .Z(n33267) );
  XOR U32936 ( .A(n33268), .B(n33269), .Z(n31453) );
  AND U32937 ( .A(n567), .B(n33270), .Z(n33269) );
  XOR U32938 ( .A(n33271), .B(n33268), .Z(n33270) );
  XNOR U32939 ( .A(n31450), .B(n33264), .Z(n33266) );
  XOR U32940 ( .A(n33272), .B(n33273), .Z(n31450) );
  AND U32941 ( .A(n564), .B(n33274), .Z(n33273) );
  XOR U32942 ( .A(n33275), .B(n33272), .Z(n33274) );
  XOR U32943 ( .A(n33276), .B(n33277), .Z(n33264) );
  AND U32944 ( .A(n33278), .B(n33279), .Z(n33277) );
  XOR U32945 ( .A(n33276), .B(n31465), .Z(n33279) );
  XOR U32946 ( .A(n33280), .B(n33281), .Z(n31465) );
  AND U32947 ( .A(n567), .B(n33282), .Z(n33281) );
  XOR U32948 ( .A(n33283), .B(n33280), .Z(n33282) );
  XNOR U32949 ( .A(n31462), .B(n33276), .Z(n33278) );
  XOR U32950 ( .A(n33284), .B(n33285), .Z(n31462) );
  AND U32951 ( .A(n564), .B(n33286), .Z(n33285) );
  XOR U32952 ( .A(n33287), .B(n33284), .Z(n33286) );
  XOR U32953 ( .A(n33288), .B(n33289), .Z(n33276) );
  AND U32954 ( .A(n33290), .B(n33291), .Z(n33289) );
  XOR U32955 ( .A(n33288), .B(n31477), .Z(n33291) );
  XOR U32956 ( .A(n33292), .B(n33293), .Z(n31477) );
  AND U32957 ( .A(n567), .B(n33294), .Z(n33293) );
  XOR U32958 ( .A(n33295), .B(n33292), .Z(n33294) );
  XNOR U32959 ( .A(n31474), .B(n33288), .Z(n33290) );
  XOR U32960 ( .A(n33296), .B(n33297), .Z(n31474) );
  AND U32961 ( .A(n564), .B(n33298), .Z(n33297) );
  XOR U32962 ( .A(n33299), .B(n33296), .Z(n33298) );
  XOR U32963 ( .A(n33300), .B(n33301), .Z(n33288) );
  AND U32964 ( .A(n33302), .B(n33303), .Z(n33301) );
  XOR U32965 ( .A(n33300), .B(n31489), .Z(n33303) );
  XOR U32966 ( .A(n33304), .B(n33305), .Z(n31489) );
  AND U32967 ( .A(n567), .B(n33306), .Z(n33305) );
  XOR U32968 ( .A(n33307), .B(n33304), .Z(n33306) );
  XNOR U32969 ( .A(n31486), .B(n33300), .Z(n33302) );
  XOR U32970 ( .A(n33308), .B(n33309), .Z(n31486) );
  AND U32971 ( .A(n564), .B(n33310), .Z(n33309) );
  XOR U32972 ( .A(n33311), .B(n33308), .Z(n33310) );
  XOR U32973 ( .A(n33312), .B(n33313), .Z(n33300) );
  AND U32974 ( .A(n33314), .B(n33315), .Z(n33313) );
  XOR U32975 ( .A(n33312), .B(n31501), .Z(n33315) );
  XOR U32976 ( .A(n33316), .B(n33317), .Z(n31501) );
  AND U32977 ( .A(n567), .B(n33318), .Z(n33317) );
  XOR U32978 ( .A(n33319), .B(n33316), .Z(n33318) );
  XNOR U32979 ( .A(n31498), .B(n33312), .Z(n33314) );
  XOR U32980 ( .A(n33320), .B(n33321), .Z(n31498) );
  AND U32981 ( .A(n564), .B(n33322), .Z(n33321) );
  XOR U32982 ( .A(n33323), .B(n33320), .Z(n33322) );
  XOR U32983 ( .A(n33324), .B(n33325), .Z(n33312) );
  AND U32984 ( .A(n33326), .B(n33327), .Z(n33325) );
  XOR U32985 ( .A(n33324), .B(n31513), .Z(n33327) );
  XOR U32986 ( .A(n33328), .B(n33329), .Z(n31513) );
  AND U32987 ( .A(n567), .B(n33330), .Z(n33329) );
  XOR U32988 ( .A(n33331), .B(n33328), .Z(n33330) );
  XNOR U32989 ( .A(n31510), .B(n33324), .Z(n33326) );
  XOR U32990 ( .A(n33332), .B(n33333), .Z(n31510) );
  AND U32991 ( .A(n564), .B(n33334), .Z(n33333) );
  XOR U32992 ( .A(n33335), .B(n33332), .Z(n33334) );
  XOR U32993 ( .A(n33336), .B(n33337), .Z(n33324) );
  AND U32994 ( .A(n33338), .B(n33339), .Z(n33337) );
  XOR U32995 ( .A(n33336), .B(n31525), .Z(n33339) );
  XOR U32996 ( .A(n33340), .B(n33341), .Z(n31525) );
  AND U32997 ( .A(n567), .B(n33342), .Z(n33341) );
  XOR U32998 ( .A(n33343), .B(n33340), .Z(n33342) );
  XNOR U32999 ( .A(n31522), .B(n33336), .Z(n33338) );
  XOR U33000 ( .A(n33344), .B(n33345), .Z(n31522) );
  AND U33001 ( .A(n564), .B(n33346), .Z(n33345) );
  XOR U33002 ( .A(n33347), .B(n33344), .Z(n33346) );
  XOR U33003 ( .A(n33348), .B(n33349), .Z(n33336) );
  AND U33004 ( .A(n33350), .B(n33351), .Z(n33349) );
  XOR U33005 ( .A(n33348), .B(n31537), .Z(n33351) );
  XOR U33006 ( .A(n33352), .B(n33353), .Z(n31537) );
  AND U33007 ( .A(n567), .B(n33354), .Z(n33353) );
  XOR U33008 ( .A(n33355), .B(n33352), .Z(n33354) );
  XNOR U33009 ( .A(n31534), .B(n33348), .Z(n33350) );
  XOR U33010 ( .A(n33356), .B(n33357), .Z(n31534) );
  AND U33011 ( .A(n564), .B(n33358), .Z(n33357) );
  XOR U33012 ( .A(n33359), .B(n33356), .Z(n33358) );
  XOR U33013 ( .A(n33360), .B(n33361), .Z(n33348) );
  AND U33014 ( .A(n33362), .B(n33363), .Z(n33361) );
  XOR U33015 ( .A(n33360), .B(n31549), .Z(n33363) );
  XOR U33016 ( .A(n33364), .B(n33365), .Z(n31549) );
  AND U33017 ( .A(n567), .B(n33366), .Z(n33365) );
  XOR U33018 ( .A(n33367), .B(n33364), .Z(n33366) );
  XNOR U33019 ( .A(n31546), .B(n33360), .Z(n33362) );
  XOR U33020 ( .A(n33368), .B(n33369), .Z(n31546) );
  AND U33021 ( .A(n564), .B(n33370), .Z(n33369) );
  XOR U33022 ( .A(n33371), .B(n33368), .Z(n33370) );
  XOR U33023 ( .A(n33372), .B(n33373), .Z(n33360) );
  AND U33024 ( .A(n33374), .B(n33375), .Z(n33373) );
  XOR U33025 ( .A(n33372), .B(n31561), .Z(n33375) );
  XOR U33026 ( .A(n33376), .B(n33377), .Z(n31561) );
  AND U33027 ( .A(n567), .B(n33378), .Z(n33377) );
  XOR U33028 ( .A(n33379), .B(n33376), .Z(n33378) );
  XNOR U33029 ( .A(n31558), .B(n33372), .Z(n33374) );
  XOR U33030 ( .A(n33380), .B(n33381), .Z(n31558) );
  AND U33031 ( .A(n564), .B(n33382), .Z(n33381) );
  XOR U33032 ( .A(n33383), .B(n33380), .Z(n33382) );
  XOR U33033 ( .A(n33384), .B(n33385), .Z(n33372) );
  AND U33034 ( .A(n33386), .B(n33387), .Z(n33385) );
  XOR U33035 ( .A(n33384), .B(n31573), .Z(n33387) );
  XOR U33036 ( .A(n33388), .B(n33389), .Z(n31573) );
  AND U33037 ( .A(n567), .B(n33390), .Z(n33389) );
  XOR U33038 ( .A(n33391), .B(n33388), .Z(n33390) );
  XNOR U33039 ( .A(n31570), .B(n33384), .Z(n33386) );
  XOR U33040 ( .A(n33392), .B(n33393), .Z(n31570) );
  AND U33041 ( .A(n564), .B(n33394), .Z(n33393) );
  XOR U33042 ( .A(n33395), .B(n33392), .Z(n33394) );
  XOR U33043 ( .A(n33396), .B(n33397), .Z(n33384) );
  AND U33044 ( .A(n33398), .B(n33399), .Z(n33397) );
  XOR U33045 ( .A(n33396), .B(n31585), .Z(n33399) );
  XOR U33046 ( .A(n33400), .B(n33401), .Z(n31585) );
  AND U33047 ( .A(n567), .B(n33402), .Z(n33401) );
  XOR U33048 ( .A(n33403), .B(n33400), .Z(n33402) );
  XNOR U33049 ( .A(n31582), .B(n33396), .Z(n33398) );
  XOR U33050 ( .A(n33404), .B(n33405), .Z(n31582) );
  AND U33051 ( .A(n564), .B(n33406), .Z(n33405) );
  XOR U33052 ( .A(n33407), .B(n33404), .Z(n33406) );
  XOR U33053 ( .A(n33408), .B(n33409), .Z(n33396) );
  AND U33054 ( .A(n33410), .B(n33411), .Z(n33409) );
  XOR U33055 ( .A(n33408), .B(n31597), .Z(n33411) );
  XOR U33056 ( .A(n33412), .B(n33413), .Z(n31597) );
  AND U33057 ( .A(n567), .B(n33414), .Z(n33413) );
  XOR U33058 ( .A(n33415), .B(n33412), .Z(n33414) );
  XNOR U33059 ( .A(n31594), .B(n33408), .Z(n33410) );
  XOR U33060 ( .A(n33416), .B(n33417), .Z(n31594) );
  AND U33061 ( .A(n564), .B(n33418), .Z(n33417) );
  XOR U33062 ( .A(n33419), .B(n33416), .Z(n33418) );
  XOR U33063 ( .A(n33420), .B(n33421), .Z(n33408) );
  AND U33064 ( .A(n33422), .B(n33423), .Z(n33421) );
  XOR U33065 ( .A(n33420), .B(n31609), .Z(n33423) );
  XOR U33066 ( .A(n33424), .B(n33425), .Z(n31609) );
  AND U33067 ( .A(n567), .B(n33426), .Z(n33425) );
  XOR U33068 ( .A(n33427), .B(n33424), .Z(n33426) );
  XNOR U33069 ( .A(n31606), .B(n33420), .Z(n33422) );
  XOR U33070 ( .A(n33428), .B(n33429), .Z(n31606) );
  AND U33071 ( .A(n564), .B(n33430), .Z(n33429) );
  XOR U33072 ( .A(n33431), .B(n33428), .Z(n33430) );
  XOR U33073 ( .A(n33432), .B(n33433), .Z(n33420) );
  AND U33074 ( .A(n33434), .B(n33435), .Z(n33433) );
  XOR U33075 ( .A(n33432), .B(n31621), .Z(n33435) );
  XOR U33076 ( .A(n33436), .B(n33437), .Z(n31621) );
  AND U33077 ( .A(n567), .B(n33438), .Z(n33437) );
  XOR U33078 ( .A(n33439), .B(n33436), .Z(n33438) );
  XNOR U33079 ( .A(n31618), .B(n33432), .Z(n33434) );
  XOR U33080 ( .A(n33440), .B(n33441), .Z(n31618) );
  AND U33081 ( .A(n564), .B(n33442), .Z(n33441) );
  XOR U33082 ( .A(n33443), .B(n33440), .Z(n33442) );
  XOR U33083 ( .A(n33444), .B(n33445), .Z(n33432) );
  AND U33084 ( .A(n33446), .B(n33447), .Z(n33445) );
  XOR U33085 ( .A(n33444), .B(n31633), .Z(n33447) );
  XOR U33086 ( .A(n33448), .B(n33449), .Z(n31633) );
  AND U33087 ( .A(n567), .B(n33450), .Z(n33449) );
  XOR U33088 ( .A(n33451), .B(n33448), .Z(n33450) );
  XNOR U33089 ( .A(n31630), .B(n33444), .Z(n33446) );
  XOR U33090 ( .A(n33452), .B(n33453), .Z(n31630) );
  AND U33091 ( .A(n564), .B(n33454), .Z(n33453) );
  XOR U33092 ( .A(n33455), .B(n33452), .Z(n33454) );
  XOR U33093 ( .A(n33456), .B(n33457), .Z(n33444) );
  AND U33094 ( .A(n33458), .B(n33459), .Z(n33457) );
  XOR U33095 ( .A(n33456), .B(n31645), .Z(n33459) );
  XOR U33096 ( .A(n33460), .B(n33461), .Z(n31645) );
  AND U33097 ( .A(n567), .B(n33462), .Z(n33461) );
  XOR U33098 ( .A(n33463), .B(n33460), .Z(n33462) );
  XNOR U33099 ( .A(n31642), .B(n33456), .Z(n33458) );
  XOR U33100 ( .A(n33464), .B(n33465), .Z(n31642) );
  AND U33101 ( .A(n564), .B(n33466), .Z(n33465) );
  XOR U33102 ( .A(n33467), .B(n33464), .Z(n33466) );
  XOR U33103 ( .A(n33468), .B(n33469), .Z(n33456) );
  AND U33104 ( .A(n33470), .B(n33471), .Z(n33469) );
  XOR U33105 ( .A(n33468), .B(n31657), .Z(n33471) );
  XOR U33106 ( .A(n33472), .B(n33473), .Z(n31657) );
  AND U33107 ( .A(n567), .B(n33474), .Z(n33473) );
  XOR U33108 ( .A(n33475), .B(n33472), .Z(n33474) );
  XNOR U33109 ( .A(n31654), .B(n33468), .Z(n33470) );
  XOR U33110 ( .A(n33476), .B(n33477), .Z(n31654) );
  AND U33111 ( .A(n564), .B(n33478), .Z(n33477) );
  XOR U33112 ( .A(n33479), .B(n33476), .Z(n33478) );
  XOR U33113 ( .A(n33480), .B(n33481), .Z(n33468) );
  AND U33114 ( .A(n33482), .B(n33483), .Z(n33481) );
  XOR U33115 ( .A(n33480), .B(n31669), .Z(n33483) );
  XOR U33116 ( .A(n33484), .B(n33485), .Z(n31669) );
  AND U33117 ( .A(n567), .B(n33486), .Z(n33485) );
  XOR U33118 ( .A(n33487), .B(n33484), .Z(n33486) );
  XNOR U33119 ( .A(n31666), .B(n33480), .Z(n33482) );
  XOR U33120 ( .A(n33488), .B(n33489), .Z(n31666) );
  AND U33121 ( .A(n564), .B(n33490), .Z(n33489) );
  XOR U33122 ( .A(n33491), .B(n33488), .Z(n33490) );
  XOR U33123 ( .A(n33492), .B(n33493), .Z(n33480) );
  AND U33124 ( .A(n33494), .B(n33495), .Z(n33493) );
  XOR U33125 ( .A(n33492), .B(n31681), .Z(n33495) );
  XOR U33126 ( .A(n33496), .B(n33497), .Z(n31681) );
  AND U33127 ( .A(n567), .B(n33498), .Z(n33497) );
  XOR U33128 ( .A(n33499), .B(n33496), .Z(n33498) );
  XNOR U33129 ( .A(n31678), .B(n33492), .Z(n33494) );
  XOR U33130 ( .A(n33500), .B(n33501), .Z(n31678) );
  AND U33131 ( .A(n564), .B(n33502), .Z(n33501) );
  XOR U33132 ( .A(n33503), .B(n33500), .Z(n33502) );
  XOR U33133 ( .A(n33504), .B(n33505), .Z(n33492) );
  AND U33134 ( .A(n33506), .B(n33507), .Z(n33505) );
  XOR U33135 ( .A(n33504), .B(n31693), .Z(n33507) );
  XOR U33136 ( .A(n33508), .B(n33509), .Z(n31693) );
  AND U33137 ( .A(n567), .B(n33510), .Z(n33509) );
  XOR U33138 ( .A(n33511), .B(n33508), .Z(n33510) );
  XNOR U33139 ( .A(n31690), .B(n33504), .Z(n33506) );
  XOR U33140 ( .A(n33512), .B(n33513), .Z(n31690) );
  AND U33141 ( .A(n564), .B(n33514), .Z(n33513) );
  XOR U33142 ( .A(n33515), .B(n33512), .Z(n33514) );
  XOR U33143 ( .A(n33516), .B(n33517), .Z(n33504) );
  AND U33144 ( .A(n33518), .B(n33519), .Z(n33517) );
  XOR U33145 ( .A(n33516), .B(n31705), .Z(n33519) );
  XOR U33146 ( .A(n33520), .B(n33521), .Z(n31705) );
  AND U33147 ( .A(n567), .B(n33522), .Z(n33521) );
  XOR U33148 ( .A(n33523), .B(n33520), .Z(n33522) );
  XNOR U33149 ( .A(n31702), .B(n33516), .Z(n33518) );
  XOR U33150 ( .A(n33524), .B(n33525), .Z(n31702) );
  AND U33151 ( .A(n564), .B(n33526), .Z(n33525) );
  XOR U33152 ( .A(n33527), .B(n33524), .Z(n33526) );
  XOR U33153 ( .A(n33528), .B(n33529), .Z(n33516) );
  AND U33154 ( .A(n33530), .B(n33531), .Z(n33529) );
  XOR U33155 ( .A(n33528), .B(n31717), .Z(n33531) );
  XOR U33156 ( .A(n33532), .B(n33533), .Z(n31717) );
  AND U33157 ( .A(n567), .B(n33534), .Z(n33533) );
  XOR U33158 ( .A(n33535), .B(n33532), .Z(n33534) );
  XNOR U33159 ( .A(n31714), .B(n33528), .Z(n33530) );
  XOR U33160 ( .A(n33536), .B(n33537), .Z(n31714) );
  AND U33161 ( .A(n564), .B(n33538), .Z(n33537) );
  XOR U33162 ( .A(n33539), .B(n33536), .Z(n33538) );
  XOR U33163 ( .A(n33540), .B(n33541), .Z(n33528) );
  AND U33164 ( .A(n33542), .B(n33543), .Z(n33541) );
  XOR U33165 ( .A(n33540), .B(n31729), .Z(n33543) );
  XOR U33166 ( .A(n33544), .B(n33545), .Z(n31729) );
  AND U33167 ( .A(n567), .B(n33546), .Z(n33545) );
  XOR U33168 ( .A(n33547), .B(n33544), .Z(n33546) );
  XNOR U33169 ( .A(n31726), .B(n33540), .Z(n33542) );
  XOR U33170 ( .A(n33548), .B(n33549), .Z(n31726) );
  AND U33171 ( .A(n564), .B(n33550), .Z(n33549) );
  XOR U33172 ( .A(n33551), .B(n33548), .Z(n33550) );
  XOR U33173 ( .A(n33552), .B(n33553), .Z(n33540) );
  AND U33174 ( .A(n33554), .B(n33555), .Z(n33553) );
  XOR U33175 ( .A(n33552), .B(n31741), .Z(n33555) );
  XOR U33176 ( .A(n33556), .B(n33557), .Z(n31741) );
  AND U33177 ( .A(n567), .B(n33558), .Z(n33557) );
  XOR U33178 ( .A(n33559), .B(n33556), .Z(n33558) );
  XNOR U33179 ( .A(n31738), .B(n33552), .Z(n33554) );
  XOR U33180 ( .A(n33560), .B(n33561), .Z(n31738) );
  AND U33181 ( .A(n564), .B(n33562), .Z(n33561) );
  XOR U33182 ( .A(n33563), .B(n33560), .Z(n33562) );
  XOR U33183 ( .A(n33564), .B(n33565), .Z(n33552) );
  AND U33184 ( .A(n33566), .B(n33567), .Z(n33565) );
  XOR U33185 ( .A(n33564), .B(n31753), .Z(n33567) );
  XOR U33186 ( .A(n33568), .B(n33569), .Z(n31753) );
  AND U33187 ( .A(n567), .B(n33570), .Z(n33569) );
  XOR U33188 ( .A(n33571), .B(n33568), .Z(n33570) );
  XNOR U33189 ( .A(n31750), .B(n33564), .Z(n33566) );
  XOR U33190 ( .A(n33572), .B(n33573), .Z(n31750) );
  AND U33191 ( .A(n564), .B(n33574), .Z(n33573) );
  XOR U33192 ( .A(n33575), .B(n33572), .Z(n33574) );
  XOR U33193 ( .A(n33576), .B(n33577), .Z(n33564) );
  AND U33194 ( .A(n33578), .B(n33579), .Z(n33577) );
  XOR U33195 ( .A(n33576), .B(n31765), .Z(n33579) );
  XOR U33196 ( .A(n33580), .B(n33581), .Z(n31765) );
  AND U33197 ( .A(n567), .B(n33582), .Z(n33581) );
  XOR U33198 ( .A(n33583), .B(n33580), .Z(n33582) );
  XNOR U33199 ( .A(n31762), .B(n33576), .Z(n33578) );
  XOR U33200 ( .A(n33584), .B(n33585), .Z(n31762) );
  AND U33201 ( .A(n564), .B(n33586), .Z(n33585) );
  XOR U33202 ( .A(n33587), .B(n33584), .Z(n33586) );
  XOR U33203 ( .A(n33588), .B(n33589), .Z(n33576) );
  AND U33204 ( .A(n33590), .B(n33591), .Z(n33589) );
  XOR U33205 ( .A(n33588), .B(n31777), .Z(n33591) );
  XOR U33206 ( .A(n33592), .B(n33593), .Z(n31777) );
  AND U33207 ( .A(n567), .B(n33594), .Z(n33593) );
  XOR U33208 ( .A(n33595), .B(n33592), .Z(n33594) );
  XNOR U33209 ( .A(n31774), .B(n33588), .Z(n33590) );
  XOR U33210 ( .A(n33596), .B(n33597), .Z(n31774) );
  AND U33211 ( .A(n564), .B(n33598), .Z(n33597) );
  XOR U33212 ( .A(n33599), .B(n33596), .Z(n33598) );
  XOR U33213 ( .A(n33600), .B(n33601), .Z(n33588) );
  AND U33214 ( .A(n33602), .B(n33603), .Z(n33601) );
  XOR U33215 ( .A(n33600), .B(n31789), .Z(n33603) );
  XOR U33216 ( .A(n33604), .B(n33605), .Z(n31789) );
  AND U33217 ( .A(n567), .B(n33606), .Z(n33605) );
  XOR U33218 ( .A(n33607), .B(n33604), .Z(n33606) );
  XNOR U33219 ( .A(n31786), .B(n33600), .Z(n33602) );
  XOR U33220 ( .A(n33608), .B(n33609), .Z(n31786) );
  AND U33221 ( .A(n564), .B(n33610), .Z(n33609) );
  XOR U33222 ( .A(n33611), .B(n33608), .Z(n33610) );
  XOR U33223 ( .A(n33612), .B(n33613), .Z(n33600) );
  AND U33224 ( .A(n33614), .B(n33615), .Z(n33613) );
  XNOR U33225 ( .A(n33616), .B(n31802), .Z(n33615) );
  XOR U33226 ( .A(n33617), .B(n33618), .Z(n31802) );
  AND U33227 ( .A(n567), .B(n33619), .Z(n33618) );
  XOR U33228 ( .A(n33617), .B(n33620), .Z(n33619) );
  XNOR U33229 ( .A(n31799), .B(n33612), .Z(n33614) );
  XOR U33230 ( .A(n33621), .B(n33622), .Z(n31799) );
  AND U33231 ( .A(n564), .B(n33623), .Z(n33622) );
  XOR U33232 ( .A(n33621), .B(n33624), .Z(n33623) );
  IV U33233 ( .A(n33616), .Z(n33612) );
  AND U33234 ( .A(n33248), .B(n33251), .Z(n33616) );
  XNOR U33235 ( .A(n33625), .B(n33626), .Z(n33251) );
  AND U33236 ( .A(n567), .B(n33627), .Z(n33626) );
  XNOR U33237 ( .A(n33628), .B(n33625), .Z(n33627) );
  XOR U33238 ( .A(n33629), .B(n33630), .Z(n567) );
  AND U33239 ( .A(n33631), .B(n33632), .Z(n33630) );
  XOR U33240 ( .A(n33259), .B(n33629), .Z(n33632) );
  IV U33241 ( .A(n33633), .Z(n33259) );
  AND U33242 ( .A(p_input[3839]), .B(p_input[3807]), .Z(n33633) );
  XOR U33243 ( .A(n33629), .B(n33256), .Z(n33631) );
  AND U33244 ( .A(p_input[3743]), .B(p_input[3775]), .Z(n33256) );
  XOR U33245 ( .A(n33634), .B(n33635), .Z(n33629) );
  AND U33246 ( .A(n33636), .B(n33637), .Z(n33635) );
  XOR U33247 ( .A(n33634), .B(n33271), .Z(n33637) );
  XNOR U33248 ( .A(p_input[3806]), .B(n33638), .Z(n33271) );
  AND U33249 ( .A(n703), .B(n33639), .Z(n33638) );
  XOR U33250 ( .A(p_input[3838]), .B(p_input[3806]), .Z(n33639) );
  XNOR U33251 ( .A(n33268), .B(n33634), .Z(n33636) );
  XOR U33252 ( .A(n33640), .B(n33641), .Z(n33268) );
  AND U33253 ( .A(n701), .B(n33642), .Z(n33641) );
  XOR U33254 ( .A(p_input[3774]), .B(p_input[3742]), .Z(n33642) );
  XOR U33255 ( .A(n33643), .B(n33644), .Z(n33634) );
  AND U33256 ( .A(n33645), .B(n33646), .Z(n33644) );
  XOR U33257 ( .A(n33643), .B(n33283), .Z(n33646) );
  XNOR U33258 ( .A(p_input[3805]), .B(n33647), .Z(n33283) );
  AND U33259 ( .A(n703), .B(n33648), .Z(n33647) );
  XOR U33260 ( .A(p_input[3837]), .B(p_input[3805]), .Z(n33648) );
  XNOR U33261 ( .A(n33280), .B(n33643), .Z(n33645) );
  XOR U33262 ( .A(n33649), .B(n33650), .Z(n33280) );
  AND U33263 ( .A(n701), .B(n33651), .Z(n33650) );
  XOR U33264 ( .A(p_input[3773]), .B(p_input[3741]), .Z(n33651) );
  XOR U33265 ( .A(n33652), .B(n33653), .Z(n33643) );
  AND U33266 ( .A(n33654), .B(n33655), .Z(n33653) );
  XOR U33267 ( .A(n33652), .B(n33295), .Z(n33655) );
  XNOR U33268 ( .A(p_input[3804]), .B(n33656), .Z(n33295) );
  AND U33269 ( .A(n703), .B(n33657), .Z(n33656) );
  XOR U33270 ( .A(p_input[3836]), .B(p_input[3804]), .Z(n33657) );
  XNOR U33271 ( .A(n33292), .B(n33652), .Z(n33654) );
  XOR U33272 ( .A(n33658), .B(n33659), .Z(n33292) );
  AND U33273 ( .A(n701), .B(n33660), .Z(n33659) );
  XOR U33274 ( .A(p_input[3772]), .B(p_input[3740]), .Z(n33660) );
  XOR U33275 ( .A(n33661), .B(n33662), .Z(n33652) );
  AND U33276 ( .A(n33663), .B(n33664), .Z(n33662) );
  XOR U33277 ( .A(n33661), .B(n33307), .Z(n33664) );
  XNOR U33278 ( .A(p_input[3803]), .B(n33665), .Z(n33307) );
  AND U33279 ( .A(n703), .B(n33666), .Z(n33665) );
  XOR U33280 ( .A(p_input[3835]), .B(p_input[3803]), .Z(n33666) );
  XNOR U33281 ( .A(n33304), .B(n33661), .Z(n33663) );
  XOR U33282 ( .A(n33667), .B(n33668), .Z(n33304) );
  AND U33283 ( .A(n701), .B(n33669), .Z(n33668) );
  XOR U33284 ( .A(p_input[3771]), .B(p_input[3739]), .Z(n33669) );
  XOR U33285 ( .A(n33670), .B(n33671), .Z(n33661) );
  AND U33286 ( .A(n33672), .B(n33673), .Z(n33671) );
  XOR U33287 ( .A(n33670), .B(n33319), .Z(n33673) );
  XNOR U33288 ( .A(p_input[3802]), .B(n33674), .Z(n33319) );
  AND U33289 ( .A(n703), .B(n33675), .Z(n33674) );
  XOR U33290 ( .A(p_input[3834]), .B(p_input[3802]), .Z(n33675) );
  XNOR U33291 ( .A(n33316), .B(n33670), .Z(n33672) );
  XOR U33292 ( .A(n33676), .B(n33677), .Z(n33316) );
  AND U33293 ( .A(n701), .B(n33678), .Z(n33677) );
  XOR U33294 ( .A(p_input[3770]), .B(p_input[3738]), .Z(n33678) );
  XOR U33295 ( .A(n33679), .B(n33680), .Z(n33670) );
  AND U33296 ( .A(n33681), .B(n33682), .Z(n33680) );
  XOR U33297 ( .A(n33679), .B(n33331), .Z(n33682) );
  XNOR U33298 ( .A(p_input[3801]), .B(n33683), .Z(n33331) );
  AND U33299 ( .A(n703), .B(n33684), .Z(n33683) );
  XOR U33300 ( .A(p_input[3833]), .B(p_input[3801]), .Z(n33684) );
  XNOR U33301 ( .A(n33328), .B(n33679), .Z(n33681) );
  XOR U33302 ( .A(n33685), .B(n33686), .Z(n33328) );
  AND U33303 ( .A(n701), .B(n33687), .Z(n33686) );
  XOR U33304 ( .A(p_input[3769]), .B(p_input[3737]), .Z(n33687) );
  XOR U33305 ( .A(n33688), .B(n33689), .Z(n33679) );
  AND U33306 ( .A(n33690), .B(n33691), .Z(n33689) );
  XOR U33307 ( .A(n33688), .B(n33343), .Z(n33691) );
  XNOR U33308 ( .A(p_input[3800]), .B(n33692), .Z(n33343) );
  AND U33309 ( .A(n703), .B(n33693), .Z(n33692) );
  XOR U33310 ( .A(p_input[3832]), .B(p_input[3800]), .Z(n33693) );
  XNOR U33311 ( .A(n33340), .B(n33688), .Z(n33690) );
  XOR U33312 ( .A(n33694), .B(n33695), .Z(n33340) );
  AND U33313 ( .A(n701), .B(n33696), .Z(n33695) );
  XOR U33314 ( .A(p_input[3768]), .B(p_input[3736]), .Z(n33696) );
  XOR U33315 ( .A(n33697), .B(n33698), .Z(n33688) );
  AND U33316 ( .A(n33699), .B(n33700), .Z(n33698) );
  XOR U33317 ( .A(n33697), .B(n33355), .Z(n33700) );
  XNOR U33318 ( .A(p_input[3799]), .B(n33701), .Z(n33355) );
  AND U33319 ( .A(n703), .B(n33702), .Z(n33701) );
  XOR U33320 ( .A(p_input[3831]), .B(p_input[3799]), .Z(n33702) );
  XNOR U33321 ( .A(n33352), .B(n33697), .Z(n33699) );
  XOR U33322 ( .A(n33703), .B(n33704), .Z(n33352) );
  AND U33323 ( .A(n701), .B(n33705), .Z(n33704) );
  XOR U33324 ( .A(p_input[3767]), .B(p_input[3735]), .Z(n33705) );
  XOR U33325 ( .A(n33706), .B(n33707), .Z(n33697) );
  AND U33326 ( .A(n33708), .B(n33709), .Z(n33707) );
  XOR U33327 ( .A(n33706), .B(n33367), .Z(n33709) );
  XNOR U33328 ( .A(p_input[3798]), .B(n33710), .Z(n33367) );
  AND U33329 ( .A(n703), .B(n33711), .Z(n33710) );
  XOR U33330 ( .A(p_input[3830]), .B(p_input[3798]), .Z(n33711) );
  XNOR U33331 ( .A(n33364), .B(n33706), .Z(n33708) );
  XOR U33332 ( .A(n33712), .B(n33713), .Z(n33364) );
  AND U33333 ( .A(n701), .B(n33714), .Z(n33713) );
  XOR U33334 ( .A(p_input[3766]), .B(p_input[3734]), .Z(n33714) );
  XOR U33335 ( .A(n33715), .B(n33716), .Z(n33706) );
  AND U33336 ( .A(n33717), .B(n33718), .Z(n33716) );
  XOR U33337 ( .A(n33715), .B(n33379), .Z(n33718) );
  XNOR U33338 ( .A(p_input[3797]), .B(n33719), .Z(n33379) );
  AND U33339 ( .A(n703), .B(n33720), .Z(n33719) );
  XOR U33340 ( .A(p_input[3829]), .B(p_input[3797]), .Z(n33720) );
  XNOR U33341 ( .A(n33376), .B(n33715), .Z(n33717) );
  XOR U33342 ( .A(n33721), .B(n33722), .Z(n33376) );
  AND U33343 ( .A(n701), .B(n33723), .Z(n33722) );
  XOR U33344 ( .A(p_input[3765]), .B(p_input[3733]), .Z(n33723) );
  XOR U33345 ( .A(n33724), .B(n33725), .Z(n33715) );
  AND U33346 ( .A(n33726), .B(n33727), .Z(n33725) );
  XOR U33347 ( .A(n33724), .B(n33391), .Z(n33727) );
  XNOR U33348 ( .A(p_input[3796]), .B(n33728), .Z(n33391) );
  AND U33349 ( .A(n703), .B(n33729), .Z(n33728) );
  XOR U33350 ( .A(p_input[3828]), .B(p_input[3796]), .Z(n33729) );
  XNOR U33351 ( .A(n33388), .B(n33724), .Z(n33726) );
  XOR U33352 ( .A(n33730), .B(n33731), .Z(n33388) );
  AND U33353 ( .A(n701), .B(n33732), .Z(n33731) );
  XOR U33354 ( .A(p_input[3764]), .B(p_input[3732]), .Z(n33732) );
  XOR U33355 ( .A(n33733), .B(n33734), .Z(n33724) );
  AND U33356 ( .A(n33735), .B(n33736), .Z(n33734) );
  XOR U33357 ( .A(n33733), .B(n33403), .Z(n33736) );
  XNOR U33358 ( .A(p_input[3795]), .B(n33737), .Z(n33403) );
  AND U33359 ( .A(n703), .B(n33738), .Z(n33737) );
  XOR U33360 ( .A(p_input[3827]), .B(p_input[3795]), .Z(n33738) );
  XNOR U33361 ( .A(n33400), .B(n33733), .Z(n33735) );
  XOR U33362 ( .A(n33739), .B(n33740), .Z(n33400) );
  AND U33363 ( .A(n701), .B(n33741), .Z(n33740) );
  XOR U33364 ( .A(p_input[3763]), .B(p_input[3731]), .Z(n33741) );
  XOR U33365 ( .A(n33742), .B(n33743), .Z(n33733) );
  AND U33366 ( .A(n33744), .B(n33745), .Z(n33743) );
  XOR U33367 ( .A(n33742), .B(n33415), .Z(n33745) );
  XNOR U33368 ( .A(p_input[3794]), .B(n33746), .Z(n33415) );
  AND U33369 ( .A(n703), .B(n33747), .Z(n33746) );
  XOR U33370 ( .A(p_input[3826]), .B(p_input[3794]), .Z(n33747) );
  XNOR U33371 ( .A(n33412), .B(n33742), .Z(n33744) );
  XOR U33372 ( .A(n33748), .B(n33749), .Z(n33412) );
  AND U33373 ( .A(n701), .B(n33750), .Z(n33749) );
  XOR U33374 ( .A(p_input[3762]), .B(p_input[3730]), .Z(n33750) );
  XOR U33375 ( .A(n33751), .B(n33752), .Z(n33742) );
  AND U33376 ( .A(n33753), .B(n33754), .Z(n33752) );
  XOR U33377 ( .A(n33751), .B(n33427), .Z(n33754) );
  XNOR U33378 ( .A(p_input[3793]), .B(n33755), .Z(n33427) );
  AND U33379 ( .A(n703), .B(n33756), .Z(n33755) );
  XOR U33380 ( .A(p_input[3825]), .B(p_input[3793]), .Z(n33756) );
  XNOR U33381 ( .A(n33424), .B(n33751), .Z(n33753) );
  XOR U33382 ( .A(n33757), .B(n33758), .Z(n33424) );
  AND U33383 ( .A(n701), .B(n33759), .Z(n33758) );
  XOR U33384 ( .A(p_input[3761]), .B(p_input[3729]), .Z(n33759) );
  XOR U33385 ( .A(n33760), .B(n33761), .Z(n33751) );
  AND U33386 ( .A(n33762), .B(n33763), .Z(n33761) );
  XOR U33387 ( .A(n33760), .B(n33439), .Z(n33763) );
  XNOR U33388 ( .A(p_input[3792]), .B(n33764), .Z(n33439) );
  AND U33389 ( .A(n703), .B(n33765), .Z(n33764) );
  XOR U33390 ( .A(p_input[3824]), .B(p_input[3792]), .Z(n33765) );
  XNOR U33391 ( .A(n33436), .B(n33760), .Z(n33762) );
  XOR U33392 ( .A(n33766), .B(n33767), .Z(n33436) );
  AND U33393 ( .A(n701), .B(n33768), .Z(n33767) );
  XOR U33394 ( .A(p_input[3760]), .B(p_input[3728]), .Z(n33768) );
  XOR U33395 ( .A(n33769), .B(n33770), .Z(n33760) );
  AND U33396 ( .A(n33771), .B(n33772), .Z(n33770) );
  XOR U33397 ( .A(n33769), .B(n33451), .Z(n33772) );
  XNOR U33398 ( .A(p_input[3791]), .B(n33773), .Z(n33451) );
  AND U33399 ( .A(n703), .B(n33774), .Z(n33773) );
  XOR U33400 ( .A(p_input[3823]), .B(p_input[3791]), .Z(n33774) );
  XNOR U33401 ( .A(n33448), .B(n33769), .Z(n33771) );
  XOR U33402 ( .A(n33775), .B(n33776), .Z(n33448) );
  AND U33403 ( .A(n701), .B(n33777), .Z(n33776) );
  XOR U33404 ( .A(p_input[3759]), .B(p_input[3727]), .Z(n33777) );
  XOR U33405 ( .A(n33778), .B(n33779), .Z(n33769) );
  AND U33406 ( .A(n33780), .B(n33781), .Z(n33779) );
  XOR U33407 ( .A(n33778), .B(n33463), .Z(n33781) );
  XNOR U33408 ( .A(p_input[3790]), .B(n33782), .Z(n33463) );
  AND U33409 ( .A(n703), .B(n33783), .Z(n33782) );
  XOR U33410 ( .A(p_input[3822]), .B(p_input[3790]), .Z(n33783) );
  XNOR U33411 ( .A(n33460), .B(n33778), .Z(n33780) );
  XOR U33412 ( .A(n33784), .B(n33785), .Z(n33460) );
  AND U33413 ( .A(n701), .B(n33786), .Z(n33785) );
  XOR U33414 ( .A(p_input[3758]), .B(p_input[3726]), .Z(n33786) );
  XOR U33415 ( .A(n33787), .B(n33788), .Z(n33778) );
  AND U33416 ( .A(n33789), .B(n33790), .Z(n33788) );
  XOR U33417 ( .A(n33787), .B(n33475), .Z(n33790) );
  XNOR U33418 ( .A(p_input[3789]), .B(n33791), .Z(n33475) );
  AND U33419 ( .A(n703), .B(n33792), .Z(n33791) );
  XOR U33420 ( .A(p_input[3821]), .B(p_input[3789]), .Z(n33792) );
  XNOR U33421 ( .A(n33472), .B(n33787), .Z(n33789) );
  XOR U33422 ( .A(n33793), .B(n33794), .Z(n33472) );
  AND U33423 ( .A(n701), .B(n33795), .Z(n33794) );
  XOR U33424 ( .A(p_input[3757]), .B(p_input[3725]), .Z(n33795) );
  XOR U33425 ( .A(n33796), .B(n33797), .Z(n33787) );
  AND U33426 ( .A(n33798), .B(n33799), .Z(n33797) );
  XOR U33427 ( .A(n33796), .B(n33487), .Z(n33799) );
  XNOR U33428 ( .A(p_input[3788]), .B(n33800), .Z(n33487) );
  AND U33429 ( .A(n703), .B(n33801), .Z(n33800) );
  XOR U33430 ( .A(p_input[3820]), .B(p_input[3788]), .Z(n33801) );
  XNOR U33431 ( .A(n33484), .B(n33796), .Z(n33798) );
  XOR U33432 ( .A(n33802), .B(n33803), .Z(n33484) );
  AND U33433 ( .A(n701), .B(n33804), .Z(n33803) );
  XOR U33434 ( .A(p_input[3756]), .B(p_input[3724]), .Z(n33804) );
  XOR U33435 ( .A(n33805), .B(n33806), .Z(n33796) );
  AND U33436 ( .A(n33807), .B(n33808), .Z(n33806) );
  XOR U33437 ( .A(n33805), .B(n33499), .Z(n33808) );
  XNOR U33438 ( .A(p_input[3787]), .B(n33809), .Z(n33499) );
  AND U33439 ( .A(n703), .B(n33810), .Z(n33809) );
  XOR U33440 ( .A(p_input[3819]), .B(p_input[3787]), .Z(n33810) );
  XNOR U33441 ( .A(n33496), .B(n33805), .Z(n33807) );
  XOR U33442 ( .A(n33811), .B(n33812), .Z(n33496) );
  AND U33443 ( .A(n701), .B(n33813), .Z(n33812) );
  XOR U33444 ( .A(p_input[3755]), .B(p_input[3723]), .Z(n33813) );
  XOR U33445 ( .A(n33814), .B(n33815), .Z(n33805) );
  AND U33446 ( .A(n33816), .B(n33817), .Z(n33815) );
  XOR U33447 ( .A(n33814), .B(n33511), .Z(n33817) );
  XNOR U33448 ( .A(p_input[3786]), .B(n33818), .Z(n33511) );
  AND U33449 ( .A(n703), .B(n33819), .Z(n33818) );
  XOR U33450 ( .A(p_input[3818]), .B(p_input[3786]), .Z(n33819) );
  XNOR U33451 ( .A(n33508), .B(n33814), .Z(n33816) );
  XOR U33452 ( .A(n33820), .B(n33821), .Z(n33508) );
  AND U33453 ( .A(n701), .B(n33822), .Z(n33821) );
  XOR U33454 ( .A(p_input[3754]), .B(p_input[3722]), .Z(n33822) );
  XOR U33455 ( .A(n33823), .B(n33824), .Z(n33814) );
  AND U33456 ( .A(n33825), .B(n33826), .Z(n33824) );
  XOR U33457 ( .A(n33823), .B(n33523), .Z(n33826) );
  XNOR U33458 ( .A(p_input[3785]), .B(n33827), .Z(n33523) );
  AND U33459 ( .A(n703), .B(n33828), .Z(n33827) );
  XOR U33460 ( .A(p_input[3817]), .B(p_input[3785]), .Z(n33828) );
  XNOR U33461 ( .A(n33520), .B(n33823), .Z(n33825) );
  XOR U33462 ( .A(n33829), .B(n33830), .Z(n33520) );
  AND U33463 ( .A(n701), .B(n33831), .Z(n33830) );
  XOR U33464 ( .A(p_input[3753]), .B(p_input[3721]), .Z(n33831) );
  XOR U33465 ( .A(n33832), .B(n33833), .Z(n33823) );
  AND U33466 ( .A(n33834), .B(n33835), .Z(n33833) );
  XOR U33467 ( .A(n33832), .B(n33535), .Z(n33835) );
  XNOR U33468 ( .A(p_input[3784]), .B(n33836), .Z(n33535) );
  AND U33469 ( .A(n703), .B(n33837), .Z(n33836) );
  XOR U33470 ( .A(p_input[3816]), .B(p_input[3784]), .Z(n33837) );
  XNOR U33471 ( .A(n33532), .B(n33832), .Z(n33834) );
  XOR U33472 ( .A(n33838), .B(n33839), .Z(n33532) );
  AND U33473 ( .A(n701), .B(n33840), .Z(n33839) );
  XOR U33474 ( .A(p_input[3752]), .B(p_input[3720]), .Z(n33840) );
  XOR U33475 ( .A(n33841), .B(n33842), .Z(n33832) );
  AND U33476 ( .A(n33843), .B(n33844), .Z(n33842) );
  XOR U33477 ( .A(n33841), .B(n33547), .Z(n33844) );
  XNOR U33478 ( .A(p_input[3783]), .B(n33845), .Z(n33547) );
  AND U33479 ( .A(n703), .B(n33846), .Z(n33845) );
  XOR U33480 ( .A(p_input[3815]), .B(p_input[3783]), .Z(n33846) );
  XNOR U33481 ( .A(n33544), .B(n33841), .Z(n33843) );
  XOR U33482 ( .A(n33847), .B(n33848), .Z(n33544) );
  AND U33483 ( .A(n701), .B(n33849), .Z(n33848) );
  XOR U33484 ( .A(p_input[3751]), .B(p_input[3719]), .Z(n33849) );
  XOR U33485 ( .A(n33850), .B(n33851), .Z(n33841) );
  AND U33486 ( .A(n33852), .B(n33853), .Z(n33851) );
  XOR U33487 ( .A(n33850), .B(n33559), .Z(n33853) );
  XNOR U33488 ( .A(p_input[3782]), .B(n33854), .Z(n33559) );
  AND U33489 ( .A(n703), .B(n33855), .Z(n33854) );
  XOR U33490 ( .A(p_input[3814]), .B(p_input[3782]), .Z(n33855) );
  XNOR U33491 ( .A(n33556), .B(n33850), .Z(n33852) );
  XOR U33492 ( .A(n33856), .B(n33857), .Z(n33556) );
  AND U33493 ( .A(n701), .B(n33858), .Z(n33857) );
  XOR U33494 ( .A(p_input[3750]), .B(p_input[3718]), .Z(n33858) );
  XOR U33495 ( .A(n33859), .B(n33860), .Z(n33850) );
  AND U33496 ( .A(n33861), .B(n33862), .Z(n33860) );
  XOR U33497 ( .A(n33859), .B(n33571), .Z(n33862) );
  XNOR U33498 ( .A(p_input[3781]), .B(n33863), .Z(n33571) );
  AND U33499 ( .A(n703), .B(n33864), .Z(n33863) );
  XOR U33500 ( .A(p_input[3813]), .B(p_input[3781]), .Z(n33864) );
  XNOR U33501 ( .A(n33568), .B(n33859), .Z(n33861) );
  XOR U33502 ( .A(n33865), .B(n33866), .Z(n33568) );
  AND U33503 ( .A(n701), .B(n33867), .Z(n33866) );
  XOR U33504 ( .A(p_input[3749]), .B(p_input[3717]), .Z(n33867) );
  XOR U33505 ( .A(n33868), .B(n33869), .Z(n33859) );
  AND U33506 ( .A(n33870), .B(n33871), .Z(n33869) );
  XOR U33507 ( .A(n33868), .B(n33583), .Z(n33871) );
  XNOR U33508 ( .A(p_input[3780]), .B(n33872), .Z(n33583) );
  AND U33509 ( .A(n703), .B(n33873), .Z(n33872) );
  XOR U33510 ( .A(p_input[3812]), .B(p_input[3780]), .Z(n33873) );
  XNOR U33511 ( .A(n33580), .B(n33868), .Z(n33870) );
  XOR U33512 ( .A(n33874), .B(n33875), .Z(n33580) );
  AND U33513 ( .A(n701), .B(n33876), .Z(n33875) );
  XOR U33514 ( .A(p_input[3748]), .B(p_input[3716]), .Z(n33876) );
  XOR U33515 ( .A(n33877), .B(n33878), .Z(n33868) );
  AND U33516 ( .A(n33879), .B(n33880), .Z(n33878) );
  XOR U33517 ( .A(n33877), .B(n33595), .Z(n33880) );
  XNOR U33518 ( .A(p_input[3779]), .B(n33881), .Z(n33595) );
  AND U33519 ( .A(n703), .B(n33882), .Z(n33881) );
  XOR U33520 ( .A(p_input[3811]), .B(p_input[3779]), .Z(n33882) );
  XNOR U33521 ( .A(n33592), .B(n33877), .Z(n33879) );
  XOR U33522 ( .A(n33883), .B(n33884), .Z(n33592) );
  AND U33523 ( .A(n701), .B(n33885), .Z(n33884) );
  XOR U33524 ( .A(p_input[3747]), .B(p_input[3715]), .Z(n33885) );
  XOR U33525 ( .A(n33886), .B(n33887), .Z(n33877) );
  AND U33526 ( .A(n33888), .B(n33889), .Z(n33887) );
  XOR U33527 ( .A(n33886), .B(n33607), .Z(n33889) );
  XNOR U33528 ( .A(p_input[3778]), .B(n33890), .Z(n33607) );
  AND U33529 ( .A(n703), .B(n33891), .Z(n33890) );
  XOR U33530 ( .A(p_input[3810]), .B(p_input[3778]), .Z(n33891) );
  XNOR U33531 ( .A(n33604), .B(n33886), .Z(n33888) );
  XOR U33532 ( .A(n33892), .B(n33893), .Z(n33604) );
  AND U33533 ( .A(n701), .B(n33894), .Z(n33893) );
  XOR U33534 ( .A(p_input[3746]), .B(p_input[3714]), .Z(n33894) );
  XOR U33535 ( .A(n33895), .B(n33896), .Z(n33886) );
  AND U33536 ( .A(n33897), .B(n33898), .Z(n33896) );
  XNOR U33537 ( .A(n33899), .B(n33620), .Z(n33898) );
  XNOR U33538 ( .A(p_input[3777]), .B(n33900), .Z(n33620) );
  AND U33539 ( .A(n703), .B(n33901), .Z(n33900) );
  XNOR U33540 ( .A(p_input[3809]), .B(n33902), .Z(n33901) );
  IV U33541 ( .A(p_input[3777]), .Z(n33902) );
  XNOR U33542 ( .A(n33617), .B(n33895), .Z(n33897) );
  XNOR U33543 ( .A(p_input[3713]), .B(n33903), .Z(n33617) );
  AND U33544 ( .A(n701), .B(n33904), .Z(n33903) );
  XOR U33545 ( .A(p_input[3745]), .B(p_input[3713]), .Z(n33904) );
  IV U33546 ( .A(n33899), .Z(n33895) );
  AND U33547 ( .A(n33625), .B(n33628), .Z(n33899) );
  XOR U33548 ( .A(p_input[3776]), .B(n33905), .Z(n33628) );
  AND U33549 ( .A(n703), .B(n33906), .Z(n33905) );
  XOR U33550 ( .A(p_input[3808]), .B(p_input[3776]), .Z(n33906) );
  XOR U33551 ( .A(n33907), .B(n33908), .Z(n703) );
  AND U33552 ( .A(n33909), .B(n33910), .Z(n33908) );
  XNOR U33553 ( .A(p_input[3839]), .B(n33907), .Z(n33910) );
  XOR U33554 ( .A(n33907), .B(p_input[3807]), .Z(n33909) );
  XOR U33555 ( .A(n33911), .B(n33912), .Z(n33907) );
  AND U33556 ( .A(n33913), .B(n33914), .Z(n33912) );
  XNOR U33557 ( .A(p_input[3838]), .B(n33911), .Z(n33914) );
  XOR U33558 ( .A(n33911), .B(p_input[3806]), .Z(n33913) );
  XOR U33559 ( .A(n33915), .B(n33916), .Z(n33911) );
  AND U33560 ( .A(n33917), .B(n33918), .Z(n33916) );
  XNOR U33561 ( .A(p_input[3837]), .B(n33915), .Z(n33918) );
  XOR U33562 ( .A(n33915), .B(p_input[3805]), .Z(n33917) );
  XOR U33563 ( .A(n33919), .B(n33920), .Z(n33915) );
  AND U33564 ( .A(n33921), .B(n33922), .Z(n33920) );
  XNOR U33565 ( .A(p_input[3836]), .B(n33919), .Z(n33922) );
  XOR U33566 ( .A(n33919), .B(p_input[3804]), .Z(n33921) );
  XOR U33567 ( .A(n33923), .B(n33924), .Z(n33919) );
  AND U33568 ( .A(n33925), .B(n33926), .Z(n33924) );
  XNOR U33569 ( .A(p_input[3835]), .B(n33923), .Z(n33926) );
  XOR U33570 ( .A(n33923), .B(p_input[3803]), .Z(n33925) );
  XOR U33571 ( .A(n33927), .B(n33928), .Z(n33923) );
  AND U33572 ( .A(n33929), .B(n33930), .Z(n33928) );
  XNOR U33573 ( .A(p_input[3834]), .B(n33927), .Z(n33930) );
  XOR U33574 ( .A(n33927), .B(p_input[3802]), .Z(n33929) );
  XOR U33575 ( .A(n33931), .B(n33932), .Z(n33927) );
  AND U33576 ( .A(n33933), .B(n33934), .Z(n33932) );
  XNOR U33577 ( .A(p_input[3833]), .B(n33931), .Z(n33934) );
  XOR U33578 ( .A(n33931), .B(p_input[3801]), .Z(n33933) );
  XOR U33579 ( .A(n33935), .B(n33936), .Z(n33931) );
  AND U33580 ( .A(n33937), .B(n33938), .Z(n33936) );
  XNOR U33581 ( .A(p_input[3832]), .B(n33935), .Z(n33938) );
  XOR U33582 ( .A(n33935), .B(p_input[3800]), .Z(n33937) );
  XOR U33583 ( .A(n33939), .B(n33940), .Z(n33935) );
  AND U33584 ( .A(n33941), .B(n33942), .Z(n33940) );
  XNOR U33585 ( .A(p_input[3831]), .B(n33939), .Z(n33942) );
  XOR U33586 ( .A(n33939), .B(p_input[3799]), .Z(n33941) );
  XOR U33587 ( .A(n33943), .B(n33944), .Z(n33939) );
  AND U33588 ( .A(n33945), .B(n33946), .Z(n33944) );
  XNOR U33589 ( .A(p_input[3830]), .B(n33943), .Z(n33946) );
  XOR U33590 ( .A(n33943), .B(p_input[3798]), .Z(n33945) );
  XOR U33591 ( .A(n33947), .B(n33948), .Z(n33943) );
  AND U33592 ( .A(n33949), .B(n33950), .Z(n33948) );
  XNOR U33593 ( .A(p_input[3829]), .B(n33947), .Z(n33950) );
  XOR U33594 ( .A(n33947), .B(p_input[3797]), .Z(n33949) );
  XOR U33595 ( .A(n33951), .B(n33952), .Z(n33947) );
  AND U33596 ( .A(n33953), .B(n33954), .Z(n33952) );
  XNOR U33597 ( .A(p_input[3828]), .B(n33951), .Z(n33954) );
  XOR U33598 ( .A(n33951), .B(p_input[3796]), .Z(n33953) );
  XOR U33599 ( .A(n33955), .B(n33956), .Z(n33951) );
  AND U33600 ( .A(n33957), .B(n33958), .Z(n33956) );
  XNOR U33601 ( .A(p_input[3827]), .B(n33955), .Z(n33958) );
  XOR U33602 ( .A(n33955), .B(p_input[3795]), .Z(n33957) );
  XOR U33603 ( .A(n33959), .B(n33960), .Z(n33955) );
  AND U33604 ( .A(n33961), .B(n33962), .Z(n33960) );
  XNOR U33605 ( .A(p_input[3826]), .B(n33959), .Z(n33962) );
  XOR U33606 ( .A(n33959), .B(p_input[3794]), .Z(n33961) );
  XOR U33607 ( .A(n33963), .B(n33964), .Z(n33959) );
  AND U33608 ( .A(n33965), .B(n33966), .Z(n33964) );
  XNOR U33609 ( .A(p_input[3825]), .B(n33963), .Z(n33966) );
  XOR U33610 ( .A(n33963), .B(p_input[3793]), .Z(n33965) );
  XOR U33611 ( .A(n33967), .B(n33968), .Z(n33963) );
  AND U33612 ( .A(n33969), .B(n33970), .Z(n33968) );
  XNOR U33613 ( .A(p_input[3824]), .B(n33967), .Z(n33970) );
  XOR U33614 ( .A(n33967), .B(p_input[3792]), .Z(n33969) );
  XOR U33615 ( .A(n33971), .B(n33972), .Z(n33967) );
  AND U33616 ( .A(n33973), .B(n33974), .Z(n33972) );
  XNOR U33617 ( .A(p_input[3823]), .B(n33971), .Z(n33974) );
  XOR U33618 ( .A(n33971), .B(p_input[3791]), .Z(n33973) );
  XOR U33619 ( .A(n33975), .B(n33976), .Z(n33971) );
  AND U33620 ( .A(n33977), .B(n33978), .Z(n33976) );
  XNOR U33621 ( .A(p_input[3822]), .B(n33975), .Z(n33978) );
  XOR U33622 ( .A(n33975), .B(p_input[3790]), .Z(n33977) );
  XOR U33623 ( .A(n33979), .B(n33980), .Z(n33975) );
  AND U33624 ( .A(n33981), .B(n33982), .Z(n33980) );
  XNOR U33625 ( .A(p_input[3821]), .B(n33979), .Z(n33982) );
  XOR U33626 ( .A(n33979), .B(p_input[3789]), .Z(n33981) );
  XOR U33627 ( .A(n33983), .B(n33984), .Z(n33979) );
  AND U33628 ( .A(n33985), .B(n33986), .Z(n33984) );
  XNOR U33629 ( .A(p_input[3820]), .B(n33983), .Z(n33986) );
  XOR U33630 ( .A(n33983), .B(p_input[3788]), .Z(n33985) );
  XOR U33631 ( .A(n33987), .B(n33988), .Z(n33983) );
  AND U33632 ( .A(n33989), .B(n33990), .Z(n33988) );
  XNOR U33633 ( .A(p_input[3819]), .B(n33987), .Z(n33990) );
  XOR U33634 ( .A(n33987), .B(p_input[3787]), .Z(n33989) );
  XOR U33635 ( .A(n33991), .B(n33992), .Z(n33987) );
  AND U33636 ( .A(n33993), .B(n33994), .Z(n33992) );
  XNOR U33637 ( .A(p_input[3818]), .B(n33991), .Z(n33994) );
  XOR U33638 ( .A(n33991), .B(p_input[3786]), .Z(n33993) );
  XOR U33639 ( .A(n33995), .B(n33996), .Z(n33991) );
  AND U33640 ( .A(n33997), .B(n33998), .Z(n33996) );
  XNOR U33641 ( .A(p_input[3817]), .B(n33995), .Z(n33998) );
  XOR U33642 ( .A(n33995), .B(p_input[3785]), .Z(n33997) );
  XOR U33643 ( .A(n33999), .B(n34000), .Z(n33995) );
  AND U33644 ( .A(n34001), .B(n34002), .Z(n34000) );
  XNOR U33645 ( .A(p_input[3816]), .B(n33999), .Z(n34002) );
  XOR U33646 ( .A(n33999), .B(p_input[3784]), .Z(n34001) );
  XOR U33647 ( .A(n34003), .B(n34004), .Z(n33999) );
  AND U33648 ( .A(n34005), .B(n34006), .Z(n34004) );
  XNOR U33649 ( .A(p_input[3815]), .B(n34003), .Z(n34006) );
  XOR U33650 ( .A(n34003), .B(p_input[3783]), .Z(n34005) );
  XOR U33651 ( .A(n34007), .B(n34008), .Z(n34003) );
  AND U33652 ( .A(n34009), .B(n34010), .Z(n34008) );
  XNOR U33653 ( .A(p_input[3814]), .B(n34007), .Z(n34010) );
  XOR U33654 ( .A(n34007), .B(p_input[3782]), .Z(n34009) );
  XOR U33655 ( .A(n34011), .B(n34012), .Z(n34007) );
  AND U33656 ( .A(n34013), .B(n34014), .Z(n34012) );
  XNOR U33657 ( .A(p_input[3813]), .B(n34011), .Z(n34014) );
  XOR U33658 ( .A(n34011), .B(p_input[3781]), .Z(n34013) );
  XOR U33659 ( .A(n34015), .B(n34016), .Z(n34011) );
  AND U33660 ( .A(n34017), .B(n34018), .Z(n34016) );
  XNOR U33661 ( .A(p_input[3812]), .B(n34015), .Z(n34018) );
  XOR U33662 ( .A(n34015), .B(p_input[3780]), .Z(n34017) );
  XOR U33663 ( .A(n34019), .B(n34020), .Z(n34015) );
  AND U33664 ( .A(n34021), .B(n34022), .Z(n34020) );
  XNOR U33665 ( .A(p_input[3811]), .B(n34019), .Z(n34022) );
  XOR U33666 ( .A(n34019), .B(p_input[3779]), .Z(n34021) );
  XOR U33667 ( .A(n34023), .B(n34024), .Z(n34019) );
  AND U33668 ( .A(n34025), .B(n34026), .Z(n34024) );
  XNOR U33669 ( .A(p_input[3810]), .B(n34023), .Z(n34026) );
  XOR U33670 ( .A(n34023), .B(p_input[3778]), .Z(n34025) );
  XNOR U33671 ( .A(n34027), .B(n34028), .Z(n34023) );
  AND U33672 ( .A(n34029), .B(n34030), .Z(n34028) );
  XOR U33673 ( .A(p_input[3809]), .B(n34027), .Z(n34030) );
  XNOR U33674 ( .A(p_input[3777]), .B(n34027), .Z(n34029) );
  AND U33675 ( .A(p_input[3808]), .B(n34031), .Z(n34027) );
  IV U33676 ( .A(p_input[3776]), .Z(n34031) );
  XNOR U33677 ( .A(p_input[3712]), .B(n34032), .Z(n33625) );
  AND U33678 ( .A(n701), .B(n34033), .Z(n34032) );
  XOR U33679 ( .A(p_input[3744]), .B(p_input[3712]), .Z(n34033) );
  XOR U33680 ( .A(n34034), .B(n34035), .Z(n701) );
  AND U33681 ( .A(n34036), .B(n34037), .Z(n34035) );
  XNOR U33682 ( .A(p_input[3775]), .B(n34034), .Z(n34037) );
  XOR U33683 ( .A(n34034), .B(p_input[3743]), .Z(n34036) );
  XOR U33684 ( .A(n34038), .B(n34039), .Z(n34034) );
  AND U33685 ( .A(n34040), .B(n34041), .Z(n34039) );
  XNOR U33686 ( .A(p_input[3774]), .B(n34038), .Z(n34041) );
  XNOR U33687 ( .A(n34038), .B(n33640), .Z(n34040) );
  IV U33688 ( .A(p_input[3742]), .Z(n33640) );
  XOR U33689 ( .A(n34042), .B(n34043), .Z(n34038) );
  AND U33690 ( .A(n34044), .B(n34045), .Z(n34043) );
  XNOR U33691 ( .A(p_input[3773]), .B(n34042), .Z(n34045) );
  XNOR U33692 ( .A(n34042), .B(n33649), .Z(n34044) );
  IV U33693 ( .A(p_input[3741]), .Z(n33649) );
  XOR U33694 ( .A(n34046), .B(n34047), .Z(n34042) );
  AND U33695 ( .A(n34048), .B(n34049), .Z(n34047) );
  XNOR U33696 ( .A(p_input[3772]), .B(n34046), .Z(n34049) );
  XNOR U33697 ( .A(n34046), .B(n33658), .Z(n34048) );
  IV U33698 ( .A(p_input[3740]), .Z(n33658) );
  XOR U33699 ( .A(n34050), .B(n34051), .Z(n34046) );
  AND U33700 ( .A(n34052), .B(n34053), .Z(n34051) );
  XNOR U33701 ( .A(p_input[3771]), .B(n34050), .Z(n34053) );
  XNOR U33702 ( .A(n34050), .B(n33667), .Z(n34052) );
  IV U33703 ( .A(p_input[3739]), .Z(n33667) );
  XOR U33704 ( .A(n34054), .B(n34055), .Z(n34050) );
  AND U33705 ( .A(n34056), .B(n34057), .Z(n34055) );
  XNOR U33706 ( .A(p_input[3770]), .B(n34054), .Z(n34057) );
  XNOR U33707 ( .A(n34054), .B(n33676), .Z(n34056) );
  IV U33708 ( .A(p_input[3738]), .Z(n33676) );
  XOR U33709 ( .A(n34058), .B(n34059), .Z(n34054) );
  AND U33710 ( .A(n34060), .B(n34061), .Z(n34059) );
  XNOR U33711 ( .A(p_input[3769]), .B(n34058), .Z(n34061) );
  XNOR U33712 ( .A(n34058), .B(n33685), .Z(n34060) );
  IV U33713 ( .A(p_input[3737]), .Z(n33685) );
  XOR U33714 ( .A(n34062), .B(n34063), .Z(n34058) );
  AND U33715 ( .A(n34064), .B(n34065), .Z(n34063) );
  XNOR U33716 ( .A(p_input[3768]), .B(n34062), .Z(n34065) );
  XNOR U33717 ( .A(n34062), .B(n33694), .Z(n34064) );
  IV U33718 ( .A(p_input[3736]), .Z(n33694) );
  XOR U33719 ( .A(n34066), .B(n34067), .Z(n34062) );
  AND U33720 ( .A(n34068), .B(n34069), .Z(n34067) );
  XNOR U33721 ( .A(p_input[3767]), .B(n34066), .Z(n34069) );
  XNOR U33722 ( .A(n34066), .B(n33703), .Z(n34068) );
  IV U33723 ( .A(p_input[3735]), .Z(n33703) );
  XOR U33724 ( .A(n34070), .B(n34071), .Z(n34066) );
  AND U33725 ( .A(n34072), .B(n34073), .Z(n34071) );
  XNOR U33726 ( .A(p_input[3766]), .B(n34070), .Z(n34073) );
  XNOR U33727 ( .A(n34070), .B(n33712), .Z(n34072) );
  IV U33728 ( .A(p_input[3734]), .Z(n33712) );
  XOR U33729 ( .A(n34074), .B(n34075), .Z(n34070) );
  AND U33730 ( .A(n34076), .B(n34077), .Z(n34075) );
  XNOR U33731 ( .A(p_input[3765]), .B(n34074), .Z(n34077) );
  XNOR U33732 ( .A(n34074), .B(n33721), .Z(n34076) );
  IV U33733 ( .A(p_input[3733]), .Z(n33721) );
  XOR U33734 ( .A(n34078), .B(n34079), .Z(n34074) );
  AND U33735 ( .A(n34080), .B(n34081), .Z(n34079) );
  XNOR U33736 ( .A(p_input[3764]), .B(n34078), .Z(n34081) );
  XNOR U33737 ( .A(n34078), .B(n33730), .Z(n34080) );
  IV U33738 ( .A(p_input[3732]), .Z(n33730) );
  XOR U33739 ( .A(n34082), .B(n34083), .Z(n34078) );
  AND U33740 ( .A(n34084), .B(n34085), .Z(n34083) );
  XNOR U33741 ( .A(p_input[3763]), .B(n34082), .Z(n34085) );
  XNOR U33742 ( .A(n34082), .B(n33739), .Z(n34084) );
  IV U33743 ( .A(p_input[3731]), .Z(n33739) );
  XOR U33744 ( .A(n34086), .B(n34087), .Z(n34082) );
  AND U33745 ( .A(n34088), .B(n34089), .Z(n34087) );
  XNOR U33746 ( .A(p_input[3762]), .B(n34086), .Z(n34089) );
  XNOR U33747 ( .A(n34086), .B(n33748), .Z(n34088) );
  IV U33748 ( .A(p_input[3730]), .Z(n33748) );
  XOR U33749 ( .A(n34090), .B(n34091), .Z(n34086) );
  AND U33750 ( .A(n34092), .B(n34093), .Z(n34091) );
  XNOR U33751 ( .A(p_input[3761]), .B(n34090), .Z(n34093) );
  XNOR U33752 ( .A(n34090), .B(n33757), .Z(n34092) );
  IV U33753 ( .A(p_input[3729]), .Z(n33757) );
  XOR U33754 ( .A(n34094), .B(n34095), .Z(n34090) );
  AND U33755 ( .A(n34096), .B(n34097), .Z(n34095) );
  XNOR U33756 ( .A(p_input[3760]), .B(n34094), .Z(n34097) );
  XNOR U33757 ( .A(n34094), .B(n33766), .Z(n34096) );
  IV U33758 ( .A(p_input[3728]), .Z(n33766) );
  XOR U33759 ( .A(n34098), .B(n34099), .Z(n34094) );
  AND U33760 ( .A(n34100), .B(n34101), .Z(n34099) );
  XNOR U33761 ( .A(p_input[3759]), .B(n34098), .Z(n34101) );
  XNOR U33762 ( .A(n34098), .B(n33775), .Z(n34100) );
  IV U33763 ( .A(p_input[3727]), .Z(n33775) );
  XOR U33764 ( .A(n34102), .B(n34103), .Z(n34098) );
  AND U33765 ( .A(n34104), .B(n34105), .Z(n34103) );
  XNOR U33766 ( .A(p_input[3758]), .B(n34102), .Z(n34105) );
  XNOR U33767 ( .A(n34102), .B(n33784), .Z(n34104) );
  IV U33768 ( .A(p_input[3726]), .Z(n33784) );
  XOR U33769 ( .A(n34106), .B(n34107), .Z(n34102) );
  AND U33770 ( .A(n34108), .B(n34109), .Z(n34107) );
  XNOR U33771 ( .A(p_input[3757]), .B(n34106), .Z(n34109) );
  XNOR U33772 ( .A(n34106), .B(n33793), .Z(n34108) );
  IV U33773 ( .A(p_input[3725]), .Z(n33793) );
  XOR U33774 ( .A(n34110), .B(n34111), .Z(n34106) );
  AND U33775 ( .A(n34112), .B(n34113), .Z(n34111) );
  XNOR U33776 ( .A(p_input[3756]), .B(n34110), .Z(n34113) );
  XNOR U33777 ( .A(n34110), .B(n33802), .Z(n34112) );
  IV U33778 ( .A(p_input[3724]), .Z(n33802) );
  XOR U33779 ( .A(n34114), .B(n34115), .Z(n34110) );
  AND U33780 ( .A(n34116), .B(n34117), .Z(n34115) );
  XNOR U33781 ( .A(p_input[3755]), .B(n34114), .Z(n34117) );
  XNOR U33782 ( .A(n34114), .B(n33811), .Z(n34116) );
  IV U33783 ( .A(p_input[3723]), .Z(n33811) );
  XOR U33784 ( .A(n34118), .B(n34119), .Z(n34114) );
  AND U33785 ( .A(n34120), .B(n34121), .Z(n34119) );
  XNOR U33786 ( .A(p_input[3754]), .B(n34118), .Z(n34121) );
  XNOR U33787 ( .A(n34118), .B(n33820), .Z(n34120) );
  IV U33788 ( .A(p_input[3722]), .Z(n33820) );
  XOR U33789 ( .A(n34122), .B(n34123), .Z(n34118) );
  AND U33790 ( .A(n34124), .B(n34125), .Z(n34123) );
  XNOR U33791 ( .A(p_input[3753]), .B(n34122), .Z(n34125) );
  XNOR U33792 ( .A(n34122), .B(n33829), .Z(n34124) );
  IV U33793 ( .A(p_input[3721]), .Z(n33829) );
  XOR U33794 ( .A(n34126), .B(n34127), .Z(n34122) );
  AND U33795 ( .A(n34128), .B(n34129), .Z(n34127) );
  XNOR U33796 ( .A(p_input[3752]), .B(n34126), .Z(n34129) );
  XNOR U33797 ( .A(n34126), .B(n33838), .Z(n34128) );
  IV U33798 ( .A(p_input[3720]), .Z(n33838) );
  XOR U33799 ( .A(n34130), .B(n34131), .Z(n34126) );
  AND U33800 ( .A(n34132), .B(n34133), .Z(n34131) );
  XNOR U33801 ( .A(p_input[3751]), .B(n34130), .Z(n34133) );
  XNOR U33802 ( .A(n34130), .B(n33847), .Z(n34132) );
  IV U33803 ( .A(p_input[3719]), .Z(n33847) );
  XOR U33804 ( .A(n34134), .B(n34135), .Z(n34130) );
  AND U33805 ( .A(n34136), .B(n34137), .Z(n34135) );
  XNOR U33806 ( .A(p_input[3750]), .B(n34134), .Z(n34137) );
  XNOR U33807 ( .A(n34134), .B(n33856), .Z(n34136) );
  IV U33808 ( .A(p_input[3718]), .Z(n33856) );
  XOR U33809 ( .A(n34138), .B(n34139), .Z(n34134) );
  AND U33810 ( .A(n34140), .B(n34141), .Z(n34139) );
  XNOR U33811 ( .A(p_input[3749]), .B(n34138), .Z(n34141) );
  XNOR U33812 ( .A(n34138), .B(n33865), .Z(n34140) );
  IV U33813 ( .A(p_input[3717]), .Z(n33865) );
  XOR U33814 ( .A(n34142), .B(n34143), .Z(n34138) );
  AND U33815 ( .A(n34144), .B(n34145), .Z(n34143) );
  XNOR U33816 ( .A(p_input[3748]), .B(n34142), .Z(n34145) );
  XNOR U33817 ( .A(n34142), .B(n33874), .Z(n34144) );
  IV U33818 ( .A(p_input[3716]), .Z(n33874) );
  XOR U33819 ( .A(n34146), .B(n34147), .Z(n34142) );
  AND U33820 ( .A(n34148), .B(n34149), .Z(n34147) );
  XNOR U33821 ( .A(p_input[3747]), .B(n34146), .Z(n34149) );
  XNOR U33822 ( .A(n34146), .B(n33883), .Z(n34148) );
  IV U33823 ( .A(p_input[3715]), .Z(n33883) );
  XOR U33824 ( .A(n34150), .B(n34151), .Z(n34146) );
  AND U33825 ( .A(n34152), .B(n34153), .Z(n34151) );
  XNOR U33826 ( .A(p_input[3746]), .B(n34150), .Z(n34153) );
  XNOR U33827 ( .A(n34150), .B(n33892), .Z(n34152) );
  IV U33828 ( .A(p_input[3714]), .Z(n33892) );
  XNOR U33829 ( .A(n34154), .B(n34155), .Z(n34150) );
  AND U33830 ( .A(n34156), .B(n34157), .Z(n34155) );
  XOR U33831 ( .A(p_input[3745]), .B(n34154), .Z(n34157) );
  XNOR U33832 ( .A(p_input[3713]), .B(n34154), .Z(n34156) );
  AND U33833 ( .A(p_input[3744]), .B(n34158), .Z(n34154) );
  IV U33834 ( .A(p_input[3712]), .Z(n34158) );
  XOR U33835 ( .A(n34159), .B(n34160), .Z(n33248) );
  AND U33836 ( .A(n564), .B(n34161), .Z(n34160) );
  XNOR U33837 ( .A(n34162), .B(n34159), .Z(n34161) );
  XOR U33838 ( .A(n34163), .B(n34164), .Z(n564) );
  AND U33839 ( .A(n34165), .B(n34166), .Z(n34164) );
  XNOR U33840 ( .A(n33263), .B(n34163), .Z(n34166) );
  AND U33841 ( .A(p_input[3711]), .B(p_input[3679]), .Z(n33263) );
  XNOR U33842 ( .A(n34163), .B(n33260), .Z(n34165) );
  IV U33843 ( .A(n34167), .Z(n33260) );
  AND U33844 ( .A(p_input[3615]), .B(p_input[3647]), .Z(n34167) );
  XOR U33845 ( .A(n34168), .B(n34169), .Z(n34163) );
  AND U33846 ( .A(n34170), .B(n34171), .Z(n34169) );
  XOR U33847 ( .A(n34168), .B(n33275), .Z(n34171) );
  XNOR U33848 ( .A(p_input[3678]), .B(n34172), .Z(n33275) );
  AND U33849 ( .A(n707), .B(n34173), .Z(n34172) );
  XOR U33850 ( .A(p_input[3710]), .B(p_input[3678]), .Z(n34173) );
  XNOR U33851 ( .A(n33272), .B(n34168), .Z(n34170) );
  XOR U33852 ( .A(n34174), .B(n34175), .Z(n33272) );
  AND U33853 ( .A(n704), .B(n34176), .Z(n34175) );
  XOR U33854 ( .A(p_input[3646]), .B(p_input[3614]), .Z(n34176) );
  XOR U33855 ( .A(n34177), .B(n34178), .Z(n34168) );
  AND U33856 ( .A(n34179), .B(n34180), .Z(n34178) );
  XOR U33857 ( .A(n34177), .B(n33287), .Z(n34180) );
  XNOR U33858 ( .A(p_input[3677]), .B(n34181), .Z(n33287) );
  AND U33859 ( .A(n707), .B(n34182), .Z(n34181) );
  XOR U33860 ( .A(p_input[3709]), .B(p_input[3677]), .Z(n34182) );
  XNOR U33861 ( .A(n33284), .B(n34177), .Z(n34179) );
  XOR U33862 ( .A(n34183), .B(n34184), .Z(n33284) );
  AND U33863 ( .A(n704), .B(n34185), .Z(n34184) );
  XOR U33864 ( .A(p_input[3645]), .B(p_input[3613]), .Z(n34185) );
  XOR U33865 ( .A(n34186), .B(n34187), .Z(n34177) );
  AND U33866 ( .A(n34188), .B(n34189), .Z(n34187) );
  XOR U33867 ( .A(n34186), .B(n33299), .Z(n34189) );
  XNOR U33868 ( .A(p_input[3676]), .B(n34190), .Z(n33299) );
  AND U33869 ( .A(n707), .B(n34191), .Z(n34190) );
  XOR U33870 ( .A(p_input[3708]), .B(p_input[3676]), .Z(n34191) );
  XNOR U33871 ( .A(n33296), .B(n34186), .Z(n34188) );
  XOR U33872 ( .A(n34192), .B(n34193), .Z(n33296) );
  AND U33873 ( .A(n704), .B(n34194), .Z(n34193) );
  XOR U33874 ( .A(p_input[3644]), .B(p_input[3612]), .Z(n34194) );
  XOR U33875 ( .A(n34195), .B(n34196), .Z(n34186) );
  AND U33876 ( .A(n34197), .B(n34198), .Z(n34196) );
  XOR U33877 ( .A(n34195), .B(n33311), .Z(n34198) );
  XNOR U33878 ( .A(p_input[3675]), .B(n34199), .Z(n33311) );
  AND U33879 ( .A(n707), .B(n34200), .Z(n34199) );
  XOR U33880 ( .A(p_input[3707]), .B(p_input[3675]), .Z(n34200) );
  XNOR U33881 ( .A(n33308), .B(n34195), .Z(n34197) );
  XOR U33882 ( .A(n34201), .B(n34202), .Z(n33308) );
  AND U33883 ( .A(n704), .B(n34203), .Z(n34202) );
  XOR U33884 ( .A(p_input[3643]), .B(p_input[3611]), .Z(n34203) );
  XOR U33885 ( .A(n34204), .B(n34205), .Z(n34195) );
  AND U33886 ( .A(n34206), .B(n34207), .Z(n34205) );
  XOR U33887 ( .A(n34204), .B(n33323), .Z(n34207) );
  XNOR U33888 ( .A(p_input[3674]), .B(n34208), .Z(n33323) );
  AND U33889 ( .A(n707), .B(n34209), .Z(n34208) );
  XOR U33890 ( .A(p_input[3706]), .B(p_input[3674]), .Z(n34209) );
  XNOR U33891 ( .A(n33320), .B(n34204), .Z(n34206) );
  XOR U33892 ( .A(n34210), .B(n34211), .Z(n33320) );
  AND U33893 ( .A(n704), .B(n34212), .Z(n34211) );
  XOR U33894 ( .A(p_input[3642]), .B(p_input[3610]), .Z(n34212) );
  XOR U33895 ( .A(n34213), .B(n34214), .Z(n34204) );
  AND U33896 ( .A(n34215), .B(n34216), .Z(n34214) );
  XOR U33897 ( .A(n34213), .B(n33335), .Z(n34216) );
  XNOR U33898 ( .A(p_input[3673]), .B(n34217), .Z(n33335) );
  AND U33899 ( .A(n707), .B(n34218), .Z(n34217) );
  XOR U33900 ( .A(p_input[3705]), .B(p_input[3673]), .Z(n34218) );
  XNOR U33901 ( .A(n33332), .B(n34213), .Z(n34215) );
  XOR U33902 ( .A(n34219), .B(n34220), .Z(n33332) );
  AND U33903 ( .A(n704), .B(n34221), .Z(n34220) );
  XOR U33904 ( .A(p_input[3641]), .B(p_input[3609]), .Z(n34221) );
  XOR U33905 ( .A(n34222), .B(n34223), .Z(n34213) );
  AND U33906 ( .A(n34224), .B(n34225), .Z(n34223) );
  XOR U33907 ( .A(n34222), .B(n33347), .Z(n34225) );
  XNOR U33908 ( .A(p_input[3672]), .B(n34226), .Z(n33347) );
  AND U33909 ( .A(n707), .B(n34227), .Z(n34226) );
  XOR U33910 ( .A(p_input[3704]), .B(p_input[3672]), .Z(n34227) );
  XNOR U33911 ( .A(n33344), .B(n34222), .Z(n34224) );
  XOR U33912 ( .A(n34228), .B(n34229), .Z(n33344) );
  AND U33913 ( .A(n704), .B(n34230), .Z(n34229) );
  XOR U33914 ( .A(p_input[3640]), .B(p_input[3608]), .Z(n34230) );
  XOR U33915 ( .A(n34231), .B(n34232), .Z(n34222) );
  AND U33916 ( .A(n34233), .B(n34234), .Z(n34232) );
  XOR U33917 ( .A(n34231), .B(n33359), .Z(n34234) );
  XNOR U33918 ( .A(p_input[3671]), .B(n34235), .Z(n33359) );
  AND U33919 ( .A(n707), .B(n34236), .Z(n34235) );
  XOR U33920 ( .A(p_input[3703]), .B(p_input[3671]), .Z(n34236) );
  XNOR U33921 ( .A(n33356), .B(n34231), .Z(n34233) );
  XOR U33922 ( .A(n34237), .B(n34238), .Z(n33356) );
  AND U33923 ( .A(n704), .B(n34239), .Z(n34238) );
  XOR U33924 ( .A(p_input[3639]), .B(p_input[3607]), .Z(n34239) );
  XOR U33925 ( .A(n34240), .B(n34241), .Z(n34231) );
  AND U33926 ( .A(n34242), .B(n34243), .Z(n34241) );
  XOR U33927 ( .A(n34240), .B(n33371), .Z(n34243) );
  XNOR U33928 ( .A(p_input[3670]), .B(n34244), .Z(n33371) );
  AND U33929 ( .A(n707), .B(n34245), .Z(n34244) );
  XOR U33930 ( .A(p_input[3702]), .B(p_input[3670]), .Z(n34245) );
  XNOR U33931 ( .A(n33368), .B(n34240), .Z(n34242) );
  XOR U33932 ( .A(n34246), .B(n34247), .Z(n33368) );
  AND U33933 ( .A(n704), .B(n34248), .Z(n34247) );
  XOR U33934 ( .A(p_input[3638]), .B(p_input[3606]), .Z(n34248) );
  XOR U33935 ( .A(n34249), .B(n34250), .Z(n34240) );
  AND U33936 ( .A(n34251), .B(n34252), .Z(n34250) );
  XOR U33937 ( .A(n34249), .B(n33383), .Z(n34252) );
  XNOR U33938 ( .A(p_input[3669]), .B(n34253), .Z(n33383) );
  AND U33939 ( .A(n707), .B(n34254), .Z(n34253) );
  XOR U33940 ( .A(p_input[3701]), .B(p_input[3669]), .Z(n34254) );
  XNOR U33941 ( .A(n33380), .B(n34249), .Z(n34251) );
  XOR U33942 ( .A(n34255), .B(n34256), .Z(n33380) );
  AND U33943 ( .A(n704), .B(n34257), .Z(n34256) );
  XOR U33944 ( .A(p_input[3637]), .B(p_input[3605]), .Z(n34257) );
  XOR U33945 ( .A(n34258), .B(n34259), .Z(n34249) );
  AND U33946 ( .A(n34260), .B(n34261), .Z(n34259) );
  XOR U33947 ( .A(n34258), .B(n33395), .Z(n34261) );
  XNOR U33948 ( .A(p_input[3668]), .B(n34262), .Z(n33395) );
  AND U33949 ( .A(n707), .B(n34263), .Z(n34262) );
  XOR U33950 ( .A(p_input[3700]), .B(p_input[3668]), .Z(n34263) );
  XNOR U33951 ( .A(n33392), .B(n34258), .Z(n34260) );
  XOR U33952 ( .A(n34264), .B(n34265), .Z(n33392) );
  AND U33953 ( .A(n704), .B(n34266), .Z(n34265) );
  XOR U33954 ( .A(p_input[3636]), .B(p_input[3604]), .Z(n34266) );
  XOR U33955 ( .A(n34267), .B(n34268), .Z(n34258) );
  AND U33956 ( .A(n34269), .B(n34270), .Z(n34268) );
  XOR U33957 ( .A(n34267), .B(n33407), .Z(n34270) );
  XNOR U33958 ( .A(p_input[3667]), .B(n34271), .Z(n33407) );
  AND U33959 ( .A(n707), .B(n34272), .Z(n34271) );
  XOR U33960 ( .A(p_input[3699]), .B(p_input[3667]), .Z(n34272) );
  XNOR U33961 ( .A(n33404), .B(n34267), .Z(n34269) );
  XOR U33962 ( .A(n34273), .B(n34274), .Z(n33404) );
  AND U33963 ( .A(n704), .B(n34275), .Z(n34274) );
  XOR U33964 ( .A(p_input[3635]), .B(p_input[3603]), .Z(n34275) );
  XOR U33965 ( .A(n34276), .B(n34277), .Z(n34267) );
  AND U33966 ( .A(n34278), .B(n34279), .Z(n34277) );
  XOR U33967 ( .A(n34276), .B(n33419), .Z(n34279) );
  XNOR U33968 ( .A(p_input[3666]), .B(n34280), .Z(n33419) );
  AND U33969 ( .A(n707), .B(n34281), .Z(n34280) );
  XOR U33970 ( .A(p_input[3698]), .B(p_input[3666]), .Z(n34281) );
  XNOR U33971 ( .A(n33416), .B(n34276), .Z(n34278) );
  XOR U33972 ( .A(n34282), .B(n34283), .Z(n33416) );
  AND U33973 ( .A(n704), .B(n34284), .Z(n34283) );
  XOR U33974 ( .A(p_input[3634]), .B(p_input[3602]), .Z(n34284) );
  XOR U33975 ( .A(n34285), .B(n34286), .Z(n34276) );
  AND U33976 ( .A(n34287), .B(n34288), .Z(n34286) );
  XOR U33977 ( .A(n34285), .B(n33431), .Z(n34288) );
  XNOR U33978 ( .A(p_input[3665]), .B(n34289), .Z(n33431) );
  AND U33979 ( .A(n707), .B(n34290), .Z(n34289) );
  XOR U33980 ( .A(p_input[3697]), .B(p_input[3665]), .Z(n34290) );
  XNOR U33981 ( .A(n33428), .B(n34285), .Z(n34287) );
  XOR U33982 ( .A(n34291), .B(n34292), .Z(n33428) );
  AND U33983 ( .A(n704), .B(n34293), .Z(n34292) );
  XOR U33984 ( .A(p_input[3633]), .B(p_input[3601]), .Z(n34293) );
  XOR U33985 ( .A(n34294), .B(n34295), .Z(n34285) );
  AND U33986 ( .A(n34296), .B(n34297), .Z(n34295) );
  XOR U33987 ( .A(n34294), .B(n33443), .Z(n34297) );
  XNOR U33988 ( .A(p_input[3664]), .B(n34298), .Z(n33443) );
  AND U33989 ( .A(n707), .B(n34299), .Z(n34298) );
  XOR U33990 ( .A(p_input[3696]), .B(p_input[3664]), .Z(n34299) );
  XNOR U33991 ( .A(n33440), .B(n34294), .Z(n34296) );
  XOR U33992 ( .A(n34300), .B(n34301), .Z(n33440) );
  AND U33993 ( .A(n704), .B(n34302), .Z(n34301) );
  XOR U33994 ( .A(p_input[3632]), .B(p_input[3600]), .Z(n34302) );
  XOR U33995 ( .A(n34303), .B(n34304), .Z(n34294) );
  AND U33996 ( .A(n34305), .B(n34306), .Z(n34304) );
  XOR U33997 ( .A(n34303), .B(n33455), .Z(n34306) );
  XNOR U33998 ( .A(p_input[3663]), .B(n34307), .Z(n33455) );
  AND U33999 ( .A(n707), .B(n34308), .Z(n34307) );
  XOR U34000 ( .A(p_input[3695]), .B(p_input[3663]), .Z(n34308) );
  XNOR U34001 ( .A(n33452), .B(n34303), .Z(n34305) );
  XOR U34002 ( .A(n34309), .B(n34310), .Z(n33452) );
  AND U34003 ( .A(n704), .B(n34311), .Z(n34310) );
  XOR U34004 ( .A(p_input[3631]), .B(p_input[3599]), .Z(n34311) );
  XOR U34005 ( .A(n34312), .B(n34313), .Z(n34303) );
  AND U34006 ( .A(n34314), .B(n34315), .Z(n34313) );
  XOR U34007 ( .A(n34312), .B(n33467), .Z(n34315) );
  XNOR U34008 ( .A(p_input[3662]), .B(n34316), .Z(n33467) );
  AND U34009 ( .A(n707), .B(n34317), .Z(n34316) );
  XOR U34010 ( .A(p_input[3694]), .B(p_input[3662]), .Z(n34317) );
  XNOR U34011 ( .A(n33464), .B(n34312), .Z(n34314) );
  XOR U34012 ( .A(n34318), .B(n34319), .Z(n33464) );
  AND U34013 ( .A(n704), .B(n34320), .Z(n34319) );
  XOR U34014 ( .A(p_input[3630]), .B(p_input[3598]), .Z(n34320) );
  XOR U34015 ( .A(n34321), .B(n34322), .Z(n34312) );
  AND U34016 ( .A(n34323), .B(n34324), .Z(n34322) );
  XOR U34017 ( .A(n34321), .B(n33479), .Z(n34324) );
  XNOR U34018 ( .A(p_input[3661]), .B(n34325), .Z(n33479) );
  AND U34019 ( .A(n707), .B(n34326), .Z(n34325) );
  XOR U34020 ( .A(p_input[3693]), .B(p_input[3661]), .Z(n34326) );
  XNOR U34021 ( .A(n33476), .B(n34321), .Z(n34323) );
  XOR U34022 ( .A(n34327), .B(n34328), .Z(n33476) );
  AND U34023 ( .A(n704), .B(n34329), .Z(n34328) );
  XOR U34024 ( .A(p_input[3629]), .B(p_input[3597]), .Z(n34329) );
  XOR U34025 ( .A(n34330), .B(n34331), .Z(n34321) );
  AND U34026 ( .A(n34332), .B(n34333), .Z(n34331) );
  XOR U34027 ( .A(n34330), .B(n33491), .Z(n34333) );
  XNOR U34028 ( .A(p_input[3660]), .B(n34334), .Z(n33491) );
  AND U34029 ( .A(n707), .B(n34335), .Z(n34334) );
  XOR U34030 ( .A(p_input[3692]), .B(p_input[3660]), .Z(n34335) );
  XNOR U34031 ( .A(n33488), .B(n34330), .Z(n34332) );
  XOR U34032 ( .A(n34336), .B(n34337), .Z(n33488) );
  AND U34033 ( .A(n704), .B(n34338), .Z(n34337) );
  XOR U34034 ( .A(p_input[3628]), .B(p_input[3596]), .Z(n34338) );
  XOR U34035 ( .A(n34339), .B(n34340), .Z(n34330) );
  AND U34036 ( .A(n34341), .B(n34342), .Z(n34340) );
  XOR U34037 ( .A(n34339), .B(n33503), .Z(n34342) );
  XNOR U34038 ( .A(p_input[3659]), .B(n34343), .Z(n33503) );
  AND U34039 ( .A(n707), .B(n34344), .Z(n34343) );
  XOR U34040 ( .A(p_input[3691]), .B(p_input[3659]), .Z(n34344) );
  XNOR U34041 ( .A(n33500), .B(n34339), .Z(n34341) );
  XOR U34042 ( .A(n34345), .B(n34346), .Z(n33500) );
  AND U34043 ( .A(n704), .B(n34347), .Z(n34346) );
  XOR U34044 ( .A(p_input[3627]), .B(p_input[3595]), .Z(n34347) );
  XOR U34045 ( .A(n34348), .B(n34349), .Z(n34339) );
  AND U34046 ( .A(n34350), .B(n34351), .Z(n34349) );
  XOR U34047 ( .A(n34348), .B(n33515), .Z(n34351) );
  XNOR U34048 ( .A(p_input[3658]), .B(n34352), .Z(n33515) );
  AND U34049 ( .A(n707), .B(n34353), .Z(n34352) );
  XOR U34050 ( .A(p_input[3690]), .B(p_input[3658]), .Z(n34353) );
  XNOR U34051 ( .A(n33512), .B(n34348), .Z(n34350) );
  XOR U34052 ( .A(n34354), .B(n34355), .Z(n33512) );
  AND U34053 ( .A(n704), .B(n34356), .Z(n34355) );
  XOR U34054 ( .A(p_input[3626]), .B(p_input[3594]), .Z(n34356) );
  XOR U34055 ( .A(n34357), .B(n34358), .Z(n34348) );
  AND U34056 ( .A(n34359), .B(n34360), .Z(n34358) );
  XOR U34057 ( .A(n34357), .B(n33527), .Z(n34360) );
  XNOR U34058 ( .A(p_input[3657]), .B(n34361), .Z(n33527) );
  AND U34059 ( .A(n707), .B(n34362), .Z(n34361) );
  XOR U34060 ( .A(p_input[3689]), .B(p_input[3657]), .Z(n34362) );
  XNOR U34061 ( .A(n33524), .B(n34357), .Z(n34359) );
  XOR U34062 ( .A(n34363), .B(n34364), .Z(n33524) );
  AND U34063 ( .A(n704), .B(n34365), .Z(n34364) );
  XOR U34064 ( .A(p_input[3625]), .B(p_input[3593]), .Z(n34365) );
  XOR U34065 ( .A(n34366), .B(n34367), .Z(n34357) );
  AND U34066 ( .A(n34368), .B(n34369), .Z(n34367) );
  XOR U34067 ( .A(n34366), .B(n33539), .Z(n34369) );
  XNOR U34068 ( .A(p_input[3656]), .B(n34370), .Z(n33539) );
  AND U34069 ( .A(n707), .B(n34371), .Z(n34370) );
  XOR U34070 ( .A(p_input[3688]), .B(p_input[3656]), .Z(n34371) );
  XNOR U34071 ( .A(n33536), .B(n34366), .Z(n34368) );
  XOR U34072 ( .A(n34372), .B(n34373), .Z(n33536) );
  AND U34073 ( .A(n704), .B(n34374), .Z(n34373) );
  XOR U34074 ( .A(p_input[3624]), .B(p_input[3592]), .Z(n34374) );
  XOR U34075 ( .A(n34375), .B(n34376), .Z(n34366) );
  AND U34076 ( .A(n34377), .B(n34378), .Z(n34376) );
  XOR U34077 ( .A(n34375), .B(n33551), .Z(n34378) );
  XNOR U34078 ( .A(p_input[3655]), .B(n34379), .Z(n33551) );
  AND U34079 ( .A(n707), .B(n34380), .Z(n34379) );
  XOR U34080 ( .A(p_input[3687]), .B(p_input[3655]), .Z(n34380) );
  XNOR U34081 ( .A(n33548), .B(n34375), .Z(n34377) );
  XOR U34082 ( .A(n34381), .B(n34382), .Z(n33548) );
  AND U34083 ( .A(n704), .B(n34383), .Z(n34382) );
  XOR U34084 ( .A(p_input[3623]), .B(p_input[3591]), .Z(n34383) );
  XOR U34085 ( .A(n34384), .B(n34385), .Z(n34375) );
  AND U34086 ( .A(n34386), .B(n34387), .Z(n34385) );
  XOR U34087 ( .A(n34384), .B(n33563), .Z(n34387) );
  XNOR U34088 ( .A(p_input[3654]), .B(n34388), .Z(n33563) );
  AND U34089 ( .A(n707), .B(n34389), .Z(n34388) );
  XOR U34090 ( .A(p_input[3686]), .B(p_input[3654]), .Z(n34389) );
  XNOR U34091 ( .A(n33560), .B(n34384), .Z(n34386) );
  XOR U34092 ( .A(n34390), .B(n34391), .Z(n33560) );
  AND U34093 ( .A(n704), .B(n34392), .Z(n34391) );
  XOR U34094 ( .A(p_input[3622]), .B(p_input[3590]), .Z(n34392) );
  XOR U34095 ( .A(n34393), .B(n34394), .Z(n34384) );
  AND U34096 ( .A(n34395), .B(n34396), .Z(n34394) );
  XOR U34097 ( .A(n34393), .B(n33575), .Z(n34396) );
  XNOR U34098 ( .A(p_input[3653]), .B(n34397), .Z(n33575) );
  AND U34099 ( .A(n707), .B(n34398), .Z(n34397) );
  XOR U34100 ( .A(p_input[3685]), .B(p_input[3653]), .Z(n34398) );
  XNOR U34101 ( .A(n33572), .B(n34393), .Z(n34395) );
  XOR U34102 ( .A(n34399), .B(n34400), .Z(n33572) );
  AND U34103 ( .A(n704), .B(n34401), .Z(n34400) );
  XOR U34104 ( .A(p_input[3621]), .B(p_input[3589]), .Z(n34401) );
  XOR U34105 ( .A(n34402), .B(n34403), .Z(n34393) );
  AND U34106 ( .A(n34404), .B(n34405), .Z(n34403) );
  XOR U34107 ( .A(n34402), .B(n33587), .Z(n34405) );
  XNOR U34108 ( .A(p_input[3652]), .B(n34406), .Z(n33587) );
  AND U34109 ( .A(n707), .B(n34407), .Z(n34406) );
  XOR U34110 ( .A(p_input[3684]), .B(p_input[3652]), .Z(n34407) );
  XNOR U34111 ( .A(n33584), .B(n34402), .Z(n34404) );
  XOR U34112 ( .A(n34408), .B(n34409), .Z(n33584) );
  AND U34113 ( .A(n704), .B(n34410), .Z(n34409) );
  XOR U34114 ( .A(p_input[3620]), .B(p_input[3588]), .Z(n34410) );
  XOR U34115 ( .A(n34411), .B(n34412), .Z(n34402) );
  AND U34116 ( .A(n34413), .B(n34414), .Z(n34412) );
  XOR U34117 ( .A(n34411), .B(n33599), .Z(n34414) );
  XNOR U34118 ( .A(p_input[3651]), .B(n34415), .Z(n33599) );
  AND U34119 ( .A(n707), .B(n34416), .Z(n34415) );
  XOR U34120 ( .A(p_input[3683]), .B(p_input[3651]), .Z(n34416) );
  XNOR U34121 ( .A(n33596), .B(n34411), .Z(n34413) );
  XOR U34122 ( .A(n34417), .B(n34418), .Z(n33596) );
  AND U34123 ( .A(n704), .B(n34419), .Z(n34418) );
  XOR U34124 ( .A(p_input[3619]), .B(p_input[3587]), .Z(n34419) );
  XOR U34125 ( .A(n34420), .B(n34421), .Z(n34411) );
  AND U34126 ( .A(n34422), .B(n34423), .Z(n34421) );
  XOR U34127 ( .A(n34420), .B(n33611), .Z(n34423) );
  XNOR U34128 ( .A(p_input[3650]), .B(n34424), .Z(n33611) );
  AND U34129 ( .A(n707), .B(n34425), .Z(n34424) );
  XOR U34130 ( .A(p_input[3682]), .B(p_input[3650]), .Z(n34425) );
  XNOR U34131 ( .A(n33608), .B(n34420), .Z(n34422) );
  XOR U34132 ( .A(n34426), .B(n34427), .Z(n33608) );
  AND U34133 ( .A(n704), .B(n34428), .Z(n34427) );
  XOR U34134 ( .A(p_input[3618]), .B(p_input[3586]), .Z(n34428) );
  XOR U34135 ( .A(n34429), .B(n34430), .Z(n34420) );
  AND U34136 ( .A(n34431), .B(n34432), .Z(n34430) );
  XNOR U34137 ( .A(n34433), .B(n33624), .Z(n34432) );
  XNOR U34138 ( .A(p_input[3649]), .B(n34434), .Z(n33624) );
  AND U34139 ( .A(n707), .B(n34435), .Z(n34434) );
  XNOR U34140 ( .A(p_input[3681]), .B(n34436), .Z(n34435) );
  IV U34141 ( .A(p_input[3649]), .Z(n34436) );
  XNOR U34142 ( .A(n33621), .B(n34429), .Z(n34431) );
  XNOR U34143 ( .A(p_input[3585]), .B(n34437), .Z(n33621) );
  AND U34144 ( .A(n704), .B(n34438), .Z(n34437) );
  XOR U34145 ( .A(p_input[3617]), .B(p_input[3585]), .Z(n34438) );
  IV U34146 ( .A(n34433), .Z(n34429) );
  AND U34147 ( .A(n34159), .B(n34162), .Z(n34433) );
  XOR U34148 ( .A(p_input[3648]), .B(n34439), .Z(n34162) );
  AND U34149 ( .A(n707), .B(n34440), .Z(n34439) );
  XOR U34150 ( .A(p_input[3680]), .B(p_input[3648]), .Z(n34440) );
  XOR U34151 ( .A(n34441), .B(n34442), .Z(n707) );
  AND U34152 ( .A(n34443), .B(n34444), .Z(n34442) );
  XNOR U34153 ( .A(p_input[3711]), .B(n34441), .Z(n34444) );
  XOR U34154 ( .A(n34441), .B(p_input[3679]), .Z(n34443) );
  XOR U34155 ( .A(n34445), .B(n34446), .Z(n34441) );
  AND U34156 ( .A(n34447), .B(n34448), .Z(n34446) );
  XNOR U34157 ( .A(p_input[3710]), .B(n34445), .Z(n34448) );
  XOR U34158 ( .A(n34445), .B(p_input[3678]), .Z(n34447) );
  XOR U34159 ( .A(n34449), .B(n34450), .Z(n34445) );
  AND U34160 ( .A(n34451), .B(n34452), .Z(n34450) );
  XNOR U34161 ( .A(p_input[3709]), .B(n34449), .Z(n34452) );
  XOR U34162 ( .A(n34449), .B(p_input[3677]), .Z(n34451) );
  XOR U34163 ( .A(n34453), .B(n34454), .Z(n34449) );
  AND U34164 ( .A(n34455), .B(n34456), .Z(n34454) );
  XNOR U34165 ( .A(p_input[3708]), .B(n34453), .Z(n34456) );
  XOR U34166 ( .A(n34453), .B(p_input[3676]), .Z(n34455) );
  XOR U34167 ( .A(n34457), .B(n34458), .Z(n34453) );
  AND U34168 ( .A(n34459), .B(n34460), .Z(n34458) );
  XNOR U34169 ( .A(p_input[3707]), .B(n34457), .Z(n34460) );
  XOR U34170 ( .A(n34457), .B(p_input[3675]), .Z(n34459) );
  XOR U34171 ( .A(n34461), .B(n34462), .Z(n34457) );
  AND U34172 ( .A(n34463), .B(n34464), .Z(n34462) );
  XNOR U34173 ( .A(p_input[3706]), .B(n34461), .Z(n34464) );
  XOR U34174 ( .A(n34461), .B(p_input[3674]), .Z(n34463) );
  XOR U34175 ( .A(n34465), .B(n34466), .Z(n34461) );
  AND U34176 ( .A(n34467), .B(n34468), .Z(n34466) );
  XNOR U34177 ( .A(p_input[3705]), .B(n34465), .Z(n34468) );
  XOR U34178 ( .A(n34465), .B(p_input[3673]), .Z(n34467) );
  XOR U34179 ( .A(n34469), .B(n34470), .Z(n34465) );
  AND U34180 ( .A(n34471), .B(n34472), .Z(n34470) );
  XNOR U34181 ( .A(p_input[3704]), .B(n34469), .Z(n34472) );
  XOR U34182 ( .A(n34469), .B(p_input[3672]), .Z(n34471) );
  XOR U34183 ( .A(n34473), .B(n34474), .Z(n34469) );
  AND U34184 ( .A(n34475), .B(n34476), .Z(n34474) );
  XNOR U34185 ( .A(p_input[3703]), .B(n34473), .Z(n34476) );
  XOR U34186 ( .A(n34473), .B(p_input[3671]), .Z(n34475) );
  XOR U34187 ( .A(n34477), .B(n34478), .Z(n34473) );
  AND U34188 ( .A(n34479), .B(n34480), .Z(n34478) );
  XNOR U34189 ( .A(p_input[3702]), .B(n34477), .Z(n34480) );
  XOR U34190 ( .A(n34477), .B(p_input[3670]), .Z(n34479) );
  XOR U34191 ( .A(n34481), .B(n34482), .Z(n34477) );
  AND U34192 ( .A(n34483), .B(n34484), .Z(n34482) );
  XNOR U34193 ( .A(p_input[3701]), .B(n34481), .Z(n34484) );
  XOR U34194 ( .A(n34481), .B(p_input[3669]), .Z(n34483) );
  XOR U34195 ( .A(n34485), .B(n34486), .Z(n34481) );
  AND U34196 ( .A(n34487), .B(n34488), .Z(n34486) );
  XNOR U34197 ( .A(p_input[3700]), .B(n34485), .Z(n34488) );
  XOR U34198 ( .A(n34485), .B(p_input[3668]), .Z(n34487) );
  XOR U34199 ( .A(n34489), .B(n34490), .Z(n34485) );
  AND U34200 ( .A(n34491), .B(n34492), .Z(n34490) );
  XNOR U34201 ( .A(p_input[3699]), .B(n34489), .Z(n34492) );
  XOR U34202 ( .A(n34489), .B(p_input[3667]), .Z(n34491) );
  XOR U34203 ( .A(n34493), .B(n34494), .Z(n34489) );
  AND U34204 ( .A(n34495), .B(n34496), .Z(n34494) );
  XNOR U34205 ( .A(p_input[3698]), .B(n34493), .Z(n34496) );
  XOR U34206 ( .A(n34493), .B(p_input[3666]), .Z(n34495) );
  XOR U34207 ( .A(n34497), .B(n34498), .Z(n34493) );
  AND U34208 ( .A(n34499), .B(n34500), .Z(n34498) );
  XNOR U34209 ( .A(p_input[3697]), .B(n34497), .Z(n34500) );
  XOR U34210 ( .A(n34497), .B(p_input[3665]), .Z(n34499) );
  XOR U34211 ( .A(n34501), .B(n34502), .Z(n34497) );
  AND U34212 ( .A(n34503), .B(n34504), .Z(n34502) );
  XNOR U34213 ( .A(p_input[3696]), .B(n34501), .Z(n34504) );
  XOR U34214 ( .A(n34501), .B(p_input[3664]), .Z(n34503) );
  XOR U34215 ( .A(n34505), .B(n34506), .Z(n34501) );
  AND U34216 ( .A(n34507), .B(n34508), .Z(n34506) );
  XNOR U34217 ( .A(p_input[3695]), .B(n34505), .Z(n34508) );
  XOR U34218 ( .A(n34505), .B(p_input[3663]), .Z(n34507) );
  XOR U34219 ( .A(n34509), .B(n34510), .Z(n34505) );
  AND U34220 ( .A(n34511), .B(n34512), .Z(n34510) );
  XNOR U34221 ( .A(p_input[3694]), .B(n34509), .Z(n34512) );
  XOR U34222 ( .A(n34509), .B(p_input[3662]), .Z(n34511) );
  XOR U34223 ( .A(n34513), .B(n34514), .Z(n34509) );
  AND U34224 ( .A(n34515), .B(n34516), .Z(n34514) );
  XNOR U34225 ( .A(p_input[3693]), .B(n34513), .Z(n34516) );
  XOR U34226 ( .A(n34513), .B(p_input[3661]), .Z(n34515) );
  XOR U34227 ( .A(n34517), .B(n34518), .Z(n34513) );
  AND U34228 ( .A(n34519), .B(n34520), .Z(n34518) );
  XNOR U34229 ( .A(p_input[3692]), .B(n34517), .Z(n34520) );
  XOR U34230 ( .A(n34517), .B(p_input[3660]), .Z(n34519) );
  XOR U34231 ( .A(n34521), .B(n34522), .Z(n34517) );
  AND U34232 ( .A(n34523), .B(n34524), .Z(n34522) );
  XNOR U34233 ( .A(p_input[3691]), .B(n34521), .Z(n34524) );
  XOR U34234 ( .A(n34521), .B(p_input[3659]), .Z(n34523) );
  XOR U34235 ( .A(n34525), .B(n34526), .Z(n34521) );
  AND U34236 ( .A(n34527), .B(n34528), .Z(n34526) );
  XNOR U34237 ( .A(p_input[3690]), .B(n34525), .Z(n34528) );
  XOR U34238 ( .A(n34525), .B(p_input[3658]), .Z(n34527) );
  XOR U34239 ( .A(n34529), .B(n34530), .Z(n34525) );
  AND U34240 ( .A(n34531), .B(n34532), .Z(n34530) );
  XNOR U34241 ( .A(p_input[3689]), .B(n34529), .Z(n34532) );
  XOR U34242 ( .A(n34529), .B(p_input[3657]), .Z(n34531) );
  XOR U34243 ( .A(n34533), .B(n34534), .Z(n34529) );
  AND U34244 ( .A(n34535), .B(n34536), .Z(n34534) );
  XNOR U34245 ( .A(p_input[3688]), .B(n34533), .Z(n34536) );
  XOR U34246 ( .A(n34533), .B(p_input[3656]), .Z(n34535) );
  XOR U34247 ( .A(n34537), .B(n34538), .Z(n34533) );
  AND U34248 ( .A(n34539), .B(n34540), .Z(n34538) );
  XNOR U34249 ( .A(p_input[3687]), .B(n34537), .Z(n34540) );
  XOR U34250 ( .A(n34537), .B(p_input[3655]), .Z(n34539) );
  XOR U34251 ( .A(n34541), .B(n34542), .Z(n34537) );
  AND U34252 ( .A(n34543), .B(n34544), .Z(n34542) );
  XNOR U34253 ( .A(p_input[3686]), .B(n34541), .Z(n34544) );
  XOR U34254 ( .A(n34541), .B(p_input[3654]), .Z(n34543) );
  XOR U34255 ( .A(n34545), .B(n34546), .Z(n34541) );
  AND U34256 ( .A(n34547), .B(n34548), .Z(n34546) );
  XNOR U34257 ( .A(p_input[3685]), .B(n34545), .Z(n34548) );
  XOR U34258 ( .A(n34545), .B(p_input[3653]), .Z(n34547) );
  XOR U34259 ( .A(n34549), .B(n34550), .Z(n34545) );
  AND U34260 ( .A(n34551), .B(n34552), .Z(n34550) );
  XNOR U34261 ( .A(p_input[3684]), .B(n34549), .Z(n34552) );
  XOR U34262 ( .A(n34549), .B(p_input[3652]), .Z(n34551) );
  XOR U34263 ( .A(n34553), .B(n34554), .Z(n34549) );
  AND U34264 ( .A(n34555), .B(n34556), .Z(n34554) );
  XNOR U34265 ( .A(p_input[3683]), .B(n34553), .Z(n34556) );
  XOR U34266 ( .A(n34553), .B(p_input[3651]), .Z(n34555) );
  XOR U34267 ( .A(n34557), .B(n34558), .Z(n34553) );
  AND U34268 ( .A(n34559), .B(n34560), .Z(n34558) );
  XNOR U34269 ( .A(p_input[3682]), .B(n34557), .Z(n34560) );
  XOR U34270 ( .A(n34557), .B(p_input[3650]), .Z(n34559) );
  XNOR U34271 ( .A(n34561), .B(n34562), .Z(n34557) );
  AND U34272 ( .A(n34563), .B(n34564), .Z(n34562) );
  XOR U34273 ( .A(p_input[3681]), .B(n34561), .Z(n34564) );
  XNOR U34274 ( .A(p_input[3649]), .B(n34561), .Z(n34563) );
  AND U34275 ( .A(p_input[3680]), .B(n34565), .Z(n34561) );
  IV U34276 ( .A(p_input[3648]), .Z(n34565) );
  XNOR U34277 ( .A(p_input[3584]), .B(n34566), .Z(n34159) );
  AND U34278 ( .A(n704), .B(n34567), .Z(n34566) );
  XOR U34279 ( .A(p_input[3616]), .B(p_input[3584]), .Z(n34567) );
  XOR U34280 ( .A(n34568), .B(n34569), .Z(n704) );
  AND U34281 ( .A(n34570), .B(n34571), .Z(n34569) );
  XNOR U34282 ( .A(p_input[3647]), .B(n34568), .Z(n34571) );
  XOR U34283 ( .A(n34568), .B(p_input[3615]), .Z(n34570) );
  XOR U34284 ( .A(n34572), .B(n34573), .Z(n34568) );
  AND U34285 ( .A(n34574), .B(n34575), .Z(n34573) );
  XNOR U34286 ( .A(p_input[3646]), .B(n34572), .Z(n34575) );
  XNOR U34287 ( .A(n34572), .B(n34174), .Z(n34574) );
  IV U34288 ( .A(p_input[3614]), .Z(n34174) );
  XOR U34289 ( .A(n34576), .B(n34577), .Z(n34572) );
  AND U34290 ( .A(n34578), .B(n34579), .Z(n34577) );
  XNOR U34291 ( .A(p_input[3645]), .B(n34576), .Z(n34579) );
  XNOR U34292 ( .A(n34576), .B(n34183), .Z(n34578) );
  IV U34293 ( .A(p_input[3613]), .Z(n34183) );
  XOR U34294 ( .A(n34580), .B(n34581), .Z(n34576) );
  AND U34295 ( .A(n34582), .B(n34583), .Z(n34581) );
  XNOR U34296 ( .A(p_input[3644]), .B(n34580), .Z(n34583) );
  XNOR U34297 ( .A(n34580), .B(n34192), .Z(n34582) );
  IV U34298 ( .A(p_input[3612]), .Z(n34192) );
  XOR U34299 ( .A(n34584), .B(n34585), .Z(n34580) );
  AND U34300 ( .A(n34586), .B(n34587), .Z(n34585) );
  XNOR U34301 ( .A(p_input[3643]), .B(n34584), .Z(n34587) );
  XNOR U34302 ( .A(n34584), .B(n34201), .Z(n34586) );
  IV U34303 ( .A(p_input[3611]), .Z(n34201) );
  XOR U34304 ( .A(n34588), .B(n34589), .Z(n34584) );
  AND U34305 ( .A(n34590), .B(n34591), .Z(n34589) );
  XNOR U34306 ( .A(p_input[3642]), .B(n34588), .Z(n34591) );
  XNOR U34307 ( .A(n34588), .B(n34210), .Z(n34590) );
  IV U34308 ( .A(p_input[3610]), .Z(n34210) );
  XOR U34309 ( .A(n34592), .B(n34593), .Z(n34588) );
  AND U34310 ( .A(n34594), .B(n34595), .Z(n34593) );
  XNOR U34311 ( .A(p_input[3641]), .B(n34592), .Z(n34595) );
  XNOR U34312 ( .A(n34592), .B(n34219), .Z(n34594) );
  IV U34313 ( .A(p_input[3609]), .Z(n34219) );
  XOR U34314 ( .A(n34596), .B(n34597), .Z(n34592) );
  AND U34315 ( .A(n34598), .B(n34599), .Z(n34597) );
  XNOR U34316 ( .A(p_input[3640]), .B(n34596), .Z(n34599) );
  XNOR U34317 ( .A(n34596), .B(n34228), .Z(n34598) );
  IV U34318 ( .A(p_input[3608]), .Z(n34228) );
  XOR U34319 ( .A(n34600), .B(n34601), .Z(n34596) );
  AND U34320 ( .A(n34602), .B(n34603), .Z(n34601) );
  XNOR U34321 ( .A(p_input[3639]), .B(n34600), .Z(n34603) );
  XNOR U34322 ( .A(n34600), .B(n34237), .Z(n34602) );
  IV U34323 ( .A(p_input[3607]), .Z(n34237) );
  XOR U34324 ( .A(n34604), .B(n34605), .Z(n34600) );
  AND U34325 ( .A(n34606), .B(n34607), .Z(n34605) );
  XNOR U34326 ( .A(p_input[3638]), .B(n34604), .Z(n34607) );
  XNOR U34327 ( .A(n34604), .B(n34246), .Z(n34606) );
  IV U34328 ( .A(p_input[3606]), .Z(n34246) );
  XOR U34329 ( .A(n34608), .B(n34609), .Z(n34604) );
  AND U34330 ( .A(n34610), .B(n34611), .Z(n34609) );
  XNOR U34331 ( .A(p_input[3637]), .B(n34608), .Z(n34611) );
  XNOR U34332 ( .A(n34608), .B(n34255), .Z(n34610) );
  IV U34333 ( .A(p_input[3605]), .Z(n34255) );
  XOR U34334 ( .A(n34612), .B(n34613), .Z(n34608) );
  AND U34335 ( .A(n34614), .B(n34615), .Z(n34613) );
  XNOR U34336 ( .A(p_input[3636]), .B(n34612), .Z(n34615) );
  XNOR U34337 ( .A(n34612), .B(n34264), .Z(n34614) );
  IV U34338 ( .A(p_input[3604]), .Z(n34264) );
  XOR U34339 ( .A(n34616), .B(n34617), .Z(n34612) );
  AND U34340 ( .A(n34618), .B(n34619), .Z(n34617) );
  XNOR U34341 ( .A(p_input[3635]), .B(n34616), .Z(n34619) );
  XNOR U34342 ( .A(n34616), .B(n34273), .Z(n34618) );
  IV U34343 ( .A(p_input[3603]), .Z(n34273) );
  XOR U34344 ( .A(n34620), .B(n34621), .Z(n34616) );
  AND U34345 ( .A(n34622), .B(n34623), .Z(n34621) );
  XNOR U34346 ( .A(p_input[3634]), .B(n34620), .Z(n34623) );
  XNOR U34347 ( .A(n34620), .B(n34282), .Z(n34622) );
  IV U34348 ( .A(p_input[3602]), .Z(n34282) );
  XOR U34349 ( .A(n34624), .B(n34625), .Z(n34620) );
  AND U34350 ( .A(n34626), .B(n34627), .Z(n34625) );
  XNOR U34351 ( .A(p_input[3633]), .B(n34624), .Z(n34627) );
  XNOR U34352 ( .A(n34624), .B(n34291), .Z(n34626) );
  IV U34353 ( .A(p_input[3601]), .Z(n34291) );
  XOR U34354 ( .A(n34628), .B(n34629), .Z(n34624) );
  AND U34355 ( .A(n34630), .B(n34631), .Z(n34629) );
  XNOR U34356 ( .A(p_input[3632]), .B(n34628), .Z(n34631) );
  XNOR U34357 ( .A(n34628), .B(n34300), .Z(n34630) );
  IV U34358 ( .A(p_input[3600]), .Z(n34300) );
  XOR U34359 ( .A(n34632), .B(n34633), .Z(n34628) );
  AND U34360 ( .A(n34634), .B(n34635), .Z(n34633) );
  XNOR U34361 ( .A(p_input[3631]), .B(n34632), .Z(n34635) );
  XNOR U34362 ( .A(n34632), .B(n34309), .Z(n34634) );
  IV U34363 ( .A(p_input[3599]), .Z(n34309) );
  XOR U34364 ( .A(n34636), .B(n34637), .Z(n34632) );
  AND U34365 ( .A(n34638), .B(n34639), .Z(n34637) );
  XNOR U34366 ( .A(p_input[3630]), .B(n34636), .Z(n34639) );
  XNOR U34367 ( .A(n34636), .B(n34318), .Z(n34638) );
  IV U34368 ( .A(p_input[3598]), .Z(n34318) );
  XOR U34369 ( .A(n34640), .B(n34641), .Z(n34636) );
  AND U34370 ( .A(n34642), .B(n34643), .Z(n34641) );
  XNOR U34371 ( .A(p_input[3629]), .B(n34640), .Z(n34643) );
  XNOR U34372 ( .A(n34640), .B(n34327), .Z(n34642) );
  IV U34373 ( .A(p_input[3597]), .Z(n34327) );
  XOR U34374 ( .A(n34644), .B(n34645), .Z(n34640) );
  AND U34375 ( .A(n34646), .B(n34647), .Z(n34645) );
  XNOR U34376 ( .A(p_input[3628]), .B(n34644), .Z(n34647) );
  XNOR U34377 ( .A(n34644), .B(n34336), .Z(n34646) );
  IV U34378 ( .A(p_input[3596]), .Z(n34336) );
  XOR U34379 ( .A(n34648), .B(n34649), .Z(n34644) );
  AND U34380 ( .A(n34650), .B(n34651), .Z(n34649) );
  XNOR U34381 ( .A(p_input[3627]), .B(n34648), .Z(n34651) );
  XNOR U34382 ( .A(n34648), .B(n34345), .Z(n34650) );
  IV U34383 ( .A(p_input[3595]), .Z(n34345) );
  XOR U34384 ( .A(n34652), .B(n34653), .Z(n34648) );
  AND U34385 ( .A(n34654), .B(n34655), .Z(n34653) );
  XNOR U34386 ( .A(p_input[3626]), .B(n34652), .Z(n34655) );
  XNOR U34387 ( .A(n34652), .B(n34354), .Z(n34654) );
  IV U34388 ( .A(p_input[3594]), .Z(n34354) );
  XOR U34389 ( .A(n34656), .B(n34657), .Z(n34652) );
  AND U34390 ( .A(n34658), .B(n34659), .Z(n34657) );
  XNOR U34391 ( .A(p_input[3625]), .B(n34656), .Z(n34659) );
  XNOR U34392 ( .A(n34656), .B(n34363), .Z(n34658) );
  IV U34393 ( .A(p_input[3593]), .Z(n34363) );
  XOR U34394 ( .A(n34660), .B(n34661), .Z(n34656) );
  AND U34395 ( .A(n34662), .B(n34663), .Z(n34661) );
  XNOR U34396 ( .A(p_input[3624]), .B(n34660), .Z(n34663) );
  XNOR U34397 ( .A(n34660), .B(n34372), .Z(n34662) );
  IV U34398 ( .A(p_input[3592]), .Z(n34372) );
  XOR U34399 ( .A(n34664), .B(n34665), .Z(n34660) );
  AND U34400 ( .A(n34666), .B(n34667), .Z(n34665) );
  XNOR U34401 ( .A(p_input[3623]), .B(n34664), .Z(n34667) );
  XNOR U34402 ( .A(n34664), .B(n34381), .Z(n34666) );
  IV U34403 ( .A(p_input[3591]), .Z(n34381) );
  XOR U34404 ( .A(n34668), .B(n34669), .Z(n34664) );
  AND U34405 ( .A(n34670), .B(n34671), .Z(n34669) );
  XNOR U34406 ( .A(p_input[3622]), .B(n34668), .Z(n34671) );
  XNOR U34407 ( .A(n34668), .B(n34390), .Z(n34670) );
  IV U34408 ( .A(p_input[3590]), .Z(n34390) );
  XOR U34409 ( .A(n34672), .B(n34673), .Z(n34668) );
  AND U34410 ( .A(n34674), .B(n34675), .Z(n34673) );
  XNOR U34411 ( .A(p_input[3621]), .B(n34672), .Z(n34675) );
  XNOR U34412 ( .A(n34672), .B(n34399), .Z(n34674) );
  IV U34413 ( .A(p_input[3589]), .Z(n34399) );
  XOR U34414 ( .A(n34676), .B(n34677), .Z(n34672) );
  AND U34415 ( .A(n34678), .B(n34679), .Z(n34677) );
  XNOR U34416 ( .A(p_input[3620]), .B(n34676), .Z(n34679) );
  XNOR U34417 ( .A(n34676), .B(n34408), .Z(n34678) );
  IV U34418 ( .A(p_input[3588]), .Z(n34408) );
  XOR U34419 ( .A(n34680), .B(n34681), .Z(n34676) );
  AND U34420 ( .A(n34682), .B(n34683), .Z(n34681) );
  XNOR U34421 ( .A(p_input[3619]), .B(n34680), .Z(n34683) );
  XNOR U34422 ( .A(n34680), .B(n34417), .Z(n34682) );
  IV U34423 ( .A(p_input[3587]), .Z(n34417) );
  XOR U34424 ( .A(n34684), .B(n34685), .Z(n34680) );
  AND U34425 ( .A(n34686), .B(n34687), .Z(n34685) );
  XNOR U34426 ( .A(p_input[3618]), .B(n34684), .Z(n34687) );
  XNOR U34427 ( .A(n34684), .B(n34426), .Z(n34686) );
  IV U34428 ( .A(p_input[3586]), .Z(n34426) );
  XNOR U34429 ( .A(n34688), .B(n34689), .Z(n34684) );
  AND U34430 ( .A(n34690), .B(n34691), .Z(n34689) );
  XOR U34431 ( .A(p_input[3617]), .B(n34688), .Z(n34691) );
  XNOR U34432 ( .A(p_input[3585]), .B(n34688), .Z(n34690) );
  AND U34433 ( .A(p_input[3616]), .B(n34692), .Z(n34688) );
  IV U34434 ( .A(p_input[3584]), .Z(n34692) );
  XOR U34435 ( .A(n34693), .B(n34694), .Z(n31049) );
  AND U34436 ( .A(n1025), .B(n34695), .Z(n34694) );
  XNOR U34437 ( .A(n34696), .B(n34693), .Z(n34695) );
  XOR U34438 ( .A(n34697), .B(n34698), .Z(n1025) );
  AND U34439 ( .A(n34699), .B(n34700), .Z(n34698) );
  XOR U34440 ( .A(n34697), .B(n31064), .Z(n34700) );
  XOR U34441 ( .A(n34701), .B(n34702), .Z(n31064) );
  AND U34442 ( .A(n879), .B(n34703), .Z(n34702) );
  XOR U34443 ( .A(n34704), .B(n34701), .Z(n34703) );
  XNOR U34444 ( .A(n31061), .B(n34697), .Z(n34699) );
  XOR U34445 ( .A(n34705), .B(n34706), .Z(n31061) );
  AND U34446 ( .A(n876), .B(n34707), .Z(n34706) );
  XOR U34447 ( .A(n34708), .B(n34705), .Z(n34707) );
  XOR U34448 ( .A(n34709), .B(n34710), .Z(n34697) );
  AND U34449 ( .A(n34711), .B(n34712), .Z(n34710) );
  XOR U34450 ( .A(n34709), .B(n31076), .Z(n34712) );
  XOR U34451 ( .A(n34713), .B(n34714), .Z(n31076) );
  AND U34452 ( .A(n879), .B(n34715), .Z(n34714) );
  XOR U34453 ( .A(n34716), .B(n34713), .Z(n34715) );
  XNOR U34454 ( .A(n31073), .B(n34709), .Z(n34711) );
  XOR U34455 ( .A(n34717), .B(n34718), .Z(n31073) );
  AND U34456 ( .A(n876), .B(n34719), .Z(n34718) );
  XOR U34457 ( .A(n34720), .B(n34717), .Z(n34719) );
  XOR U34458 ( .A(n34721), .B(n34722), .Z(n34709) );
  AND U34459 ( .A(n34723), .B(n34724), .Z(n34722) );
  XOR U34460 ( .A(n34721), .B(n31088), .Z(n34724) );
  XOR U34461 ( .A(n34725), .B(n34726), .Z(n31088) );
  AND U34462 ( .A(n879), .B(n34727), .Z(n34726) );
  XOR U34463 ( .A(n34728), .B(n34725), .Z(n34727) );
  XNOR U34464 ( .A(n31085), .B(n34721), .Z(n34723) );
  XOR U34465 ( .A(n34729), .B(n34730), .Z(n31085) );
  AND U34466 ( .A(n876), .B(n34731), .Z(n34730) );
  XOR U34467 ( .A(n34732), .B(n34729), .Z(n34731) );
  XOR U34468 ( .A(n34733), .B(n34734), .Z(n34721) );
  AND U34469 ( .A(n34735), .B(n34736), .Z(n34734) );
  XOR U34470 ( .A(n34733), .B(n31100), .Z(n34736) );
  XOR U34471 ( .A(n34737), .B(n34738), .Z(n31100) );
  AND U34472 ( .A(n879), .B(n34739), .Z(n34738) );
  XOR U34473 ( .A(n34740), .B(n34737), .Z(n34739) );
  XNOR U34474 ( .A(n31097), .B(n34733), .Z(n34735) );
  XOR U34475 ( .A(n34741), .B(n34742), .Z(n31097) );
  AND U34476 ( .A(n876), .B(n34743), .Z(n34742) );
  XOR U34477 ( .A(n34744), .B(n34741), .Z(n34743) );
  XOR U34478 ( .A(n34745), .B(n34746), .Z(n34733) );
  AND U34479 ( .A(n34747), .B(n34748), .Z(n34746) );
  XOR U34480 ( .A(n34745), .B(n31112), .Z(n34748) );
  XOR U34481 ( .A(n34749), .B(n34750), .Z(n31112) );
  AND U34482 ( .A(n879), .B(n34751), .Z(n34750) );
  XOR U34483 ( .A(n34752), .B(n34749), .Z(n34751) );
  XNOR U34484 ( .A(n31109), .B(n34745), .Z(n34747) );
  XOR U34485 ( .A(n34753), .B(n34754), .Z(n31109) );
  AND U34486 ( .A(n876), .B(n34755), .Z(n34754) );
  XOR U34487 ( .A(n34756), .B(n34753), .Z(n34755) );
  XOR U34488 ( .A(n34757), .B(n34758), .Z(n34745) );
  AND U34489 ( .A(n34759), .B(n34760), .Z(n34758) );
  XOR U34490 ( .A(n34757), .B(n31124), .Z(n34760) );
  XOR U34491 ( .A(n34761), .B(n34762), .Z(n31124) );
  AND U34492 ( .A(n879), .B(n34763), .Z(n34762) );
  XOR U34493 ( .A(n34764), .B(n34761), .Z(n34763) );
  XNOR U34494 ( .A(n31121), .B(n34757), .Z(n34759) );
  XOR U34495 ( .A(n34765), .B(n34766), .Z(n31121) );
  AND U34496 ( .A(n876), .B(n34767), .Z(n34766) );
  XOR U34497 ( .A(n34768), .B(n34765), .Z(n34767) );
  XOR U34498 ( .A(n34769), .B(n34770), .Z(n34757) );
  AND U34499 ( .A(n34771), .B(n34772), .Z(n34770) );
  XOR U34500 ( .A(n34769), .B(n31136), .Z(n34772) );
  XOR U34501 ( .A(n34773), .B(n34774), .Z(n31136) );
  AND U34502 ( .A(n879), .B(n34775), .Z(n34774) );
  XOR U34503 ( .A(n34776), .B(n34773), .Z(n34775) );
  XNOR U34504 ( .A(n31133), .B(n34769), .Z(n34771) );
  XOR U34505 ( .A(n34777), .B(n34778), .Z(n31133) );
  AND U34506 ( .A(n876), .B(n34779), .Z(n34778) );
  XOR U34507 ( .A(n34780), .B(n34777), .Z(n34779) );
  XOR U34508 ( .A(n34781), .B(n34782), .Z(n34769) );
  AND U34509 ( .A(n34783), .B(n34784), .Z(n34782) );
  XOR U34510 ( .A(n34781), .B(n31148), .Z(n34784) );
  XOR U34511 ( .A(n34785), .B(n34786), .Z(n31148) );
  AND U34512 ( .A(n879), .B(n34787), .Z(n34786) );
  XOR U34513 ( .A(n34788), .B(n34785), .Z(n34787) );
  XNOR U34514 ( .A(n31145), .B(n34781), .Z(n34783) );
  XOR U34515 ( .A(n34789), .B(n34790), .Z(n31145) );
  AND U34516 ( .A(n876), .B(n34791), .Z(n34790) );
  XOR U34517 ( .A(n34792), .B(n34789), .Z(n34791) );
  XOR U34518 ( .A(n34793), .B(n34794), .Z(n34781) );
  AND U34519 ( .A(n34795), .B(n34796), .Z(n34794) );
  XOR U34520 ( .A(n34793), .B(n31160), .Z(n34796) );
  XOR U34521 ( .A(n34797), .B(n34798), .Z(n31160) );
  AND U34522 ( .A(n879), .B(n34799), .Z(n34798) );
  XOR U34523 ( .A(n34800), .B(n34797), .Z(n34799) );
  XNOR U34524 ( .A(n31157), .B(n34793), .Z(n34795) );
  XOR U34525 ( .A(n34801), .B(n34802), .Z(n31157) );
  AND U34526 ( .A(n876), .B(n34803), .Z(n34802) );
  XOR U34527 ( .A(n34804), .B(n34801), .Z(n34803) );
  XOR U34528 ( .A(n34805), .B(n34806), .Z(n34793) );
  AND U34529 ( .A(n34807), .B(n34808), .Z(n34806) );
  XOR U34530 ( .A(n34805), .B(n31172), .Z(n34808) );
  XOR U34531 ( .A(n34809), .B(n34810), .Z(n31172) );
  AND U34532 ( .A(n879), .B(n34811), .Z(n34810) );
  XOR U34533 ( .A(n34812), .B(n34809), .Z(n34811) );
  XNOR U34534 ( .A(n31169), .B(n34805), .Z(n34807) );
  XOR U34535 ( .A(n34813), .B(n34814), .Z(n31169) );
  AND U34536 ( .A(n876), .B(n34815), .Z(n34814) );
  XOR U34537 ( .A(n34816), .B(n34813), .Z(n34815) );
  XOR U34538 ( .A(n34817), .B(n34818), .Z(n34805) );
  AND U34539 ( .A(n34819), .B(n34820), .Z(n34818) );
  XOR U34540 ( .A(n34817), .B(n31184), .Z(n34820) );
  XOR U34541 ( .A(n34821), .B(n34822), .Z(n31184) );
  AND U34542 ( .A(n879), .B(n34823), .Z(n34822) );
  XOR U34543 ( .A(n34824), .B(n34821), .Z(n34823) );
  XNOR U34544 ( .A(n31181), .B(n34817), .Z(n34819) );
  XOR U34545 ( .A(n34825), .B(n34826), .Z(n31181) );
  AND U34546 ( .A(n876), .B(n34827), .Z(n34826) );
  XOR U34547 ( .A(n34828), .B(n34825), .Z(n34827) );
  XOR U34548 ( .A(n34829), .B(n34830), .Z(n34817) );
  AND U34549 ( .A(n34831), .B(n34832), .Z(n34830) );
  XOR U34550 ( .A(n34829), .B(n31196), .Z(n34832) );
  XOR U34551 ( .A(n34833), .B(n34834), .Z(n31196) );
  AND U34552 ( .A(n879), .B(n34835), .Z(n34834) );
  XOR U34553 ( .A(n34836), .B(n34833), .Z(n34835) );
  XNOR U34554 ( .A(n31193), .B(n34829), .Z(n34831) );
  XOR U34555 ( .A(n34837), .B(n34838), .Z(n31193) );
  AND U34556 ( .A(n876), .B(n34839), .Z(n34838) );
  XOR U34557 ( .A(n34840), .B(n34837), .Z(n34839) );
  XOR U34558 ( .A(n34841), .B(n34842), .Z(n34829) );
  AND U34559 ( .A(n34843), .B(n34844), .Z(n34842) );
  XOR U34560 ( .A(n34841), .B(n31208), .Z(n34844) );
  XOR U34561 ( .A(n34845), .B(n34846), .Z(n31208) );
  AND U34562 ( .A(n879), .B(n34847), .Z(n34846) );
  XOR U34563 ( .A(n34848), .B(n34845), .Z(n34847) );
  XNOR U34564 ( .A(n31205), .B(n34841), .Z(n34843) );
  XOR U34565 ( .A(n34849), .B(n34850), .Z(n31205) );
  AND U34566 ( .A(n876), .B(n34851), .Z(n34850) );
  XOR U34567 ( .A(n34852), .B(n34849), .Z(n34851) );
  XOR U34568 ( .A(n34853), .B(n34854), .Z(n34841) );
  AND U34569 ( .A(n34855), .B(n34856), .Z(n34854) );
  XOR U34570 ( .A(n34853), .B(n31220), .Z(n34856) );
  XOR U34571 ( .A(n34857), .B(n34858), .Z(n31220) );
  AND U34572 ( .A(n879), .B(n34859), .Z(n34858) );
  XOR U34573 ( .A(n34860), .B(n34857), .Z(n34859) );
  XNOR U34574 ( .A(n31217), .B(n34853), .Z(n34855) );
  XOR U34575 ( .A(n34861), .B(n34862), .Z(n31217) );
  AND U34576 ( .A(n876), .B(n34863), .Z(n34862) );
  XOR U34577 ( .A(n34864), .B(n34861), .Z(n34863) );
  XOR U34578 ( .A(n34865), .B(n34866), .Z(n34853) );
  AND U34579 ( .A(n34867), .B(n34868), .Z(n34866) );
  XOR U34580 ( .A(n34865), .B(n31232), .Z(n34868) );
  XOR U34581 ( .A(n34869), .B(n34870), .Z(n31232) );
  AND U34582 ( .A(n879), .B(n34871), .Z(n34870) );
  XOR U34583 ( .A(n34872), .B(n34869), .Z(n34871) );
  XNOR U34584 ( .A(n31229), .B(n34865), .Z(n34867) );
  XOR U34585 ( .A(n34873), .B(n34874), .Z(n31229) );
  AND U34586 ( .A(n876), .B(n34875), .Z(n34874) );
  XOR U34587 ( .A(n34876), .B(n34873), .Z(n34875) );
  XOR U34588 ( .A(n34877), .B(n34878), .Z(n34865) );
  AND U34589 ( .A(n34879), .B(n34880), .Z(n34878) );
  XOR U34590 ( .A(n34877), .B(n31244), .Z(n34880) );
  XOR U34591 ( .A(n34881), .B(n34882), .Z(n31244) );
  AND U34592 ( .A(n879), .B(n34883), .Z(n34882) );
  XOR U34593 ( .A(n34884), .B(n34881), .Z(n34883) );
  XNOR U34594 ( .A(n31241), .B(n34877), .Z(n34879) );
  XOR U34595 ( .A(n34885), .B(n34886), .Z(n31241) );
  AND U34596 ( .A(n876), .B(n34887), .Z(n34886) );
  XOR U34597 ( .A(n34888), .B(n34885), .Z(n34887) );
  XOR U34598 ( .A(n34889), .B(n34890), .Z(n34877) );
  AND U34599 ( .A(n34891), .B(n34892), .Z(n34890) );
  XOR U34600 ( .A(n34889), .B(n31256), .Z(n34892) );
  XOR U34601 ( .A(n34893), .B(n34894), .Z(n31256) );
  AND U34602 ( .A(n879), .B(n34895), .Z(n34894) );
  XOR U34603 ( .A(n34896), .B(n34893), .Z(n34895) );
  XNOR U34604 ( .A(n31253), .B(n34889), .Z(n34891) );
  XOR U34605 ( .A(n34897), .B(n34898), .Z(n31253) );
  AND U34606 ( .A(n876), .B(n34899), .Z(n34898) );
  XOR U34607 ( .A(n34900), .B(n34897), .Z(n34899) );
  XOR U34608 ( .A(n34901), .B(n34902), .Z(n34889) );
  AND U34609 ( .A(n34903), .B(n34904), .Z(n34902) );
  XOR U34610 ( .A(n34901), .B(n31268), .Z(n34904) );
  XOR U34611 ( .A(n34905), .B(n34906), .Z(n31268) );
  AND U34612 ( .A(n879), .B(n34907), .Z(n34906) );
  XOR U34613 ( .A(n34908), .B(n34905), .Z(n34907) );
  XNOR U34614 ( .A(n31265), .B(n34901), .Z(n34903) );
  XOR U34615 ( .A(n34909), .B(n34910), .Z(n31265) );
  AND U34616 ( .A(n876), .B(n34911), .Z(n34910) );
  XOR U34617 ( .A(n34912), .B(n34909), .Z(n34911) );
  XOR U34618 ( .A(n34913), .B(n34914), .Z(n34901) );
  AND U34619 ( .A(n34915), .B(n34916), .Z(n34914) );
  XOR U34620 ( .A(n34913), .B(n31280), .Z(n34916) );
  XOR U34621 ( .A(n34917), .B(n34918), .Z(n31280) );
  AND U34622 ( .A(n879), .B(n34919), .Z(n34918) );
  XOR U34623 ( .A(n34920), .B(n34917), .Z(n34919) );
  XNOR U34624 ( .A(n31277), .B(n34913), .Z(n34915) );
  XOR U34625 ( .A(n34921), .B(n34922), .Z(n31277) );
  AND U34626 ( .A(n876), .B(n34923), .Z(n34922) );
  XOR U34627 ( .A(n34924), .B(n34921), .Z(n34923) );
  XOR U34628 ( .A(n34925), .B(n34926), .Z(n34913) );
  AND U34629 ( .A(n34927), .B(n34928), .Z(n34926) );
  XOR U34630 ( .A(n34925), .B(n31292), .Z(n34928) );
  XOR U34631 ( .A(n34929), .B(n34930), .Z(n31292) );
  AND U34632 ( .A(n879), .B(n34931), .Z(n34930) );
  XOR U34633 ( .A(n34932), .B(n34929), .Z(n34931) );
  XNOR U34634 ( .A(n31289), .B(n34925), .Z(n34927) );
  XOR U34635 ( .A(n34933), .B(n34934), .Z(n31289) );
  AND U34636 ( .A(n876), .B(n34935), .Z(n34934) );
  XOR U34637 ( .A(n34936), .B(n34933), .Z(n34935) );
  XOR U34638 ( .A(n34937), .B(n34938), .Z(n34925) );
  AND U34639 ( .A(n34939), .B(n34940), .Z(n34938) );
  XOR U34640 ( .A(n34937), .B(n31304), .Z(n34940) );
  XOR U34641 ( .A(n34941), .B(n34942), .Z(n31304) );
  AND U34642 ( .A(n879), .B(n34943), .Z(n34942) );
  XOR U34643 ( .A(n34944), .B(n34941), .Z(n34943) );
  XNOR U34644 ( .A(n31301), .B(n34937), .Z(n34939) );
  XOR U34645 ( .A(n34945), .B(n34946), .Z(n31301) );
  AND U34646 ( .A(n876), .B(n34947), .Z(n34946) );
  XOR U34647 ( .A(n34948), .B(n34945), .Z(n34947) );
  XOR U34648 ( .A(n34949), .B(n34950), .Z(n34937) );
  AND U34649 ( .A(n34951), .B(n34952), .Z(n34950) );
  XOR U34650 ( .A(n34949), .B(n31316), .Z(n34952) );
  XOR U34651 ( .A(n34953), .B(n34954), .Z(n31316) );
  AND U34652 ( .A(n879), .B(n34955), .Z(n34954) );
  XOR U34653 ( .A(n34956), .B(n34953), .Z(n34955) );
  XNOR U34654 ( .A(n31313), .B(n34949), .Z(n34951) );
  XOR U34655 ( .A(n34957), .B(n34958), .Z(n31313) );
  AND U34656 ( .A(n876), .B(n34959), .Z(n34958) );
  XOR U34657 ( .A(n34960), .B(n34957), .Z(n34959) );
  XOR U34658 ( .A(n34961), .B(n34962), .Z(n34949) );
  AND U34659 ( .A(n34963), .B(n34964), .Z(n34962) );
  XOR U34660 ( .A(n34961), .B(n31328), .Z(n34964) );
  XOR U34661 ( .A(n34965), .B(n34966), .Z(n31328) );
  AND U34662 ( .A(n879), .B(n34967), .Z(n34966) );
  XOR U34663 ( .A(n34968), .B(n34965), .Z(n34967) );
  XNOR U34664 ( .A(n31325), .B(n34961), .Z(n34963) );
  XOR U34665 ( .A(n34969), .B(n34970), .Z(n31325) );
  AND U34666 ( .A(n876), .B(n34971), .Z(n34970) );
  XOR U34667 ( .A(n34972), .B(n34969), .Z(n34971) );
  XOR U34668 ( .A(n34973), .B(n34974), .Z(n34961) );
  AND U34669 ( .A(n34975), .B(n34976), .Z(n34974) );
  XOR U34670 ( .A(n34973), .B(n31340), .Z(n34976) );
  XOR U34671 ( .A(n34977), .B(n34978), .Z(n31340) );
  AND U34672 ( .A(n879), .B(n34979), .Z(n34978) );
  XOR U34673 ( .A(n34980), .B(n34977), .Z(n34979) );
  XNOR U34674 ( .A(n31337), .B(n34973), .Z(n34975) );
  XOR U34675 ( .A(n34981), .B(n34982), .Z(n31337) );
  AND U34676 ( .A(n876), .B(n34983), .Z(n34982) );
  XOR U34677 ( .A(n34984), .B(n34981), .Z(n34983) );
  XOR U34678 ( .A(n34985), .B(n34986), .Z(n34973) );
  AND U34679 ( .A(n34987), .B(n34988), .Z(n34986) );
  XOR U34680 ( .A(n34985), .B(n31352), .Z(n34988) );
  XOR U34681 ( .A(n34989), .B(n34990), .Z(n31352) );
  AND U34682 ( .A(n879), .B(n34991), .Z(n34990) );
  XOR U34683 ( .A(n34992), .B(n34989), .Z(n34991) );
  XNOR U34684 ( .A(n31349), .B(n34985), .Z(n34987) );
  XOR U34685 ( .A(n34993), .B(n34994), .Z(n31349) );
  AND U34686 ( .A(n876), .B(n34995), .Z(n34994) );
  XOR U34687 ( .A(n34996), .B(n34993), .Z(n34995) );
  XOR U34688 ( .A(n34997), .B(n34998), .Z(n34985) );
  AND U34689 ( .A(n34999), .B(n35000), .Z(n34998) );
  XOR U34690 ( .A(n34997), .B(n31364), .Z(n35000) );
  XOR U34691 ( .A(n35001), .B(n35002), .Z(n31364) );
  AND U34692 ( .A(n879), .B(n35003), .Z(n35002) );
  XOR U34693 ( .A(n35004), .B(n35001), .Z(n35003) );
  XNOR U34694 ( .A(n31361), .B(n34997), .Z(n34999) );
  XOR U34695 ( .A(n35005), .B(n35006), .Z(n31361) );
  AND U34696 ( .A(n876), .B(n35007), .Z(n35006) );
  XOR U34697 ( .A(n35008), .B(n35005), .Z(n35007) );
  XOR U34698 ( .A(n35009), .B(n35010), .Z(n34997) );
  AND U34699 ( .A(n35011), .B(n35012), .Z(n35010) );
  XOR U34700 ( .A(n35009), .B(n31376), .Z(n35012) );
  XOR U34701 ( .A(n35013), .B(n35014), .Z(n31376) );
  AND U34702 ( .A(n879), .B(n35015), .Z(n35014) );
  XOR U34703 ( .A(n35016), .B(n35013), .Z(n35015) );
  XNOR U34704 ( .A(n31373), .B(n35009), .Z(n35011) );
  XOR U34705 ( .A(n35017), .B(n35018), .Z(n31373) );
  AND U34706 ( .A(n876), .B(n35019), .Z(n35018) );
  XOR U34707 ( .A(n35020), .B(n35017), .Z(n35019) );
  XOR U34708 ( .A(n35021), .B(n35022), .Z(n35009) );
  AND U34709 ( .A(n35023), .B(n35024), .Z(n35022) );
  XOR U34710 ( .A(n35021), .B(n31388), .Z(n35024) );
  XOR U34711 ( .A(n35025), .B(n35026), .Z(n31388) );
  AND U34712 ( .A(n879), .B(n35027), .Z(n35026) );
  XOR U34713 ( .A(n35028), .B(n35025), .Z(n35027) );
  XNOR U34714 ( .A(n31385), .B(n35021), .Z(n35023) );
  XOR U34715 ( .A(n35029), .B(n35030), .Z(n31385) );
  AND U34716 ( .A(n876), .B(n35031), .Z(n35030) );
  XOR U34717 ( .A(n35032), .B(n35029), .Z(n35031) );
  XOR U34718 ( .A(n35033), .B(n35034), .Z(n35021) );
  AND U34719 ( .A(n35035), .B(n35036), .Z(n35034) );
  XOR U34720 ( .A(n35033), .B(n31400), .Z(n35036) );
  XOR U34721 ( .A(n35037), .B(n35038), .Z(n31400) );
  AND U34722 ( .A(n879), .B(n35039), .Z(n35038) );
  XOR U34723 ( .A(n35040), .B(n35037), .Z(n35039) );
  XNOR U34724 ( .A(n31397), .B(n35033), .Z(n35035) );
  XOR U34725 ( .A(n35041), .B(n35042), .Z(n31397) );
  AND U34726 ( .A(n876), .B(n35043), .Z(n35042) );
  XOR U34727 ( .A(n35044), .B(n35041), .Z(n35043) );
  XOR U34728 ( .A(n35045), .B(n35046), .Z(n35033) );
  AND U34729 ( .A(n35047), .B(n35048), .Z(n35046) );
  XOR U34730 ( .A(n35045), .B(n31412), .Z(n35048) );
  XOR U34731 ( .A(n35049), .B(n35050), .Z(n31412) );
  AND U34732 ( .A(n879), .B(n35051), .Z(n35050) );
  XOR U34733 ( .A(n35052), .B(n35049), .Z(n35051) );
  XNOR U34734 ( .A(n31409), .B(n35045), .Z(n35047) );
  XOR U34735 ( .A(n35053), .B(n35054), .Z(n31409) );
  AND U34736 ( .A(n876), .B(n35055), .Z(n35054) );
  XOR U34737 ( .A(n35056), .B(n35053), .Z(n35055) );
  XOR U34738 ( .A(n35057), .B(n35058), .Z(n35045) );
  AND U34739 ( .A(n35059), .B(n35060), .Z(n35058) );
  XNOR U34740 ( .A(n35061), .B(n31425), .Z(n35060) );
  XOR U34741 ( .A(n35062), .B(n35063), .Z(n31425) );
  AND U34742 ( .A(n879), .B(n35064), .Z(n35063) );
  XOR U34743 ( .A(n35062), .B(n35065), .Z(n35064) );
  XNOR U34744 ( .A(n31422), .B(n35057), .Z(n35059) );
  XOR U34745 ( .A(n35066), .B(n35067), .Z(n31422) );
  AND U34746 ( .A(n876), .B(n35068), .Z(n35067) );
  XOR U34747 ( .A(n35066), .B(n35069), .Z(n35068) );
  IV U34748 ( .A(n35061), .Z(n35057) );
  AND U34749 ( .A(n34693), .B(n34696), .Z(n35061) );
  XNOR U34750 ( .A(n35070), .B(n35071), .Z(n34696) );
  AND U34751 ( .A(n879), .B(n35072), .Z(n35071) );
  XNOR U34752 ( .A(n35073), .B(n35070), .Z(n35072) );
  XOR U34753 ( .A(n35074), .B(n35075), .Z(n879) );
  AND U34754 ( .A(n35076), .B(n35077), .Z(n35075) );
  XOR U34755 ( .A(n35074), .B(n34704), .Z(n35077) );
  XNOR U34756 ( .A(n35078), .B(n35079), .Z(n34704) );
  AND U34757 ( .A(n35080), .B(n575), .Z(n35079) );
  AND U34758 ( .A(n35078), .B(n35081), .Z(n35080) );
  XNOR U34759 ( .A(n34701), .B(n35074), .Z(n35076) );
  XOR U34760 ( .A(n35082), .B(n35083), .Z(n34701) );
  AND U34761 ( .A(n35084), .B(n573), .Z(n35083) );
  NOR U34762 ( .A(n35082), .B(n35085), .Z(n35084) );
  XOR U34763 ( .A(n35086), .B(n35087), .Z(n35074) );
  AND U34764 ( .A(n35088), .B(n35089), .Z(n35087) );
  XOR U34765 ( .A(n35086), .B(n34716), .Z(n35089) );
  XOR U34766 ( .A(n35090), .B(n35091), .Z(n34716) );
  AND U34767 ( .A(n575), .B(n35092), .Z(n35091) );
  XOR U34768 ( .A(n35093), .B(n35090), .Z(n35092) );
  XNOR U34769 ( .A(n34713), .B(n35086), .Z(n35088) );
  XOR U34770 ( .A(n35094), .B(n35095), .Z(n34713) );
  AND U34771 ( .A(n573), .B(n35096), .Z(n35095) );
  XOR U34772 ( .A(n35097), .B(n35094), .Z(n35096) );
  XOR U34773 ( .A(n35098), .B(n35099), .Z(n35086) );
  AND U34774 ( .A(n35100), .B(n35101), .Z(n35099) );
  XOR U34775 ( .A(n35098), .B(n34728), .Z(n35101) );
  XOR U34776 ( .A(n35102), .B(n35103), .Z(n34728) );
  AND U34777 ( .A(n575), .B(n35104), .Z(n35103) );
  XOR U34778 ( .A(n35105), .B(n35102), .Z(n35104) );
  XNOR U34779 ( .A(n34725), .B(n35098), .Z(n35100) );
  XOR U34780 ( .A(n35106), .B(n35107), .Z(n34725) );
  AND U34781 ( .A(n573), .B(n35108), .Z(n35107) );
  XOR U34782 ( .A(n35109), .B(n35106), .Z(n35108) );
  XOR U34783 ( .A(n35110), .B(n35111), .Z(n35098) );
  AND U34784 ( .A(n35112), .B(n35113), .Z(n35111) );
  XOR U34785 ( .A(n35110), .B(n34740), .Z(n35113) );
  XOR U34786 ( .A(n35114), .B(n35115), .Z(n34740) );
  AND U34787 ( .A(n575), .B(n35116), .Z(n35115) );
  XOR U34788 ( .A(n35117), .B(n35114), .Z(n35116) );
  XNOR U34789 ( .A(n34737), .B(n35110), .Z(n35112) );
  XOR U34790 ( .A(n35118), .B(n35119), .Z(n34737) );
  AND U34791 ( .A(n573), .B(n35120), .Z(n35119) );
  XOR U34792 ( .A(n35121), .B(n35118), .Z(n35120) );
  XOR U34793 ( .A(n35122), .B(n35123), .Z(n35110) );
  AND U34794 ( .A(n35124), .B(n35125), .Z(n35123) );
  XOR U34795 ( .A(n35122), .B(n34752), .Z(n35125) );
  XOR U34796 ( .A(n35126), .B(n35127), .Z(n34752) );
  AND U34797 ( .A(n575), .B(n35128), .Z(n35127) );
  XOR U34798 ( .A(n35129), .B(n35126), .Z(n35128) );
  XNOR U34799 ( .A(n34749), .B(n35122), .Z(n35124) );
  XOR U34800 ( .A(n35130), .B(n35131), .Z(n34749) );
  AND U34801 ( .A(n573), .B(n35132), .Z(n35131) );
  XOR U34802 ( .A(n35133), .B(n35130), .Z(n35132) );
  XOR U34803 ( .A(n35134), .B(n35135), .Z(n35122) );
  AND U34804 ( .A(n35136), .B(n35137), .Z(n35135) );
  XOR U34805 ( .A(n35134), .B(n34764), .Z(n35137) );
  XOR U34806 ( .A(n35138), .B(n35139), .Z(n34764) );
  AND U34807 ( .A(n575), .B(n35140), .Z(n35139) );
  XOR U34808 ( .A(n35141), .B(n35138), .Z(n35140) );
  XNOR U34809 ( .A(n34761), .B(n35134), .Z(n35136) );
  XOR U34810 ( .A(n35142), .B(n35143), .Z(n34761) );
  AND U34811 ( .A(n573), .B(n35144), .Z(n35143) );
  XOR U34812 ( .A(n35145), .B(n35142), .Z(n35144) );
  XOR U34813 ( .A(n35146), .B(n35147), .Z(n35134) );
  AND U34814 ( .A(n35148), .B(n35149), .Z(n35147) );
  XOR U34815 ( .A(n35146), .B(n34776), .Z(n35149) );
  XOR U34816 ( .A(n35150), .B(n35151), .Z(n34776) );
  AND U34817 ( .A(n575), .B(n35152), .Z(n35151) );
  XOR U34818 ( .A(n35153), .B(n35150), .Z(n35152) );
  XNOR U34819 ( .A(n34773), .B(n35146), .Z(n35148) );
  XOR U34820 ( .A(n35154), .B(n35155), .Z(n34773) );
  AND U34821 ( .A(n573), .B(n35156), .Z(n35155) );
  XOR U34822 ( .A(n35157), .B(n35154), .Z(n35156) );
  XOR U34823 ( .A(n35158), .B(n35159), .Z(n35146) );
  AND U34824 ( .A(n35160), .B(n35161), .Z(n35159) );
  XOR U34825 ( .A(n35158), .B(n34788), .Z(n35161) );
  XOR U34826 ( .A(n35162), .B(n35163), .Z(n34788) );
  AND U34827 ( .A(n575), .B(n35164), .Z(n35163) );
  XOR U34828 ( .A(n35165), .B(n35162), .Z(n35164) );
  XNOR U34829 ( .A(n34785), .B(n35158), .Z(n35160) );
  XOR U34830 ( .A(n35166), .B(n35167), .Z(n34785) );
  AND U34831 ( .A(n573), .B(n35168), .Z(n35167) );
  XOR U34832 ( .A(n35169), .B(n35166), .Z(n35168) );
  XOR U34833 ( .A(n35170), .B(n35171), .Z(n35158) );
  AND U34834 ( .A(n35172), .B(n35173), .Z(n35171) );
  XOR U34835 ( .A(n35170), .B(n34800), .Z(n35173) );
  XOR U34836 ( .A(n35174), .B(n35175), .Z(n34800) );
  AND U34837 ( .A(n575), .B(n35176), .Z(n35175) );
  XOR U34838 ( .A(n35177), .B(n35174), .Z(n35176) );
  XNOR U34839 ( .A(n34797), .B(n35170), .Z(n35172) );
  XOR U34840 ( .A(n35178), .B(n35179), .Z(n34797) );
  AND U34841 ( .A(n573), .B(n35180), .Z(n35179) );
  XOR U34842 ( .A(n35181), .B(n35178), .Z(n35180) );
  XOR U34843 ( .A(n35182), .B(n35183), .Z(n35170) );
  AND U34844 ( .A(n35184), .B(n35185), .Z(n35183) );
  XOR U34845 ( .A(n35182), .B(n34812), .Z(n35185) );
  XOR U34846 ( .A(n35186), .B(n35187), .Z(n34812) );
  AND U34847 ( .A(n575), .B(n35188), .Z(n35187) );
  XOR U34848 ( .A(n35189), .B(n35186), .Z(n35188) );
  XNOR U34849 ( .A(n34809), .B(n35182), .Z(n35184) );
  XOR U34850 ( .A(n35190), .B(n35191), .Z(n34809) );
  AND U34851 ( .A(n573), .B(n35192), .Z(n35191) );
  XOR U34852 ( .A(n35193), .B(n35190), .Z(n35192) );
  XOR U34853 ( .A(n35194), .B(n35195), .Z(n35182) );
  AND U34854 ( .A(n35196), .B(n35197), .Z(n35195) );
  XOR U34855 ( .A(n35194), .B(n34824), .Z(n35197) );
  XOR U34856 ( .A(n35198), .B(n35199), .Z(n34824) );
  AND U34857 ( .A(n575), .B(n35200), .Z(n35199) );
  XOR U34858 ( .A(n35201), .B(n35198), .Z(n35200) );
  XNOR U34859 ( .A(n34821), .B(n35194), .Z(n35196) );
  XOR U34860 ( .A(n35202), .B(n35203), .Z(n34821) );
  AND U34861 ( .A(n573), .B(n35204), .Z(n35203) );
  XOR U34862 ( .A(n35205), .B(n35202), .Z(n35204) );
  XOR U34863 ( .A(n35206), .B(n35207), .Z(n35194) );
  AND U34864 ( .A(n35208), .B(n35209), .Z(n35207) );
  XOR U34865 ( .A(n35206), .B(n34836), .Z(n35209) );
  XOR U34866 ( .A(n35210), .B(n35211), .Z(n34836) );
  AND U34867 ( .A(n575), .B(n35212), .Z(n35211) );
  XOR U34868 ( .A(n35213), .B(n35210), .Z(n35212) );
  XNOR U34869 ( .A(n34833), .B(n35206), .Z(n35208) );
  XOR U34870 ( .A(n35214), .B(n35215), .Z(n34833) );
  AND U34871 ( .A(n573), .B(n35216), .Z(n35215) );
  XOR U34872 ( .A(n35217), .B(n35214), .Z(n35216) );
  XOR U34873 ( .A(n35218), .B(n35219), .Z(n35206) );
  AND U34874 ( .A(n35220), .B(n35221), .Z(n35219) );
  XOR U34875 ( .A(n35218), .B(n34848), .Z(n35221) );
  XOR U34876 ( .A(n35222), .B(n35223), .Z(n34848) );
  AND U34877 ( .A(n575), .B(n35224), .Z(n35223) );
  XOR U34878 ( .A(n35225), .B(n35222), .Z(n35224) );
  XNOR U34879 ( .A(n34845), .B(n35218), .Z(n35220) );
  XOR U34880 ( .A(n35226), .B(n35227), .Z(n34845) );
  AND U34881 ( .A(n573), .B(n35228), .Z(n35227) );
  XOR U34882 ( .A(n35229), .B(n35226), .Z(n35228) );
  XOR U34883 ( .A(n35230), .B(n35231), .Z(n35218) );
  AND U34884 ( .A(n35232), .B(n35233), .Z(n35231) );
  XOR U34885 ( .A(n35230), .B(n34860), .Z(n35233) );
  XOR U34886 ( .A(n35234), .B(n35235), .Z(n34860) );
  AND U34887 ( .A(n575), .B(n35236), .Z(n35235) );
  XOR U34888 ( .A(n35237), .B(n35234), .Z(n35236) );
  XNOR U34889 ( .A(n34857), .B(n35230), .Z(n35232) );
  XOR U34890 ( .A(n35238), .B(n35239), .Z(n34857) );
  AND U34891 ( .A(n573), .B(n35240), .Z(n35239) );
  XOR U34892 ( .A(n35241), .B(n35238), .Z(n35240) );
  XOR U34893 ( .A(n35242), .B(n35243), .Z(n35230) );
  AND U34894 ( .A(n35244), .B(n35245), .Z(n35243) );
  XOR U34895 ( .A(n35242), .B(n34872), .Z(n35245) );
  XOR U34896 ( .A(n35246), .B(n35247), .Z(n34872) );
  AND U34897 ( .A(n575), .B(n35248), .Z(n35247) );
  XOR U34898 ( .A(n35249), .B(n35246), .Z(n35248) );
  XNOR U34899 ( .A(n34869), .B(n35242), .Z(n35244) );
  XOR U34900 ( .A(n35250), .B(n35251), .Z(n34869) );
  AND U34901 ( .A(n573), .B(n35252), .Z(n35251) );
  XOR U34902 ( .A(n35253), .B(n35250), .Z(n35252) );
  XOR U34903 ( .A(n35254), .B(n35255), .Z(n35242) );
  AND U34904 ( .A(n35256), .B(n35257), .Z(n35255) );
  XOR U34905 ( .A(n35254), .B(n34884), .Z(n35257) );
  XOR U34906 ( .A(n35258), .B(n35259), .Z(n34884) );
  AND U34907 ( .A(n575), .B(n35260), .Z(n35259) );
  XOR U34908 ( .A(n35261), .B(n35258), .Z(n35260) );
  XNOR U34909 ( .A(n34881), .B(n35254), .Z(n35256) );
  XOR U34910 ( .A(n35262), .B(n35263), .Z(n34881) );
  AND U34911 ( .A(n573), .B(n35264), .Z(n35263) );
  XOR U34912 ( .A(n35265), .B(n35262), .Z(n35264) );
  XOR U34913 ( .A(n35266), .B(n35267), .Z(n35254) );
  AND U34914 ( .A(n35268), .B(n35269), .Z(n35267) );
  XOR U34915 ( .A(n35266), .B(n34896), .Z(n35269) );
  XOR U34916 ( .A(n35270), .B(n35271), .Z(n34896) );
  AND U34917 ( .A(n575), .B(n35272), .Z(n35271) );
  XOR U34918 ( .A(n35273), .B(n35270), .Z(n35272) );
  XNOR U34919 ( .A(n34893), .B(n35266), .Z(n35268) );
  XOR U34920 ( .A(n35274), .B(n35275), .Z(n34893) );
  AND U34921 ( .A(n573), .B(n35276), .Z(n35275) );
  XOR U34922 ( .A(n35277), .B(n35274), .Z(n35276) );
  XOR U34923 ( .A(n35278), .B(n35279), .Z(n35266) );
  AND U34924 ( .A(n35280), .B(n35281), .Z(n35279) );
  XOR U34925 ( .A(n35278), .B(n34908), .Z(n35281) );
  XOR U34926 ( .A(n35282), .B(n35283), .Z(n34908) );
  AND U34927 ( .A(n575), .B(n35284), .Z(n35283) );
  XOR U34928 ( .A(n35285), .B(n35282), .Z(n35284) );
  XNOR U34929 ( .A(n34905), .B(n35278), .Z(n35280) );
  XOR U34930 ( .A(n35286), .B(n35287), .Z(n34905) );
  AND U34931 ( .A(n573), .B(n35288), .Z(n35287) );
  XOR U34932 ( .A(n35289), .B(n35286), .Z(n35288) );
  XOR U34933 ( .A(n35290), .B(n35291), .Z(n35278) );
  AND U34934 ( .A(n35292), .B(n35293), .Z(n35291) );
  XOR U34935 ( .A(n35290), .B(n34920), .Z(n35293) );
  XOR U34936 ( .A(n35294), .B(n35295), .Z(n34920) );
  AND U34937 ( .A(n575), .B(n35296), .Z(n35295) );
  XOR U34938 ( .A(n35297), .B(n35294), .Z(n35296) );
  XNOR U34939 ( .A(n34917), .B(n35290), .Z(n35292) );
  XOR U34940 ( .A(n35298), .B(n35299), .Z(n34917) );
  AND U34941 ( .A(n573), .B(n35300), .Z(n35299) );
  XOR U34942 ( .A(n35301), .B(n35298), .Z(n35300) );
  XOR U34943 ( .A(n35302), .B(n35303), .Z(n35290) );
  AND U34944 ( .A(n35304), .B(n35305), .Z(n35303) );
  XOR U34945 ( .A(n35302), .B(n34932), .Z(n35305) );
  XOR U34946 ( .A(n35306), .B(n35307), .Z(n34932) );
  AND U34947 ( .A(n575), .B(n35308), .Z(n35307) );
  XOR U34948 ( .A(n35309), .B(n35306), .Z(n35308) );
  XNOR U34949 ( .A(n34929), .B(n35302), .Z(n35304) );
  XOR U34950 ( .A(n35310), .B(n35311), .Z(n34929) );
  AND U34951 ( .A(n573), .B(n35312), .Z(n35311) );
  XOR U34952 ( .A(n35313), .B(n35310), .Z(n35312) );
  XOR U34953 ( .A(n35314), .B(n35315), .Z(n35302) );
  AND U34954 ( .A(n35316), .B(n35317), .Z(n35315) );
  XOR U34955 ( .A(n35314), .B(n34944), .Z(n35317) );
  XOR U34956 ( .A(n35318), .B(n35319), .Z(n34944) );
  AND U34957 ( .A(n575), .B(n35320), .Z(n35319) );
  XOR U34958 ( .A(n35321), .B(n35318), .Z(n35320) );
  XNOR U34959 ( .A(n34941), .B(n35314), .Z(n35316) );
  XOR U34960 ( .A(n35322), .B(n35323), .Z(n34941) );
  AND U34961 ( .A(n573), .B(n35324), .Z(n35323) );
  XOR U34962 ( .A(n35325), .B(n35322), .Z(n35324) );
  XOR U34963 ( .A(n35326), .B(n35327), .Z(n35314) );
  AND U34964 ( .A(n35328), .B(n35329), .Z(n35327) );
  XOR U34965 ( .A(n35326), .B(n34956), .Z(n35329) );
  XOR U34966 ( .A(n35330), .B(n35331), .Z(n34956) );
  AND U34967 ( .A(n575), .B(n35332), .Z(n35331) );
  XOR U34968 ( .A(n35333), .B(n35330), .Z(n35332) );
  XNOR U34969 ( .A(n34953), .B(n35326), .Z(n35328) );
  XOR U34970 ( .A(n35334), .B(n35335), .Z(n34953) );
  AND U34971 ( .A(n573), .B(n35336), .Z(n35335) );
  XOR U34972 ( .A(n35337), .B(n35334), .Z(n35336) );
  XOR U34973 ( .A(n35338), .B(n35339), .Z(n35326) );
  AND U34974 ( .A(n35340), .B(n35341), .Z(n35339) );
  XOR U34975 ( .A(n35338), .B(n34968), .Z(n35341) );
  XOR U34976 ( .A(n35342), .B(n35343), .Z(n34968) );
  AND U34977 ( .A(n575), .B(n35344), .Z(n35343) );
  XOR U34978 ( .A(n35345), .B(n35342), .Z(n35344) );
  XNOR U34979 ( .A(n34965), .B(n35338), .Z(n35340) );
  XOR U34980 ( .A(n35346), .B(n35347), .Z(n34965) );
  AND U34981 ( .A(n573), .B(n35348), .Z(n35347) );
  XOR U34982 ( .A(n35349), .B(n35346), .Z(n35348) );
  XOR U34983 ( .A(n35350), .B(n35351), .Z(n35338) );
  AND U34984 ( .A(n35352), .B(n35353), .Z(n35351) );
  XOR U34985 ( .A(n35350), .B(n34980), .Z(n35353) );
  XOR U34986 ( .A(n35354), .B(n35355), .Z(n34980) );
  AND U34987 ( .A(n575), .B(n35356), .Z(n35355) );
  XOR U34988 ( .A(n35357), .B(n35354), .Z(n35356) );
  XNOR U34989 ( .A(n34977), .B(n35350), .Z(n35352) );
  XOR U34990 ( .A(n35358), .B(n35359), .Z(n34977) );
  AND U34991 ( .A(n573), .B(n35360), .Z(n35359) );
  XOR U34992 ( .A(n35361), .B(n35358), .Z(n35360) );
  XOR U34993 ( .A(n35362), .B(n35363), .Z(n35350) );
  AND U34994 ( .A(n35364), .B(n35365), .Z(n35363) );
  XOR U34995 ( .A(n35362), .B(n34992), .Z(n35365) );
  XOR U34996 ( .A(n35366), .B(n35367), .Z(n34992) );
  AND U34997 ( .A(n575), .B(n35368), .Z(n35367) );
  XOR U34998 ( .A(n35369), .B(n35366), .Z(n35368) );
  XNOR U34999 ( .A(n34989), .B(n35362), .Z(n35364) );
  XOR U35000 ( .A(n35370), .B(n35371), .Z(n34989) );
  AND U35001 ( .A(n573), .B(n35372), .Z(n35371) );
  XOR U35002 ( .A(n35373), .B(n35370), .Z(n35372) );
  XOR U35003 ( .A(n35374), .B(n35375), .Z(n35362) );
  AND U35004 ( .A(n35376), .B(n35377), .Z(n35375) );
  XOR U35005 ( .A(n35374), .B(n35004), .Z(n35377) );
  XOR U35006 ( .A(n35378), .B(n35379), .Z(n35004) );
  AND U35007 ( .A(n575), .B(n35380), .Z(n35379) );
  XOR U35008 ( .A(n35381), .B(n35378), .Z(n35380) );
  XNOR U35009 ( .A(n35001), .B(n35374), .Z(n35376) );
  XOR U35010 ( .A(n35382), .B(n35383), .Z(n35001) );
  AND U35011 ( .A(n573), .B(n35384), .Z(n35383) );
  XOR U35012 ( .A(n35385), .B(n35382), .Z(n35384) );
  XOR U35013 ( .A(n35386), .B(n35387), .Z(n35374) );
  AND U35014 ( .A(n35388), .B(n35389), .Z(n35387) );
  XOR U35015 ( .A(n35386), .B(n35016), .Z(n35389) );
  XOR U35016 ( .A(n35390), .B(n35391), .Z(n35016) );
  AND U35017 ( .A(n575), .B(n35392), .Z(n35391) );
  XOR U35018 ( .A(n35393), .B(n35390), .Z(n35392) );
  XNOR U35019 ( .A(n35013), .B(n35386), .Z(n35388) );
  XOR U35020 ( .A(n35394), .B(n35395), .Z(n35013) );
  AND U35021 ( .A(n573), .B(n35396), .Z(n35395) );
  XOR U35022 ( .A(n35397), .B(n35394), .Z(n35396) );
  XOR U35023 ( .A(n35398), .B(n35399), .Z(n35386) );
  AND U35024 ( .A(n35400), .B(n35401), .Z(n35399) );
  XOR U35025 ( .A(n35398), .B(n35028), .Z(n35401) );
  XOR U35026 ( .A(n35402), .B(n35403), .Z(n35028) );
  AND U35027 ( .A(n575), .B(n35404), .Z(n35403) );
  XOR U35028 ( .A(n35405), .B(n35402), .Z(n35404) );
  XNOR U35029 ( .A(n35025), .B(n35398), .Z(n35400) );
  XOR U35030 ( .A(n35406), .B(n35407), .Z(n35025) );
  AND U35031 ( .A(n573), .B(n35408), .Z(n35407) );
  XOR U35032 ( .A(n35409), .B(n35406), .Z(n35408) );
  XOR U35033 ( .A(n35410), .B(n35411), .Z(n35398) );
  AND U35034 ( .A(n35412), .B(n35413), .Z(n35411) );
  XOR U35035 ( .A(n35410), .B(n35040), .Z(n35413) );
  XOR U35036 ( .A(n35414), .B(n35415), .Z(n35040) );
  AND U35037 ( .A(n575), .B(n35416), .Z(n35415) );
  XOR U35038 ( .A(n35417), .B(n35414), .Z(n35416) );
  XNOR U35039 ( .A(n35037), .B(n35410), .Z(n35412) );
  XOR U35040 ( .A(n35418), .B(n35419), .Z(n35037) );
  AND U35041 ( .A(n573), .B(n35420), .Z(n35419) );
  XOR U35042 ( .A(n35421), .B(n35418), .Z(n35420) );
  XOR U35043 ( .A(n35422), .B(n35423), .Z(n35410) );
  AND U35044 ( .A(n35424), .B(n35425), .Z(n35423) );
  XOR U35045 ( .A(n35422), .B(n35052), .Z(n35425) );
  XOR U35046 ( .A(n35426), .B(n35427), .Z(n35052) );
  AND U35047 ( .A(n575), .B(n35428), .Z(n35427) );
  XOR U35048 ( .A(n35429), .B(n35426), .Z(n35428) );
  XNOR U35049 ( .A(n35049), .B(n35422), .Z(n35424) );
  XOR U35050 ( .A(n35430), .B(n35431), .Z(n35049) );
  AND U35051 ( .A(n573), .B(n35432), .Z(n35431) );
  XOR U35052 ( .A(n35433), .B(n35430), .Z(n35432) );
  XOR U35053 ( .A(n35434), .B(n35435), .Z(n35422) );
  AND U35054 ( .A(n35436), .B(n35437), .Z(n35435) );
  XNOR U35055 ( .A(n35438), .B(n35065), .Z(n35437) );
  XOR U35056 ( .A(n35439), .B(n35440), .Z(n35065) );
  AND U35057 ( .A(n575), .B(n35441), .Z(n35440) );
  XOR U35058 ( .A(n35439), .B(n35442), .Z(n35441) );
  XNOR U35059 ( .A(n35062), .B(n35434), .Z(n35436) );
  XOR U35060 ( .A(n35443), .B(n35444), .Z(n35062) );
  AND U35061 ( .A(n573), .B(n35445), .Z(n35444) );
  XOR U35062 ( .A(n35443), .B(n35446), .Z(n35445) );
  IV U35063 ( .A(n35438), .Z(n35434) );
  AND U35064 ( .A(n35070), .B(n35073), .Z(n35438) );
  XNOR U35065 ( .A(n35447), .B(n35448), .Z(n35073) );
  AND U35066 ( .A(n575), .B(n35449), .Z(n35448) );
  XNOR U35067 ( .A(n35450), .B(n35447), .Z(n35449) );
  XOR U35068 ( .A(n35451), .B(n35452), .Z(n575) );
  AND U35069 ( .A(n35453), .B(n35454), .Z(n35452) );
  XOR U35070 ( .A(n35081), .B(n35451), .Z(n35454) );
  IV U35071 ( .A(n35455), .Z(n35081) );
  AND U35072 ( .A(p_input[3583]), .B(p_input[3551]), .Z(n35455) );
  XOR U35073 ( .A(n35451), .B(n35078), .Z(n35453) );
  AND U35074 ( .A(p_input[3487]), .B(p_input[3519]), .Z(n35078) );
  XOR U35075 ( .A(n35456), .B(n35457), .Z(n35451) );
  AND U35076 ( .A(n35458), .B(n35459), .Z(n35457) );
  XOR U35077 ( .A(n35456), .B(n35093), .Z(n35459) );
  XNOR U35078 ( .A(p_input[3550]), .B(n35460), .Z(n35093) );
  AND U35079 ( .A(n719), .B(n35461), .Z(n35460) );
  XOR U35080 ( .A(p_input[3582]), .B(p_input[3550]), .Z(n35461) );
  XNOR U35081 ( .A(n35090), .B(n35456), .Z(n35458) );
  XOR U35082 ( .A(n35462), .B(n35463), .Z(n35090) );
  AND U35083 ( .A(n717), .B(n35464), .Z(n35463) );
  XOR U35084 ( .A(p_input[3518]), .B(p_input[3486]), .Z(n35464) );
  XOR U35085 ( .A(n35465), .B(n35466), .Z(n35456) );
  AND U35086 ( .A(n35467), .B(n35468), .Z(n35466) );
  XOR U35087 ( .A(n35465), .B(n35105), .Z(n35468) );
  XNOR U35088 ( .A(p_input[3549]), .B(n35469), .Z(n35105) );
  AND U35089 ( .A(n719), .B(n35470), .Z(n35469) );
  XOR U35090 ( .A(p_input[3581]), .B(p_input[3549]), .Z(n35470) );
  XNOR U35091 ( .A(n35102), .B(n35465), .Z(n35467) );
  XOR U35092 ( .A(n35471), .B(n35472), .Z(n35102) );
  AND U35093 ( .A(n717), .B(n35473), .Z(n35472) );
  XOR U35094 ( .A(p_input[3517]), .B(p_input[3485]), .Z(n35473) );
  XOR U35095 ( .A(n35474), .B(n35475), .Z(n35465) );
  AND U35096 ( .A(n35476), .B(n35477), .Z(n35475) );
  XOR U35097 ( .A(n35474), .B(n35117), .Z(n35477) );
  XNOR U35098 ( .A(p_input[3548]), .B(n35478), .Z(n35117) );
  AND U35099 ( .A(n719), .B(n35479), .Z(n35478) );
  XOR U35100 ( .A(p_input[3580]), .B(p_input[3548]), .Z(n35479) );
  XNOR U35101 ( .A(n35114), .B(n35474), .Z(n35476) );
  XOR U35102 ( .A(n35480), .B(n35481), .Z(n35114) );
  AND U35103 ( .A(n717), .B(n35482), .Z(n35481) );
  XOR U35104 ( .A(p_input[3516]), .B(p_input[3484]), .Z(n35482) );
  XOR U35105 ( .A(n35483), .B(n35484), .Z(n35474) );
  AND U35106 ( .A(n35485), .B(n35486), .Z(n35484) );
  XOR U35107 ( .A(n35483), .B(n35129), .Z(n35486) );
  XNOR U35108 ( .A(p_input[3547]), .B(n35487), .Z(n35129) );
  AND U35109 ( .A(n719), .B(n35488), .Z(n35487) );
  XOR U35110 ( .A(p_input[3579]), .B(p_input[3547]), .Z(n35488) );
  XNOR U35111 ( .A(n35126), .B(n35483), .Z(n35485) );
  XOR U35112 ( .A(n35489), .B(n35490), .Z(n35126) );
  AND U35113 ( .A(n717), .B(n35491), .Z(n35490) );
  XOR U35114 ( .A(p_input[3515]), .B(p_input[3483]), .Z(n35491) );
  XOR U35115 ( .A(n35492), .B(n35493), .Z(n35483) );
  AND U35116 ( .A(n35494), .B(n35495), .Z(n35493) );
  XOR U35117 ( .A(n35492), .B(n35141), .Z(n35495) );
  XNOR U35118 ( .A(p_input[3546]), .B(n35496), .Z(n35141) );
  AND U35119 ( .A(n719), .B(n35497), .Z(n35496) );
  XOR U35120 ( .A(p_input[3578]), .B(p_input[3546]), .Z(n35497) );
  XNOR U35121 ( .A(n35138), .B(n35492), .Z(n35494) );
  XOR U35122 ( .A(n35498), .B(n35499), .Z(n35138) );
  AND U35123 ( .A(n717), .B(n35500), .Z(n35499) );
  XOR U35124 ( .A(p_input[3514]), .B(p_input[3482]), .Z(n35500) );
  XOR U35125 ( .A(n35501), .B(n35502), .Z(n35492) );
  AND U35126 ( .A(n35503), .B(n35504), .Z(n35502) );
  XOR U35127 ( .A(n35501), .B(n35153), .Z(n35504) );
  XNOR U35128 ( .A(p_input[3545]), .B(n35505), .Z(n35153) );
  AND U35129 ( .A(n719), .B(n35506), .Z(n35505) );
  XOR U35130 ( .A(p_input[3577]), .B(p_input[3545]), .Z(n35506) );
  XNOR U35131 ( .A(n35150), .B(n35501), .Z(n35503) );
  XOR U35132 ( .A(n35507), .B(n35508), .Z(n35150) );
  AND U35133 ( .A(n717), .B(n35509), .Z(n35508) );
  XOR U35134 ( .A(p_input[3513]), .B(p_input[3481]), .Z(n35509) );
  XOR U35135 ( .A(n35510), .B(n35511), .Z(n35501) );
  AND U35136 ( .A(n35512), .B(n35513), .Z(n35511) );
  XOR U35137 ( .A(n35510), .B(n35165), .Z(n35513) );
  XNOR U35138 ( .A(p_input[3544]), .B(n35514), .Z(n35165) );
  AND U35139 ( .A(n719), .B(n35515), .Z(n35514) );
  XOR U35140 ( .A(p_input[3576]), .B(p_input[3544]), .Z(n35515) );
  XNOR U35141 ( .A(n35162), .B(n35510), .Z(n35512) );
  XOR U35142 ( .A(n35516), .B(n35517), .Z(n35162) );
  AND U35143 ( .A(n717), .B(n35518), .Z(n35517) );
  XOR U35144 ( .A(p_input[3512]), .B(p_input[3480]), .Z(n35518) );
  XOR U35145 ( .A(n35519), .B(n35520), .Z(n35510) );
  AND U35146 ( .A(n35521), .B(n35522), .Z(n35520) );
  XOR U35147 ( .A(n35519), .B(n35177), .Z(n35522) );
  XNOR U35148 ( .A(p_input[3543]), .B(n35523), .Z(n35177) );
  AND U35149 ( .A(n719), .B(n35524), .Z(n35523) );
  XOR U35150 ( .A(p_input[3575]), .B(p_input[3543]), .Z(n35524) );
  XNOR U35151 ( .A(n35174), .B(n35519), .Z(n35521) );
  XOR U35152 ( .A(n35525), .B(n35526), .Z(n35174) );
  AND U35153 ( .A(n717), .B(n35527), .Z(n35526) );
  XOR U35154 ( .A(p_input[3511]), .B(p_input[3479]), .Z(n35527) );
  XOR U35155 ( .A(n35528), .B(n35529), .Z(n35519) );
  AND U35156 ( .A(n35530), .B(n35531), .Z(n35529) );
  XOR U35157 ( .A(n35528), .B(n35189), .Z(n35531) );
  XNOR U35158 ( .A(p_input[3542]), .B(n35532), .Z(n35189) );
  AND U35159 ( .A(n719), .B(n35533), .Z(n35532) );
  XOR U35160 ( .A(p_input[3574]), .B(p_input[3542]), .Z(n35533) );
  XNOR U35161 ( .A(n35186), .B(n35528), .Z(n35530) );
  XOR U35162 ( .A(n35534), .B(n35535), .Z(n35186) );
  AND U35163 ( .A(n717), .B(n35536), .Z(n35535) );
  XOR U35164 ( .A(p_input[3510]), .B(p_input[3478]), .Z(n35536) );
  XOR U35165 ( .A(n35537), .B(n35538), .Z(n35528) );
  AND U35166 ( .A(n35539), .B(n35540), .Z(n35538) );
  XOR U35167 ( .A(n35537), .B(n35201), .Z(n35540) );
  XNOR U35168 ( .A(p_input[3541]), .B(n35541), .Z(n35201) );
  AND U35169 ( .A(n719), .B(n35542), .Z(n35541) );
  XOR U35170 ( .A(p_input[3573]), .B(p_input[3541]), .Z(n35542) );
  XNOR U35171 ( .A(n35198), .B(n35537), .Z(n35539) );
  XOR U35172 ( .A(n35543), .B(n35544), .Z(n35198) );
  AND U35173 ( .A(n717), .B(n35545), .Z(n35544) );
  XOR U35174 ( .A(p_input[3509]), .B(p_input[3477]), .Z(n35545) );
  XOR U35175 ( .A(n35546), .B(n35547), .Z(n35537) );
  AND U35176 ( .A(n35548), .B(n35549), .Z(n35547) );
  XOR U35177 ( .A(n35546), .B(n35213), .Z(n35549) );
  XNOR U35178 ( .A(p_input[3540]), .B(n35550), .Z(n35213) );
  AND U35179 ( .A(n719), .B(n35551), .Z(n35550) );
  XOR U35180 ( .A(p_input[3572]), .B(p_input[3540]), .Z(n35551) );
  XNOR U35181 ( .A(n35210), .B(n35546), .Z(n35548) );
  XOR U35182 ( .A(n35552), .B(n35553), .Z(n35210) );
  AND U35183 ( .A(n717), .B(n35554), .Z(n35553) );
  XOR U35184 ( .A(p_input[3508]), .B(p_input[3476]), .Z(n35554) );
  XOR U35185 ( .A(n35555), .B(n35556), .Z(n35546) );
  AND U35186 ( .A(n35557), .B(n35558), .Z(n35556) );
  XOR U35187 ( .A(n35555), .B(n35225), .Z(n35558) );
  XNOR U35188 ( .A(p_input[3539]), .B(n35559), .Z(n35225) );
  AND U35189 ( .A(n719), .B(n35560), .Z(n35559) );
  XOR U35190 ( .A(p_input[3571]), .B(p_input[3539]), .Z(n35560) );
  XNOR U35191 ( .A(n35222), .B(n35555), .Z(n35557) );
  XOR U35192 ( .A(n35561), .B(n35562), .Z(n35222) );
  AND U35193 ( .A(n717), .B(n35563), .Z(n35562) );
  XOR U35194 ( .A(p_input[3507]), .B(p_input[3475]), .Z(n35563) );
  XOR U35195 ( .A(n35564), .B(n35565), .Z(n35555) );
  AND U35196 ( .A(n35566), .B(n35567), .Z(n35565) );
  XOR U35197 ( .A(n35564), .B(n35237), .Z(n35567) );
  XNOR U35198 ( .A(p_input[3538]), .B(n35568), .Z(n35237) );
  AND U35199 ( .A(n719), .B(n35569), .Z(n35568) );
  XOR U35200 ( .A(p_input[3570]), .B(p_input[3538]), .Z(n35569) );
  XNOR U35201 ( .A(n35234), .B(n35564), .Z(n35566) );
  XOR U35202 ( .A(n35570), .B(n35571), .Z(n35234) );
  AND U35203 ( .A(n717), .B(n35572), .Z(n35571) );
  XOR U35204 ( .A(p_input[3506]), .B(p_input[3474]), .Z(n35572) );
  XOR U35205 ( .A(n35573), .B(n35574), .Z(n35564) );
  AND U35206 ( .A(n35575), .B(n35576), .Z(n35574) );
  XOR U35207 ( .A(n35573), .B(n35249), .Z(n35576) );
  XNOR U35208 ( .A(p_input[3537]), .B(n35577), .Z(n35249) );
  AND U35209 ( .A(n719), .B(n35578), .Z(n35577) );
  XOR U35210 ( .A(p_input[3569]), .B(p_input[3537]), .Z(n35578) );
  XNOR U35211 ( .A(n35246), .B(n35573), .Z(n35575) );
  XOR U35212 ( .A(n35579), .B(n35580), .Z(n35246) );
  AND U35213 ( .A(n717), .B(n35581), .Z(n35580) );
  XOR U35214 ( .A(p_input[3505]), .B(p_input[3473]), .Z(n35581) );
  XOR U35215 ( .A(n35582), .B(n35583), .Z(n35573) );
  AND U35216 ( .A(n35584), .B(n35585), .Z(n35583) );
  XOR U35217 ( .A(n35582), .B(n35261), .Z(n35585) );
  XNOR U35218 ( .A(p_input[3536]), .B(n35586), .Z(n35261) );
  AND U35219 ( .A(n719), .B(n35587), .Z(n35586) );
  XOR U35220 ( .A(p_input[3568]), .B(p_input[3536]), .Z(n35587) );
  XNOR U35221 ( .A(n35258), .B(n35582), .Z(n35584) );
  XOR U35222 ( .A(n35588), .B(n35589), .Z(n35258) );
  AND U35223 ( .A(n717), .B(n35590), .Z(n35589) );
  XOR U35224 ( .A(p_input[3504]), .B(p_input[3472]), .Z(n35590) );
  XOR U35225 ( .A(n35591), .B(n35592), .Z(n35582) );
  AND U35226 ( .A(n35593), .B(n35594), .Z(n35592) );
  XOR U35227 ( .A(n35591), .B(n35273), .Z(n35594) );
  XNOR U35228 ( .A(p_input[3535]), .B(n35595), .Z(n35273) );
  AND U35229 ( .A(n719), .B(n35596), .Z(n35595) );
  XOR U35230 ( .A(p_input[3567]), .B(p_input[3535]), .Z(n35596) );
  XNOR U35231 ( .A(n35270), .B(n35591), .Z(n35593) );
  XOR U35232 ( .A(n35597), .B(n35598), .Z(n35270) );
  AND U35233 ( .A(n717), .B(n35599), .Z(n35598) );
  XOR U35234 ( .A(p_input[3503]), .B(p_input[3471]), .Z(n35599) );
  XOR U35235 ( .A(n35600), .B(n35601), .Z(n35591) );
  AND U35236 ( .A(n35602), .B(n35603), .Z(n35601) );
  XOR U35237 ( .A(n35600), .B(n35285), .Z(n35603) );
  XNOR U35238 ( .A(p_input[3534]), .B(n35604), .Z(n35285) );
  AND U35239 ( .A(n719), .B(n35605), .Z(n35604) );
  XOR U35240 ( .A(p_input[3566]), .B(p_input[3534]), .Z(n35605) );
  XNOR U35241 ( .A(n35282), .B(n35600), .Z(n35602) );
  XOR U35242 ( .A(n35606), .B(n35607), .Z(n35282) );
  AND U35243 ( .A(n717), .B(n35608), .Z(n35607) );
  XOR U35244 ( .A(p_input[3502]), .B(p_input[3470]), .Z(n35608) );
  XOR U35245 ( .A(n35609), .B(n35610), .Z(n35600) );
  AND U35246 ( .A(n35611), .B(n35612), .Z(n35610) );
  XOR U35247 ( .A(n35609), .B(n35297), .Z(n35612) );
  XNOR U35248 ( .A(p_input[3533]), .B(n35613), .Z(n35297) );
  AND U35249 ( .A(n719), .B(n35614), .Z(n35613) );
  XOR U35250 ( .A(p_input[3565]), .B(p_input[3533]), .Z(n35614) );
  XNOR U35251 ( .A(n35294), .B(n35609), .Z(n35611) );
  XOR U35252 ( .A(n35615), .B(n35616), .Z(n35294) );
  AND U35253 ( .A(n717), .B(n35617), .Z(n35616) );
  XOR U35254 ( .A(p_input[3501]), .B(p_input[3469]), .Z(n35617) );
  XOR U35255 ( .A(n35618), .B(n35619), .Z(n35609) );
  AND U35256 ( .A(n35620), .B(n35621), .Z(n35619) );
  XOR U35257 ( .A(n35618), .B(n35309), .Z(n35621) );
  XNOR U35258 ( .A(p_input[3532]), .B(n35622), .Z(n35309) );
  AND U35259 ( .A(n719), .B(n35623), .Z(n35622) );
  XOR U35260 ( .A(p_input[3564]), .B(p_input[3532]), .Z(n35623) );
  XNOR U35261 ( .A(n35306), .B(n35618), .Z(n35620) );
  XOR U35262 ( .A(n35624), .B(n35625), .Z(n35306) );
  AND U35263 ( .A(n717), .B(n35626), .Z(n35625) );
  XOR U35264 ( .A(p_input[3500]), .B(p_input[3468]), .Z(n35626) );
  XOR U35265 ( .A(n35627), .B(n35628), .Z(n35618) );
  AND U35266 ( .A(n35629), .B(n35630), .Z(n35628) );
  XOR U35267 ( .A(n35627), .B(n35321), .Z(n35630) );
  XNOR U35268 ( .A(p_input[3531]), .B(n35631), .Z(n35321) );
  AND U35269 ( .A(n719), .B(n35632), .Z(n35631) );
  XOR U35270 ( .A(p_input[3563]), .B(p_input[3531]), .Z(n35632) );
  XNOR U35271 ( .A(n35318), .B(n35627), .Z(n35629) );
  XOR U35272 ( .A(n35633), .B(n35634), .Z(n35318) );
  AND U35273 ( .A(n717), .B(n35635), .Z(n35634) );
  XOR U35274 ( .A(p_input[3499]), .B(p_input[3467]), .Z(n35635) );
  XOR U35275 ( .A(n35636), .B(n35637), .Z(n35627) );
  AND U35276 ( .A(n35638), .B(n35639), .Z(n35637) );
  XOR U35277 ( .A(n35636), .B(n35333), .Z(n35639) );
  XNOR U35278 ( .A(p_input[3530]), .B(n35640), .Z(n35333) );
  AND U35279 ( .A(n719), .B(n35641), .Z(n35640) );
  XOR U35280 ( .A(p_input[3562]), .B(p_input[3530]), .Z(n35641) );
  XNOR U35281 ( .A(n35330), .B(n35636), .Z(n35638) );
  XOR U35282 ( .A(n35642), .B(n35643), .Z(n35330) );
  AND U35283 ( .A(n717), .B(n35644), .Z(n35643) );
  XOR U35284 ( .A(p_input[3498]), .B(p_input[3466]), .Z(n35644) );
  XOR U35285 ( .A(n35645), .B(n35646), .Z(n35636) );
  AND U35286 ( .A(n35647), .B(n35648), .Z(n35646) );
  XOR U35287 ( .A(n35645), .B(n35345), .Z(n35648) );
  XNOR U35288 ( .A(p_input[3529]), .B(n35649), .Z(n35345) );
  AND U35289 ( .A(n719), .B(n35650), .Z(n35649) );
  XOR U35290 ( .A(p_input[3561]), .B(p_input[3529]), .Z(n35650) );
  XNOR U35291 ( .A(n35342), .B(n35645), .Z(n35647) );
  XOR U35292 ( .A(n35651), .B(n35652), .Z(n35342) );
  AND U35293 ( .A(n717), .B(n35653), .Z(n35652) );
  XOR U35294 ( .A(p_input[3497]), .B(p_input[3465]), .Z(n35653) );
  XOR U35295 ( .A(n35654), .B(n35655), .Z(n35645) );
  AND U35296 ( .A(n35656), .B(n35657), .Z(n35655) );
  XOR U35297 ( .A(n35654), .B(n35357), .Z(n35657) );
  XNOR U35298 ( .A(p_input[3528]), .B(n35658), .Z(n35357) );
  AND U35299 ( .A(n719), .B(n35659), .Z(n35658) );
  XOR U35300 ( .A(p_input[3560]), .B(p_input[3528]), .Z(n35659) );
  XNOR U35301 ( .A(n35354), .B(n35654), .Z(n35656) );
  XOR U35302 ( .A(n35660), .B(n35661), .Z(n35354) );
  AND U35303 ( .A(n717), .B(n35662), .Z(n35661) );
  XOR U35304 ( .A(p_input[3496]), .B(p_input[3464]), .Z(n35662) );
  XOR U35305 ( .A(n35663), .B(n35664), .Z(n35654) );
  AND U35306 ( .A(n35665), .B(n35666), .Z(n35664) );
  XOR U35307 ( .A(n35663), .B(n35369), .Z(n35666) );
  XNOR U35308 ( .A(p_input[3527]), .B(n35667), .Z(n35369) );
  AND U35309 ( .A(n719), .B(n35668), .Z(n35667) );
  XOR U35310 ( .A(p_input[3559]), .B(p_input[3527]), .Z(n35668) );
  XNOR U35311 ( .A(n35366), .B(n35663), .Z(n35665) );
  XOR U35312 ( .A(n35669), .B(n35670), .Z(n35366) );
  AND U35313 ( .A(n717), .B(n35671), .Z(n35670) );
  XOR U35314 ( .A(p_input[3495]), .B(p_input[3463]), .Z(n35671) );
  XOR U35315 ( .A(n35672), .B(n35673), .Z(n35663) );
  AND U35316 ( .A(n35674), .B(n35675), .Z(n35673) );
  XOR U35317 ( .A(n35672), .B(n35381), .Z(n35675) );
  XNOR U35318 ( .A(p_input[3526]), .B(n35676), .Z(n35381) );
  AND U35319 ( .A(n719), .B(n35677), .Z(n35676) );
  XOR U35320 ( .A(p_input[3558]), .B(p_input[3526]), .Z(n35677) );
  XNOR U35321 ( .A(n35378), .B(n35672), .Z(n35674) );
  XOR U35322 ( .A(n35678), .B(n35679), .Z(n35378) );
  AND U35323 ( .A(n717), .B(n35680), .Z(n35679) );
  XOR U35324 ( .A(p_input[3494]), .B(p_input[3462]), .Z(n35680) );
  XOR U35325 ( .A(n35681), .B(n35682), .Z(n35672) );
  AND U35326 ( .A(n35683), .B(n35684), .Z(n35682) );
  XOR U35327 ( .A(n35681), .B(n35393), .Z(n35684) );
  XNOR U35328 ( .A(p_input[3525]), .B(n35685), .Z(n35393) );
  AND U35329 ( .A(n719), .B(n35686), .Z(n35685) );
  XOR U35330 ( .A(p_input[3557]), .B(p_input[3525]), .Z(n35686) );
  XNOR U35331 ( .A(n35390), .B(n35681), .Z(n35683) );
  XOR U35332 ( .A(n35687), .B(n35688), .Z(n35390) );
  AND U35333 ( .A(n717), .B(n35689), .Z(n35688) );
  XOR U35334 ( .A(p_input[3493]), .B(p_input[3461]), .Z(n35689) );
  XOR U35335 ( .A(n35690), .B(n35691), .Z(n35681) );
  AND U35336 ( .A(n35692), .B(n35693), .Z(n35691) );
  XOR U35337 ( .A(n35690), .B(n35405), .Z(n35693) );
  XNOR U35338 ( .A(p_input[3524]), .B(n35694), .Z(n35405) );
  AND U35339 ( .A(n719), .B(n35695), .Z(n35694) );
  XOR U35340 ( .A(p_input[3556]), .B(p_input[3524]), .Z(n35695) );
  XNOR U35341 ( .A(n35402), .B(n35690), .Z(n35692) );
  XOR U35342 ( .A(n35696), .B(n35697), .Z(n35402) );
  AND U35343 ( .A(n717), .B(n35698), .Z(n35697) );
  XOR U35344 ( .A(p_input[3492]), .B(p_input[3460]), .Z(n35698) );
  XOR U35345 ( .A(n35699), .B(n35700), .Z(n35690) );
  AND U35346 ( .A(n35701), .B(n35702), .Z(n35700) );
  XOR U35347 ( .A(n35699), .B(n35417), .Z(n35702) );
  XNOR U35348 ( .A(p_input[3523]), .B(n35703), .Z(n35417) );
  AND U35349 ( .A(n719), .B(n35704), .Z(n35703) );
  XOR U35350 ( .A(p_input[3555]), .B(p_input[3523]), .Z(n35704) );
  XNOR U35351 ( .A(n35414), .B(n35699), .Z(n35701) );
  XOR U35352 ( .A(n35705), .B(n35706), .Z(n35414) );
  AND U35353 ( .A(n717), .B(n35707), .Z(n35706) );
  XOR U35354 ( .A(p_input[3491]), .B(p_input[3459]), .Z(n35707) );
  XOR U35355 ( .A(n35708), .B(n35709), .Z(n35699) );
  AND U35356 ( .A(n35710), .B(n35711), .Z(n35709) );
  XOR U35357 ( .A(n35708), .B(n35429), .Z(n35711) );
  XNOR U35358 ( .A(p_input[3522]), .B(n35712), .Z(n35429) );
  AND U35359 ( .A(n719), .B(n35713), .Z(n35712) );
  XOR U35360 ( .A(p_input[3554]), .B(p_input[3522]), .Z(n35713) );
  XNOR U35361 ( .A(n35426), .B(n35708), .Z(n35710) );
  XOR U35362 ( .A(n35714), .B(n35715), .Z(n35426) );
  AND U35363 ( .A(n717), .B(n35716), .Z(n35715) );
  XOR U35364 ( .A(p_input[3490]), .B(p_input[3458]), .Z(n35716) );
  XOR U35365 ( .A(n35717), .B(n35718), .Z(n35708) );
  AND U35366 ( .A(n35719), .B(n35720), .Z(n35718) );
  XNOR U35367 ( .A(n35721), .B(n35442), .Z(n35720) );
  XNOR U35368 ( .A(p_input[3521]), .B(n35722), .Z(n35442) );
  AND U35369 ( .A(n719), .B(n35723), .Z(n35722) );
  XNOR U35370 ( .A(p_input[3553]), .B(n35724), .Z(n35723) );
  IV U35371 ( .A(p_input[3521]), .Z(n35724) );
  XNOR U35372 ( .A(n35439), .B(n35717), .Z(n35719) );
  XNOR U35373 ( .A(p_input[3457]), .B(n35725), .Z(n35439) );
  AND U35374 ( .A(n717), .B(n35726), .Z(n35725) );
  XOR U35375 ( .A(p_input[3489]), .B(p_input[3457]), .Z(n35726) );
  IV U35376 ( .A(n35721), .Z(n35717) );
  AND U35377 ( .A(n35447), .B(n35450), .Z(n35721) );
  XOR U35378 ( .A(p_input[3520]), .B(n35727), .Z(n35450) );
  AND U35379 ( .A(n719), .B(n35728), .Z(n35727) );
  XOR U35380 ( .A(p_input[3552]), .B(p_input[3520]), .Z(n35728) );
  XOR U35381 ( .A(n35729), .B(n35730), .Z(n719) );
  AND U35382 ( .A(n35731), .B(n35732), .Z(n35730) );
  XNOR U35383 ( .A(p_input[3583]), .B(n35729), .Z(n35732) );
  XOR U35384 ( .A(n35729), .B(p_input[3551]), .Z(n35731) );
  XOR U35385 ( .A(n35733), .B(n35734), .Z(n35729) );
  AND U35386 ( .A(n35735), .B(n35736), .Z(n35734) );
  XNOR U35387 ( .A(p_input[3582]), .B(n35733), .Z(n35736) );
  XOR U35388 ( .A(n35733), .B(p_input[3550]), .Z(n35735) );
  XOR U35389 ( .A(n35737), .B(n35738), .Z(n35733) );
  AND U35390 ( .A(n35739), .B(n35740), .Z(n35738) );
  XNOR U35391 ( .A(p_input[3581]), .B(n35737), .Z(n35740) );
  XOR U35392 ( .A(n35737), .B(p_input[3549]), .Z(n35739) );
  XOR U35393 ( .A(n35741), .B(n35742), .Z(n35737) );
  AND U35394 ( .A(n35743), .B(n35744), .Z(n35742) );
  XNOR U35395 ( .A(p_input[3580]), .B(n35741), .Z(n35744) );
  XOR U35396 ( .A(n35741), .B(p_input[3548]), .Z(n35743) );
  XOR U35397 ( .A(n35745), .B(n35746), .Z(n35741) );
  AND U35398 ( .A(n35747), .B(n35748), .Z(n35746) );
  XNOR U35399 ( .A(p_input[3579]), .B(n35745), .Z(n35748) );
  XOR U35400 ( .A(n35745), .B(p_input[3547]), .Z(n35747) );
  XOR U35401 ( .A(n35749), .B(n35750), .Z(n35745) );
  AND U35402 ( .A(n35751), .B(n35752), .Z(n35750) );
  XNOR U35403 ( .A(p_input[3578]), .B(n35749), .Z(n35752) );
  XOR U35404 ( .A(n35749), .B(p_input[3546]), .Z(n35751) );
  XOR U35405 ( .A(n35753), .B(n35754), .Z(n35749) );
  AND U35406 ( .A(n35755), .B(n35756), .Z(n35754) );
  XNOR U35407 ( .A(p_input[3577]), .B(n35753), .Z(n35756) );
  XOR U35408 ( .A(n35753), .B(p_input[3545]), .Z(n35755) );
  XOR U35409 ( .A(n35757), .B(n35758), .Z(n35753) );
  AND U35410 ( .A(n35759), .B(n35760), .Z(n35758) );
  XNOR U35411 ( .A(p_input[3576]), .B(n35757), .Z(n35760) );
  XOR U35412 ( .A(n35757), .B(p_input[3544]), .Z(n35759) );
  XOR U35413 ( .A(n35761), .B(n35762), .Z(n35757) );
  AND U35414 ( .A(n35763), .B(n35764), .Z(n35762) );
  XNOR U35415 ( .A(p_input[3575]), .B(n35761), .Z(n35764) );
  XOR U35416 ( .A(n35761), .B(p_input[3543]), .Z(n35763) );
  XOR U35417 ( .A(n35765), .B(n35766), .Z(n35761) );
  AND U35418 ( .A(n35767), .B(n35768), .Z(n35766) );
  XNOR U35419 ( .A(p_input[3574]), .B(n35765), .Z(n35768) );
  XOR U35420 ( .A(n35765), .B(p_input[3542]), .Z(n35767) );
  XOR U35421 ( .A(n35769), .B(n35770), .Z(n35765) );
  AND U35422 ( .A(n35771), .B(n35772), .Z(n35770) );
  XNOR U35423 ( .A(p_input[3573]), .B(n35769), .Z(n35772) );
  XOR U35424 ( .A(n35769), .B(p_input[3541]), .Z(n35771) );
  XOR U35425 ( .A(n35773), .B(n35774), .Z(n35769) );
  AND U35426 ( .A(n35775), .B(n35776), .Z(n35774) );
  XNOR U35427 ( .A(p_input[3572]), .B(n35773), .Z(n35776) );
  XOR U35428 ( .A(n35773), .B(p_input[3540]), .Z(n35775) );
  XOR U35429 ( .A(n35777), .B(n35778), .Z(n35773) );
  AND U35430 ( .A(n35779), .B(n35780), .Z(n35778) );
  XNOR U35431 ( .A(p_input[3571]), .B(n35777), .Z(n35780) );
  XOR U35432 ( .A(n35777), .B(p_input[3539]), .Z(n35779) );
  XOR U35433 ( .A(n35781), .B(n35782), .Z(n35777) );
  AND U35434 ( .A(n35783), .B(n35784), .Z(n35782) );
  XNOR U35435 ( .A(p_input[3570]), .B(n35781), .Z(n35784) );
  XOR U35436 ( .A(n35781), .B(p_input[3538]), .Z(n35783) );
  XOR U35437 ( .A(n35785), .B(n35786), .Z(n35781) );
  AND U35438 ( .A(n35787), .B(n35788), .Z(n35786) );
  XNOR U35439 ( .A(p_input[3569]), .B(n35785), .Z(n35788) );
  XOR U35440 ( .A(n35785), .B(p_input[3537]), .Z(n35787) );
  XOR U35441 ( .A(n35789), .B(n35790), .Z(n35785) );
  AND U35442 ( .A(n35791), .B(n35792), .Z(n35790) );
  XNOR U35443 ( .A(p_input[3568]), .B(n35789), .Z(n35792) );
  XOR U35444 ( .A(n35789), .B(p_input[3536]), .Z(n35791) );
  XOR U35445 ( .A(n35793), .B(n35794), .Z(n35789) );
  AND U35446 ( .A(n35795), .B(n35796), .Z(n35794) );
  XNOR U35447 ( .A(p_input[3567]), .B(n35793), .Z(n35796) );
  XOR U35448 ( .A(n35793), .B(p_input[3535]), .Z(n35795) );
  XOR U35449 ( .A(n35797), .B(n35798), .Z(n35793) );
  AND U35450 ( .A(n35799), .B(n35800), .Z(n35798) );
  XNOR U35451 ( .A(p_input[3566]), .B(n35797), .Z(n35800) );
  XOR U35452 ( .A(n35797), .B(p_input[3534]), .Z(n35799) );
  XOR U35453 ( .A(n35801), .B(n35802), .Z(n35797) );
  AND U35454 ( .A(n35803), .B(n35804), .Z(n35802) );
  XNOR U35455 ( .A(p_input[3565]), .B(n35801), .Z(n35804) );
  XOR U35456 ( .A(n35801), .B(p_input[3533]), .Z(n35803) );
  XOR U35457 ( .A(n35805), .B(n35806), .Z(n35801) );
  AND U35458 ( .A(n35807), .B(n35808), .Z(n35806) );
  XNOR U35459 ( .A(p_input[3564]), .B(n35805), .Z(n35808) );
  XOR U35460 ( .A(n35805), .B(p_input[3532]), .Z(n35807) );
  XOR U35461 ( .A(n35809), .B(n35810), .Z(n35805) );
  AND U35462 ( .A(n35811), .B(n35812), .Z(n35810) );
  XNOR U35463 ( .A(p_input[3563]), .B(n35809), .Z(n35812) );
  XOR U35464 ( .A(n35809), .B(p_input[3531]), .Z(n35811) );
  XOR U35465 ( .A(n35813), .B(n35814), .Z(n35809) );
  AND U35466 ( .A(n35815), .B(n35816), .Z(n35814) );
  XNOR U35467 ( .A(p_input[3562]), .B(n35813), .Z(n35816) );
  XOR U35468 ( .A(n35813), .B(p_input[3530]), .Z(n35815) );
  XOR U35469 ( .A(n35817), .B(n35818), .Z(n35813) );
  AND U35470 ( .A(n35819), .B(n35820), .Z(n35818) );
  XNOR U35471 ( .A(p_input[3561]), .B(n35817), .Z(n35820) );
  XOR U35472 ( .A(n35817), .B(p_input[3529]), .Z(n35819) );
  XOR U35473 ( .A(n35821), .B(n35822), .Z(n35817) );
  AND U35474 ( .A(n35823), .B(n35824), .Z(n35822) );
  XNOR U35475 ( .A(p_input[3560]), .B(n35821), .Z(n35824) );
  XOR U35476 ( .A(n35821), .B(p_input[3528]), .Z(n35823) );
  XOR U35477 ( .A(n35825), .B(n35826), .Z(n35821) );
  AND U35478 ( .A(n35827), .B(n35828), .Z(n35826) );
  XNOR U35479 ( .A(p_input[3559]), .B(n35825), .Z(n35828) );
  XOR U35480 ( .A(n35825), .B(p_input[3527]), .Z(n35827) );
  XOR U35481 ( .A(n35829), .B(n35830), .Z(n35825) );
  AND U35482 ( .A(n35831), .B(n35832), .Z(n35830) );
  XNOR U35483 ( .A(p_input[3558]), .B(n35829), .Z(n35832) );
  XOR U35484 ( .A(n35829), .B(p_input[3526]), .Z(n35831) );
  XOR U35485 ( .A(n35833), .B(n35834), .Z(n35829) );
  AND U35486 ( .A(n35835), .B(n35836), .Z(n35834) );
  XNOR U35487 ( .A(p_input[3557]), .B(n35833), .Z(n35836) );
  XOR U35488 ( .A(n35833), .B(p_input[3525]), .Z(n35835) );
  XOR U35489 ( .A(n35837), .B(n35838), .Z(n35833) );
  AND U35490 ( .A(n35839), .B(n35840), .Z(n35838) );
  XNOR U35491 ( .A(p_input[3556]), .B(n35837), .Z(n35840) );
  XOR U35492 ( .A(n35837), .B(p_input[3524]), .Z(n35839) );
  XOR U35493 ( .A(n35841), .B(n35842), .Z(n35837) );
  AND U35494 ( .A(n35843), .B(n35844), .Z(n35842) );
  XNOR U35495 ( .A(p_input[3555]), .B(n35841), .Z(n35844) );
  XOR U35496 ( .A(n35841), .B(p_input[3523]), .Z(n35843) );
  XOR U35497 ( .A(n35845), .B(n35846), .Z(n35841) );
  AND U35498 ( .A(n35847), .B(n35848), .Z(n35846) );
  XNOR U35499 ( .A(p_input[3554]), .B(n35845), .Z(n35848) );
  XOR U35500 ( .A(n35845), .B(p_input[3522]), .Z(n35847) );
  XNOR U35501 ( .A(n35849), .B(n35850), .Z(n35845) );
  AND U35502 ( .A(n35851), .B(n35852), .Z(n35850) );
  XOR U35503 ( .A(p_input[3553]), .B(n35849), .Z(n35852) );
  XNOR U35504 ( .A(p_input[3521]), .B(n35849), .Z(n35851) );
  AND U35505 ( .A(p_input[3552]), .B(n35853), .Z(n35849) );
  IV U35506 ( .A(p_input[3520]), .Z(n35853) );
  XNOR U35507 ( .A(p_input[3456]), .B(n35854), .Z(n35447) );
  AND U35508 ( .A(n717), .B(n35855), .Z(n35854) );
  XOR U35509 ( .A(p_input[3488]), .B(p_input[3456]), .Z(n35855) );
  XOR U35510 ( .A(n35856), .B(n35857), .Z(n717) );
  AND U35511 ( .A(n35858), .B(n35859), .Z(n35857) );
  XNOR U35512 ( .A(p_input[3519]), .B(n35856), .Z(n35859) );
  XOR U35513 ( .A(n35856), .B(p_input[3487]), .Z(n35858) );
  XOR U35514 ( .A(n35860), .B(n35861), .Z(n35856) );
  AND U35515 ( .A(n35862), .B(n35863), .Z(n35861) );
  XNOR U35516 ( .A(p_input[3518]), .B(n35860), .Z(n35863) );
  XNOR U35517 ( .A(n35860), .B(n35462), .Z(n35862) );
  IV U35518 ( .A(p_input[3486]), .Z(n35462) );
  XOR U35519 ( .A(n35864), .B(n35865), .Z(n35860) );
  AND U35520 ( .A(n35866), .B(n35867), .Z(n35865) );
  XNOR U35521 ( .A(p_input[3517]), .B(n35864), .Z(n35867) );
  XNOR U35522 ( .A(n35864), .B(n35471), .Z(n35866) );
  IV U35523 ( .A(p_input[3485]), .Z(n35471) );
  XOR U35524 ( .A(n35868), .B(n35869), .Z(n35864) );
  AND U35525 ( .A(n35870), .B(n35871), .Z(n35869) );
  XNOR U35526 ( .A(p_input[3516]), .B(n35868), .Z(n35871) );
  XNOR U35527 ( .A(n35868), .B(n35480), .Z(n35870) );
  IV U35528 ( .A(p_input[3484]), .Z(n35480) );
  XOR U35529 ( .A(n35872), .B(n35873), .Z(n35868) );
  AND U35530 ( .A(n35874), .B(n35875), .Z(n35873) );
  XNOR U35531 ( .A(p_input[3515]), .B(n35872), .Z(n35875) );
  XNOR U35532 ( .A(n35872), .B(n35489), .Z(n35874) );
  IV U35533 ( .A(p_input[3483]), .Z(n35489) );
  XOR U35534 ( .A(n35876), .B(n35877), .Z(n35872) );
  AND U35535 ( .A(n35878), .B(n35879), .Z(n35877) );
  XNOR U35536 ( .A(p_input[3514]), .B(n35876), .Z(n35879) );
  XNOR U35537 ( .A(n35876), .B(n35498), .Z(n35878) );
  IV U35538 ( .A(p_input[3482]), .Z(n35498) );
  XOR U35539 ( .A(n35880), .B(n35881), .Z(n35876) );
  AND U35540 ( .A(n35882), .B(n35883), .Z(n35881) );
  XNOR U35541 ( .A(p_input[3513]), .B(n35880), .Z(n35883) );
  XNOR U35542 ( .A(n35880), .B(n35507), .Z(n35882) );
  IV U35543 ( .A(p_input[3481]), .Z(n35507) );
  XOR U35544 ( .A(n35884), .B(n35885), .Z(n35880) );
  AND U35545 ( .A(n35886), .B(n35887), .Z(n35885) );
  XNOR U35546 ( .A(p_input[3512]), .B(n35884), .Z(n35887) );
  XNOR U35547 ( .A(n35884), .B(n35516), .Z(n35886) );
  IV U35548 ( .A(p_input[3480]), .Z(n35516) );
  XOR U35549 ( .A(n35888), .B(n35889), .Z(n35884) );
  AND U35550 ( .A(n35890), .B(n35891), .Z(n35889) );
  XNOR U35551 ( .A(p_input[3511]), .B(n35888), .Z(n35891) );
  XNOR U35552 ( .A(n35888), .B(n35525), .Z(n35890) );
  IV U35553 ( .A(p_input[3479]), .Z(n35525) );
  XOR U35554 ( .A(n35892), .B(n35893), .Z(n35888) );
  AND U35555 ( .A(n35894), .B(n35895), .Z(n35893) );
  XNOR U35556 ( .A(p_input[3510]), .B(n35892), .Z(n35895) );
  XNOR U35557 ( .A(n35892), .B(n35534), .Z(n35894) );
  IV U35558 ( .A(p_input[3478]), .Z(n35534) );
  XOR U35559 ( .A(n35896), .B(n35897), .Z(n35892) );
  AND U35560 ( .A(n35898), .B(n35899), .Z(n35897) );
  XNOR U35561 ( .A(p_input[3509]), .B(n35896), .Z(n35899) );
  XNOR U35562 ( .A(n35896), .B(n35543), .Z(n35898) );
  IV U35563 ( .A(p_input[3477]), .Z(n35543) );
  XOR U35564 ( .A(n35900), .B(n35901), .Z(n35896) );
  AND U35565 ( .A(n35902), .B(n35903), .Z(n35901) );
  XNOR U35566 ( .A(p_input[3508]), .B(n35900), .Z(n35903) );
  XNOR U35567 ( .A(n35900), .B(n35552), .Z(n35902) );
  IV U35568 ( .A(p_input[3476]), .Z(n35552) );
  XOR U35569 ( .A(n35904), .B(n35905), .Z(n35900) );
  AND U35570 ( .A(n35906), .B(n35907), .Z(n35905) );
  XNOR U35571 ( .A(p_input[3507]), .B(n35904), .Z(n35907) );
  XNOR U35572 ( .A(n35904), .B(n35561), .Z(n35906) );
  IV U35573 ( .A(p_input[3475]), .Z(n35561) );
  XOR U35574 ( .A(n35908), .B(n35909), .Z(n35904) );
  AND U35575 ( .A(n35910), .B(n35911), .Z(n35909) );
  XNOR U35576 ( .A(p_input[3506]), .B(n35908), .Z(n35911) );
  XNOR U35577 ( .A(n35908), .B(n35570), .Z(n35910) );
  IV U35578 ( .A(p_input[3474]), .Z(n35570) );
  XOR U35579 ( .A(n35912), .B(n35913), .Z(n35908) );
  AND U35580 ( .A(n35914), .B(n35915), .Z(n35913) );
  XNOR U35581 ( .A(p_input[3505]), .B(n35912), .Z(n35915) );
  XNOR U35582 ( .A(n35912), .B(n35579), .Z(n35914) );
  IV U35583 ( .A(p_input[3473]), .Z(n35579) );
  XOR U35584 ( .A(n35916), .B(n35917), .Z(n35912) );
  AND U35585 ( .A(n35918), .B(n35919), .Z(n35917) );
  XNOR U35586 ( .A(p_input[3504]), .B(n35916), .Z(n35919) );
  XNOR U35587 ( .A(n35916), .B(n35588), .Z(n35918) );
  IV U35588 ( .A(p_input[3472]), .Z(n35588) );
  XOR U35589 ( .A(n35920), .B(n35921), .Z(n35916) );
  AND U35590 ( .A(n35922), .B(n35923), .Z(n35921) );
  XNOR U35591 ( .A(p_input[3503]), .B(n35920), .Z(n35923) );
  XNOR U35592 ( .A(n35920), .B(n35597), .Z(n35922) );
  IV U35593 ( .A(p_input[3471]), .Z(n35597) );
  XOR U35594 ( .A(n35924), .B(n35925), .Z(n35920) );
  AND U35595 ( .A(n35926), .B(n35927), .Z(n35925) );
  XNOR U35596 ( .A(p_input[3502]), .B(n35924), .Z(n35927) );
  XNOR U35597 ( .A(n35924), .B(n35606), .Z(n35926) );
  IV U35598 ( .A(p_input[3470]), .Z(n35606) );
  XOR U35599 ( .A(n35928), .B(n35929), .Z(n35924) );
  AND U35600 ( .A(n35930), .B(n35931), .Z(n35929) );
  XNOR U35601 ( .A(p_input[3501]), .B(n35928), .Z(n35931) );
  XNOR U35602 ( .A(n35928), .B(n35615), .Z(n35930) );
  IV U35603 ( .A(p_input[3469]), .Z(n35615) );
  XOR U35604 ( .A(n35932), .B(n35933), .Z(n35928) );
  AND U35605 ( .A(n35934), .B(n35935), .Z(n35933) );
  XNOR U35606 ( .A(p_input[3500]), .B(n35932), .Z(n35935) );
  XNOR U35607 ( .A(n35932), .B(n35624), .Z(n35934) );
  IV U35608 ( .A(p_input[3468]), .Z(n35624) );
  XOR U35609 ( .A(n35936), .B(n35937), .Z(n35932) );
  AND U35610 ( .A(n35938), .B(n35939), .Z(n35937) );
  XNOR U35611 ( .A(p_input[3499]), .B(n35936), .Z(n35939) );
  XNOR U35612 ( .A(n35936), .B(n35633), .Z(n35938) );
  IV U35613 ( .A(p_input[3467]), .Z(n35633) );
  XOR U35614 ( .A(n35940), .B(n35941), .Z(n35936) );
  AND U35615 ( .A(n35942), .B(n35943), .Z(n35941) );
  XNOR U35616 ( .A(p_input[3498]), .B(n35940), .Z(n35943) );
  XNOR U35617 ( .A(n35940), .B(n35642), .Z(n35942) );
  IV U35618 ( .A(p_input[3466]), .Z(n35642) );
  XOR U35619 ( .A(n35944), .B(n35945), .Z(n35940) );
  AND U35620 ( .A(n35946), .B(n35947), .Z(n35945) );
  XNOR U35621 ( .A(p_input[3497]), .B(n35944), .Z(n35947) );
  XNOR U35622 ( .A(n35944), .B(n35651), .Z(n35946) );
  IV U35623 ( .A(p_input[3465]), .Z(n35651) );
  XOR U35624 ( .A(n35948), .B(n35949), .Z(n35944) );
  AND U35625 ( .A(n35950), .B(n35951), .Z(n35949) );
  XNOR U35626 ( .A(p_input[3496]), .B(n35948), .Z(n35951) );
  XNOR U35627 ( .A(n35948), .B(n35660), .Z(n35950) );
  IV U35628 ( .A(p_input[3464]), .Z(n35660) );
  XOR U35629 ( .A(n35952), .B(n35953), .Z(n35948) );
  AND U35630 ( .A(n35954), .B(n35955), .Z(n35953) );
  XNOR U35631 ( .A(p_input[3495]), .B(n35952), .Z(n35955) );
  XNOR U35632 ( .A(n35952), .B(n35669), .Z(n35954) );
  IV U35633 ( .A(p_input[3463]), .Z(n35669) );
  XOR U35634 ( .A(n35956), .B(n35957), .Z(n35952) );
  AND U35635 ( .A(n35958), .B(n35959), .Z(n35957) );
  XNOR U35636 ( .A(p_input[3494]), .B(n35956), .Z(n35959) );
  XNOR U35637 ( .A(n35956), .B(n35678), .Z(n35958) );
  IV U35638 ( .A(p_input[3462]), .Z(n35678) );
  XOR U35639 ( .A(n35960), .B(n35961), .Z(n35956) );
  AND U35640 ( .A(n35962), .B(n35963), .Z(n35961) );
  XNOR U35641 ( .A(p_input[3493]), .B(n35960), .Z(n35963) );
  XNOR U35642 ( .A(n35960), .B(n35687), .Z(n35962) );
  IV U35643 ( .A(p_input[3461]), .Z(n35687) );
  XOR U35644 ( .A(n35964), .B(n35965), .Z(n35960) );
  AND U35645 ( .A(n35966), .B(n35967), .Z(n35965) );
  XNOR U35646 ( .A(p_input[3492]), .B(n35964), .Z(n35967) );
  XNOR U35647 ( .A(n35964), .B(n35696), .Z(n35966) );
  IV U35648 ( .A(p_input[3460]), .Z(n35696) );
  XOR U35649 ( .A(n35968), .B(n35969), .Z(n35964) );
  AND U35650 ( .A(n35970), .B(n35971), .Z(n35969) );
  XNOR U35651 ( .A(p_input[3491]), .B(n35968), .Z(n35971) );
  XNOR U35652 ( .A(n35968), .B(n35705), .Z(n35970) );
  IV U35653 ( .A(p_input[3459]), .Z(n35705) );
  XOR U35654 ( .A(n35972), .B(n35973), .Z(n35968) );
  AND U35655 ( .A(n35974), .B(n35975), .Z(n35973) );
  XNOR U35656 ( .A(p_input[3490]), .B(n35972), .Z(n35975) );
  XNOR U35657 ( .A(n35972), .B(n35714), .Z(n35974) );
  IV U35658 ( .A(p_input[3458]), .Z(n35714) );
  XNOR U35659 ( .A(n35976), .B(n35977), .Z(n35972) );
  AND U35660 ( .A(n35978), .B(n35979), .Z(n35977) );
  XOR U35661 ( .A(p_input[3489]), .B(n35976), .Z(n35979) );
  XNOR U35662 ( .A(p_input[3457]), .B(n35976), .Z(n35978) );
  AND U35663 ( .A(p_input[3488]), .B(n35980), .Z(n35976) );
  IV U35664 ( .A(p_input[3456]), .Z(n35980) );
  XOR U35665 ( .A(n35981), .B(n35982), .Z(n35070) );
  AND U35666 ( .A(n573), .B(n35983), .Z(n35982) );
  XNOR U35667 ( .A(n35984), .B(n35981), .Z(n35983) );
  XOR U35668 ( .A(n35985), .B(n35986), .Z(n573) );
  AND U35669 ( .A(n35987), .B(n35988), .Z(n35986) );
  XNOR U35670 ( .A(n35085), .B(n35985), .Z(n35988) );
  AND U35671 ( .A(p_input[3455]), .B(p_input[3423]), .Z(n35085) );
  XNOR U35672 ( .A(n35985), .B(n35082), .Z(n35987) );
  IV U35673 ( .A(n35989), .Z(n35082) );
  AND U35674 ( .A(p_input[3359]), .B(p_input[3391]), .Z(n35989) );
  XOR U35675 ( .A(n35990), .B(n35991), .Z(n35985) );
  AND U35676 ( .A(n35992), .B(n35993), .Z(n35991) );
  XOR U35677 ( .A(n35990), .B(n35097), .Z(n35993) );
  XNOR U35678 ( .A(p_input[3422]), .B(n35994), .Z(n35097) );
  AND U35679 ( .A(n723), .B(n35995), .Z(n35994) );
  XOR U35680 ( .A(p_input[3454]), .B(p_input[3422]), .Z(n35995) );
  XNOR U35681 ( .A(n35094), .B(n35990), .Z(n35992) );
  XOR U35682 ( .A(n35996), .B(n35997), .Z(n35094) );
  AND U35683 ( .A(n720), .B(n35998), .Z(n35997) );
  XOR U35684 ( .A(p_input[3390]), .B(p_input[3358]), .Z(n35998) );
  XOR U35685 ( .A(n35999), .B(n36000), .Z(n35990) );
  AND U35686 ( .A(n36001), .B(n36002), .Z(n36000) );
  XOR U35687 ( .A(n35999), .B(n35109), .Z(n36002) );
  XNOR U35688 ( .A(p_input[3421]), .B(n36003), .Z(n35109) );
  AND U35689 ( .A(n723), .B(n36004), .Z(n36003) );
  XOR U35690 ( .A(p_input[3453]), .B(p_input[3421]), .Z(n36004) );
  XNOR U35691 ( .A(n35106), .B(n35999), .Z(n36001) );
  XOR U35692 ( .A(n36005), .B(n36006), .Z(n35106) );
  AND U35693 ( .A(n720), .B(n36007), .Z(n36006) );
  XOR U35694 ( .A(p_input[3389]), .B(p_input[3357]), .Z(n36007) );
  XOR U35695 ( .A(n36008), .B(n36009), .Z(n35999) );
  AND U35696 ( .A(n36010), .B(n36011), .Z(n36009) );
  XOR U35697 ( .A(n36008), .B(n35121), .Z(n36011) );
  XNOR U35698 ( .A(p_input[3420]), .B(n36012), .Z(n35121) );
  AND U35699 ( .A(n723), .B(n36013), .Z(n36012) );
  XOR U35700 ( .A(p_input[3452]), .B(p_input[3420]), .Z(n36013) );
  XNOR U35701 ( .A(n35118), .B(n36008), .Z(n36010) );
  XOR U35702 ( .A(n36014), .B(n36015), .Z(n35118) );
  AND U35703 ( .A(n720), .B(n36016), .Z(n36015) );
  XOR U35704 ( .A(p_input[3388]), .B(p_input[3356]), .Z(n36016) );
  XOR U35705 ( .A(n36017), .B(n36018), .Z(n36008) );
  AND U35706 ( .A(n36019), .B(n36020), .Z(n36018) );
  XOR U35707 ( .A(n36017), .B(n35133), .Z(n36020) );
  XNOR U35708 ( .A(p_input[3419]), .B(n36021), .Z(n35133) );
  AND U35709 ( .A(n723), .B(n36022), .Z(n36021) );
  XOR U35710 ( .A(p_input[3451]), .B(p_input[3419]), .Z(n36022) );
  XNOR U35711 ( .A(n35130), .B(n36017), .Z(n36019) );
  XOR U35712 ( .A(n36023), .B(n36024), .Z(n35130) );
  AND U35713 ( .A(n720), .B(n36025), .Z(n36024) );
  XOR U35714 ( .A(p_input[3387]), .B(p_input[3355]), .Z(n36025) );
  XOR U35715 ( .A(n36026), .B(n36027), .Z(n36017) );
  AND U35716 ( .A(n36028), .B(n36029), .Z(n36027) );
  XOR U35717 ( .A(n36026), .B(n35145), .Z(n36029) );
  XNOR U35718 ( .A(p_input[3418]), .B(n36030), .Z(n35145) );
  AND U35719 ( .A(n723), .B(n36031), .Z(n36030) );
  XOR U35720 ( .A(p_input[3450]), .B(p_input[3418]), .Z(n36031) );
  XNOR U35721 ( .A(n35142), .B(n36026), .Z(n36028) );
  XOR U35722 ( .A(n36032), .B(n36033), .Z(n35142) );
  AND U35723 ( .A(n720), .B(n36034), .Z(n36033) );
  XOR U35724 ( .A(p_input[3386]), .B(p_input[3354]), .Z(n36034) );
  XOR U35725 ( .A(n36035), .B(n36036), .Z(n36026) );
  AND U35726 ( .A(n36037), .B(n36038), .Z(n36036) );
  XOR U35727 ( .A(n36035), .B(n35157), .Z(n36038) );
  XNOR U35728 ( .A(p_input[3417]), .B(n36039), .Z(n35157) );
  AND U35729 ( .A(n723), .B(n36040), .Z(n36039) );
  XOR U35730 ( .A(p_input[3449]), .B(p_input[3417]), .Z(n36040) );
  XNOR U35731 ( .A(n35154), .B(n36035), .Z(n36037) );
  XOR U35732 ( .A(n36041), .B(n36042), .Z(n35154) );
  AND U35733 ( .A(n720), .B(n36043), .Z(n36042) );
  XOR U35734 ( .A(p_input[3385]), .B(p_input[3353]), .Z(n36043) );
  XOR U35735 ( .A(n36044), .B(n36045), .Z(n36035) );
  AND U35736 ( .A(n36046), .B(n36047), .Z(n36045) );
  XOR U35737 ( .A(n36044), .B(n35169), .Z(n36047) );
  XNOR U35738 ( .A(p_input[3416]), .B(n36048), .Z(n35169) );
  AND U35739 ( .A(n723), .B(n36049), .Z(n36048) );
  XOR U35740 ( .A(p_input[3448]), .B(p_input[3416]), .Z(n36049) );
  XNOR U35741 ( .A(n35166), .B(n36044), .Z(n36046) );
  XOR U35742 ( .A(n36050), .B(n36051), .Z(n35166) );
  AND U35743 ( .A(n720), .B(n36052), .Z(n36051) );
  XOR U35744 ( .A(p_input[3384]), .B(p_input[3352]), .Z(n36052) );
  XOR U35745 ( .A(n36053), .B(n36054), .Z(n36044) );
  AND U35746 ( .A(n36055), .B(n36056), .Z(n36054) );
  XOR U35747 ( .A(n36053), .B(n35181), .Z(n36056) );
  XNOR U35748 ( .A(p_input[3415]), .B(n36057), .Z(n35181) );
  AND U35749 ( .A(n723), .B(n36058), .Z(n36057) );
  XOR U35750 ( .A(p_input[3447]), .B(p_input[3415]), .Z(n36058) );
  XNOR U35751 ( .A(n35178), .B(n36053), .Z(n36055) );
  XOR U35752 ( .A(n36059), .B(n36060), .Z(n35178) );
  AND U35753 ( .A(n720), .B(n36061), .Z(n36060) );
  XOR U35754 ( .A(p_input[3383]), .B(p_input[3351]), .Z(n36061) );
  XOR U35755 ( .A(n36062), .B(n36063), .Z(n36053) );
  AND U35756 ( .A(n36064), .B(n36065), .Z(n36063) );
  XOR U35757 ( .A(n36062), .B(n35193), .Z(n36065) );
  XNOR U35758 ( .A(p_input[3414]), .B(n36066), .Z(n35193) );
  AND U35759 ( .A(n723), .B(n36067), .Z(n36066) );
  XOR U35760 ( .A(p_input[3446]), .B(p_input[3414]), .Z(n36067) );
  XNOR U35761 ( .A(n35190), .B(n36062), .Z(n36064) );
  XOR U35762 ( .A(n36068), .B(n36069), .Z(n35190) );
  AND U35763 ( .A(n720), .B(n36070), .Z(n36069) );
  XOR U35764 ( .A(p_input[3382]), .B(p_input[3350]), .Z(n36070) );
  XOR U35765 ( .A(n36071), .B(n36072), .Z(n36062) );
  AND U35766 ( .A(n36073), .B(n36074), .Z(n36072) );
  XOR U35767 ( .A(n36071), .B(n35205), .Z(n36074) );
  XNOR U35768 ( .A(p_input[3413]), .B(n36075), .Z(n35205) );
  AND U35769 ( .A(n723), .B(n36076), .Z(n36075) );
  XOR U35770 ( .A(p_input[3445]), .B(p_input[3413]), .Z(n36076) );
  XNOR U35771 ( .A(n35202), .B(n36071), .Z(n36073) );
  XOR U35772 ( .A(n36077), .B(n36078), .Z(n35202) );
  AND U35773 ( .A(n720), .B(n36079), .Z(n36078) );
  XOR U35774 ( .A(p_input[3381]), .B(p_input[3349]), .Z(n36079) );
  XOR U35775 ( .A(n36080), .B(n36081), .Z(n36071) );
  AND U35776 ( .A(n36082), .B(n36083), .Z(n36081) );
  XOR U35777 ( .A(n36080), .B(n35217), .Z(n36083) );
  XNOR U35778 ( .A(p_input[3412]), .B(n36084), .Z(n35217) );
  AND U35779 ( .A(n723), .B(n36085), .Z(n36084) );
  XOR U35780 ( .A(p_input[3444]), .B(p_input[3412]), .Z(n36085) );
  XNOR U35781 ( .A(n35214), .B(n36080), .Z(n36082) );
  XOR U35782 ( .A(n36086), .B(n36087), .Z(n35214) );
  AND U35783 ( .A(n720), .B(n36088), .Z(n36087) );
  XOR U35784 ( .A(p_input[3380]), .B(p_input[3348]), .Z(n36088) );
  XOR U35785 ( .A(n36089), .B(n36090), .Z(n36080) );
  AND U35786 ( .A(n36091), .B(n36092), .Z(n36090) );
  XOR U35787 ( .A(n36089), .B(n35229), .Z(n36092) );
  XNOR U35788 ( .A(p_input[3411]), .B(n36093), .Z(n35229) );
  AND U35789 ( .A(n723), .B(n36094), .Z(n36093) );
  XOR U35790 ( .A(p_input[3443]), .B(p_input[3411]), .Z(n36094) );
  XNOR U35791 ( .A(n35226), .B(n36089), .Z(n36091) );
  XOR U35792 ( .A(n36095), .B(n36096), .Z(n35226) );
  AND U35793 ( .A(n720), .B(n36097), .Z(n36096) );
  XOR U35794 ( .A(p_input[3379]), .B(p_input[3347]), .Z(n36097) );
  XOR U35795 ( .A(n36098), .B(n36099), .Z(n36089) );
  AND U35796 ( .A(n36100), .B(n36101), .Z(n36099) );
  XOR U35797 ( .A(n36098), .B(n35241), .Z(n36101) );
  XNOR U35798 ( .A(p_input[3410]), .B(n36102), .Z(n35241) );
  AND U35799 ( .A(n723), .B(n36103), .Z(n36102) );
  XOR U35800 ( .A(p_input[3442]), .B(p_input[3410]), .Z(n36103) );
  XNOR U35801 ( .A(n35238), .B(n36098), .Z(n36100) );
  XOR U35802 ( .A(n36104), .B(n36105), .Z(n35238) );
  AND U35803 ( .A(n720), .B(n36106), .Z(n36105) );
  XOR U35804 ( .A(p_input[3378]), .B(p_input[3346]), .Z(n36106) );
  XOR U35805 ( .A(n36107), .B(n36108), .Z(n36098) );
  AND U35806 ( .A(n36109), .B(n36110), .Z(n36108) );
  XOR U35807 ( .A(n36107), .B(n35253), .Z(n36110) );
  XNOR U35808 ( .A(p_input[3409]), .B(n36111), .Z(n35253) );
  AND U35809 ( .A(n723), .B(n36112), .Z(n36111) );
  XOR U35810 ( .A(p_input[3441]), .B(p_input[3409]), .Z(n36112) );
  XNOR U35811 ( .A(n35250), .B(n36107), .Z(n36109) );
  XOR U35812 ( .A(n36113), .B(n36114), .Z(n35250) );
  AND U35813 ( .A(n720), .B(n36115), .Z(n36114) );
  XOR U35814 ( .A(p_input[3377]), .B(p_input[3345]), .Z(n36115) );
  XOR U35815 ( .A(n36116), .B(n36117), .Z(n36107) );
  AND U35816 ( .A(n36118), .B(n36119), .Z(n36117) );
  XOR U35817 ( .A(n36116), .B(n35265), .Z(n36119) );
  XNOR U35818 ( .A(p_input[3408]), .B(n36120), .Z(n35265) );
  AND U35819 ( .A(n723), .B(n36121), .Z(n36120) );
  XOR U35820 ( .A(p_input[3440]), .B(p_input[3408]), .Z(n36121) );
  XNOR U35821 ( .A(n35262), .B(n36116), .Z(n36118) );
  XOR U35822 ( .A(n36122), .B(n36123), .Z(n35262) );
  AND U35823 ( .A(n720), .B(n36124), .Z(n36123) );
  XOR U35824 ( .A(p_input[3376]), .B(p_input[3344]), .Z(n36124) );
  XOR U35825 ( .A(n36125), .B(n36126), .Z(n36116) );
  AND U35826 ( .A(n36127), .B(n36128), .Z(n36126) );
  XOR U35827 ( .A(n36125), .B(n35277), .Z(n36128) );
  XNOR U35828 ( .A(p_input[3407]), .B(n36129), .Z(n35277) );
  AND U35829 ( .A(n723), .B(n36130), .Z(n36129) );
  XOR U35830 ( .A(p_input[3439]), .B(p_input[3407]), .Z(n36130) );
  XNOR U35831 ( .A(n35274), .B(n36125), .Z(n36127) );
  XOR U35832 ( .A(n36131), .B(n36132), .Z(n35274) );
  AND U35833 ( .A(n720), .B(n36133), .Z(n36132) );
  XOR U35834 ( .A(p_input[3375]), .B(p_input[3343]), .Z(n36133) );
  XOR U35835 ( .A(n36134), .B(n36135), .Z(n36125) );
  AND U35836 ( .A(n36136), .B(n36137), .Z(n36135) );
  XOR U35837 ( .A(n36134), .B(n35289), .Z(n36137) );
  XNOR U35838 ( .A(p_input[3406]), .B(n36138), .Z(n35289) );
  AND U35839 ( .A(n723), .B(n36139), .Z(n36138) );
  XOR U35840 ( .A(p_input[3438]), .B(p_input[3406]), .Z(n36139) );
  XNOR U35841 ( .A(n35286), .B(n36134), .Z(n36136) );
  XOR U35842 ( .A(n36140), .B(n36141), .Z(n35286) );
  AND U35843 ( .A(n720), .B(n36142), .Z(n36141) );
  XOR U35844 ( .A(p_input[3374]), .B(p_input[3342]), .Z(n36142) );
  XOR U35845 ( .A(n36143), .B(n36144), .Z(n36134) );
  AND U35846 ( .A(n36145), .B(n36146), .Z(n36144) );
  XOR U35847 ( .A(n36143), .B(n35301), .Z(n36146) );
  XNOR U35848 ( .A(p_input[3405]), .B(n36147), .Z(n35301) );
  AND U35849 ( .A(n723), .B(n36148), .Z(n36147) );
  XOR U35850 ( .A(p_input[3437]), .B(p_input[3405]), .Z(n36148) );
  XNOR U35851 ( .A(n35298), .B(n36143), .Z(n36145) );
  XOR U35852 ( .A(n36149), .B(n36150), .Z(n35298) );
  AND U35853 ( .A(n720), .B(n36151), .Z(n36150) );
  XOR U35854 ( .A(p_input[3373]), .B(p_input[3341]), .Z(n36151) );
  XOR U35855 ( .A(n36152), .B(n36153), .Z(n36143) );
  AND U35856 ( .A(n36154), .B(n36155), .Z(n36153) );
  XOR U35857 ( .A(n36152), .B(n35313), .Z(n36155) );
  XNOR U35858 ( .A(p_input[3404]), .B(n36156), .Z(n35313) );
  AND U35859 ( .A(n723), .B(n36157), .Z(n36156) );
  XOR U35860 ( .A(p_input[3436]), .B(p_input[3404]), .Z(n36157) );
  XNOR U35861 ( .A(n35310), .B(n36152), .Z(n36154) );
  XOR U35862 ( .A(n36158), .B(n36159), .Z(n35310) );
  AND U35863 ( .A(n720), .B(n36160), .Z(n36159) );
  XOR U35864 ( .A(p_input[3372]), .B(p_input[3340]), .Z(n36160) );
  XOR U35865 ( .A(n36161), .B(n36162), .Z(n36152) );
  AND U35866 ( .A(n36163), .B(n36164), .Z(n36162) );
  XOR U35867 ( .A(n36161), .B(n35325), .Z(n36164) );
  XNOR U35868 ( .A(p_input[3403]), .B(n36165), .Z(n35325) );
  AND U35869 ( .A(n723), .B(n36166), .Z(n36165) );
  XOR U35870 ( .A(p_input[3435]), .B(p_input[3403]), .Z(n36166) );
  XNOR U35871 ( .A(n35322), .B(n36161), .Z(n36163) );
  XOR U35872 ( .A(n36167), .B(n36168), .Z(n35322) );
  AND U35873 ( .A(n720), .B(n36169), .Z(n36168) );
  XOR U35874 ( .A(p_input[3371]), .B(p_input[3339]), .Z(n36169) );
  XOR U35875 ( .A(n36170), .B(n36171), .Z(n36161) );
  AND U35876 ( .A(n36172), .B(n36173), .Z(n36171) );
  XOR U35877 ( .A(n36170), .B(n35337), .Z(n36173) );
  XNOR U35878 ( .A(p_input[3402]), .B(n36174), .Z(n35337) );
  AND U35879 ( .A(n723), .B(n36175), .Z(n36174) );
  XOR U35880 ( .A(p_input[3434]), .B(p_input[3402]), .Z(n36175) );
  XNOR U35881 ( .A(n35334), .B(n36170), .Z(n36172) );
  XOR U35882 ( .A(n36176), .B(n36177), .Z(n35334) );
  AND U35883 ( .A(n720), .B(n36178), .Z(n36177) );
  XOR U35884 ( .A(p_input[3370]), .B(p_input[3338]), .Z(n36178) );
  XOR U35885 ( .A(n36179), .B(n36180), .Z(n36170) );
  AND U35886 ( .A(n36181), .B(n36182), .Z(n36180) );
  XOR U35887 ( .A(n36179), .B(n35349), .Z(n36182) );
  XNOR U35888 ( .A(p_input[3401]), .B(n36183), .Z(n35349) );
  AND U35889 ( .A(n723), .B(n36184), .Z(n36183) );
  XOR U35890 ( .A(p_input[3433]), .B(p_input[3401]), .Z(n36184) );
  XNOR U35891 ( .A(n35346), .B(n36179), .Z(n36181) );
  XOR U35892 ( .A(n36185), .B(n36186), .Z(n35346) );
  AND U35893 ( .A(n720), .B(n36187), .Z(n36186) );
  XOR U35894 ( .A(p_input[3369]), .B(p_input[3337]), .Z(n36187) );
  XOR U35895 ( .A(n36188), .B(n36189), .Z(n36179) );
  AND U35896 ( .A(n36190), .B(n36191), .Z(n36189) );
  XOR U35897 ( .A(n36188), .B(n35361), .Z(n36191) );
  XNOR U35898 ( .A(p_input[3400]), .B(n36192), .Z(n35361) );
  AND U35899 ( .A(n723), .B(n36193), .Z(n36192) );
  XOR U35900 ( .A(p_input[3432]), .B(p_input[3400]), .Z(n36193) );
  XNOR U35901 ( .A(n35358), .B(n36188), .Z(n36190) );
  XOR U35902 ( .A(n36194), .B(n36195), .Z(n35358) );
  AND U35903 ( .A(n720), .B(n36196), .Z(n36195) );
  XOR U35904 ( .A(p_input[3368]), .B(p_input[3336]), .Z(n36196) );
  XOR U35905 ( .A(n36197), .B(n36198), .Z(n36188) );
  AND U35906 ( .A(n36199), .B(n36200), .Z(n36198) );
  XOR U35907 ( .A(n36197), .B(n35373), .Z(n36200) );
  XNOR U35908 ( .A(p_input[3399]), .B(n36201), .Z(n35373) );
  AND U35909 ( .A(n723), .B(n36202), .Z(n36201) );
  XOR U35910 ( .A(p_input[3431]), .B(p_input[3399]), .Z(n36202) );
  XNOR U35911 ( .A(n35370), .B(n36197), .Z(n36199) );
  XOR U35912 ( .A(n36203), .B(n36204), .Z(n35370) );
  AND U35913 ( .A(n720), .B(n36205), .Z(n36204) );
  XOR U35914 ( .A(p_input[3367]), .B(p_input[3335]), .Z(n36205) );
  XOR U35915 ( .A(n36206), .B(n36207), .Z(n36197) );
  AND U35916 ( .A(n36208), .B(n36209), .Z(n36207) );
  XOR U35917 ( .A(n36206), .B(n35385), .Z(n36209) );
  XNOR U35918 ( .A(p_input[3398]), .B(n36210), .Z(n35385) );
  AND U35919 ( .A(n723), .B(n36211), .Z(n36210) );
  XOR U35920 ( .A(p_input[3430]), .B(p_input[3398]), .Z(n36211) );
  XNOR U35921 ( .A(n35382), .B(n36206), .Z(n36208) );
  XOR U35922 ( .A(n36212), .B(n36213), .Z(n35382) );
  AND U35923 ( .A(n720), .B(n36214), .Z(n36213) );
  XOR U35924 ( .A(p_input[3366]), .B(p_input[3334]), .Z(n36214) );
  XOR U35925 ( .A(n36215), .B(n36216), .Z(n36206) );
  AND U35926 ( .A(n36217), .B(n36218), .Z(n36216) );
  XOR U35927 ( .A(n36215), .B(n35397), .Z(n36218) );
  XNOR U35928 ( .A(p_input[3397]), .B(n36219), .Z(n35397) );
  AND U35929 ( .A(n723), .B(n36220), .Z(n36219) );
  XOR U35930 ( .A(p_input[3429]), .B(p_input[3397]), .Z(n36220) );
  XNOR U35931 ( .A(n35394), .B(n36215), .Z(n36217) );
  XOR U35932 ( .A(n36221), .B(n36222), .Z(n35394) );
  AND U35933 ( .A(n720), .B(n36223), .Z(n36222) );
  XOR U35934 ( .A(p_input[3365]), .B(p_input[3333]), .Z(n36223) );
  XOR U35935 ( .A(n36224), .B(n36225), .Z(n36215) );
  AND U35936 ( .A(n36226), .B(n36227), .Z(n36225) );
  XOR U35937 ( .A(n36224), .B(n35409), .Z(n36227) );
  XNOR U35938 ( .A(p_input[3396]), .B(n36228), .Z(n35409) );
  AND U35939 ( .A(n723), .B(n36229), .Z(n36228) );
  XOR U35940 ( .A(p_input[3428]), .B(p_input[3396]), .Z(n36229) );
  XNOR U35941 ( .A(n35406), .B(n36224), .Z(n36226) );
  XOR U35942 ( .A(n36230), .B(n36231), .Z(n35406) );
  AND U35943 ( .A(n720), .B(n36232), .Z(n36231) );
  XOR U35944 ( .A(p_input[3364]), .B(p_input[3332]), .Z(n36232) );
  XOR U35945 ( .A(n36233), .B(n36234), .Z(n36224) );
  AND U35946 ( .A(n36235), .B(n36236), .Z(n36234) );
  XOR U35947 ( .A(n36233), .B(n35421), .Z(n36236) );
  XNOR U35948 ( .A(p_input[3395]), .B(n36237), .Z(n35421) );
  AND U35949 ( .A(n723), .B(n36238), .Z(n36237) );
  XOR U35950 ( .A(p_input[3427]), .B(p_input[3395]), .Z(n36238) );
  XNOR U35951 ( .A(n35418), .B(n36233), .Z(n36235) );
  XOR U35952 ( .A(n36239), .B(n36240), .Z(n35418) );
  AND U35953 ( .A(n720), .B(n36241), .Z(n36240) );
  XOR U35954 ( .A(p_input[3363]), .B(p_input[3331]), .Z(n36241) );
  XOR U35955 ( .A(n36242), .B(n36243), .Z(n36233) );
  AND U35956 ( .A(n36244), .B(n36245), .Z(n36243) );
  XOR U35957 ( .A(n36242), .B(n35433), .Z(n36245) );
  XNOR U35958 ( .A(p_input[3394]), .B(n36246), .Z(n35433) );
  AND U35959 ( .A(n723), .B(n36247), .Z(n36246) );
  XOR U35960 ( .A(p_input[3426]), .B(p_input[3394]), .Z(n36247) );
  XNOR U35961 ( .A(n35430), .B(n36242), .Z(n36244) );
  XOR U35962 ( .A(n36248), .B(n36249), .Z(n35430) );
  AND U35963 ( .A(n720), .B(n36250), .Z(n36249) );
  XOR U35964 ( .A(p_input[3362]), .B(p_input[3330]), .Z(n36250) );
  XOR U35965 ( .A(n36251), .B(n36252), .Z(n36242) );
  AND U35966 ( .A(n36253), .B(n36254), .Z(n36252) );
  XNOR U35967 ( .A(n36255), .B(n35446), .Z(n36254) );
  XNOR U35968 ( .A(p_input[3393]), .B(n36256), .Z(n35446) );
  AND U35969 ( .A(n723), .B(n36257), .Z(n36256) );
  XNOR U35970 ( .A(p_input[3425]), .B(n36258), .Z(n36257) );
  IV U35971 ( .A(p_input[3393]), .Z(n36258) );
  XNOR U35972 ( .A(n35443), .B(n36251), .Z(n36253) );
  XNOR U35973 ( .A(p_input[3329]), .B(n36259), .Z(n35443) );
  AND U35974 ( .A(n720), .B(n36260), .Z(n36259) );
  XOR U35975 ( .A(p_input[3361]), .B(p_input[3329]), .Z(n36260) );
  IV U35976 ( .A(n36255), .Z(n36251) );
  AND U35977 ( .A(n35981), .B(n35984), .Z(n36255) );
  XOR U35978 ( .A(p_input[3392]), .B(n36261), .Z(n35984) );
  AND U35979 ( .A(n723), .B(n36262), .Z(n36261) );
  XOR U35980 ( .A(p_input[3424]), .B(p_input[3392]), .Z(n36262) );
  XOR U35981 ( .A(n36263), .B(n36264), .Z(n723) );
  AND U35982 ( .A(n36265), .B(n36266), .Z(n36264) );
  XNOR U35983 ( .A(p_input[3455]), .B(n36263), .Z(n36266) );
  XOR U35984 ( .A(n36263), .B(p_input[3423]), .Z(n36265) );
  XOR U35985 ( .A(n36267), .B(n36268), .Z(n36263) );
  AND U35986 ( .A(n36269), .B(n36270), .Z(n36268) );
  XNOR U35987 ( .A(p_input[3454]), .B(n36267), .Z(n36270) );
  XOR U35988 ( .A(n36267), .B(p_input[3422]), .Z(n36269) );
  XOR U35989 ( .A(n36271), .B(n36272), .Z(n36267) );
  AND U35990 ( .A(n36273), .B(n36274), .Z(n36272) );
  XNOR U35991 ( .A(p_input[3453]), .B(n36271), .Z(n36274) );
  XOR U35992 ( .A(n36271), .B(p_input[3421]), .Z(n36273) );
  XOR U35993 ( .A(n36275), .B(n36276), .Z(n36271) );
  AND U35994 ( .A(n36277), .B(n36278), .Z(n36276) );
  XNOR U35995 ( .A(p_input[3452]), .B(n36275), .Z(n36278) );
  XOR U35996 ( .A(n36275), .B(p_input[3420]), .Z(n36277) );
  XOR U35997 ( .A(n36279), .B(n36280), .Z(n36275) );
  AND U35998 ( .A(n36281), .B(n36282), .Z(n36280) );
  XNOR U35999 ( .A(p_input[3451]), .B(n36279), .Z(n36282) );
  XOR U36000 ( .A(n36279), .B(p_input[3419]), .Z(n36281) );
  XOR U36001 ( .A(n36283), .B(n36284), .Z(n36279) );
  AND U36002 ( .A(n36285), .B(n36286), .Z(n36284) );
  XNOR U36003 ( .A(p_input[3450]), .B(n36283), .Z(n36286) );
  XOR U36004 ( .A(n36283), .B(p_input[3418]), .Z(n36285) );
  XOR U36005 ( .A(n36287), .B(n36288), .Z(n36283) );
  AND U36006 ( .A(n36289), .B(n36290), .Z(n36288) );
  XNOR U36007 ( .A(p_input[3449]), .B(n36287), .Z(n36290) );
  XOR U36008 ( .A(n36287), .B(p_input[3417]), .Z(n36289) );
  XOR U36009 ( .A(n36291), .B(n36292), .Z(n36287) );
  AND U36010 ( .A(n36293), .B(n36294), .Z(n36292) );
  XNOR U36011 ( .A(p_input[3448]), .B(n36291), .Z(n36294) );
  XOR U36012 ( .A(n36291), .B(p_input[3416]), .Z(n36293) );
  XOR U36013 ( .A(n36295), .B(n36296), .Z(n36291) );
  AND U36014 ( .A(n36297), .B(n36298), .Z(n36296) );
  XNOR U36015 ( .A(p_input[3447]), .B(n36295), .Z(n36298) );
  XOR U36016 ( .A(n36295), .B(p_input[3415]), .Z(n36297) );
  XOR U36017 ( .A(n36299), .B(n36300), .Z(n36295) );
  AND U36018 ( .A(n36301), .B(n36302), .Z(n36300) );
  XNOR U36019 ( .A(p_input[3446]), .B(n36299), .Z(n36302) );
  XOR U36020 ( .A(n36299), .B(p_input[3414]), .Z(n36301) );
  XOR U36021 ( .A(n36303), .B(n36304), .Z(n36299) );
  AND U36022 ( .A(n36305), .B(n36306), .Z(n36304) );
  XNOR U36023 ( .A(p_input[3445]), .B(n36303), .Z(n36306) );
  XOR U36024 ( .A(n36303), .B(p_input[3413]), .Z(n36305) );
  XOR U36025 ( .A(n36307), .B(n36308), .Z(n36303) );
  AND U36026 ( .A(n36309), .B(n36310), .Z(n36308) );
  XNOR U36027 ( .A(p_input[3444]), .B(n36307), .Z(n36310) );
  XOR U36028 ( .A(n36307), .B(p_input[3412]), .Z(n36309) );
  XOR U36029 ( .A(n36311), .B(n36312), .Z(n36307) );
  AND U36030 ( .A(n36313), .B(n36314), .Z(n36312) );
  XNOR U36031 ( .A(p_input[3443]), .B(n36311), .Z(n36314) );
  XOR U36032 ( .A(n36311), .B(p_input[3411]), .Z(n36313) );
  XOR U36033 ( .A(n36315), .B(n36316), .Z(n36311) );
  AND U36034 ( .A(n36317), .B(n36318), .Z(n36316) );
  XNOR U36035 ( .A(p_input[3442]), .B(n36315), .Z(n36318) );
  XOR U36036 ( .A(n36315), .B(p_input[3410]), .Z(n36317) );
  XOR U36037 ( .A(n36319), .B(n36320), .Z(n36315) );
  AND U36038 ( .A(n36321), .B(n36322), .Z(n36320) );
  XNOR U36039 ( .A(p_input[3441]), .B(n36319), .Z(n36322) );
  XOR U36040 ( .A(n36319), .B(p_input[3409]), .Z(n36321) );
  XOR U36041 ( .A(n36323), .B(n36324), .Z(n36319) );
  AND U36042 ( .A(n36325), .B(n36326), .Z(n36324) );
  XNOR U36043 ( .A(p_input[3440]), .B(n36323), .Z(n36326) );
  XOR U36044 ( .A(n36323), .B(p_input[3408]), .Z(n36325) );
  XOR U36045 ( .A(n36327), .B(n36328), .Z(n36323) );
  AND U36046 ( .A(n36329), .B(n36330), .Z(n36328) );
  XNOR U36047 ( .A(p_input[3439]), .B(n36327), .Z(n36330) );
  XOR U36048 ( .A(n36327), .B(p_input[3407]), .Z(n36329) );
  XOR U36049 ( .A(n36331), .B(n36332), .Z(n36327) );
  AND U36050 ( .A(n36333), .B(n36334), .Z(n36332) );
  XNOR U36051 ( .A(p_input[3438]), .B(n36331), .Z(n36334) );
  XOR U36052 ( .A(n36331), .B(p_input[3406]), .Z(n36333) );
  XOR U36053 ( .A(n36335), .B(n36336), .Z(n36331) );
  AND U36054 ( .A(n36337), .B(n36338), .Z(n36336) );
  XNOR U36055 ( .A(p_input[3437]), .B(n36335), .Z(n36338) );
  XOR U36056 ( .A(n36335), .B(p_input[3405]), .Z(n36337) );
  XOR U36057 ( .A(n36339), .B(n36340), .Z(n36335) );
  AND U36058 ( .A(n36341), .B(n36342), .Z(n36340) );
  XNOR U36059 ( .A(p_input[3436]), .B(n36339), .Z(n36342) );
  XOR U36060 ( .A(n36339), .B(p_input[3404]), .Z(n36341) );
  XOR U36061 ( .A(n36343), .B(n36344), .Z(n36339) );
  AND U36062 ( .A(n36345), .B(n36346), .Z(n36344) );
  XNOR U36063 ( .A(p_input[3435]), .B(n36343), .Z(n36346) );
  XOR U36064 ( .A(n36343), .B(p_input[3403]), .Z(n36345) );
  XOR U36065 ( .A(n36347), .B(n36348), .Z(n36343) );
  AND U36066 ( .A(n36349), .B(n36350), .Z(n36348) );
  XNOR U36067 ( .A(p_input[3434]), .B(n36347), .Z(n36350) );
  XOR U36068 ( .A(n36347), .B(p_input[3402]), .Z(n36349) );
  XOR U36069 ( .A(n36351), .B(n36352), .Z(n36347) );
  AND U36070 ( .A(n36353), .B(n36354), .Z(n36352) );
  XNOR U36071 ( .A(p_input[3433]), .B(n36351), .Z(n36354) );
  XOR U36072 ( .A(n36351), .B(p_input[3401]), .Z(n36353) );
  XOR U36073 ( .A(n36355), .B(n36356), .Z(n36351) );
  AND U36074 ( .A(n36357), .B(n36358), .Z(n36356) );
  XNOR U36075 ( .A(p_input[3432]), .B(n36355), .Z(n36358) );
  XOR U36076 ( .A(n36355), .B(p_input[3400]), .Z(n36357) );
  XOR U36077 ( .A(n36359), .B(n36360), .Z(n36355) );
  AND U36078 ( .A(n36361), .B(n36362), .Z(n36360) );
  XNOR U36079 ( .A(p_input[3431]), .B(n36359), .Z(n36362) );
  XOR U36080 ( .A(n36359), .B(p_input[3399]), .Z(n36361) );
  XOR U36081 ( .A(n36363), .B(n36364), .Z(n36359) );
  AND U36082 ( .A(n36365), .B(n36366), .Z(n36364) );
  XNOR U36083 ( .A(p_input[3430]), .B(n36363), .Z(n36366) );
  XOR U36084 ( .A(n36363), .B(p_input[3398]), .Z(n36365) );
  XOR U36085 ( .A(n36367), .B(n36368), .Z(n36363) );
  AND U36086 ( .A(n36369), .B(n36370), .Z(n36368) );
  XNOR U36087 ( .A(p_input[3429]), .B(n36367), .Z(n36370) );
  XOR U36088 ( .A(n36367), .B(p_input[3397]), .Z(n36369) );
  XOR U36089 ( .A(n36371), .B(n36372), .Z(n36367) );
  AND U36090 ( .A(n36373), .B(n36374), .Z(n36372) );
  XNOR U36091 ( .A(p_input[3428]), .B(n36371), .Z(n36374) );
  XOR U36092 ( .A(n36371), .B(p_input[3396]), .Z(n36373) );
  XOR U36093 ( .A(n36375), .B(n36376), .Z(n36371) );
  AND U36094 ( .A(n36377), .B(n36378), .Z(n36376) );
  XNOR U36095 ( .A(p_input[3427]), .B(n36375), .Z(n36378) );
  XOR U36096 ( .A(n36375), .B(p_input[3395]), .Z(n36377) );
  XOR U36097 ( .A(n36379), .B(n36380), .Z(n36375) );
  AND U36098 ( .A(n36381), .B(n36382), .Z(n36380) );
  XNOR U36099 ( .A(p_input[3426]), .B(n36379), .Z(n36382) );
  XOR U36100 ( .A(n36379), .B(p_input[3394]), .Z(n36381) );
  XNOR U36101 ( .A(n36383), .B(n36384), .Z(n36379) );
  AND U36102 ( .A(n36385), .B(n36386), .Z(n36384) );
  XOR U36103 ( .A(p_input[3425]), .B(n36383), .Z(n36386) );
  XNOR U36104 ( .A(p_input[3393]), .B(n36383), .Z(n36385) );
  AND U36105 ( .A(p_input[3424]), .B(n36387), .Z(n36383) );
  IV U36106 ( .A(p_input[3392]), .Z(n36387) );
  XNOR U36107 ( .A(p_input[3328]), .B(n36388), .Z(n35981) );
  AND U36108 ( .A(n720), .B(n36389), .Z(n36388) );
  XOR U36109 ( .A(p_input[3360]), .B(p_input[3328]), .Z(n36389) );
  XOR U36110 ( .A(n36390), .B(n36391), .Z(n720) );
  AND U36111 ( .A(n36392), .B(n36393), .Z(n36391) );
  XNOR U36112 ( .A(p_input[3391]), .B(n36390), .Z(n36393) );
  XOR U36113 ( .A(n36390), .B(p_input[3359]), .Z(n36392) );
  XOR U36114 ( .A(n36394), .B(n36395), .Z(n36390) );
  AND U36115 ( .A(n36396), .B(n36397), .Z(n36395) );
  XNOR U36116 ( .A(p_input[3390]), .B(n36394), .Z(n36397) );
  XNOR U36117 ( .A(n36394), .B(n35996), .Z(n36396) );
  IV U36118 ( .A(p_input[3358]), .Z(n35996) );
  XOR U36119 ( .A(n36398), .B(n36399), .Z(n36394) );
  AND U36120 ( .A(n36400), .B(n36401), .Z(n36399) );
  XNOR U36121 ( .A(p_input[3389]), .B(n36398), .Z(n36401) );
  XNOR U36122 ( .A(n36398), .B(n36005), .Z(n36400) );
  IV U36123 ( .A(p_input[3357]), .Z(n36005) );
  XOR U36124 ( .A(n36402), .B(n36403), .Z(n36398) );
  AND U36125 ( .A(n36404), .B(n36405), .Z(n36403) );
  XNOR U36126 ( .A(p_input[3388]), .B(n36402), .Z(n36405) );
  XNOR U36127 ( .A(n36402), .B(n36014), .Z(n36404) );
  IV U36128 ( .A(p_input[3356]), .Z(n36014) );
  XOR U36129 ( .A(n36406), .B(n36407), .Z(n36402) );
  AND U36130 ( .A(n36408), .B(n36409), .Z(n36407) );
  XNOR U36131 ( .A(p_input[3387]), .B(n36406), .Z(n36409) );
  XNOR U36132 ( .A(n36406), .B(n36023), .Z(n36408) );
  IV U36133 ( .A(p_input[3355]), .Z(n36023) );
  XOR U36134 ( .A(n36410), .B(n36411), .Z(n36406) );
  AND U36135 ( .A(n36412), .B(n36413), .Z(n36411) );
  XNOR U36136 ( .A(p_input[3386]), .B(n36410), .Z(n36413) );
  XNOR U36137 ( .A(n36410), .B(n36032), .Z(n36412) );
  IV U36138 ( .A(p_input[3354]), .Z(n36032) );
  XOR U36139 ( .A(n36414), .B(n36415), .Z(n36410) );
  AND U36140 ( .A(n36416), .B(n36417), .Z(n36415) );
  XNOR U36141 ( .A(p_input[3385]), .B(n36414), .Z(n36417) );
  XNOR U36142 ( .A(n36414), .B(n36041), .Z(n36416) );
  IV U36143 ( .A(p_input[3353]), .Z(n36041) );
  XOR U36144 ( .A(n36418), .B(n36419), .Z(n36414) );
  AND U36145 ( .A(n36420), .B(n36421), .Z(n36419) );
  XNOR U36146 ( .A(p_input[3384]), .B(n36418), .Z(n36421) );
  XNOR U36147 ( .A(n36418), .B(n36050), .Z(n36420) );
  IV U36148 ( .A(p_input[3352]), .Z(n36050) );
  XOR U36149 ( .A(n36422), .B(n36423), .Z(n36418) );
  AND U36150 ( .A(n36424), .B(n36425), .Z(n36423) );
  XNOR U36151 ( .A(p_input[3383]), .B(n36422), .Z(n36425) );
  XNOR U36152 ( .A(n36422), .B(n36059), .Z(n36424) );
  IV U36153 ( .A(p_input[3351]), .Z(n36059) );
  XOR U36154 ( .A(n36426), .B(n36427), .Z(n36422) );
  AND U36155 ( .A(n36428), .B(n36429), .Z(n36427) );
  XNOR U36156 ( .A(p_input[3382]), .B(n36426), .Z(n36429) );
  XNOR U36157 ( .A(n36426), .B(n36068), .Z(n36428) );
  IV U36158 ( .A(p_input[3350]), .Z(n36068) );
  XOR U36159 ( .A(n36430), .B(n36431), .Z(n36426) );
  AND U36160 ( .A(n36432), .B(n36433), .Z(n36431) );
  XNOR U36161 ( .A(p_input[3381]), .B(n36430), .Z(n36433) );
  XNOR U36162 ( .A(n36430), .B(n36077), .Z(n36432) );
  IV U36163 ( .A(p_input[3349]), .Z(n36077) );
  XOR U36164 ( .A(n36434), .B(n36435), .Z(n36430) );
  AND U36165 ( .A(n36436), .B(n36437), .Z(n36435) );
  XNOR U36166 ( .A(p_input[3380]), .B(n36434), .Z(n36437) );
  XNOR U36167 ( .A(n36434), .B(n36086), .Z(n36436) );
  IV U36168 ( .A(p_input[3348]), .Z(n36086) );
  XOR U36169 ( .A(n36438), .B(n36439), .Z(n36434) );
  AND U36170 ( .A(n36440), .B(n36441), .Z(n36439) );
  XNOR U36171 ( .A(p_input[3379]), .B(n36438), .Z(n36441) );
  XNOR U36172 ( .A(n36438), .B(n36095), .Z(n36440) );
  IV U36173 ( .A(p_input[3347]), .Z(n36095) );
  XOR U36174 ( .A(n36442), .B(n36443), .Z(n36438) );
  AND U36175 ( .A(n36444), .B(n36445), .Z(n36443) );
  XNOR U36176 ( .A(p_input[3378]), .B(n36442), .Z(n36445) );
  XNOR U36177 ( .A(n36442), .B(n36104), .Z(n36444) );
  IV U36178 ( .A(p_input[3346]), .Z(n36104) );
  XOR U36179 ( .A(n36446), .B(n36447), .Z(n36442) );
  AND U36180 ( .A(n36448), .B(n36449), .Z(n36447) );
  XNOR U36181 ( .A(p_input[3377]), .B(n36446), .Z(n36449) );
  XNOR U36182 ( .A(n36446), .B(n36113), .Z(n36448) );
  IV U36183 ( .A(p_input[3345]), .Z(n36113) );
  XOR U36184 ( .A(n36450), .B(n36451), .Z(n36446) );
  AND U36185 ( .A(n36452), .B(n36453), .Z(n36451) );
  XNOR U36186 ( .A(p_input[3376]), .B(n36450), .Z(n36453) );
  XNOR U36187 ( .A(n36450), .B(n36122), .Z(n36452) );
  IV U36188 ( .A(p_input[3344]), .Z(n36122) );
  XOR U36189 ( .A(n36454), .B(n36455), .Z(n36450) );
  AND U36190 ( .A(n36456), .B(n36457), .Z(n36455) );
  XNOR U36191 ( .A(p_input[3375]), .B(n36454), .Z(n36457) );
  XNOR U36192 ( .A(n36454), .B(n36131), .Z(n36456) );
  IV U36193 ( .A(p_input[3343]), .Z(n36131) );
  XOR U36194 ( .A(n36458), .B(n36459), .Z(n36454) );
  AND U36195 ( .A(n36460), .B(n36461), .Z(n36459) );
  XNOR U36196 ( .A(p_input[3374]), .B(n36458), .Z(n36461) );
  XNOR U36197 ( .A(n36458), .B(n36140), .Z(n36460) );
  IV U36198 ( .A(p_input[3342]), .Z(n36140) );
  XOR U36199 ( .A(n36462), .B(n36463), .Z(n36458) );
  AND U36200 ( .A(n36464), .B(n36465), .Z(n36463) );
  XNOR U36201 ( .A(p_input[3373]), .B(n36462), .Z(n36465) );
  XNOR U36202 ( .A(n36462), .B(n36149), .Z(n36464) );
  IV U36203 ( .A(p_input[3341]), .Z(n36149) );
  XOR U36204 ( .A(n36466), .B(n36467), .Z(n36462) );
  AND U36205 ( .A(n36468), .B(n36469), .Z(n36467) );
  XNOR U36206 ( .A(p_input[3372]), .B(n36466), .Z(n36469) );
  XNOR U36207 ( .A(n36466), .B(n36158), .Z(n36468) );
  IV U36208 ( .A(p_input[3340]), .Z(n36158) );
  XOR U36209 ( .A(n36470), .B(n36471), .Z(n36466) );
  AND U36210 ( .A(n36472), .B(n36473), .Z(n36471) );
  XNOR U36211 ( .A(p_input[3371]), .B(n36470), .Z(n36473) );
  XNOR U36212 ( .A(n36470), .B(n36167), .Z(n36472) );
  IV U36213 ( .A(p_input[3339]), .Z(n36167) );
  XOR U36214 ( .A(n36474), .B(n36475), .Z(n36470) );
  AND U36215 ( .A(n36476), .B(n36477), .Z(n36475) );
  XNOR U36216 ( .A(p_input[3370]), .B(n36474), .Z(n36477) );
  XNOR U36217 ( .A(n36474), .B(n36176), .Z(n36476) );
  IV U36218 ( .A(p_input[3338]), .Z(n36176) );
  XOR U36219 ( .A(n36478), .B(n36479), .Z(n36474) );
  AND U36220 ( .A(n36480), .B(n36481), .Z(n36479) );
  XNOR U36221 ( .A(p_input[3369]), .B(n36478), .Z(n36481) );
  XNOR U36222 ( .A(n36478), .B(n36185), .Z(n36480) );
  IV U36223 ( .A(p_input[3337]), .Z(n36185) );
  XOR U36224 ( .A(n36482), .B(n36483), .Z(n36478) );
  AND U36225 ( .A(n36484), .B(n36485), .Z(n36483) );
  XNOR U36226 ( .A(p_input[3368]), .B(n36482), .Z(n36485) );
  XNOR U36227 ( .A(n36482), .B(n36194), .Z(n36484) );
  IV U36228 ( .A(p_input[3336]), .Z(n36194) );
  XOR U36229 ( .A(n36486), .B(n36487), .Z(n36482) );
  AND U36230 ( .A(n36488), .B(n36489), .Z(n36487) );
  XNOR U36231 ( .A(p_input[3367]), .B(n36486), .Z(n36489) );
  XNOR U36232 ( .A(n36486), .B(n36203), .Z(n36488) );
  IV U36233 ( .A(p_input[3335]), .Z(n36203) );
  XOR U36234 ( .A(n36490), .B(n36491), .Z(n36486) );
  AND U36235 ( .A(n36492), .B(n36493), .Z(n36491) );
  XNOR U36236 ( .A(p_input[3366]), .B(n36490), .Z(n36493) );
  XNOR U36237 ( .A(n36490), .B(n36212), .Z(n36492) );
  IV U36238 ( .A(p_input[3334]), .Z(n36212) );
  XOR U36239 ( .A(n36494), .B(n36495), .Z(n36490) );
  AND U36240 ( .A(n36496), .B(n36497), .Z(n36495) );
  XNOR U36241 ( .A(p_input[3365]), .B(n36494), .Z(n36497) );
  XNOR U36242 ( .A(n36494), .B(n36221), .Z(n36496) );
  IV U36243 ( .A(p_input[3333]), .Z(n36221) );
  XOR U36244 ( .A(n36498), .B(n36499), .Z(n36494) );
  AND U36245 ( .A(n36500), .B(n36501), .Z(n36499) );
  XNOR U36246 ( .A(p_input[3364]), .B(n36498), .Z(n36501) );
  XNOR U36247 ( .A(n36498), .B(n36230), .Z(n36500) );
  IV U36248 ( .A(p_input[3332]), .Z(n36230) );
  XOR U36249 ( .A(n36502), .B(n36503), .Z(n36498) );
  AND U36250 ( .A(n36504), .B(n36505), .Z(n36503) );
  XNOR U36251 ( .A(p_input[3363]), .B(n36502), .Z(n36505) );
  XNOR U36252 ( .A(n36502), .B(n36239), .Z(n36504) );
  IV U36253 ( .A(p_input[3331]), .Z(n36239) );
  XOR U36254 ( .A(n36506), .B(n36507), .Z(n36502) );
  AND U36255 ( .A(n36508), .B(n36509), .Z(n36507) );
  XNOR U36256 ( .A(p_input[3362]), .B(n36506), .Z(n36509) );
  XNOR U36257 ( .A(n36506), .B(n36248), .Z(n36508) );
  IV U36258 ( .A(p_input[3330]), .Z(n36248) );
  XNOR U36259 ( .A(n36510), .B(n36511), .Z(n36506) );
  AND U36260 ( .A(n36512), .B(n36513), .Z(n36511) );
  XOR U36261 ( .A(p_input[3361]), .B(n36510), .Z(n36513) );
  XNOR U36262 ( .A(p_input[3329]), .B(n36510), .Z(n36512) );
  AND U36263 ( .A(p_input[3360]), .B(n36514), .Z(n36510) );
  IV U36264 ( .A(p_input[3328]), .Z(n36514) );
  XOR U36265 ( .A(n36515), .B(n36516), .Z(n34693) );
  AND U36266 ( .A(n876), .B(n36517), .Z(n36516) );
  XNOR U36267 ( .A(n36518), .B(n36515), .Z(n36517) );
  XOR U36268 ( .A(n36519), .B(n36520), .Z(n876) );
  AND U36269 ( .A(n36521), .B(n36522), .Z(n36520) );
  XOR U36270 ( .A(n36519), .B(n34708), .Z(n36522) );
  XNOR U36271 ( .A(n36523), .B(n36524), .Z(n34708) );
  AND U36272 ( .A(n36525), .B(n579), .Z(n36524) );
  AND U36273 ( .A(n36523), .B(n36526), .Z(n36525) );
  XNOR U36274 ( .A(n34705), .B(n36519), .Z(n36521) );
  XOR U36275 ( .A(n36527), .B(n36528), .Z(n34705) );
  AND U36276 ( .A(n36529), .B(n576), .Z(n36528) );
  NOR U36277 ( .A(n36527), .B(n36530), .Z(n36529) );
  XOR U36278 ( .A(n36531), .B(n36532), .Z(n36519) );
  AND U36279 ( .A(n36533), .B(n36534), .Z(n36532) );
  XOR U36280 ( .A(n36531), .B(n34720), .Z(n36534) );
  XOR U36281 ( .A(n36535), .B(n36536), .Z(n34720) );
  AND U36282 ( .A(n579), .B(n36537), .Z(n36536) );
  XOR U36283 ( .A(n36538), .B(n36535), .Z(n36537) );
  XNOR U36284 ( .A(n34717), .B(n36531), .Z(n36533) );
  XOR U36285 ( .A(n36539), .B(n36540), .Z(n34717) );
  AND U36286 ( .A(n576), .B(n36541), .Z(n36540) );
  XOR U36287 ( .A(n36542), .B(n36539), .Z(n36541) );
  XOR U36288 ( .A(n36543), .B(n36544), .Z(n36531) );
  AND U36289 ( .A(n36545), .B(n36546), .Z(n36544) );
  XOR U36290 ( .A(n36543), .B(n34732), .Z(n36546) );
  XOR U36291 ( .A(n36547), .B(n36548), .Z(n34732) );
  AND U36292 ( .A(n579), .B(n36549), .Z(n36548) );
  XOR U36293 ( .A(n36550), .B(n36547), .Z(n36549) );
  XNOR U36294 ( .A(n34729), .B(n36543), .Z(n36545) );
  XOR U36295 ( .A(n36551), .B(n36552), .Z(n34729) );
  AND U36296 ( .A(n576), .B(n36553), .Z(n36552) );
  XOR U36297 ( .A(n36554), .B(n36551), .Z(n36553) );
  XOR U36298 ( .A(n36555), .B(n36556), .Z(n36543) );
  AND U36299 ( .A(n36557), .B(n36558), .Z(n36556) );
  XOR U36300 ( .A(n36555), .B(n34744), .Z(n36558) );
  XOR U36301 ( .A(n36559), .B(n36560), .Z(n34744) );
  AND U36302 ( .A(n579), .B(n36561), .Z(n36560) );
  XOR U36303 ( .A(n36562), .B(n36559), .Z(n36561) );
  XNOR U36304 ( .A(n34741), .B(n36555), .Z(n36557) );
  XOR U36305 ( .A(n36563), .B(n36564), .Z(n34741) );
  AND U36306 ( .A(n576), .B(n36565), .Z(n36564) );
  XOR U36307 ( .A(n36566), .B(n36563), .Z(n36565) );
  XOR U36308 ( .A(n36567), .B(n36568), .Z(n36555) );
  AND U36309 ( .A(n36569), .B(n36570), .Z(n36568) );
  XOR U36310 ( .A(n36567), .B(n34756), .Z(n36570) );
  XOR U36311 ( .A(n36571), .B(n36572), .Z(n34756) );
  AND U36312 ( .A(n579), .B(n36573), .Z(n36572) );
  XOR U36313 ( .A(n36574), .B(n36571), .Z(n36573) );
  XNOR U36314 ( .A(n34753), .B(n36567), .Z(n36569) );
  XOR U36315 ( .A(n36575), .B(n36576), .Z(n34753) );
  AND U36316 ( .A(n576), .B(n36577), .Z(n36576) );
  XOR U36317 ( .A(n36578), .B(n36575), .Z(n36577) );
  XOR U36318 ( .A(n36579), .B(n36580), .Z(n36567) );
  AND U36319 ( .A(n36581), .B(n36582), .Z(n36580) );
  XOR U36320 ( .A(n36579), .B(n34768), .Z(n36582) );
  XOR U36321 ( .A(n36583), .B(n36584), .Z(n34768) );
  AND U36322 ( .A(n579), .B(n36585), .Z(n36584) );
  XOR U36323 ( .A(n36586), .B(n36583), .Z(n36585) );
  XNOR U36324 ( .A(n34765), .B(n36579), .Z(n36581) );
  XOR U36325 ( .A(n36587), .B(n36588), .Z(n34765) );
  AND U36326 ( .A(n576), .B(n36589), .Z(n36588) );
  XOR U36327 ( .A(n36590), .B(n36587), .Z(n36589) );
  XOR U36328 ( .A(n36591), .B(n36592), .Z(n36579) );
  AND U36329 ( .A(n36593), .B(n36594), .Z(n36592) );
  XOR U36330 ( .A(n36591), .B(n34780), .Z(n36594) );
  XOR U36331 ( .A(n36595), .B(n36596), .Z(n34780) );
  AND U36332 ( .A(n579), .B(n36597), .Z(n36596) );
  XOR U36333 ( .A(n36598), .B(n36595), .Z(n36597) );
  XNOR U36334 ( .A(n34777), .B(n36591), .Z(n36593) );
  XOR U36335 ( .A(n36599), .B(n36600), .Z(n34777) );
  AND U36336 ( .A(n576), .B(n36601), .Z(n36600) );
  XOR U36337 ( .A(n36602), .B(n36599), .Z(n36601) );
  XOR U36338 ( .A(n36603), .B(n36604), .Z(n36591) );
  AND U36339 ( .A(n36605), .B(n36606), .Z(n36604) );
  XOR U36340 ( .A(n36603), .B(n34792), .Z(n36606) );
  XOR U36341 ( .A(n36607), .B(n36608), .Z(n34792) );
  AND U36342 ( .A(n579), .B(n36609), .Z(n36608) );
  XOR U36343 ( .A(n36610), .B(n36607), .Z(n36609) );
  XNOR U36344 ( .A(n34789), .B(n36603), .Z(n36605) );
  XOR U36345 ( .A(n36611), .B(n36612), .Z(n34789) );
  AND U36346 ( .A(n576), .B(n36613), .Z(n36612) );
  XOR U36347 ( .A(n36614), .B(n36611), .Z(n36613) );
  XOR U36348 ( .A(n36615), .B(n36616), .Z(n36603) );
  AND U36349 ( .A(n36617), .B(n36618), .Z(n36616) );
  XOR U36350 ( .A(n36615), .B(n34804), .Z(n36618) );
  XOR U36351 ( .A(n36619), .B(n36620), .Z(n34804) );
  AND U36352 ( .A(n579), .B(n36621), .Z(n36620) );
  XOR U36353 ( .A(n36622), .B(n36619), .Z(n36621) );
  XNOR U36354 ( .A(n34801), .B(n36615), .Z(n36617) );
  XOR U36355 ( .A(n36623), .B(n36624), .Z(n34801) );
  AND U36356 ( .A(n576), .B(n36625), .Z(n36624) );
  XOR U36357 ( .A(n36626), .B(n36623), .Z(n36625) );
  XOR U36358 ( .A(n36627), .B(n36628), .Z(n36615) );
  AND U36359 ( .A(n36629), .B(n36630), .Z(n36628) );
  XOR U36360 ( .A(n36627), .B(n34816), .Z(n36630) );
  XOR U36361 ( .A(n36631), .B(n36632), .Z(n34816) );
  AND U36362 ( .A(n579), .B(n36633), .Z(n36632) );
  XOR U36363 ( .A(n36634), .B(n36631), .Z(n36633) );
  XNOR U36364 ( .A(n34813), .B(n36627), .Z(n36629) );
  XOR U36365 ( .A(n36635), .B(n36636), .Z(n34813) );
  AND U36366 ( .A(n576), .B(n36637), .Z(n36636) );
  XOR U36367 ( .A(n36638), .B(n36635), .Z(n36637) );
  XOR U36368 ( .A(n36639), .B(n36640), .Z(n36627) );
  AND U36369 ( .A(n36641), .B(n36642), .Z(n36640) );
  XOR U36370 ( .A(n36639), .B(n34828), .Z(n36642) );
  XOR U36371 ( .A(n36643), .B(n36644), .Z(n34828) );
  AND U36372 ( .A(n579), .B(n36645), .Z(n36644) );
  XOR U36373 ( .A(n36646), .B(n36643), .Z(n36645) );
  XNOR U36374 ( .A(n34825), .B(n36639), .Z(n36641) );
  XOR U36375 ( .A(n36647), .B(n36648), .Z(n34825) );
  AND U36376 ( .A(n576), .B(n36649), .Z(n36648) );
  XOR U36377 ( .A(n36650), .B(n36647), .Z(n36649) );
  XOR U36378 ( .A(n36651), .B(n36652), .Z(n36639) );
  AND U36379 ( .A(n36653), .B(n36654), .Z(n36652) );
  XOR U36380 ( .A(n36651), .B(n34840), .Z(n36654) );
  XOR U36381 ( .A(n36655), .B(n36656), .Z(n34840) );
  AND U36382 ( .A(n579), .B(n36657), .Z(n36656) );
  XOR U36383 ( .A(n36658), .B(n36655), .Z(n36657) );
  XNOR U36384 ( .A(n34837), .B(n36651), .Z(n36653) );
  XOR U36385 ( .A(n36659), .B(n36660), .Z(n34837) );
  AND U36386 ( .A(n576), .B(n36661), .Z(n36660) );
  XOR U36387 ( .A(n36662), .B(n36659), .Z(n36661) );
  XOR U36388 ( .A(n36663), .B(n36664), .Z(n36651) );
  AND U36389 ( .A(n36665), .B(n36666), .Z(n36664) );
  XOR U36390 ( .A(n36663), .B(n34852), .Z(n36666) );
  XOR U36391 ( .A(n36667), .B(n36668), .Z(n34852) );
  AND U36392 ( .A(n579), .B(n36669), .Z(n36668) );
  XOR U36393 ( .A(n36670), .B(n36667), .Z(n36669) );
  XNOR U36394 ( .A(n34849), .B(n36663), .Z(n36665) );
  XOR U36395 ( .A(n36671), .B(n36672), .Z(n34849) );
  AND U36396 ( .A(n576), .B(n36673), .Z(n36672) );
  XOR U36397 ( .A(n36674), .B(n36671), .Z(n36673) );
  XOR U36398 ( .A(n36675), .B(n36676), .Z(n36663) );
  AND U36399 ( .A(n36677), .B(n36678), .Z(n36676) );
  XOR U36400 ( .A(n36675), .B(n34864), .Z(n36678) );
  XOR U36401 ( .A(n36679), .B(n36680), .Z(n34864) );
  AND U36402 ( .A(n579), .B(n36681), .Z(n36680) );
  XOR U36403 ( .A(n36682), .B(n36679), .Z(n36681) );
  XNOR U36404 ( .A(n34861), .B(n36675), .Z(n36677) );
  XOR U36405 ( .A(n36683), .B(n36684), .Z(n34861) );
  AND U36406 ( .A(n576), .B(n36685), .Z(n36684) );
  XOR U36407 ( .A(n36686), .B(n36683), .Z(n36685) );
  XOR U36408 ( .A(n36687), .B(n36688), .Z(n36675) );
  AND U36409 ( .A(n36689), .B(n36690), .Z(n36688) );
  XOR U36410 ( .A(n36687), .B(n34876), .Z(n36690) );
  XOR U36411 ( .A(n36691), .B(n36692), .Z(n34876) );
  AND U36412 ( .A(n579), .B(n36693), .Z(n36692) );
  XOR U36413 ( .A(n36694), .B(n36691), .Z(n36693) );
  XNOR U36414 ( .A(n34873), .B(n36687), .Z(n36689) );
  XOR U36415 ( .A(n36695), .B(n36696), .Z(n34873) );
  AND U36416 ( .A(n576), .B(n36697), .Z(n36696) );
  XOR U36417 ( .A(n36698), .B(n36695), .Z(n36697) );
  XOR U36418 ( .A(n36699), .B(n36700), .Z(n36687) );
  AND U36419 ( .A(n36701), .B(n36702), .Z(n36700) );
  XOR U36420 ( .A(n36699), .B(n34888), .Z(n36702) );
  XOR U36421 ( .A(n36703), .B(n36704), .Z(n34888) );
  AND U36422 ( .A(n579), .B(n36705), .Z(n36704) );
  XOR U36423 ( .A(n36706), .B(n36703), .Z(n36705) );
  XNOR U36424 ( .A(n34885), .B(n36699), .Z(n36701) );
  XOR U36425 ( .A(n36707), .B(n36708), .Z(n34885) );
  AND U36426 ( .A(n576), .B(n36709), .Z(n36708) );
  XOR U36427 ( .A(n36710), .B(n36707), .Z(n36709) );
  XOR U36428 ( .A(n36711), .B(n36712), .Z(n36699) );
  AND U36429 ( .A(n36713), .B(n36714), .Z(n36712) );
  XOR U36430 ( .A(n36711), .B(n34900), .Z(n36714) );
  XOR U36431 ( .A(n36715), .B(n36716), .Z(n34900) );
  AND U36432 ( .A(n579), .B(n36717), .Z(n36716) );
  XOR U36433 ( .A(n36718), .B(n36715), .Z(n36717) );
  XNOR U36434 ( .A(n34897), .B(n36711), .Z(n36713) );
  XOR U36435 ( .A(n36719), .B(n36720), .Z(n34897) );
  AND U36436 ( .A(n576), .B(n36721), .Z(n36720) );
  XOR U36437 ( .A(n36722), .B(n36719), .Z(n36721) );
  XOR U36438 ( .A(n36723), .B(n36724), .Z(n36711) );
  AND U36439 ( .A(n36725), .B(n36726), .Z(n36724) );
  XOR U36440 ( .A(n36723), .B(n34912), .Z(n36726) );
  XOR U36441 ( .A(n36727), .B(n36728), .Z(n34912) );
  AND U36442 ( .A(n579), .B(n36729), .Z(n36728) );
  XOR U36443 ( .A(n36730), .B(n36727), .Z(n36729) );
  XNOR U36444 ( .A(n34909), .B(n36723), .Z(n36725) );
  XOR U36445 ( .A(n36731), .B(n36732), .Z(n34909) );
  AND U36446 ( .A(n576), .B(n36733), .Z(n36732) );
  XOR U36447 ( .A(n36734), .B(n36731), .Z(n36733) );
  XOR U36448 ( .A(n36735), .B(n36736), .Z(n36723) );
  AND U36449 ( .A(n36737), .B(n36738), .Z(n36736) );
  XOR U36450 ( .A(n36735), .B(n34924), .Z(n36738) );
  XOR U36451 ( .A(n36739), .B(n36740), .Z(n34924) );
  AND U36452 ( .A(n579), .B(n36741), .Z(n36740) );
  XOR U36453 ( .A(n36742), .B(n36739), .Z(n36741) );
  XNOR U36454 ( .A(n34921), .B(n36735), .Z(n36737) );
  XOR U36455 ( .A(n36743), .B(n36744), .Z(n34921) );
  AND U36456 ( .A(n576), .B(n36745), .Z(n36744) );
  XOR U36457 ( .A(n36746), .B(n36743), .Z(n36745) );
  XOR U36458 ( .A(n36747), .B(n36748), .Z(n36735) );
  AND U36459 ( .A(n36749), .B(n36750), .Z(n36748) );
  XOR U36460 ( .A(n36747), .B(n34936), .Z(n36750) );
  XOR U36461 ( .A(n36751), .B(n36752), .Z(n34936) );
  AND U36462 ( .A(n579), .B(n36753), .Z(n36752) );
  XOR U36463 ( .A(n36754), .B(n36751), .Z(n36753) );
  XNOR U36464 ( .A(n34933), .B(n36747), .Z(n36749) );
  XOR U36465 ( .A(n36755), .B(n36756), .Z(n34933) );
  AND U36466 ( .A(n576), .B(n36757), .Z(n36756) );
  XOR U36467 ( .A(n36758), .B(n36755), .Z(n36757) );
  XOR U36468 ( .A(n36759), .B(n36760), .Z(n36747) );
  AND U36469 ( .A(n36761), .B(n36762), .Z(n36760) );
  XOR U36470 ( .A(n36759), .B(n34948), .Z(n36762) );
  XOR U36471 ( .A(n36763), .B(n36764), .Z(n34948) );
  AND U36472 ( .A(n579), .B(n36765), .Z(n36764) );
  XOR U36473 ( .A(n36766), .B(n36763), .Z(n36765) );
  XNOR U36474 ( .A(n34945), .B(n36759), .Z(n36761) );
  XOR U36475 ( .A(n36767), .B(n36768), .Z(n34945) );
  AND U36476 ( .A(n576), .B(n36769), .Z(n36768) );
  XOR U36477 ( .A(n36770), .B(n36767), .Z(n36769) );
  XOR U36478 ( .A(n36771), .B(n36772), .Z(n36759) );
  AND U36479 ( .A(n36773), .B(n36774), .Z(n36772) );
  XOR U36480 ( .A(n36771), .B(n34960), .Z(n36774) );
  XOR U36481 ( .A(n36775), .B(n36776), .Z(n34960) );
  AND U36482 ( .A(n579), .B(n36777), .Z(n36776) );
  XOR U36483 ( .A(n36778), .B(n36775), .Z(n36777) );
  XNOR U36484 ( .A(n34957), .B(n36771), .Z(n36773) );
  XOR U36485 ( .A(n36779), .B(n36780), .Z(n34957) );
  AND U36486 ( .A(n576), .B(n36781), .Z(n36780) );
  XOR U36487 ( .A(n36782), .B(n36779), .Z(n36781) );
  XOR U36488 ( .A(n36783), .B(n36784), .Z(n36771) );
  AND U36489 ( .A(n36785), .B(n36786), .Z(n36784) );
  XOR U36490 ( .A(n36783), .B(n34972), .Z(n36786) );
  XOR U36491 ( .A(n36787), .B(n36788), .Z(n34972) );
  AND U36492 ( .A(n579), .B(n36789), .Z(n36788) );
  XOR U36493 ( .A(n36790), .B(n36787), .Z(n36789) );
  XNOR U36494 ( .A(n34969), .B(n36783), .Z(n36785) );
  XOR U36495 ( .A(n36791), .B(n36792), .Z(n34969) );
  AND U36496 ( .A(n576), .B(n36793), .Z(n36792) );
  XOR U36497 ( .A(n36794), .B(n36791), .Z(n36793) );
  XOR U36498 ( .A(n36795), .B(n36796), .Z(n36783) );
  AND U36499 ( .A(n36797), .B(n36798), .Z(n36796) );
  XOR U36500 ( .A(n36795), .B(n34984), .Z(n36798) );
  XOR U36501 ( .A(n36799), .B(n36800), .Z(n34984) );
  AND U36502 ( .A(n579), .B(n36801), .Z(n36800) );
  XOR U36503 ( .A(n36802), .B(n36799), .Z(n36801) );
  XNOR U36504 ( .A(n34981), .B(n36795), .Z(n36797) );
  XOR U36505 ( .A(n36803), .B(n36804), .Z(n34981) );
  AND U36506 ( .A(n576), .B(n36805), .Z(n36804) );
  XOR U36507 ( .A(n36806), .B(n36803), .Z(n36805) );
  XOR U36508 ( .A(n36807), .B(n36808), .Z(n36795) );
  AND U36509 ( .A(n36809), .B(n36810), .Z(n36808) );
  XOR U36510 ( .A(n36807), .B(n34996), .Z(n36810) );
  XOR U36511 ( .A(n36811), .B(n36812), .Z(n34996) );
  AND U36512 ( .A(n579), .B(n36813), .Z(n36812) );
  XOR U36513 ( .A(n36814), .B(n36811), .Z(n36813) );
  XNOR U36514 ( .A(n34993), .B(n36807), .Z(n36809) );
  XOR U36515 ( .A(n36815), .B(n36816), .Z(n34993) );
  AND U36516 ( .A(n576), .B(n36817), .Z(n36816) );
  XOR U36517 ( .A(n36818), .B(n36815), .Z(n36817) );
  XOR U36518 ( .A(n36819), .B(n36820), .Z(n36807) );
  AND U36519 ( .A(n36821), .B(n36822), .Z(n36820) );
  XOR U36520 ( .A(n36819), .B(n35008), .Z(n36822) );
  XOR U36521 ( .A(n36823), .B(n36824), .Z(n35008) );
  AND U36522 ( .A(n579), .B(n36825), .Z(n36824) );
  XOR U36523 ( .A(n36826), .B(n36823), .Z(n36825) );
  XNOR U36524 ( .A(n35005), .B(n36819), .Z(n36821) );
  XOR U36525 ( .A(n36827), .B(n36828), .Z(n35005) );
  AND U36526 ( .A(n576), .B(n36829), .Z(n36828) );
  XOR U36527 ( .A(n36830), .B(n36827), .Z(n36829) );
  XOR U36528 ( .A(n36831), .B(n36832), .Z(n36819) );
  AND U36529 ( .A(n36833), .B(n36834), .Z(n36832) );
  XOR U36530 ( .A(n36831), .B(n35020), .Z(n36834) );
  XOR U36531 ( .A(n36835), .B(n36836), .Z(n35020) );
  AND U36532 ( .A(n579), .B(n36837), .Z(n36836) );
  XOR U36533 ( .A(n36838), .B(n36835), .Z(n36837) );
  XNOR U36534 ( .A(n35017), .B(n36831), .Z(n36833) );
  XOR U36535 ( .A(n36839), .B(n36840), .Z(n35017) );
  AND U36536 ( .A(n576), .B(n36841), .Z(n36840) );
  XOR U36537 ( .A(n36842), .B(n36839), .Z(n36841) );
  XOR U36538 ( .A(n36843), .B(n36844), .Z(n36831) );
  AND U36539 ( .A(n36845), .B(n36846), .Z(n36844) );
  XOR U36540 ( .A(n36843), .B(n35032), .Z(n36846) );
  XOR U36541 ( .A(n36847), .B(n36848), .Z(n35032) );
  AND U36542 ( .A(n579), .B(n36849), .Z(n36848) );
  XOR U36543 ( .A(n36850), .B(n36847), .Z(n36849) );
  XNOR U36544 ( .A(n35029), .B(n36843), .Z(n36845) );
  XOR U36545 ( .A(n36851), .B(n36852), .Z(n35029) );
  AND U36546 ( .A(n576), .B(n36853), .Z(n36852) );
  XOR U36547 ( .A(n36854), .B(n36851), .Z(n36853) );
  XOR U36548 ( .A(n36855), .B(n36856), .Z(n36843) );
  AND U36549 ( .A(n36857), .B(n36858), .Z(n36856) );
  XOR U36550 ( .A(n36855), .B(n35044), .Z(n36858) );
  XOR U36551 ( .A(n36859), .B(n36860), .Z(n35044) );
  AND U36552 ( .A(n579), .B(n36861), .Z(n36860) );
  XOR U36553 ( .A(n36862), .B(n36859), .Z(n36861) );
  XNOR U36554 ( .A(n35041), .B(n36855), .Z(n36857) );
  XOR U36555 ( .A(n36863), .B(n36864), .Z(n35041) );
  AND U36556 ( .A(n576), .B(n36865), .Z(n36864) );
  XOR U36557 ( .A(n36866), .B(n36863), .Z(n36865) );
  XOR U36558 ( .A(n36867), .B(n36868), .Z(n36855) );
  AND U36559 ( .A(n36869), .B(n36870), .Z(n36868) );
  XOR U36560 ( .A(n36867), .B(n35056), .Z(n36870) );
  XOR U36561 ( .A(n36871), .B(n36872), .Z(n35056) );
  AND U36562 ( .A(n579), .B(n36873), .Z(n36872) );
  XOR U36563 ( .A(n36874), .B(n36871), .Z(n36873) );
  XNOR U36564 ( .A(n35053), .B(n36867), .Z(n36869) );
  XOR U36565 ( .A(n36875), .B(n36876), .Z(n35053) );
  AND U36566 ( .A(n576), .B(n36877), .Z(n36876) );
  XOR U36567 ( .A(n36878), .B(n36875), .Z(n36877) );
  XOR U36568 ( .A(n36879), .B(n36880), .Z(n36867) );
  AND U36569 ( .A(n36881), .B(n36882), .Z(n36880) );
  XNOR U36570 ( .A(n36883), .B(n35069), .Z(n36882) );
  XOR U36571 ( .A(n36884), .B(n36885), .Z(n35069) );
  AND U36572 ( .A(n579), .B(n36886), .Z(n36885) );
  XOR U36573 ( .A(n36884), .B(n36887), .Z(n36886) );
  XNOR U36574 ( .A(n35066), .B(n36879), .Z(n36881) );
  XOR U36575 ( .A(n36888), .B(n36889), .Z(n35066) );
  AND U36576 ( .A(n576), .B(n36890), .Z(n36889) );
  XOR U36577 ( .A(n36888), .B(n36891), .Z(n36890) );
  IV U36578 ( .A(n36883), .Z(n36879) );
  AND U36579 ( .A(n36515), .B(n36518), .Z(n36883) );
  XNOR U36580 ( .A(n36892), .B(n36893), .Z(n36518) );
  AND U36581 ( .A(n579), .B(n36894), .Z(n36893) );
  XNOR U36582 ( .A(n36895), .B(n36892), .Z(n36894) );
  XOR U36583 ( .A(n36896), .B(n36897), .Z(n579) );
  AND U36584 ( .A(n36898), .B(n36899), .Z(n36897) );
  XOR U36585 ( .A(n36526), .B(n36896), .Z(n36899) );
  IV U36586 ( .A(n36900), .Z(n36526) );
  AND U36587 ( .A(p_input[3327]), .B(p_input[3295]), .Z(n36900) );
  XOR U36588 ( .A(n36896), .B(n36523), .Z(n36898) );
  AND U36589 ( .A(p_input[3231]), .B(p_input[3263]), .Z(n36523) );
  XOR U36590 ( .A(n36901), .B(n36902), .Z(n36896) );
  AND U36591 ( .A(n36903), .B(n36904), .Z(n36902) );
  XOR U36592 ( .A(n36901), .B(n36538), .Z(n36904) );
  XNOR U36593 ( .A(p_input[3294]), .B(n36905), .Z(n36538) );
  AND U36594 ( .A(n731), .B(n36906), .Z(n36905) );
  XOR U36595 ( .A(p_input[3326]), .B(p_input[3294]), .Z(n36906) );
  XNOR U36596 ( .A(n36535), .B(n36901), .Z(n36903) );
  XOR U36597 ( .A(n36907), .B(n36908), .Z(n36535) );
  AND U36598 ( .A(n729), .B(n36909), .Z(n36908) );
  XOR U36599 ( .A(p_input[3262]), .B(p_input[3230]), .Z(n36909) );
  XOR U36600 ( .A(n36910), .B(n36911), .Z(n36901) );
  AND U36601 ( .A(n36912), .B(n36913), .Z(n36911) );
  XOR U36602 ( .A(n36910), .B(n36550), .Z(n36913) );
  XNOR U36603 ( .A(p_input[3293]), .B(n36914), .Z(n36550) );
  AND U36604 ( .A(n731), .B(n36915), .Z(n36914) );
  XOR U36605 ( .A(p_input[3325]), .B(p_input[3293]), .Z(n36915) );
  XNOR U36606 ( .A(n36547), .B(n36910), .Z(n36912) );
  XOR U36607 ( .A(n36916), .B(n36917), .Z(n36547) );
  AND U36608 ( .A(n729), .B(n36918), .Z(n36917) );
  XOR U36609 ( .A(p_input[3261]), .B(p_input[3229]), .Z(n36918) );
  XOR U36610 ( .A(n36919), .B(n36920), .Z(n36910) );
  AND U36611 ( .A(n36921), .B(n36922), .Z(n36920) );
  XOR U36612 ( .A(n36919), .B(n36562), .Z(n36922) );
  XNOR U36613 ( .A(p_input[3292]), .B(n36923), .Z(n36562) );
  AND U36614 ( .A(n731), .B(n36924), .Z(n36923) );
  XOR U36615 ( .A(p_input[3324]), .B(p_input[3292]), .Z(n36924) );
  XNOR U36616 ( .A(n36559), .B(n36919), .Z(n36921) );
  XOR U36617 ( .A(n36925), .B(n36926), .Z(n36559) );
  AND U36618 ( .A(n729), .B(n36927), .Z(n36926) );
  XOR U36619 ( .A(p_input[3260]), .B(p_input[3228]), .Z(n36927) );
  XOR U36620 ( .A(n36928), .B(n36929), .Z(n36919) );
  AND U36621 ( .A(n36930), .B(n36931), .Z(n36929) );
  XOR U36622 ( .A(n36928), .B(n36574), .Z(n36931) );
  XNOR U36623 ( .A(p_input[3291]), .B(n36932), .Z(n36574) );
  AND U36624 ( .A(n731), .B(n36933), .Z(n36932) );
  XOR U36625 ( .A(p_input[3323]), .B(p_input[3291]), .Z(n36933) );
  XNOR U36626 ( .A(n36571), .B(n36928), .Z(n36930) );
  XOR U36627 ( .A(n36934), .B(n36935), .Z(n36571) );
  AND U36628 ( .A(n729), .B(n36936), .Z(n36935) );
  XOR U36629 ( .A(p_input[3259]), .B(p_input[3227]), .Z(n36936) );
  XOR U36630 ( .A(n36937), .B(n36938), .Z(n36928) );
  AND U36631 ( .A(n36939), .B(n36940), .Z(n36938) );
  XOR U36632 ( .A(n36937), .B(n36586), .Z(n36940) );
  XNOR U36633 ( .A(p_input[3290]), .B(n36941), .Z(n36586) );
  AND U36634 ( .A(n731), .B(n36942), .Z(n36941) );
  XOR U36635 ( .A(p_input[3322]), .B(p_input[3290]), .Z(n36942) );
  XNOR U36636 ( .A(n36583), .B(n36937), .Z(n36939) );
  XOR U36637 ( .A(n36943), .B(n36944), .Z(n36583) );
  AND U36638 ( .A(n729), .B(n36945), .Z(n36944) );
  XOR U36639 ( .A(p_input[3258]), .B(p_input[3226]), .Z(n36945) );
  XOR U36640 ( .A(n36946), .B(n36947), .Z(n36937) );
  AND U36641 ( .A(n36948), .B(n36949), .Z(n36947) );
  XOR U36642 ( .A(n36946), .B(n36598), .Z(n36949) );
  XNOR U36643 ( .A(p_input[3289]), .B(n36950), .Z(n36598) );
  AND U36644 ( .A(n731), .B(n36951), .Z(n36950) );
  XOR U36645 ( .A(p_input[3321]), .B(p_input[3289]), .Z(n36951) );
  XNOR U36646 ( .A(n36595), .B(n36946), .Z(n36948) );
  XOR U36647 ( .A(n36952), .B(n36953), .Z(n36595) );
  AND U36648 ( .A(n729), .B(n36954), .Z(n36953) );
  XOR U36649 ( .A(p_input[3257]), .B(p_input[3225]), .Z(n36954) );
  XOR U36650 ( .A(n36955), .B(n36956), .Z(n36946) );
  AND U36651 ( .A(n36957), .B(n36958), .Z(n36956) );
  XOR U36652 ( .A(n36955), .B(n36610), .Z(n36958) );
  XNOR U36653 ( .A(p_input[3288]), .B(n36959), .Z(n36610) );
  AND U36654 ( .A(n731), .B(n36960), .Z(n36959) );
  XOR U36655 ( .A(p_input[3320]), .B(p_input[3288]), .Z(n36960) );
  XNOR U36656 ( .A(n36607), .B(n36955), .Z(n36957) );
  XOR U36657 ( .A(n36961), .B(n36962), .Z(n36607) );
  AND U36658 ( .A(n729), .B(n36963), .Z(n36962) );
  XOR U36659 ( .A(p_input[3256]), .B(p_input[3224]), .Z(n36963) );
  XOR U36660 ( .A(n36964), .B(n36965), .Z(n36955) );
  AND U36661 ( .A(n36966), .B(n36967), .Z(n36965) );
  XOR U36662 ( .A(n36964), .B(n36622), .Z(n36967) );
  XNOR U36663 ( .A(p_input[3287]), .B(n36968), .Z(n36622) );
  AND U36664 ( .A(n731), .B(n36969), .Z(n36968) );
  XOR U36665 ( .A(p_input[3319]), .B(p_input[3287]), .Z(n36969) );
  XNOR U36666 ( .A(n36619), .B(n36964), .Z(n36966) );
  XOR U36667 ( .A(n36970), .B(n36971), .Z(n36619) );
  AND U36668 ( .A(n729), .B(n36972), .Z(n36971) );
  XOR U36669 ( .A(p_input[3255]), .B(p_input[3223]), .Z(n36972) );
  XOR U36670 ( .A(n36973), .B(n36974), .Z(n36964) );
  AND U36671 ( .A(n36975), .B(n36976), .Z(n36974) );
  XOR U36672 ( .A(n36973), .B(n36634), .Z(n36976) );
  XNOR U36673 ( .A(p_input[3286]), .B(n36977), .Z(n36634) );
  AND U36674 ( .A(n731), .B(n36978), .Z(n36977) );
  XOR U36675 ( .A(p_input[3318]), .B(p_input[3286]), .Z(n36978) );
  XNOR U36676 ( .A(n36631), .B(n36973), .Z(n36975) );
  XOR U36677 ( .A(n36979), .B(n36980), .Z(n36631) );
  AND U36678 ( .A(n729), .B(n36981), .Z(n36980) );
  XOR U36679 ( .A(p_input[3254]), .B(p_input[3222]), .Z(n36981) );
  XOR U36680 ( .A(n36982), .B(n36983), .Z(n36973) );
  AND U36681 ( .A(n36984), .B(n36985), .Z(n36983) );
  XOR U36682 ( .A(n36982), .B(n36646), .Z(n36985) );
  XNOR U36683 ( .A(p_input[3285]), .B(n36986), .Z(n36646) );
  AND U36684 ( .A(n731), .B(n36987), .Z(n36986) );
  XOR U36685 ( .A(p_input[3317]), .B(p_input[3285]), .Z(n36987) );
  XNOR U36686 ( .A(n36643), .B(n36982), .Z(n36984) );
  XOR U36687 ( .A(n36988), .B(n36989), .Z(n36643) );
  AND U36688 ( .A(n729), .B(n36990), .Z(n36989) );
  XOR U36689 ( .A(p_input[3253]), .B(p_input[3221]), .Z(n36990) );
  XOR U36690 ( .A(n36991), .B(n36992), .Z(n36982) );
  AND U36691 ( .A(n36993), .B(n36994), .Z(n36992) );
  XOR U36692 ( .A(n36991), .B(n36658), .Z(n36994) );
  XNOR U36693 ( .A(p_input[3284]), .B(n36995), .Z(n36658) );
  AND U36694 ( .A(n731), .B(n36996), .Z(n36995) );
  XOR U36695 ( .A(p_input[3316]), .B(p_input[3284]), .Z(n36996) );
  XNOR U36696 ( .A(n36655), .B(n36991), .Z(n36993) );
  XOR U36697 ( .A(n36997), .B(n36998), .Z(n36655) );
  AND U36698 ( .A(n729), .B(n36999), .Z(n36998) );
  XOR U36699 ( .A(p_input[3252]), .B(p_input[3220]), .Z(n36999) );
  XOR U36700 ( .A(n37000), .B(n37001), .Z(n36991) );
  AND U36701 ( .A(n37002), .B(n37003), .Z(n37001) );
  XOR U36702 ( .A(n37000), .B(n36670), .Z(n37003) );
  XNOR U36703 ( .A(p_input[3283]), .B(n37004), .Z(n36670) );
  AND U36704 ( .A(n731), .B(n37005), .Z(n37004) );
  XOR U36705 ( .A(p_input[3315]), .B(p_input[3283]), .Z(n37005) );
  XNOR U36706 ( .A(n36667), .B(n37000), .Z(n37002) );
  XOR U36707 ( .A(n37006), .B(n37007), .Z(n36667) );
  AND U36708 ( .A(n729), .B(n37008), .Z(n37007) );
  XOR U36709 ( .A(p_input[3251]), .B(p_input[3219]), .Z(n37008) );
  XOR U36710 ( .A(n37009), .B(n37010), .Z(n37000) );
  AND U36711 ( .A(n37011), .B(n37012), .Z(n37010) );
  XOR U36712 ( .A(n37009), .B(n36682), .Z(n37012) );
  XNOR U36713 ( .A(p_input[3282]), .B(n37013), .Z(n36682) );
  AND U36714 ( .A(n731), .B(n37014), .Z(n37013) );
  XOR U36715 ( .A(p_input[3314]), .B(p_input[3282]), .Z(n37014) );
  XNOR U36716 ( .A(n36679), .B(n37009), .Z(n37011) );
  XOR U36717 ( .A(n37015), .B(n37016), .Z(n36679) );
  AND U36718 ( .A(n729), .B(n37017), .Z(n37016) );
  XOR U36719 ( .A(p_input[3250]), .B(p_input[3218]), .Z(n37017) );
  XOR U36720 ( .A(n37018), .B(n37019), .Z(n37009) );
  AND U36721 ( .A(n37020), .B(n37021), .Z(n37019) );
  XOR U36722 ( .A(n37018), .B(n36694), .Z(n37021) );
  XNOR U36723 ( .A(p_input[3281]), .B(n37022), .Z(n36694) );
  AND U36724 ( .A(n731), .B(n37023), .Z(n37022) );
  XOR U36725 ( .A(p_input[3313]), .B(p_input[3281]), .Z(n37023) );
  XNOR U36726 ( .A(n36691), .B(n37018), .Z(n37020) );
  XOR U36727 ( .A(n37024), .B(n37025), .Z(n36691) );
  AND U36728 ( .A(n729), .B(n37026), .Z(n37025) );
  XOR U36729 ( .A(p_input[3249]), .B(p_input[3217]), .Z(n37026) );
  XOR U36730 ( .A(n37027), .B(n37028), .Z(n37018) );
  AND U36731 ( .A(n37029), .B(n37030), .Z(n37028) );
  XOR U36732 ( .A(n37027), .B(n36706), .Z(n37030) );
  XNOR U36733 ( .A(p_input[3280]), .B(n37031), .Z(n36706) );
  AND U36734 ( .A(n731), .B(n37032), .Z(n37031) );
  XOR U36735 ( .A(p_input[3312]), .B(p_input[3280]), .Z(n37032) );
  XNOR U36736 ( .A(n36703), .B(n37027), .Z(n37029) );
  XOR U36737 ( .A(n37033), .B(n37034), .Z(n36703) );
  AND U36738 ( .A(n729), .B(n37035), .Z(n37034) );
  XOR U36739 ( .A(p_input[3248]), .B(p_input[3216]), .Z(n37035) );
  XOR U36740 ( .A(n37036), .B(n37037), .Z(n37027) );
  AND U36741 ( .A(n37038), .B(n37039), .Z(n37037) );
  XOR U36742 ( .A(n37036), .B(n36718), .Z(n37039) );
  XNOR U36743 ( .A(p_input[3279]), .B(n37040), .Z(n36718) );
  AND U36744 ( .A(n731), .B(n37041), .Z(n37040) );
  XOR U36745 ( .A(p_input[3311]), .B(p_input[3279]), .Z(n37041) );
  XNOR U36746 ( .A(n36715), .B(n37036), .Z(n37038) );
  XOR U36747 ( .A(n37042), .B(n37043), .Z(n36715) );
  AND U36748 ( .A(n729), .B(n37044), .Z(n37043) );
  XOR U36749 ( .A(p_input[3247]), .B(p_input[3215]), .Z(n37044) );
  XOR U36750 ( .A(n37045), .B(n37046), .Z(n37036) );
  AND U36751 ( .A(n37047), .B(n37048), .Z(n37046) );
  XOR U36752 ( .A(n37045), .B(n36730), .Z(n37048) );
  XNOR U36753 ( .A(p_input[3278]), .B(n37049), .Z(n36730) );
  AND U36754 ( .A(n731), .B(n37050), .Z(n37049) );
  XOR U36755 ( .A(p_input[3310]), .B(p_input[3278]), .Z(n37050) );
  XNOR U36756 ( .A(n36727), .B(n37045), .Z(n37047) );
  XOR U36757 ( .A(n37051), .B(n37052), .Z(n36727) );
  AND U36758 ( .A(n729), .B(n37053), .Z(n37052) );
  XOR U36759 ( .A(p_input[3246]), .B(p_input[3214]), .Z(n37053) );
  XOR U36760 ( .A(n37054), .B(n37055), .Z(n37045) );
  AND U36761 ( .A(n37056), .B(n37057), .Z(n37055) );
  XOR U36762 ( .A(n37054), .B(n36742), .Z(n37057) );
  XNOR U36763 ( .A(p_input[3277]), .B(n37058), .Z(n36742) );
  AND U36764 ( .A(n731), .B(n37059), .Z(n37058) );
  XOR U36765 ( .A(p_input[3309]), .B(p_input[3277]), .Z(n37059) );
  XNOR U36766 ( .A(n36739), .B(n37054), .Z(n37056) );
  XOR U36767 ( .A(n37060), .B(n37061), .Z(n36739) );
  AND U36768 ( .A(n729), .B(n37062), .Z(n37061) );
  XOR U36769 ( .A(p_input[3245]), .B(p_input[3213]), .Z(n37062) );
  XOR U36770 ( .A(n37063), .B(n37064), .Z(n37054) );
  AND U36771 ( .A(n37065), .B(n37066), .Z(n37064) );
  XOR U36772 ( .A(n37063), .B(n36754), .Z(n37066) );
  XNOR U36773 ( .A(p_input[3276]), .B(n37067), .Z(n36754) );
  AND U36774 ( .A(n731), .B(n37068), .Z(n37067) );
  XOR U36775 ( .A(p_input[3308]), .B(p_input[3276]), .Z(n37068) );
  XNOR U36776 ( .A(n36751), .B(n37063), .Z(n37065) );
  XOR U36777 ( .A(n37069), .B(n37070), .Z(n36751) );
  AND U36778 ( .A(n729), .B(n37071), .Z(n37070) );
  XOR U36779 ( .A(p_input[3244]), .B(p_input[3212]), .Z(n37071) );
  XOR U36780 ( .A(n37072), .B(n37073), .Z(n37063) );
  AND U36781 ( .A(n37074), .B(n37075), .Z(n37073) );
  XOR U36782 ( .A(n37072), .B(n36766), .Z(n37075) );
  XNOR U36783 ( .A(p_input[3275]), .B(n37076), .Z(n36766) );
  AND U36784 ( .A(n731), .B(n37077), .Z(n37076) );
  XOR U36785 ( .A(p_input[3307]), .B(p_input[3275]), .Z(n37077) );
  XNOR U36786 ( .A(n36763), .B(n37072), .Z(n37074) );
  XOR U36787 ( .A(n37078), .B(n37079), .Z(n36763) );
  AND U36788 ( .A(n729), .B(n37080), .Z(n37079) );
  XOR U36789 ( .A(p_input[3243]), .B(p_input[3211]), .Z(n37080) );
  XOR U36790 ( .A(n37081), .B(n37082), .Z(n37072) );
  AND U36791 ( .A(n37083), .B(n37084), .Z(n37082) );
  XOR U36792 ( .A(n37081), .B(n36778), .Z(n37084) );
  XNOR U36793 ( .A(p_input[3274]), .B(n37085), .Z(n36778) );
  AND U36794 ( .A(n731), .B(n37086), .Z(n37085) );
  XOR U36795 ( .A(p_input[3306]), .B(p_input[3274]), .Z(n37086) );
  XNOR U36796 ( .A(n36775), .B(n37081), .Z(n37083) );
  XOR U36797 ( .A(n37087), .B(n37088), .Z(n36775) );
  AND U36798 ( .A(n729), .B(n37089), .Z(n37088) );
  XOR U36799 ( .A(p_input[3242]), .B(p_input[3210]), .Z(n37089) );
  XOR U36800 ( .A(n37090), .B(n37091), .Z(n37081) );
  AND U36801 ( .A(n37092), .B(n37093), .Z(n37091) );
  XOR U36802 ( .A(n37090), .B(n36790), .Z(n37093) );
  XNOR U36803 ( .A(p_input[3273]), .B(n37094), .Z(n36790) );
  AND U36804 ( .A(n731), .B(n37095), .Z(n37094) );
  XOR U36805 ( .A(p_input[3305]), .B(p_input[3273]), .Z(n37095) );
  XNOR U36806 ( .A(n36787), .B(n37090), .Z(n37092) );
  XOR U36807 ( .A(n37096), .B(n37097), .Z(n36787) );
  AND U36808 ( .A(n729), .B(n37098), .Z(n37097) );
  XOR U36809 ( .A(p_input[3241]), .B(p_input[3209]), .Z(n37098) );
  XOR U36810 ( .A(n37099), .B(n37100), .Z(n37090) );
  AND U36811 ( .A(n37101), .B(n37102), .Z(n37100) );
  XOR U36812 ( .A(n37099), .B(n36802), .Z(n37102) );
  XNOR U36813 ( .A(p_input[3272]), .B(n37103), .Z(n36802) );
  AND U36814 ( .A(n731), .B(n37104), .Z(n37103) );
  XOR U36815 ( .A(p_input[3304]), .B(p_input[3272]), .Z(n37104) );
  XNOR U36816 ( .A(n36799), .B(n37099), .Z(n37101) );
  XOR U36817 ( .A(n37105), .B(n37106), .Z(n36799) );
  AND U36818 ( .A(n729), .B(n37107), .Z(n37106) );
  XOR U36819 ( .A(p_input[3240]), .B(p_input[3208]), .Z(n37107) );
  XOR U36820 ( .A(n37108), .B(n37109), .Z(n37099) );
  AND U36821 ( .A(n37110), .B(n37111), .Z(n37109) );
  XOR U36822 ( .A(n37108), .B(n36814), .Z(n37111) );
  XNOR U36823 ( .A(p_input[3271]), .B(n37112), .Z(n36814) );
  AND U36824 ( .A(n731), .B(n37113), .Z(n37112) );
  XOR U36825 ( .A(p_input[3303]), .B(p_input[3271]), .Z(n37113) );
  XNOR U36826 ( .A(n36811), .B(n37108), .Z(n37110) );
  XOR U36827 ( .A(n37114), .B(n37115), .Z(n36811) );
  AND U36828 ( .A(n729), .B(n37116), .Z(n37115) );
  XOR U36829 ( .A(p_input[3239]), .B(p_input[3207]), .Z(n37116) );
  XOR U36830 ( .A(n37117), .B(n37118), .Z(n37108) );
  AND U36831 ( .A(n37119), .B(n37120), .Z(n37118) );
  XOR U36832 ( .A(n37117), .B(n36826), .Z(n37120) );
  XNOR U36833 ( .A(p_input[3270]), .B(n37121), .Z(n36826) );
  AND U36834 ( .A(n731), .B(n37122), .Z(n37121) );
  XOR U36835 ( .A(p_input[3302]), .B(p_input[3270]), .Z(n37122) );
  XNOR U36836 ( .A(n36823), .B(n37117), .Z(n37119) );
  XOR U36837 ( .A(n37123), .B(n37124), .Z(n36823) );
  AND U36838 ( .A(n729), .B(n37125), .Z(n37124) );
  XOR U36839 ( .A(p_input[3238]), .B(p_input[3206]), .Z(n37125) );
  XOR U36840 ( .A(n37126), .B(n37127), .Z(n37117) );
  AND U36841 ( .A(n37128), .B(n37129), .Z(n37127) );
  XOR U36842 ( .A(n37126), .B(n36838), .Z(n37129) );
  XNOR U36843 ( .A(p_input[3269]), .B(n37130), .Z(n36838) );
  AND U36844 ( .A(n731), .B(n37131), .Z(n37130) );
  XOR U36845 ( .A(p_input[3301]), .B(p_input[3269]), .Z(n37131) );
  XNOR U36846 ( .A(n36835), .B(n37126), .Z(n37128) );
  XOR U36847 ( .A(n37132), .B(n37133), .Z(n36835) );
  AND U36848 ( .A(n729), .B(n37134), .Z(n37133) );
  XOR U36849 ( .A(p_input[3237]), .B(p_input[3205]), .Z(n37134) );
  XOR U36850 ( .A(n37135), .B(n37136), .Z(n37126) );
  AND U36851 ( .A(n37137), .B(n37138), .Z(n37136) );
  XOR U36852 ( .A(n37135), .B(n36850), .Z(n37138) );
  XNOR U36853 ( .A(p_input[3268]), .B(n37139), .Z(n36850) );
  AND U36854 ( .A(n731), .B(n37140), .Z(n37139) );
  XOR U36855 ( .A(p_input[3300]), .B(p_input[3268]), .Z(n37140) );
  XNOR U36856 ( .A(n36847), .B(n37135), .Z(n37137) );
  XOR U36857 ( .A(n37141), .B(n37142), .Z(n36847) );
  AND U36858 ( .A(n729), .B(n37143), .Z(n37142) );
  XOR U36859 ( .A(p_input[3236]), .B(p_input[3204]), .Z(n37143) );
  XOR U36860 ( .A(n37144), .B(n37145), .Z(n37135) );
  AND U36861 ( .A(n37146), .B(n37147), .Z(n37145) );
  XOR U36862 ( .A(n37144), .B(n36862), .Z(n37147) );
  XNOR U36863 ( .A(p_input[3267]), .B(n37148), .Z(n36862) );
  AND U36864 ( .A(n731), .B(n37149), .Z(n37148) );
  XOR U36865 ( .A(p_input[3299]), .B(p_input[3267]), .Z(n37149) );
  XNOR U36866 ( .A(n36859), .B(n37144), .Z(n37146) );
  XOR U36867 ( .A(n37150), .B(n37151), .Z(n36859) );
  AND U36868 ( .A(n729), .B(n37152), .Z(n37151) );
  XOR U36869 ( .A(p_input[3235]), .B(p_input[3203]), .Z(n37152) );
  XOR U36870 ( .A(n37153), .B(n37154), .Z(n37144) );
  AND U36871 ( .A(n37155), .B(n37156), .Z(n37154) );
  XOR U36872 ( .A(n37153), .B(n36874), .Z(n37156) );
  XNOR U36873 ( .A(p_input[3266]), .B(n37157), .Z(n36874) );
  AND U36874 ( .A(n731), .B(n37158), .Z(n37157) );
  XOR U36875 ( .A(p_input[3298]), .B(p_input[3266]), .Z(n37158) );
  XNOR U36876 ( .A(n36871), .B(n37153), .Z(n37155) );
  XOR U36877 ( .A(n37159), .B(n37160), .Z(n36871) );
  AND U36878 ( .A(n729), .B(n37161), .Z(n37160) );
  XOR U36879 ( .A(p_input[3234]), .B(p_input[3202]), .Z(n37161) );
  XOR U36880 ( .A(n37162), .B(n37163), .Z(n37153) );
  AND U36881 ( .A(n37164), .B(n37165), .Z(n37163) );
  XNOR U36882 ( .A(n37166), .B(n36887), .Z(n37165) );
  XNOR U36883 ( .A(p_input[3265]), .B(n37167), .Z(n36887) );
  AND U36884 ( .A(n731), .B(n37168), .Z(n37167) );
  XNOR U36885 ( .A(p_input[3297]), .B(n37169), .Z(n37168) );
  IV U36886 ( .A(p_input[3265]), .Z(n37169) );
  XNOR U36887 ( .A(n36884), .B(n37162), .Z(n37164) );
  XNOR U36888 ( .A(p_input[3201]), .B(n37170), .Z(n36884) );
  AND U36889 ( .A(n729), .B(n37171), .Z(n37170) );
  XOR U36890 ( .A(p_input[3233]), .B(p_input[3201]), .Z(n37171) );
  IV U36891 ( .A(n37166), .Z(n37162) );
  AND U36892 ( .A(n36892), .B(n36895), .Z(n37166) );
  XOR U36893 ( .A(p_input[3264]), .B(n37172), .Z(n36895) );
  AND U36894 ( .A(n731), .B(n37173), .Z(n37172) );
  XOR U36895 ( .A(p_input[3296]), .B(p_input[3264]), .Z(n37173) );
  XOR U36896 ( .A(n37174), .B(n37175), .Z(n731) );
  AND U36897 ( .A(n37176), .B(n37177), .Z(n37175) );
  XNOR U36898 ( .A(p_input[3327]), .B(n37174), .Z(n37177) );
  XOR U36899 ( .A(n37174), .B(p_input[3295]), .Z(n37176) );
  XOR U36900 ( .A(n37178), .B(n37179), .Z(n37174) );
  AND U36901 ( .A(n37180), .B(n37181), .Z(n37179) );
  XNOR U36902 ( .A(p_input[3326]), .B(n37178), .Z(n37181) );
  XOR U36903 ( .A(n37178), .B(p_input[3294]), .Z(n37180) );
  XOR U36904 ( .A(n37182), .B(n37183), .Z(n37178) );
  AND U36905 ( .A(n37184), .B(n37185), .Z(n37183) );
  XNOR U36906 ( .A(p_input[3325]), .B(n37182), .Z(n37185) );
  XOR U36907 ( .A(n37182), .B(p_input[3293]), .Z(n37184) );
  XOR U36908 ( .A(n37186), .B(n37187), .Z(n37182) );
  AND U36909 ( .A(n37188), .B(n37189), .Z(n37187) );
  XNOR U36910 ( .A(p_input[3324]), .B(n37186), .Z(n37189) );
  XOR U36911 ( .A(n37186), .B(p_input[3292]), .Z(n37188) );
  XOR U36912 ( .A(n37190), .B(n37191), .Z(n37186) );
  AND U36913 ( .A(n37192), .B(n37193), .Z(n37191) );
  XNOR U36914 ( .A(p_input[3323]), .B(n37190), .Z(n37193) );
  XOR U36915 ( .A(n37190), .B(p_input[3291]), .Z(n37192) );
  XOR U36916 ( .A(n37194), .B(n37195), .Z(n37190) );
  AND U36917 ( .A(n37196), .B(n37197), .Z(n37195) );
  XNOR U36918 ( .A(p_input[3322]), .B(n37194), .Z(n37197) );
  XOR U36919 ( .A(n37194), .B(p_input[3290]), .Z(n37196) );
  XOR U36920 ( .A(n37198), .B(n37199), .Z(n37194) );
  AND U36921 ( .A(n37200), .B(n37201), .Z(n37199) );
  XNOR U36922 ( .A(p_input[3321]), .B(n37198), .Z(n37201) );
  XOR U36923 ( .A(n37198), .B(p_input[3289]), .Z(n37200) );
  XOR U36924 ( .A(n37202), .B(n37203), .Z(n37198) );
  AND U36925 ( .A(n37204), .B(n37205), .Z(n37203) );
  XNOR U36926 ( .A(p_input[3320]), .B(n37202), .Z(n37205) );
  XOR U36927 ( .A(n37202), .B(p_input[3288]), .Z(n37204) );
  XOR U36928 ( .A(n37206), .B(n37207), .Z(n37202) );
  AND U36929 ( .A(n37208), .B(n37209), .Z(n37207) );
  XNOR U36930 ( .A(p_input[3319]), .B(n37206), .Z(n37209) );
  XOR U36931 ( .A(n37206), .B(p_input[3287]), .Z(n37208) );
  XOR U36932 ( .A(n37210), .B(n37211), .Z(n37206) );
  AND U36933 ( .A(n37212), .B(n37213), .Z(n37211) );
  XNOR U36934 ( .A(p_input[3318]), .B(n37210), .Z(n37213) );
  XOR U36935 ( .A(n37210), .B(p_input[3286]), .Z(n37212) );
  XOR U36936 ( .A(n37214), .B(n37215), .Z(n37210) );
  AND U36937 ( .A(n37216), .B(n37217), .Z(n37215) );
  XNOR U36938 ( .A(p_input[3317]), .B(n37214), .Z(n37217) );
  XOR U36939 ( .A(n37214), .B(p_input[3285]), .Z(n37216) );
  XOR U36940 ( .A(n37218), .B(n37219), .Z(n37214) );
  AND U36941 ( .A(n37220), .B(n37221), .Z(n37219) );
  XNOR U36942 ( .A(p_input[3316]), .B(n37218), .Z(n37221) );
  XOR U36943 ( .A(n37218), .B(p_input[3284]), .Z(n37220) );
  XOR U36944 ( .A(n37222), .B(n37223), .Z(n37218) );
  AND U36945 ( .A(n37224), .B(n37225), .Z(n37223) );
  XNOR U36946 ( .A(p_input[3315]), .B(n37222), .Z(n37225) );
  XOR U36947 ( .A(n37222), .B(p_input[3283]), .Z(n37224) );
  XOR U36948 ( .A(n37226), .B(n37227), .Z(n37222) );
  AND U36949 ( .A(n37228), .B(n37229), .Z(n37227) );
  XNOR U36950 ( .A(p_input[3314]), .B(n37226), .Z(n37229) );
  XOR U36951 ( .A(n37226), .B(p_input[3282]), .Z(n37228) );
  XOR U36952 ( .A(n37230), .B(n37231), .Z(n37226) );
  AND U36953 ( .A(n37232), .B(n37233), .Z(n37231) );
  XNOR U36954 ( .A(p_input[3313]), .B(n37230), .Z(n37233) );
  XOR U36955 ( .A(n37230), .B(p_input[3281]), .Z(n37232) );
  XOR U36956 ( .A(n37234), .B(n37235), .Z(n37230) );
  AND U36957 ( .A(n37236), .B(n37237), .Z(n37235) );
  XNOR U36958 ( .A(p_input[3312]), .B(n37234), .Z(n37237) );
  XOR U36959 ( .A(n37234), .B(p_input[3280]), .Z(n37236) );
  XOR U36960 ( .A(n37238), .B(n37239), .Z(n37234) );
  AND U36961 ( .A(n37240), .B(n37241), .Z(n37239) );
  XNOR U36962 ( .A(p_input[3311]), .B(n37238), .Z(n37241) );
  XOR U36963 ( .A(n37238), .B(p_input[3279]), .Z(n37240) );
  XOR U36964 ( .A(n37242), .B(n37243), .Z(n37238) );
  AND U36965 ( .A(n37244), .B(n37245), .Z(n37243) );
  XNOR U36966 ( .A(p_input[3310]), .B(n37242), .Z(n37245) );
  XOR U36967 ( .A(n37242), .B(p_input[3278]), .Z(n37244) );
  XOR U36968 ( .A(n37246), .B(n37247), .Z(n37242) );
  AND U36969 ( .A(n37248), .B(n37249), .Z(n37247) );
  XNOR U36970 ( .A(p_input[3309]), .B(n37246), .Z(n37249) );
  XOR U36971 ( .A(n37246), .B(p_input[3277]), .Z(n37248) );
  XOR U36972 ( .A(n37250), .B(n37251), .Z(n37246) );
  AND U36973 ( .A(n37252), .B(n37253), .Z(n37251) );
  XNOR U36974 ( .A(p_input[3308]), .B(n37250), .Z(n37253) );
  XOR U36975 ( .A(n37250), .B(p_input[3276]), .Z(n37252) );
  XOR U36976 ( .A(n37254), .B(n37255), .Z(n37250) );
  AND U36977 ( .A(n37256), .B(n37257), .Z(n37255) );
  XNOR U36978 ( .A(p_input[3307]), .B(n37254), .Z(n37257) );
  XOR U36979 ( .A(n37254), .B(p_input[3275]), .Z(n37256) );
  XOR U36980 ( .A(n37258), .B(n37259), .Z(n37254) );
  AND U36981 ( .A(n37260), .B(n37261), .Z(n37259) );
  XNOR U36982 ( .A(p_input[3306]), .B(n37258), .Z(n37261) );
  XOR U36983 ( .A(n37258), .B(p_input[3274]), .Z(n37260) );
  XOR U36984 ( .A(n37262), .B(n37263), .Z(n37258) );
  AND U36985 ( .A(n37264), .B(n37265), .Z(n37263) );
  XNOR U36986 ( .A(p_input[3305]), .B(n37262), .Z(n37265) );
  XOR U36987 ( .A(n37262), .B(p_input[3273]), .Z(n37264) );
  XOR U36988 ( .A(n37266), .B(n37267), .Z(n37262) );
  AND U36989 ( .A(n37268), .B(n37269), .Z(n37267) );
  XNOR U36990 ( .A(p_input[3304]), .B(n37266), .Z(n37269) );
  XOR U36991 ( .A(n37266), .B(p_input[3272]), .Z(n37268) );
  XOR U36992 ( .A(n37270), .B(n37271), .Z(n37266) );
  AND U36993 ( .A(n37272), .B(n37273), .Z(n37271) );
  XNOR U36994 ( .A(p_input[3303]), .B(n37270), .Z(n37273) );
  XOR U36995 ( .A(n37270), .B(p_input[3271]), .Z(n37272) );
  XOR U36996 ( .A(n37274), .B(n37275), .Z(n37270) );
  AND U36997 ( .A(n37276), .B(n37277), .Z(n37275) );
  XNOR U36998 ( .A(p_input[3302]), .B(n37274), .Z(n37277) );
  XOR U36999 ( .A(n37274), .B(p_input[3270]), .Z(n37276) );
  XOR U37000 ( .A(n37278), .B(n37279), .Z(n37274) );
  AND U37001 ( .A(n37280), .B(n37281), .Z(n37279) );
  XNOR U37002 ( .A(p_input[3301]), .B(n37278), .Z(n37281) );
  XOR U37003 ( .A(n37278), .B(p_input[3269]), .Z(n37280) );
  XOR U37004 ( .A(n37282), .B(n37283), .Z(n37278) );
  AND U37005 ( .A(n37284), .B(n37285), .Z(n37283) );
  XNOR U37006 ( .A(p_input[3300]), .B(n37282), .Z(n37285) );
  XOR U37007 ( .A(n37282), .B(p_input[3268]), .Z(n37284) );
  XOR U37008 ( .A(n37286), .B(n37287), .Z(n37282) );
  AND U37009 ( .A(n37288), .B(n37289), .Z(n37287) );
  XNOR U37010 ( .A(p_input[3299]), .B(n37286), .Z(n37289) );
  XOR U37011 ( .A(n37286), .B(p_input[3267]), .Z(n37288) );
  XOR U37012 ( .A(n37290), .B(n37291), .Z(n37286) );
  AND U37013 ( .A(n37292), .B(n37293), .Z(n37291) );
  XNOR U37014 ( .A(p_input[3298]), .B(n37290), .Z(n37293) );
  XOR U37015 ( .A(n37290), .B(p_input[3266]), .Z(n37292) );
  XNOR U37016 ( .A(n37294), .B(n37295), .Z(n37290) );
  AND U37017 ( .A(n37296), .B(n37297), .Z(n37295) );
  XOR U37018 ( .A(p_input[3297]), .B(n37294), .Z(n37297) );
  XNOR U37019 ( .A(p_input[3265]), .B(n37294), .Z(n37296) );
  AND U37020 ( .A(p_input[3296]), .B(n37298), .Z(n37294) );
  IV U37021 ( .A(p_input[3264]), .Z(n37298) );
  XNOR U37022 ( .A(p_input[3200]), .B(n37299), .Z(n36892) );
  AND U37023 ( .A(n729), .B(n37300), .Z(n37299) );
  XOR U37024 ( .A(p_input[3232]), .B(p_input[3200]), .Z(n37300) );
  XOR U37025 ( .A(n37301), .B(n37302), .Z(n729) );
  AND U37026 ( .A(n37303), .B(n37304), .Z(n37302) );
  XNOR U37027 ( .A(p_input[3263]), .B(n37301), .Z(n37304) );
  XOR U37028 ( .A(n37301), .B(p_input[3231]), .Z(n37303) );
  XOR U37029 ( .A(n37305), .B(n37306), .Z(n37301) );
  AND U37030 ( .A(n37307), .B(n37308), .Z(n37306) );
  XNOR U37031 ( .A(p_input[3262]), .B(n37305), .Z(n37308) );
  XNOR U37032 ( .A(n37305), .B(n36907), .Z(n37307) );
  IV U37033 ( .A(p_input[3230]), .Z(n36907) );
  XOR U37034 ( .A(n37309), .B(n37310), .Z(n37305) );
  AND U37035 ( .A(n37311), .B(n37312), .Z(n37310) );
  XNOR U37036 ( .A(p_input[3261]), .B(n37309), .Z(n37312) );
  XNOR U37037 ( .A(n37309), .B(n36916), .Z(n37311) );
  IV U37038 ( .A(p_input[3229]), .Z(n36916) );
  XOR U37039 ( .A(n37313), .B(n37314), .Z(n37309) );
  AND U37040 ( .A(n37315), .B(n37316), .Z(n37314) );
  XNOR U37041 ( .A(p_input[3260]), .B(n37313), .Z(n37316) );
  XNOR U37042 ( .A(n37313), .B(n36925), .Z(n37315) );
  IV U37043 ( .A(p_input[3228]), .Z(n36925) );
  XOR U37044 ( .A(n37317), .B(n37318), .Z(n37313) );
  AND U37045 ( .A(n37319), .B(n37320), .Z(n37318) );
  XNOR U37046 ( .A(p_input[3259]), .B(n37317), .Z(n37320) );
  XNOR U37047 ( .A(n37317), .B(n36934), .Z(n37319) );
  IV U37048 ( .A(p_input[3227]), .Z(n36934) );
  XOR U37049 ( .A(n37321), .B(n37322), .Z(n37317) );
  AND U37050 ( .A(n37323), .B(n37324), .Z(n37322) );
  XNOR U37051 ( .A(p_input[3258]), .B(n37321), .Z(n37324) );
  XNOR U37052 ( .A(n37321), .B(n36943), .Z(n37323) );
  IV U37053 ( .A(p_input[3226]), .Z(n36943) );
  XOR U37054 ( .A(n37325), .B(n37326), .Z(n37321) );
  AND U37055 ( .A(n37327), .B(n37328), .Z(n37326) );
  XNOR U37056 ( .A(p_input[3257]), .B(n37325), .Z(n37328) );
  XNOR U37057 ( .A(n37325), .B(n36952), .Z(n37327) );
  IV U37058 ( .A(p_input[3225]), .Z(n36952) );
  XOR U37059 ( .A(n37329), .B(n37330), .Z(n37325) );
  AND U37060 ( .A(n37331), .B(n37332), .Z(n37330) );
  XNOR U37061 ( .A(p_input[3256]), .B(n37329), .Z(n37332) );
  XNOR U37062 ( .A(n37329), .B(n36961), .Z(n37331) );
  IV U37063 ( .A(p_input[3224]), .Z(n36961) );
  XOR U37064 ( .A(n37333), .B(n37334), .Z(n37329) );
  AND U37065 ( .A(n37335), .B(n37336), .Z(n37334) );
  XNOR U37066 ( .A(p_input[3255]), .B(n37333), .Z(n37336) );
  XNOR U37067 ( .A(n37333), .B(n36970), .Z(n37335) );
  IV U37068 ( .A(p_input[3223]), .Z(n36970) );
  XOR U37069 ( .A(n37337), .B(n37338), .Z(n37333) );
  AND U37070 ( .A(n37339), .B(n37340), .Z(n37338) );
  XNOR U37071 ( .A(p_input[3254]), .B(n37337), .Z(n37340) );
  XNOR U37072 ( .A(n37337), .B(n36979), .Z(n37339) );
  IV U37073 ( .A(p_input[3222]), .Z(n36979) );
  XOR U37074 ( .A(n37341), .B(n37342), .Z(n37337) );
  AND U37075 ( .A(n37343), .B(n37344), .Z(n37342) );
  XNOR U37076 ( .A(p_input[3253]), .B(n37341), .Z(n37344) );
  XNOR U37077 ( .A(n37341), .B(n36988), .Z(n37343) );
  IV U37078 ( .A(p_input[3221]), .Z(n36988) );
  XOR U37079 ( .A(n37345), .B(n37346), .Z(n37341) );
  AND U37080 ( .A(n37347), .B(n37348), .Z(n37346) );
  XNOR U37081 ( .A(p_input[3252]), .B(n37345), .Z(n37348) );
  XNOR U37082 ( .A(n37345), .B(n36997), .Z(n37347) );
  IV U37083 ( .A(p_input[3220]), .Z(n36997) );
  XOR U37084 ( .A(n37349), .B(n37350), .Z(n37345) );
  AND U37085 ( .A(n37351), .B(n37352), .Z(n37350) );
  XNOR U37086 ( .A(p_input[3251]), .B(n37349), .Z(n37352) );
  XNOR U37087 ( .A(n37349), .B(n37006), .Z(n37351) );
  IV U37088 ( .A(p_input[3219]), .Z(n37006) );
  XOR U37089 ( .A(n37353), .B(n37354), .Z(n37349) );
  AND U37090 ( .A(n37355), .B(n37356), .Z(n37354) );
  XNOR U37091 ( .A(p_input[3250]), .B(n37353), .Z(n37356) );
  XNOR U37092 ( .A(n37353), .B(n37015), .Z(n37355) );
  IV U37093 ( .A(p_input[3218]), .Z(n37015) );
  XOR U37094 ( .A(n37357), .B(n37358), .Z(n37353) );
  AND U37095 ( .A(n37359), .B(n37360), .Z(n37358) );
  XNOR U37096 ( .A(p_input[3249]), .B(n37357), .Z(n37360) );
  XNOR U37097 ( .A(n37357), .B(n37024), .Z(n37359) );
  IV U37098 ( .A(p_input[3217]), .Z(n37024) );
  XOR U37099 ( .A(n37361), .B(n37362), .Z(n37357) );
  AND U37100 ( .A(n37363), .B(n37364), .Z(n37362) );
  XNOR U37101 ( .A(p_input[3248]), .B(n37361), .Z(n37364) );
  XNOR U37102 ( .A(n37361), .B(n37033), .Z(n37363) );
  IV U37103 ( .A(p_input[3216]), .Z(n37033) );
  XOR U37104 ( .A(n37365), .B(n37366), .Z(n37361) );
  AND U37105 ( .A(n37367), .B(n37368), .Z(n37366) );
  XNOR U37106 ( .A(p_input[3247]), .B(n37365), .Z(n37368) );
  XNOR U37107 ( .A(n37365), .B(n37042), .Z(n37367) );
  IV U37108 ( .A(p_input[3215]), .Z(n37042) );
  XOR U37109 ( .A(n37369), .B(n37370), .Z(n37365) );
  AND U37110 ( .A(n37371), .B(n37372), .Z(n37370) );
  XNOR U37111 ( .A(p_input[3246]), .B(n37369), .Z(n37372) );
  XNOR U37112 ( .A(n37369), .B(n37051), .Z(n37371) );
  IV U37113 ( .A(p_input[3214]), .Z(n37051) );
  XOR U37114 ( .A(n37373), .B(n37374), .Z(n37369) );
  AND U37115 ( .A(n37375), .B(n37376), .Z(n37374) );
  XNOR U37116 ( .A(p_input[3245]), .B(n37373), .Z(n37376) );
  XNOR U37117 ( .A(n37373), .B(n37060), .Z(n37375) );
  IV U37118 ( .A(p_input[3213]), .Z(n37060) );
  XOR U37119 ( .A(n37377), .B(n37378), .Z(n37373) );
  AND U37120 ( .A(n37379), .B(n37380), .Z(n37378) );
  XNOR U37121 ( .A(p_input[3244]), .B(n37377), .Z(n37380) );
  XNOR U37122 ( .A(n37377), .B(n37069), .Z(n37379) );
  IV U37123 ( .A(p_input[3212]), .Z(n37069) );
  XOR U37124 ( .A(n37381), .B(n37382), .Z(n37377) );
  AND U37125 ( .A(n37383), .B(n37384), .Z(n37382) );
  XNOR U37126 ( .A(p_input[3243]), .B(n37381), .Z(n37384) );
  XNOR U37127 ( .A(n37381), .B(n37078), .Z(n37383) );
  IV U37128 ( .A(p_input[3211]), .Z(n37078) );
  XOR U37129 ( .A(n37385), .B(n37386), .Z(n37381) );
  AND U37130 ( .A(n37387), .B(n37388), .Z(n37386) );
  XNOR U37131 ( .A(p_input[3242]), .B(n37385), .Z(n37388) );
  XNOR U37132 ( .A(n37385), .B(n37087), .Z(n37387) );
  IV U37133 ( .A(p_input[3210]), .Z(n37087) );
  XOR U37134 ( .A(n37389), .B(n37390), .Z(n37385) );
  AND U37135 ( .A(n37391), .B(n37392), .Z(n37390) );
  XNOR U37136 ( .A(p_input[3241]), .B(n37389), .Z(n37392) );
  XNOR U37137 ( .A(n37389), .B(n37096), .Z(n37391) );
  IV U37138 ( .A(p_input[3209]), .Z(n37096) );
  XOR U37139 ( .A(n37393), .B(n37394), .Z(n37389) );
  AND U37140 ( .A(n37395), .B(n37396), .Z(n37394) );
  XNOR U37141 ( .A(p_input[3240]), .B(n37393), .Z(n37396) );
  XNOR U37142 ( .A(n37393), .B(n37105), .Z(n37395) );
  IV U37143 ( .A(p_input[3208]), .Z(n37105) );
  XOR U37144 ( .A(n37397), .B(n37398), .Z(n37393) );
  AND U37145 ( .A(n37399), .B(n37400), .Z(n37398) );
  XNOR U37146 ( .A(p_input[3239]), .B(n37397), .Z(n37400) );
  XNOR U37147 ( .A(n37397), .B(n37114), .Z(n37399) );
  IV U37148 ( .A(p_input[3207]), .Z(n37114) );
  XOR U37149 ( .A(n37401), .B(n37402), .Z(n37397) );
  AND U37150 ( .A(n37403), .B(n37404), .Z(n37402) );
  XNOR U37151 ( .A(p_input[3238]), .B(n37401), .Z(n37404) );
  XNOR U37152 ( .A(n37401), .B(n37123), .Z(n37403) );
  IV U37153 ( .A(p_input[3206]), .Z(n37123) );
  XOR U37154 ( .A(n37405), .B(n37406), .Z(n37401) );
  AND U37155 ( .A(n37407), .B(n37408), .Z(n37406) );
  XNOR U37156 ( .A(p_input[3237]), .B(n37405), .Z(n37408) );
  XNOR U37157 ( .A(n37405), .B(n37132), .Z(n37407) );
  IV U37158 ( .A(p_input[3205]), .Z(n37132) );
  XOR U37159 ( .A(n37409), .B(n37410), .Z(n37405) );
  AND U37160 ( .A(n37411), .B(n37412), .Z(n37410) );
  XNOR U37161 ( .A(p_input[3236]), .B(n37409), .Z(n37412) );
  XNOR U37162 ( .A(n37409), .B(n37141), .Z(n37411) );
  IV U37163 ( .A(p_input[3204]), .Z(n37141) );
  XOR U37164 ( .A(n37413), .B(n37414), .Z(n37409) );
  AND U37165 ( .A(n37415), .B(n37416), .Z(n37414) );
  XNOR U37166 ( .A(p_input[3235]), .B(n37413), .Z(n37416) );
  XNOR U37167 ( .A(n37413), .B(n37150), .Z(n37415) );
  IV U37168 ( .A(p_input[3203]), .Z(n37150) );
  XOR U37169 ( .A(n37417), .B(n37418), .Z(n37413) );
  AND U37170 ( .A(n37419), .B(n37420), .Z(n37418) );
  XNOR U37171 ( .A(p_input[3234]), .B(n37417), .Z(n37420) );
  XNOR U37172 ( .A(n37417), .B(n37159), .Z(n37419) );
  IV U37173 ( .A(p_input[3202]), .Z(n37159) );
  XNOR U37174 ( .A(n37421), .B(n37422), .Z(n37417) );
  AND U37175 ( .A(n37423), .B(n37424), .Z(n37422) );
  XOR U37176 ( .A(p_input[3233]), .B(n37421), .Z(n37424) );
  XNOR U37177 ( .A(p_input[3201]), .B(n37421), .Z(n37423) );
  AND U37178 ( .A(p_input[3232]), .B(n37425), .Z(n37421) );
  IV U37179 ( .A(p_input[3200]), .Z(n37425) );
  XOR U37180 ( .A(n37426), .B(n37427), .Z(n36515) );
  AND U37181 ( .A(n576), .B(n37428), .Z(n37427) );
  XNOR U37182 ( .A(n37429), .B(n37426), .Z(n37428) );
  XOR U37183 ( .A(n37430), .B(n37431), .Z(n576) );
  AND U37184 ( .A(n37432), .B(n37433), .Z(n37431) );
  XNOR U37185 ( .A(n36530), .B(n37430), .Z(n37433) );
  AND U37186 ( .A(p_input[3199]), .B(p_input[3167]), .Z(n36530) );
  XNOR U37187 ( .A(n37430), .B(n36527), .Z(n37432) );
  IV U37188 ( .A(n37434), .Z(n36527) );
  AND U37189 ( .A(p_input[3103]), .B(p_input[3135]), .Z(n37434) );
  XOR U37190 ( .A(n37435), .B(n37436), .Z(n37430) );
  AND U37191 ( .A(n37437), .B(n37438), .Z(n37436) );
  XOR U37192 ( .A(n37435), .B(n36542), .Z(n37438) );
  XNOR U37193 ( .A(p_input[3166]), .B(n37439), .Z(n36542) );
  AND U37194 ( .A(n735), .B(n37440), .Z(n37439) );
  XOR U37195 ( .A(p_input[3198]), .B(p_input[3166]), .Z(n37440) );
  XNOR U37196 ( .A(n36539), .B(n37435), .Z(n37437) );
  XOR U37197 ( .A(n37441), .B(n37442), .Z(n36539) );
  AND U37198 ( .A(n732), .B(n37443), .Z(n37442) );
  XOR U37199 ( .A(p_input[3134]), .B(p_input[3102]), .Z(n37443) );
  XOR U37200 ( .A(n37444), .B(n37445), .Z(n37435) );
  AND U37201 ( .A(n37446), .B(n37447), .Z(n37445) );
  XOR U37202 ( .A(n37444), .B(n36554), .Z(n37447) );
  XNOR U37203 ( .A(p_input[3165]), .B(n37448), .Z(n36554) );
  AND U37204 ( .A(n735), .B(n37449), .Z(n37448) );
  XOR U37205 ( .A(p_input[3197]), .B(p_input[3165]), .Z(n37449) );
  XNOR U37206 ( .A(n36551), .B(n37444), .Z(n37446) );
  XOR U37207 ( .A(n37450), .B(n37451), .Z(n36551) );
  AND U37208 ( .A(n732), .B(n37452), .Z(n37451) );
  XOR U37209 ( .A(p_input[3133]), .B(p_input[3101]), .Z(n37452) );
  XOR U37210 ( .A(n37453), .B(n37454), .Z(n37444) );
  AND U37211 ( .A(n37455), .B(n37456), .Z(n37454) );
  XOR U37212 ( .A(n37453), .B(n36566), .Z(n37456) );
  XNOR U37213 ( .A(p_input[3164]), .B(n37457), .Z(n36566) );
  AND U37214 ( .A(n735), .B(n37458), .Z(n37457) );
  XOR U37215 ( .A(p_input[3196]), .B(p_input[3164]), .Z(n37458) );
  XNOR U37216 ( .A(n36563), .B(n37453), .Z(n37455) );
  XOR U37217 ( .A(n37459), .B(n37460), .Z(n36563) );
  AND U37218 ( .A(n732), .B(n37461), .Z(n37460) );
  XOR U37219 ( .A(p_input[3132]), .B(p_input[3100]), .Z(n37461) );
  XOR U37220 ( .A(n37462), .B(n37463), .Z(n37453) );
  AND U37221 ( .A(n37464), .B(n37465), .Z(n37463) );
  XOR U37222 ( .A(n37462), .B(n36578), .Z(n37465) );
  XNOR U37223 ( .A(p_input[3163]), .B(n37466), .Z(n36578) );
  AND U37224 ( .A(n735), .B(n37467), .Z(n37466) );
  XOR U37225 ( .A(p_input[3195]), .B(p_input[3163]), .Z(n37467) );
  XNOR U37226 ( .A(n36575), .B(n37462), .Z(n37464) );
  XOR U37227 ( .A(n37468), .B(n37469), .Z(n36575) );
  AND U37228 ( .A(n732), .B(n37470), .Z(n37469) );
  XOR U37229 ( .A(p_input[3131]), .B(p_input[3099]), .Z(n37470) );
  XOR U37230 ( .A(n37471), .B(n37472), .Z(n37462) );
  AND U37231 ( .A(n37473), .B(n37474), .Z(n37472) );
  XOR U37232 ( .A(n37471), .B(n36590), .Z(n37474) );
  XNOR U37233 ( .A(p_input[3162]), .B(n37475), .Z(n36590) );
  AND U37234 ( .A(n735), .B(n37476), .Z(n37475) );
  XOR U37235 ( .A(p_input[3194]), .B(p_input[3162]), .Z(n37476) );
  XNOR U37236 ( .A(n36587), .B(n37471), .Z(n37473) );
  XOR U37237 ( .A(n37477), .B(n37478), .Z(n36587) );
  AND U37238 ( .A(n732), .B(n37479), .Z(n37478) );
  XOR U37239 ( .A(p_input[3130]), .B(p_input[3098]), .Z(n37479) );
  XOR U37240 ( .A(n37480), .B(n37481), .Z(n37471) );
  AND U37241 ( .A(n37482), .B(n37483), .Z(n37481) );
  XOR U37242 ( .A(n37480), .B(n36602), .Z(n37483) );
  XNOR U37243 ( .A(p_input[3161]), .B(n37484), .Z(n36602) );
  AND U37244 ( .A(n735), .B(n37485), .Z(n37484) );
  XOR U37245 ( .A(p_input[3193]), .B(p_input[3161]), .Z(n37485) );
  XNOR U37246 ( .A(n36599), .B(n37480), .Z(n37482) );
  XOR U37247 ( .A(n37486), .B(n37487), .Z(n36599) );
  AND U37248 ( .A(n732), .B(n37488), .Z(n37487) );
  XOR U37249 ( .A(p_input[3129]), .B(p_input[3097]), .Z(n37488) );
  XOR U37250 ( .A(n37489), .B(n37490), .Z(n37480) );
  AND U37251 ( .A(n37491), .B(n37492), .Z(n37490) );
  XOR U37252 ( .A(n37489), .B(n36614), .Z(n37492) );
  XNOR U37253 ( .A(p_input[3160]), .B(n37493), .Z(n36614) );
  AND U37254 ( .A(n735), .B(n37494), .Z(n37493) );
  XOR U37255 ( .A(p_input[3192]), .B(p_input[3160]), .Z(n37494) );
  XNOR U37256 ( .A(n36611), .B(n37489), .Z(n37491) );
  XOR U37257 ( .A(n37495), .B(n37496), .Z(n36611) );
  AND U37258 ( .A(n732), .B(n37497), .Z(n37496) );
  XOR U37259 ( .A(p_input[3128]), .B(p_input[3096]), .Z(n37497) );
  XOR U37260 ( .A(n37498), .B(n37499), .Z(n37489) );
  AND U37261 ( .A(n37500), .B(n37501), .Z(n37499) );
  XOR U37262 ( .A(n37498), .B(n36626), .Z(n37501) );
  XNOR U37263 ( .A(p_input[3159]), .B(n37502), .Z(n36626) );
  AND U37264 ( .A(n735), .B(n37503), .Z(n37502) );
  XOR U37265 ( .A(p_input[3191]), .B(p_input[3159]), .Z(n37503) );
  XNOR U37266 ( .A(n36623), .B(n37498), .Z(n37500) );
  XOR U37267 ( .A(n37504), .B(n37505), .Z(n36623) );
  AND U37268 ( .A(n732), .B(n37506), .Z(n37505) );
  XOR U37269 ( .A(p_input[3127]), .B(p_input[3095]), .Z(n37506) );
  XOR U37270 ( .A(n37507), .B(n37508), .Z(n37498) );
  AND U37271 ( .A(n37509), .B(n37510), .Z(n37508) );
  XOR U37272 ( .A(n37507), .B(n36638), .Z(n37510) );
  XNOR U37273 ( .A(p_input[3158]), .B(n37511), .Z(n36638) );
  AND U37274 ( .A(n735), .B(n37512), .Z(n37511) );
  XOR U37275 ( .A(p_input[3190]), .B(p_input[3158]), .Z(n37512) );
  XNOR U37276 ( .A(n36635), .B(n37507), .Z(n37509) );
  XOR U37277 ( .A(n37513), .B(n37514), .Z(n36635) );
  AND U37278 ( .A(n732), .B(n37515), .Z(n37514) );
  XOR U37279 ( .A(p_input[3126]), .B(p_input[3094]), .Z(n37515) );
  XOR U37280 ( .A(n37516), .B(n37517), .Z(n37507) );
  AND U37281 ( .A(n37518), .B(n37519), .Z(n37517) );
  XOR U37282 ( .A(n37516), .B(n36650), .Z(n37519) );
  XNOR U37283 ( .A(p_input[3157]), .B(n37520), .Z(n36650) );
  AND U37284 ( .A(n735), .B(n37521), .Z(n37520) );
  XOR U37285 ( .A(p_input[3189]), .B(p_input[3157]), .Z(n37521) );
  XNOR U37286 ( .A(n36647), .B(n37516), .Z(n37518) );
  XOR U37287 ( .A(n37522), .B(n37523), .Z(n36647) );
  AND U37288 ( .A(n732), .B(n37524), .Z(n37523) );
  XOR U37289 ( .A(p_input[3125]), .B(p_input[3093]), .Z(n37524) );
  XOR U37290 ( .A(n37525), .B(n37526), .Z(n37516) );
  AND U37291 ( .A(n37527), .B(n37528), .Z(n37526) );
  XOR U37292 ( .A(n37525), .B(n36662), .Z(n37528) );
  XNOR U37293 ( .A(p_input[3156]), .B(n37529), .Z(n36662) );
  AND U37294 ( .A(n735), .B(n37530), .Z(n37529) );
  XOR U37295 ( .A(p_input[3188]), .B(p_input[3156]), .Z(n37530) );
  XNOR U37296 ( .A(n36659), .B(n37525), .Z(n37527) );
  XOR U37297 ( .A(n37531), .B(n37532), .Z(n36659) );
  AND U37298 ( .A(n732), .B(n37533), .Z(n37532) );
  XOR U37299 ( .A(p_input[3124]), .B(p_input[3092]), .Z(n37533) );
  XOR U37300 ( .A(n37534), .B(n37535), .Z(n37525) );
  AND U37301 ( .A(n37536), .B(n37537), .Z(n37535) );
  XOR U37302 ( .A(n37534), .B(n36674), .Z(n37537) );
  XNOR U37303 ( .A(p_input[3155]), .B(n37538), .Z(n36674) );
  AND U37304 ( .A(n735), .B(n37539), .Z(n37538) );
  XOR U37305 ( .A(p_input[3187]), .B(p_input[3155]), .Z(n37539) );
  XNOR U37306 ( .A(n36671), .B(n37534), .Z(n37536) );
  XOR U37307 ( .A(n37540), .B(n37541), .Z(n36671) );
  AND U37308 ( .A(n732), .B(n37542), .Z(n37541) );
  XOR U37309 ( .A(p_input[3123]), .B(p_input[3091]), .Z(n37542) );
  XOR U37310 ( .A(n37543), .B(n37544), .Z(n37534) );
  AND U37311 ( .A(n37545), .B(n37546), .Z(n37544) );
  XOR U37312 ( .A(n37543), .B(n36686), .Z(n37546) );
  XNOR U37313 ( .A(p_input[3154]), .B(n37547), .Z(n36686) );
  AND U37314 ( .A(n735), .B(n37548), .Z(n37547) );
  XOR U37315 ( .A(p_input[3186]), .B(p_input[3154]), .Z(n37548) );
  XNOR U37316 ( .A(n36683), .B(n37543), .Z(n37545) );
  XOR U37317 ( .A(n37549), .B(n37550), .Z(n36683) );
  AND U37318 ( .A(n732), .B(n37551), .Z(n37550) );
  XOR U37319 ( .A(p_input[3122]), .B(p_input[3090]), .Z(n37551) );
  XOR U37320 ( .A(n37552), .B(n37553), .Z(n37543) );
  AND U37321 ( .A(n37554), .B(n37555), .Z(n37553) );
  XOR U37322 ( .A(n37552), .B(n36698), .Z(n37555) );
  XNOR U37323 ( .A(p_input[3153]), .B(n37556), .Z(n36698) );
  AND U37324 ( .A(n735), .B(n37557), .Z(n37556) );
  XOR U37325 ( .A(p_input[3185]), .B(p_input[3153]), .Z(n37557) );
  XNOR U37326 ( .A(n36695), .B(n37552), .Z(n37554) );
  XOR U37327 ( .A(n37558), .B(n37559), .Z(n36695) );
  AND U37328 ( .A(n732), .B(n37560), .Z(n37559) );
  XOR U37329 ( .A(p_input[3121]), .B(p_input[3089]), .Z(n37560) );
  XOR U37330 ( .A(n37561), .B(n37562), .Z(n37552) );
  AND U37331 ( .A(n37563), .B(n37564), .Z(n37562) );
  XOR U37332 ( .A(n37561), .B(n36710), .Z(n37564) );
  XNOR U37333 ( .A(p_input[3152]), .B(n37565), .Z(n36710) );
  AND U37334 ( .A(n735), .B(n37566), .Z(n37565) );
  XOR U37335 ( .A(p_input[3184]), .B(p_input[3152]), .Z(n37566) );
  XNOR U37336 ( .A(n36707), .B(n37561), .Z(n37563) );
  XOR U37337 ( .A(n37567), .B(n37568), .Z(n36707) );
  AND U37338 ( .A(n732), .B(n37569), .Z(n37568) );
  XOR U37339 ( .A(p_input[3120]), .B(p_input[3088]), .Z(n37569) );
  XOR U37340 ( .A(n37570), .B(n37571), .Z(n37561) );
  AND U37341 ( .A(n37572), .B(n37573), .Z(n37571) );
  XOR U37342 ( .A(n37570), .B(n36722), .Z(n37573) );
  XNOR U37343 ( .A(p_input[3151]), .B(n37574), .Z(n36722) );
  AND U37344 ( .A(n735), .B(n37575), .Z(n37574) );
  XOR U37345 ( .A(p_input[3183]), .B(p_input[3151]), .Z(n37575) );
  XNOR U37346 ( .A(n36719), .B(n37570), .Z(n37572) );
  XOR U37347 ( .A(n37576), .B(n37577), .Z(n36719) );
  AND U37348 ( .A(n732), .B(n37578), .Z(n37577) );
  XOR U37349 ( .A(p_input[3119]), .B(p_input[3087]), .Z(n37578) );
  XOR U37350 ( .A(n37579), .B(n37580), .Z(n37570) );
  AND U37351 ( .A(n37581), .B(n37582), .Z(n37580) );
  XOR U37352 ( .A(n37579), .B(n36734), .Z(n37582) );
  XNOR U37353 ( .A(p_input[3150]), .B(n37583), .Z(n36734) );
  AND U37354 ( .A(n735), .B(n37584), .Z(n37583) );
  XOR U37355 ( .A(p_input[3182]), .B(p_input[3150]), .Z(n37584) );
  XNOR U37356 ( .A(n36731), .B(n37579), .Z(n37581) );
  XOR U37357 ( .A(n37585), .B(n37586), .Z(n36731) );
  AND U37358 ( .A(n732), .B(n37587), .Z(n37586) );
  XOR U37359 ( .A(p_input[3118]), .B(p_input[3086]), .Z(n37587) );
  XOR U37360 ( .A(n37588), .B(n37589), .Z(n37579) );
  AND U37361 ( .A(n37590), .B(n37591), .Z(n37589) );
  XOR U37362 ( .A(n37588), .B(n36746), .Z(n37591) );
  XNOR U37363 ( .A(p_input[3149]), .B(n37592), .Z(n36746) );
  AND U37364 ( .A(n735), .B(n37593), .Z(n37592) );
  XOR U37365 ( .A(p_input[3181]), .B(p_input[3149]), .Z(n37593) );
  XNOR U37366 ( .A(n36743), .B(n37588), .Z(n37590) );
  XOR U37367 ( .A(n37594), .B(n37595), .Z(n36743) );
  AND U37368 ( .A(n732), .B(n37596), .Z(n37595) );
  XOR U37369 ( .A(p_input[3117]), .B(p_input[3085]), .Z(n37596) );
  XOR U37370 ( .A(n37597), .B(n37598), .Z(n37588) );
  AND U37371 ( .A(n37599), .B(n37600), .Z(n37598) );
  XOR U37372 ( .A(n37597), .B(n36758), .Z(n37600) );
  XNOR U37373 ( .A(p_input[3148]), .B(n37601), .Z(n36758) );
  AND U37374 ( .A(n735), .B(n37602), .Z(n37601) );
  XOR U37375 ( .A(p_input[3180]), .B(p_input[3148]), .Z(n37602) );
  XNOR U37376 ( .A(n36755), .B(n37597), .Z(n37599) );
  XOR U37377 ( .A(n37603), .B(n37604), .Z(n36755) );
  AND U37378 ( .A(n732), .B(n37605), .Z(n37604) );
  XOR U37379 ( .A(p_input[3116]), .B(p_input[3084]), .Z(n37605) );
  XOR U37380 ( .A(n37606), .B(n37607), .Z(n37597) );
  AND U37381 ( .A(n37608), .B(n37609), .Z(n37607) );
  XOR U37382 ( .A(n37606), .B(n36770), .Z(n37609) );
  XNOR U37383 ( .A(p_input[3147]), .B(n37610), .Z(n36770) );
  AND U37384 ( .A(n735), .B(n37611), .Z(n37610) );
  XOR U37385 ( .A(p_input[3179]), .B(p_input[3147]), .Z(n37611) );
  XNOR U37386 ( .A(n36767), .B(n37606), .Z(n37608) );
  XOR U37387 ( .A(n37612), .B(n37613), .Z(n36767) );
  AND U37388 ( .A(n732), .B(n37614), .Z(n37613) );
  XOR U37389 ( .A(p_input[3115]), .B(p_input[3083]), .Z(n37614) );
  XOR U37390 ( .A(n37615), .B(n37616), .Z(n37606) );
  AND U37391 ( .A(n37617), .B(n37618), .Z(n37616) );
  XOR U37392 ( .A(n37615), .B(n36782), .Z(n37618) );
  XNOR U37393 ( .A(p_input[3146]), .B(n37619), .Z(n36782) );
  AND U37394 ( .A(n735), .B(n37620), .Z(n37619) );
  XOR U37395 ( .A(p_input[3178]), .B(p_input[3146]), .Z(n37620) );
  XNOR U37396 ( .A(n36779), .B(n37615), .Z(n37617) );
  XOR U37397 ( .A(n37621), .B(n37622), .Z(n36779) );
  AND U37398 ( .A(n732), .B(n37623), .Z(n37622) );
  XOR U37399 ( .A(p_input[3114]), .B(p_input[3082]), .Z(n37623) );
  XOR U37400 ( .A(n37624), .B(n37625), .Z(n37615) );
  AND U37401 ( .A(n37626), .B(n37627), .Z(n37625) );
  XOR U37402 ( .A(n37624), .B(n36794), .Z(n37627) );
  XNOR U37403 ( .A(p_input[3145]), .B(n37628), .Z(n36794) );
  AND U37404 ( .A(n735), .B(n37629), .Z(n37628) );
  XOR U37405 ( .A(p_input[3177]), .B(p_input[3145]), .Z(n37629) );
  XNOR U37406 ( .A(n36791), .B(n37624), .Z(n37626) );
  XOR U37407 ( .A(n37630), .B(n37631), .Z(n36791) );
  AND U37408 ( .A(n732), .B(n37632), .Z(n37631) );
  XOR U37409 ( .A(p_input[3113]), .B(p_input[3081]), .Z(n37632) );
  XOR U37410 ( .A(n37633), .B(n37634), .Z(n37624) );
  AND U37411 ( .A(n37635), .B(n37636), .Z(n37634) );
  XOR U37412 ( .A(n37633), .B(n36806), .Z(n37636) );
  XNOR U37413 ( .A(p_input[3144]), .B(n37637), .Z(n36806) );
  AND U37414 ( .A(n735), .B(n37638), .Z(n37637) );
  XOR U37415 ( .A(p_input[3176]), .B(p_input[3144]), .Z(n37638) );
  XNOR U37416 ( .A(n36803), .B(n37633), .Z(n37635) );
  XOR U37417 ( .A(n37639), .B(n37640), .Z(n36803) );
  AND U37418 ( .A(n732), .B(n37641), .Z(n37640) );
  XOR U37419 ( .A(p_input[3112]), .B(p_input[3080]), .Z(n37641) );
  XOR U37420 ( .A(n37642), .B(n37643), .Z(n37633) );
  AND U37421 ( .A(n37644), .B(n37645), .Z(n37643) );
  XOR U37422 ( .A(n37642), .B(n36818), .Z(n37645) );
  XNOR U37423 ( .A(p_input[3143]), .B(n37646), .Z(n36818) );
  AND U37424 ( .A(n735), .B(n37647), .Z(n37646) );
  XOR U37425 ( .A(p_input[3175]), .B(p_input[3143]), .Z(n37647) );
  XNOR U37426 ( .A(n36815), .B(n37642), .Z(n37644) );
  XOR U37427 ( .A(n37648), .B(n37649), .Z(n36815) );
  AND U37428 ( .A(n732), .B(n37650), .Z(n37649) );
  XOR U37429 ( .A(p_input[3111]), .B(p_input[3079]), .Z(n37650) );
  XOR U37430 ( .A(n37651), .B(n37652), .Z(n37642) );
  AND U37431 ( .A(n37653), .B(n37654), .Z(n37652) );
  XOR U37432 ( .A(n37651), .B(n36830), .Z(n37654) );
  XNOR U37433 ( .A(p_input[3142]), .B(n37655), .Z(n36830) );
  AND U37434 ( .A(n735), .B(n37656), .Z(n37655) );
  XOR U37435 ( .A(p_input[3174]), .B(p_input[3142]), .Z(n37656) );
  XNOR U37436 ( .A(n36827), .B(n37651), .Z(n37653) );
  XOR U37437 ( .A(n37657), .B(n37658), .Z(n36827) );
  AND U37438 ( .A(n732), .B(n37659), .Z(n37658) );
  XOR U37439 ( .A(p_input[3110]), .B(p_input[3078]), .Z(n37659) );
  XOR U37440 ( .A(n37660), .B(n37661), .Z(n37651) );
  AND U37441 ( .A(n37662), .B(n37663), .Z(n37661) );
  XOR U37442 ( .A(n37660), .B(n36842), .Z(n37663) );
  XNOR U37443 ( .A(p_input[3141]), .B(n37664), .Z(n36842) );
  AND U37444 ( .A(n735), .B(n37665), .Z(n37664) );
  XOR U37445 ( .A(p_input[3173]), .B(p_input[3141]), .Z(n37665) );
  XNOR U37446 ( .A(n36839), .B(n37660), .Z(n37662) );
  XOR U37447 ( .A(n37666), .B(n37667), .Z(n36839) );
  AND U37448 ( .A(n732), .B(n37668), .Z(n37667) );
  XOR U37449 ( .A(p_input[3109]), .B(p_input[3077]), .Z(n37668) );
  XOR U37450 ( .A(n37669), .B(n37670), .Z(n37660) );
  AND U37451 ( .A(n37671), .B(n37672), .Z(n37670) );
  XOR U37452 ( .A(n37669), .B(n36854), .Z(n37672) );
  XNOR U37453 ( .A(p_input[3140]), .B(n37673), .Z(n36854) );
  AND U37454 ( .A(n735), .B(n37674), .Z(n37673) );
  XOR U37455 ( .A(p_input[3172]), .B(p_input[3140]), .Z(n37674) );
  XNOR U37456 ( .A(n36851), .B(n37669), .Z(n37671) );
  XOR U37457 ( .A(n37675), .B(n37676), .Z(n36851) );
  AND U37458 ( .A(n732), .B(n37677), .Z(n37676) );
  XOR U37459 ( .A(p_input[3108]), .B(p_input[3076]), .Z(n37677) );
  XOR U37460 ( .A(n37678), .B(n37679), .Z(n37669) );
  AND U37461 ( .A(n37680), .B(n37681), .Z(n37679) );
  XOR U37462 ( .A(n37678), .B(n36866), .Z(n37681) );
  XNOR U37463 ( .A(p_input[3139]), .B(n37682), .Z(n36866) );
  AND U37464 ( .A(n735), .B(n37683), .Z(n37682) );
  XOR U37465 ( .A(p_input[3171]), .B(p_input[3139]), .Z(n37683) );
  XNOR U37466 ( .A(n36863), .B(n37678), .Z(n37680) );
  XOR U37467 ( .A(n37684), .B(n37685), .Z(n36863) );
  AND U37468 ( .A(n732), .B(n37686), .Z(n37685) );
  XOR U37469 ( .A(p_input[3107]), .B(p_input[3075]), .Z(n37686) );
  XOR U37470 ( .A(n37687), .B(n37688), .Z(n37678) );
  AND U37471 ( .A(n37689), .B(n37690), .Z(n37688) );
  XOR U37472 ( .A(n37687), .B(n36878), .Z(n37690) );
  XNOR U37473 ( .A(p_input[3138]), .B(n37691), .Z(n36878) );
  AND U37474 ( .A(n735), .B(n37692), .Z(n37691) );
  XOR U37475 ( .A(p_input[3170]), .B(p_input[3138]), .Z(n37692) );
  XNOR U37476 ( .A(n36875), .B(n37687), .Z(n37689) );
  XOR U37477 ( .A(n37693), .B(n37694), .Z(n36875) );
  AND U37478 ( .A(n732), .B(n37695), .Z(n37694) );
  XOR U37479 ( .A(p_input[3106]), .B(p_input[3074]), .Z(n37695) );
  XOR U37480 ( .A(n37696), .B(n37697), .Z(n37687) );
  AND U37481 ( .A(n37698), .B(n37699), .Z(n37697) );
  XNOR U37482 ( .A(n37700), .B(n36891), .Z(n37699) );
  XNOR U37483 ( .A(p_input[3137]), .B(n37701), .Z(n36891) );
  AND U37484 ( .A(n735), .B(n37702), .Z(n37701) );
  XNOR U37485 ( .A(p_input[3169]), .B(n37703), .Z(n37702) );
  IV U37486 ( .A(p_input[3137]), .Z(n37703) );
  XNOR U37487 ( .A(n36888), .B(n37696), .Z(n37698) );
  XNOR U37488 ( .A(p_input[3073]), .B(n37704), .Z(n36888) );
  AND U37489 ( .A(n732), .B(n37705), .Z(n37704) );
  XOR U37490 ( .A(p_input[3105]), .B(p_input[3073]), .Z(n37705) );
  IV U37491 ( .A(n37700), .Z(n37696) );
  AND U37492 ( .A(n37426), .B(n37429), .Z(n37700) );
  XOR U37493 ( .A(p_input[3136]), .B(n37706), .Z(n37429) );
  AND U37494 ( .A(n735), .B(n37707), .Z(n37706) );
  XOR U37495 ( .A(p_input[3168]), .B(p_input[3136]), .Z(n37707) );
  XOR U37496 ( .A(n37708), .B(n37709), .Z(n735) );
  AND U37497 ( .A(n37710), .B(n37711), .Z(n37709) );
  XNOR U37498 ( .A(p_input[3199]), .B(n37708), .Z(n37711) );
  XOR U37499 ( .A(n37708), .B(p_input[3167]), .Z(n37710) );
  XOR U37500 ( .A(n37712), .B(n37713), .Z(n37708) );
  AND U37501 ( .A(n37714), .B(n37715), .Z(n37713) );
  XNOR U37502 ( .A(p_input[3198]), .B(n37712), .Z(n37715) );
  XOR U37503 ( .A(n37712), .B(p_input[3166]), .Z(n37714) );
  XOR U37504 ( .A(n37716), .B(n37717), .Z(n37712) );
  AND U37505 ( .A(n37718), .B(n37719), .Z(n37717) );
  XNOR U37506 ( .A(p_input[3197]), .B(n37716), .Z(n37719) );
  XOR U37507 ( .A(n37716), .B(p_input[3165]), .Z(n37718) );
  XOR U37508 ( .A(n37720), .B(n37721), .Z(n37716) );
  AND U37509 ( .A(n37722), .B(n37723), .Z(n37721) );
  XNOR U37510 ( .A(p_input[3196]), .B(n37720), .Z(n37723) );
  XOR U37511 ( .A(n37720), .B(p_input[3164]), .Z(n37722) );
  XOR U37512 ( .A(n37724), .B(n37725), .Z(n37720) );
  AND U37513 ( .A(n37726), .B(n37727), .Z(n37725) );
  XNOR U37514 ( .A(p_input[3195]), .B(n37724), .Z(n37727) );
  XOR U37515 ( .A(n37724), .B(p_input[3163]), .Z(n37726) );
  XOR U37516 ( .A(n37728), .B(n37729), .Z(n37724) );
  AND U37517 ( .A(n37730), .B(n37731), .Z(n37729) );
  XNOR U37518 ( .A(p_input[3194]), .B(n37728), .Z(n37731) );
  XOR U37519 ( .A(n37728), .B(p_input[3162]), .Z(n37730) );
  XOR U37520 ( .A(n37732), .B(n37733), .Z(n37728) );
  AND U37521 ( .A(n37734), .B(n37735), .Z(n37733) );
  XNOR U37522 ( .A(p_input[3193]), .B(n37732), .Z(n37735) );
  XOR U37523 ( .A(n37732), .B(p_input[3161]), .Z(n37734) );
  XOR U37524 ( .A(n37736), .B(n37737), .Z(n37732) );
  AND U37525 ( .A(n37738), .B(n37739), .Z(n37737) );
  XNOR U37526 ( .A(p_input[3192]), .B(n37736), .Z(n37739) );
  XOR U37527 ( .A(n37736), .B(p_input[3160]), .Z(n37738) );
  XOR U37528 ( .A(n37740), .B(n37741), .Z(n37736) );
  AND U37529 ( .A(n37742), .B(n37743), .Z(n37741) );
  XNOR U37530 ( .A(p_input[3191]), .B(n37740), .Z(n37743) );
  XOR U37531 ( .A(n37740), .B(p_input[3159]), .Z(n37742) );
  XOR U37532 ( .A(n37744), .B(n37745), .Z(n37740) );
  AND U37533 ( .A(n37746), .B(n37747), .Z(n37745) );
  XNOR U37534 ( .A(p_input[3190]), .B(n37744), .Z(n37747) );
  XOR U37535 ( .A(n37744), .B(p_input[3158]), .Z(n37746) );
  XOR U37536 ( .A(n37748), .B(n37749), .Z(n37744) );
  AND U37537 ( .A(n37750), .B(n37751), .Z(n37749) );
  XNOR U37538 ( .A(p_input[3189]), .B(n37748), .Z(n37751) );
  XOR U37539 ( .A(n37748), .B(p_input[3157]), .Z(n37750) );
  XOR U37540 ( .A(n37752), .B(n37753), .Z(n37748) );
  AND U37541 ( .A(n37754), .B(n37755), .Z(n37753) );
  XNOR U37542 ( .A(p_input[3188]), .B(n37752), .Z(n37755) );
  XOR U37543 ( .A(n37752), .B(p_input[3156]), .Z(n37754) );
  XOR U37544 ( .A(n37756), .B(n37757), .Z(n37752) );
  AND U37545 ( .A(n37758), .B(n37759), .Z(n37757) );
  XNOR U37546 ( .A(p_input[3187]), .B(n37756), .Z(n37759) );
  XOR U37547 ( .A(n37756), .B(p_input[3155]), .Z(n37758) );
  XOR U37548 ( .A(n37760), .B(n37761), .Z(n37756) );
  AND U37549 ( .A(n37762), .B(n37763), .Z(n37761) );
  XNOR U37550 ( .A(p_input[3186]), .B(n37760), .Z(n37763) );
  XOR U37551 ( .A(n37760), .B(p_input[3154]), .Z(n37762) );
  XOR U37552 ( .A(n37764), .B(n37765), .Z(n37760) );
  AND U37553 ( .A(n37766), .B(n37767), .Z(n37765) );
  XNOR U37554 ( .A(p_input[3185]), .B(n37764), .Z(n37767) );
  XOR U37555 ( .A(n37764), .B(p_input[3153]), .Z(n37766) );
  XOR U37556 ( .A(n37768), .B(n37769), .Z(n37764) );
  AND U37557 ( .A(n37770), .B(n37771), .Z(n37769) );
  XNOR U37558 ( .A(p_input[3184]), .B(n37768), .Z(n37771) );
  XOR U37559 ( .A(n37768), .B(p_input[3152]), .Z(n37770) );
  XOR U37560 ( .A(n37772), .B(n37773), .Z(n37768) );
  AND U37561 ( .A(n37774), .B(n37775), .Z(n37773) );
  XNOR U37562 ( .A(p_input[3183]), .B(n37772), .Z(n37775) );
  XOR U37563 ( .A(n37772), .B(p_input[3151]), .Z(n37774) );
  XOR U37564 ( .A(n37776), .B(n37777), .Z(n37772) );
  AND U37565 ( .A(n37778), .B(n37779), .Z(n37777) );
  XNOR U37566 ( .A(p_input[3182]), .B(n37776), .Z(n37779) );
  XOR U37567 ( .A(n37776), .B(p_input[3150]), .Z(n37778) );
  XOR U37568 ( .A(n37780), .B(n37781), .Z(n37776) );
  AND U37569 ( .A(n37782), .B(n37783), .Z(n37781) );
  XNOR U37570 ( .A(p_input[3181]), .B(n37780), .Z(n37783) );
  XOR U37571 ( .A(n37780), .B(p_input[3149]), .Z(n37782) );
  XOR U37572 ( .A(n37784), .B(n37785), .Z(n37780) );
  AND U37573 ( .A(n37786), .B(n37787), .Z(n37785) );
  XNOR U37574 ( .A(p_input[3180]), .B(n37784), .Z(n37787) );
  XOR U37575 ( .A(n37784), .B(p_input[3148]), .Z(n37786) );
  XOR U37576 ( .A(n37788), .B(n37789), .Z(n37784) );
  AND U37577 ( .A(n37790), .B(n37791), .Z(n37789) );
  XNOR U37578 ( .A(p_input[3179]), .B(n37788), .Z(n37791) );
  XOR U37579 ( .A(n37788), .B(p_input[3147]), .Z(n37790) );
  XOR U37580 ( .A(n37792), .B(n37793), .Z(n37788) );
  AND U37581 ( .A(n37794), .B(n37795), .Z(n37793) );
  XNOR U37582 ( .A(p_input[3178]), .B(n37792), .Z(n37795) );
  XOR U37583 ( .A(n37792), .B(p_input[3146]), .Z(n37794) );
  XOR U37584 ( .A(n37796), .B(n37797), .Z(n37792) );
  AND U37585 ( .A(n37798), .B(n37799), .Z(n37797) );
  XNOR U37586 ( .A(p_input[3177]), .B(n37796), .Z(n37799) );
  XOR U37587 ( .A(n37796), .B(p_input[3145]), .Z(n37798) );
  XOR U37588 ( .A(n37800), .B(n37801), .Z(n37796) );
  AND U37589 ( .A(n37802), .B(n37803), .Z(n37801) );
  XNOR U37590 ( .A(p_input[3176]), .B(n37800), .Z(n37803) );
  XOR U37591 ( .A(n37800), .B(p_input[3144]), .Z(n37802) );
  XOR U37592 ( .A(n37804), .B(n37805), .Z(n37800) );
  AND U37593 ( .A(n37806), .B(n37807), .Z(n37805) );
  XNOR U37594 ( .A(p_input[3175]), .B(n37804), .Z(n37807) );
  XOR U37595 ( .A(n37804), .B(p_input[3143]), .Z(n37806) );
  XOR U37596 ( .A(n37808), .B(n37809), .Z(n37804) );
  AND U37597 ( .A(n37810), .B(n37811), .Z(n37809) );
  XNOR U37598 ( .A(p_input[3174]), .B(n37808), .Z(n37811) );
  XOR U37599 ( .A(n37808), .B(p_input[3142]), .Z(n37810) );
  XOR U37600 ( .A(n37812), .B(n37813), .Z(n37808) );
  AND U37601 ( .A(n37814), .B(n37815), .Z(n37813) );
  XNOR U37602 ( .A(p_input[3173]), .B(n37812), .Z(n37815) );
  XOR U37603 ( .A(n37812), .B(p_input[3141]), .Z(n37814) );
  XOR U37604 ( .A(n37816), .B(n37817), .Z(n37812) );
  AND U37605 ( .A(n37818), .B(n37819), .Z(n37817) );
  XNOR U37606 ( .A(p_input[3172]), .B(n37816), .Z(n37819) );
  XOR U37607 ( .A(n37816), .B(p_input[3140]), .Z(n37818) );
  XOR U37608 ( .A(n37820), .B(n37821), .Z(n37816) );
  AND U37609 ( .A(n37822), .B(n37823), .Z(n37821) );
  XNOR U37610 ( .A(p_input[3171]), .B(n37820), .Z(n37823) );
  XOR U37611 ( .A(n37820), .B(p_input[3139]), .Z(n37822) );
  XOR U37612 ( .A(n37824), .B(n37825), .Z(n37820) );
  AND U37613 ( .A(n37826), .B(n37827), .Z(n37825) );
  XNOR U37614 ( .A(p_input[3170]), .B(n37824), .Z(n37827) );
  XOR U37615 ( .A(n37824), .B(p_input[3138]), .Z(n37826) );
  XNOR U37616 ( .A(n37828), .B(n37829), .Z(n37824) );
  AND U37617 ( .A(n37830), .B(n37831), .Z(n37829) );
  XOR U37618 ( .A(p_input[3169]), .B(n37828), .Z(n37831) );
  XNOR U37619 ( .A(p_input[3137]), .B(n37828), .Z(n37830) );
  AND U37620 ( .A(p_input[3168]), .B(n37832), .Z(n37828) );
  IV U37621 ( .A(p_input[3136]), .Z(n37832) );
  XNOR U37622 ( .A(p_input[3072]), .B(n37833), .Z(n37426) );
  AND U37623 ( .A(n732), .B(n37834), .Z(n37833) );
  XOR U37624 ( .A(p_input[3104]), .B(p_input[3072]), .Z(n37834) );
  XOR U37625 ( .A(n37835), .B(n37836), .Z(n732) );
  AND U37626 ( .A(n37837), .B(n37838), .Z(n37836) );
  XNOR U37627 ( .A(p_input[3135]), .B(n37835), .Z(n37838) );
  XOR U37628 ( .A(n37835), .B(p_input[3103]), .Z(n37837) );
  XOR U37629 ( .A(n37839), .B(n37840), .Z(n37835) );
  AND U37630 ( .A(n37841), .B(n37842), .Z(n37840) );
  XNOR U37631 ( .A(p_input[3134]), .B(n37839), .Z(n37842) );
  XNOR U37632 ( .A(n37839), .B(n37441), .Z(n37841) );
  IV U37633 ( .A(p_input[3102]), .Z(n37441) );
  XOR U37634 ( .A(n37843), .B(n37844), .Z(n37839) );
  AND U37635 ( .A(n37845), .B(n37846), .Z(n37844) );
  XNOR U37636 ( .A(p_input[3133]), .B(n37843), .Z(n37846) );
  XNOR U37637 ( .A(n37843), .B(n37450), .Z(n37845) );
  IV U37638 ( .A(p_input[3101]), .Z(n37450) );
  XOR U37639 ( .A(n37847), .B(n37848), .Z(n37843) );
  AND U37640 ( .A(n37849), .B(n37850), .Z(n37848) );
  XNOR U37641 ( .A(p_input[3132]), .B(n37847), .Z(n37850) );
  XNOR U37642 ( .A(n37847), .B(n37459), .Z(n37849) );
  IV U37643 ( .A(p_input[3100]), .Z(n37459) );
  XOR U37644 ( .A(n37851), .B(n37852), .Z(n37847) );
  AND U37645 ( .A(n37853), .B(n37854), .Z(n37852) );
  XNOR U37646 ( .A(p_input[3131]), .B(n37851), .Z(n37854) );
  XNOR U37647 ( .A(n37851), .B(n37468), .Z(n37853) );
  IV U37648 ( .A(p_input[3099]), .Z(n37468) );
  XOR U37649 ( .A(n37855), .B(n37856), .Z(n37851) );
  AND U37650 ( .A(n37857), .B(n37858), .Z(n37856) );
  XNOR U37651 ( .A(p_input[3130]), .B(n37855), .Z(n37858) );
  XNOR U37652 ( .A(n37855), .B(n37477), .Z(n37857) );
  IV U37653 ( .A(p_input[3098]), .Z(n37477) );
  XOR U37654 ( .A(n37859), .B(n37860), .Z(n37855) );
  AND U37655 ( .A(n37861), .B(n37862), .Z(n37860) );
  XNOR U37656 ( .A(p_input[3129]), .B(n37859), .Z(n37862) );
  XNOR U37657 ( .A(n37859), .B(n37486), .Z(n37861) );
  IV U37658 ( .A(p_input[3097]), .Z(n37486) );
  XOR U37659 ( .A(n37863), .B(n37864), .Z(n37859) );
  AND U37660 ( .A(n37865), .B(n37866), .Z(n37864) );
  XNOR U37661 ( .A(p_input[3128]), .B(n37863), .Z(n37866) );
  XNOR U37662 ( .A(n37863), .B(n37495), .Z(n37865) );
  IV U37663 ( .A(p_input[3096]), .Z(n37495) );
  XOR U37664 ( .A(n37867), .B(n37868), .Z(n37863) );
  AND U37665 ( .A(n37869), .B(n37870), .Z(n37868) );
  XNOR U37666 ( .A(p_input[3127]), .B(n37867), .Z(n37870) );
  XNOR U37667 ( .A(n37867), .B(n37504), .Z(n37869) );
  IV U37668 ( .A(p_input[3095]), .Z(n37504) );
  XOR U37669 ( .A(n37871), .B(n37872), .Z(n37867) );
  AND U37670 ( .A(n37873), .B(n37874), .Z(n37872) );
  XNOR U37671 ( .A(p_input[3126]), .B(n37871), .Z(n37874) );
  XNOR U37672 ( .A(n37871), .B(n37513), .Z(n37873) );
  IV U37673 ( .A(p_input[3094]), .Z(n37513) );
  XOR U37674 ( .A(n37875), .B(n37876), .Z(n37871) );
  AND U37675 ( .A(n37877), .B(n37878), .Z(n37876) );
  XNOR U37676 ( .A(p_input[3125]), .B(n37875), .Z(n37878) );
  XNOR U37677 ( .A(n37875), .B(n37522), .Z(n37877) );
  IV U37678 ( .A(p_input[3093]), .Z(n37522) );
  XOR U37679 ( .A(n37879), .B(n37880), .Z(n37875) );
  AND U37680 ( .A(n37881), .B(n37882), .Z(n37880) );
  XNOR U37681 ( .A(p_input[3124]), .B(n37879), .Z(n37882) );
  XNOR U37682 ( .A(n37879), .B(n37531), .Z(n37881) );
  IV U37683 ( .A(p_input[3092]), .Z(n37531) );
  XOR U37684 ( .A(n37883), .B(n37884), .Z(n37879) );
  AND U37685 ( .A(n37885), .B(n37886), .Z(n37884) );
  XNOR U37686 ( .A(p_input[3123]), .B(n37883), .Z(n37886) );
  XNOR U37687 ( .A(n37883), .B(n37540), .Z(n37885) );
  IV U37688 ( .A(p_input[3091]), .Z(n37540) );
  XOR U37689 ( .A(n37887), .B(n37888), .Z(n37883) );
  AND U37690 ( .A(n37889), .B(n37890), .Z(n37888) );
  XNOR U37691 ( .A(p_input[3122]), .B(n37887), .Z(n37890) );
  XNOR U37692 ( .A(n37887), .B(n37549), .Z(n37889) );
  IV U37693 ( .A(p_input[3090]), .Z(n37549) );
  XOR U37694 ( .A(n37891), .B(n37892), .Z(n37887) );
  AND U37695 ( .A(n37893), .B(n37894), .Z(n37892) );
  XNOR U37696 ( .A(p_input[3121]), .B(n37891), .Z(n37894) );
  XNOR U37697 ( .A(n37891), .B(n37558), .Z(n37893) );
  IV U37698 ( .A(p_input[3089]), .Z(n37558) );
  XOR U37699 ( .A(n37895), .B(n37896), .Z(n37891) );
  AND U37700 ( .A(n37897), .B(n37898), .Z(n37896) );
  XNOR U37701 ( .A(p_input[3120]), .B(n37895), .Z(n37898) );
  XNOR U37702 ( .A(n37895), .B(n37567), .Z(n37897) );
  IV U37703 ( .A(p_input[3088]), .Z(n37567) );
  XOR U37704 ( .A(n37899), .B(n37900), .Z(n37895) );
  AND U37705 ( .A(n37901), .B(n37902), .Z(n37900) );
  XNOR U37706 ( .A(p_input[3119]), .B(n37899), .Z(n37902) );
  XNOR U37707 ( .A(n37899), .B(n37576), .Z(n37901) );
  IV U37708 ( .A(p_input[3087]), .Z(n37576) );
  XOR U37709 ( .A(n37903), .B(n37904), .Z(n37899) );
  AND U37710 ( .A(n37905), .B(n37906), .Z(n37904) );
  XNOR U37711 ( .A(p_input[3118]), .B(n37903), .Z(n37906) );
  XNOR U37712 ( .A(n37903), .B(n37585), .Z(n37905) );
  IV U37713 ( .A(p_input[3086]), .Z(n37585) );
  XOR U37714 ( .A(n37907), .B(n37908), .Z(n37903) );
  AND U37715 ( .A(n37909), .B(n37910), .Z(n37908) );
  XNOR U37716 ( .A(p_input[3117]), .B(n37907), .Z(n37910) );
  XNOR U37717 ( .A(n37907), .B(n37594), .Z(n37909) );
  IV U37718 ( .A(p_input[3085]), .Z(n37594) );
  XOR U37719 ( .A(n37911), .B(n37912), .Z(n37907) );
  AND U37720 ( .A(n37913), .B(n37914), .Z(n37912) );
  XNOR U37721 ( .A(p_input[3116]), .B(n37911), .Z(n37914) );
  XNOR U37722 ( .A(n37911), .B(n37603), .Z(n37913) );
  IV U37723 ( .A(p_input[3084]), .Z(n37603) );
  XOR U37724 ( .A(n37915), .B(n37916), .Z(n37911) );
  AND U37725 ( .A(n37917), .B(n37918), .Z(n37916) );
  XNOR U37726 ( .A(p_input[3115]), .B(n37915), .Z(n37918) );
  XNOR U37727 ( .A(n37915), .B(n37612), .Z(n37917) );
  IV U37728 ( .A(p_input[3083]), .Z(n37612) );
  XOR U37729 ( .A(n37919), .B(n37920), .Z(n37915) );
  AND U37730 ( .A(n37921), .B(n37922), .Z(n37920) );
  XNOR U37731 ( .A(p_input[3114]), .B(n37919), .Z(n37922) );
  XNOR U37732 ( .A(n37919), .B(n37621), .Z(n37921) );
  IV U37733 ( .A(p_input[3082]), .Z(n37621) );
  XOR U37734 ( .A(n37923), .B(n37924), .Z(n37919) );
  AND U37735 ( .A(n37925), .B(n37926), .Z(n37924) );
  XNOR U37736 ( .A(p_input[3113]), .B(n37923), .Z(n37926) );
  XNOR U37737 ( .A(n37923), .B(n37630), .Z(n37925) );
  IV U37738 ( .A(p_input[3081]), .Z(n37630) );
  XOR U37739 ( .A(n37927), .B(n37928), .Z(n37923) );
  AND U37740 ( .A(n37929), .B(n37930), .Z(n37928) );
  XNOR U37741 ( .A(p_input[3112]), .B(n37927), .Z(n37930) );
  XNOR U37742 ( .A(n37927), .B(n37639), .Z(n37929) );
  IV U37743 ( .A(p_input[3080]), .Z(n37639) );
  XOR U37744 ( .A(n37931), .B(n37932), .Z(n37927) );
  AND U37745 ( .A(n37933), .B(n37934), .Z(n37932) );
  XNOR U37746 ( .A(p_input[3111]), .B(n37931), .Z(n37934) );
  XNOR U37747 ( .A(n37931), .B(n37648), .Z(n37933) );
  IV U37748 ( .A(p_input[3079]), .Z(n37648) );
  XOR U37749 ( .A(n37935), .B(n37936), .Z(n37931) );
  AND U37750 ( .A(n37937), .B(n37938), .Z(n37936) );
  XNOR U37751 ( .A(p_input[3110]), .B(n37935), .Z(n37938) );
  XNOR U37752 ( .A(n37935), .B(n37657), .Z(n37937) );
  IV U37753 ( .A(p_input[3078]), .Z(n37657) );
  XOR U37754 ( .A(n37939), .B(n37940), .Z(n37935) );
  AND U37755 ( .A(n37941), .B(n37942), .Z(n37940) );
  XNOR U37756 ( .A(p_input[3109]), .B(n37939), .Z(n37942) );
  XNOR U37757 ( .A(n37939), .B(n37666), .Z(n37941) );
  IV U37758 ( .A(p_input[3077]), .Z(n37666) );
  XOR U37759 ( .A(n37943), .B(n37944), .Z(n37939) );
  AND U37760 ( .A(n37945), .B(n37946), .Z(n37944) );
  XNOR U37761 ( .A(p_input[3108]), .B(n37943), .Z(n37946) );
  XNOR U37762 ( .A(n37943), .B(n37675), .Z(n37945) );
  IV U37763 ( .A(p_input[3076]), .Z(n37675) );
  XOR U37764 ( .A(n37947), .B(n37948), .Z(n37943) );
  AND U37765 ( .A(n37949), .B(n37950), .Z(n37948) );
  XNOR U37766 ( .A(p_input[3107]), .B(n37947), .Z(n37950) );
  XNOR U37767 ( .A(n37947), .B(n37684), .Z(n37949) );
  IV U37768 ( .A(p_input[3075]), .Z(n37684) );
  XOR U37769 ( .A(n37951), .B(n37952), .Z(n37947) );
  AND U37770 ( .A(n37953), .B(n37954), .Z(n37952) );
  XNOR U37771 ( .A(p_input[3106]), .B(n37951), .Z(n37954) );
  XNOR U37772 ( .A(n37951), .B(n37693), .Z(n37953) );
  IV U37773 ( .A(p_input[3074]), .Z(n37693) );
  XNOR U37774 ( .A(n37955), .B(n37956), .Z(n37951) );
  AND U37775 ( .A(n37957), .B(n37958), .Z(n37956) );
  XOR U37776 ( .A(p_input[3105]), .B(n37955), .Z(n37958) );
  XNOR U37777 ( .A(p_input[3073]), .B(n37955), .Z(n37957) );
  AND U37778 ( .A(p_input[3104]), .B(n37959), .Z(n37955) );
  IV U37779 ( .A(p_input[3072]), .Z(n37959) );
  XOR U37780 ( .A(n37960), .B(n37961), .Z(n30672) );
  AND U37781 ( .A(n1097), .B(n37962), .Z(n37961) );
  XNOR U37782 ( .A(n37963), .B(n37960), .Z(n37962) );
  XOR U37783 ( .A(n37964), .B(n37965), .Z(n1097) );
  AND U37784 ( .A(n37966), .B(n37967), .Z(n37965) );
  XOR U37785 ( .A(n37964), .B(n30687), .Z(n37967) );
  XOR U37786 ( .A(n37968), .B(n37969), .Z(n30687) );
  AND U37787 ( .A(n1031), .B(n37970), .Z(n37969) );
  XOR U37788 ( .A(n37971), .B(n37968), .Z(n37970) );
  XNOR U37789 ( .A(n30684), .B(n37964), .Z(n37966) );
  XOR U37790 ( .A(n37972), .B(n37973), .Z(n30684) );
  AND U37791 ( .A(n1028), .B(n37974), .Z(n37973) );
  XOR U37792 ( .A(n37975), .B(n37972), .Z(n37974) );
  XOR U37793 ( .A(n37976), .B(n37977), .Z(n37964) );
  AND U37794 ( .A(n37978), .B(n37979), .Z(n37977) );
  XOR U37795 ( .A(n37976), .B(n30699), .Z(n37979) );
  XOR U37796 ( .A(n37980), .B(n37981), .Z(n30699) );
  AND U37797 ( .A(n1031), .B(n37982), .Z(n37981) );
  XOR U37798 ( .A(n37983), .B(n37980), .Z(n37982) );
  XNOR U37799 ( .A(n30696), .B(n37976), .Z(n37978) );
  XOR U37800 ( .A(n37984), .B(n37985), .Z(n30696) );
  AND U37801 ( .A(n1028), .B(n37986), .Z(n37985) );
  XOR U37802 ( .A(n37987), .B(n37984), .Z(n37986) );
  XOR U37803 ( .A(n37988), .B(n37989), .Z(n37976) );
  AND U37804 ( .A(n37990), .B(n37991), .Z(n37989) );
  XOR U37805 ( .A(n37988), .B(n30711), .Z(n37991) );
  XOR U37806 ( .A(n37992), .B(n37993), .Z(n30711) );
  AND U37807 ( .A(n1031), .B(n37994), .Z(n37993) );
  XOR U37808 ( .A(n37995), .B(n37992), .Z(n37994) );
  XNOR U37809 ( .A(n30708), .B(n37988), .Z(n37990) );
  XOR U37810 ( .A(n37996), .B(n37997), .Z(n30708) );
  AND U37811 ( .A(n1028), .B(n37998), .Z(n37997) );
  XOR U37812 ( .A(n37999), .B(n37996), .Z(n37998) );
  XOR U37813 ( .A(n38000), .B(n38001), .Z(n37988) );
  AND U37814 ( .A(n38002), .B(n38003), .Z(n38001) );
  XOR U37815 ( .A(n38000), .B(n30723), .Z(n38003) );
  XOR U37816 ( .A(n38004), .B(n38005), .Z(n30723) );
  AND U37817 ( .A(n1031), .B(n38006), .Z(n38005) );
  XOR U37818 ( .A(n38007), .B(n38004), .Z(n38006) );
  XNOR U37819 ( .A(n30720), .B(n38000), .Z(n38002) );
  XOR U37820 ( .A(n38008), .B(n38009), .Z(n30720) );
  AND U37821 ( .A(n1028), .B(n38010), .Z(n38009) );
  XOR U37822 ( .A(n38011), .B(n38008), .Z(n38010) );
  XOR U37823 ( .A(n38012), .B(n38013), .Z(n38000) );
  AND U37824 ( .A(n38014), .B(n38015), .Z(n38013) );
  XOR U37825 ( .A(n38012), .B(n30735), .Z(n38015) );
  XOR U37826 ( .A(n38016), .B(n38017), .Z(n30735) );
  AND U37827 ( .A(n1031), .B(n38018), .Z(n38017) );
  XOR U37828 ( .A(n38019), .B(n38016), .Z(n38018) );
  XNOR U37829 ( .A(n30732), .B(n38012), .Z(n38014) );
  XOR U37830 ( .A(n38020), .B(n38021), .Z(n30732) );
  AND U37831 ( .A(n1028), .B(n38022), .Z(n38021) );
  XOR U37832 ( .A(n38023), .B(n38020), .Z(n38022) );
  XOR U37833 ( .A(n38024), .B(n38025), .Z(n38012) );
  AND U37834 ( .A(n38026), .B(n38027), .Z(n38025) );
  XOR U37835 ( .A(n38024), .B(n30747), .Z(n38027) );
  XOR U37836 ( .A(n38028), .B(n38029), .Z(n30747) );
  AND U37837 ( .A(n1031), .B(n38030), .Z(n38029) );
  XOR U37838 ( .A(n38031), .B(n38028), .Z(n38030) );
  XNOR U37839 ( .A(n30744), .B(n38024), .Z(n38026) );
  XOR U37840 ( .A(n38032), .B(n38033), .Z(n30744) );
  AND U37841 ( .A(n1028), .B(n38034), .Z(n38033) );
  XOR U37842 ( .A(n38035), .B(n38032), .Z(n38034) );
  XOR U37843 ( .A(n38036), .B(n38037), .Z(n38024) );
  AND U37844 ( .A(n38038), .B(n38039), .Z(n38037) );
  XOR U37845 ( .A(n38036), .B(n30759), .Z(n38039) );
  XOR U37846 ( .A(n38040), .B(n38041), .Z(n30759) );
  AND U37847 ( .A(n1031), .B(n38042), .Z(n38041) );
  XOR U37848 ( .A(n38043), .B(n38040), .Z(n38042) );
  XNOR U37849 ( .A(n30756), .B(n38036), .Z(n38038) );
  XOR U37850 ( .A(n38044), .B(n38045), .Z(n30756) );
  AND U37851 ( .A(n1028), .B(n38046), .Z(n38045) );
  XOR U37852 ( .A(n38047), .B(n38044), .Z(n38046) );
  XOR U37853 ( .A(n38048), .B(n38049), .Z(n38036) );
  AND U37854 ( .A(n38050), .B(n38051), .Z(n38049) );
  XOR U37855 ( .A(n38048), .B(n30771), .Z(n38051) );
  XOR U37856 ( .A(n38052), .B(n38053), .Z(n30771) );
  AND U37857 ( .A(n1031), .B(n38054), .Z(n38053) );
  XOR U37858 ( .A(n38055), .B(n38052), .Z(n38054) );
  XNOR U37859 ( .A(n30768), .B(n38048), .Z(n38050) );
  XOR U37860 ( .A(n38056), .B(n38057), .Z(n30768) );
  AND U37861 ( .A(n1028), .B(n38058), .Z(n38057) );
  XOR U37862 ( .A(n38059), .B(n38056), .Z(n38058) );
  XOR U37863 ( .A(n38060), .B(n38061), .Z(n38048) );
  AND U37864 ( .A(n38062), .B(n38063), .Z(n38061) );
  XOR U37865 ( .A(n38060), .B(n30783), .Z(n38063) );
  XOR U37866 ( .A(n38064), .B(n38065), .Z(n30783) );
  AND U37867 ( .A(n1031), .B(n38066), .Z(n38065) );
  XOR U37868 ( .A(n38067), .B(n38064), .Z(n38066) );
  XNOR U37869 ( .A(n30780), .B(n38060), .Z(n38062) );
  XOR U37870 ( .A(n38068), .B(n38069), .Z(n30780) );
  AND U37871 ( .A(n1028), .B(n38070), .Z(n38069) );
  XOR U37872 ( .A(n38071), .B(n38068), .Z(n38070) );
  XOR U37873 ( .A(n38072), .B(n38073), .Z(n38060) );
  AND U37874 ( .A(n38074), .B(n38075), .Z(n38073) );
  XOR U37875 ( .A(n38072), .B(n30795), .Z(n38075) );
  XOR U37876 ( .A(n38076), .B(n38077), .Z(n30795) );
  AND U37877 ( .A(n1031), .B(n38078), .Z(n38077) );
  XOR U37878 ( .A(n38079), .B(n38076), .Z(n38078) );
  XNOR U37879 ( .A(n30792), .B(n38072), .Z(n38074) );
  XOR U37880 ( .A(n38080), .B(n38081), .Z(n30792) );
  AND U37881 ( .A(n1028), .B(n38082), .Z(n38081) );
  XOR U37882 ( .A(n38083), .B(n38080), .Z(n38082) );
  XOR U37883 ( .A(n38084), .B(n38085), .Z(n38072) );
  AND U37884 ( .A(n38086), .B(n38087), .Z(n38085) );
  XOR U37885 ( .A(n38084), .B(n30807), .Z(n38087) );
  XOR U37886 ( .A(n38088), .B(n38089), .Z(n30807) );
  AND U37887 ( .A(n1031), .B(n38090), .Z(n38089) );
  XOR U37888 ( .A(n38091), .B(n38088), .Z(n38090) );
  XNOR U37889 ( .A(n30804), .B(n38084), .Z(n38086) );
  XOR U37890 ( .A(n38092), .B(n38093), .Z(n30804) );
  AND U37891 ( .A(n1028), .B(n38094), .Z(n38093) );
  XOR U37892 ( .A(n38095), .B(n38092), .Z(n38094) );
  XOR U37893 ( .A(n38096), .B(n38097), .Z(n38084) );
  AND U37894 ( .A(n38098), .B(n38099), .Z(n38097) );
  XOR U37895 ( .A(n38096), .B(n30819), .Z(n38099) );
  XOR U37896 ( .A(n38100), .B(n38101), .Z(n30819) );
  AND U37897 ( .A(n1031), .B(n38102), .Z(n38101) );
  XOR U37898 ( .A(n38103), .B(n38100), .Z(n38102) );
  XNOR U37899 ( .A(n30816), .B(n38096), .Z(n38098) );
  XOR U37900 ( .A(n38104), .B(n38105), .Z(n30816) );
  AND U37901 ( .A(n1028), .B(n38106), .Z(n38105) );
  XOR U37902 ( .A(n38107), .B(n38104), .Z(n38106) );
  XOR U37903 ( .A(n38108), .B(n38109), .Z(n38096) );
  AND U37904 ( .A(n38110), .B(n38111), .Z(n38109) );
  XOR U37905 ( .A(n38108), .B(n30831), .Z(n38111) );
  XOR U37906 ( .A(n38112), .B(n38113), .Z(n30831) );
  AND U37907 ( .A(n1031), .B(n38114), .Z(n38113) );
  XOR U37908 ( .A(n38115), .B(n38112), .Z(n38114) );
  XNOR U37909 ( .A(n30828), .B(n38108), .Z(n38110) );
  XOR U37910 ( .A(n38116), .B(n38117), .Z(n30828) );
  AND U37911 ( .A(n1028), .B(n38118), .Z(n38117) );
  XOR U37912 ( .A(n38119), .B(n38116), .Z(n38118) );
  XOR U37913 ( .A(n38120), .B(n38121), .Z(n38108) );
  AND U37914 ( .A(n38122), .B(n38123), .Z(n38121) );
  XOR U37915 ( .A(n38120), .B(n30843), .Z(n38123) );
  XOR U37916 ( .A(n38124), .B(n38125), .Z(n30843) );
  AND U37917 ( .A(n1031), .B(n38126), .Z(n38125) );
  XOR U37918 ( .A(n38127), .B(n38124), .Z(n38126) );
  XNOR U37919 ( .A(n30840), .B(n38120), .Z(n38122) );
  XOR U37920 ( .A(n38128), .B(n38129), .Z(n30840) );
  AND U37921 ( .A(n1028), .B(n38130), .Z(n38129) );
  XOR U37922 ( .A(n38131), .B(n38128), .Z(n38130) );
  XOR U37923 ( .A(n38132), .B(n38133), .Z(n38120) );
  AND U37924 ( .A(n38134), .B(n38135), .Z(n38133) );
  XOR U37925 ( .A(n38132), .B(n30855), .Z(n38135) );
  XOR U37926 ( .A(n38136), .B(n38137), .Z(n30855) );
  AND U37927 ( .A(n1031), .B(n38138), .Z(n38137) );
  XOR U37928 ( .A(n38139), .B(n38136), .Z(n38138) );
  XNOR U37929 ( .A(n30852), .B(n38132), .Z(n38134) );
  XOR U37930 ( .A(n38140), .B(n38141), .Z(n30852) );
  AND U37931 ( .A(n1028), .B(n38142), .Z(n38141) );
  XOR U37932 ( .A(n38143), .B(n38140), .Z(n38142) );
  XOR U37933 ( .A(n38144), .B(n38145), .Z(n38132) );
  AND U37934 ( .A(n38146), .B(n38147), .Z(n38145) );
  XOR U37935 ( .A(n38144), .B(n30867), .Z(n38147) );
  XOR U37936 ( .A(n38148), .B(n38149), .Z(n30867) );
  AND U37937 ( .A(n1031), .B(n38150), .Z(n38149) );
  XOR U37938 ( .A(n38151), .B(n38148), .Z(n38150) );
  XNOR U37939 ( .A(n30864), .B(n38144), .Z(n38146) );
  XOR U37940 ( .A(n38152), .B(n38153), .Z(n30864) );
  AND U37941 ( .A(n1028), .B(n38154), .Z(n38153) );
  XOR U37942 ( .A(n38155), .B(n38152), .Z(n38154) );
  XOR U37943 ( .A(n38156), .B(n38157), .Z(n38144) );
  AND U37944 ( .A(n38158), .B(n38159), .Z(n38157) );
  XOR U37945 ( .A(n38156), .B(n30879), .Z(n38159) );
  XOR U37946 ( .A(n38160), .B(n38161), .Z(n30879) );
  AND U37947 ( .A(n1031), .B(n38162), .Z(n38161) );
  XOR U37948 ( .A(n38163), .B(n38160), .Z(n38162) );
  XNOR U37949 ( .A(n30876), .B(n38156), .Z(n38158) );
  XOR U37950 ( .A(n38164), .B(n38165), .Z(n30876) );
  AND U37951 ( .A(n1028), .B(n38166), .Z(n38165) );
  XOR U37952 ( .A(n38167), .B(n38164), .Z(n38166) );
  XOR U37953 ( .A(n38168), .B(n38169), .Z(n38156) );
  AND U37954 ( .A(n38170), .B(n38171), .Z(n38169) );
  XOR U37955 ( .A(n38168), .B(n30891), .Z(n38171) );
  XOR U37956 ( .A(n38172), .B(n38173), .Z(n30891) );
  AND U37957 ( .A(n1031), .B(n38174), .Z(n38173) );
  XOR U37958 ( .A(n38175), .B(n38172), .Z(n38174) );
  XNOR U37959 ( .A(n30888), .B(n38168), .Z(n38170) );
  XOR U37960 ( .A(n38176), .B(n38177), .Z(n30888) );
  AND U37961 ( .A(n1028), .B(n38178), .Z(n38177) );
  XOR U37962 ( .A(n38179), .B(n38176), .Z(n38178) );
  XOR U37963 ( .A(n38180), .B(n38181), .Z(n38168) );
  AND U37964 ( .A(n38182), .B(n38183), .Z(n38181) );
  XOR U37965 ( .A(n38180), .B(n30903), .Z(n38183) );
  XOR U37966 ( .A(n38184), .B(n38185), .Z(n30903) );
  AND U37967 ( .A(n1031), .B(n38186), .Z(n38185) );
  XOR U37968 ( .A(n38187), .B(n38184), .Z(n38186) );
  XNOR U37969 ( .A(n30900), .B(n38180), .Z(n38182) );
  XOR U37970 ( .A(n38188), .B(n38189), .Z(n30900) );
  AND U37971 ( .A(n1028), .B(n38190), .Z(n38189) );
  XOR U37972 ( .A(n38191), .B(n38188), .Z(n38190) );
  XOR U37973 ( .A(n38192), .B(n38193), .Z(n38180) );
  AND U37974 ( .A(n38194), .B(n38195), .Z(n38193) );
  XOR U37975 ( .A(n38192), .B(n30915), .Z(n38195) );
  XOR U37976 ( .A(n38196), .B(n38197), .Z(n30915) );
  AND U37977 ( .A(n1031), .B(n38198), .Z(n38197) );
  XOR U37978 ( .A(n38199), .B(n38196), .Z(n38198) );
  XNOR U37979 ( .A(n30912), .B(n38192), .Z(n38194) );
  XOR U37980 ( .A(n38200), .B(n38201), .Z(n30912) );
  AND U37981 ( .A(n1028), .B(n38202), .Z(n38201) );
  XOR U37982 ( .A(n38203), .B(n38200), .Z(n38202) );
  XOR U37983 ( .A(n38204), .B(n38205), .Z(n38192) );
  AND U37984 ( .A(n38206), .B(n38207), .Z(n38205) );
  XOR U37985 ( .A(n38204), .B(n30927), .Z(n38207) );
  XOR U37986 ( .A(n38208), .B(n38209), .Z(n30927) );
  AND U37987 ( .A(n1031), .B(n38210), .Z(n38209) );
  XOR U37988 ( .A(n38211), .B(n38208), .Z(n38210) );
  XNOR U37989 ( .A(n30924), .B(n38204), .Z(n38206) );
  XOR U37990 ( .A(n38212), .B(n38213), .Z(n30924) );
  AND U37991 ( .A(n1028), .B(n38214), .Z(n38213) );
  XOR U37992 ( .A(n38215), .B(n38212), .Z(n38214) );
  XOR U37993 ( .A(n38216), .B(n38217), .Z(n38204) );
  AND U37994 ( .A(n38218), .B(n38219), .Z(n38217) );
  XOR U37995 ( .A(n38216), .B(n30939), .Z(n38219) );
  XOR U37996 ( .A(n38220), .B(n38221), .Z(n30939) );
  AND U37997 ( .A(n1031), .B(n38222), .Z(n38221) );
  XOR U37998 ( .A(n38223), .B(n38220), .Z(n38222) );
  XNOR U37999 ( .A(n30936), .B(n38216), .Z(n38218) );
  XOR U38000 ( .A(n38224), .B(n38225), .Z(n30936) );
  AND U38001 ( .A(n1028), .B(n38226), .Z(n38225) );
  XOR U38002 ( .A(n38227), .B(n38224), .Z(n38226) );
  XOR U38003 ( .A(n38228), .B(n38229), .Z(n38216) );
  AND U38004 ( .A(n38230), .B(n38231), .Z(n38229) );
  XOR U38005 ( .A(n38228), .B(n30951), .Z(n38231) );
  XOR U38006 ( .A(n38232), .B(n38233), .Z(n30951) );
  AND U38007 ( .A(n1031), .B(n38234), .Z(n38233) );
  XOR U38008 ( .A(n38235), .B(n38232), .Z(n38234) );
  XNOR U38009 ( .A(n30948), .B(n38228), .Z(n38230) );
  XOR U38010 ( .A(n38236), .B(n38237), .Z(n30948) );
  AND U38011 ( .A(n1028), .B(n38238), .Z(n38237) );
  XOR U38012 ( .A(n38239), .B(n38236), .Z(n38238) );
  XOR U38013 ( .A(n38240), .B(n38241), .Z(n38228) );
  AND U38014 ( .A(n38242), .B(n38243), .Z(n38241) );
  XOR U38015 ( .A(n38240), .B(n30963), .Z(n38243) );
  XOR U38016 ( .A(n38244), .B(n38245), .Z(n30963) );
  AND U38017 ( .A(n1031), .B(n38246), .Z(n38245) );
  XOR U38018 ( .A(n38247), .B(n38244), .Z(n38246) );
  XNOR U38019 ( .A(n30960), .B(n38240), .Z(n38242) );
  XOR U38020 ( .A(n38248), .B(n38249), .Z(n30960) );
  AND U38021 ( .A(n1028), .B(n38250), .Z(n38249) );
  XOR U38022 ( .A(n38251), .B(n38248), .Z(n38250) );
  XOR U38023 ( .A(n38252), .B(n38253), .Z(n38240) );
  AND U38024 ( .A(n38254), .B(n38255), .Z(n38253) );
  XOR U38025 ( .A(n38252), .B(n30975), .Z(n38255) );
  XOR U38026 ( .A(n38256), .B(n38257), .Z(n30975) );
  AND U38027 ( .A(n1031), .B(n38258), .Z(n38257) );
  XOR U38028 ( .A(n38259), .B(n38256), .Z(n38258) );
  XNOR U38029 ( .A(n30972), .B(n38252), .Z(n38254) );
  XOR U38030 ( .A(n38260), .B(n38261), .Z(n30972) );
  AND U38031 ( .A(n1028), .B(n38262), .Z(n38261) );
  XOR U38032 ( .A(n38263), .B(n38260), .Z(n38262) );
  XOR U38033 ( .A(n38264), .B(n38265), .Z(n38252) );
  AND U38034 ( .A(n38266), .B(n38267), .Z(n38265) );
  XOR U38035 ( .A(n38264), .B(n30987), .Z(n38267) );
  XOR U38036 ( .A(n38268), .B(n38269), .Z(n30987) );
  AND U38037 ( .A(n1031), .B(n38270), .Z(n38269) );
  XOR U38038 ( .A(n38271), .B(n38268), .Z(n38270) );
  XNOR U38039 ( .A(n30984), .B(n38264), .Z(n38266) );
  XOR U38040 ( .A(n38272), .B(n38273), .Z(n30984) );
  AND U38041 ( .A(n1028), .B(n38274), .Z(n38273) );
  XOR U38042 ( .A(n38275), .B(n38272), .Z(n38274) );
  XOR U38043 ( .A(n38276), .B(n38277), .Z(n38264) );
  AND U38044 ( .A(n38278), .B(n38279), .Z(n38277) );
  XOR U38045 ( .A(n38276), .B(n30999), .Z(n38279) );
  XOR U38046 ( .A(n38280), .B(n38281), .Z(n30999) );
  AND U38047 ( .A(n1031), .B(n38282), .Z(n38281) );
  XOR U38048 ( .A(n38283), .B(n38280), .Z(n38282) );
  XNOR U38049 ( .A(n30996), .B(n38276), .Z(n38278) );
  XOR U38050 ( .A(n38284), .B(n38285), .Z(n30996) );
  AND U38051 ( .A(n1028), .B(n38286), .Z(n38285) );
  XOR U38052 ( .A(n38287), .B(n38284), .Z(n38286) );
  XOR U38053 ( .A(n38288), .B(n38289), .Z(n38276) );
  AND U38054 ( .A(n38290), .B(n38291), .Z(n38289) );
  XOR U38055 ( .A(n38288), .B(n31011), .Z(n38291) );
  XOR U38056 ( .A(n38292), .B(n38293), .Z(n31011) );
  AND U38057 ( .A(n1031), .B(n38294), .Z(n38293) );
  XOR U38058 ( .A(n38295), .B(n38292), .Z(n38294) );
  XNOR U38059 ( .A(n31008), .B(n38288), .Z(n38290) );
  XOR U38060 ( .A(n38296), .B(n38297), .Z(n31008) );
  AND U38061 ( .A(n1028), .B(n38298), .Z(n38297) );
  XOR U38062 ( .A(n38299), .B(n38296), .Z(n38298) );
  XOR U38063 ( .A(n38300), .B(n38301), .Z(n38288) );
  AND U38064 ( .A(n38302), .B(n38303), .Z(n38301) );
  XOR U38065 ( .A(n38300), .B(n31023), .Z(n38303) );
  XOR U38066 ( .A(n38304), .B(n38305), .Z(n31023) );
  AND U38067 ( .A(n1031), .B(n38306), .Z(n38305) );
  XOR U38068 ( .A(n38307), .B(n38304), .Z(n38306) );
  XNOR U38069 ( .A(n31020), .B(n38300), .Z(n38302) );
  XOR U38070 ( .A(n38308), .B(n38309), .Z(n31020) );
  AND U38071 ( .A(n1028), .B(n38310), .Z(n38309) );
  XOR U38072 ( .A(n38311), .B(n38308), .Z(n38310) );
  XOR U38073 ( .A(n38312), .B(n38313), .Z(n38300) );
  AND U38074 ( .A(n38314), .B(n38315), .Z(n38313) );
  XOR U38075 ( .A(n38312), .B(n31035), .Z(n38315) );
  XOR U38076 ( .A(n38316), .B(n38317), .Z(n31035) );
  AND U38077 ( .A(n1031), .B(n38318), .Z(n38317) );
  XOR U38078 ( .A(n38319), .B(n38316), .Z(n38318) );
  XNOR U38079 ( .A(n31032), .B(n38312), .Z(n38314) );
  XOR U38080 ( .A(n38320), .B(n38321), .Z(n31032) );
  AND U38081 ( .A(n1028), .B(n38322), .Z(n38321) );
  XOR U38082 ( .A(n38323), .B(n38320), .Z(n38322) );
  XOR U38083 ( .A(n38324), .B(n38325), .Z(n38312) );
  AND U38084 ( .A(n38326), .B(n38327), .Z(n38325) );
  XNOR U38085 ( .A(n38328), .B(n31048), .Z(n38327) );
  XOR U38086 ( .A(n38329), .B(n38330), .Z(n31048) );
  AND U38087 ( .A(n1031), .B(n38331), .Z(n38330) );
  XOR U38088 ( .A(n38329), .B(n38332), .Z(n38331) );
  XNOR U38089 ( .A(n31045), .B(n38324), .Z(n38326) );
  XOR U38090 ( .A(n38333), .B(n38334), .Z(n31045) );
  AND U38091 ( .A(n1028), .B(n38335), .Z(n38334) );
  XOR U38092 ( .A(n38333), .B(n38336), .Z(n38335) );
  IV U38093 ( .A(n38328), .Z(n38324) );
  AND U38094 ( .A(n37960), .B(n37963), .Z(n38328) );
  XNOR U38095 ( .A(n38337), .B(n38338), .Z(n37963) );
  AND U38096 ( .A(n1031), .B(n38339), .Z(n38338) );
  XNOR U38097 ( .A(n38340), .B(n38337), .Z(n38339) );
  XOR U38098 ( .A(n38341), .B(n38342), .Z(n1031) );
  AND U38099 ( .A(n38343), .B(n38344), .Z(n38342) );
  XOR U38100 ( .A(n38341), .B(n37971), .Z(n38344) );
  XOR U38101 ( .A(n38345), .B(n38346), .Z(n37971) );
  AND U38102 ( .A(n887), .B(n38347), .Z(n38346) );
  XOR U38103 ( .A(n38348), .B(n38345), .Z(n38347) );
  XNOR U38104 ( .A(n37968), .B(n38341), .Z(n38343) );
  XOR U38105 ( .A(n38349), .B(n38350), .Z(n37968) );
  AND U38106 ( .A(n885), .B(n38351), .Z(n38350) );
  XOR U38107 ( .A(n38352), .B(n38349), .Z(n38351) );
  XOR U38108 ( .A(n38353), .B(n38354), .Z(n38341) );
  AND U38109 ( .A(n38355), .B(n38356), .Z(n38354) );
  XOR U38110 ( .A(n38353), .B(n37983), .Z(n38356) );
  XOR U38111 ( .A(n38357), .B(n38358), .Z(n37983) );
  AND U38112 ( .A(n887), .B(n38359), .Z(n38358) );
  XOR U38113 ( .A(n38360), .B(n38357), .Z(n38359) );
  XNOR U38114 ( .A(n37980), .B(n38353), .Z(n38355) );
  XOR U38115 ( .A(n38361), .B(n38362), .Z(n37980) );
  AND U38116 ( .A(n885), .B(n38363), .Z(n38362) );
  XOR U38117 ( .A(n38364), .B(n38361), .Z(n38363) );
  XOR U38118 ( .A(n38365), .B(n38366), .Z(n38353) );
  AND U38119 ( .A(n38367), .B(n38368), .Z(n38366) );
  XOR U38120 ( .A(n38365), .B(n37995), .Z(n38368) );
  XOR U38121 ( .A(n38369), .B(n38370), .Z(n37995) );
  AND U38122 ( .A(n887), .B(n38371), .Z(n38370) );
  XOR U38123 ( .A(n38372), .B(n38369), .Z(n38371) );
  XNOR U38124 ( .A(n37992), .B(n38365), .Z(n38367) );
  XOR U38125 ( .A(n38373), .B(n38374), .Z(n37992) );
  AND U38126 ( .A(n885), .B(n38375), .Z(n38374) );
  XOR U38127 ( .A(n38376), .B(n38373), .Z(n38375) );
  XOR U38128 ( .A(n38377), .B(n38378), .Z(n38365) );
  AND U38129 ( .A(n38379), .B(n38380), .Z(n38378) );
  XOR U38130 ( .A(n38377), .B(n38007), .Z(n38380) );
  XOR U38131 ( .A(n38381), .B(n38382), .Z(n38007) );
  AND U38132 ( .A(n887), .B(n38383), .Z(n38382) );
  XOR U38133 ( .A(n38384), .B(n38381), .Z(n38383) );
  XNOR U38134 ( .A(n38004), .B(n38377), .Z(n38379) );
  XOR U38135 ( .A(n38385), .B(n38386), .Z(n38004) );
  AND U38136 ( .A(n885), .B(n38387), .Z(n38386) );
  XOR U38137 ( .A(n38388), .B(n38385), .Z(n38387) );
  XOR U38138 ( .A(n38389), .B(n38390), .Z(n38377) );
  AND U38139 ( .A(n38391), .B(n38392), .Z(n38390) );
  XOR U38140 ( .A(n38389), .B(n38019), .Z(n38392) );
  XOR U38141 ( .A(n38393), .B(n38394), .Z(n38019) );
  AND U38142 ( .A(n887), .B(n38395), .Z(n38394) );
  XOR U38143 ( .A(n38396), .B(n38393), .Z(n38395) );
  XNOR U38144 ( .A(n38016), .B(n38389), .Z(n38391) );
  XOR U38145 ( .A(n38397), .B(n38398), .Z(n38016) );
  AND U38146 ( .A(n885), .B(n38399), .Z(n38398) );
  XOR U38147 ( .A(n38400), .B(n38397), .Z(n38399) );
  XOR U38148 ( .A(n38401), .B(n38402), .Z(n38389) );
  AND U38149 ( .A(n38403), .B(n38404), .Z(n38402) );
  XOR U38150 ( .A(n38401), .B(n38031), .Z(n38404) );
  XOR U38151 ( .A(n38405), .B(n38406), .Z(n38031) );
  AND U38152 ( .A(n887), .B(n38407), .Z(n38406) );
  XOR U38153 ( .A(n38408), .B(n38405), .Z(n38407) );
  XNOR U38154 ( .A(n38028), .B(n38401), .Z(n38403) );
  XOR U38155 ( .A(n38409), .B(n38410), .Z(n38028) );
  AND U38156 ( .A(n885), .B(n38411), .Z(n38410) );
  XOR U38157 ( .A(n38412), .B(n38409), .Z(n38411) );
  XOR U38158 ( .A(n38413), .B(n38414), .Z(n38401) );
  AND U38159 ( .A(n38415), .B(n38416), .Z(n38414) );
  XOR U38160 ( .A(n38413), .B(n38043), .Z(n38416) );
  XOR U38161 ( .A(n38417), .B(n38418), .Z(n38043) );
  AND U38162 ( .A(n887), .B(n38419), .Z(n38418) );
  XOR U38163 ( .A(n38420), .B(n38417), .Z(n38419) );
  XNOR U38164 ( .A(n38040), .B(n38413), .Z(n38415) );
  XOR U38165 ( .A(n38421), .B(n38422), .Z(n38040) );
  AND U38166 ( .A(n885), .B(n38423), .Z(n38422) );
  XOR U38167 ( .A(n38424), .B(n38421), .Z(n38423) );
  XOR U38168 ( .A(n38425), .B(n38426), .Z(n38413) );
  AND U38169 ( .A(n38427), .B(n38428), .Z(n38426) );
  XOR U38170 ( .A(n38425), .B(n38055), .Z(n38428) );
  XOR U38171 ( .A(n38429), .B(n38430), .Z(n38055) );
  AND U38172 ( .A(n887), .B(n38431), .Z(n38430) );
  XOR U38173 ( .A(n38432), .B(n38429), .Z(n38431) );
  XNOR U38174 ( .A(n38052), .B(n38425), .Z(n38427) );
  XOR U38175 ( .A(n38433), .B(n38434), .Z(n38052) );
  AND U38176 ( .A(n885), .B(n38435), .Z(n38434) );
  XOR U38177 ( .A(n38436), .B(n38433), .Z(n38435) );
  XOR U38178 ( .A(n38437), .B(n38438), .Z(n38425) );
  AND U38179 ( .A(n38439), .B(n38440), .Z(n38438) );
  XOR U38180 ( .A(n38437), .B(n38067), .Z(n38440) );
  XOR U38181 ( .A(n38441), .B(n38442), .Z(n38067) );
  AND U38182 ( .A(n887), .B(n38443), .Z(n38442) );
  XOR U38183 ( .A(n38444), .B(n38441), .Z(n38443) );
  XNOR U38184 ( .A(n38064), .B(n38437), .Z(n38439) );
  XOR U38185 ( .A(n38445), .B(n38446), .Z(n38064) );
  AND U38186 ( .A(n885), .B(n38447), .Z(n38446) );
  XOR U38187 ( .A(n38448), .B(n38445), .Z(n38447) );
  XOR U38188 ( .A(n38449), .B(n38450), .Z(n38437) );
  AND U38189 ( .A(n38451), .B(n38452), .Z(n38450) );
  XOR U38190 ( .A(n38449), .B(n38079), .Z(n38452) );
  XOR U38191 ( .A(n38453), .B(n38454), .Z(n38079) );
  AND U38192 ( .A(n887), .B(n38455), .Z(n38454) );
  XOR U38193 ( .A(n38456), .B(n38453), .Z(n38455) );
  XNOR U38194 ( .A(n38076), .B(n38449), .Z(n38451) );
  XOR U38195 ( .A(n38457), .B(n38458), .Z(n38076) );
  AND U38196 ( .A(n885), .B(n38459), .Z(n38458) );
  XOR U38197 ( .A(n38460), .B(n38457), .Z(n38459) );
  XOR U38198 ( .A(n38461), .B(n38462), .Z(n38449) );
  AND U38199 ( .A(n38463), .B(n38464), .Z(n38462) );
  XOR U38200 ( .A(n38461), .B(n38091), .Z(n38464) );
  XOR U38201 ( .A(n38465), .B(n38466), .Z(n38091) );
  AND U38202 ( .A(n887), .B(n38467), .Z(n38466) );
  XOR U38203 ( .A(n38468), .B(n38465), .Z(n38467) );
  XNOR U38204 ( .A(n38088), .B(n38461), .Z(n38463) );
  XOR U38205 ( .A(n38469), .B(n38470), .Z(n38088) );
  AND U38206 ( .A(n885), .B(n38471), .Z(n38470) );
  XOR U38207 ( .A(n38472), .B(n38469), .Z(n38471) );
  XOR U38208 ( .A(n38473), .B(n38474), .Z(n38461) );
  AND U38209 ( .A(n38475), .B(n38476), .Z(n38474) );
  XOR U38210 ( .A(n38473), .B(n38103), .Z(n38476) );
  XOR U38211 ( .A(n38477), .B(n38478), .Z(n38103) );
  AND U38212 ( .A(n887), .B(n38479), .Z(n38478) );
  XOR U38213 ( .A(n38480), .B(n38477), .Z(n38479) );
  XNOR U38214 ( .A(n38100), .B(n38473), .Z(n38475) );
  XOR U38215 ( .A(n38481), .B(n38482), .Z(n38100) );
  AND U38216 ( .A(n885), .B(n38483), .Z(n38482) );
  XOR U38217 ( .A(n38484), .B(n38481), .Z(n38483) );
  XOR U38218 ( .A(n38485), .B(n38486), .Z(n38473) );
  AND U38219 ( .A(n38487), .B(n38488), .Z(n38486) );
  XOR U38220 ( .A(n38485), .B(n38115), .Z(n38488) );
  XOR U38221 ( .A(n38489), .B(n38490), .Z(n38115) );
  AND U38222 ( .A(n887), .B(n38491), .Z(n38490) );
  XOR U38223 ( .A(n38492), .B(n38489), .Z(n38491) );
  XNOR U38224 ( .A(n38112), .B(n38485), .Z(n38487) );
  XOR U38225 ( .A(n38493), .B(n38494), .Z(n38112) );
  AND U38226 ( .A(n885), .B(n38495), .Z(n38494) );
  XOR U38227 ( .A(n38496), .B(n38493), .Z(n38495) );
  XOR U38228 ( .A(n38497), .B(n38498), .Z(n38485) );
  AND U38229 ( .A(n38499), .B(n38500), .Z(n38498) );
  XOR U38230 ( .A(n38497), .B(n38127), .Z(n38500) );
  XOR U38231 ( .A(n38501), .B(n38502), .Z(n38127) );
  AND U38232 ( .A(n887), .B(n38503), .Z(n38502) );
  XOR U38233 ( .A(n38504), .B(n38501), .Z(n38503) );
  XNOR U38234 ( .A(n38124), .B(n38497), .Z(n38499) );
  XOR U38235 ( .A(n38505), .B(n38506), .Z(n38124) );
  AND U38236 ( .A(n885), .B(n38507), .Z(n38506) );
  XOR U38237 ( .A(n38508), .B(n38505), .Z(n38507) );
  XOR U38238 ( .A(n38509), .B(n38510), .Z(n38497) );
  AND U38239 ( .A(n38511), .B(n38512), .Z(n38510) );
  XOR U38240 ( .A(n38509), .B(n38139), .Z(n38512) );
  XOR U38241 ( .A(n38513), .B(n38514), .Z(n38139) );
  AND U38242 ( .A(n887), .B(n38515), .Z(n38514) );
  XOR U38243 ( .A(n38516), .B(n38513), .Z(n38515) );
  XNOR U38244 ( .A(n38136), .B(n38509), .Z(n38511) );
  XOR U38245 ( .A(n38517), .B(n38518), .Z(n38136) );
  AND U38246 ( .A(n885), .B(n38519), .Z(n38518) );
  XOR U38247 ( .A(n38520), .B(n38517), .Z(n38519) );
  XOR U38248 ( .A(n38521), .B(n38522), .Z(n38509) );
  AND U38249 ( .A(n38523), .B(n38524), .Z(n38522) );
  XOR U38250 ( .A(n38521), .B(n38151), .Z(n38524) );
  XOR U38251 ( .A(n38525), .B(n38526), .Z(n38151) );
  AND U38252 ( .A(n887), .B(n38527), .Z(n38526) );
  XOR U38253 ( .A(n38528), .B(n38525), .Z(n38527) );
  XNOR U38254 ( .A(n38148), .B(n38521), .Z(n38523) );
  XOR U38255 ( .A(n38529), .B(n38530), .Z(n38148) );
  AND U38256 ( .A(n885), .B(n38531), .Z(n38530) );
  XOR U38257 ( .A(n38532), .B(n38529), .Z(n38531) );
  XOR U38258 ( .A(n38533), .B(n38534), .Z(n38521) );
  AND U38259 ( .A(n38535), .B(n38536), .Z(n38534) );
  XOR U38260 ( .A(n38533), .B(n38163), .Z(n38536) );
  XOR U38261 ( .A(n38537), .B(n38538), .Z(n38163) );
  AND U38262 ( .A(n887), .B(n38539), .Z(n38538) );
  XOR U38263 ( .A(n38540), .B(n38537), .Z(n38539) );
  XNOR U38264 ( .A(n38160), .B(n38533), .Z(n38535) );
  XOR U38265 ( .A(n38541), .B(n38542), .Z(n38160) );
  AND U38266 ( .A(n885), .B(n38543), .Z(n38542) );
  XOR U38267 ( .A(n38544), .B(n38541), .Z(n38543) );
  XOR U38268 ( .A(n38545), .B(n38546), .Z(n38533) );
  AND U38269 ( .A(n38547), .B(n38548), .Z(n38546) );
  XOR U38270 ( .A(n38545), .B(n38175), .Z(n38548) );
  XOR U38271 ( .A(n38549), .B(n38550), .Z(n38175) );
  AND U38272 ( .A(n887), .B(n38551), .Z(n38550) );
  XOR U38273 ( .A(n38552), .B(n38549), .Z(n38551) );
  XNOR U38274 ( .A(n38172), .B(n38545), .Z(n38547) );
  XOR U38275 ( .A(n38553), .B(n38554), .Z(n38172) );
  AND U38276 ( .A(n885), .B(n38555), .Z(n38554) );
  XOR U38277 ( .A(n38556), .B(n38553), .Z(n38555) );
  XOR U38278 ( .A(n38557), .B(n38558), .Z(n38545) );
  AND U38279 ( .A(n38559), .B(n38560), .Z(n38558) );
  XOR U38280 ( .A(n38557), .B(n38187), .Z(n38560) );
  XOR U38281 ( .A(n38561), .B(n38562), .Z(n38187) );
  AND U38282 ( .A(n887), .B(n38563), .Z(n38562) );
  XOR U38283 ( .A(n38564), .B(n38561), .Z(n38563) );
  XNOR U38284 ( .A(n38184), .B(n38557), .Z(n38559) );
  XOR U38285 ( .A(n38565), .B(n38566), .Z(n38184) );
  AND U38286 ( .A(n885), .B(n38567), .Z(n38566) );
  XOR U38287 ( .A(n38568), .B(n38565), .Z(n38567) );
  XOR U38288 ( .A(n38569), .B(n38570), .Z(n38557) );
  AND U38289 ( .A(n38571), .B(n38572), .Z(n38570) );
  XOR U38290 ( .A(n38569), .B(n38199), .Z(n38572) );
  XOR U38291 ( .A(n38573), .B(n38574), .Z(n38199) );
  AND U38292 ( .A(n887), .B(n38575), .Z(n38574) );
  XOR U38293 ( .A(n38576), .B(n38573), .Z(n38575) );
  XNOR U38294 ( .A(n38196), .B(n38569), .Z(n38571) );
  XOR U38295 ( .A(n38577), .B(n38578), .Z(n38196) );
  AND U38296 ( .A(n885), .B(n38579), .Z(n38578) );
  XOR U38297 ( .A(n38580), .B(n38577), .Z(n38579) );
  XOR U38298 ( .A(n38581), .B(n38582), .Z(n38569) );
  AND U38299 ( .A(n38583), .B(n38584), .Z(n38582) );
  XOR U38300 ( .A(n38581), .B(n38211), .Z(n38584) );
  XOR U38301 ( .A(n38585), .B(n38586), .Z(n38211) );
  AND U38302 ( .A(n887), .B(n38587), .Z(n38586) );
  XOR U38303 ( .A(n38588), .B(n38585), .Z(n38587) );
  XNOR U38304 ( .A(n38208), .B(n38581), .Z(n38583) );
  XOR U38305 ( .A(n38589), .B(n38590), .Z(n38208) );
  AND U38306 ( .A(n885), .B(n38591), .Z(n38590) );
  XOR U38307 ( .A(n38592), .B(n38589), .Z(n38591) );
  XOR U38308 ( .A(n38593), .B(n38594), .Z(n38581) );
  AND U38309 ( .A(n38595), .B(n38596), .Z(n38594) );
  XOR U38310 ( .A(n38593), .B(n38223), .Z(n38596) );
  XOR U38311 ( .A(n38597), .B(n38598), .Z(n38223) );
  AND U38312 ( .A(n887), .B(n38599), .Z(n38598) );
  XOR U38313 ( .A(n38600), .B(n38597), .Z(n38599) );
  XNOR U38314 ( .A(n38220), .B(n38593), .Z(n38595) );
  XOR U38315 ( .A(n38601), .B(n38602), .Z(n38220) );
  AND U38316 ( .A(n885), .B(n38603), .Z(n38602) );
  XOR U38317 ( .A(n38604), .B(n38601), .Z(n38603) );
  XOR U38318 ( .A(n38605), .B(n38606), .Z(n38593) );
  AND U38319 ( .A(n38607), .B(n38608), .Z(n38606) );
  XOR U38320 ( .A(n38605), .B(n38235), .Z(n38608) );
  XOR U38321 ( .A(n38609), .B(n38610), .Z(n38235) );
  AND U38322 ( .A(n887), .B(n38611), .Z(n38610) );
  XOR U38323 ( .A(n38612), .B(n38609), .Z(n38611) );
  XNOR U38324 ( .A(n38232), .B(n38605), .Z(n38607) );
  XOR U38325 ( .A(n38613), .B(n38614), .Z(n38232) );
  AND U38326 ( .A(n885), .B(n38615), .Z(n38614) );
  XOR U38327 ( .A(n38616), .B(n38613), .Z(n38615) );
  XOR U38328 ( .A(n38617), .B(n38618), .Z(n38605) );
  AND U38329 ( .A(n38619), .B(n38620), .Z(n38618) );
  XOR U38330 ( .A(n38617), .B(n38247), .Z(n38620) );
  XOR U38331 ( .A(n38621), .B(n38622), .Z(n38247) );
  AND U38332 ( .A(n887), .B(n38623), .Z(n38622) );
  XOR U38333 ( .A(n38624), .B(n38621), .Z(n38623) );
  XNOR U38334 ( .A(n38244), .B(n38617), .Z(n38619) );
  XOR U38335 ( .A(n38625), .B(n38626), .Z(n38244) );
  AND U38336 ( .A(n885), .B(n38627), .Z(n38626) );
  XOR U38337 ( .A(n38628), .B(n38625), .Z(n38627) );
  XOR U38338 ( .A(n38629), .B(n38630), .Z(n38617) );
  AND U38339 ( .A(n38631), .B(n38632), .Z(n38630) );
  XOR U38340 ( .A(n38629), .B(n38259), .Z(n38632) );
  XOR U38341 ( .A(n38633), .B(n38634), .Z(n38259) );
  AND U38342 ( .A(n887), .B(n38635), .Z(n38634) );
  XOR U38343 ( .A(n38636), .B(n38633), .Z(n38635) );
  XNOR U38344 ( .A(n38256), .B(n38629), .Z(n38631) );
  XOR U38345 ( .A(n38637), .B(n38638), .Z(n38256) );
  AND U38346 ( .A(n885), .B(n38639), .Z(n38638) );
  XOR U38347 ( .A(n38640), .B(n38637), .Z(n38639) );
  XOR U38348 ( .A(n38641), .B(n38642), .Z(n38629) );
  AND U38349 ( .A(n38643), .B(n38644), .Z(n38642) );
  XOR U38350 ( .A(n38641), .B(n38271), .Z(n38644) );
  XOR U38351 ( .A(n38645), .B(n38646), .Z(n38271) );
  AND U38352 ( .A(n887), .B(n38647), .Z(n38646) );
  XOR U38353 ( .A(n38648), .B(n38645), .Z(n38647) );
  XNOR U38354 ( .A(n38268), .B(n38641), .Z(n38643) );
  XOR U38355 ( .A(n38649), .B(n38650), .Z(n38268) );
  AND U38356 ( .A(n885), .B(n38651), .Z(n38650) );
  XOR U38357 ( .A(n38652), .B(n38649), .Z(n38651) );
  XOR U38358 ( .A(n38653), .B(n38654), .Z(n38641) );
  AND U38359 ( .A(n38655), .B(n38656), .Z(n38654) );
  XOR U38360 ( .A(n38653), .B(n38283), .Z(n38656) );
  XOR U38361 ( .A(n38657), .B(n38658), .Z(n38283) );
  AND U38362 ( .A(n887), .B(n38659), .Z(n38658) );
  XOR U38363 ( .A(n38660), .B(n38657), .Z(n38659) );
  XNOR U38364 ( .A(n38280), .B(n38653), .Z(n38655) );
  XOR U38365 ( .A(n38661), .B(n38662), .Z(n38280) );
  AND U38366 ( .A(n885), .B(n38663), .Z(n38662) );
  XOR U38367 ( .A(n38664), .B(n38661), .Z(n38663) );
  XOR U38368 ( .A(n38665), .B(n38666), .Z(n38653) );
  AND U38369 ( .A(n38667), .B(n38668), .Z(n38666) );
  XOR U38370 ( .A(n38665), .B(n38295), .Z(n38668) );
  XOR U38371 ( .A(n38669), .B(n38670), .Z(n38295) );
  AND U38372 ( .A(n887), .B(n38671), .Z(n38670) );
  XOR U38373 ( .A(n38672), .B(n38669), .Z(n38671) );
  XNOR U38374 ( .A(n38292), .B(n38665), .Z(n38667) );
  XOR U38375 ( .A(n38673), .B(n38674), .Z(n38292) );
  AND U38376 ( .A(n885), .B(n38675), .Z(n38674) );
  XOR U38377 ( .A(n38676), .B(n38673), .Z(n38675) );
  XOR U38378 ( .A(n38677), .B(n38678), .Z(n38665) );
  AND U38379 ( .A(n38679), .B(n38680), .Z(n38678) );
  XOR U38380 ( .A(n38677), .B(n38307), .Z(n38680) );
  XOR U38381 ( .A(n38681), .B(n38682), .Z(n38307) );
  AND U38382 ( .A(n887), .B(n38683), .Z(n38682) );
  XOR U38383 ( .A(n38684), .B(n38681), .Z(n38683) );
  XNOR U38384 ( .A(n38304), .B(n38677), .Z(n38679) );
  XOR U38385 ( .A(n38685), .B(n38686), .Z(n38304) );
  AND U38386 ( .A(n885), .B(n38687), .Z(n38686) );
  XOR U38387 ( .A(n38688), .B(n38685), .Z(n38687) );
  XOR U38388 ( .A(n38689), .B(n38690), .Z(n38677) );
  AND U38389 ( .A(n38691), .B(n38692), .Z(n38690) );
  XOR U38390 ( .A(n38689), .B(n38319), .Z(n38692) );
  XOR U38391 ( .A(n38693), .B(n38694), .Z(n38319) );
  AND U38392 ( .A(n887), .B(n38695), .Z(n38694) );
  XOR U38393 ( .A(n38696), .B(n38693), .Z(n38695) );
  XNOR U38394 ( .A(n38316), .B(n38689), .Z(n38691) );
  XOR U38395 ( .A(n38697), .B(n38698), .Z(n38316) );
  AND U38396 ( .A(n885), .B(n38699), .Z(n38698) );
  XOR U38397 ( .A(n38700), .B(n38697), .Z(n38699) );
  XOR U38398 ( .A(n38701), .B(n38702), .Z(n38689) );
  AND U38399 ( .A(n38703), .B(n38704), .Z(n38702) );
  XNOR U38400 ( .A(n38705), .B(n38332), .Z(n38704) );
  XOR U38401 ( .A(n38706), .B(n38707), .Z(n38332) );
  AND U38402 ( .A(n887), .B(n38708), .Z(n38707) );
  XOR U38403 ( .A(n38706), .B(n38709), .Z(n38708) );
  XNOR U38404 ( .A(n38329), .B(n38701), .Z(n38703) );
  XOR U38405 ( .A(n38710), .B(n38711), .Z(n38329) );
  AND U38406 ( .A(n885), .B(n38712), .Z(n38711) );
  XOR U38407 ( .A(n38710), .B(n38713), .Z(n38712) );
  IV U38408 ( .A(n38705), .Z(n38701) );
  AND U38409 ( .A(n38337), .B(n38340), .Z(n38705) );
  XNOR U38410 ( .A(n38714), .B(n38715), .Z(n38340) );
  AND U38411 ( .A(n887), .B(n38716), .Z(n38715) );
  XNOR U38412 ( .A(n38717), .B(n38714), .Z(n38716) );
  XOR U38413 ( .A(n38718), .B(n38719), .Z(n887) );
  AND U38414 ( .A(n38720), .B(n38721), .Z(n38719) );
  XOR U38415 ( .A(n38718), .B(n38348), .Z(n38721) );
  XNOR U38416 ( .A(n38722), .B(n38723), .Z(n38348) );
  AND U38417 ( .A(n38724), .B(n591), .Z(n38723) );
  AND U38418 ( .A(n38722), .B(n38725), .Z(n38724) );
  XNOR U38419 ( .A(n38345), .B(n38718), .Z(n38720) );
  XOR U38420 ( .A(n38726), .B(n38727), .Z(n38345) );
  AND U38421 ( .A(n38728), .B(n589), .Z(n38727) );
  NOR U38422 ( .A(n38726), .B(n38729), .Z(n38728) );
  XOR U38423 ( .A(n38730), .B(n38731), .Z(n38718) );
  AND U38424 ( .A(n38732), .B(n38733), .Z(n38731) );
  XOR U38425 ( .A(n38730), .B(n38360), .Z(n38733) );
  XOR U38426 ( .A(n38734), .B(n38735), .Z(n38360) );
  AND U38427 ( .A(n591), .B(n38736), .Z(n38735) );
  XOR U38428 ( .A(n38737), .B(n38734), .Z(n38736) );
  XNOR U38429 ( .A(n38357), .B(n38730), .Z(n38732) );
  XOR U38430 ( .A(n38738), .B(n38739), .Z(n38357) );
  AND U38431 ( .A(n589), .B(n38740), .Z(n38739) );
  XOR U38432 ( .A(n38741), .B(n38738), .Z(n38740) );
  XOR U38433 ( .A(n38742), .B(n38743), .Z(n38730) );
  AND U38434 ( .A(n38744), .B(n38745), .Z(n38743) );
  XOR U38435 ( .A(n38742), .B(n38372), .Z(n38745) );
  XOR U38436 ( .A(n38746), .B(n38747), .Z(n38372) );
  AND U38437 ( .A(n591), .B(n38748), .Z(n38747) );
  XOR U38438 ( .A(n38749), .B(n38746), .Z(n38748) );
  XNOR U38439 ( .A(n38369), .B(n38742), .Z(n38744) );
  XOR U38440 ( .A(n38750), .B(n38751), .Z(n38369) );
  AND U38441 ( .A(n589), .B(n38752), .Z(n38751) );
  XOR U38442 ( .A(n38753), .B(n38750), .Z(n38752) );
  XOR U38443 ( .A(n38754), .B(n38755), .Z(n38742) );
  AND U38444 ( .A(n38756), .B(n38757), .Z(n38755) );
  XOR U38445 ( .A(n38754), .B(n38384), .Z(n38757) );
  XOR U38446 ( .A(n38758), .B(n38759), .Z(n38384) );
  AND U38447 ( .A(n591), .B(n38760), .Z(n38759) );
  XOR U38448 ( .A(n38761), .B(n38758), .Z(n38760) );
  XNOR U38449 ( .A(n38381), .B(n38754), .Z(n38756) );
  XOR U38450 ( .A(n38762), .B(n38763), .Z(n38381) );
  AND U38451 ( .A(n589), .B(n38764), .Z(n38763) );
  XOR U38452 ( .A(n38765), .B(n38762), .Z(n38764) );
  XOR U38453 ( .A(n38766), .B(n38767), .Z(n38754) );
  AND U38454 ( .A(n38768), .B(n38769), .Z(n38767) );
  XOR U38455 ( .A(n38766), .B(n38396), .Z(n38769) );
  XOR U38456 ( .A(n38770), .B(n38771), .Z(n38396) );
  AND U38457 ( .A(n591), .B(n38772), .Z(n38771) );
  XOR U38458 ( .A(n38773), .B(n38770), .Z(n38772) );
  XNOR U38459 ( .A(n38393), .B(n38766), .Z(n38768) );
  XOR U38460 ( .A(n38774), .B(n38775), .Z(n38393) );
  AND U38461 ( .A(n589), .B(n38776), .Z(n38775) );
  XOR U38462 ( .A(n38777), .B(n38774), .Z(n38776) );
  XOR U38463 ( .A(n38778), .B(n38779), .Z(n38766) );
  AND U38464 ( .A(n38780), .B(n38781), .Z(n38779) );
  XOR U38465 ( .A(n38778), .B(n38408), .Z(n38781) );
  XOR U38466 ( .A(n38782), .B(n38783), .Z(n38408) );
  AND U38467 ( .A(n591), .B(n38784), .Z(n38783) );
  XOR U38468 ( .A(n38785), .B(n38782), .Z(n38784) );
  XNOR U38469 ( .A(n38405), .B(n38778), .Z(n38780) );
  XOR U38470 ( .A(n38786), .B(n38787), .Z(n38405) );
  AND U38471 ( .A(n589), .B(n38788), .Z(n38787) );
  XOR U38472 ( .A(n38789), .B(n38786), .Z(n38788) );
  XOR U38473 ( .A(n38790), .B(n38791), .Z(n38778) );
  AND U38474 ( .A(n38792), .B(n38793), .Z(n38791) );
  XOR U38475 ( .A(n38790), .B(n38420), .Z(n38793) );
  XOR U38476 ( .A(n38794), .B(n38795), .Z(n38420) );
  AND U38477 ( .A(n591), .B(n38796), .Z(n38795) );
  XOR U38478 ( .A(n38797), .B(n38794), .Z(n38796) );
  XNOR U38479 ( .A(n38417), .B(n38790), .Z(n38792) );
  XOR U38480 ( .A(n38798), .B(n38799), .Z(n38417) );
  AND U38481 ( .A(n589), .B(n38800), .Z(n38799) );
  XOR U38482 ( .A(n38801), .B(n38798), .Z(n38800) );
  XOR U38483 ( .A(n38802), .B(n38803), .Z(n38790) );
  AND U38484 ( .A(n38804), .B(n38805), .Z(n38803) );
  XOR U38485 ( .A(n38802), .B(n38432), .Z(n38805) );
  XOR U38486 ( .A(n38806), .B(n38807), .Z(n38432) );
  AND U38487 ( .A(n591), .B(n38808), .Z(n38807) );
  XOR U38488 ( .A(n38809), .B(n38806), .Z(n38808) );
  XNOR U38489 ( .A(n38429), .B(n38802), .Z(n38804) );
  XOR U38490 ( .A(n38810), .B(n38811), .Z(n38429) );
  AND U38491 ( .A(n589), .B(n38812), .Z(n38811) );
  XOR U38492 ( .A(n38813), .B(n38810), .Z(n38812) );
  XOR U38493 ( .A(n38814), .B(n38815), .Z(n38802) );
  AND U38494 ( .A(n38816), .B(n38817), .Z(n38815) );
  XOR U38495 ( .A(n38814), .B(n38444), .Z(n38817) );
  XOR U38496 ( .A(n38818), .B(n38819), .Z(n38444) );
  AND U38497 ( .A(n591), .B(n38820), .Z(n38819) );
  XOR U38498 ( .A(n38821), .B(n38818), .Z(n38820) );
  XNOR U38499 ( .A(n38441), .B(n38814), .Z(n38816) );
  XOR U38500 ( .A(n38822), .B(n38823), .Z(n38441) );
  AND U38501 ( .A(n589), .B(n38824), .Z(n38823) );
  XOR U38502 ( .A(n38825), .B(n38822), .Z(n38824) );
  XOR U38503 ( .A(n38826), .B(n38827), .Z(n38814) );
  AND U38504 ( .A(n38828), .B(n38829), .Z(n38827) );
  XOR U38505 ( .A(n38826), .B(n38456), .Z(n38829) );
  XOR U38506 ( .A(n38830), .B(n38831), .Z(n38456) );
  AND U38507 ( .A(n591), .B(n38832), .Z(n38831) );
  XOR U38508 ( .A(n38833), .B(n38830), .Z(n38832) );
  XNOR U38509 ( .A(n38453), .B(n38826), .Z(n38828) );
  XOR U38510 ( .A(n38834), .B(n38835), .Z(n38453) );
  AND U38511 ( .A(n589), .B(n38836), .Z(n38835) );
  XOR U38512 ( .A(n38837), .B(n38834), .Z(n38836) );
  XOR U38513 ( .A(n38838), .B(n38839), .Z(n38826) );
  AND U38514 ( .A(n38840), .B(n38841), .Z(n38839) );
  XOR U38515 ( .A(n38838), .B(n38468), .Z(n38841) );
  XOR U38516 ( .A(n38842), .B(n38843), .Z(n38468) );
  AND U38517 ( .A(n591), .B(n38844), .Z(n38843) );
  XOR U38518 ( .A(n38845), .B(n38842), .Z(n38844) );
  XNOR U38519 ( .A(n38465), .B(n38838), .Z(n38840) );
  XOR U38520 ( .A(n38846), .B(n38847), .Z(n38465) );
  AND U38521 ( .A(n589), .B(n38848), .Z(n38847) );
  XOR U38522 ( .A(n38849), .B(n38846), .Z(n38848) );
  XOR U38523 ( .A(n38850), .B(n38851), .Z(n38838) );
  AND U38524 ( .A(n38852), .B(n38853), .Z(n38851) );
  XOR U38525 ( .A(n38850), .B(n38480), .Z(n38853) );
  XOR U38526 ( .A(n38854), .B(n38855), .Z(n38480) );
  AND U38527 ( .A(n591), .B(n38856), .Z(n38855) );
  XOR U38528 ( .A(n38857), .B(n38854), .Z(n38856) );
  XNOR U38529 ( .A(n38477), .B(n38850), .Z(n38852) );
  XOR U38530 ( .A(n38858), .B(n38859), .Z(n38477) );
  AND U38531 ( .A(n589), .B(n38860), .Z(n38859) );
  XOR U38532 ( .A(n38861), .B(n38858), .Z(n38860) );
  XOR U38533 ( .A(n38862), .B(n38863), .Z(n38850) );
  AND U38534 ( .A(n38864), .B(n38865), .Z(n38863) );
  XOR U38535 ( .A(n38862), .B(n38492), .Z(n38865) );
  XOR U38536 ( .A(n38866), .B(n38867), .Z(n38492) );
  AND U38537 ( .A(n591), .B(n38868), .Z(n38867) );
  XOR U38538 ( .A(n38869), .B(n38866), .Z(n38868) );
  XNOR U38539 ( .A(n38489), .B(n38862), .Z(n38864) );
  XOR U38540 ( .A(n38870), .B(n38871), .Z(n38489) );
  AND U38541 ( .A(n589), .B(n38872), .Z(n38871) );
  XOR U38542 ( .A(n38873), .B(n38870), .Z(n38872) );
  XOR U38543 ( .A(n38874), .B(n38875), .Z(n38862) );
  AND U38544 ( .A(n38876), .B(n38877), .Z(n38875) );
  XOR U38545 ( .A(n38874), .B(n38504), .Z(n38877) );
  XOR U38546 ( .A(n38878), .B(n38879), .Z(n38504) );
  AND U38547 ( .A(n591), .B(n38880), .Z(n38879) );
  XOR U38548 ( .A(n38881), .B(n38878), .Z(n38880) );
  XNOR U38549 ( .A(n38501), .B(n38874), .Z(n38876) );
  XOR U38550 ( .A(n38882), .B(n38883), .Z(n38501) );
  AND U38551 ( .A(n589), .B(n38884), .Z(n38883) );
  XOR U38552 ( .A(n38885), .B(n38882), .Z(n38884) );
  XOR U38553 ( .A(n38886), .B(n38887), .Z(n38874) );
  AND U38554 ( .A(n38888), .B(n38889), .Z(n38887) );
  XOR U38555 ( .A(n38886), .B(n38516), .Z(n38889) );
  XOR U38556 ( .A(n38890), .B(n38891), .Z(n38516) );
  AND U38557 ( .A(n591), .B(n38892), .Z(n38891) );
  XOR U38558 ( .A(n38893), .B(n38890), .Z(n38892) );
  XNOR U38559 ( .A(n38513), .B(n38886), .Z(n38888) );
  XOR U38560 ( .A(n38894), .B(n38895), .Z(n38513) );
  AND U38561 ( .A(n589), .B(n38896), .Z(n38895) );
  XOR U38562 ( .A(n38897), .B(n38894), .Z(n38896) );
  XOR U38563 ( .A(n38898), .B(n38899), .Z(n38886) );
  AND U38564 ( .A(n38900), .B(n38901), .Z(n38899) );
  XOR U38565 ( .A(n38898), .B(n38528), .Z(n38901) );
  XOR U38566 ( .A(n38902), .B(n38903), .Z(n38528) );
  AND U38567 ( .A(n591), .B(n38904), .Z(n38903) );
  XOR U38568 ( .A(n38905), .B(n38902), .Z(n38904) );
  XNOR U38569 ( .A(n38525), .B(n38898), .Z(n38900) );
  XOR U38570 ( .A(n38906), .B(n38907), .Z(n38525) );
  AND U38571 ( .A(n589), .B(n38908), .Z(n38907) );
  XOR U38572 ( .A(n38909), .B(n38906), .Z(n38908) );
  XOR U38573 ( .A(n38910), .B(n38911), .Z(n38898) );
  AND U38574 ( .A(n38912), .B(n38913), .Z(n38911) );
  XOR U38575 ( .A(n38910), .B(n38540), .Z(n38913) );
  XOR U38576 ( .A(n38914), .B(n38915), .Z(n38540) );
  AND U38577 ( .A(n591), .B(n38916), .Z(n38915) );
  XOR U38578 ( .A(n38917), .B(n38914), .Z(n38916) );
  XNOR U38579 ( .A(n38537), .B(n38910), .Z(n38912) );
  XOR U38580 ( .A(n38918), .B(n38919), .Z(n38537) );
  AND U38581 ( .A(n589), .B(n38920), .Z(n38919) );
  XOR U38582 ( .A(n38921), .B(n38918), .Z(n38920) );
  XOR U38583 ( .A(n38922), .B(n38923), .Z(n38910) );
  AND U38584 ( .A(n38924), .B(n38925), .Z(n38923) );
  XOR U38585 ( .A(n38922), .B(n38552), .Z(n38925) );
  XOR U38586 ( .A(n38926), .B(n38927), .Z(n38552) );
  AND U38587 ( .A(n591), .B(n38928), .Z(n38927) );
  XOR U38588 ( .A(n38929), .B(n38926), .Z(n38928) );
  XNOR U38589 ( .A(n38549), .B(n38922), .Z(n38924) );
  XOR U38590 ( .A(n38930), .B(n38931), .Z(n38549) );
  AND U38591 ( .A(n589), .B(n38932), .Z(n38931) );
  XOR U38592 ( .A(n38933), .B(n38930), .Z(n38932) );
  XOR U38593 ( .A(n38934), .B(n38935), .Z(n38922) );
  AND U38594 ( .A(n38936), .B(n38937), .Z(n38935) );
  XOR U38595 ( .A(n38934), .B(n38564), .Z(n38937) );
  XOR U38596 ( .A(n38938), .B(n38939), .Z(n38564) );
  AND U38597 ( .A(n591), .B(n38940), .Z(n38939) );
  XOR U38598 ( .A(n38941), .B(n38938), .Z(n38940) );
  XNOR U38599 ( .A(n38561), .B(n38934), .Z(n38936) );
  XOR U38600 ( .A(n38942), .B(n38943), .Z(n38561) );
  AND U38601 ( .A(n589), .B(n38944), .Z(n38943) );
  XOR U38602 ( .A(n38945), .B(n38942), .Z(n38944) );
  XOR U38603 ( .A(n38946), .B(n38947), .Z(n38934) );
  AND U38604 ( .A(n38948), .B(n38949), .Z(n38947) );
  XOR U38605 ( .A(n38946), .B(n38576), .Z(n38949) );
  XOR U38606 ( .A(n38950), .B(n38951), .Z(n38576) );
  AND U38607 ( .A(n591), .B(n38952), .Z(n38951) );
  XOR U38608 ( .A(n38953), .B(n38950), .Z(n38952) );
  XNOR U38609 ( .A(n38573), .B(n38946), .Z(n38948) );
  XOR U38610 ( .A(n38954), .B(n38955), .Z(n38573) );
  AND U38611 ( .A(n589), .B(n38956), .Z(n38955) );
  XOR U38612 ( .A(n38957), .B(n38954), .Z(n38956) );
  XOR U38613 ( .A(n38958), .B(n38959), .Z(n38946) );
  AND U38614 ( .A(n38960), .B(n38961), .Z(n38959) );
  XOR U38615 ( .A(n38958), .B(n38588), .Z(n38961) );
  XOR U38616 ( .A(n38962), .B(n38963), .Z(n38588) );
  AND U38617 ( .A(n591), .B(n38964), .Z(n38963) );
  XOR U38618 ( .A(n38965), .B(n38962), .Z(n38964) );
  XNOR U38619 ( .A(n38585), .B(n38958), .Z(n38960) );
  XOR U38620 ( .A(n38966), .B(n38967), .Z(n38585) );
  AND U38621 ( .A(n589), .B(n38968), .Z(n38967) );
  XOR U38622 ( .A(n38969), .B(n38966), .Z(n38968) );
  XOR U38623 ( .A(n38970), .B(n38971), .Z(n38958) );
  AND U38624 ( .A(n38972), .B(n38973), .Z(n38971) );
  XOR U38625 ( .A(n38970), .B(n38600), .Z(n38973) );
  XOR U38626 ( .A(n38974), .B(n38975), .Z(n38600) );
  AND U38627 ( .A(n591), .B(n38976), .Z(n38975) );
  XOR U38628 ( .A(n38977), .B(n38974), .Z(n38976) );
  XNOR U38629 ( .A(n38597), .B(n38970), .Z(n38972) );
  XOR U38630 ( .A(n38978), .B(n38979), .Z(n38597) );
  AND U38631 ( .A(n589), .B(n38980), .Z(n38979) );
  XOR U38632 ( .A(n38981), .B(n38978), .Z(n38980) );
  XOR U38633 ( .A(n38982), .B(n38983), .Z(n38970) );
  AND U38634 ( .A(n38984), .B(n38985), .Z(n38983) );
  XOR U38635 ( .A(n38982), .B(n38612), .Z(n38985) );
  XOR U38636 ( .A(n38986), .B(n38987), .Z(n38612) );
  AND U38637 ( .A(n591), .B(n38988), .Z(n38987) );
  XOR U38638 ( .A(n38989), .B(n38986), .Z(n38988) );
  XNOR U38639 ( .A(n38609), .B(n38982), .Z(n38984) );
  XOR U38640 ( .A(n38990), .B(n38991), .Z(n38609) );
  AND U38641 ( .A(n589), .B(n38992), .Z(n38991) );
  XOR U38642 ( .A(n38993), .B(n38990), .Z(n38992) );
  XOR U38643 ( .A(n38994), .B(n38995), .Z(n38982) );
  AND U38644 ( .A(n38996), .B(n38997), .Z(n38995) );
  XOR U38645 ( .A(n38994), .B(n38624), .Z(n38997) );
  XOR U38646 ( .A(n38998), .B(n38999), .Z(n38624) );
  AND U38647 ( .A(n591), .B(n39000), .Z(n38999) );
  XOR U38648 ( .A(n39001), .B(n38998), .Z(n39000) );
  XNOR U38649 ( .A(n38621), .B(n38994), .Z(n38996) );
  XOR U38650 ( .A(n39002), .B(n39003), .Z(n38621) );
  AND U38651 ( .A(n589), .B(n39004), .Z(n39003) );
  XOR U38652 ( .A(n39005), .B(n39002), .Z(n39004) );
  XOR U38653 ( .A(n39006), .B(n39007), .Z(n38994) );
  AND U38654 ( .A(n39008), .B(n39009), .Z(n39007) );
  XOR U38655 ( .A(n39006), .B(n38636), .Z(n39009) );
  XOR U38656 ( .A(n39010), .B(n39011), .Z(n38636) );
  AND U38657 ( .A(n591), .B(n39012), .Z(n39011) );
  XOR U38658 ( .A(n39013), .B(n39010), .Z(n39012) );
  XNOR U38659 ( .A(n38633), .B(n39006), .Z(n39008) );
  XOR U38660 ( .A(n39014), .B(n39015), .Z(n38633) );
  AND U38661 ( .A(n589), .B(n39016), .Z(n39015) );
  XOR U38662 ( .A(n39017), .B(n39014), .Z(n39016) );
  XOR U38663 ( .A(n39018), .B(n39019), .Z(n39006) );
  AND U38664 ( .A(n39020), .B(n39021), .Z(n39019) );
  XOR U38665 ( .A(n39018), .B(n38648), .Z(n39021) );
  XOR U38666 ( .A(n39022), .B(n39023), .Z(n38648) );
  AND U38667 ( .A(n591), .B(n39024), .Z(n39023) );
  XOR U38668 ( .A(n39025), .B(n39022), .Z(n39024) );
  XNOR U38669 ( .A(n38645), .B(n39018), .Z(n39020) );
  XOR U38670 ( .A(n39026), .B(n39027), .Z(n38645) );
  AND U38671 ( .A(n589), .B(n39028), .Z(n39027) );
  XOR U38672 ( .A(n39029), .B(n39026), .Z(n39028) );
  XOR U38673 ( .A(n39030), .B(n39031), .Z(n39018) );
  AND U38674 ( .A(n39032), .B(n39033), .Z(n39031) );
  XOR U38675 ( .A(n39030), .B(n38660), .Z(n39033) );
  XOR U38676 ( .A(n39034), .B(n39035), .Z(n38660) );
  AND U38677 ( .A(n591), .B(n39036), .Z(n39035) );
  XOR U38678 ( .A(n39037), .B(n39034), .Z(n39036) );
  XNOR U38679 ( .A(n38657), .B(n39030), .Z(n39032) );
  XOR U38680 ( .A(n39038), .B(n39039), .Z(n38657) );
  AND U38681 ( .A(n589), .B(n39040), .Z(n39039) );
  XOR U38682 ( .A(n39041), .B(n39038), .Z(n39040) );
  XOR U38683 ( .A(n39042), .B(n39043), .Z(n39030) );
  AND U38684 ( .A(n39044), .B(n39045), .Z(n39043) );
  XOR U38685 ( .A(n39042), .B(n38672), .Z(n39045) );
  XOR U38686 ( .A(n39046), .B(n39047), .Z(n38672) );
  AND U38687 ( .A(n591), .B(n39048), .Z(n39047) );
  XOR U38688 ( .A(n39049), .B(n39046), .Z(n39048) );
  XNOR U38689 ( .A(n38669), .B(n39042), .Z(n39044) );
  XOR U38690 ( .A(n39050), .B(n39051), .Z(n38669) );
  AND U38691 ( .A(n589), .B(n39052), .Z(n39051) );
  XOR U38692 ( .A(n39053), .B(n39050), .Z(n39052) );
  XOR U38693 ( .A(n39054), .B(n39055), .Z(n39042) );
  AND U38694 ( .A(n39056), .B(n39057), .Z(n39055) );
  XOR U38695 ( .A(n39054), .B(n38684), .Z(n39057) );
  XOR U38696 ( .A(n39058), .B(n39059), .Z(n38684) );
  AND U38697 ( .A(n591), .B(n39060), .Z(n39059) );
  XOR U38698 ( .A(n39061), .B(n39058), .Z(n39060) );
  XNOR U38699 ( .A(n38681), .B(n39054), .Z(n39056) );
  XOR U38700 ( .A(n39062), .B(n39063), .Z(n38681) );
  AND U38701 ( .A(n589), .B(n39064), .Z(n39063) );
  XOR U38702 ( .A(n39065), .B(n39062), .Z(n39064) );
  XOR U38703 ( .A(n39066), .B(n39067), .Z(n39054) );
  AND U38704 ( .A(n39068), .B(n39069), .Z(n39067) );
  XOR U38705 ( .A(n39066), .B(n38696), .Z(n39069) );
  XOR U38706 ( .A(n39070), .B(n39071), .Z(n38696) );
  AND U38707 ( .A(n591), .B(n39072), .Z(n39071) );
  XOR U38708 ( .A(n39073), .B(n39070), .Z(n39072) );
  XNOR U38709 ( .A(n38693), .B(n39066), .Z(n39068) );
  XOR U38710 ( .A(n39074), .B(n39075), .Z(n38693) );
  AND U38711 ( .A(n589), .B(n39076), .Z(n39075) );
  XOR U38712 ( .A(n39077), .B(n39074), .Z(n39076) );
  XOR U38713 ( .A(n39078), .B(n39079), .Z(n39066) );
  AND U38714 ( .A(n39080), .B(n39081), .Z(n39079) );
  XNOR U38715 ( .A(n39082), .B(n38709), .Z(n39081) );
  XOR U38716 ( .A(n39083), .B(n39084), .Z(n38709) );
  AND U38717 ( .A(n591), .B(n39085), .Z(n39084) );
  XOR U38718 ( .A(n39083), .B(n39086), .Z(n39085) );
  XNOR U38719 ( .A(n38706), .B(n39078), .Z(n39080) );
  XOR U38720 ( .A(n39087), .B(n39088), .Z(n38706) );
  AND U38721 ( .A(n589), .B(n39089), .Z(n39088) );
  XOR U38722 ( .A(n39087), .B(n39090), .Z(n39089) );
  IV U38723 ( .A(n39082), .Z(n39078) );
  AND U38724 ( .A(n38714), .B(n38717), .Z(n39082) );
  XNOR U38725 ( .A(n39091), .B(n39092), .Z(n38717) );
  AND U38726 ( .A(n591), .B(n39093), .Z(n39092) );
  XNOR U38727 ( .A(n39094), .B(n39091), .Z(n39093) );
  XOR U38728 ( .A(n39095), .B(n39096), .Z(n591) );
  AND U38729 ( .A(n39097), .B(n39098), .Z(n39096) );
  XOR U38730 ( .A(n38725), .B(n39095), .Z(n39098) );
  IV U38731 ( .A(n39099), .Z(n38725) );
  AND U38732 ( .A(p_input[3071]), .B(p_input[3039]), .Z(n39099) );
  XOR U38733 ( .A(n39095), .B(n38722), .Z(n39097) );
  AND U38734 ( .A(p_input[2975]), .B(p_input[3007]), .Z(n38722) );
  XOR U38735 ( .A(n39100), .B(n39101), .Z(n39095) );
  AND U38736 ( .A(n39102), .B(n39103), .Z(n39101) );
  XOR U38737 ( .A(n39100), .B(n38737), .Z(n39103) );
  XNOR U38738 ( .A(p_input[3038]), .B(n39104), .Z(n38737) );
  AND U38739 ( .A(n751), .B(n39105), .Z(n39104) );
  XOR U38740 ( .A(p_input[3070]), .B(p_input[3038]), .Z(n39105) );
  XNOR U38741 ( .A(n38734), .B(n39100), .Z(n39102) );
  XOR U38742 ( .A(n39106), .B(n39107), .Z(n38734) );
  AND U38743 ( .A(n749), .B(n39108), .Z(n39107) );
  XOR U38744 ( .A(p_input[3006]), .B(p_input[2974]), .Z(n39108) );
  XOR U38745 ( .A(n39109), .B(n39110), .Z(n39100) );
  AND U38746 ( .A(n39111), .B(n39112), .Z(n39110) );
  XOR U38747 ( .A(n39109), .B(n38749), .Z(n39112) );
  XNOR U38748 ( .A(p_input[3037]), .B(n39113), .Z(n38749) );
  AND U38749 ( .A(n751), .B(n39114), .Z(n39113) );
  XOR U38750 ( .A(p_input[3069]), .B(p_input[3037]), .Z(n39114) );
  XNOR U38751 ( .A(n38746), .B(n39109), .Z(n39111) );
  XOR U38752 ( .A(n39115), .B(n39116), .Z(n38746) );
  AND U38753 ( .A(n749), .B(n39117), .Z(n39116) );
  XOR U38754 ( .A(p_input[3005]), .B(p_input[2973]), .Z(n39117) );
  XOR U38755 ( .A(n39118), .B(n39119), .Z(n39109) );
  AND U38756 ( .A(n39120), .B(n39121), .Z(n39119) );
  XOR U38757 ( .A(n39118), .B(n38761), .Z(n39121) );
  XNOR U38758 ( .A(p_input[3036]), .B(n39122), .Z(n38761) );
  AND U38759 ( .A(n751), .B(n39123), .Z(n39122) );
  XOR U38760 ( .A(p_input[3068]), .B(p_input[3036]), .Z(n39123) );
  XNOR U38761 ( .A(n38758), .B(n39118), .Z(n39120) );
  XOR U38762 ( .A(n39124), .B(n39125), .Z(n38758) );
  AND U38763 ( .A(n749), .B(n39126), .Z(n39125) );
  XOR U38764 ( .A(p_input[3004]), .B(p_input[2972]), .Z(n39126) );
  XOR U38765 ( .A(n39127), .B(n39128), .Z(n39118) );
  AND U38766 ( .A(n39129), .B(n39130), .Z(n39128) );
  XOR U38767 ( .A(n39127), .B(n38773), .Z(n39130) );
  XNOR U38768 ( .A(p_input[3035]), .B(n39131), .Z(n38773) );
  AND U38769 ( .A(n751), .B(n39132), .Z(n39131) );
  XOR U38770 ( .A(p_input[3067]), .B(p_input[3035]), .Z(n39132) );
  XNOR U38771 ( .A(n38770), .B(n39127), .Z(n39129) );
  XOR U38772 ( .A(n39133), .B(n39134), .Z(n38770) );
  AND U38773 ( .A(n749), .B(n39135), .Z(n39134) );
  XOR U38774 ( .A(p_input[3003]), .B(p_input[2971]), .Z(n39135) );
  XOR U38775 ( .A(n39136), .B(n39137), .Z(n39127) );
  AND U38776 ( .A(n39138), .B(n39139), .Z(n39137) );
  XOR U38777 ( .A(n39136), .B(n38785), .Z(n39139) );
  XNOR U38778 ( .A(p_input[3034]), .B(n39140), .Z(n38785) );
  AND U38779 ( .A(n751), .B(n39141), .Z(n39140) );
  XOR U38780 ( .A(p_input[3066]), .B(p_input[3034]), .Z(n39141) );
  XNOR U38781 ( .A(n38782), .B(n39136), .Z(n39138) );
  XOR U38782 ( .A(n39142), .B(n39143), .Z(n38782) );
  AND U38783 ( .A(n749), .B(n39144), .Z(n39143) );
  XOR U38784 ( .A(p_input[3002]), .B(p_input[2970]), .Z(n39144) );
  XOR U38785 ( .A(n39145), .B(n39146), .Z(n39136) );
  AND U38786 ( .A(n39147), .B(n39148), .Z(n39146) );
  XOR U38787 ( .A(n39145), .B(n38797), .Z(n39148) );
  XNOR U38788 ( .A(p_input[3033]), .B(n39149), .Z(n38797) );
  AND U38789 ( .A(n751), .B(n39150), .Z(n39149) );
  XOR U38790 ( .A(p_input[3065]), .B(p_input[3033]), .Z(n39150) );
  XNOR U38791 ( .A(n38794), .B(n39145), .Z(n39147) );
  XOR U38792 ( .A(n39151), .B(n39152), .Z(n38794) );
  AND U38793 ( .A(n749), .B(n39153), .Z(n39152) );
  XOR U38794 ( .A(p_input[3001]), .B(p_input[2969]), .Z(n39153) );
  XOR U38795 ( .A(n39154), .B(n39155), .Z(n39145) );
  AND U38796 ( .A(n39156), .B(n39157), .Z(n39155) );
  XOR U38797 ( .A(n39154), .B(n38809), .Z(n39157) );
  XNOR U38798 ( .A(p_input[3032]), .B(n39158), .Z(n38809) );
  AND U38799 ( .A(n751), .B(n39159), .Z(n39158) );
  XOR U38800 ( .A(p_input[3064]), .B(p_input[3032]), .Z(n39159) );
  XNOR U38801 ( .A(n38806), .B(n39154), .Z(n39156) );
  XOR U38802 ( .A(n39160), .B(n39161), .Z(n38806) );
  AND U38803 ( .A(n749), .B(n39162), .Z(n39161) );
  XOR U38804 ( .A(p_input[3000]), .B(p_input[2968]), .Z(n39162) );
  XOR U38805 ( .A(n39163), .B(n39164), .Z(n39154) );
  AND U38806 ( .A(n39165), .B(n39166), .Z(n39164) );
  XOR U38807 ( .A(n39163), .B(n38821), .Z(n39166) );
  XNOR U38808 ( .A(p_input[3031]), .B(n39167), .Z(n38821) );
  AND U38809 ( .A(n751), .B(n39168), .Z(n39167) );
  XOR U38810 ( .A(p_input[3063]), .B(p_input[3031]), .Z(n39168) );
  XNOR U38811 ( .A(n38818), .B(n39163), .Z(n39165) );
  XOR U38812 ( .A(n39169), .B(n39170), .Z(n38818) );
  AND U38813 ( .A(n749), .B(n39171), .Z(n39170) );
  XOR U38814 ( .A(p_input[2999]), .B(p_input[2967]), .Z(n39171) );
  XOR U38815 ( .A(n39172), .B(n39173), .Z(n39163) );
  AND U38816 ( .A(n39174), .B(n39175), .Z(n39173) );
  XOR U38817 ( .A(n39172), .B(n38833), .Z(n39175) );
  XNOR U38818 ( .A(p_input[3030]), .B(n39176), .Z(n38833) );
  AND U38819 ( .A(n751), .B(n39177), .Z(n39176) );
  XOR U38820 ( .A(p_input[3062]), .B(p_input[3030]), .Z(n39177) );
  XNOR U38821 ( .A(n38830), .B(n39172), .Z(n39174) );
  XOR U38822 ( .A(n39178), .B(n39179), .Z(n38830) );
  AND U38823 ( .A(n749), .B(n39180), .Z(n39179) );
  XOR U38824 ( .A(p_input[2998]), .B(p_input[2966]), .Z(n39180) );
  XOR U38825 ( .A(n39181), .B(n39182), .Z(n39172) );
  AND U38826 ( .A(n39183), .B(n39184), .Z(n39182) );
  XOR U38827 ( .A(n39181), .B(n38845), .Z(n39184) );
  XNOR U38828 ( .A(p_input[3029]), .B(n39185), .Z(n38845) );
  AND U38829 ( .A(n751), .B(n39186), .Z(n39185) );
  XOR U38830 ( .A(p_input[3061]), .B(p_input[3029]), .Z(n39186) );
  XNOR U38831 ( .A(n38842), .B(n39181), .Z(n39183) );
  XOR U38832 ( .A(n39187), .B(n39188), .Z(n38842) );
  AND U38833 ( .A(n749), .B(n39189), .Z(n39188) );
  XOR U38834 ( .A(p_input[2997]), .B(p_input[2965]), .Z(n39189) );
  XOR U38835 ( .A(n39190), .B(n39191), .Z(n39181) );
  AND U38836 ( .A(n39192), .B(n39193), .Z(n39191) );
  XOR U38837 ( .A(n39190), .B(n38857), .Z(n39193) );
  XNOR U38838 ( .A(p_input[3028]), .B(n39194), .Z(n38857) );
  AND U38839 ( .A(n751), .B(n39195), .Z(n39194) );
  XOR U38840 ( .A(p_input[3060]), .B(p_input[3028]), .Z(n39195) );
  XNOR U38841 ( .A(n38854), .B(n39190), .Z(n39192) );
  XOR U38842 ( .A(n39196), .B(n39197), .Z(n38854) );
  AND U38843 ( .A(n749), .B(n39198), .Z(n39197) );
  XOR U38844 ( .A(p_input[2996]), .B(p_input[2964]), .Z(n39198) );
  XOR U38845 ( .A(n39199), .B(n39200), .Z(n39190) );
  AND U38846 ( .A(n39201), .B(n39202), .Z(n39200) );
  XOR U38847 ( .A(n39199), .B(n38869), .Z(n39202) );
  XNOR U38848 ( .A(p_input[3027]), .B(n39203), .Z(n38869) );
  AND U38849 ( .A(n751), .B(n39204), .Z(n39203) );
  XOR U38850 ( .A(p_input[3059]), .B(p_input[3027]), .Z(n39204) );
  XNOR U38851 ( .A(n38866), .B(n39199), .Z(n39201) );
  XOR U38852 ( .A(n39205), .B(n39206), .Z(n38866) );
  AND U38853 ( .A(n749), .B(n39207), .Z(n39206) );
  XOR U38854 ( .A(p_input[2995]), .B(p_input[2963]), .Z(n39207) );
  XOR U38855 ( .A(n39208), .B(n39209), .Z(n39199) );
  AND U38856 ( .A(n39210), .B(n39211), .Z(n39209) );
  XOR U38857 ( .A(n39208), .B(n38881), .Z(n39211) );
  XNOR U38858 ( .A(p_input[3026]), .B(n39212), .Z(n38881) );
  AND U38859 ( .A(n751), .B(n39213), .Z(n39212) );
  XOR U38860 ( .A(p_input[3058]), .B(p_input[3026]), .Z(n39213) );
  XNOR U38861 ( .A(n38878), .B(n39208), .Z(n39210) );
  XOR U38862 ( .A(n39214), .B(n39215), .Z(n38878) );
  AND U38863 ( .A(n749), .B(n39216), .Z(n39215) );
  XOR U38864 ( .A(p_input[2994]), .B(p_input[2962]), .Z(n39216) );
  XOR U38865 ( .A(n39217), .B(n39218), .Z(n39208) );
  AND U38866 ( .A(n39219), .B(n39220), .Z(n39218) );
  XOR U38867 ( .A(n39217), .B(n38893), .Z(n39220) );
  XNOR U38868 ( .A(p_input[3025]), .B(n39221), .Z(n38893) );
  AND U38869 ( .A(n751), .B(n39222), .Z(n39221) );
  XOR U38870 ( .A(p_input[3057]), .B(p_input[3025]), .Z(n39222) );
  XNOR U38871 ( .A(n38890), .B(n39217), .Z(n39219) );
  XOR U38872 ( .A(n39223), .B(n39224), .Z(n38890) );
  AND U38873 ( .A(n749), .B(n39225), .Z(n39224) );
  XOR U38874 ( .A(p_input[2993]), .B(p_input[2961]), .Z(n39225) );
  XOR U38875 ( .A(n39226), .B(n39227), .Z(n39217) );
  AND U38876 ( .A(n39228), .B(n39229), .Z(n39227) );
  XOR U38877 ( .A(n39226), .B(n38905), .Z(n39229) );
  XNOR U38878 ( .A(p_input[3024]), .B(n39230), .Z(n38905) );
  AND U38879 ( .A(n751), .B(n39231), .Z(n39230) );
  XOR U38880 ( .A(p_input[3056]), .B(p_input[3024]), .Z(n39231) );
  XNOR U38881 ( .A(n38902), .B(n39226), .Z(n39228) );
  XOR U38882 ( .A(n39232), .B(n39233), .Z(n38902) );
  AND U38883 ( .A(n749), .B(n39234), .Z(n39233) );
  XOR U38884 ( .A(p_input[2992]), .B(p_input[2960]), .Z(n39234) );
  XOR U38885 ( .A(n39235), .B(n39236), .Z(n39226) );
  AND U38886 ( .A(n39237), .B(n39238), .Z(n39236) );
  XOR U38887 ( .A(n39235), .B(n38917), .Z(n39238) );
  XNOR U38888 ( .A(p_input[3023]), .B(n39239), .Z(n38917) );
  AND U38889 ( .A(n751), .B(n39240), .Z(n39239) );
  XOR U38890 ( .A(p_input[3055]), .B(p_input[3023]), .Z(n39240) );
  XNOR U38891 ( .A(n38914), .B(n39235), .Z(n39237) );
  XOR U38892 ( .A(n39241), .B(n39242), .Z(n38914) );
  AND U38893 ( .A(n749), .B(n39243), .Z(n39242) );
  XOR U38894 ( .A(p_input[2991]), .B(p_input[2959]), .Z(n39243) );
  XOR U38895 ( .A(n39244), .B(n39245), .Z(n39235) );
  AND U38896 ( .A(n39246), .B(n39247), .Z(n39245) );
  XOR U38897 ( .A(n39244), .B(n38929), .Z(n39247) );
  XNOR U38898 ( .A(p_input[3022]), .B(n39248), .Z(n38929) );
  AND U38899 ( .A(n751), .B(n39249), .Z(n39248) );
  XOR U38900 ( .A(p_input[3054]), .B(p_input[3022]), .Z(n39249) );
  XNOR U38901 ( .A(n38926), .B(n39244), .Z(n39246) );
  XOR U38902 ( .A(n39250), .B(n39251), .Z(n38926) );
  AND U38903 ( .A(n749), .B(n39252), .Z(n39251) );
  XOR U38904 ( .A(p_input[2990]), .B(p_input[2958]), .Z(n39252) );
  XOR U38905 ( .A(n39253), .B(n39254), .Z(n39244) );
  AND U38906 ( .A(n39255), .B(n39256), .Z(n39254) );
  XOR U38907 ( .A(n39253), .B(n38941), .Z(n39256) );
  XNOR U38908 ( .A(p_input[3021]), .B(n39257), .Z(n38941) );
  AND U38909 ( .A(n751), .B(n39258), .Z(n39257) );
  XOR U38910 ( .A(p_input[3053]), .B(p_input[3021]), .Z(n39258) );
  XNOR U38911 ( .A(n38938), .B(n39253), .Z(n39255) );
  XOR U38912 ( .A(n39259), .B(n39260), .Z(n38938) );
  AND U38913 ( .A(n749), .B(n39261), .Z(n39260) );
  XOR U38914 ( .A(p_input[2989]), .B(p_input[2957]), .Z(n39261) );
  XOR U38915 ( .A(n39262), .B(n39263), .Z(n39253) );
  AND U38916 ( .A(n39264), .B(n39265), .Z(n39263) );
  XOR U38917 ( .A(n39262), .B(n38953), .Z(n39265) );
  XNOR U38918 ( .A(p_input[3020]), .B(n39266), .Z(n38953) );
  AND U38919 ( .A(n751), .B(n39267), .Z(n39266) );
  XOR U38920 ( .A(p_input[3052]), .B(p_input[3020]), .Z(n39267) );
  XNOR U38921 ( .A(n38950), .B(n39262), .Z(n39264) );
  XOR U38922 ( .A(n39268), .B(n39269), .Z(n38950) );
  AND U38923 ( .A(n749), .B(n39270), .Z(n39269) );
  XOR U38924 ( .A(p_input[2988]), .B(p_input[2956]), .Z(n39270) );
  XOR U38925 ( .A(n39271), .B(n39272), .Z(n39262) );
  AND U38926 ( .A(n39273), .B(n39274), .Z(n39272) );
  XOR U38927 ( .A(n39271), .B(n38965), .Z(n39274) );
  XNOR U38928 ( .A(p_input[3019]), .B(n39275), .Z(n38965) );
  AND U38929 ( .A(n751), .B(n39276), .Z(n39275) );
  XOR U38930 ( .A(p_input[3051]), .B(p_input[3019]), .Z(n39276) );
  XNOR U38931 ( .A(n38962), .B(n39271), .Z(n39273) );
  XOR U38932 ( .A(n39277), .B(n39278), .Z(n38962) );
  AND U38933 ( .A(n749), .B(n39279), .Z(n39278) );
  XOR U38934 ( .A(p_input[2987]), .B(p_input[2955]), .Z(n39279) );
  XOR U38935 ( .A(n39280), .B(n39281), .Z(n39271) );
  AND U38936 ( .A(n39282), .B(n39283), .Z(n39281) );
  XOR U38937 ( .A(n39280), .B(n38977), .Z(n39283) );
  XNOR U38938 ( .A(p_input[3018]), .B(n39284), .Z(n38977) );
  AND U38939 ( .A(n751), .B(n39285), .Z(n39284) );
  XOR U38940 ( .A(p_input[3050]), .B(p_input[3018]), .Z(n39285) );
  XNOR U38941 ( .A(n38974), .B(n39280), .Z(n39282) );
  XOR U38942 ( .A(n39286), .B(n39287), .Z(n38974) );
  AND U38943 ( .A(n749), .B(n39288), .Z(n39287) );
  XOR U38944 ( .A(p_input[2986]), .B(p_input[2954]), .Z(n39288) );
  XOR U38945 ( .A(n39289), .B(n39290), .Z(n39280) );
  AND U38946 ( .A(n39291), .B(n39292), .Z(n39290) );
  XOR U38947 ( .A(n39289), .B(n38989), .Z(n39292) );
  XNOR U38948 ( .A(p_input[3017]), .B(n39293), .Z(n38989) );
  AND U38949 ( .A(n751), .B(n39294), .Z(n39293) );
  XOR U38950 ( .A(p_input[3049]), .B(p_input[3017]), .Z(n39294) );
  XNOR U38951 ( .A(n38986), .B(n39289), .Z(n39291) );
  XOR U38952 ( .A(n39295), .B(n39296), .Z(n38986) );
  AND U38953 ( .A(n749), .B(n39297), .Z(n39296) );
  XOR U38954 ( .A(p_input[2985]), .B(p_input[2953]), .Z(n39297) );
  XOR U38955 ( .A(n39298), .B(n39299), .Z(n39289) );
  AND U38956 ( .A(n39300), .B(n39301), .Z(n39299) );
  XOR U38957 ( .A(n39298), .B(n39001), .Z(n39301) );
  XNOR U38958 ( .A(p_input[3016]), .B(n39302), .Z(n39001) );
  AND U38959 ( .A(n751), .B(n39303), .Z(n39302) );
  XOR U38960 ( .A(p_input[3048]), .B(p_input[3016]), .Z(n39303) );
  XNOR U38961 ( .A(n38998), .B(n39298), .Z(n39300) );
  XOR U38962 ( .A(n39304), .B(n39305), .Z(n38998) );
  AND U38963 ( .A(n749), .B(n39306), .Z(n39305) );
  XOR U38964 ( .A(p_input[2984]), .B(p_input[2952]), .Z(n39306) );
  XOR U38965 ( .A(n39307), .B(n39308), .Z(n39298) );
  AND U38966 ( .A(n39309), .B(n39310), .Z(n39308) );
  XOR U38967 ( .A(n39307), .B(n39013), .Z(n39310) );
  XNOR U38968 ( .A(p_input[3015]), .B(n39311), .Z(n39013) );
  AND U38969 ( .A(n751), .B(n39312), .Z(n39311) );
  XOR U38970 ( .A(p_input[3047]), .B(p_input[3015]), .Z(n39312) );
  XNOR U38971 ( .A(n39010), .B(n39307), .Z(n39309) );
  XOR U38972 ( .A(n39313), .B(n39314), .Z(n39010) );
  AND U38973 ( .A(n749), .B(n39315), .Z(n39314) );
  XOR U38974 ( .A(p_input[2983]), .B(p_input[2951]), .Z(n39315) );
  XOR U38975 ( .A(n39316), .B(n39317), .Z(n39307) );
  AND U38976 ( .A(n39318), .B(n39319), .Z(n39317) );
  XOR U38977 ( .A(n39316), .B(n39025), .Z(n39319) );
  XNOR U38978 ( .A(p_input[3014]), .B(n39320), .Z(n39025) );
  AND U38979 ( .A(n751), .B(n39321), .Z(n39320) );
  XOR U38980 ( .A(p_input[3046]), .B(p_input[3014]), .Z(n39321) );
  XNOR U38981 ( .A(n39022), .B(n39316), .Z(n39318) );
  XOR U38982 ( .A(n39322), .B(n39323), .Z(n39022) );
  AND U38983 ( .A(n749), .B(n39324), .Z(n39323) );
  XOR U38984 ( .A(p_input[2982]), .B(p_input[2950]), .Z(n39324) );
  XOR U38985 ( .A(n39325), .B(n39326), .Z(n39316) );
  AND U38986 ( .A(n39327), .B(n39328), .Z(n39326) );
  XOR U38987 ( .A(n39325), .B(n39037), .Z(n39328) );
  XNOR U38988 ( .A(p_input[3013]), .B(n39329), .Z(n39037) );
  AND U38989 ( .A(n751), .B(n39330), .Z(n39329) );
  XOR U38990 ( .A(p_input[3045]), .B(p_input[3013]), .Z(n39330) );
  XNOR U38991 ( .A(n39034), .B(n39325), .Z(n39327) );
  XOR U38992 ( .A(n39331), .B(n39332), .Z(n39034) );
  AND U38993 ( .A(n749), .B(n39333), .Z(n39332) );
  XOR U38994 ( .A(p_input[2981]), .B(p_input[2949]), .Z(n39333) );
  XOR U38995 ( .A(n39334), .B(n39335), .Z(n39325) );
  AND U38996 ( .A(n39336), .B(n39337), .Z(n39335) );
  XOR U38997 ( .A(n39334), .B(n39049), .Z(n39337) );
  XNOR U38998 ( .A(p_input[3012]), .B(n39338), .Z(n39049) );
  AND U38999 ( .A(n751), .B(n39339), .Z(n39338) );
  XOR U39000 ( .A(p_input[3044]), .B(p_input[3012]), .Z(n39339) );
  XNOR U39001 ( .A(n39046), .B(n39334), .Z(n39336) );
  XOR U39002 ( .A(n39340), .B(n39341), .Z(n39046) );
  AND U39003 ( .A(n749), .B(n39342), .Z(n39341) );
  XOR U39004 ( .A(p_input[2980]), .B(p_input[2948]), .Z(n39342) );
  XOR U39005 ( .A(n39343), .B(n39344), .Z(n39334) );
  AND U39006 ( .A(n39345), .B(n39346), .Z(n39344) );
  XOR U39007 ( .A(n39343), .B(n39061), .Z(n39346) );
  XNOR U39008 ( .A(p_input[3011]), .B(n39347), .Z(n39061) );
  AND U39009 ( .A(n751), .B(n39348), .Z(n39347) );
  XOR U39010 ( .A(p_input[3043]), .B(p_input[3011]), .Z(n39348) );
  XNOR U39011 ( .A(n39058), .B(n39343), .Z(n39345) );
  XOR U39012 ( .A(n39349), .B(n39350), .Z(n39058) );
  AND U39013 ( .A(n749), .B(n39351), .Z(n39350) );
  XOR U39014 ( .A(p_input[2979]), .B(p_input[2947]), .Z(n39351) );
  XOR U39015 ( .A(n39352), .B(n39353), .Z(n39343) );
  AND U39016 ( .A(n39354), .B(n39355), .Z(n39353) );
  XOR U39017 ( .A(n39352), .B(n39073), .Z(n39355) );
  XNOR U39018 ( .A(p_input[3010]), .B(n39356), .Z(n39073) );
  AND U39019 ( .A(n751), .B(n39357), .Z(n39356) );
  XOR U39020 ( .A(p_input[3042]), .B(p_input[3010]), .Z(n39357) );
  XNOR U39021 ( .A(n39070), .B(n39352), .Z(n39354) );
  XOR U39022 ( .A(n39358), .B(n39359), .Z(n39070) );
  AND U39023 ( .A(n749), .B(n39360), .Z(n39359) );
  XOR U39024 ( .A(p_input[2978]), .B(p_input[2946]), .Z(n39360) );
  XOR U39025 ( .A(n39361), .B(n39362), .Z(n39352) );
  AND U39026 ( .A(n39363), .B(n39364), .Z(n39362) );
  XNOR U39027 ( .A(n39365), .B(n39086), .Z(n39364) );
  XNOR U39028 ( .A(p_input[3009]), .B(n39366), .Z(n39086) );
  AND U39029 ( .A(n751), .B(n39367), .Z(n39366) );
  XNOR U39030 ( .A(p_input[3041]), .B(n39368), .Z(n39367) );
  IV U39031 ( .A(p_input[3009]), .Z(n39368) );
  XNOR U39032 ( .A(n39083), .B(n39361), .Z(n39363) );
  XNOR U39033 ( .A(p_input[2945]), .B(n39369), .Z(n39083) );
  AND U39034 ( .A(n749), .B(n39370), .Z(n39369) );
  XOR U39035 ( .A(p_input[2977]), .B(p_input[2945]), .Z(n39370) );
  IV U39036 ( .A(n39365), .Z(n39361) );
  AND U39037 ( .A(n39091), .B(n39094), .Z(n39365) );
  XOR U39038 ( .A(p_input[3008]), .B(n39371), .Z(n39094) );
  AND U39039 ( .A(n751), .B(n39372), .Z(n39371) );
  XOR U39040 ( .A(p_input[3040]), .B(p_input[3008]), .Z(n39372) );
  XOR U39041 ( .A(n39373), .B(n39374), .Z(n751) );
  AND U39042 ( .A(n39375), .B(n39376), .Z(n39374) );
  XNOR U39043 ( .A(p_input[3071]), .B(n39373), .Z(n39376) );
  XOR U39044 ( .A(n39373), .B(p_input[3039]), .Z(n39375) );
  XOR U39045 ( .A(n39377), .B(n39378), .Z(n39373) );
  AND U39046 ( .A(n39379), .B(n39380), .Z(n39378) );
  XNOR U39047 ( .A(p_input[3070]), .B(n39377), .Z(n39380) );
  XOR U39048 ( .A(n39377), .B(p_input[3038]), .Z(n39379) );
  XOR U39049 ( .A(n39381), .B(n39382), .Z(n39377) );
  AND U39050 ( .A(n39383), .B(n39384), .Z(n39382) );
  XNOR U39051 ( .A(p_input[3069]), .B(n39381), .Z(n39384) );
  XOR U39052 ( .A(n39381), .B(p_input[3037]), .Z(n39383) );
  XOR U39053 ( .A(n39385), .B(n39386), .Z(n39381) );
  AND U39054 ( .A(n39387), .B(n39388), .Z(n39386) );
  XNOR U39055 ( .A(p_input[3068]), .B(n39385), .Z(n39388) );
  XOR U39056 ( .A(n39385), .B(p_input[3036]), .Z(n39387) );
  XOR U39057 ( .A(n39389), .B(n39390), .Z(n39385) );
  AND U39058 ( .A(n39391), .B(n39392), .Z(n39390) );
  XNOR U39059 ( .A(p_input[3067]), .B(n39389), .Z(n39392) );
  XOR U39060 ( .A(n39389), .B(p_input[3035]), .Z(n39391) );
  XOR U39061 ( .A(n39393), .B(n39394), .Z(n39389) );
  AND U39062 ( .A(n39395), .B(n39396), .Z(n39394) );
  XNOR U39063 ( .A(p_input[3066]), .B(n39393), .Z(n39396) );
  XOR U39064 ( .A(n39393), .B(p_input[3034]), .Z(n39395) );
  XOR U39065 ( .A(n39397), .B(n39398), .Z(n39393) );
  AND U39066 ( .A(n39399), .B(n39400), .Z(n39398) );
  XNOR U39067 ( .A(p_input[3065]), .B(n39397), .Z(n39400) );
  XOR U39068 ( .A(n39397), .B(p_input[3033]), .Z(n39399) );
  XOR U39069 ( .A(n39401), .B(n39402), .Z(n39397) );
  AND U39070 ( .A(n39403), .B(n39404), .Z(n39402) );
  XNOR U39071 ( .A(p_input[3064]), .B(n39401), .Z(n39404) );
  XOR U39072 ( .A(n39401), .B(p_input[3032]), .Z(n39403) );
  XOR U39073 ( .A(n39405), .B(n39406), .Z(n39401) );
  AND U39074 ( .A(n39407), .B(n39408), .Z(n39406) );
  XNOR U39075 ( .A(p_input[3063]), .B(n39405), .Z(n39408) );
  XOR U39076 ( .A(n39405), .B(p_input[3031]), .Z(n39407) );
  XOR U39077 ( .A(n39409), .B(n39410), .Z(n39405) );
  AND U39078 ( .A(n39411), .B(n39412), .Z(n39410) );
  XNOR U39079 ( .A(p_input[3062]), .B(n39409), .Z(n39412) );
  XOR U39080 ( .A(n39409), .B(p_input[3030]), .Z(n39411) );
  XOR U39081 ( .A(n39413), .B(n39414), .Z(n39409) );
  AND U39082 ( .A(n39415), .B(n39416), .Z(n39414) );
  XNOR U39083 ( .A(p_input[3061]), .B(n39413), .Z(n39416) );
  XOR U39084 ( .A(n39413), .B(p_input[3029]), .Z(n39415) );
  XOR U39085 ( .A(n39417), .B(n39418), .Z(n39413) );
  AND U39086 ( .A(n39419), .B(n39420), .Z(n39418) );
  XNOR U39087 ( .A(p_input[3060]), .B(n39417), .Z(n39420) );
  XOR U39088 ( .A(n39417), .B(p_input[3028]), .Z(n39419) );
  XOR U39089 ( .A(n39421), .B(n39422), .Z(n39417) );
  AND U39090 ( .A(n39423), .B(n39424), .Z(n39422) );
  XNOR U39091 ( .A(p_input[3059]), .B(n39421), .Z(n39424) );
  XOR U39092 ( .A(n39421), .B(p_input[3027]), .Z(n39423) );
  XOR U39093 ( .A(n39425), .B(n39426), .Z(n39421) );
  AND U39094 ( .A(n39427), .B(n39428), .Z(n39426) );
  XNOR U39095 ( .A(p_input[3058]), .B(n39425), .Z(n39428) );
  XOR U39096 ( .A(n39425), .B(p_input[3026]), .Z(n39427) );
  XOR U39097 ( .A(n39429), .B(n39430), .Z(n39425) );
  AND U39098 ( .A(n39431), .B(n39432), .Z(n39430) );
  XNOR U39099 ( .A(p_input[3057]), .B(n39429), .Z(n39432) );
  XOR U39100 ( .A(n39429), .B(p_input[3025]), .Z(n39431) );
  XOR U39101 ( .A(n39433), .B(n39434), .Z(n39429) );
  AND U39102 ( .A(n39435), .B(n39436), .Z(n39434) );
  XNOR U39103 ( .A(p_input[3056]), .B(n39433), .Z(n39436) );
  XOR U39104 ( .A(n39433), .B(p_input[3024]), .Z(n39435) );
  XOR U39105 ( .A(n39437), .B(n39438), .Z(n39433) );
  AND U39106 ( .A(n39439), .B(n39440), .Z(n39438) );
  XNOR U39107 ( .A(p_input[3055]), .B(n39437), .Z(n39440) );
  XOR U39108 ( .A(n39437), .B(p_input[3023]), .Z(n39439) );
  XOR U39109 ( .A(n39441), .B(n39442), .Z(n39437) );
  AND U39110 ( .A(n39443), .B(n39444), .Z(n39442) );
  XNOR U39111 ( .A(p_input[3054]), .B(n39441), .Z(n39444) );
  XOR U39112 ( .A(n39441), .B(p_input[3022]), .Z(n39443) );
  XOR U39113 ( .A(n39445), .B(n39446), .Z(n39441) );
  AND U39114 ( .A(n39447), .B(n39448), .Z(n39446) );
  XNOR U39115 ( .A(p_input[3053]), .B(n39445), .Z(n39448) );
  XOR U39116 ( .A(n39445), .B(p_input[3021]), .Z(n39447) );
  XOR U39117 ( .A(n39449), .B(n39450), .Z(n39445) );
  AND U39118 ( .A(n39451), .B(n39452), .Z(n39450) );
  XNOR U39119 ( .A(p_input[3052]), .B(n39449), .Z(n39452) );
  XOR U39120 ( .A(n39449), .B(p_input[3020]), .Z(n39451) );
  XOR U39121 ( .A(n39453), .B(n39454), .Z(n39449) );
  AND U39122 ( .A(n39455), .B(n39456), .Z(n39454) );
  XNOR U39123 ( .A(p_input[3051]), .B(n39453), .Z(n39456) );
  XOR U39124 ( .A(n39453), .B(p_input[3019]), .Z(n39455) );
  XOR U39125 ( .A(n39457), .B(n39458), .Z(n39453) );
  AND U39126 ( .A(n39459), .B(n39460), .Z(n39458) );
  XNOR U39127 ( .A(p_input[3050]), .B(n39457), .Z(n39460) );
  XOR U39128 ( .A(n39457), .B(p_input[3018]), .Z(n39459) );
  XOR U39129 ( .A(n39461), .B(n39462), .Z(n39457) );
  AND U39130 ( .A(n39463), .B(n39464), .Z(n39462) );
  XNOR U39131 ( .A(p_input[3049]), .B(n39461), .Z(n39464) );
  XOR U39132 ( .A(n39461), .B(p_input[3017]), .Z(n39463) );
  XOR U39133 ( .A(n39465), .B(n39466), .Z(n39461) );
  AND U39134 ( .A(n39467), .B(n39468), .Z(n39466) );
  XNOR U39135 ( .A(p_input[3048]), .B(n39465), .Z(n39468) );
  XOR U39136 ( .A(n39465), .B(p_input[3016]), .Z(n39467) );
  XOR U39137 ( .A(n39469), .B(n39470), .Z(n39465) );
  AND U39138 ( .A(n39471), .B(n39472), .Z(n39470) );
  XNOR U39139 ( .A(p_input[3047]), .B(n39469), .Z(n39472) );
  XOR U39140 ( .A(n39469), .B(p_input[3015]), .Z(n39471) );
  XOR U39141 ( .A(n39473), .B(n39474), .Z(n39469) );
  AND U39142 ( .A(n39475), .B(n39476), .Z(n39474) );
  XNOR U39143 ( .A(p_input[3046]), .B(n39473), .Z(n39476) );
  XOR U39144 ( .A(n39473), .B(p_input[3014]), .Z(n39475) );
  XOR U39145 ( .A(n39477), .B(n39478), .Z(n39473) );
  AND U39146 ( .A(n39479), .B(n39480), .Z(n39478) );
  XNOR U39147 ( .A(p_input[3045]), .B(n39477), .Z(n39480) );
  XOR U39148 ( .A(n39477), .B(p_input[3013]), .Z(n39479) );
  XOR U39149 ( .A(n39481), .B(n39482), .Z(n39477) );
  AND U39150 ( .A(n39483), .B(n39484), .Z(n39482) );
  XNOR U39151 ( .A(p_input[3044]), .B(n39481), .Z(n39484) );
  XOR U39152 ( .A(n39481), .B(p_input[3012]), .Z(n39483) );
  XOR U39153 ( .A(n39485), .B(n39486), .Z(n39481) );
  AND U39154 ( .A(n39487), .B(n39488), .Z(n39486) );
  XNOR U39155 ( .A(p_input[3043]), .B(n39485), .Z(n39488) );
  XOR U39156 ( .A(n39485), .B(p_input[3011]), .Z(n39487) );
  XOR U39157 ( .A(n39489), .B(n39490), .Z(n39485) );
  AND U39158 ( .A(n39491), .B(n39492), .Z(n39490) );
  XNOR U39159 ( .A(p_input[3042]), .B(n39489), .Z(n39492) );
  XOR U39160 ( .A(n39489), .B(p_input[3010]), .Z(n39491) );
  XNOR U39161 ( .A(n39493), .B(n39494), .Z(n39489) );
  AND U39162 ( .A(n39495), .B(n39496), .Z(n39494) );
  XOR U39163 ( .A(p_input[3041]), .B(n39493), .Z(n39496) );
  XNOR U39164 ( .A(p_input[3009]), .B(n39493), .Z(n39495) );
  AND U39165 ( .A(p_input[3040]), .B(n39497), .Z(n39493) );
  IV U39166 ( .A(p_input[3008]), .Z(n39497) );
  XNOR U39167 ( .A(p_input[2944]), .B(n39498), .Z(n39091) );
  AND U39168 ( .A(n749), .B(n39499), .Z(n39498) );
  XOR U39169 ( .A(p_input[2976]), .B(p_input[2944]), .Z(n39499) );
  XOR U39170 ( .A(n39500), .B(n39501), .Z(n749) );
  AND U39171 ( .A(n39502), .B(n39503), .Z(n39501) );
  XNOR U39172 ( .A(p_input[3007]), .B(n39500), .Z(n39503) );
  XOR U39173 ( .A(n39500), .B(p_input[2975]), .Z(n39502) );
  XOR U39174 ( .A(n39504), .B(n39505), .Z(n39500) );
  AND U39175 ( .A(n39506), .B(n39507), .Z(n39505) );
  XNOR U39176 ( .A(p_input[3006]), .B(n39504), .Z(n39507) );
  XNOR U39177 ( .A(n39504), .B(n39106), .Z(n39506) );
  IV U39178 ( .A(p_input[2974]), .Z(n39106) );
  XOR U39179 ( .A(n39508), .B(n39509), .Z(n39504) );
  AND U39180 ( .A(n39510), .B(n39511), .Z(n39509) );
  XNOR U39181 ( .A(p_input[3005]), .B(n39508), .Z(n39511) );
  XNOR U39182 ( .A(n39508), .B(n39115), .Z(n39510) );
  IV U39183 ( .A(p_input[2973]), .Z(n39115) );
  XOR U39184 ( .A(n39512), .B(n39513), .Z(n39508) );
  AND U39185 ( .A(n39514), .B(n39515), .Z(n39513) );
  XNOR U39186 ( .A(p_input[3004]), .B(n39512), .Z(n39515) );
  XNOR U39187 ( .A(n39512), .B(n39124), .Z(n39514) );
  IV U39188 ( .A(p_input[2972]), .Z(n39124) );
  XOR U39189 ( .A(n39516), .B(n39517), .Z(n39512) );
  AND U39190 ( .A(n39518), .B(n39519), .Z(n39517) );
  XNOR U39191 ( .A(p_input[3003]), .B(n39516), .Z(n39519) );
  XNOR U39192 ( .A(n39516), .B(n39133), .Z(n39518) );
  IV U39193 ( .A(p_input[2971]), .Z(n39133) );
  XOR U39194 ( .A(n39520), .B(n39521), .Z(n39516) );
  AND U39195 ( .A(n39522), .B(n39523), .Z(n39521) );
  XNOR U39196 ( .A(p_input[3002]), .B(n39520), .Z(n39523) );
  XNOR U39197 ( .A(n39520), .B(n39142), .Z(n39522) );
  IV U39198 ( .A(p_input[2970]), .Z(n39142) );
  XOR U39199 ( .A(n39524), .B(n39525), .Z(n39520) );
  AND U39200 ( .A(n39526), .B(n39527), .Z(n39525) );
  XNOR U39201 ( .A(p_input[3001]), .B(n39524), .Z(n39527) );
  XNOR U39202 ( .A(n39524), .B(n39151), .Z(n39526) );
  IV U39203 ( .A(p_input[2969]), .Z(n39151) );
  XOR U39204 ( .A(n39528), .B(n39529), .Z(n39524) );
  AND U39205 ( .A(n39530), .B(n39531), .Z(n39529) );
  XNOR U39206 ( .A(p_input[3000]), .B(n39528), .Z(n39531) );
  XNOR U39207 ( .A(n39528), .B(n39160), .Z(n39530) );
  IV U39208 ( .A(p_input[2968]), .Z(n39160) );
  XOR U39209 ( .A(n39532), .B(n39533), .Z(n39528) );
  AND U39210 ( .A(n39534), .B(n39535), .Z(n39533) );
  XNOR U39211 ( .A(p_input[2999]), .B(n39532), .Z(n39535) );
  XNOR U39212 ( .A(n39532), .B(n39169), .Z(n39534) );
  IV U39213 ( .A(p_input[2967]), .Z(n39169) );
  XOR U39214 ( .A(n39536), .B(n39537), .Z(n39532) );
  AND U39215 ( .A(n39538), .B(n39539), .Z(n39537) );
  XNOR U39216 ( .A(p_input[2998]), .B(n39536), .Z(n39539) );
  XNOR U39217 ( .A(n39536), .B(n39178), .Z(n39538) );
  IV U39218 ( .A(p_input[2966]), .Z(n39178) );
  XOR U39219 ( .A(n39540), .B(n39541), .Z(n39536) );
  AND U39220 ( .A(n39542), .B(n39543), .Z(n39541) );
  XNOR U39221 ( .A(p_input[2997]), .B(n39540), .Z(n39543) );
  XNOR U39222 ( .A(n39540), .B(n39187), .Z(n39542) );
  IV U39223 ( .A(p_input[2965]), .Z(n39187) );
  XOR U39224 ( .A(n39544), .B(n39545), .Z(n39540) );
  AND U39225 ( .A(n39546), .B(n39547), .Z(n39545) );
  XNOR U39226 ( .A(p_input[2996]), .B(n39544), .Z(n39547) );
  XNOR U39227 ( .A(n39544), .B(n39196), .Z(n39546) );
  IV U39228 ( .A(p_input[2964]), .Z(n39196) );
  XOR U39229 ( .A(n39548), .B(n39549), .Z(n39544) );
  AND U39230 ( .A(n39550), .B(n39551), .Z(n39549) );
  XNOR U39231 ( .A(p_input[2995]), .B(n39548), .Z(n39551) );
  XNOR U39232 ( .A(n39548), .B(n39205), .Z(n39550) );
  IV U39233 ( .A(p_input[2963]), .Z(n39205) );
  XOR U39234 ( .A(n39552), .B(n39553), .Z(n39548) );
  AND U39235 ( .A(n39554), .B(n39555), .Z(n39553) );
  XNOR U39236 ( .A(p_input[2994]), .B(n39552), .Z(n39555) );
  XNOR U39237 ( .A(n39552), .B(n39214), .Z(n39554) );
  IV U39238 ( .A(p_input[2962]), .Z(n39214) );
  XOR U39239 ( .A(n39556), .B(n39557), .Z(n39552) );
  AND U39240 ( .A(n39558), .B(n39559), .Z(n39557) );
  XNOR U39241 ( .A(p_input[2993]), .B(n39556), .Z(n39559) );
  XNOR U39242 ( .A(n39556), .B(n39223), .Z(n39558) );
  IV U39243 ( .A(p_input[2961]), .Z(n39223) );
  XOR U39244 ( .A(n39560), .B(n39561), .Z(n39556) );
  AND U39245 ( .A(n39562), .B(n39563), .Z(n39561) );
  XNOR U39246 ( .A(p_input[2992]), .B(n39560), .Z(n39563) );
  XNOR U39247 ( .A(n39560), .B(n39232), .Z(n39562) );
  IV U39248 ( .A(p_input[2960]), .Z(n39232) );
  XOR U39249 ( .A(n39564), .B(n39565), .Z(n39560) );
  AND U39250 ( .A(n39566), .B(n39567), .Z(n39565) );
  XNOR U39251 ( .A(p_input[2991]), .B(n39564), .Z(n39567) );
  XNOR U39252 ( .A(n39564), .B(n39241), .Z(n39566) );
  IV U39253 ( .A(p_input[2959]), .Z(n39241) );
  XOR U39254 ( .A(n39568), .B(n39569), .Z(n39564) );
  AND U39255 ( .A(n39570), .B(n39571), .Z(n39569) );
  XNOR U39256 ( .A(p_input[2990]), .B(n39568), .Z(n39571) );
  XNOR U39257 ( .A(n39568), .B(n39250), .Z(n39570) );
  IV U39258 ( .A(p_input[2958]), .Z(n39250) );
  XOR U39259 ( .A(n39572), .B(n39573), .Z(n39568) );
  AND U39260 ( .A(n39574), .B(n39575), .Z(n39573) );
  XNOR U39261 ( .A(p_input[2989]), .B(n39572), .Z(n39575) );
  XNOR U39262 ( .A(n39572), .B(n39259), .Z(n39574) );
  IV U39263 ( .A(p_input[2957]), .Z(n39259) );
  XOR U39264 ( .A(n39576), .B(n39577), .Z(n39572) );
  AND U39265 ( .A(n39578), .B(n39579), .Z(n39577) );
  XNOR U39266 ( .A(p_input[2988]), .B(n39576), .Z(n39579) );
  XNOR U39267 ( .A(n39576), .B(n39268), .Z(n39578) );
  IV U39268 ( .A(p_input[2956]), .Z(n39268) );
  XOR U39269 ( .A(n39580), .B(n39581), .Z(n39576) );
  AND U39270 ( .A(n39582), .B(n39583), .Z(n39581) );
  XNOR U39271 ( .A(p_input[2987]), .B(n39580), .Z(n39583) );
  XNOR U39272 ( .A(n39580), .B(n39277), .Z(n39582) );
  IV U39273 ( .A(p_input[2955]), .Z(n39277) );
  XOR U39274 ( .A(n39584), .B(n39585), .Z(n39580) );
  AND U39275 ( .A(n39586), .B(n39587), .Z(n39585) );
  XNOR U39276 ( .A(p_input[2986]), .B(n39584), .Z(n39587) );
  XNOR U39277 ( .A(n39584), .B(n39286), .Z(n39586) );
  IV U39278 ( .A(p_input[2954]), .Z(n39286) );
  XOR U39279 ( .A(n39588), .B(n39589), .Z(n39584) );
  AND U39280 ( .A(n39590), .B(n39591), .Z(n39589) );
  XNOR U39281 ( .A(p_input[2985]), .B(n39588), .Z(n39591) );
  XNOR U39282 ( .A(n39588), .B(n39295), .Z(n39590) );
  IV U39283 ( .A(p_input[2953]), .Z(n39295) );
  XOR U39284 ( .A(n39592), .B(n39593), .Z(n39588) );
  AND U39285 ( .A(n39594), .B(n39595), .Z(n39593) );
  XNOR U39286 ( .A(p_input[2984]), .B(n39592), .Z(n39595) );
  XNOR U39287 ( .A(n39592), .B(n39304), .Z(n39594) );
  IV U39288 ( .A(p_input[2952]), .Z(n39304) );
  XOR U39289 ( .A(n39596), .B(n39597), .Z(n39592) );
  AND U39290 ( .A(n39598), .B(n39599), .Z(n39597) );
  XNOR U39291 ( .A(p_input[2983]), .B(n39596), .Z(n39599) );
  XNOR U39292 ( .A(n39596), .B(n39313), .Z(n39598) );
  IV U39293 ( .A(p_input[2951]), .Z(n39313) );
  XOR U39294 ( .A(n39600), .B(n39601), .Z(n39596) );
  AND U39295 ( .A(n39602), .B(n39603), .Z(n39601) );
  XNOR U39296 ( .A(p_input[2982]), .B(n39600), .Z(n39603) );
  XNOR U39297 ( .A(n39600), .B(n39322), .Z(n39602) );
  IV U39298 ( .A(p_input[2950]), .Z(n39322) );
  XOR U39299 ( .A(n39604), .B(n39605), .Z(n39600) );
  AND U39300 ( .A(n39606), .B(n39607), .Z(n39605) );
  XNOR U39301 ( .A(p_input[2981]), .B(n39604), .Z(n39607) );
  XNOR U39302 ( .A(n39604), .B(n39331), .Z(n39606) );
  IV U39303 ( .A(p_input[2949]), .Z(n39331) );
  XOR U39304 ( .A(n39608), .B(n39609), .Z(n39604) );
  AND U39305 ( .A(n39610), .B(n39611), .Z(n39609) );
  XNOR U39306 ( .A(p_input[2980]), .B(n39608), .Z(n39611) );
  XNOR U39307 ( .A(n39608), .B(n39340), .Z(n39610) );
  IV U39308 ( .A(p_input[2948]), .Z(n39340) );
  XOR U39309 ( .A(n39612), .B(n39613), .Z(n39608) );
  AND U39310 ( .A(n39614), .B(n39615), .Z(n39613) );
  XNOR U39311 ( .A(p_input[2979]), .B(n39612), .Z(n39615) );
  XNOR U39312 ( .A(n39612), .B(n39349), .Z(n39614) );
  IV U39313 ( .A(p_input[2947]), .Z(n39349) );
  XOR U39314 ( .A(n39616), .B(n39617), .Z(n39612) );
  AND U39315 ( .A(n39618), .B(n39619), .Z(n39617) );
  XNOR U39316 ( .A(p_input[2978]), .B(n39616), .Z(n39619) );
  XNOR U39317 ( .A(n39616), .B(n39358), .Z(n39618) );
  IV U39318 ( .A(p_input[2946]), .Z(n39358) );
  XNOR U39319 ( .A(n39620), .B(n39621), .Z(n39616) );
  AND U39320 ( .A(n39622), .B(n39623), .Z(n39621) );
  XOR U39321 ( .A(p_input[2977]), .B(n39620), .Z(n39623) );
  XNOR U39322 ( .A(p_input[2945]), .B(n39620), .Z(n39622) );
  AND U39323 ( .A(p_input[2976]), .B(n39624), .Z(n39620) );
  IV U39324 ( .A(p_input[2944]), .Z(n39624) );
  XOR U39325 ( .A(n39625), .B(n39626), .Z(n38714) );
  AND U39326 ( .A(n589), .B(n39627), .Z(n39626) );
  XNOR U39327 ( .A(n39628), .B(n39625), .Z(n39627) );
  XOR U39328 ( .A(n39629), .B(n39630), .Z(n589) );
  AND U39329 ( .A(n39631), .B(n39632), .Z(n39630) );
  XNOR U39330 ( .A(n38729), .B(n39629), .Z(n39632) );
  AND U39331 ( .A(p_input[2943]), .B(p_input[2911]), .Z(n38729) );
  XNOR U39332 ( .A(n39629), .B(n38726), .Z(n39631) );
  IV U39333 ( .A(n39633), .Z(n38726) );
  AND U39334 ( .A(p_input[2847]), .B(p_input[2879]), .Z(n39633) );
  XOR U39335 ( .A(n39634), .B(n39635), .Z(n39629) );
  AND U39336 ( .A(n39636), .B(n39637), .Z(n39635) );
  XOR U39337 ( .A(n39634), .B(n38741), .Z(n39637) );
  XNOR U39338 ( .A(p_input[2910]), .B(n39638), .Z(n38741) );
  AND U39339 ( .A(n755), .B(n39639), .Z(n39638) );
  XOR U39340 ( .A(p_input[2942]), .B(p_input[2910]), .Z(n39639) );
  XNOR U39341 ( .A(n38738), .B(n39634), .Z(n39636) );
  XOR U39342 ( .A(n39640), .B(n39641), .Z(n38738) );
  AND U39343 ( .A(n752), .B(n39642), .Z(n39641) );
  XOR U39344 ( .A(p_input[2878]), .B(p_input[2846]), .Z(n39642) );
  XOR U39345 ( .A(n39643), .B(n39644), .Z(n39634) );
  AND U39346 ( .A(n39645), .B(n39646), .Z(n39644) );
  XOR U39347 ( .A(n39643), .B(n38753), .Z(n39646) );
  XNOR U39348 ( .A(p_input[2909]), .B(n39647), .Z(n38753) );
  AND U39349 ( .A(n755), .B(n39648), .Z(n39647) );
  XOR U39350 ( .A(p_input[2941]), .B(p_input[2909]), .Z(n39648) );
  XNOR U39351 ( .A(n38750), .B(n39643), .Z(n39645) );
  XOR U39352 ( .A(n39649), .B(n39650), .Z(n38750) );
  AND U39353 ( .A(n752), .B(n39651), .Z(n39650) );
  XOR U39354 ( .A(p_input[2877]), .B(p_input[2845]), .Z(n39651) );
  XOR U39355 ( .A(n39652), .B(n39653), .Z(n39643) );
  AND U39356 ( .A(n39654), .B(n39655), .Z(n39653) );
  XOR U39357 ( .A(n39652), .B(n38765), .Z(n39655) );
  XNOR U39358 ( .A(p_input[2908]), .B(n39656), .Z(n38765) );
  AND U39359 ( .A(n755), .B(n39657), .Z(n39656) );
  XOR U39360 ( .A(p_input[2940]), .B(p_input[2908]), .Z(n39657) );
  XNOR U39361 ( .A(n38762), .B(n39652), .Z(n39654) );
  XOR U39362 ( .A(n39658), .B(n39659), .Z(n38762) );
  AND U39363 ( .A(n752), .B(n39660), .Z(n39659) );
  XOR U39364 ( .A(p_input[2876]), .B(p_input[2844]), .Z(n39660) );
  XOR U39365 ( .A(n39661), .B(n39662), .Z(n39652) );
  AND U39366 ( .A(n39663), .B(n39664), .Z(n39662) );
  XOR U39367 ( .A(n39661), .B(n38777), .Z(n39664) );
  XNOR U39368 ( .A(p_input[2907]), .B(n39665), .Z(n38777) );
  AND U39369 ( .A(n755), .B(n39666), .Z(n39665) );
  XOR U39370 ( .A(p_input[2939]), .B(p_input[2907]), .Z(n39666) );
  XNOR U39371 ( .A(n38774), .B(n39661), .Z(n39663) );
  XOR U39372 ( .A(n39667), .B(n39668), .Z(n38774) );
  AND U39373 ( .A(n752), .B(n39669), .Z(n39668) );
  XOR U39374 ( .A(p_input[2875]), .B(p_input[2843]), .Z(n39669) );
  XOR U39375 ( .A(n39670), .B(n39671), .Z(n39661) );
  AND U39376 ( .A(n39672), .B(n39673), .Z(n39671) );
  XOR U39377 ( .A(n39670), .B(n38789), .Z(n39673) );
  XNOR U39378 ( .A(p_input[2906]), .B(n39674), .Z(n38789) );
  AND U39379 ( .A(n755), .B(n39675), .Z(n39674) );
  XOR U39380 ( .A(p_input[2938]), .B(p_input[2906]), .Z(n39675) );
  XNOR U39381 ( .A(n38786), .B(n39670), .Z(n39672) );
  XOR U39382 ( .A(n39676), .B(n39677), .Z(n38786) );
  AND U39383 ( .A(n752), .B(n39678), .Z(n39677) );
  XOR U39384 ( .A(p_input[2874]), .B(p_input[2842]), .Z(n39678) );
  XOR U39385 ( .A(n39679), .B(n39680), .Z(n39670) );
  AND U39386 ( .A(n39681), .B(n39682), .Z(n39680) );
  XOR U39387 ( .A(n39679), .B(n38801), .Z(n39682) );
  XNOR U39388 ( .A(p_input[2905]), .B(n39683), .Z(n38801) );
  AND U39389 ( .A(n755), .B(n39684), .Z(n39683) );
  XOR U39390 ( .A(p_input[2937]), .B(p_input[2905]), .Z(n39684) );
  XNOR U39391 ( .A(n38798), .B(n39679), .Z(n39681) );
  XOR U39392 ( .A(n39685), .B(n39686), .Z(n38798) );
  AND U39393 ( .A(n752), .B(n39687), .Z(n39686) );
  XOR U39394 ( .A(p_input[2873]), .B(p_input[2841]), .Z(n39687) );
  XOR U39395 ( .A(n39688), .B(n39689), .Z(n39679) );
  AND U39396 ( .A(n39690), .B(n39691), .Z(n39689) );
  XOR U39397 ( .A(n39688), .B(n38813), .Z(n39691) );
  XNOR U39398 ( .A(p_input[2904]), .B(n39692), .Z(n38813) );
  AND U39399 ( .A(n755), .B(n39693), .Z(n39692) );
  XOR U39400 ( .A(p_input[2936]), .B(p_input[2904]), .Z(n39693) );
  XNOR U39401 ( .A(n38810), .B(n39688), .Z(n39690) );
  XOR U39402 ( .A(n39694), .B(n39695), .Z(n38810) );
  AND U39403 ( .A(n752), .B(n39696), .Z(n39695) );
  XOR U39404 ( .A(p_input[2872]), .B(p_input[2840]), .Z(n39696) );
  XOR U39405 ( .A(n39697), .B(n39698), .Z(n39688) );
  AND U39406 ( .A(n39699), .B(n39700), .Z(n39698) );
  XOR U39407 ( .A(n39697), .B(n38825), .Z(n39700) );
  XNOR U39408 ( .A(p_input[2903]), .B(n39701), .Z(n38825) );
  AND U39409 ( .A(n755), .B(n39702), .Z(n39701) );
  XOR U39410 ( .A(p_input[2935]), .B(p_input[2903]), .Z(n39702) );
  XNOR U39411 ( .A(n38822), .B(n39697), .Z(n39699) );
  XOR U39412 ( .A(n39703), .B(n39704), .Z(n38822) );
  AND U39413 ( .A(n752), .B(n39705), .Z(n39704) );
  XOR U39414 ( .A(p_input[2871]), .B(p_input[2839]), .Z(n39705) );
  XOR U39415 ( .A(n39706), .B(n39707), .Z(n39697) );
  AND U39416 ( .A(n39708), .B(n39709), .Z(n39707) );
  XOR U39417 ( .A(n39706), .B(n38837), .Z(n39709) );
  XNOR U39418 ( .A(p_input[2902]), .B(n39710), .Z(n38837) );
  AND U39419 ( .A(n755), .B(n39711), .Z(n39710) );
  XOR U39420 ( .A(p_input[2934]), .B(p_input[2902]), .Z(n39711) );
  XNOR U39421 ( .A(n38834), .B(n39706), .Z(n39708) );
  XOR U39422 ( .A(n39712), .B(n39713), .Z(n38834) );
  AND U39423 ( .A(n752), .B(n39714), .Z(n39713) );
  XOR U39424 ( .A(p_input[2870]), .B(p_input[2838]), .Z(n39714) );
  XOR U39425 ( .A(n39715), .B(n39716), .Z(n39706) );
  AND U39426 ( .A(n39717), .B(n39718), .Z(n39716) );
  XOR U39427 ( .A(n39715), .B(n38849), .Z(n39718) );
  XNOR U39428 ( .A(p_input[2901]), .B(n39719), .Z(n38849) );
  AND U39429 ( .A(n755), .B(n39720), .Z(n39719) );
  XOR U39430 ( .A(p_input[2933]), .B(p_input[2901]), .Z(n39720) );
  XNOR U39431 ( .A(n38846), .B(n39715), .Z(n39717) );
  XOR U39432 ( .A(n39721), .B(n39722), .Z(n38846) );
  AND U39433 ( .A(n752), .B(n39723), .Z(n39722) );
  XOR U39434 ( .A(p_input[2869]), .B(p_input[2837]), .Z(n39723) );
  XOR U39435 ( .A(n39724), .B(n39725), .Z(n39715) );
  AND U39436 ( .A(n39726), .B(n39727), .Z(n39725) );
  XOR U39437 ( .A(n39724), .B(n38861), .Z(n39727) );
  XNOR U39438 ( .A(p_input[2900]), .B(n39728), .Z(n38861) );
  AND U39439 ( .A(n755), .B(n39729), .Z(n39728) );
  XOR U39440 ( .A(p_input[2932]), .B(p_input[2900]), .Z(n39729) );
  XNOR U39441 ( .A(n38858), .B(n39724), .Z(n39726) );
  XOR U39442 ( .A(n39730), .B(n39731), .Z(n38858) );
  AND U39443 ( .A(n752), .B(n39732), .Z(n39731) );
  XOR U39444 ( .A(p_input[2868]), .B(p_input[2836]), .Z(n39732) );
  XOR U39445 ( .A(n39733), .B(n39734), .Z(n39724) );
  AND U39446 ( .A(n39735), .B(n39736), .Z(n39734) );
  XOR U39447 ( .A(n39733), .B(n38873), .Z(n39736) );
  XNOR U39448 ( .A(p_input[2899]), .B(n39737), .Z(n38873) );
  AND U39449 ( .A(n755), .B(n39738), .Z(n39737) );
  XOR U39450 ( .A(p_input[2931]), .B(p_input[2899]), .Z(n39738) );
  XNOR U39451 ( .A(n38870), .B(n39733), .Z(n39735) );
  XOR U39452 ( .A(n39739), .B(n39740), .Z(n38870) );
  AND U39453 ( .A(n752), .B(n39741), .Z(n39740) );
  XOR U39454 ( .A(p_input[2867]), .B(p_input[2835]), .Z(n39741) );
  XOR U39455 ( .A(n39742), .B(n39743), .Z(n39733) );
  AND U39456 ( .A(n39744), .B(n39745), .Z(n39743) );
  XOR U39457 ( .A(n39742), .B(n38885), .Z(n39745) );
  XNOR U39458 ( .A(p_input[2898]), .B(n39746), .Z(n38885) );
  AND U39459 ( .A(n755), .B(n39747), .Z(n39746) );
  XOR U39460 ( .A(p_input[2930]), .B(p_input[2898]), .Z(n39747) );
  XNOR U39461 ( .A(n38882), .B(n39742), .Z(n39744) );
  XOR U39462 ( .A(n39748), .B(n39749), .Z(n38882) );
  AND U39463 ( .A(n752), .B(n39750), .Z(n39749) );
  XOR U39464 ( .A(p_input[2866]), .B(p_input[2834]), .Z(n39750) );
  XOR U39465 ( .A(n39751), .B(n39752), .Z(n39742) );
  AND U39466 ( .A(n39753), .B(n39754), .Z(n39752) );
  XOR U39467 ( .A(n39751), .B(n38897), .Z(n39754) );
  XNOR U39468 ( .A(p_input[2897]), .B(n39755), .Z(n38897) );
  AND U39469 ( .A(n755), .B(n39756), .Z(n39755) );
  XOR U39470 ( .A(p_input[2929]), .B(p_input[2897]), .Z(n39756) );
  XNOR U39471 ( .A(n38894), .B(n39751), .Z(n39753) );
  XOR U39472 ( .A(n39757), .B(n39758), .Z(n38894) );
  AND U39473 ( .A(n752), .B(n39759), .Z(n39758) );
  XOR U39474 ( .A(p_input[2865]), .B(p_input[2833]), .Z(n39759) );
  XOR U39475 ( .A(n39760), .B(n39761), .Z(n39751) );
  AND U39476 ( .A(n39762), .B(n39763), .Z(n39761) );
  XOR U39477 ( .A(n39760), .B(n38909), .Z(n39763) );
  XNOR U39478 ( .A(p_input[2896]), .B(n39764), .Z(n38909) );
  AND U39479 ( .A(n755), .B(n39765), .Z(n39764) );
  XOR U39480 ( .A(p_input[2928]), .B(p_input[2896]), .Z(n39765) );
  XNOR U39481 ( .A(n38906), .B(n39760), .Z(n39762) );
  XOR U39482 ( .A(n39766), .B(n39767), .Z(n38906) );
  AND U39483 ( .A(n752), .B(n39768), .Z(n39767) );
  XOR U39484 ( .A(p_input[2864]), .B(p_input[2832]), .Z(n39768) );
  XOR U39485 ( .A(n39769), .B(n39770), .Z(n39760) );
  AND U39486 ( .A(n39771), .B(n39772), .Z(n39770) );
  XOR U39487 ( .A(n39769), .B(n38921), .Z(n39772) );
  XNOR U39488 ( .A(p_input[2895]), .B(n39773), .Z(n38921) );
  AND U39489 ( .A(n755), .B(n39774), .Z(n39773) );
  XOR U39490 ( .A(p_input[2927]), .B(p_input[2895]), .Z(n39774) );
  XNOR U39491 ( .A(n38918), .B(n39769), .Z(n39771) );
  XOR U39492 ( .A(n39775), .B(n39776), .Z(n38918) );
  AND U39493 ( .A(n752), .B(n39777), .Z(n39776) );
  XOR U39494 ( .A(p_input[2863]), .B(p_input[2831]), .Z(n39777) );
  XOR U39495 ( .A(n39778), .B(n39779), .Z(n39769) );
  AND U39496 ( .A(n39780), .B(n39781), .Z(n39779) );
  XOR U39497 ( .A(n39778), .B(n38933), .Z(n39781) );
  XNOR U39498 ( .A(p_input[2894]), .B(n39782), .Z(n38933) );
  AND U39499 ( .A(n755), .B(n39783), .Z(n39782) );
  XOR U39500 ( .A(p_input[2926]), .B(p_input[2894]), .Z(n39783) );
  XNOR U39501 ( .A(n38930), .B(n39778), .Z(n39780) );
  XOR U39502 ( .A(n39784), .B(n39785), .Z(n38930) );
  AND U39503 ( .A(n752), .B(n39786), .Z(n39785) );
  XOR U39504 ( .A(p_input[2862]), .B(p_input[2830]), .Z(n39786) );
  XOR U39505 ( .A(n39787), .B(n39788), .Z(n39778) );
  AND U39506 ( .A(n39789), .B(n39790), .Z(n39788) );
  XOR U39507 ( .A(n39787), .B(n38945), .Z(n39790) );
  XNOR U39508 ( .A(p_input[2893]), .B(n39791), .Z(n38945) );
  AND U39509 ( .A(n755), .B(n39792), .Z(n39791) );
  XOR U39510 ( .A(p_input[2925]), .B(p_input[2893]), .Z(n39792) );
  XNOR U39511 ( .A(n38942), .B(n39787), .Z(n39789) );
  XOR U39512 ( .A(n39793), .B(n39794), .Z(n38942) );
  AND U39513 ( .A(n752), .B(n39795), .Z(n39794) );
  XOR U39514 ( .A(p_input[2861]), .B(p_input[2829]), .Z(n39795) );
  XOR U39515 ( .A(n39796), .B(n39797), .Z(n39787) );
  AND U39516 ( .A(n39798), .B(n39799), .Z(n39797) );
  XOR U39517 ( .A(n39796), .B(n38957), .Z(n39799) );
  XNOR U39518 ( .A(p_input[2892]), .B(n39800), .Z(n38957) );
  AND U39519 ( .A(n755), .B(n39801), .Z(n39800) );
  XOR U39520 ( .A(p_input[2924]), .B(p_input[2892]), .Z(n39801) );
  XNOR U39521 ( .A(n38954), .B(n39796), .Z(n39798) );
  XOR U39522 ( .A(n39802), .B(n39803), .Z(n38954) );
  AND U39523 ( .A(n752), .B(n39804), .Z(n39803) );
  XOR U39524 ( .A(p_input[2860]), .B(p_input[2828]), .Z(n39804) );
  XOR U39525 ( .A(n39805), .B(n39806), .Z(n39796) );
  AND U39526 ( .A(n39807), .B(n39808), .Z(n39806) );
  XOR U39527 ( .A(n39805), .B(n38969), .Z(n39808) );
  XNOR U39528 ( .A(p_input[2891]), .B(n39809), .Z(n38969) );
  AND U39529 ( .A(n755), .B(n39810), .Z(n39809) );
  XOR U39530 ( .A(p_input[2923]), .B(p_input[2891]), .Z(n39810) );
  XNOR U39531 ( .A(n38966), .B(n39805), .Z(n39807) );
  XOR U39532 ( .A(n39811), .B(n39812), .Z(n38966) );
  AND U39533 ( .A(n752), .B(n39813), .Z(n39812) );
  XOR U39534 ( .A(p_input[2859]), .B(p_input[2827]), .Z(n39813) );
  XOR U39535 ( .A(n39814), .B(n39815), .Z(n39805) );
  AND U39536 ( .A(n39816), .B(n39817), .Z(n39815) );
  XOR U39537 ( .A(n39814), .B(n38981), .Z(n39817) );
  XNOR U39538 ( .A(p_input[2890]), .B(n39818), .Z(n38981) );
  AND U39539 ( .A(n755), .B(n39819), .Z(n39818) );
  XOR U39540 ( .A(p_input[2922]), .B(p_input[2890]), .Z(n39819) );
  XNOR U39541 ( .A(n38978), .B(n39814), .Z(n39816) );
  XOR U39542 ( .A(n39820), .B(n39821), .Z(n38978) );
  AND U39543 ( .A(n752), .B(n39822), .Z(n39821) );
  XOR U39544 ( .A(p_input[2858]), .B(p_input[2826]), .Z(n39822) );
  XOR U39545 ( .A(n39823), .B(n39824), .Z(n39814) );
  AND U39546 ( .A(n39825), .B(n39826), .Z(n39824) );
  XOR U39547 ( .A(n39823), .B(n38993), .Z(n39826) );
  XNOR U39548 ( .A(p_input[2889]), .B(n39827), .Z(n38993) );
  AND U39549 ( .A(n755), .B(n39828), .Z(n39827) );
  XOR U39550 ( .A(p_input[2921]), .B(p_input[2889]), .Z(n39828) );
  XNOR U39551 ( .A(n38990), .B(n39823), .Z(n39825) );
  XOR U39552 ( .A(n39829), .B(n39830), .Z(n38990) );
  AND U39553 ( .A(n752), .B(n39831), .Z(n39830) );
  XOR U39554 ( .A(p_input[2857]), .B(p_input[2825]), .Z(n39831) );
  XOR U39555 ( .A(n39832), .B(n39833), .Z(n39823) );
  AND U39556 ( .A(n39834), .B(n39835), .Z(n39833) );
  XOR U39557 ( .A(n39832), .B(n39005), .Z(n39835) );
  XNOR U39558 ( .A(p_input[2888]), .B(n39836), .Z(n39005) );
  AND U39559 ( .A(n755), .B(n39837), .Z(n39836) );
  XOR U39560 ( .A(p_input[2920]), .B(p_input[2888]), .Z(n39837) );
  XNOR U39561 ( .A(n39002), .B(n39832), .Z(n39834) );
  XOR U39562 ( .A(n39838), .B(n39839), .Z(n39002) );
  AND U39563 ( .A(n752), .B(n39840), .Z(n39839) );
  XOR U39564 ( .A(p_input[2856]), .B(p_input[2824]), .Z(n39840) );
  XOR U39565 ( .A(n39841), .B(n39842), .Z(n39832) );
  AND U39566 ( .A(n39843), .B(n39844), .Z(n39842) );
  XOR U39567 ( .A(n39841), .B(n39017), .Z(n39844) );
  XNOR U39568 ( .A(p_input[2887]), .B(n39845), .Z(n39017) );
  AND U39569 ( .A(n755), .B(n39846), .Z(n39845) );
  XOR U39570 ( .A(p_input[2919]), .B(p_input[2887]), .Z(n39846) );
  XNOR U39571 ( .A(n39014), .B(n39841), .Z(n39843) );
  XOR U39572 ( .A(n39847), .B(n39848), .Z(n39014) );
  AND U39573 ( .A(n752), .B(n39849), .Z(n39848) );
  XOR U39574 ( .A(p_input[2855]), .B(p_input[2823]), .Z(n39849) );
  XOR U39575 ( .A(n39850), .B(n39851), .Z(n39841) );
  AND U39576 ( .A(n39852), .B(n39853), .Z(n39851) );
  XOR U39577 ( .A(n39850), .B(n39029), .Z(n39853) );
  XNOR U39578 ( .A(p_input[2886]), .B(n39854), .Z(n39029) );
  AND U39579 ( .A(n755), .B(n39855), .Z(n39854) );
  XOR U39580 ( .A(p_input[2918]), .B(p_input[2886]), .Z(n39855) );
  XNOR U39581 ( .A(n39026), .B(n39850), .Z(n39852) );
  XOR U39582 ( .A(n39856), .B(n39857), .Z(n39026) );
  AND U39583 ( .A(n752), .B(n39858), .Z(n39857) );
  XOR U39584 ( .A(p_input[2854]), .B(p_input[2822]), .Z(n39858) );
  XOR U39585 ( .A(n39859), .B(n39860), .Z(n39850) );
  AND U39586 ( .A(n39861), .B(n39862), .Z(n39860) );
  XOR U39587 ( .A(n39859), .B(n39041), .Z(n39862) );
  XNOR U39588 ( .A(p_input[2885]), .B(n39863), .Z(n39041) );
  AND U39589 ( .A(n755), .B(n39864), .Z(n39863) );
  XOR U39590 ( .A(p_input[2917]), .B(p_input[2885]), .Z(n39864) );
  XNOR U39591 ( .A(n39038), .B(n39859), .Z(n39861) );
  XOR U39592 ( .A(n39865), .B(n39866), .Z(n39038) );
  AND U39593 ( .A(n752), .B(n39867), .Z(n39866) );
  XOR U39594 ( .A(p_input[2853]), .B(p_input[2821]), .Z(n39867) );
  XOR U39595 ( .A(n39868), .B(n39869), .Z(n39859) );
  AND U39596 ( .A(n39870), .B(n39871), .Z(n39869) );
  XOR U39597 ( .A(n39868), .B(n39053), .Z(n39871) );
  XNOR U39598 ( .A(p_input[2884]), .B(n39872), .Z(n39053) );
  AND U39599 ( .A(n755), .B(n39873), .Z(n39872) );
  XOR U39600 ( .A(p_input[2916]), .B(p_input[2884]), .Z(n39873) );
  XNOR U39601 ( .A(n39050), .B(n39868), .Z(n39870) );
  XOR U39602 ( .A(n39874), .B(n39875), .Z(n39050) );
  AND U39603 ( .A(n752), .B(n39876), .Z(n39875) );
  XOR U39604 ( .A(p_input[2852]), .B(p_input[2820]), .Z(n39876) );
  XOR U39605 ( .A(n39877), .B(n39878), .Z(n39868) );
  AND U39606 ( .A(n39879), .B(n39880), .Z(n39878) );
  XOR U39607 ( .A(n39877), .B(n39065), .Z(n39880) );
  XNOR U39608 ( .A(p_input[2883]), .B(n39881), .Z(n39065) );
  AND U39609 ( .A(n755), .B(n39882), .Z(n39881) );
  XOR U39610 ( .A(p_input[2915]), .B(p_input[2883]), .Z(n39882) );
  XNOR U39611 ( .A(n39062), .B(n39877), .Z(n39879) );
  XOR U39612 ( .A(n39883), .B(n39884), .Z(n39062) );
  AND U39613 ( .A(n752), .B(n39885), .Z(n39884) );
  XOR U39614 ( .A(p_input[2851]), .B(p_input[2819]), .Z(n39885) );
  XOR U39615 ( .A(n39886), .B(n39887), .Z(n39877) );
  AND U39616 ( .A(n39888), .B(n39889), .Z(n39887) );
  XOR U39617 ( .A(n39886), .B(n39077), .Z(n39889) );
  XNOR U39618 ( .A(p_input[2882]), .B(n39890), .Z(n39077) );
  AND U39619 ( .A(n755), .B(n39891), .Z(n39890) );
  XOR U39620 ( .A(p_input[2914]), .B(p_input[2882]), .Z(n39891) );
  XNOR U39621 ( .A(n39074), .B(n39886), .Z(n39888) );
  XOR U39622 ( .A(n39892), .B(n39893), .Z(n39074) );
  AND U39623 ( .A(n752), .B(n39894), .Z(n39893) );
  XOR U39624 ( .A(p_input[2850]), .B(p_input[2818]), .Z(n39894) );
  XOR U39625 ( .A(n39895), .B(n39896), .Z(n39886) );
  AND U39626 ( .A(n39897), .B(n39898), .Z(n39896) );
  XNOR U39627 ( .A(n39899), .B(n39090), .Z(n39898) );
  XNOR U39628 ( .A(p_input[2881]), .B(n39900), .Z(n39090) );
  AND U39629 ( .A(n755), .B(n39901), .Z(n39900) );
  XNOR U39630 ( .A(p_input[2913]), .B(n39902), .Z(n39901) );
  IV U39631 ( .A(p_input[2881]), .Z(n39902) );
  XNOR U39632 ( .A(n39087), .B(n39895), .Z(n39897) );
  XNOR U39633 ( .A(p_input[2817]), .B(n39903), .Z(n39087) );
  AND U39634 ( .A(n752), .B(n39904), .Z(n39903) );
  XOR U39635 ( .A(p_input[2849]), .B(p_input[2817]), .Z(n39904) );
  IV U39636 ( .A(n39899), .Z(n39895) );
  AND U39637 ( .A(n39625), .B(n39628), .Z(n39899) );
  XOR U39638 ( .A(p_input[2880]), .B(n39905), .Z(n39628) );
  AND U39639 ( .A(n755), .B(n39906), .Z(n39905) );
  XOR U39640 ( .A(p_input[2912]), .B(p_input[2880]), .Z(n39906) );
  XOR U39641 ( .A(n39907), .B(n39908), .Z(n755) );
  AND U39642 ( .A(n39909), .B(n39910), .Z(n39908) );
  XNOR U39643 ( .A(p_input[2943]), .B(n39907), .Z(n39910) );
  XOR U39644 ( .A(n39907), .B(p_input[2911]), .Z(n39909) );
  XOR U39645 ( .A(n39911), .B(n39912), .Z(n39907) );
  AND U39646 ( .A(n39913), .B(n39914), .Z(n39912) );
  XNOR U39647 ( .A(p_input[2942]), .B(n39911), .Z(n39914) );
  XOR U39648 ( .A(n39911), .B(p_input[2910]), .Z(n39913) );
  XOR U39649 ( .A(n39915), .B(n39916), .Z(n39911) );
  AND U39650 ( .A(n39917), .B(n39918), .Z(n39916) );
  XNOR U39651 ( .A(p_input[2941]), .B(n39915), .Z(n39918) );
  XOR U39652 ( .A(n39915), .B(p_input[2909]), .Z(n39917) );
  XOR U39653 ( .A(n39919), .B(n39920), .Z(n39915) );
  AND U39654 ( .A(n39921), .B(n39922), .Z(n39920) );
  XNOR U39655 ( .A(p_input[2940]), .B(n39919), .Z(n39922) );
  XOR U39656 ( .A(n39919), .B(p_input[2908]), .Z(n39921) );
  XOR U39657 ( .A(n39923), .B(n39924), .Z(n39919) );
  AND U39658 ( .A(n39925), .B(n39926), .Z(n39924) );
  XNOR U39659 ( .A(p_input[2939]), .B(n39923), .Z(n39926) );
  XOR U39660 ( .A(n39923), .B(p_input[2907]), .Z(n39925) );
  XOR U39661 ( .A(n39927), .B(n39928), .Z(n39923) );
  AND U39662 ( .A(n39929), .B(n39930), .Z(n39928) );
  XNOR U39663 ( .A(p_input[2938]), .B(n39927), .Z(n39930) );
  XOR U39664 ( .A(n39927), .B(p_input[2906]), .Z(n39929) );
  XOR U39665 ( .A(n39931), .B(n39932), .Z(n39927) );
  AND U39666 ( .A(n39933), .B(n39934), .Z(n39932) );
  XNOR U39667 ( .A(p_input[2937]), .B(n39931), .Z(n39934) );
  XOR U39668 ( .A(n39931), .B(p_input[2905]), .Z(n39933) );
  XOR U39669 ( .A(n39935), .B(n39936), .Z(n39931) );
  AND U39670 ( .A(n39937), .B(n39938), .Z(n39936) );
  XNOR U39671 ( .A(p_input[2936]), .B(n39935), .Z(n39938) );
  XOR U39672 ( .A(n39935), .B(p_input[2904]), .Z(n39937) );
  XOR U39673 ( .A(n39939), .B(n39940), .Z(n39935) );
  AND U39674 ( .A(n39941), .B(n39942), .Z(n39940) );
  XNOR U39675 ( .A(p_input[2935]), .B(n39939), .Z(n39942) );
  XOR U39676 ( .A(n39939), .B(p_input[2903]), .Z(n39941) );
  XOR U39677 ( .A(n39943), .B(n39944), .Z(n39939) );
  AND U39678 ( .A(n39945), .B(n39946), .Z(n39944) );
  XNOR U39679 ( .A(p_input[2934]), .B(n39943), .Z(n39946) );
  XOR U39680 ( .A(n39943), .B(p_input[2902]), .Z(n39945) );
  XOR U39681 ( .A(n39947), .B(n39948), .Z(n39943) );
  AND U39682 ( .A(n39949), .B(n39950), .Z(n39948) );
  XNOR U39683 ( .A(p_input[2933]), .B(n39947), .Z(n39950) );
  XOR U39684 ( .A(n39947), .B(p_input[2901]), .Z(n39949) );
  XOR U39685 ( .A(n39951), .B(n39952), .Z(n39947) );
  AND U39686 ( .A(n39953), .B(n39954), .Z(n39952) );
  XNOR U39687 ( .A(p_input[2932]), .B(n39951), .Z(n39954) );
  XOR U39688 ( .A(n39951), .B(p_input[2900]), .Z(n39953) );
  XOR U39689 ( .A(n39955), .B(n39956), .Z(n39951) );
  AND U39690 ( .A(n39957), .B(n39958), .Z(n39956) );
  XNOR U39691 ( .A(p_input[2931]), .B(n39955), .Z(n39958) );
  XOR U39692 ( .A(n39955), .B(p_input[2899]), .Z(n39957) );
  XOR U39693 ( .A(n39959), .B(n39960), .Z(n39955) );
  AND U39694 ( .A(n39961), .B(n39962), .Z(n39960) );
  XNOR U39695 ( .A(p_input[2930]), .B(n39959), .Z(n39962) );
  XOR U39696 ( .A(n39959), .B(p_input[2898]), .Z(n39961) );
  XOR U39697 ( .A(n39963), .B(n39964), .Z(n39959) );
  AND U39698 ( .A(n39965), .B(n39966), .Z(n39964) );
  XNOR U39699 ( .A(p_input[2929]), .B(n39963), .Z(n39966) );
  XOR U39700 ( .A(n39963), .B(p_input[2897]), .Z(n39965) );
  XOR U39701 ( .A(n39967), .B(n39968), .Z(n39963) );
  AND U39702 ( .A(n39969), .B(n39970), .Z(n39968) );
  XNOR U39703 ( .A(p_input[2928]), .B(n39967), .Z(n39970) );
  XOR U39704 ( .A(n39967), .B(p_input[2896]), .Z(n39969) );
  XOR U39705 ( .A(n39971), .B(n39972), .Z(n39967) );
  AND U39706 ( .A(n39973), .B(n39974), .Z(n39972) );
  XNOR U39707 ( .A(p_input[2927]), .B(n39971), .Z(n39974) );
  XOR U39708 ( .A(n39971), .B(p_input[2895]), .Z(n39973) );
  XOR U39709 ( .A(n39975), .B(n39976), .Z(n39971) );
  AND U39710 ( .A(n39977), .B(n39978), .Z(n39976) );
  XNOR U39711 ( .A(p_input[2926]), .B(n39975), .Z(n39978) );
  XOR U39712 ( .A(n39975), .B(p_input[2894]), .Z(n39977) );
  XOR U39713 ( .A(n39979), .B(n39980), .Z(n39975) );
  AND U39714 ( .A(n39981), .B(n39982), .Z(n39980) );
  XNOR U39715 ( .A(p_input[2925]), .B(n39979), .Z(n39982) );
  XOR U39716 ( .A(n39979), .B(p_input[2893]), .Z(n39981) );
  XOR U39717 ( .A(n39983), .B(n39984), .Z(n39979) );
  AND U39718 ( .A(n39985), .B(n39986), .Z(n39984) );
  XNOR U39719 ( .A(p_input[2924]), .B(n39983), .Z(n39986) );
  XOR U39720 ( .A(n39983), .B(p_input[2892]), .Z(n39985) );
  XOR U39721 ( .A(n39987), .B(n39988), .Z(n39983) );
  AND U39722 ( .A(n39989), .B(n39990), .Z(n39988) );
  XNOR U39723 ( .A(p_input[2923]), .B(n39987), .Z(n39990) );
  XOR U39724 ( .A(n39987), .B(p_input[2891]), .Z(n39989) );
  XOR U39725 ( .A(n39991), .B(n39992), .Z(n39987) );
  AND U39726 ( .A(n39993), .B(n39994), .Z(n39992) );
  XNOR U39727 ( .A(p_input[2922]), .B(n39991), .Z(n39994) );
  XOR U39728 ( .A(n39991), .B(p_input[2890]), .Z(n39993) );
  XOR U39729 ( .A(n39995), .B(n39996), .Z(n39991) );
  AND U39730 ( .A(n39997), .B(n39998), .Z(n39996) );
  XNOR U39731 ( .A(p_input[2921]), .B(n39995), .Z(n39998) );
  XOR U39732 ( .A(n39995), .B(p_input[2889]), .Z(n39997) );
  XOR U39733 ( .A(n39999), .B(n40000), .Z(n39995) );
  AND U39734 ( .A(n40001), .B(n40002), .Z(n40000) );
  XNOR U39735 ( .A(p_input[2920]), .B(n39999), .Z(n40002) );
  XOR U39736 ( .A(n39999), .B(p_input[2888]), .Z(n40001) );
  XOR U39737 ( .A(n40003), .B(n40004), .Z(n39999) );
  AND U39738 ( .A(n40005), .B(n40006), .Z(n40004) );
  XNOR U39739 ( .A(p_input[2919]), .B(n40003), .Z(n40006) );
  XOR U39740 ( .A(n40003), .B(p_input[2887]), .Z(n40005) );
  XOR U39741 ( .A(n40007), .B(n40008), .Z(n40003) );
  AND U39742 ( .A(n40009), .B(n40010), .Z(n40008) );
  XNOR U39743 ( .A(p_input[2918]), .B(n40007), .Z(n40010) );
  XOR U39744 ( .A(n40007), .B(p_input[2886]), .Z(n40009) );
  XOR U39745 ( .A(n40011), .B(n40012), .Z(n40007) );
  AND U39746 ( .A(n40013), .B(n40014), .Z(n40012) );
  XNOR U39747 ( .A(p_input[2917]), .B(n40011), .Z(n40014) );
  XOR U39748 ( .A(n40011), .B(p_input[2885]), .Z(n40013) );
  XOR U39749 ( .A(n40015), .B(n40016), .Z(n40011) );
  AND U39750 ( .A(n40017), .B(n40018), .Z(n40016) );
  XNOR U39751 ( .A(p_input[2916]), .B(n40015), .Z(n40018) );
  XOR U39752 ( .A(n40015), .B(p_input[2884]), .Z(n40017) );
  XOR U39753 ( .A(n40019), .B(n40020), .Z(n40015) );
  AND U39754 ( .A(n40021), .B(n40022), .Z(n40020) );
  XNOR U39755 ( .A(p_input[2915]), .B(n40019), .Z(n40022) );
  XOR U39756 ( .A(n40019), .B(p_input[2883]), .Z(n40021) );
  XOR U39757 ( .A(n40023), .B(n40024), .Z(n40019) );
  AND U39758 ( .A(n40025), .B(n40026), .Z(n40024) );
  XNOR U39759 ( .A(p_input[2914]), .B(n40023), .Z(n40026) );
  XOR U39760 ( .A(n40023), .B(p_input[2882]), .Z(n40025) );
  XNOR U39761 ( .A(n40027), .B(n40028), .Z(n40023) );
  AND U39762 ( .A(n40029), .B(n40030), .Z(n40028) );
  XOR U39763 ( .A(p_input[2913]), .B(n40027), .Z(n40030) );
  XNOR U39764 ( .A(p_input[2881]), .B(n40027), .Z(n40029) );
  AND U39765 ( .A(p_input[2912]), .B(n40031), .Z(n40027) );
  IV U39766 ( .A(p_input[2880]), .Z(n40031) );
  XNOR U39767 ( .A(p_input[2816]), .B(n40032), .Z(n39625) );
  AND U39768 ( .A(n752), .B(n40033), .Z(n40032) );
  XOR U39769 ( .A(p_input[2848]), .B(p_input[2816]), .Z(n40033) );
  XOR U39770 ( .A(n40034), .B(n40035), .Z(n752) );
  AND U39771 ( .A(n40036), .B(n40037), .Z(n40035) );
  XNOR U39772 ( .A(p_input[2879]), .B(n40034), .Z(n40037) );
  XOR U39773 ( .A(n40034), .B(p_input[2847]), .Z(n40036) );
  XOR U39774 ( .A(n40038), .B(n40039), .Z(n40034) );
  AND U39775 ( .A(n40040), .B(n40041), .Z(n40039) );
  XNOR U39776 ( .A(p_input[2878]), .B(n40038), .Z(n40041) );
  XNOR U39777 ( .A(n40038), .B(n39640), .Z(n40040) );
  IV U39778 ( .A(p_input[2846]), .Z(n39640) );
  XOR U39779 ( .A(n40042), .B(n40043), .Z(n40038) );
  AND U39780 ( .A(n40044), .B(n40045), .Z(n40043) );
  XNOR U39781 ( .A(p_input[2877]), .B(n40042), .Z(n40045) );
  XNOR U39782 ( .A(n40042), .B(n39649), .Z(n40044) );
  IV U39783 ( .A(p_input[2845]), .Z(n39649) );
  XOR U39784 ( .A(n40046), .B(n40047), .Z(n40042) );
  AND U39785 ( .A(n40048), .B(n40049), .Z(n40047) );
  XNOR U39786 ( .A(p_input[2876]), .B(n40046), .Z(n40049) );
  XNOR U39787 ( .A(n40046), .B(n39658), .Z(n40048) );
  IV U39788 ( .A(p_input[2844]), .Z(n39658) );
  XOR U39789 ( .A(n40050), .B(n40051), .Z(n40046) );
  AND U39790 ( .A(n40052), .B(n40053), .Z(n40051) );
  XNOR U39791 ( .A(p_input[2875]), .B(n40050), .Z(n40053) );
  XNOR U39792 ( .A(n40050), .B(n39667), .Z(n40052) );
  IV U39793 ( .A(p_input[2843]), .Z(n39667) );
  XOR U39794 ( .A(n40054), .B(n40055), .Z(n40050) );
  AND U39795 ( .A(n40056), .B(n40057), .Z(n40055) );
  XNOR U39796 ( .A(p_input[2874]), .B(n40054), .Z(n40057) );
  XNOR U39797 ( .A(n40054), .B(n39676), .Z(n40056) );
  IV U39798 ( .A(p_input[2842]), .Z(n39676) );
  XOR U39799 ( .A(n40058), .B(n40059), .Z(n40054) );
  AND U39800 ( .A(n40060), .B(n40061), .Z(n40059) );
  XNOR U39801 ( .A(p_input[2873]), .B(n40058), .Z(n40061) );
  XNOR U39802 ( .A(n40058), .B(n39685), .Z(n40060) );
  IV U39803 ( .A(p_input[2841]), .Z(n39685) );
  XOR U39804 ( .A(n40062), .B(n40063), .Z(n40058) );
  AND U39805 ( .A(n40064), .B(n40065), .Z(n40063) );
  XNOR U39806 ( .A(p_input[2872]), .B(n40062), .Z(n40065) );
  XNOR U39807 ( .A(n40062), .B(n39694), .Z(n40064) );
  IV U39808 ( .A(p_input[2840]), .Z(n39694) );
  XOR U39809 ( .A(n40066), .B(n40067), .Z(n40062) );
  AND U39810 ( .A(n40068), .B(n40069), .Z(n40067) );
  XNOR U39811 ( .A(p_input[2871]), .B(n40066), .Z(n40069) );
  XNOR U39812 ( .A(n40066), .B(n39703), .Z(n40068) );
  IV U39813 ( .A(p_input[2839]), .Z(n39703) );
  XOR U39814 ( .A(n40070), .B(n40071), .Z(n40066) );
  AND U39815 ( .A(n40072), .B(n40073), .Z(n40071) );
  XNOR U39816 ( .A(p_input[2870]), .B(n40070), .Z(n40073) );
  XNOR U39817 ( .A(n40070), .B(n39712), .Z(n40072) );
  IV U39818 ( .A(p_input[2838]), .Z(n39712) );
  XOR U39819 ( .A(n40074), .B(n40075), .Z(n40070) );
  AND U39820 ( .A(n40076), .B(n40077), .Z(n40075) );
  XNOR U39821 ( .A(p_input[2869]), .B(n40074), .Z(n40077) );
  XNOR U39822 ( .A(n40074), .B(n39721), .Z(n40076) );
  IV U39823 ( .A(p_input[2837]), .Z(n39721) );
  XOR U39824 ( .A(n40078), .B(n40079), .Z(n40074) );
  AND U39825 ( .A(n40080), .B(n40081), .Z(n40079) );
  XNOR U39826 ( .A(p_input[2868]), .B(n40078), .Z(n40081) );
  XNOR U39827 ( .A(n40078), .B(n39730), .Z(n40080) );
  IV U39828 ( .A(p_input[2836]), .Z(n39730) );
  XOR U39829 ( .A(n40082), .B(n40083), .Z(n40078) );
  AND U39830 ( .A(n40084), .B(n40085), .Z(n40083) );
  XNOR U39831 ( .A(p_input[2867]), .B(n40082), .Z(n40085) );
  XNOR U39832 ( .A(n40082), .B(n39739), .Z(n40084) );
  IV U39833 ( .A(p_input[2835]), .Z(n39739) );
  XOR U39834 ( .A(n40086), .B(n40087), .Z(n40082) );
  AND U39835 ( .A(n40088), .B(n40089), .Z(n40087) );
  XNOR U39836 ( .A(p_input[2866]), .B(n40086), .Z(n40089) );
  XNOR U39837 ( .A(n40086), .B(n39748), .Z(n40088) );
  IV U39838 ( .A(p_input[2834]), .Z(n39748) );
  XOR U39839 ( .A(n40090), .B(n40091), .Z(n40086) );
  AND U39840 ( .A(n40092), .B(n40093), .Z(n40091) );
  XNOR U39841 ( .A(p_input[2865]), .B(n40090), .Z(n40093) );
  XNOR U39842 ( .A(n40090), .B(n39757), .Z(n40092) );
  IV U39843 ( .A(p_input[2833]), .Z(n39757) );
  XOR U39844 ( .A(n40094), .B(n40095), .Z(n40090) );
  AND U39845 ( .A(n40096), .B(n40097), .Z(n40095) );
  XNOR U39846 ( .A(p_input[2864]), .B(n40094), .Z(n40097) );
  XNOR U39847 ( .A(n40094), .B(n39766), .Z(n40096) );
  IV U39848 ( .A(p_input[2832]), .Z(n39766) );
  XOR U39849 ( .A(n40098), .B(n40099), .Z(n40094) );
  AND U39850 ( .A(n40100), .B(n40101), .Z(n40099) );
  XNOR U39851 ( .A(p_input[2863]), .B(n40098), .Z(n40101) );
  XNOR U39852 ( .A(n40098), .B(n39775), .Z(n40100) );
  IV U39853 ( .A(p_input[2831]), .Z(n39775) );
  XOR U39854 ( .A(n40102), .B(n40103), .Z(n40098) );
  AND U39855 ( .A(n40104), .B(n40105), .Z(n40103) );
  XNOR U39856 ( .A(p_input[2862]), .B(n40102), .Z(n40105) );
  XNOR U39857 ( .A(n40102), .B(n39784), .Z(n40104) );
  IV U39858 ( .A(p_input[2830]), .Z(n39784) );
  XOR U39859 ( .A(n40106), .B(n40107), .Z(n40102) );
  AND U39860 ( .A(n40108), .B(n40109), .Z(n40107) );
  XNOR U39861 ( .A(p_input[2861]), .B(n40106), .Z(n40109) );
  XNOR U39862 ( .A(n40106), .B(n39793), .Z(n40108) );
  IV U39863 ( .A(p_input[2829]), .Z(n39793) );
  XOR U39864 ( .A(n40110), .B(n40111), .Z(n40106) );
  AND U39865 ( .A(n40112), .B(n40113), .Z(n40111) );
  XNOR U39866 ( .A(p_input[2860]), .B(n40110), .Z(n40113) );
  XNOR U39867 ( .A(n40110), .B(n39802), .Z(n40112) );
  IV U39868 ( .A(p_input[2828]), .Z(n39802) );
  XOR U39869 ( .A(n40114), .B(n40115), .Z(n40110) );
  AND U39870 ( .A(n40116), .B(n40117), .Z(n40115) );
  XNOR U39871 ( .A(p_input[2859]), .B(n40114), .Z(n40117) );
  XNOR U39872 ( .A(n40114), .B(n39811), .Z(n40116) );
  IV U39873 ( .A(p_input[2827]), .Z(n39811) );
  XOR U39874 ( .A(n40118), .B(n40119), .Z(n40114) );
  AND U39875 ( .A(n40120), .B(n40121), .Z(n40119) );
  XNOR U39876 ( .A(p_input[2858]), .B(n40118), .Z(n40121) );
  XNOR U39877 ( .A(n40118), .B(n39820), .Z(n40120) );
  IV U39878 ( .A(p_input[2826]), .Z(n39820) );
  XOR U39879 ( .A(n40122), .B(n40123), .Z(n40118) );
  AND U39880 ( .A(n40124), .B(n40125), .Z(n40123) );
  XNOR U39881 ( .A(p_input[2857]), .B(n40122), .Z(n40125) );
  XNOR U39882 ( .A(n40122), .B(n39829), .Z(n40124) );
  IV U39883 ( .A(p_input[2825]), .Z(n39829) );
  XOR U39884 ( .A(n40126), .B(n40127), .Z(n40122) );
  AND U39885 ( .A(n40128), .B(n40129), .Z(n40127) );
  XNOR U39886 ( .A(p_input[2856]), .B(n40126), .Z(n40129) );
  XNOR U39887 ( .A(n40126), .B(n39838), .Z(n40128) );
  IV U39888 ( .A(p_input[2824]), .Z(n39838) );
  XOR U39889 ( .A(n40130), .B(n40131), .Z(n40126) );
  AND U39890 ( .A(n40132), .B(n40133), .Z(n40131) );
  XNOR U39891 ( .A(p_input[2855]), .B(n40130), .Z(n40133) );
  XNOR U39892 ( .A(n40130), .B(n39847), .Z(n40132) );
  IV U39893 ( .A(p_input[2823]), .Z(n39847) );
  XOR U39894 ( .A(n40134), .B(n40135), .Z(n40130) );
  AND U39895 ( .A(n40136), .B(n40137), .Z(n40135) );
  XNOR U39896 ( .A(p_input[2854]), .B(n40134), .Z(n40137) );
  XNOR U39897 ( .A(n40134), .B(n39856), .Z(n40136) );
  IV U39898 ( .A(p_input[2822]), .Z(n39856) );
  XOR U39899 ( .A(n40138), .B(n40139), .Z(n40134) );
  AND U39900 ( .A(n40140), .B(n40141), .Z(n40139) );
  XNOR U39901 ( .A(p_input[2853]), .B(n40138), .Z(n40141) );
  XNOR U39902 ( .A(n40138), .B(n39865), .Z(n40140) );
  IV U39903 ( .A(p_input[2821]), .Z(n39865) );
  XOR U39904 ( .A(n40142), .B(n40143), .Z(n40138) );
  AND U39905 ( .A(n40144), .B(n40145), .Z(n40143) );
  XNOR U39906 ( .A(p_input[2852]), .B(n40142), .Z(n40145) );
  XNOR U39907 ( .A(n40142), .B(n39874), .Z(n40144) );
  IV U39908 ( .A(p_input[2820]), .Z(n39874) );
  XOR U39909 ( .A(n40146), .B(n40147), .Z(n40142) );
  AND U39910 ( .A(n40148), .B(n40149), .Z(n40147) );
  XNOR U39911 ( .A(p_input[2851]), .B(n40146), .Z(n40149) );
  XNOR U39912 ( .A(n40146), .B(n39883), .Z(n40148) );
  IV U39913 ( .A(p_input[2819]), .Z(n39883) );
  XOR U39914 ( .A(n40150), .B(n40151), .Z(n40146) );
  AND U39915 ( .A(n40152), .B(n40153), .Z(n40151) );
  XNOR U39916 ( .A(p_input[2850]), .B(n40150), .Z(n40153) );
  XNOR U39917 ( .A(n40150), .B(n39892), .Z(n40152) );
  IV U39918 ( .A(p_input[2818]), .Z(n39892) );
  XNOR U39919 ( .A(n40154), .B(n40155), .Z(n40150) );
  AND U39920 ( .A(n40156), .B(n40157), .Z(n40155) );
  XOR U39921 ( .A(p_input[2849]), .B(n40154), .Z(n40157) );
  XNOR U39922 ( .A(p_input[2817]), .B(n40154), .Z(n40156) );
  AND U39923 ( .A(p_input[2848]), .B(n40158), .Z(n40154) );
  IV U39924 ( .A(p_input[2816]), .Z(n40158) );
  XOR U39925 ( .A(n40159), .B(n40160), .Z(n38337) );
  AND U39926 ( .A(n885), .B(n40161), .Z(n40160) );
  XNOR U39927 ( .A(n40162), .B(n40159), .Z(n40161) );
  XOR U39928 ( .A(n40163), .B(n40164), .Z(n885) );
  AND U39929 ( .A(n40165), .B(n40166), .Z(n40164) );
  XOR U39930 ( .A(n40163), .B(n38352), .Z(n40166) );
  XNOR U39931 ( .A(n40167), .B(n40168), .Z(n38352) );
  AND U39932 ( .A(n40169), .B(n595), .Z(n40168) );
  AND U39933 ( .A(n40167), .B(n40170), .Z(n40169) );
  XNOR U39934 ( .A(n38349), .B(n40163), .Z(n40165) );
  XOR U39935 ( .A(n40171), .B(n40172), .Z(n38349) );
  AND U39936 ( .A(n40173), .B(n592), .Z(n40172) );
  NOR U39937 ( .A(n40171), .B(n40174), .Z(n40173) );
  XOR U39938 ( .A(n40175), .B(n40176), .Z(n40163) );
  AND U39939 ( .A(n40177), .B(n40178), .Z(n40176) );
  XOR U39940 ( .A(n40175), .B(n38364), .Z(n40178) );
  XOR U39941 ( .A(n40179), .B(n40180), .Z(n38364) );
  AND U39942 ( .A(n595), .B(n40181), .Z(n40180) );
  XOR U39943 ( .A(n40182), .B(n40179), .Z(n40181) );
  XNOR U39944 ( .A(n38361), .B(n40175), .Z(n40177) );
  XOR U39945 ( .A(n40183), .B(n40184), .Z(n38361) );
  AND U39946 ( .A(n592), .B(n40185), .Z(n40184) );
  XOR U39947 ( .A(n40186), .B(n40183), .Z(n40185) );
  XOR U39948 ( .A(n40187), .B(n40188), .Z(n40175) );
  AND U39949 ( .A(n40189), .B(n40190), .Z(n40188) );
  XOR U39950 ( .A(n40187), .B(n38376), .Z(n40190) );
  XOR U39951 ( .A(n40191), .B(n40192), .Z(n38376) );
  AND U39952 ( .A(n595), .B(n40193), .Z(n40192) );
  XOR U39953 ( .A(n40194), .B(n40191), .Z(n40193) );
  XNOR U39954 ( .A(n38373), .B(n40187), .Z(n40189) );
  XOR U39955 ( .A(n40195), .B(n40196), .Z(n38373) );
  AND U39956 ( .A(n592), .B(n40197), .Z(n40196) );
  XOR U39957 ( .A(n40198), .B(n40195), .Z(n40197) );
  XOR U39958 ( .A(n40199), .B(n40200), .Z(n40187) );
  AND U39959 ( .A(n40201), .B(n40202), .Z(n40200) );
  XOR U39960 ( .A(n40199), .B(n38388), .Z(n40202) );
  XOR U39961 ( .A(n40203), .B(n40204), .Z(n38388) );
  AND U39962 ( .A(n595), .B(n40205), .Z(n40204) );
  XOR U39963 ( .A(n40206), .B(n40203), .Z(n40205) );
  XNOR U39964 ( .A(n38385), .B(n40199), .Z(n40201) );
  XOR U39965 ( .A(n40207), .B(n40208), .Z(n38385) );
  AND U39966 ( .A(n592), .B(n40209), .Z(n40208) );
  XOR U39967 ( .A(n40210), .B(n40207), .Z(n40209) );
  XOR U39968 ( .A(n40211), .B(n40212), .Z(n40199) );
  AND U39969 ( .A(n40213), .B(n40214), .Z(n40212) );
  XOR U39970 ( .A(n40211), .B(n38400), .Z(n40214) );
  XOR U39971 ( .A(n40215), .B(n40216), .Z(n38400) );
  AND U39972 ( .A(n595), .B(n40217), .Z(n40216) );
  XOR U39973 ( .A(n40218), .B(n40215), .Z(n40217) );
  XNOR U39974 ( .A(n38397), .B(n40211), .Z(n40213) );
  XOR U39975 ( .A(n40219), .B(n40220), .Z(n38397) );
  AND U39976 ( .A(n592), .B(n40221), .Z(n40220) );
  XOR U39977 ( .A(n40222), .B(n40219), .Z(n40221) );
  XOR U39978 ( .A(n40223), .B(n40224), .Z(n40211) );
  AND U39979 ( .A(n40225), .B(n40226), .Z(n40224) );
  XOR U39980 ( .A(n40223), .B(n38412), .Z(n40226) );
  XOR U39981 ( .A(n40227), .B(n40228), .Z(n38412) );
  AND U39982 ( .A(n595), .B(n40229), .Z(n40228) );
  XOR U39983 ( .A(n40230), .B(n40227), .Z(n40229) );
  XNOR U39984 ( .A(n38409), .B(n40223), .Z(n40225) );
  XOR U39985 ( .A(n40231), .B(n40232), .Z(n38409) );
  AND U39986 ( .A(n592), .B(n40233), .Z(n40232) );
  XOR U39987 ( .A(n40234), .B(n40231), .Z(n40233) );
  XOR U39988 ( .A(n40235), .B(n40236), .Z(n40223) );
  AND U39989 ( .A(n40237), .B(n40238), .Z(n40236) );
  XOR U39990 ( .A(n40235), .B(n38424), .Z(n40238) );
  XOR U39991 ( .A(n40239), .B(n40240), .Z(n38424) );
  AND U39992 ( .A(n595), .B(n40241), .Z(n40240) );
  XOR U39993 ( .A(n40242), .B(n40239), .Z(n40241) );
  XNOR U39994 ( .A(n38421), .B(n40235), .Z(n40237) );
  XOR U39995 ( .A(n40243), .B(n40244), .Z(n38421) );
  AND U39996 ( .A(n592), .B(n40245), .Z(n40244) );
  XOR U39997 ( .A(n40246), .B(n40243), .Z(n40245) );
  XOR U39998 ( .A(n40247), .B(n40248), .Z(n40235) );
  AND U39999 ( .A(n40249), .B(n40250), .Z(n40248) );
  XOR U40000 ( .A(n40247), .B(n38436), .Z(n40250) );
  XOR U40001 ( .A(n40251), .B(n40252), .Z(n38436) );
  AND U40002 ( .A(n595), .B(n40253), .Z(n40252) );
  XOR U40003 ( .A(n40254), .B(n40251), .Z(n40253) );
  XNOR U40004 ( .A(n38433), .B(n40247), .Z(n40249) );
  XOR U40005 ( .A(n40255), .B(n40256), .Z(n38433) );
  AND U40006 ( .A(n592), .B(n40257), .Z(n40256) );
  XOR U40007 ( .A(n40258), .B(n40255), .Z(n40257) );
  XOR U40008 ( .A(n40259), .B(n40260), .Z(n40247) );
  AND U40009 ( .A(n40261), .B(n40262), .Z(n40260) );
  XOR U40010 ( .A(n40259), .B(n38448), .Z(n40262) );
  XOR U40011 ( .A(n40263), .B(n40264), .Z(n38448) );
  AND U40012 ( .A(n595), .B(n40265), .Z(n40264) );
  XOR U40013 ( .A(n40266), .B(n40263), .Z(n40265) );
  XNOR U40014 ( .A(n38445), .B(n40259), .Z(n40261) );
  XOR U40015 ( .A(n40267), .B(n40268), .Z(n38445) );
  AND U40016 ( .A(n592), .B(n40269), .Z(n40268) );
  XOR U40017 ( .A(n40270), .B(n40267), .Z(n40269) );
  XOR U40018 ( .A(n40271), .B(n40272), .Z(n40259) );
  AND U40019 ( .A(n40273), .B(n40274), .Z(n40272) );
  XOR U40020 ( .A(n40271), .B(n38460), .Z(n40274) );
  XOR U40021 ( .A(n40275), .B(n40276), .Z(n38460) );
  AND U40022 ( .A(n595), .B(n40277), .Z(n40276) );
  XOR U40023 ( .A(n40278), .B(n40275), .Z(n40277) );
  XNOR U40024 ( .A(n38457), .B(n40271), .Z(n40273) );
  XOR U40025 ( .A(n40279), .B(n40280), .Z(n38457) );
  AND U40026 ( .A(n592), .B(n40281), .Z(n40280) );
  XOR U40027 ( .A(n40282), .B(n40279), .Z(n40281) );
  XOR U40028 ( .A(n40283), .B(n40284), .Z(n40271) );
  AND U40029 ( .A(n40285), .B(n40286), .Z(n40284) );
  XOR U40030 ( .A(n40283), .B(n38472), .Z(n40286) );
  XOR U40031 ( .A(n40287), .B(n40288), .Z(n38472) );
  AND U40032 ( .A(n595), .B(n40289), .Z(n40288) );
  XOR U40033 ( .A(n40290), .B(n40287), .Z(n40289) );
  XNOR U40034 ( .A(n38469), .B(n40283), .Z(n40285) );
  XOR U40035 ( .A(n40291), .B(n40292), .Z(n38469) );
  AND U40036 ( .A(n592), .B(n40293), .Z(n40292) );
  XOR U40037 ( .A(n40294), .B(n40291), .Z(n40293) );
  XOR U40038 ( .A(n40295), .B(n40296), .Z(n40283) );
  AND U40039 ( .A(n40297), .B(n40298), .Z(n40296) );
  XOR U40040 ( .A(n40295), .B(n38484), .Z(n40298) );
  XOR U40041 ( .A(n40299), .B(n40300), .Z(n38484) );
  AND U40042 ( .A(n595), .B(n40301), .Z(n40300) );
  XOR U40043 ( .A(n40302), .B(n40299), .Z(n40301) );
  XNOR U40044 ( .A(n38481), .B(n40295), .Z(n40297) );
  XOR U40045 ( .A(n40303), .B(n40304), .Z(n38481) );
  AND U40046 ( .A(n592), .B(n40305), .Z(n40304) );
  XOR U40047 ( .A(n40306), .B(n40303), .Z(n40305) );
  XOR U40048 ( .A(n40307), .B(n40308), .Z(n40295) );
  AND U40049 ( .A(n40309), .B(n40310), .Z(n40308) );
  XOR U40050 ( .A(n40307), .B(n38496), .Z(n40310) );
  XOR U40051 ( .A(n40311), .B(n40312), .Z(n38496) );
  AND U40052 ( .A(n595), .B(n40313), .Z(n40312) );
  XOR U40053 ( .A(n40314), .B(n40311), .Z(n40313) );
  XNOR U40054 ( .A(n38493), .B(n40307), .Z(n40309) );
  XOR U40055 ( .A(n40315), .B(n40316), .Z(n38493) );
  AND U40056 ( .A(n592), .B(n40317), .Z(n40316) );
  XOR U40057 ( .A(n40318), .B(n40315), .Z(n40317) );
  XOR U40058 ( .A(n40319), .B(n40320), .Z(n40307) );
  AND U40059 ( .A(n40321), .B(n40322), .Z(n40320) );
  XOR U40060 ( .A(n40319), .B(n38508), .Z(n40322) );
  XOR U40061 ( .A(n40323), .B(n40324), .Z(n38508) );
  AND U40062 ( .A(n595), .B(n40325), .Z(n40324) );
  XOR U40063 ( .A(n40326), .B(n40323), .Z(n40325) );
  XNOR U40064 ( .A(n38505), .B(n40319), .Z(n40321) );
  XOR U40065 ( .A(n40327), .B(n40328), .Z(n38505) );
  AND U40066 ( .A(n592), .B(n40329), .Z(n40328) );
  XOR U40067 ( .A(n40330), .B(n40327), .Z(n40329) );
  XOR U40068 ( .A(n40331), .B(n40332), .Z(n40319) );
  AND U40069 ( .A(n40333), .B(n40334), .Z(n40332) );
  XOR U40070 ( .A(n40331), .B(n38520), .Z(n40334) );
  XOR U40071 ( .A(n40335), .B(n40336), .Z(n38520) );
  AND U40072 ( .A(n595), .B(n40337), .Z(n40336) );
  XOR U40073 ( .A(n40338), .B(n40335), .Z(n40337) );
  XNOR U40074 ( .A(n38517), .B(n40331), .Z(n40333) );
  XOR U40075 ( .A(n40339), .B(n40340), .Z(n38517) );
  AND U40076 ( .A(n592), .B(n40341), .Z(n40340) );
  XOR U40077 ( .A(n40342), .B(n40339), .Z(n40341) );
  XOR U40078 ( .A(n40343), .B(n40344), .Z(n40331) );
  AND U40079 ( .A(n40345), .B(n40346), .Z(n40344) );
  XOR U40080 ( .A(n40343), .B(n38532), .Z(n40346) );
  XOR U40081 ( .A(n40347), .B(n40348), .Z(n38532) );
  AND U40082 ( .A(n595), .B(n40349), .Z(n40348) );
  XOR U40083 ( .A(n40350), .B(n40347), .Z(n40349) );
  XNOR U40084 ( .A(n38529), .B(n40343), .Z(n40345) );
  XOR U40085 ( .A(n40351), .B(n40352), .Z(n38529) );
  AND U40086 ( .A(n592), .B(n40353), .Z(n40352) );
  XOR U40087 ( .A(n40354), .B(n40351), .Z(n40353) );
  XOR U40088 ( .A(n40355), .B(n40356), .Z(n40343) );
  AND U40089 ( .A(n40357), .B(n40358), .Z(n40356) );
  XOR U40090 ( .A(n40355), .B(n38544), .Z(n40358) );
  XOR U40091 ( .A(n40359), .B(n40360), .Z(n38544) );
  AND U40092 ( .A(n595), .B(n40361), .Z(n40360) );
  XOR U40093 ( .A(n40362), .B(n40359), .Z(n40361) );
  XNOR U40094 ( .A(n38541), .B(n40355), .Z(n40357) );
  XOR U40095 ( .A(n40363), .B(n40364), .Z(n38541) );
  AND U40096 ( .A(n592), .B(n40365), .Z(n40364) );
  XOR U40097 ( .A(n40366), .B(n40363), .Z(n40365) );
  XOR U40098 ( .A(n40367), .B(n40368), .Z(n40355) );
  AND U40099 ( .A(n40369), .B(n40370), .Z(n40368) );
  XOR U40100 ( .A(n40367), .B(n38556), .Z(n40370) );
  XOR U40101 ( .A(n40371), .B(n40372), .Z(n38556) );
  AND U40102 ( .A(n595), .B(n40373), .Z(n40372) );
  XOR U40103 ( .A(n40374), .B(n40371), .Z(n40373) );
  XNOR U40104 ( .A(n38553), .B(n40367), .Z(n40369) );
  XOR U40105 ( .A(n40375), .B(n40376), .Z(n38553) );
  AND U40106 ( .A(n592), .B(n40377), .Z(n40376) );
  XOR U40107 ( .A(n40378), .B(n40375), .Z(n40377) );
  XOR U40108 ( .A(n40379), .B(n40380), .Z(n40367) );
  AND U40109 ( .A(n40381), .B(n40382), .Z(n40380) );
  XOR U40110 ( .A(n40379), .B(n38568), .Z(n40382) );
  XOR U40111 ( .A(n40383), .B(n40384), .Z(n38568) );
  AND U40112 ( .A(n595), .B(n40385), .Z(n40384) );
  XOR U40113 ( .A(n40386), .B(n40383), .Z(n40385) );
  XNOR U40114 ( .A(n38565), .B(n40379), .Z(n40381) );
  XOR U40115 ( .A(n40387), .B(n40388), .Z(n38565) );
  AND U40116 ( .A(n592), .B(n40389), .Z(n40388) );
  XOR U40117 ( .A(n40390), .B(n40387), .Z(n40389) );
  XOR U40118 ( .A(n40391), .B(n40392), .Z(n40379) );
  AND U40119 ( .A(n40393), .B(n40394), .Z(n40392) );
  XOR U40120 ( .A(n40391), .B(n38580), .Z(n40394) );
  XOR U40121 ( .A(n40395), .B(n40396), .Z(n38580) );
  AND U40122 ( .A(n595), .B(n40397), .Z(n40396) );
  XOR U40123 ( .A(n40398), .B(n40395), .Z(n40397) );
  XNOR U40124 ( .A(n38577), .B(n40391), .Z(n40393) );
  XOR U40125 ( .A(n40399), .B(n40400), .Z(n38577) );
  AND U40126 ( .A(n592), .B(n40401), .Z(n40400) );
  XOR U40127 ( .A(n40402), .B(n40399), .Z(n40401) );
  XOR U40128 ( .A(n40403), .B(n40404), .Z(n40391) );
  AND U40129 ( .A(n40405), .B(n40406), .Z(n40404) );
  XOR U40130 ( .A(n40403), .B(n38592), .Z(n40406) );
  XOR U40131 ( .A(n40407), .B(n40408), .Z(n38592) );
  AND U40132 ( .A(n595), .B(n40409), .Z(n40408) );
  XOR U40133 ( .A(n40410), .B(n40407), .Z(n40409) );
  XNOR U40134 ( .A(n38589), .B(n40403), .Z(n40405) );
  XOR U40135 ( .A(n40411), .B(n40412), .Z(n38589) );
  AND U40136 ( .A(n592), .B(n40413), .Z(n40412) );
  XOR U40137 ( .A(n40414), .B(n40411), .Z(n40413) );
  XOR U40138 ( .A(n40415), .B(n40416), .Z(n40403) );
  AND U40139 ( .A(n40417), .B(n40418), .Z(n40416) );
  XOR U40140 ( .A(n40415), .B(n38604), .Z(n40418) );
  XOR U40141 ( .A(n40419), .B(n40420), .Z(n38604) );
  AND U40142 ( .A(n595), .B(n40421), .Z(n40420) );
  XOR U40143 ( .A(n40422), .B(n40419), .Z(n40421) );
  XNOR U40144 ( .A(n38601), .B(n40415), .Z(n40417) );
  XOR U40145 ( .A(n40423), .B(n40424), .Z(n38601) );
  AND U40146 ( .A(n592), .B(n40425), .Z(n40424) );
  XOR U40147 ( .A(n40426), .B(n40423), .Z(n40425) );
  XOR U40148 ( .A(n40427), .B(n40428), .Z(n40415) );
  AND U40149 ( .A(n40429), .B(n40430), .Z(n40428) );
  XOR U40150 ( .A(n40427), .B(n38616), .Z(n40430) );
  XOR U40151 ( .A(n40431), .B(n40432), .Z(n38616) );
  AND U40152 ( .A(n595), .B(n40433), .Z(n40432) );
  XOR U40153 ( .A(n40434), .B(n40431), .Z(n40433) );
  XNOR U40154 ( .A(n38613), .B(n40427), .Z(n40429) );
  XOR U40155 ( .A(n40435), .B(n40436), .Z(n38613) );
  AND U40156 ( .A(n592), .B(n40437), .Z(n40436) );
  XOR U40157 ( .A(n40438), .B(n40435), .Z(n40437) );
  XOR U40158 ( .A(n40439), .B(n40440), .Z(n40427) );
  AND U40159 ( .A(n40441), .B(n40442), .Z(n40440) );
  XOR U40160 ( .A(n40439), .B(n38628), .Z(n40442) );
  XOR U40161 ( .A(n40443), .B(n40444), .Z(n38628) );
  AND U40162 ( .A(n595), .B(n40445), .Z(n40444) );
  XOR U40163 ( .A(n40446), .B(n40443), .Z(n40445) );
  XNOR U40164 ( .A(n38625), .B(n40439), .Z(n40441) );
  XOR U40165 ( .A(n40447), .B(n40448), .Z(n38625) );
  AND U40166 ( .A(n592), .B(n40449), .Z(n40448) );
  XOR U40167 ( .A(n40450), .B(n40447), .Z(n40449) );
  XOR U40168 ( .A(n40451), .B(n40452), .Z(n40439) );
  AND U40169 ( .A(n40453), .B(n40454), .Z(n40452) );
  XOR U40170 ( .A(n40451), .B(n38640), .Z(n40454) );
  XOR U40171 ( .A(n40455), .B(n40456), .Z(n38640) );
  AND U40172 ( .A(n595), .B(n40457), .Z(n40456) );
  XOR U40173 ( .A(n40458), .B(n40455), .Z(n40457) );
  XNOR U40174 ( .A(n38637), .B(n40451), .Z(n40453) );
  XOR U40175 ( .A(n40459), .B(n40460), .Z(n38637) );
  AND U40176 ( .A(n592), .B(n40461), .Z(n40460) );
  XOR U40177 ( .A(n40462), .B(n40459), .Z(n40461) );
  XOR U40178 ( .A(n40463), .B(n40464), .Z(n40451) );
  AND U40179 ( .A(n40465), .B(n40466), .Z(n40464) );
  XOR U40180 ( .A(n40463), .B(n38652), .Z(n40466) );
  XOR U40181 ( .A(n40467), .B(n40468), .Z(n38652) );
  AND U40182 ( .A(n595), .B(n40469), .Z(n40468) );
  XOR U40183 ( .A(n40470), .B(n40467), .Z(n40469) );
  XNOR U40184 ( .A(n38649), .B(n40463), .Z(n40465) );
  XOR U40185 ( .A(n40471), .B(n40472), .Z(n38649) );
  AND U40186 ( .A(n592), .B(n40473), .Z(n40472) );
  XOR U40187 ( .A(n40474), .B(n40471), .Z(n40473) );
  XOR U40188 ( .A(n40475), .B(n40476), .Z(n40463) );
  AND U40189 ( .A(n40477), .B(n40478), .Z(n40476) );
  XOR U40190 ( .A(n40475), .B(n38664), .Z(n40478) );
  XOR U40191 ( .A(n40479), .B(n40480), .Z(n38664) );
  AND U40192 ( .A(n595), .B(n40481), .Z(n40480) );
  XOR U40193 ( .A(n40482), .B(n40479), .Z(n40481) );
  XNOR U40194 ( .A(n38661), .B(n40475), .Z(n40477) );
  XOR U40195 ( .A(n40483), .B(n40484), .Z(n38661) );
  AND U40196 ( .A(n592), .B(n40485), .Z(n40484) );
  XOR U40197 ( .A(n40486), .B(n40483), .Z(n40485) );
  XOR U40198 ( .A(n40487), .B(n40488), .Z(n40475) );
  AND U40199 ( .A(n40489), .B(n40490), .Z(n40488) );
  XOR U40200 ( .A(n40487), .B(n38676), .Z(n40490) );
  XOR U40201 ( .A(n40491), .B(n40492), .Z(n38676) );
  AND U40202 ( .A(n595), .B(n40493), .Z(n40492) );
  XOR U40203 ( .A(n40494), .B(n40491), .Z(n40493) );
  XNOR U40204 ( .A(n38673), .B(n40487), .Z(n40489) );
  XOR U40205 ( .A(n40495), .B(n40496), .Z(n38673) );
  AND U40206 ( .A(n592), .B(n40497), .Z(n40496) );
  XOR U40207 ( .A(n40498), .B(n40495), .Z(n40497) );
  XOR U40208 ( .A(n40499), .B(n40500), .Z(n40487) );
  AND U40209 ( .A(n40501), .B(n40502), .Z(n40500) );
  XOR U40210 ( .A(n40499), .B(n38688), .Z(n40502) );
  XOR U40211 ( .A(n40503), .B(n40504), .Z(n38688) );
  AND U40212 ( .A(n595), .B(n40505), .Z(n40504) );
  XOR U40213 ( .A(n40506), .B(n40503), .Z(n40505) );
  XNOR U40214 ( .A(n38685), .B(n40499), .Z(n40501) );
  XOR U40215 ( .A(n40507), .B(n40508), .Z(n38685) );
  AND U40216 ( .A(n592), .B(n40509), .Z(n40508) );
  XOR U40217 ( .A(n40510), .B(n40507), .Z(n40509) );
  XOR U40218 ( .A(n40511), .B(n40512), .Z(n40499) );
  AND U40219 ( .A(n40513), .B(n40514), .Z(n40512) );
  XOR U40220 ( .A(n40511), .B(n38700), .Z(n40514) );
  XOR U40221 ( .A(n40515), .B(n40516), .Z(n38700) );
  AND U40222 ( .A(n595), .B(n40517), .Z(n40516) );
  XOR U40223 ( .A(n40518), .B(n40515), .Z(n40517) );
  XNOR U40224 ( .A(n38697), .B(n40511), .Z(n40513) );
  XOR U40225 ( .A(n40519), .B(n40520), .Z(n38697) );
  AND U40226 ( .A(n592), .B(n40521), .Z(n40520) );
  XOR U40227 ( .A(n40522), .B(n40519), .Z(n40521) );
  XOR U40228 ( .A(n40523), .B(n40524), .Z(n40511) );
  AND U40229 ( .A(n40525), .B(n40526), .Z(n40524) );
  XNOR U40230 ( .A(n40527), .B(n38713), .Z(n40526) );
  XOR U40231 ( .A(n40528), .B(n40529), .Z(n38713) );
  AND U40232 ( .A(n595), .B(n40530), .Z(n40529) );
  XOR U40233 ( .A(n40528), .B(n40531), .Z(n40530) );
  XNOR U40234 ( .A(n38710), .B(n40523), .Z(n40525) );
  XOR U40235 ( .A(n40532), .B(n40533), .Z(n38710) );
  AND U40236 ( .A(n592), .B(n40534), .Z(n40533) );
  XOR U40237 ( .A(n40532), .B(n40535), .Z(n40534) );
  IV U40238 ( .A(n40527), .Z(n40523) );
  AND U40239 ( .A(n40159), .B(n40162), .Z(n40527) );
  XNOR U40240 ( .A(n40536), .B(n40537), .Z(n40162) );
  AND U40241 ( .A(n595), .B(n40538), .Z(n40537) );
  XNOR U40242 ( .A(n40539), .B(n40536), .Z(n40538) );
  XOR U40243 ( .A(n40540), .B(n40541), .Z(n595) );
  AND U40244 ( .A(n40542), .B(n40543), .Z(n40541) );
  XOR U40245 ( .A(n40170), .B(n40540), .Z(n40543) );
  IV U40246 ( .A(n40544), .Z(n40170) );
  AND U40247 ( .A(p_input[2815]), .B(p_input[2783]), .Z(n40544) );
  XOR U40248 ( .A(n40540), .B(n40167), .Z(n40542) );
  AND U40249 ( .A(p_input[2719]), .B(p_input[2751]), .Z(n40167) );
  XOR U40250 ( .A(n40545), .B(n40546), .Z(n40540) );
  AND U40251 ( .A(n40547), .B(n40548), .Z(n40546) );
  XOR U40252 ( .A(n40545), .B(n40182), .Z(n40548) );
  XNOR U40253 ( .A(p_input[2782]), .B(n40549), .Z(n40182) );
  AND U40254 ( .A(n763), .B(n40550), .Z(n40549) );
  XOR U40255 ( .A(p_input[2814]), .B(p_input[2782]), .Z(n40550) );
  XNOR U40256 ( .A(n40179), .B(n40545), .Z(n40547) );
  XOR U40257 ( .A(n40551), .B(n40552), .Z(n40179) );
  AND U40258 ( .A(n761), .B(n40553), .Z(n40552) );
  XOR U40259 ( .A(p_input[2750]), .B(p_input[2718]), .Z(n40553) );
  XOR U40260 ( .A(n40554), .B(n40555), .Z(n40545) );
  AND U40261 ( .A(n40556), .B(n40557), .Z(n40555) );
  XOR U40262 ( .A(n40554), .B(n40194), .Z(n40557) );
  XNOR U40263 ( .A(p_input[2781]), .B(n40558), .Z(n40194) );
  AND U40264 ( .A(n763), .B(n40559), .Z(n40558) );
  XOR U40265 ( .A(p_input[2813]), .B(p_input[2781]), .Z(n40559) );
  XNOR U40266 ( .A(n40191), .B(n40554), .Z(n40556) );
  XOR U40267 ( .A(n40560), .B(n40561), .Z(n40191) );
  AND U40268 ( .A(n761), .B(n40562), .Z(n40561) );
  XOR U40269 ( .A(p_input[2749]), .B(p_input[2717]), .Z(n40562) );
  XOR U40270 ( .A(n40563), .B(n40564), .Z(n40554) );
  AND U40271 ( .A(n40565), .B(n40566), .Z(n40564) );
  XOR U40272 ( .A(n40563), .B(n40206), .Z(n40566) );
  XNOR U40273 ( .A(p_input[2780]), .B(n40567), .Z(n40206) );
  AND U40274 ( .A(n763), .B(n40568), .Z(n40567) );
  XOR U40275 ( .A(p_input[2812]), .B(p_input[2780]), .Z(n40568) );
  XNOR U40276 ( .A(n40203), .B(n40563), .Z(n40565) );
  XOR U40277 ( .A(n40569), .B(n40570), .Z(n40203) );
  AND U40278 ( .A(n761), .B(n40571), .Z(n40570) );
  XOR U40279 ( .A(p_input[2748]), .B(p_input[2716]), .Z(n40571) );
  XOR U40280 ( .A(n40572), .B(n40573), .Z(n40563) );
  AND U40281 ( .A(n40574), .B(n40575), .Z(n40573) );
  XOR U40282 ( .A(n40572), .B(n40218), .Z(n40575) );
  XNOR U40283 ( .A(p_input[2779]), .B(n40576), .Z(n40218) );
  AND U40284 ( .A(n763), .B(n40577), .Z(n40576) );
  XOR U40285 ( .A(p_input[2811]), .B(p_input[2779]), .Z(n40577) );
  XNOR U40286 ( .A(n40215), .B(n40572), .Z(n40574) );
  XOR U40287 ( .A(n40578), .B(n40579), .Z(n40215) );
  AND U40288 ( .A(n761), .B(n40580), .Z(n40579) );
  XOR U40289 ( .A(p_input[2747]), .B(p_input[2715]), .Z(n40580) );
  XOR U40290 ( .A(n40581), .B(n40582), .Z(n40572) );
  AND U40291 ( .A(n40583), .B(n40584), .Z(n40582) );
  XOR U40292 ( .A(n40581), .B(n40230), .Z(n40584) );
  XNOR U40293 ( .A(p_input[2778]), .B(n40585), .Z(n40230) );
  AND U40294 ( .A(n763), .B(n40586), .Z(n40585) );
  XOR U40295 ( .A(p_input[2810]), .B(p_input[2778]), .Z(n40586) );
  XNOR U40296 ( .A(n40227), .B(n40581), .Z(n40583) );
  XOR U40297 ( .A(n40587), .B(n40588), .Z(n40227) );
  AND U40298 ( .A(n761), .B(n40589), .Z(n40588) );
  XOR U40299 ( .A(p_input[2746]), .B(p_input[2714]), .Z(n40589) );
  XOR U40300 ( .A(n40590), .B(n40591), .Z(n40581) );
  AND U40301 ( .A(n40592), .B(n40593), .Z(n40591) );
  XOR U40302 ( .A(n40590), .B(n40242), .Z(n40593) );
  XNOR U40303 ( .A(p_input[2777]), .B(n40594), .Z(n40242) );
  AND U40304 ( .A(n763), .B(n40595), .Z(n40594) );
  XOR U40305 ( .A(p_input[2809]), .B(p_input[2777]), .Z(n40595) );
  XNOR U40306 ( .A(n40239), .B(n40590), .Z(n40592) );
  XOR U40307 ( .A(n40596), .B(n40597), .Z(n40239) );
  AND U40308 ( .A(n761), .B(n40598), .Z(n40597) );
  XOR U40309 ( .A(p_input[2745]), .B(p_input[2713]), .Z(n40598) );
  XOR U40310 ( .A(n40599), .B(n40600), .Z(n40590) );
  AND U40311 ( .A(n40601), .B(n40602), .Z(n40600) );
  XOR U40312 ( .A(n40599), .B(n40254), .Z(n40602) );
  XNOR U40313 ( .A(p_input[2776]), .B(n40603), .Z(n40254) );
  AND U40314 ( .A(n763), .B(n40604), .Z(n40603) );
  XOR U40315 ( .A(p_input[2808]), .B(p_input[2776]), .Z(n40604) );
  XNOR U40316 ( .A(n40251), .B(n40599), .Z(n40601) );
  XOR U40317 ( .A(n40605), .B(n40606), .Z(n40251) );
  AND U40318 ( .A(n761), .B(n40607), .Z(n40606) );
  XOR U40319 ( .A(p_input[2744]), .B(p_input[2712]), .Z(n40607) );
  XOR U40320 ( .A(n40608), .B(n40609), .Z(n40599) );
  AND U40321 ( .A(n40610), .B(n40611), .Z(n40609) );
  XOR U40322 ( .A(n40608), .B(n40266), .Z(n40611) );
  XNOR U40323 ( .A(p_input[2775]), .B(n40612), .Z(n40266) );
  AND U40324 ( .A(n763), .B(n40613), .Z(n40612) );
  XOR U40325 ( .A(p_input[2807]), .B(p_input[2775]), .Z(n40613) );
  XNOR U40326 ( .A(n40263), .B(n40608), .Z(n40610) );
  XOR U40327 ( .A(n40614), .B(n40615), .Z(n40263) );
  AND U40328 ( .A(n761), .B(n40616), .Z(n40615) );
  XOR U40329 ( .A(p_input[2743]), .B(p_input[2711]), .Z(n40616) );
  XOR U40330 ( .A(n40617), .B(n40618), .Z(n40608) );
  AND U40331 ( .A(n40619), .B(n40620), .Z(n40618) );
  XOR U40332 ( .A(n40617), .B(n40278), .Z(n40620) );
  XNOR U40333 ( .A(p_input[2774]), .B(n40621), .Z(n40278) );
  AND U40334 ( .A(n763), .B(n40622), .Z(n40621) );
  XOR U40335 ( .A(p_input[2806]), .B(p_input[2774]), .Z(n40622) );
  XNOR U40336 ( .A(n40275), .B(n40617), .Z(n40619) );
  XOR U40337 ( .A(n40623), .B(n40624), .Z(n40275) );
  AND U40338 ( .A(n761), .B(n40625), .Z(n40624) );
  XOR U40339 ( .A(p_input[2742]), .B(p_input[2710]), .Z(n40625) );
  XOR U40340 ( .A(n40626), .B(n40627), .Z(n40617) );
  AND U40341 ( .A(n40628), .B(n40629), .Z(n40627) );
  XOR U40342 ( .A(n40626), .B(n40290), .Z(n40629) );
  XNOR U40343 ( .A(p_input[2773]), .B(n40630), .Z(n40290) );
  AND U40344 ( .A(n763), .B(n40631), .Z(n40630) );
  XOR U40345 ( .A(p_input[2805]), .B(p_input[2773]), .Z(n40631) );
  XNOR U40346 ( .A(n40287), .B(n40626), .Z(n40628) );
  XOR U40347 ( .A(n40632), .B(n40633), .Z(n40287) );
  AND U40348 ( .A(n761), .B(n40634), .Z(n40633) );
  XOR U40349 ( .A(p_input[2741]), .B(p_input[2709]), .Z(n40634) );
  XOR U40350 ( .A(n40635), .B(n40636), .Z(n40626) );
  AND U40351 ( .A(n40637), .B(n40638), .Z(n40636) );
  XOR U40352 ( .A(n40635), .B(n40302), .Z(n40638) );
  XNOR U40353 ( .A(p_input[2772]), .B(n40639), .Z(n40302) );
  AND U40354 ( .A(n763), .B(n40640), .Z(n40639) );
  XOR U40355 ( .A(p_input[2804]), .B(p_input[2772]), .Z(n40640) );
  XNOR U40356 ( .A(n40299), .B(n40635), .Z(n40637) );
  XOR U40357 ( .A(n40641), .B(n40642), .Z(n40299) );
  AND U40358 ( .A(n761), .B(n40643), .Z(n40642) );
  XOR U40359 ( .A(p_input[2740]), .B(p_input[2708]), .Z(n40643) );
  XOR U40360 ( .A(n40644), .B(n40645), .Z(n40635) );
  AND U40361 ( .A(n40646), .B(n40647), .Z(n40645) );
  XOR U40362 ( .A(n40644), .B(n40314), .Z(n40647) );
  XNOR U40363 ( .A(p_input[2771]), .B(n40648), .Z(n40314) );
  AND U40364 ( .A(n763), .B(n40649), .Z(n40648) );
  XOR U40365 ( .A(p_input[2803]), .B(p_input[2771]), .Z(n40649) );
  XNOR U40366 ( .A(n40311), .B(n40644), .Z(n40646) );
  XOR U40367 ( .A(n40650), .B(n40651), .Z(n40311) );
  AND U40368 ( .A(n761), .B(n40652), .Z(n40651) );
  XOR U40369 ( .A(p_input[2739]), .B(p_input[2707]), .Z(n40652) );
  XOR U40370 ( .A(n40653), .B(n40654), .Z(n40644) );
  AND U40371 ( .A(n40655), .B(n40656), .Z(n40654) );
  XOR U40372 ( .A(n40653), .B(n40326), .Z(n40656) );
  XNOR U40373 ( .A(p_input[2770]), .B(n40657), .Z(n40326) );
  AND U40374 ( .A(n763), .B(n40658), .Z(n40657) );
  XOR U40375 ( .A(p_input[2802]), .B(p_input[2770]), .Z(n40658) );
  XNOR U40376 ( .A(n40323), .B(n40653), .Z(n40655) );
  XOR U40377 ( .A(n40659), .B(n40660), .Z(n40323) );
  AND U40378 ( .A(n761), .B(n40661), .Z(n40660) );
  XOR U40379 ( .A(p_input[2738]), .B(p_input[2706]), .Z(n40661) );
  XOR U40380 ( .A(n40662), .B(n40663), .Z(n40653) );
  AND U40381 ( .A(n40664), .B(n40665), .Z(n40663) );
  XOR U40382 ( .A(n40662), .B(n40338), .Z(n40665) );
  XNOR U40383 ( .A(p_input[2769]), .B(n40666), .Z(n40338) );
  AND U40384 ( .A(n763), .B(n40667), .Z(n40666) );
  XOR U40385 ( .A(p_input[2801]), .B(p_input[2769]), .Z(n40667) );
  XNOR U40386 ( .A(n40335), .B(n40662), .Z(n40664) );
  XOR U40387 ( .A(n40668), .B(n40669), .Z(n40335) );
  AND U40388 ( .A(n761), .B(n40670), .Z(n40669) );
  XOR U40389 ( .A(p_input[2737]), .B(p_input[2705]), .Z(n40670) );
  XOR U40390 ( .A(n40671), .B(n40672), .Z(n40662) );
  AND U40391 ( .A(n40673), .B(n40674), .Z(n40672) );
  XOR U40392 ( .A(n40671), .B(n40350), .Z(n40674) );
  XNOR U40393 ( .A(p_input[2768]), .B(n40675), .Z(n40350) );
  AND U40394 ( .A(n763), .B(n40676), .Z(n40675) );
  XOR U40395 ( .A(p_input[2800]), .B(p_input[2768]), .Z(n40676) );
  XNOR U40396 ( .A(n40347), .B(n40671), .Z(n40673) );
  XOR U40397 ( .A(n40677), .B(n40678), .Z(n40347) );
  AND U40398 ( .A(n761), .B(n40679), .Z(n40678) );
  XOR U40399 ( .A(p_input[2736]), .B(p_input[2704]), .Z(n40679) );
  XOR U40400 ( .A(n40680), .B(n40681), .Z(n40671) );
  AND U40401 ( .A(n40682), .B(n40683), .Z(n40681) );
  XOR U40402 ( .A(n40680), .B(n40362), .Z(n40683) );
  XNOR U40403 ( .A(p_input[2767]), .B(n40684), .Z(n40362) );
  AND U40404 ( .A(n763), .B(n40685), .Z(n40684) );
  XOR U40405 ( .A(p_input[2799]), .B(p_input[2767]), .Z(n40685) );
  XNOR U40406 ( .A(n40359), .B(n40680), .Z(n40682) );
  XOR U40407 ( .A(n40686), .B(n40687), .Z(n40359) );
  AND U40408 ( .A(n761), .B(n40688), .Z(n40687) );
  XOR U40409 ( .A(p_input[2735]), .B(p_input[2703]), .Z(n40688) );
  XOR U40410 ( .A(n40689), .B(n40690), .Z(n40680) );
  AND U40411 ( .A(n40691), .B(n40692), .Z(n40690) );
  XOR U40412 ( .A(n40689), .B(n40374), .Z(n40692) );
  XNOR U40413 ( .A(p_input[2766]), .B(n40693), .Z(n40374) );
  AND U40414 ( .A(n763), .B(n40694), .Z(n40693) );
  XOR U40415 ( .A(p_input[2798]), .B(p_input[2766]), .Z(n40694) );
  XNOR U40416 ( .A(n40371), .B(n40689), .Z(n40691) );
  XOR U40417 ( .A(n40695), .B(n40696), .Z(n40371) );
  AND U40418 ( .A(n761), .B(n40697), .Z(n40696) );
  XOR U40419 ( .A(p_input[2734]), .B(p_input[2702]), .Z(n40697) );
  XOR U40420 ( .A(n40698), .B(n40699), .Z(n40689) );
  AND U40421 ( .A(n40700), .B(n40701), .Z(n40699) );
  XOR U40422 ( .A(n40698), .B(n40386), .Z(n40701) );
  XNOR U40423 ( .A(p_input[2765]), .B(n40702), .Z(n40386) );
  AND U40424 ( .A(n763), .B(n40703), .Z(n40702) );
  XOR U40425 ( .A(p_input[2797]), .B(p_input[2765]), .Z(n40703) );
  XNOR U40426 ( .A(n40383), .B(n40698), .Z(n40700) );
  XOR U40427 ( .A(n40704), .B(n40705), .Z(n40383) );
  AND U40428 ( .A(n761), .B(n40706), .Z(n40705) );
  XOR U40429 ( .A(p_input[2733]), .B(p_input[2701]), .Z(n40706) );
  XOR U40430 ( .A(n40707), .B(n40708), .Z(n40698) );
  AND U40431 ( .A(n40709), .B(n40710), .Z(n40708) );
  XOR U40432 ( .A(n40707), .B(n40398), .Z(n40710) );
  XNOR U40433 ( .A(p_input[2764]), .B(n40711), .Z(n40398) );
  AND U40434 ( .A(n763), .B(n40712), .Z(n40711) );
  XOR U40435 ( .A(p_input[2796]), .B(p_input[2764]), .Z(n40712) );
  XNOR U40436 ( .A(n40395), .B(n40707), .Z(n40709) );
  XOR U40437 ( .A(n40713), .B(n40714), .Z(n40395) );
  AND U40438 ( .A(n761), .B(n40715), .Z(n40714) );
  XOR U40439 ( .A(p_input[2732]), .B(p_input[2700]), .Z(n40715) );
  XOR U40440 ( .A(n40716), .B(n40717), .Z(n40707) );
  AND U40441 ( .A(n40718), .B(n40719), .Z(n40717) );
  XOR U40442 ( .A(n40716), .B(n40410), .Z(n40719) );
  XNOR U40443 ( .A(p_input[2763]), .B(n40720), .Z(n40410) );
  AND U40444 ( .A(n763), .B(n40721), .Z(n40720) );
  XOR U40445 ( .A(p_input[2795]), .B(p_input[2763]), .Z(n40721) );
  XNOR U40446 ( .A(n40407), .B(n40716), .Z(n40718) );
  XOR U40447 ( .A(n40722), .B(n40723), .Z(n40407) );
  AND U40448 ( .A(n761), .B(n40724), .Z(n40723) );
  XOR U40449 ( .A(p_input[2731]), .B(p_input[2699]), .Z(n40724) );
  XOR U40450 ( .A(n40725), .B(n40726), .Z(n40716) );
  AND U40451 ( .A(n40727), .B(n40728), .Z(n40726) );
  XOR U40452 ( .A(n40725), .B(n40422), .Z(n40728) );
  XNOR U40453 ( .A(p_input[2762]), .B(n40729), .Z(n40422) );
  AND U40454 ( .A(n763), .B(n40730), .Z(n40729) );
  XOR U40455 ( .A(p_input[2794]), .B(p_input[2762]), .Z(n40730) );
  XNOR U40456 ( .A(n40419), .B(n40725), .Z(n40727) );
  XOR U40457 ( .A(n40731), .B(n40732), .Z(n40419) );
  AND U40458 ( .A(n761), .B(n40733), .Z(n40732) );
  XOR U40459 ( .A(p_input[2730]), .B(p_input[2698]), .Z(n40733) );
  XOR U40460 ( .A(n40734), .B(n40735), .Z(n40725) );
  AND U40461 ( .A(n40736), .B(n40737), .Z(n40735) );
  XOR U40462 ( .A(n40734), .B(n40434), .Z(n40737) );
  XNOR U40463 ( .A(p_input[2761]), .B(n40738), .Z(n40434) );
  AND U40464 ( .A(n763), .B(n40739), .Z(n40738) );
  XOR U40465 ( .A(p_input[2793]), .B(p_input[2761]), .Z(n40739) );
  XNOR U40466 ( .A(n40431), .B(n40734), .Z(n40736) );
  XOR U40467 ( .A(n40740), .B(n40741), .Z(n40431) );
  AND U40468 ( .A(n761), .B(n40742), .Z(n40741) );
  XOR U40469 ( .A(p_input[2729]), .B(p_input[2697]), .Z(n40742) );
  XOR U40470 ( .A(n40743), .B(n40744), .Z(n40734) );
  AND U40471 ( .A(n40745), .B(n40746), .Z(n40744) );
  XOR U40472 ( .A(n40743), .B(n40446), .Z(n40746) );
  XNOR U40473 ( .A(p_input[2760]), .B(n40747), .Z(n40446) );
  AND U40474 ( .A(n763), .B(n40748), .Z(n40747) );
  XOR U40475 ( .A(p_input[2792]), .B(p_input[2760]), .Z(n40748) );
  XNOR U40476 ( .A(n40443), .B(n40743), .Z(n40745) );
  XOR U40477 ( .A(n40749), .B(n40750), .Z(n40443) );
  AND U40478 ( .A(n761), .B(n40751), .Z(n40750) );
  XOR U40479 ( .A(p_input[2728]), .B(p_input[2696]), .Z(n40751) );
  XOR U40480 ( .A(n40752), .B(n40753), .Z(n40743) );
  AND U40481 ( .A(n40754), .B(n40755), .Z(n40753) );
  XOR U40482 ( .A(n40752), .B(n40458), .Z(n40755) );
  XNOR U40483 ( .A(p_input[2759]), .B(n40756), .Z(n40458) );
  AND U40484 ( .A(n763), .B(n40757), .Z(n40756) );
  XOR U40485 ( .A(p_input[2791]), .B(p_input[2759]), .Z(n40757) );
  XNOR U40486 ( .A(n40455), .B(n40752), .Z(n40754) );
  XOR U40487 ( .A(n40758), .B(n40759), .Z(n40455) );
  AND U40488 ( .A(n761), .B(n40760), .Z(n40759) );
  XOR U40489 ( .A(p_input[2727]), .B(p_input[2695]), .Z(n40760) );
  XOR U40490 ( .A(n40761), .B(n40762), .Z(n40752) );
  AND U40491 ( .A(n40763), .B(n40764), .Z(n40762) );
  XOR U40492 ( .A(n40761), .B(n40470), .Z(n40764) );
  XNOR U40493 ( .A(p_input[2758]), .B(n40765), .Z(n40470) );
  AND U40494 ( .A(n763), .B(n40766), .Z(n40765) );
  XOR U40495 ( .A(p_input[2790]), .B(p_input[2758]), .Z(n40766) );
  XNOR U40496 ( .A(n40467), .B(n40761), .Z(n40763) );
  XOR U40497 ( .A(n40767), .B(n40768), .Z(n40467) );
  AND U40498 ( .A(n761), .B(n40769), .Z(n40768) );
  XOR U40499 ( .A(p_input[2726]), .B(p_input[2694]), .Z(n40769) );
  XOR U40500 ( .A(n40770), .B(n40771), .Z(n40761) );
  AND U40501 ( .A(n40772), .B(n40773), .Z(n40771) );
  XOR U40502 ( .A(n40770), .B(n40482), .Z(n40773) );
  XNOR U40503 ( .A(p_input[2757]), .B(n40774), .Z(n40482) );
  AND U40504 ( .A(n763), .B(n40775), .Z(n40774) );
  XOR U40505 ( .A(p_input[2789]), .B(p_input[2757]), .Z(n40775) );
  XNOR U40506 ( .A(n40479), .B(n40770), .Z(n40772) );
  XOR U40507 ( .A(n40776), .B(n40777), .Z(n40479) );
  AND U40508 ( .A(n761), .B(n40778), .Z(n40777) );
  XOR U40509 ( .A(p_input[2725]), .B(p_input[2693]), .Z(n40778) );
  XOR U40510 ( .A(n40779), .B(n40780), .Z(n40770) );
  AND U40511 ( .A(n40781), .B(n40782), .Z(n40780) );
  XOR U40512 ( .A(n40779), .B(n40494), .Z(n40782) );
  XNOR U40513 ( .A(p_input[2756]), .B(n40783), .Z(n40494) );
  AND U40514 ( .A(n763), .B(n40784), .Z(n40783) );
  XOR U40515 ( .A(p_input[2788]), .B(p_input[2756]), .Z(n40784) );
  XNOR U40516 ( .A(n40491), .B(n40779), .Z(n40781) );
  XOR U40517 ( .A(n40785), .B(n40786), .Z(n40491) );
  AND U40518 ( .A(n761), .B(n40787), .Z(n40786) );
  XOR U40519 ( .A(p_input[2724]), .B(p_input[2692]), .Z(n40787) );
  XOR U40520 ( .A(n40788), .B(n40789), .Z(n40779) );
  AND U40521 ( .A(n40790), .B(n40791), .Z(n40789) );
  XOR U40522 ( .A(n40788), .B(n40506), .Z(n40791) );
  XNOR U40523 ( .A(p_input[2755]), .B(n40792), .Z(n40506) );
  AND U40524 ( .A(n763), .B(n40793), .Z(n40792) );
  XOR U40525 ( .A(p_input[2787]), .B(p_input[2755]), .Z(n40793) );
  XNOR U40526 ( .A(n40503), .B(n40788), .Z(n40790) );
  XOR U40527 ( .A(n40794), .B(n40795), .Z(n40503) );
  AND U40528 ( .A(n761), .B(n40796), .Z(n40795) );
  XOR U40529 ( .A(p_input[2723]), .B(p_input[2691]), .Z(n40796) );
  XOR U40530 ( .A(n40797), .B(n40798), .Z(n40788) );
  AND U40531 ( .A(n40799), .B(n40800), .Z(n40798) );
  XOR U40532 ( .A(n40797), .B(n40518), .Z(n40800) );
  XNOR U40533 ( .A(p_input[2754]), .B(n40801), .Z(n40518) );
  AND U40534 ( .A(n763), .B(n40802), .Z(n40801) );
  XOR U40535 ( .A(p_input[2786]), .B(p_input[2754]), .Z(n40802) );
  XNOR U40536 ( .A(n40515), .B(n40797), .Z(n40799) );
  XOR U40537 ( .A(n40803), .B(n40804), .Z(n40515) );
  AND U40538 ( .A(n761), .B(n40805), .Z(n40804) );
  XOR U40539 ( .A(p_input[2722]), .B(p_input[2690]), .Z(n40805) );
  XOR U40540 ( .A(n40806), .B(n40807), .Z(n40797) );
  AND U40541 ( .A(n40808), .B(n40809), .Z(n40807) );
  XNOR U40542 ( .A(n40810), .B(n40531), .Z(n40809) );
  XNOR U40543 ( .A(p_input[2753]), .B(n40811), .Z(n40531) );
  AND U40544 ( .A(n763), .B(n40812), .Z(n40811) );
  XNOR U40545 ( .A(p_input[2785]), .B(n40813), .Z(n40812) );
  IV U40546 ( .A(p_input[2753]), .Z(n40813) );
  XNOR U40547 ( .A(n40528), .B(n40806), .Z(n40808) );
  XNOR U40548 ( .A(p_input[2689]), .B(n40814), .Z(n40528) );
  AND U40549 ( .A(n761), .B(n40815), .Z(n40814) );
  XOR U40550 ( .A(p_input[2721]), .B(p_input[2689]), .Z(n40815) );
  IV U40551 ( .A(n40810), .Z(n40806) );
  AND U40552 ( .A(n40536), .B(n40539), .Z(n40810) );
  XOR U40553 ( .A(p_input[2752]), .B(n40816), .Z(n40539) );
  AND U40554 ( .A(n763), .B(n40817), .Z(n40816) );
  XOR U40555 ( .A(p_input[2784]), .B(p_input[2752]), .Z(n40817) );
  XOR U40556 ( .A(n40818), .B(n40819), .Z(n763) );
  AND U40557 ( .A(n40820), .B(n40821), .Z(n40819) );
  XNOR U40558 ( .A(p_input[2815]), .B(n40818), .Z(n40821) );
  XOR U40559 ( .A(n40818), .B(p_input[2783]), .Z(n40820) );
  XOR U40560 ( .A(n40822), .B(n40823), .Z(n40818) );
  AND U40561 ( .A(n40824), .B(n40825), .Z(n40823) );
  XNOR U40562 ( .A(p_input[2814]), .B(n40822), .Z(n40825) );
  XOR U40563 ( .A(n40822), .B(p_input[2782]), .Z(n40824) );
  XOR U40564 ( .A(n40826), .B(n40827), .Z(n40822) );
  AND U40565 ( .A(n40828), .B(n40829), .Z(n40827) );
  XNOR U40566 ( .A(p_input[2813]), .B(n40826), .Z(n40829) );
  XOR U40567 ( .A(n40826), .B(p_input[2781]), .Z(n40828) );
  XOR U40568 ( .A(n40830), .B(n40831), .Z(n40826) );
  AND U40569 ( .A(n40832), .B(n40833), .Z(n40831) );
  XNOR U40570 ( .A(p_input[2812]), .B(n40830), .Z(n40833) );
  XOR U40571 ( .A(n40830), .B(p_input[2780]), .Z(n40832) );
  XOR U40572 ( .A(n40834), .B(n40835), .Z(n40830) );
  AND U40573 ( .A(n40836), .B(n40837), .Z(n40835) );
  XNOR U40574 ( .A(p_input[2811]), .B(n40834), .Z(n40837) );
  XOR U40575 ( .A(n40834), .B(p_input[2779]), .Z(n40836) );
  XOR U40576 ( .A(n40838), .B(n40839), .Z(n40834) );
  AND U40577 ( .A(n40840), .B(n40841), .Z(n40839) );
  XNOR U40578 ( .A(p_input[2810]), .B(n40838), .Z(n40841) );
  XOR U40579 ( .A(n40838), .B(p_input[2778]), .Z(n40840) );
  XOR U40580 ( .A(n40842), .B(n40843), .Z(n40838) );
  AND U40581 ( .A(n40844), .B(n40845), .Z(n40843) );
  XNOR U40582 ( .A(p_input[2809]), .B(n40842), .Z(n40845) );
  XOR U40583 ( .A(n40842), .B(p_input[2777]), .Z(n40844) );
  XOR U40584 ( .A(n40846), .B(n40847), .Z(n40842) );
  AND U40585 ( .A(n40848), .B(n40849), .Z(n40847) );
  XNOR U40586 ( .A(p_input[2808]), .B(n40846), .Z(n40849) );
  XOR U40587 ( .A(n40846), .B(p_input[2776]), .Z(n40848) );
  XOR U40588 ( .A(n40850), .B(n40851), .Z(n40846) );
  AND U40589 ( .A(n40852), .B(n40853), .Z(n40851) );
  XNOR U40590 ( .A(p_input[2807]), .B(n40850), .Z(n40853) );
  XOR U40591 ( .A(n40850), .B(p_input[2775]), .Z(n40852) );
  XOR U40592 ( .A(n40854), .B(n40855), .Z(n40850) );
  AND U40593 ( .A(n40856), .B(n40857), .Z(n40855) );
  XNOR U40594 ( .A(p_input[2806]), .B(n40854), .Z(n40857) );
  XOR U40595 ( .A(n40854), .B(p_input[2774]), .Z(n40856) );
  XOR U40596 ( .A(n40858), .B(n40859), .Z(n40854) );
  AND U40597 ( .A(n40860), .B(n40861), .Z(n40859) );
  XNOR U40598 ( .A(p_input[2805]), .B(n40858), .Z(n40861) );
  XOR U40599 ( .A(n40858), .B(p_input[2773]), .Z(n40860) );
  XOR U40600 ( .A(n40862), .B(n40863), .Z(n40858) );
  AND U40601 ( .A(n40864), .B(n40865), .Z(n40863) );
  XNOR U40602 ( .A(p_input[2804]), .B(n40862), .Z(n40865) );
  XOR U40603 ( .A(n40862), .B(p_input[2772]), .Z(n40864) );
  XOR U40604 ( .A(n40866), .B(n40867), .Z(n40862) );
  AND U40605 ( .A(n40868), .B(n40869), .Z(n40867) );
  XNOR U40606 ( .A(p_input[2803]), .B(n40866), .Z(n40869) );
  XOR U40607 ( .A(n40866), .B(p_input[2771]), .Z(n40868) );
  XOR U40608 ( .A(n40870), .B(n40871), .Z(n40866) );
  AND U40609 ( .A(n40872), .B(n40873), .Z(n40871) );
  XNOR U40610 ( .A(p_input[2802]), .B(n40870), .Z(n40873) );
  XOR U40611 ( .A(n40870), .B(p_input[2770]), .Z(n40872) );
  XOR U40612 ( .A(n40874), .B(n40875), .Z(n40870) );
  AND U40613 ( .A(n40876), .B(n40877), .Z(n40875) );
  XNOR U40614 ( .A(p_input[2801]), .B(n40874), .Z(n40877) );
  XOR U40615 ( .A(n40874), .B(p_input[2769]), .Z(n40876) );
  XOR U40616 ( .A(n40878), .B(n40879), .Z(n40874) );
  AND U40617 ( .A(n40880), .B(n40881), .Z(n40879) );
  XNOR U40618 ( .A(p_input[2800]), .B(n40878), .Z(n40881) );
  XOR U40619 ( .A(n40878), .B(p_input[2768]), .Z(n40880) );
  XOR U40620 ( .A(n40882), .B(n40883), .Z(n40878) );
  AND U40621 ( .A(n40884), .B(n40885), .Z(n40883) );
  XNOR U40622 ( .A(p_input[2799]), .B(n40882), .Z(n40885) );
  XOR U40623 ( .A(n40882), .B(p_input[2767]), .Z(n40884) );
  XOR U40624 ( .A(n40886), .B(n40887), .Z(n40882) );
  AND U40625 ( .A(n40888), .B(n40889), .Z(n40887) );
  XNOR U40626 ( .A(p_input[2798]), .B(n40886), .Z(n40889) );
  XOR U40627 ( .A(n40886), .B(p_input[2766]), .Z(n40888) );
  XOR U40628 ( .A(n40890), .B(n40891), .Z(n40886) );
  AND U40629 ( .A(n40892), .B(n40893), .Z(n40891) );
  XNOR U40630 ( .A(p_input[2797]), .B(n40890), .Z(n40893) );
  XOR U40631 ( .A(n40890), .B(p_input[2765]), .Z(n40892) );
  XOR U40632 ( .A(n40894), .B(n40895), .Z(n40890) );
  AND U40633 ( .A(n40896), .B(n40897), .Z(n40895) );
  XNOR U40634 ( .A(p_input[2796]), .B(n40894), .Z(n40897) );
  XOR U40635 ( .A(n40894), .B(p_input[2764]), .Z(n40896) );
  XOR U40636 ( .A(n40898), .B(n40899), .Z(n40894) );
  AND U40637 ( .A(n40900), .B(n40901), .Z(n40899) );
  XNOR U40638 ( .A(p_input[2795]), .B(n40898), .Z(n40901) );
  XOR U40639 ( .A(n40898), .B(p_input[2763]), .Z(n40900) );
  XOR U40640 ( .A(n40902), .B(n40903), .Z(n40898) );
  AND U40641 ( .A(n40904), .B(n40905), .Z(n40903) );
  XNOR U40642 ( .A(p_input[2794]), .B(n40902), .Z(n40905) );
  XOR U40643 ( .A(n40902), .B(p_input[2762]), .Z(n40904) );
  XOR U40644 ( .A(n40906), .B(n40907), .Z(n40902) );
  AND U40645 ( .A(n40908), .B(n40909), .Z(n40907) );
  XNOR U40646 ( .A(p_input[2793]), .B(n40906), .Z(n40909) );
  XOR U40647 ( .A(n40906), .B(p_input[2761]), .Z(n40908) );
  XOR U40648 ( .A(n40910), .B(n40911), .Z(n40906) );
  AND U40649 ( .A(n40912), .B(n40913), .Z(n40911) );
  XNOR U40650 ( .A(p_input[2792]), .B(n40910), .Z(n40913) );
  XOR U40651 ( .A(n40910), .B(p_input[2760]), .Z(n40912) );
  XOR U40652 ( .A(n40914), .B(n40915), .Z(n40910) );
  AND U40653 ( .A(n40916), .B(n40917), .Z(n40915) );
  XNOR U40654 ( .A(p_input[2791]), .B(n40914), .Z(n40917) );
  XOR U40655 ( .A(n40914), .B(p_input[2759]), .Z(n40916) );
  XOR U40656 ( .A(n40918), .B(n40919), .Z(n40914) );
  AND U40657 ( .A(n40920), .B(n40921), .Z(n40919) );
  XNOR U40658 ( .A(p_input[2790]), .B(n40918), .Z(n40921) );
  XOR U40659 ( .A(n40918), .B(p_input[2758]), .Z(n40920) );
  XOR U40660 ( .A(n40922), .B(n40923), .Z(n40918) );
  AND U40661 ( .A(n40924), .B(n40925), .Z(n40923) );
  XNOR U40662 ( .A(p_input[2789]), .B(n40922), .Z(n40925) );
  XOR U40663 ( .A(n40922), .B(p_input[2757]), .Z(n40924) );
  XOR U40664 ( .A(n40926), .B(n40927), .Z(n40922) );
  AND U40665 ( .A(n40928), .B(n40929), .Z(n40927) );
  XNOR U40666 ( .A(p_input[2788]), .B(n40926), .Z(n40929) );
  XOR U40667 ( .A(n40926), .B(p_input[2756]), .Z(n40928) );
  XOR U40668 ( .A(n40930), .B(n40931), .Z(n40926) );
  AND U40669 ( .A(n40932), .B(n40933), .Z(n40931) );
  XNOR U40670 ( .A(p_input[2787]), .B(n40930), .Z(n40933) );
  XOR U40671 ( .A(n40930), .B(p_input[2755]), .Z(n40932) );
  XOR U40672 ( .A(n40934), .B(n40935), .Z(n40930) );
  AND U40673 ( .A(n40936), .B(n40937), .Z(n40935) );
  XNOR U40674 ( .A(p_input[2786]), .B(n40934), .Z(n40937) );
  XOR U40675 ( .A(n40934), .B(p_input[2754]), .Z(n40936) );
  XNOR U40676 ( .A(n40938), .B(n40939), .Z(n40934) );
  AND U40677 ( .A(n40940), .B(n40941), .Z(n40939) );
  XOR U40678 ( .A(p_input[2785]), .B(n40938), .Z(n40941) );
  XNOR U40679 ( .A(p_input[2753]), .B(n40938), .Z(n40940) );
  AND U40680 ( .A(p_input[2784]), .B(n40942), .Z(n40938) );
  IV U40681 ( .A(p_input[2752]), .Z(n40942) );
  XNOR U40682 ( .A(p_input[2688]), .B(n40943), .Z(n40536) );
  AND U40683 ( .A(n761), .B(n40944), .Z(n40943) );
  XOR U40684 ( .A(p_input[2720]), .B(p_input[2688]), .Z(n40944) );
  XOR U40685 ( .A(n40945), .B(n40946), .Z(n761) );
  AND U40686 ( .A(n40947), .B(n40948), .Z(n40946) );
  XNOR U40687 ( .A(p_input[2751]), .B(n40945), .Z(n40948) );
  XOR U40688 ( .A(n40945), .B(p_input[2719]), .Z(n40947) );
  XOR U40689 ( .A(n40949), .B(n40950), .Z(n40945) );
  AND U40690 ( .A(n40951), .B(n40952), .Z(n40950) );
  XNOR U40691 ( .A(p_input[2750]), .B(n40949), .Z(n40952) );
  XNOR U40692 ( .A(n40949), .B(n40551), .Z(n40951) );
  IV U40693 ( .A(p_input[2718]), .Z(n40551) );
  XOR U40694 ( .A(n40953), .B(n40954), .Z(n40949) );
  AND U40695 ( .A(n40955), .B(n40956), .Z(n40954) );
  XNOR U40696 ( .A(p_input[2749]), .B(n40953), .Z(n40956) );
  XNOR U40697 ( .A(n40953), .B(n40560), .Z(n40955) );
  IV U40698 ( .A(p_input[2717]), .Z(n40560) );
  XOR U40699 ( .A(n40957), .B(n40958), .Z(n40953) );
  AND U40700 ( .A(n40959), .B(n40960), .Z(n40958) );
  XNOR U40701 ( .A(p_input[2748]), .B(n40957), .Z(n40960) );
  XNOR U40702 ( .A(n40957), .B(n40569), .Z(n40959) );
  IV U40703 ( .A(p_input[2716]), .Z(n40569) );
  XOR U40704 ( .A(n40961), .B(n40962), .Z(n40957) );
  AND U40705 ( .A(n40963), .B(n40964), .Z(n40962) );
  XNOR U40706 ( .A(p_input[2747]), .B(n40961), .Z(n40964) );
  XNOR U40707 ( .A(n40961), .B(n40578), .Z(n40963) );
  IV U40708 ( .A(p_input[2715]), .Z(n40578) );
  XOR U40709 ( .A(n40965), .B(n40966), .Z(n40961) );
  AND U40710 ( .A(n40967), .B(n40968), .Z(n40966) );
  XNOR U40711 ( .A(p_input[2746]), .B(n40965), .Z(n40968) );
  XNOR U40712 ( .A(n40965), .B(n40587), .Z(n40967) );
  IV U40713 ( .A(p_input[2714]), .Z(n40587) );
  XOR U40714 ( .A(n40969), .B(n40970), .Z(n40965) );
  AND U40715 ( .A(n40971), .B(n40972), .Z(n40970) );
  XNOR U40716 ( .A(p_input[2745]), .B(n40969), .Z(n40972) );
  XNOR U40717 ( .A(n40969), .B(n40596), .Z(n40971) );
  IV U40718 ( .A(p_input[2713]), .Z(n40596) );
  XOR U40719 ( .A(n40973), .B(n40974), .Z(n40969) );
  AND U40720 ( .A(n40975), .B(n40976), .Z(n40974) );
  XNOR U40721 ( .A(p_input[2744]), .B(n40973), .Z(n40976) );
  XNOR U40722 ( .A(n40973), .B(n40605), .Z(n40975) );
  IV U40723 ( .A(p_input[2712]), .Z(n40605) );
  XOR U40724 ( .A(n40977), .B(n40978), .Z(n40973) );
  AND U40725 ( .A(n40979), .B(n40980), .Z(n40978) );
  XNOR U40726 ( .A(p_input[2743]), .B(n40977), .Z(n40980) );
  XNOR U40727 ( .A(n40977), .B(n40614), .Z(n40979) );
  IV U40728 ( .A(p_input[2711]), .Z(n40614) );
  XOR U40729 ( .A(n40981), .B(n40982), .Z(n40977) );
  AND U40730 ( .A(n40983), .B(n40984), .Z(n40982) );
  XNOR U40731 ( .A(p_input[2742]), .B(n40981), .Z(n40984) );
  XNOR U40732 ( .A(n40981), .B(n40623), .Z(n40983) );
  IV U40733 ( .A(p_input[2710]), .Z(n40623) );
  XOR U40734 ( .A(n40985), .B(n40986), .Z(n40981) );
  AND U40735 ( .A(n40987), .B(n40988), .Z(n40986) );
  XNOR U40736 ( .A(p_input[2741]), .B(n40985), .Z(n40988) );
  XNOR U40737 ( .A(n40985), .B(n40632), .Z(n40987) );
  IV U40738 ( .A(p_input[2709]), .Z(n40632) );
  XOR U40739 ( .A(n40989), .B(n40990), .Z(n40985) );
  AND U40740 ( .A(n40991), .B(n40992), .Z(n40990) );
  XNOR U40741 ( .A(p_input[2740]), .B(n40989), .Z(n40992) );
  XNOR U40742 ( .A(n40989), .B(n40641), .Z(n40991) );
  IV U40743 ( .A(p_input[2708]), .Z(n40641) );
  XOR U40744 ( .A(n40993), .B(n40994), .Z(n40989) );
  AND U40745 ( .A(n40995), .B(n40996), .Z(n40994) );
  XNOR U40746 ( .A(p_input[2739]), .B(n40993), .Z(n40996) );
  XNOR U40747 ( .A(n40993), .B(n40650), .Z(n40995) );
  IV U40748 ( .A(p_input[2707]), .Z(n40650) );
  XOR U40749 ( .A(n40997), .B(n40998), .Z(n40993) );
  AND U40750 ( .A(n40999), .B(n41000), .Z(n40998) );
  XNOR U40751 ( .A(p_input[2738]), .B(n40997), .Z(n41000) );
  XNOR U40752 ( .A(n40997), .B(n40659), .Z(n40999) );
  IV U40753 ( .A(p_input[2706]), .Z(n40659) );
  XOR U40754 ( .A(n41001), .B(n41002), .Z(n40997) );
  AND U40755 ( .A(n41003), .B(n41004), .Z(n41002) );
  XNOR U40756 ( .A(p_input[2737]), .B(n41001), .Z(n41004) );
  XNOR U40757 ( .A(n41001), .B(n40668), .Z(n41003) );
  IV U40758 ( .A(p_input[2705]), .Z(n40668) );
  XOR U40759 ( .A(n41005), .B(n41006), .Z(n41001) );
  AND U40760 ( .A(n41007), .B(n41008), .Z(n41006) );
  XNOR U40761 ( .A(p_input[2736]), .B(n41005), .Z(n41008) );
  XNOR U40762 ( .A(n41005), .B(n40677), .Z(n41007) );
  IV U40763 ( .A(p_input[2704]), .Z(n40677) );
  XOR U40764 ( .A(n41009), .B(n41010), .Z(n41005) );
  AND U40765 ( .A(n41011), .B(n41012), .Z(n41010) );
  XNOR U40766 ( .A(p_input[2735]), .B(n41009), .Z(n41012) );
  XNOR U40767 ( .A(n41009), .B(n40686), .Z(n41011) );
  IV U40768 ( .A(p_input[2703]), .Z(n40686) );
  XOR U40769 ( .A(n41013), .B(n41014), .Z(n41009) );
  AND U40770 ( .A(n41015), .B(n41016), .Z(n41014) );
  XNOR U40771 ( .A(p_input[2734]), .B(n41013), .Z(n41016) );
  XNOR U40772 ( .A(n41013), .B(n40695), .Z(n41015) );
  IV U40773 ( .A(p_input[2702]), .Z(n40695) );
  XOR U40774 ( .A(n41017), .B(n41018), .Z(n41013) );
  AND U40775 ( .A(n41019), .B(n41020), .Z(n41018) );
  XNOR U40776 ( .A(p_input[2733]), .B(n41017), .Z(n41020) );
  XNOR U40777 ( .A(n41017), .B(n40704), .Z(n41019) );
  IV U40778 ( .A(p_input[2701]), .Z(n40704) );
  XOR U40779 ( .A(n41021), .B(n41022), .Z(n41017) );
  AND U40780 ( .A(n41023), .B(n41024), .Z(n41022) );
  XNOR U40781 ( .A(p_input[2732]), .B(n41021), .Z(n41024) );
  XNOR U40782 ( .A(n41021), .B(n40713), .Z(n41023) );
  IV U40783 ( .A(p_input[2700]), .Z(n40713) );
  XOR U40784 ( .A(n41025), .B(n41026), .Z(n41021) );
  AND U40785 ( .A(n41027), .B(n41028), .Z(n41026) );
  XNOR U40786 ( .A(p_input[2731]), .B(n41025), .Z(n41028) );
  XNOR U40787 ( .A(n41025), .B(n40722), .Z(n41027) );
  IV U40788 ( .A(p_input[2699]), .Z(n40722) );
  XOR U40789 ( .A(n41029), .B(n41030), .Z(n41025) );
  AND U40790 ( .A(n41031), .B(n41032), .Z(n41030) );
  XNOR U40791 ( .A(p_input[2730]), .B(n41029), .Z(n41032) );
  XNOR U40792 ( .A(n41029), .B(n40731), .Z(n41031) );
  IV U40793 ( .A(p_input[2698]), .Z(n40731) );
  XOR U40794 ( .A(n41033), .B(n41034), .Z(n41029) );
  AND U40795 ( .A(n41035), .B(n41036), .Z(n41034) );
  XNOR U40796 ( .A(p_input[2729]), .B(n41033), .Z(n41036) );
  XNOR U40797 ( .A(n41033), .B(n40740), .Z(n41035) );
  IV U40798 ( .A(p_input[2697]), .Z(n40740) );
  XOR U40799 ( .A(n41037), .B(n41038), .Z(n41033) );
  AND U40800 ( .A(n41039), .B(n41040), .Z(n41038) );
  XNOR U40801 ( .A(p_input[2728]), .B(n41037), .Z(n41040) );
  XNOR U40802 ( .A(n41037), .B(n40749), .Z(n41039) );
  IV U40803 ( .A(p_input[2696]), .Z(n40749) );
  XOR U40804 ( .A(n41041), .B(n41042), .Z(n41037) );
  AND U40805 ( .A(n41043), .B(n41044), .Z(n41042) );
  XNOR U40806 ( .A(p_input[2727]), .B(n41041), .Z(n41044) );
  XNOR U40807 ( .A(n41041), .B(n40758), .Z(n41043) );
  IV U40808 ( .A(p_input[2695]), .Z(n40758) );
  XOR U40809 ( .A(n41045), .B(n41046), .Z(n41041) );
  AND U40810 ( .A(n41047), .B(n41048), .Z(n41046) );
  XNOR U40811 ( .A(p_input[2726]), .B(n41045), .Z(n41048) );
  XNOR U40812 ( .A(n41045), .B(n40767), .Z(n41047) );
  IV U40813 ( .A(p_input[2694]), .Z(n40767) );
  XOR U40814 ( .A(n41049), .B(n41050), .Z(n41045) );
  AND U40815 ( .A(n41051), .B(n41052), .Z(n41050) );
  XNOR U40816 ( .A(p_input[2725]), .B(n41049), .Z(n41052) );
  XNOR U40817 ( .A(n41049), .B(n40776), .Z(n41051) );
  IV U40818 ( .A(p_input[2693]), .Z(n40776) );
  XOR U40819 ( .A(n41053), .B(n41054), .Z(n41049) );
  AND U40820 ( .A(n41055), .B(n41056), .Z(n41054) );
  XNOR U40821 ( .A(p_input[2724]), .B(n41053), .Z(n41056) );
  XNOR U40822 ( .A(n41053), .B(n40785), .Z(n41055) );
  IV U40823 ( .A(p_input[2692]), .Z(n40785) );
  XOR U40824 ( .A(n41057), .B(n41058), .Z(n41053) );
  AND U40825 ( .A(n41059), .B(n41060), .Z(n41058) );
  XNOR U40826 ( .A(p_input[2723]), .B(n41057), .Z(n41060) );
  XNOR U40827 ( .A(n41057), .B(n40794), .Z(n41059) );
  IV U40828 ( .A(p_input[2691]), .Z(n40794) );
  XOR U40829 ( .A(n41061), .B(n41062), .Z(n41057) );
  AND U40830 ( .A(n41063), .B(n41064), .Z(n41062) );
  XNOR U40831 ( .A(p_input[2722]), .B(n41061), .Z(n41064) );
  XNOR U40832 ( .A(n41061), .B(n40803), .Z(n41063) );
  IV U40833 ( .A(p_input[2690]), .Z(n40803) );
  XNOR U40834 ( .A(n41065), .B(n41066), .Z(n41061) );
  AND U40835 ( .A(n41067), .B(n41068), .Z(n41066) );
  XOR U40836 ( .A(p_input[2721]), .B(n41065), .Z(n41068) );
  XNOR U40837 ( .A(p_input[2689]), .B(n41065), .Z(n41067) );
  AND U40838 ( .A(p_input[2720]), .B(n41069), .Z(n41065) );
  IV U40839 ( .A(p_input[2688]), .Z(n41069) );
  XOR U40840 ( .A(n41070), .B(n41071), .Z(n40159) );
  AND U40841 ( .A(n592), .B(n41072), .Z(n41071) );
  XNOR U40842 ( .A(n41073), .B(n41070), .Z(n41072) );
  XOR U40843 ( .A(n41074), .B(n41075), .Z(n592) );
  AND U40844 ( .A(n41076), .B(n41077), .Z(n41075) );
  XNOR U40845 ( .A(n40174), .B(n41074), .Z(n41077) );
  AND U40846 ( .A(p_input[2687]), .B(p_input[2655]), .Z(n40174) );
  XNOR U40847 ( .A(n41074), .B(n40171), .Z(n41076) );
  IV U40848 ( .A(n41078), .Z(n40171) );
  AND U40849 ( .A(p_input[2591]), .B(p_input[2623]), .Z(n41078) );
  XOR U40850 ( .A(n41079), .B(n41080), .Z(n41074) );
  AND U40851 ( .A(n41081), .B(n41082), .Z(n41080) );
  XOR U40852 ( .A(n41079), .B(n40186), .Z(n41082) );
  XNOR U40853 ( .A(p_input[2654]), .B(n41083), .Z(n40186) );
  AND U40854 ( .A(n767), .B(n41084), .Z(n41083) );
  XOR U40855 ( .A(p_input[2686]), .B(p_input[2654]), .Z(n41084) );
  XNOR U40856 ( .A(n40183), .B(n41079), .Z(n41081) );
  XOR U40857 ( .A(n41085), .B(n41086), .Z(n40183) );
  AND U40858 ( .A(n764), .B(n41087), .Z(n41086) );
  XOR U40859 ( .A(p_input[2622]), .B(p_input[2590]), .Z(n41087) );
  XOR U40860 ( .A(n41088), .B(n41089), .Z(n41079) );
  AND U40861 ( .A(n41090), .B(n41091), .Z(n41089) );
  XOR U40862 ( .A(n41088), .B(n40198), .Z(n41091) );
  XNOR U40863 ( .A(p_input[2653]), .B(n41092), .Z(n40198) );
  AND U40864 ( .A(n767), .B(n41093), .Z(n41092) );
  XOR U40865 ( .A(p_input[2685]), .B(p_input[2653]), .Z(n41093) );
  XNOR U40866 ( .A(n40195), .B(n41088), .Z(n41090) );
  XOR U40867 ( .A(n41094), .B(n41095), .Z(n40195) );
  AND U40868 ( .A(n764), .B(n41096), .Z(n41095) );
  XOR U40869 ( .A(p_input[2621]), .B(p_input[2589]), .Z(n41096) );
  XOR U40870 ( .A(n41097), .B(n41098), .Z(n41088) );
  AND U40871 ( .A(n41099), .B(n41100), .Z(n41098) );
  XOR U40872 ( .A(n41097), .B(n40210), .Z(n41100) );
  XNOR U40873 ( .A(p_input[2652]), .B(n41101), .Z(n40210) );
  AND U40874 ( .A(n767), .B(n41102), .Z(n41101) );
  XOR U40875 ( .A(p_input[2684]), .B(p_input[2652]), .Z(n41102) );
  XNOR U40876 ( .A(n40207), .B(n41097), .Z(n41099) );
  XOR U40877 ( .A(n41103), .B(n41104), .Z(n40207) );
  AND U40878 ( .A(n764), .B(n41105), .Z(n41104) );
  XOR U40879 ( .A(p_input[2620]), .B(p_input[2588]), .Z(n41105) );
  XOR U40880 ( .A(n41106), .B(n41107), .Z(n41097) );
  AND U40881 ( .A(n41108), .B(n41109), .Z(n41107) );
  XOR U40882 ( .A(n41106), .B(n40222), .Z(n41109) );
  XNOR U40883 ( .A(p_input[2651]), .B(n41110), .Z(n40222) );
  AND U40884 ( .A(n767), .B(n41111), .Z(n41110) );
  XOR U40885 ( .A(p_input[2683]), .B(p_input[2651]), .Z(n41111) );
  XNOR U40886 ( .A(n40219), .B(n41106), .Z(n41108) );
  XOR U40887 ( .A(n41112), .B(n41113), .Z(n40219) );
  AND U40888 ( .A(n764), .B(n41114), .Z(n41113) );
  XOR U40889 ( .A(p_input[2619]), .B(p_input[2587]), .Z(n41114) );
  XOR U40890 ( .A(n41115), .B(n41116), .Z(n41106) );
  AND U40891 ( .A(n41117), .B(n41118), .Z(n41116) );
  XOR U40892 ( .A(n41115), .B(n40234), .Z(n41118) );
  XNOR U40893 ( .A(p_input[2650]), .B(n41119), .Z(n40234) );
  AND U40894 ( .A(n767), .B(n41120), .Z(n41119) );
  XOR U40895 ( .A(p_input[2682]), .B(p_input[2650]), .Z(n41120) );
  XNOR U40896 ( .A(n40231), .B(n41115), .Z(n41117) );
  XOR U40897 ( .A(n41121), .B(n41122), .Z(n40231) );
  AND U40898 ( .A(n764), .B(n41123), .Z(n41122) );
  XOR U40899 ( .A(p_input[2618]), .B(p_input[2586]), .Z(n41123) );
  XOR U40900 ( .A(n41124), .B(n41125), .Z(n41115) );
  AND U40901 ( .A(n41126), .B(n41127), .Z(n41125) );
  XOR U40902 ( .A(n41124), .B(n40246), .Z(n41127) );
  XNOR U40903 ( .A(p_input[2649]), .B(n41128), .Z(n40246) );
  AND U40904 ( .A(n767), .B(n41129), .Z(n41128) );
  XOR U40905 ( .A(p_input[2681]), .B(p_input[2649]), .Z(n41129) );
  XNOR U40906 ( .A(n40243), .B(n41124), .Z(n41126) );
  XOR U40907 ( .A(n41130), .B(n41131), .Z(n40243) );
  AND U40908 ( .A(n764), .B(n41132), .Z(n41131) );
  XOR U40909 ( .A(p_input[2617]), .B(p_input[2585]), .Z(n41132) );
  XOR U40910 ( .A(n41133), .B(n41134), .Z(n41124) );
  AND U40911 ( .A(n41135), .B(n41136), .Z(n41134) );
  XOR U40912 ( .A(n41133), .B(n40258), .Z(n41136) );
  XNOR U40913 ( .A(p_input[2648]), .B(n41137), .Z(n40258) );
  AND U40914 ( .A(n767), .B(n41138), .Z(n41137) );
  XOR U40915 ( .A(p_input[2680]), .B(p_input[2648]), .Z(n41138) );
  XNOR U40916 ( .A(n40255), .B(n41133), .Z(n41135) );
  XOR U40917 ( .A(n41139), .B(n41140), .Z(n40255) );
  AND U40918 ( .A(n764), .B(n41141), .Z(n41140) );
  XOR U40919 ( .A(p_input[2616]), .B(p_input[2584]), .Z(n41141) );
  XOR U40920 ( .A(n41142), .B(n41143), .Z(n41133) );
  AND U40921 ( .A(n41144), .B(n41145), .Z(n41143) );
  XOR U40922 ( .A(n41142), .B(n40270), .Z(n41145) );
  XNOR U40923 ( .A(p_input[2647]), .B(n41146), .Z(n40270) );
  AND U40924 ( .A(n767), .B(n41147), .Z(n41146) );
  XOR U40925 ( .A(p_input[2679]), .B(p_input[2647]), .Z(n41147) );
  XNOR U40926 ( .A(n40267), .B(n41142), .Z(n41144) );
  XOR U40927 ( .A(n41148), .B(n41149), .Z(n40267) );
  AND U40928 ( .A(n764), .B(n41150), .Z(n41149) );
  XOR U40929 ( .A(p_input[2615]), .B(p_input[2583]), .Z(n41150) );
  XOR U40930 ( .A(n41151), .B(n41152), .Z(n41142) );
  AND U40931 ( .A(n41153), .B(n41154), .Z(n41152) );
  XOR U40932 ( .A(n41151), .B(n40282), .Z(n41154) );
  XNOR U40933 ( .A(p_input[2646]), .B(n41155), .Z(n40282) );
  AND U40934 ( .A(n767), .B(n41156), .Z(n41155) );
  XOR U40935 ( .A(p_input[2678]), .B(p_input[2646]), .Z(n41156) );
  XNOR U40936 ( .A(n40279), .B(n41151), .Z(n41153) );
  XOR U40937 ( .A(n41157), .B(n41158), .Z(n40279) );
  AND U40938 ( .A(n764), .B(n41159), .Z(n41158) );
  XOR U40939 ( .A(p_input[2614]), .B(p_input[2582]), .Z(n41159) );
  XOR U40940 ( .A(n41160), .B(n41161), .Z(n41151) );
  AND U40941 ( .A(n41162), .B(n41163), .Z(n41161) );
  XOR U40942 ( .A(n41160), .B(n40294), .Z(n41163) );
  XNOR U40943 ( .A(p_input[2645]), .B(n41164), .Z(n40294) );
  AND U40944 ( .A(n767), .B(n41165), .Z(n41164) );
  XOR U40945 ( .A(p_input[2677]), .B(p_input[2645]), .Z(n41165) );
  XNOR U40946 ( .A(n40291), .B(n41160), .Z(n41162) );
  XOR U40947 ( .A(n41166), .B(n41167), .Z(n40291) );
  AND U40948 ( .A(n764), .B(n41168), .Z(n41167) );
  XOR U40949 ( .A(p_input[2613]), .B(p_input[2581]), .Z(n41168) );
  XOR U40950 ( .A(n41169), .B(n41170), .Z(n41160) );
  AND U40951 ( .A(n41171), .B(n41172), .Z(n41170) );
  XOR U40952 ( .A(n41169), .B(n40306), .Z(n41172) );
  XNOR U40953 ( .A(p_input[2644]), .B(n41173), .Z(n40306) );
  AND U40954 ( .A(n767), .B(n41174), .Z(n41173) );
  XOR U40955 ( .A(p_input[2676]), .B(p_input[2644]), .Z(n41174) );
  XNOR U40956 ( .A(n40303), .B(n41169), .Z(n41171) );
  XOR U40957 ( .A(n41175), .B(n41176), .Z(n40303) );
  AND U40958 ( .A(n764), .B(n41177), .Z(n41176) );
  XOR U40959 ( .A(p_input[2612]), .B(p_input[2580]), .Z(n41177) );
  XOR U40960 ( .A(n41178), .B(n41179), .Z(n41169) );
  AND U40961 ( .A(n41180), .B(n41181), .Z(n41179) );
  XOR U40962 ( .A(n41178), .B(n40318), .Z(n41181) );
  XNOR U40963 ( .A(p_input[2643]), .B(n41182), .Z(n40318) );
  AND U40964 ( .A(n767), .B(n41183), .Z(n41182) );
  XOR U40965 ( .A(p_input[2675]), .B(p_input[2643]), .Z(n41183) );
  XNOR U40966 ( .A(n40315), .B(n41178), .Z(n41180) );
  XOR U40967 ( .A(n41184), .B(n41185), .Z(n40315) );
  AND U40968 ( .A(n764), .B(n41186), .Z(n41185) );
  XOR U40969 ( .A(p_input[2611]), .B(p_input[2579]), .Z(n41186) );
  XOR U40970 ( .A(n41187), .B(n41188), .Z(n41178) );
  AND U40971 ( .A(n41189), .B(n41190), .Z(n41188) );
  XOR U40972 ( .A(n41187), .B(n40330), .Z(n41190) );
  XNOR U40973 ( .A(p_input[2642]), .B(n41191), .Z(n40330) );
  AND U40974 ( .A(n767), .B(n41192), .Z(n41191) );
  XOR U40975 ( .A(p_input[2674]), .B(p_input[2642]), .Z(n41192) );
  XNOR U40976 ( .A(n40327), .B(n41187), .Z(n41189) );
  XOR U40977 ( .A(n41193), .B(n41194), .Z(n40327) );
  AND U40978 ( .A(n764), .B(n41195), .Z(n41194) );
  XOR U40979 ( .A(p_input[2610]), .B(p_input[2578]), .Z(n41195) );
  XOR U40980 ( .A(n41196), .B(n41197), .Z(n41187) );
  AND U40981 ( .A(n41198), .B(n41199), .Z(n41197) );
  XOR U40982 ( .A(n41196), .B(n40342), .Z(n41199) );
  XNOR U40983 ( .A(p_input[2641]), .B(n41200), .Z(n40342) );
  AND U40984 ( .A(n767), .B(n41201), .Z(n41200) );
  XOR U40985 ( .A(p_input[2673]), .B(p_input[2641]), .Z(n41201) );
  XNOR U40986 ( .A(n40339), .B(n41196), .Z(n41198) );
  XOR U40987 ( .A(n41202), .B(n41203), .Z(n40339) );
  AND U40988 ( .A(n764), .B(n41204), .Z(n41203) );
  XOR U40989 ( .A(p_input[2609]), .B(p_input[2577]), .Z(n41204) );
  XOR U40990 ( .A(n41205), .B(n41206), .Z(n41196) );
  AND U40991 ( .A(n41207), .B(n41208), .Z(n41206) );
  XOR U40992 ( .A(n41205), .B(n40354), .Z(n41208) );
  XNOR U40993 ( .A(p_input[2640]), .B(n41209), .Z(n40354) );
  AND U40994 ( .A(n767), .B(n41210), .Z(n41209) );
  XOR U40995 ( .A(p_input[2672]), .B(p_input[2640]), .Z(n41210) );
  XNOR U40996 ( .A(n40351), .B(n41205), .Z(n41207) );
  XOR U40997 ( .A(n41211), .B(n41212), .Z(n40351) );
  AND U40998 ( .A(n764), .B(n41213), .Z(n41212) );
  XOR U40999 ( .A(p_input[2608]), .B(p_input[2576]), .Z(n41213) );
  XOR U41000 ( .A(n41214), .B(n41215), .Z(n41205) );
  AND U41001 ( .A(n41216), .B(n41217), .Z(n41215) );
  XOR U41002 ( .A(n41214), .B(n40366), .Z(n41217) );
  XNOR U41003 ( .A(p_input[2639]), .B(n41218), .Z(n40366) );
  AND U41004 ( .A(n767), .B(n41219), .Z(n41218) );
  XOR U41005 ( .A(p_input[2671]), .B(p_input[2639]), .Z(n41219) );
  XNOR U41006 ( .A(n40363), .B(n41214), .Z(n41216) );
  XOR U41007 ( .A(n41220), .B(n41221), .Z(n40363) );
  AND U41008 ( .A(n764), .B(n41222), .Z(n41221) );
  XOR U41009 ( .A(p_input[2607]), .B(p_input[2575]), .Z(n41222) );
  XOR U41010 ( .A(n41223), .B(n41224), .Z(n41214) );
  AND U41011 ( .A(n41225), .B(n41226), .Z(n41224) );
  XOR U41012 ( .A(n41223), .B(n40378), .Z(n41226) );
  XNOR U41013 ( .A(p_input[2638]), .B(n41227), .Z(n40378) );
  AND U41014 ( .A(n767), .B(n41228), .Z(n41227) );
  XOR U41015 ( .A(p_input[2670]), .B(p_input[2638]), .Z(n41228) );
  XNOR U41016 ( .A(n40375), .B(n41223), .Z(n41225) );
  XOR U41017 ( .A(n41229), .B(n41230), .Z(n40375) );
  AND U41018 ( .A(n764), .B(n41231), .Z(n41230) );
  XOR U41019 ( .A(p_input[2606]), .B(p_input[2574]), .Z(n41231) );
  XOR U41020 ( .A(n41232), .B(n41233), .Z(n41223) );
  AND U41021 ( .A(n41234), .B(n41235), .Z(n41233) );
  XOR U41022 ( .A(n41232), .B(n40390), .Z(n41235) );
  XNOR U41023 ( .A(p_input[2637]), .B(n41236), .Z(n40390) );
  AND U41024 ( .A(n767), .B(n41237), .Z(n41236) );
  XOR U41025 ( .A(p_input[2669]), .B(p_input[2637]), .Z(n41237) );
  XNOR U41026 ( .A(n40387), .B(n41232), .Z(n41234) );
  XOR U41027 ( .A(n41238), .B(n41239), .Z(n40387) );
  AND U41028 ( .A(n764), .B(n41240), .Z(n41239) );
  XOR U41029 ( .A(p_input[2605]), .B(p_input[2573]), .Z(n41240) );
  XOR U41030 ( .A(n41241), .B(n41242), .Z(n41232) );
  AND U41031 ( .A(n41243), .B(n41244), .Z(n41242) );
  XOR U41032 ( .A(n41241), .B(n40402), .Z(n41244) );
  XNOR U41033 ( .A(p_input[2636]), .B(n41245), .Z(n40402) );
  AND U41034 ( .A(n767), .B(n41246), .Z(n41245) );
  XOR U41035 ( .A(p_input[2668]), .B(p_input[2636]), .Z(n41246) );
  XNOR U41036 ( .A(n40399), .B(n41241), .Z(n41243) );
  XOR U41037 ( .A(n41247), .B(n41248), .Z(n40399) );
  AND U41038 ( .A(n764), .B(n41249), .Z(n41248) );
  XOR U41039 ( .A(p_input[2604]), .B(p_input[2572]), .Z(n41249) );
  XOR U41040 ( .A(n41250), .B(n41251), .Z(n41241) );
  AND U41041 ( .A(n41252), .B(n41253), .Z(n41251) );
  XOR U41042 ( .A(n41250), .B(n40414), .Z(n41253) );
  XNOR U41043 ( .A(p_input[2635]), .B(n41254), .Z(n40414) );
  AND U41044 ( .A(n767), .B(n41255), .Z(n41254) );
  XOR U41045 ( .A(p_input[2667]), .B(p_input[2635]), .Z(n41255) );
  XNOR U41046 ( .A(n40411), .B(n41250), .Z(n41252) );
  XOR U41047 ( .A(n41256), .B(n41257), .Z(n40411) );
  AND U41048 ( .A(n764), .B(n41258), .Z(n41257) );
  XOR U41049 ( .A(p_input[2603]), .B(p_input[2571]), .Z(n41258) );
  XOR U41050 ( .A(n41259), .B(n41260), .Z(n41250) );
  AND U41051 ( .A(n41261), .B(n41262), .Z(n41260) );
  XOR U41052 ( .A(n41259), .B(n40426), .Z(n41262) );
  XNOR U41053 ( .A(p_input[2634]), .B(n41263), .Z(n40426) );
  AND U41054 ( .A(n767), .B(n41264), .Z(n41263) );
  XOR U41055 ( .A(p_input[2666]), .B(p_input[2634]), .Z(n41264) );
  XNOR U41056 ( .A(n40423), .B(n41259), .Z(n41261) );
  XOR U41057 ( .A(n41265), .B(n41266), .Z(n40423) );
  AND U41058 ( .A(n764), .B(n41267), .Z(n41266) );
  XOR U41059 ( .A(p_input[2602]), .B(p_input[2570]), .Z(n41267) );
  XOR U41060 ( .A(n41268), .B(n41269), .Z(n41259) );
  AND U41061 ( .A(n41270), .B(n41271), .Z(n41269) );
  XOR U41062 ( .A(n41268), .B(n40438), .Z(n41271) );
  XNOR U41063 ( .A(p_input[2633]), .B(n41272), .Z(n40438) );
  AND U41064 ( .A(n767), .B(n41273), .Z(n41272) );
  XOR U41065 ( .A(p_input[2665]), .B(p_input[2633]), .Z(n41273) );
  XNOR U41066 ( .A(n40435), .B(n41268), .Z(n41270) );
  XOR U41067 ( .A(n41274), .B(n41275), .Z(n40435) );
  AND U41068 ( .A(n764), .B(n41276), .Z(n41275) );
  XOR U41069 ( .A(p_input[2601]), .B(p_input[2569]), .Z(n41276) );
  XOR U41070 ( .A(n41277), .B(n41278), .Z(n41268) );
  AND U41071 ( .A(n41279), .B(n41280), .Z(n41278) );
  XOR U41072 ( .A(n41277), .B(n40450), .Z(n41280) );
  XNOR U41073 ( .A(p_input[2632]), .B(n41281), .Z(n40450) );
  AND U41074 ( .A(n767), .B(n41282), .Z(n41281) );
  XOR U41075 ( .A(p_input[2664]), .B(p_input[2632]), .Z(n41282) );
  XNOR U41076 ( .A(n40447), .B(n41277), .Z(n41279) );
  XOR U41077 ( .A(n41283), .B(n41284), .Z(n40447) );
  AND U41078 ( .A(n764), .B(n41285), .Z(n41284) );
  XOR U41079 ( .A(p_input[2600]), .B(p_input[2568]), .Z(n41285) );
  XOR U41080 ( .A(n41286), .B(n41287), .Z(n41277) );
  AND U41081 ( .A(n41288), .B(n41289), .Z(n41287) );
  XOR U41082 ( .A(n41286), .B(n40462), .Z(n41289) );
  XNOR U41083 ( .A(p_input[2631]), .B(n41290), .Z(n40462) );
  AND U41084 ( .A(n767), .B(n41291), .Z(n41290) );
  XOR U41085 ( .A(p_input[2663]), .B(p_input[2631]), .Z(n41291) );
  XNOR U41086 ( .A(n40459), .B(n41286), .Z(n41288) );
  XOR U41087 ( .A(n41292), .B(n41293), .Z(n40459) );
  AND U41088 ( .A(n764), .B(n41294), .Z(n41293) );
  XOR U41089 ( .A(p_input[2599]), .B(p_input[2567]), .Z(n41294) );
  XOR U41090 ( .A(n41295), .B(n41296), .Z(n41286) );
  AND U41091 ( .A(n41297), .B(n41298), .Z(n41296) );
  XOR U41092 ( .A(n41295), .B(n40474), .Z(n41298) );
  XNOR U41093 ( .A(p_input[2630]), .B(n41299), .Z(n40474) );
  AND U41094 ( .A(n767), .B(n41300), .Z(n41299) );
  XOR U41095 ( .A(p_input[2662]), .B(p_input[2630]), .Z(n41300) );
  XNOR U41096 ( .A(n40471), .B(n41295), .Z(n41297) );
  XOR U41097 ( .A(n41301), .B(n41302), .Z(n40471) );
  AND U41098 ( .A(n764), .B(n41303), .Z(n41302) );
  XOR U41099 ( .A(p_input[2598]), .B(p_input[2566]), .Z(n41303) );
  XOR U41100 ( .A(n41304), .B(n41305), .Z(n41295) );
  AND U41101 ( .A(n41306), .B(n41307), .Z(n41305) );
  XOR U41102 ( .A(n41304), .B(n40486), .Z(n41307) );
  XNOR U41103 ( .A(p_input[2629]), .B(n41308), .Z(n40486) );
  AND U41104 ( .A(n767), .B(n41309), .Z(n41308) );
  XOR U41105 ( .A(p_input[2661]), .B(p_input[2629]), .Z(n41309) );
  XNOR U41106 ( .A(n40483), .B(n41304), .Z(n41306) );
  XOR U41107 ( .A(n41310), .B(n41311), .Z(n40483) );
  AND U41108 ( .A(n764), .B(n41312), .Z(n41311) );
  XOR U41109 ( .A(p_input[2597]), .B(p_input[2565]), .Z(n41312) );
  XOR U41110 ( .A(n41313), .B(n41314), .Z(n41304) );
  AND U41111 ( .A(n41315), .B(n41316), .Z(n41314) );
  XOR U41112 ( .A(n41313), .B(n40498), .Z(n41316) );
  XNOR U41113 ( .A(p_input[2628]), .B(n41317), .Z(n40498) );
  AND U41114 ( .A(n767), .B(n41318), .Z(n41317) );
  XOR U41115 ( .A(p_input[2660]), .B(p_input[2628]), .Z(n41318) );
  XNOR U41116 ( .A(n40495), .B(n41313), .Z(n41315) );
  XOR U41117 ( .A(n41319), .B(n41320), .Z(n40495) );
  AND U41118 ( .A(n764), .B(n41321), .Z(n41320) );
  XOR U41119 ( .A(p_input[2596]), .B(p_input[2564]), .Z(n41321) );
  XOR U41120 ( .A(n41322), .B(n41323), .Z(n41313) );
  AND U41121 ( .A(n41324), .B(n41325), .Z(n41323) );
  XOR U41122 ( .A(n41322), .B(n40510), .Z(n41325) );
  XNOR U41123 ( .A(p_input[2627]), .B(n41326), .Z(n40510) );
  AND U41124 ( .A(n767), .B(n41327), .Z(n41326) );
  XOR U41125 ( .A(p_input[2659]), .B(p_input[2627]), .Z(n41327) );
  XNOR U41126 ( .A(n40507), .B(n41322), .Z(n41324) );
  XOR U41127 ( .A(n41328), .B(n41329), .Z(n40507) );
  AND U41128 ( .A(n764), .B(n41330), .Z(n41329) );
  XOR U41129 ( .A(p_input[2595]), .B(p_input[2563]), .Z(n41330) );
  XOR U41130 ( .A(n41331), .B(n41332), .Z(n41322) );
  AND U41131 ( .A(n41333), .B(n41334), .Z(n41332) );
  XOR U41132 ( .A(n41331), .B(n40522), .Z(n41334) );
  XNOR U41133 ( .A(p_input[2626]), .B(n41335), .Z(n40522) );
  AND U41134 ( .A(n767), .B(n41336), .Z(n41335) );
  XOR U41135 ( .A(p_input[2658]), .B(p_input[2626]), .Z(n41336) );
  XNOR U41136 ( .A(n40519), .B(n41331), .Z(n41333) );
  XOR U41137 ( .A(n41337), .B(n41338), .Z(n40519) );
  AND U41138 ( .A(n764), .B(n41339), .Z(n41338) );
  XOR U41139 ( .A(p_input[2594]), .B(p_input[2562]), .Z(n41339) );
  XOR U41140 ( .A(n41340), .B(n41341), .Z(n41331) );
  AND U41141 ( .A(n41342), .B(n41343), .Z(n41341) );
  XNOR U41142 ( .A(n41344), .B(n40535), .Z(n41343) );
  XNOR U41143 ( .A(p_input[2625]), .B(n41345), .Z(n40535) );
  AND U41144 ( .A(n767), .B(n41346), .Z(n41345) );
  XNOR U41145 ( .A(p_input[2657]), .B(n41347), .Z(n41346) );
  IV U41146 ( .A(p_input[2625]), .Z(n41347) );
  XNOR U41147 ( .A(n40532), .B(n41340), .Z(n41342) );
  XNOR U41148 ( .A(p_input[2561]), .B(n41348), .Z(n40532) );
  AND U41149 ( .A(n764), .B(n41349), .Z(n41348) );
  XOR U41150 ( .A(p_input[2593]), .B(p_input[2561]), .Z(n41349) );
  IV U41151 ( .A(n41344), .Z(n41340) );
  AND U41152 ( .A(n41070), .B(n41073), .Z(n41344) );
  XOR U41153 ( .A(p_input[2624]), .B(n41350), .Z(n41073) );
  AND U41154 ( .A(n767), .B(n41351), .Z(n41350) );
  XOR U41155 ( .A(p_input[2656]), .B(p_input[2624]), .Z(n41351) );
  XOR U41156 ( .A(n41352), .B(n41353), .Z(n767) );
  AND U41157 ( .A(n41354), .B(n41355), .Z(n41353) );
  XNOR U41158 ( .A(p_input[2687]), .B(n41352), .Z(n41355) );
  XOR U41159 ( .A(n41352), .B(p_input[2655]), .Z(n41354) );
  XOR U41160 ( .A(n41356), .B(n41357), .Z(n41352) );
  AND U41161 ( .A(n41358), .B(n41359), .Z(n41357) );
  XNOR U41162 ( .A(p_input[2686]), .B(n41356), .Z(n41359) );
  XOR U41163 ( .A(n41356), .B(p_input[2654]), .Z(n41358) );
  XOR U41164 ( .A(n41360), .B(n41361), .Z(n41356) );
  AND U41165 ( .A(n41362), .B(n41363), .Z(n41361) );
  XNOR U41166 ( .A(p_input[2685]), .B(n41360), .Z(n41363) );
  XOR U41167 ( .A(n41360), .B(p_input[2653]), .Z(n41362) );
  XOR U41168 ( .A(n41364), .B(n41365), .Z(n41360) );
  AND U41169 ( .A(n41366), .B(n41367), .Z(n41365) );
  XNOR U41170 ( .A(p_input[2684]), .B(n41364), .Z(n41367) );
  XOR U41171 ( .A(n41364), .B(p_input[2652]), .Z(n41366) );
  XOR U41172 ( .A(n41368), .B(n41369), .Z(n41364) );
  AND U41173 ( .A(n41370), .B(n41371), .Z(n41369) );
  XNOR U41174 ( .A(p_input[2683]), .B(n41368), .Z(n41371) );
  XOR U41175 ( .A(n41368), .B(p_input[2651]), .Z(n41370) );
  XOR U41176 ( .A(n41372), .B(n41373), .Z(n41368) );
  AND U41177 ( .A(n41374), .B(n41375), .Z(n41373) );
  XNOR U41178 ( .A(p_input[2682]), .B(n41372), .Z(n41375) );
  XOR U41179 ( .A(n41372), .B(p_input[2650]), .Z(n41374) );
  XOR U41180 ( .A(n41376), .B(n41377), .Z(n41372) );
  AND U41181 ( .A(n41378), .B(n41379), .Z(n41377) );
  XNOR U41182 ( .A(p_input[2681]), .B(n41376), .Z(n41379) );
  XOR U41183 ( .A(n41376), .B(p_input[2649]), .Z(n41378) );
  XOR U41184 ( .A(n41380), .B(n41381), .Z(n41376) );
  AND U41185 ( .A(n41382), .B(n41383), .Z(n41381) );
  XNOR U41186 ( .A(p_input[2680]), .B(n41380), .Z(n41383) );
  XOR U41187 ( .A(n41380), .B(p_input[2648]), .Z(n41382) );
  XOR U41188 ( .A(n41384), .B(n41385), .Z(n41380) );
  AND U41189 ( .A(n41386), .B(n41387), .Z(n41385) );
  XNOR U41190 ( .A(p_input[2679]), .B(n41384), .Z(n41387) );
  XOR U41191 ( .A(n41384), .B(p_input[2647]), .Z(n41386) );
  XOR U41192 ( .A(n41388), .B(n41389), .Z(n41384) );
  AND U41193 ( .A(n41390), .B(n41391), .Z(n41389) );
  XNOR U41194 ( .A(p_input[2678]), .B(n41388), .Z(n41391) );
  XOR U41195 ( .A(n41388), .B(p_input[2646]), .Z(n41390) );
  XOR U41196 ( .A(n41392), .B(n41393), .Z(n41388) );
  AND U41197 ( .A(n41394), .B(n41395), .Z(n41393) );
  XNOR U41198 ( .A(p_input[2677]), .B(n41392), .Z(n41395) );
  XOR U41199 ( .A(n41392), .B(p_input[2645]), .Z(n41394) );
  XOR U41200 ( .A(n41396), .B(n41397), .Z(n41392) );
  AND U41201 ( .A(n41398), .B(n41399), .Z(n41397) );
  XNOR U41202 ( .A(p_input[2676]), .B(n41396), .Z(n41399) );
  XOR U41203 ( .A(n41396), .B(p_input[2644]), .Z(n41398) );
  XOR U41204 ( .A(n41400), .B(n41401), .Z(n41396) );
  AND U41205 ( .A(n41402), .B(n41403), .Z(n41401) );
  XNOR U41206 ( .A(p_input[2675]), .B(n41400), .Z(n41403) );
  XOR U41207 ( .A(n41400), .B(p_input[2643]), .Z(n41402) );
  XOR U41208 ( .A(n41404), .B(n41405), .Z(n41400) );
  AND U41209 ( .A(n41406), .B(n41407), .Z(n41405) );
  XNOR U41210 ( .A(p_input[2674]), .B(n41404), .Z(n41407) );
  XOR U41211 ( .A(n41404), .B(p_input[2642]), .Z(n41406) );
  XOR U41212 ( .A(n41408), .B(n41409), .Z(n41404) );
  AND U41213 ( .A(n41410), .B(n41411), .Z(n41409) );
  XNOR U41214 ( .A(p_input[2673]), .B(n41408), .Z(n41411) );
  XOR U41215 ( .A(n41408), .B(p_input[2641]), .Z(n41410) );
  XOR U41216 ( .A(n41412), .B(n41413), .Z(n41408) );
  AND U41217 ( .A(n41414), .B(n41415), .Z(n41413) );
  XNOR U41218 ( .A(p_input[2672]), .B(n41412), .Z(n41415) );
  XOR U41219 ( .A(n41412), .B(p_input[2640]), .Z(n41414) );
  XOR U41220 ( .A(n41416), .B(n41417), .Z(n41412) );
  AND U41221 ( .A(n41418), .B(n41419), .Z(n41417) );
  XNOR U41222 ( .A(p_input[2671]), .B(n41416), .Z(n41419) );
  XOR U41223 ( .A(n41416), .B(p_input[2639]), .Z(n41418) );
  XOR U41224 ( .A(n41420), .B(n41421), .Z(n41416) );
  AND U41225 ( .A(n41422), .B(n41423), .Z(n41421) );
  XNOR U41226 ( .A(p_input[2670]), .B(n41420), .Z(n41423) );
  XOR U41227 ( .A(n41420), .B(p_input[2638]), .Z(n41422) );
  XOR U41228 ( .A(n41424), .B(n41425), .Z(n41420) );
  AND U41229 ( .A(n41426), .B(n41427), .Z(n41425) );
  XNOR U41230 ( .A(p_input[2669]), .B(n41424), .Z(n41427) );
  XOR U41231 ( .A(n41424), .B(p_input[2637]), .Z(n41426) );
  XOR U41232 ( .A(n41428), .B(n41429), .Z(n41424) );
  AND U41233 ( .A(n41430), .B(n41431), .Z(n41429) );
  XNOR U41234 ( .A(p_input[2668]), .B(n41428), .Z(n41431) );
  XOR U41235 ( .A(n41428), .B(p_input[2636]), .Z(n41430) );
  XOR U41236 ( .A(n41432), .B(n41433), .Z(n41428) );
  AND U41237 ( .A(n41434), .B(n41435), .Z(n41433) );
  XNOR U41238 ( .A(p_input[2667]), .B(n41432), .Z(n41435) );
  XOR U41239 ( .A(n41432), .B(p_input[2635]), .Z(n41434) );
  XOR U41240 ( .A(n41436), .B(n41437), .Z(n41432) );
  AND U41241 ( .A(n41438), .B(n41439), .Z(n41437) );
  XNOR U41242 ( .A(p_input[2666]), .B(n41436), .Z(n41439) );
  XOR U41243 ( .A(n41436), .B(p_input[2634]), .Z(n41438) );
  XOR U41244 ( .A(n41440), .B(n41441), .Z(n41436) );
  AND U41245 ( .A(n41442), .B(n41443), .Z(n41441) );
  XNOR U41246 ( .A(p_input[2665]), .B(n41440), .Z(n41443) );
  XOR U41247 ( .A(n41440), .B(p_input[2633]), .Z(n41442) );
  XOR U41248 ( .A(n41444), .B(n41445), .Z(n41440) );
  AND U41249 ( .A(n41446), .B(n41447), .Z(n41445) );
  XNOR U41250 ( .A(p_input[2664]), .B(n41444), .Z(n41447) );
  XOR U41251 ( .A(n41444), .B(p_input[2632]), .Z(n41446) );
  XOR U41252 ( .A(n41448), .B(n41449), .Z(n41444) );
  AND U41253 ( .A(n41450), .B(n41451), .Z(n41449) );
  XNOR U41254 ( .A(p_input[2663]), .B(n41448), .Z(n41451) );
  XOR U41255 ( .A(n41448), .B(p_input[2631]), .Z(n41450) );
  XOR U41256 ( .A(n41452), .B(n41453), .Z(n41448) );
  AND U41257 ( .A(n41454), .B(n41455), .Z(n41453) );
  XNOR U41258 ( .A(p_input[2662]), .B(n41452), .Z(n41455) );
  XOR U41259 ( .A(n41452), .B(p_input[2630]), .Z(n41454) );
  XOR U41260 ( .A(n41456), .B(n41457), .Z(n41452) );
  AND U41261 ( .A(n41458), .B(n41459), .Z(n41457) );
  XNOR U41262 ( .A(p_input[2661]), .B(n41456), .Z(n41459) );
  XOR U41263 ( .A(n41456), .B(p_input[2629]), .Z(n41458) );
  XOR U41264 ( .A(n41460), .B(n41461), .Z(n41456) );
  AND U41265 ( .A(n41462), .B(n41463), .Z(n41461) );
  XNOR U41266 ( .A(p_input[2660]), .B(n41460), .Z(n41463) );
  XOR U41267 ( .A(n41460), .B(p_input[2628]), .Z(n41462) );
  XOR U41268 ( .A(n41464), .B(n41465), .Z(n41460) );
  AND U41269 ( .A(n41466), .B(n41467), .Z(n41465) );
  XNOR U41270 ( .A(p_input[2659]), .B(n41464), .Z(n41467) );
  XOR U41271 ( .A(n41464), .B(p_input[2627]), .Z(n41466) );
  XOR U41272 ( .A(n41468), .B(n41469), .Z(n41464) );
  AND U41273 ( .A(n41470), .B(n41471), .Z(n41469) );
  XNOR U41274 ( .A(p_input[2658]), .B(n41468), .Z(n41471) );
  XOR U41275 ( .A(n41468), .B(p_input[2626]), .Z(n41470) );
  XNOR U41276 ( .A(n41472), .B(n41473), .Z(n41468) );
  AND U41277 ( .A(n41474), .B(n41475), .Z(n41473) );
  XOR U41278 ( .A(p_input[2657]), .B(n41472), .Z(n41475) );
  XNOR U41279 ( .A(p_input[2625]), .B(n41472), .Z(n41474) );
  AND U41280 ( .A(p_input[2656]), .B(n41476), .Z(n41472) );
  IV U41281 ( .A(p_input[2624]), .Z(n41476) );
  XNOR U41282 ( .A(p_input[2560]), .B(n41477), .Z(n41070) );
  AND U41283 ( .A(n764), .B(n41478), .Z(n41477) );
  XOR U41284 ( .A(p_input[2592]), .B(p_input[2560]), .Z(n41478) );
  XOR U41285 ( .A(n41479), .B(n41480), .Z(n764) );
  AND U41286 ( .A(n41481), .B(n41482), .Z(n41480) );
  XNOR U41287 ( .A(p_input[2623]), .B(n41479), .Z(n41482) );
  XOR U41288 ( .A(n41479), .B(p_input[2591]), .Z(n41481) );
  XOR U41289 ( .A(n41483), .B(n41484), .Z(n41479) );
  AND U41290 ( .A(n41485), .B(n41486), .Z(n41484) );
  XNOR U41291 ( .A(p_input[2622]), .B(n41483), .Z(n41486) );
  XNOR U41292 ( .A(n41483), .B(n41085), .Z(n41485) );
  IV U41293 ( .A(p_input[2590]), .Z(n41085) );
  XOR U41294 ( .A(n41487), .B(n41488), .Z(n41483) );
  AND U41295 ( .A(n41489), .B(n41490), .Z(n41488) );
  XNOR U41296 ( .A(p_input[2621]), .B(n41487), .Z(n41490) );
  XNOR U41297 ( .A(n41487), .B(n41094), .Z(n41489) );
  IV U41298 ( .A(p_input[2589]), .Z(n41094) );
  XOR U41299 ( .A(n41491), .B(n41492), .Z(n41487) );
  AND U41300 ( .A(n41493), .B(n41494), .Z(n41492) );
  XNOR U41301 ( .A(p_input[2620]), .B(n41491), .Z(n41494) );
  XNOR U41302 ( .A(n41491), .B(n41103), .Z(n41493) );
  IV U41303 ( .A(p_input[2588]), .Z(n41103) );
  XOR U41304 ( .A(n41495), .B(n41496), .Z(n41491) );
  AND U41305 ( .A(n41497), .B(n41498), .Z(n41496) );
  XNOR U41306 ( .A(p_input[2619]), .B(n41495), .Z(n41498) );
  XNOR U41307 ( .A(n41495), .B(n41112), .Z(n41497) );
  IV U41308 ( .A(p_input[2587]), .Z(n41112) );
  XOR U41309 ( .A(n41499), .B(n41500), .Z(n41495) );
  AND U41310 ( .A(n41501), .B(n41502), .Z(n41500) );
  XNOR U41311 ( .A(p_input[2618]), .B(n41499), .Z(n41502) );
  XNOR U41312 ( .A(n41499), .B(n41121), .Z(n41501) );
  IV U41313 ( .A(p_input[2586]), .Z(n41121) );
  XOR U41314 ( .A(n41503), .B(n41504), .Z(n41499) );
  AND U41315 ( .A(n41505), .B(n41506), .Z(n41504) );
  XNOR U41316 ( .A(p_input[2617]), .B(n41503), .Z(n41506) );
  XNOR U41317 ( .A(n41503), .B(n41130), .Z(n41505) );
  IV U41318 ( .A(p_input[2585]), .Z(n41130) );
  XOR U41319 ( .A(n41507), .B(n41508), .Z(n41503) );
  AND U41320 ( .A(n41509), .B(n41510), .Z(n41508) );
  XNOR U41321 ( .A(p_input[2616]), .B(n41507), .Z(n41510) );
  XNOR U41322 ( .A(n41507), .B(n41139), .Z(n41509) );
  IV U41323 ( .A(p_input[2584]), .Z(n41139) );
  XOR U41324 ( .A(n41511), .B(n41512), .Z(n41507) );
  AND U41325 ( .A(n41513), .B(n41514), .Z(n41512) );
  XNOR U41326 ( .A(p_input[2615]), .B(n41511), .Z(n41514) );
  XNOR U41327 ( .A(n41511), .B(n41148), .Z(n41513) );
  IV U41328 ( .A(p_input[2583]), .Z(n41148) );
  XOR U41329 ( .A(n41515), .B(n41516), .Z(n41511) );
  AND U41330 ( .A(n41517), .B(n41518), .Z(n41516) );
  XNOR U41331 ( .A(p_input[2614]), .B(n41515), .Z(n41518) );
  XNOR U41332 ( .A(n41515), .B(n41157), .Z(n41517) );
  IV U41333 ( .A(p_input[2582]), .Z(n41157) );
  XOR U41334 ( .A(n41519), .B(n41520), .Z(n41515) );
  AND U41335 ( .A(n41521), .B(n41522), .Z(n41520) );
  XNOR U41336 ( .A(p_input[2613]), .B(n41519), .Z(n41522) );
  XNOR U41337 ( .A(n41519), .B(n41166), .Z(n41521) );
  IV U41338 ( .A(p_input[2581]), .Z(n41166) );
  XOR U41339 ( .A(n41523), .B(n41524), .Z(n41519) );
  AND U41340 ( .A(n41525), .B(n41526), .Z(n41524) );
  XNOR U41341 ( .A(p_input[2612]), .B(n41523), .Z(n41526) );
  XNOR U41342 ( .A(n41523), .B(n41175), .Z(n41525) );
  IV U41343 ( .A(p_input[2580]), .Z(n41175) );
  XOR U41344 ( .A(n41527), .B(n41528), .Z(n41523) );
  AND U41345 ( .A(n41529), .B(n41530), .Z(n41528) );
  XNOR U41346 ( .A(p_input[2611]), .B(n41527), .Z(n41530) );
  XNOR U41347 ( .A(n41527), .B(n41184), .Z(n41529) );
  IV U41348 ( .A(p_input[2579]), .Z(n41184) );
  XOR U41349 ( .A(n41531), .B(n41532), .Z(n41527) );
  AND U41350 ( .A(n41533), .B(n41534), .Z(n41532) );
  XNOR U41351 ( .A(p_input[2610]), .B(n41531), .Z(n41534) );
  XNOR U41352 ( .A(n41531), .B(n41193), .Z(n41533) );
  IV U41353 ( .A(p_input[2578]), .Z(n41193) );
  XOR U41354 ( .A(n41535), .B(n41536), .Z(n41531) );
  AND U41355 ( .A(n41537), .B(n41538), .Z(n41536) );
  XNOR U41356 ( .A(p_input[2609]), .B(n41535), .Z(n41538) );
  XNOR U41357 ( .A(n41535), .B(n41202), .Z(n41537) );
  IV U41358 ( .A(p_input[2577]), .Z(n41202) );
  XOR U41359 ( .A(n41539), .B(n41540), .Z(n41535) );
  AND U41360 ( .A(n41541), .B(n41542), .Z(n41540) );
  XNOR U41361 ( .A(p_input[2608]), .B(n41539), .Z(n41542) );
  XNOR U41362 ( .A(n41539), .B(n41211), .Z(n41541) );
  IV U41363 ( .A(p_input[2576]), .Z(n41211) );
  XOR U41364 ( .A(n41543), .B(n41544), .Z(n41539) );
  AND U41365 ( .A(n41545), .B(n41546), .Z(n41544) );
  XNOR U41366 ( .A(p_input[2607]), .B(n41543), .Z(n41546) );
  XNOR U41367 ( .A(n41543), .B(n41220), .Z(n41545) );
  IV U41368 ( .A(p_input[2575]), .Z(n41220) );
  XOR U41369 ( .A(n41547), .B(n41548), .Z(n41543) );
  AND U41370 ( .A(n41549), .B(n41550), .Z(n41548) );
  XNOR U41371 ( .A(p_input[2606]), .B(n41547), .Z(n41550) );
  XNOR U41372 ( .A(n41547), .B(n41229), .Z(n41549) );
  IV U41373 ( .A(p_input[2574]), .Z(n41229) );
  XOR U41374 ( .A(n41551), .B(n41552), .Z(n41547) );
  AND U41375 ( .A(n41553), .B(n41554), .Z(n41552) );
  XNOR U41376 ( .A(p_input[2605]), .B(n41551), .Z(n41554) );
  XNOR U41377 ( .A(n41551), .B(n41238), .Z(n41553) );
  IV U41378 ( .A(p_input[2573]), .Z(n41238) );
  XOR U41379 ( .A(n41555), .B(n41556), .Z(n41551) );
  AND U41380 ( .A(n41557), .B(n41558), .Z(n41556) );
  XNOR U41381 ( .A(p_input[2604]), .B(n41555), .Z(n41558) );
  XNOR U41382 ( .A(n41555), .B(n41247), .Z(n41557) );
  IV U41383 ( .A(p_input[2572]), .Z(n41247) );
  XOR U41384 ( .A(n41559), .B(n41560), .Z(n41555) );
  AND U41385 ( .A(n41561), .B(n41562), .Z(n41560) );
  XNOR U41386 ( .A(p_input[2603]), .B(n41559), .Z(n41562) );
  XNOR U41387 ( .A(n41559), .B(n41256), .Z(n41561) );
  IV U41388 ( .A(p_input[2571]), .Z(n41256) );
  XOR U41389 ( .A(n41563), .B(n41564), .Z(n41559) );
  AND U41390 ( .A(n41565), .B(n41566), .Z(n41564) );
  XNOR U41391 ( .A(p_input[2602]), .B(n41563), .Z(n41566) );
  XNOR U41392 ( .A(n41563), .B(n41265), .Z(n41565) );
  IV U41393 ( .A(p_input[2570]), .Z(n41265) );
  XOR U41394 ( .A(n41567), .B(n41568), .Z(n41563) );
  AND U41395 ( .A(n41569), .B(n41570), .Z(n41568) );
  XNOR U41396 ( .A(p_input[2601]), .B(n41567), .Z(n41570) );
  XNOR U41397 ( .A(n41567), .B(n41274), .Z(n41569) );
  IV U41398 ( .A(p_input[2569]), .Z(n41274) );
  XOR U41399 ( .A(n41571), .B(n41572), .Z(n41567) );
  AND U41400 ( .A(n41573), .B(n41574), .Z(n41572) );
  XNOR U41401 ( .A(p_input[2600]), .B(n41571), .Z(n41574) );
  XNOR U41402 ( .A(n41571), .B(n41283), .Z(n41573) );
  IV U41403 ( .A(p_input[2568]), .Z(n41283) );
  XOR U41404 ( .A(n41575), .B(n41576), .Z(n41571) );
  AND U41405 ( .A(n41577), .B(n41578), .Z(n41576) );
  XNOR U41406 ( .A(p_input[2599]), .B(n41575), .Z(n41578) );
  XNOR U41407 ( .A(n41575), .B(n41292), .Z(n41577) );
  IV U41408 ( .A(p_input[2567]), .Z(n41292) );
  XOR U41409 ( .A(n41579), .B(n41580), .Z(n41575) );
  AND U41410 ( .A(n41581), .B(n41582), .Z(n41580) );
  XNOR U41411 ( .A(p_input[2598]), .B(n41579), .Z(n41582) );
  XNOR U41412 ( .A(n41579), .B(n41301), .Z(n41581) );
  IV U41413 ( .A(p_input[2566]), .Z(n41301) );
  XOR U41414 ( .A(n41583), .B(n41584), .Z(n41579) );
  AND U41415 ( .A(n41585), .B(n41586), .Z(n41584) );
  XNOR U41416 ( .A(p_input[2597]), .B(n41583), .Z(n41586) );
  XNOR U41417 ( .A(n41583), .B(n41310), .Z(n41585) );
  IV U41418 ( .A(p_input[2565]), .Z(n41310) );
  XOR U41419 ( .A(n41587), .B(n41588), .Z(n41583) );
  AND U41420 ( .A(n41589), .B(n41590), .Z(n41588) );
  XNOR U41421 ( .A(p_input[2596]), .B(n41587), .Z(n41590) );
  XNOR U41422 ( .A(n41587), .B(n41319), .Z(n41589) );
  IV U41423 ( .A(p_input[2564]), .Z(n41319) );
  XOR U41424 ( .A(n41591), .B(n41592), .Z(n41587) );
  AND U41425 ( .A(n41593), .B(n41594), .Z(n41592) );
  XNOR U41426 ( .A(p_input[2595]), .B(n41591), .Z(n41594) );
  XNOR U41427 ( .A(n41591), .B(n41328), .Z(n41593) );
  IV U41428 ( .A(p_input[2563]), .Z(n41328) );
  XOR U41429 ( .A(n41595), .B(n41596), .Z(n41591) );
  AND U41430 ( .A(n41597), .B(n41598), .Z(n41596) );
  XNOR U41431 ( .A(p_input[2594]), .B(n41595), .Z(n41598) );
  XNOR U41432 ( .A(n41595), .B(n41337), .Z(n41597) );
  IV U41433 ( .A(p_input[2562]), .Z(n41337) );
  XNOR U41434 ( .A(n41599), .B(n41600), .Z(n41595) );
  AND U41435 ( .A(n41601), .B(n41602), .Z(n41600) );
  XOR U41436 ( .A(p_input[2593]), .B(n41599), .Z(n41602) );
  XNOR U41437 ( .A(p_input[2561]), .B(n41599), .Z(n41601) );
  AND U41438 ( .A(p_input[2592]), .B(n41603), .Z(n41599) );
  IV U41439 ( .A(p_input[2560]), .Z(n41603) );
  XOR U41440 ( .A(n41604), .B(n41605), .Z(n37960) );
  AND U41441 ( .A(n1028), .B(n41606), .Z(n41605) );
  XNOR U41442 ( .A(n41607), .B(n41604), .Z(n41606) );
  XOR U41443 ( .A(n41608), .B(n41609), .Z(n1028) );
  AND U41444 ( .A(n41610), .B(n41611), .Z(n41609) );
  XOR U41445 ( .A(n41608), .B(n37975), .Z(n41611) );
  XOR U41446 ( .A(n41612), .B(n41613), .Z(n37975) );
  AND U41447 ( .A(n891), .B(n41614), .Z(n41613) );
  XOR U41448 ( .A(n41615), .B(n41612), .Z(n41614) );
  XNOR U41449 ( .A(n37972), .B(n41608), .Z(n41610) );
  XOR U41450 ( .A(n41616), .B(n41617), .Z(n37972) );
  AND U41451 ( .A(n888), .B(n41618), .Z(n41617) );
  XOR U41452 ( .A(n41619), .B(n41616), .Z(n41618) );
  XOR U41453 ( .A(n41620), .B(n41621), .Z(n41608) );
  AND U41454 ( .A(n41622), .B(n41623), .Z(n41621) );
  XOR U41455 ( .A(n41620), .B(n37987), .Z(n41623) );
  XOR U41456 ( .A(n41624), .B(n41625), .Z(n37987) );
  AND U41457 ( .A(n891), .B(n41626), .Z(n41625) );
  XOR U41458 ( .A(n41627), .B(n41624), .Z(n41626) );
  XNOR U41459 ( .A(n37984), .B(n41620), .Z(n41622) );
  XOR U41460 ( .A(n41628), .B(n41629), .Z(n37984) );
  AND U41461 ( .A(n888), .B(n41630), .Z(n41629) );
  XOR U41462 ( .A(n41631), .B(n41628), .Z(n41630) );
  XOR U41463 ( .A(n41632), .B(n41633), .Z(n41620) );
  AND U41464 ( .A(n41634), .B(n41635), .Z(n41633) );
  XOR U41465 ( .A(n41632), .B(n37999), .Z(n41635) );
  XOR U41466 ( .A(n41636), .B(n41637), .Z(n37999) );
  AND U41467 ( .A(n891), .B(n41638), .Z(n41637) );
  XOR U41468 ( .A(n41639), .B(n41636), .Z(n41638) );
  XNOR U41469 ( .A(n37996), .B(n41632), .Z(n41634) );
  XOR U41470 ( .A(n41640), .B(n41641), .Z(n37996) );
  AND U41471 ( .A(n888), .B(n41642), .Z(n41641) );
  XOR U41472 ( .A(n41643), .B(n41640), .Z(n41642) );
  XOR U41473 ( .A(n41644), .B(n41645), .Z(n41632) );
  AND U41474 ( .A(n41646), .B(n41647), .Z(n41645) );
  XOR U41475 ( .A(n41644), .B(n38011), .Z(n41647) );
  XOR U41476 ( .A(n41648), .B(n41649), .Z(n38011) );
  AND U41477 ( .A(n891), .B(n41650), .Z(n41649) );
  XOR U41478 ( .A(n41651), .B(n41648), .Z(n41650) );
  XNOR U41479 ( .A(n38008), .B(n41644), .Z(n41646) );
  XOR U41480 ( .A(n41652), .B(n41653), .Z(n38008) );
  AND U41481 ( .A(n888), .B(n41654), .Z(n41653) );
  XOR U41482 ( .A(n41655), .B(n41652), .Z(n41654) );
  XOR U41483 ( .A(n41656), .B(n41657), .Z(n41644) );
  AND U41484 ( .A(n41658), .B(n41659), .Z(n41657) );
  XOR U41485 ( .A(n41656), .B(n38023), .Z(n41659) );
  XOR U41486 ( .A(n41660), .B(n41661), .Z(n38023) );
  AND U41487 ( .A(n891), .B(n41662), .Z(n41661) );
  XOR U41488 ( .A(n41663), .B(n41660), .Z(n41662) );
  XNOR U41489 ( .A(n38020), .B(n41656), .Z(n41658) );
  XOR U41490 ( .A(n41664), .B(n41665), .Z(n38020) );
  AND U41491 ( .A(n888), .B(n41666), .Z(n41665) );
  XOR U41492 ( .A(n41667), .B(n41664), .Z(n41666) );
  XOR U41493 ( .A(n41668), .B(n41669), .Z(n41656) );
  AND U41494 ( .A(n41670), .B(n41671), .Z(n41669) );
  XOR U41495 ( .A(n41668), .B(n38035), .Z(n41671) );
  XOR U41496 ( .A(n41672), .B(n41673), .Z(n38035) );
  AND U41497 ( .A(n891), .B(n41674), .Z(n41673) );
  XOR U41498 ( .A(n41675), .B(n41672), .Z(n41674) );
  XNOR U41499 ( .A(n38032), .B(n41668), .Z(n41670) );
  XOR U41500 ( .A(n41676), .B(n41677), .Z(n38032) );
  AND U41501 ( .A(n888), .B(n41678), .Z(n41677) );
  XOR U41502 ( .A(n41679), .B(n41676), .Z(n41678) );
  XOR U41503 ( .A(n41680), .B(n41681), .Z(n41668) );
  AND U41504 ( .A(n41682), .B(n41683), .Z(n41681) );
  XOR U41505 ( .A(n41680), .B(n38047), .Z(n41683) );
  XOR U41506 ( .A(n41684), .B(n41685), .Z(n38047) );
  AND U41507 ( .A(n891), .B(n41686), .Z(n41685) );
  XOR U41508 ( .A(n41687), .B(n41684), .Z(n41686) );
  XNOR U41509 ( .A(n38044), .B(n41680), .Z(n41682) );
  XOR U41510 ( .A(n41688), .B(n41689), .Z(n38044) );
  AND U41511 ( .A(n888), .B(n41690), .Z(n41689) );
  XOR U41512 ( .A(n41691), .B(n41688), .Z(n41690) );
  XOR U41513 ( .A(n41692), .B(n41693), .Z(n41680) );
  AND U41514 ( .A(n41694), .B(n41695), .Z(n41693) );
  XOR U41515 ( .A(n41692), .B(n38059), .Z(n41695) );
  XOR U41516 ( .A(n41696), .B(n41697), .Z(n38059) );
  AND U41517 ( .A(n891), .B(n41698), .Z(n41697) );
  XOR U41518 ( .A(n41699), .B(n41696), .Z(n41698) );
  XNOR U41519 ( .A(n38056), .B(n41692), .Z(n41694) );
  XOR U41520 ( .A(n41700), .B(n41701), .Z(n38056) );
  AND U41521 ( .A(n888), .B(n41702), .Z(n41701) );
  XOR U41522 ( .A(n41703), .B(n41700), .Z(n41702) );
  XOR U41523 ( .A(n41704), .B(n41705), .Z(n41692) );
  AND U41524 ( .A(n41706), .B(n41707), .Z(n41705) );
  XOR U41525 ( .A(n41704), .B(n38071), .Z(n41707) );
  XOR U41526 ( .A(n41708), .B(n41709), .Z(n38071) );
  AND U41527 ( .A(n891), .B(n41710), .Z(n41709) );
  XOR U41528 ( .A(n41711), .B(n41708), .Z(n41710) );
  XNOR U41529 ( .A(n38068), .B(n41704), .Z(n41706) );
  XOR U41530 ( .A(n41712), .B(n41713), .Z(n38068) );
  AND U41531 ( .A(n888), .B(n41714), .Z(n41713) );
  XOR U41532 ( .A(n41715), .B(n41712), .Z(n41714) );
  XOR U41533 ( .A(n41716), .B(n41717), .Z(n41704) );
  AND U41534 ( .A(n41718), .B(n41719), .Z(n41717) );
  XOR U41535 ( .A(n41716), .B(n38083), .Z(n41719) );
  XOR U41536 ( .A(n41720), .B(n41721), .Z(n38083) );
  AND U41537 ( .A(n891), .B(n41722), .Z(n41721) );
  XOR U41538 ( .A(n41723), .B(n41720), .Z(n41722) );
  XNOR U41539 ( .A(n38080), .B(n41716), .Z(n41718) );
  XOR U41540 ( .A(n41724), .B(n41725), .Z(n38080) );
  AND U41541 ( .A(n888), .B(n41726), .Z(n41725) );
  XOR U41542 ( .A(n41727), .B(n41724), .Z(n41726) );
  XOR U41543 ( .A(n41728), .B(n41729), .Z(n41716) );
  AND U41544 ( .A(n41730), .B(n41731), .Z(n41729) );
  XOR U41545 ( .A(n41728), .B(n38095), .Z(n41731) );
  XOR U41546 ( .A(n41732), .B(n41733), .Z(n38095) );
  AND U41547 ( .A(n891), .B(n41734), .Z(n41733) );
  XOR U41548 ( .A(n41735), .B(n41732), .Z(n41734) );
  XNOR U41549 ( .A(n38092), .B(n41728), .Z(n41730) );
  XOR U41550 ( .A(n41736), .B(n41737), .Z(n38092) );
  AND U41551 ( .A(n888), .B(n41738), .Z(n41737) );
  XOR U41552 ( .A(n41739), .B(n41736), .Z(n41738) );
  XOR U41553 ( .A(n41740), .B(n41741), .Z(n41728) );
  AND U41554 ( .A(n41742), .B(n41743), .Z(n41741) );
  XOR U41555 ( .A(n41740), .B(n38107), .Z(n41743) );
  XOR U41556 ( .A(n41744), .B(n41745), .Z(n38107) );
  AND U41557 ( .A(n891), .B(n41746), .Z(n41745) );
  XOR U41558 ( .A(n41747), .B(n41744), .Z(n41746) );
  XNOR U41559 ( .A(n38104), .B(n41740), .Z(n41742) );
  XOR U41560 ( .A(n41748), .B(n41749), .Z(n38104) );
  AND U41561 ( .A(n888), .B(n41750), .Z(n41749) );
  XOR U41562 ( .A(n41751), .B(n41748), .Z(n41750) );
  XOR U41563 ( .A(n41752), .B(n41753), .Z(n41740) );
  AND U41564 ( .A(n41754), .B(n41755), .Z(n41753) );
  XOR U41565 ( .A(n41752), .B(n38119), .Z(n41755) );
  XOR U41566 ( .A(n41756), .B(n41757), .Z(n38119) );
  AND U41567 ( .A(n891), .B(n41758), .Z(n41757) );
  XOR U41568 ( .A(n41759), .B(n41756), .Z(n41758) );
  XNOR U41569 ( .A(n38116), .B(n41752), .Z(n41754) );
  XOR U41570 ( .A(n41760), .B(n41761), .Z(n38116) );
  AND U41571 ( .A(n888), .B(n41762), .Z(n41761) );
  XOR U41572 ( .A(n41763), .B(n41760), .Z(n41762) );
  XOR U41573 ( .A(n41764), .B(n41765), .Z(n41752) );
  AND U41574 ( .A(n41766), .B(n41767), .Z(n41765) );
  XOR U41575 ( .A(n41764), .B(n38131), .Z(n41767) );
  XOR U41576 ( .A(n41768), .B(n41769), .Z(n38131) );
  AND U41577 ( .A(n891), .B(n41770), .Z(n41769) );
  XOR U41578 ( .A(n41771), .B(n41768), .Z(n41770) );
  XNOR U41579 ( .A(n38128), .B(n41764), .Z(n41766) );
  XOR U41580 ( .A(n41772), .B(n41773), .Z(n38128) );
  AND U41581 ( .A(n888), .B(n41774), .Z(n41773) );
  XOR U41582 ( .A(n41775), .B(n41772), .Z(n41774) );
  XOR U41583 ( .A(n41776), .B(n41777), .Z(n41764) );
  AND U41584 ( .A(n41778), .B(n41779), .Z(n41777) );
  XOR U41585 ( .A(n41776), .B(n38143), .Z(n41779) );
  XOR U41586 ( .A(n41780), .B(n41781), .Z(n38143) );
  AND U41587 ( .A(n891), .B(n41782), .Z(n41781) );
  XOR U41588 ( .A(n41783), .B(n41780), .Z(n41782) );
  XNOR U41589 ( .A(n38140), .B(n41776), .Z(n41778) );
  XOR U41590 ( .A(n41784), .B(n41785), .Z(n38140) );
  AND U41591 ( .A(n888), .B(n41786), .Z(n41785) );
  XOR U41592 ( .A(n41787), .B(n41784), .Z(n41786) );
  XOR U41593 ( .A(n41788), .B(n41789), .Z(n41776) );
  AND U41594 ( .A(n41790), .B(n41791), .Z(n41789) );
  XOR U41595 ( .A(n41788), .B(n38155), .Z(n41791) );
  XOR U41596 ( .A(n41792), .B(n41793), .Z(n38155) );
  AND U41597 ( .A(n891), .B(n41794), .Z(n41793) );
  XOR U41598 ( .A(n41795), .B(n41792), .Z(n41794) );
  XNOR U41599 ( .A(n38152), .B(n41788), .Z(n41790) );
  XOR U41600 ( .A(n41796), .B(n41797), .Z(n38152) );
  AND U41601 ( .A(n888), .B(n41798), .Z(n41797) );
  XOR U41602 ( .A(n41799), .B(n41796), .Z(n41798) );
  XOR U41603 ( .A(n41800), .B(n41801), .Z(n41788) );
  AND U41604 ( .A(n41802), .B(n41803), .Z(n41801) );
  XOR U41605 ( .A(n41800), .B(n38167), .Z(n41803) );
  XOR U41606 ( .A(n41804), .B(n41805), .Z(n38167) );
  AND U41607 ( .A(n891), .B(n41806), .Z(n41805) );
  XOR U41608 ( .A(n41807), .B(n41804), .Z(n41806) );
  XNOR U41609 ( .A(n38164), .B(n41800), .Z(n41802) );
  XOR U41610 ( .A(n41808), .B(n41809), .Z(n38164) );
  AND U41611 ( .A(n888), .B(n41810), .Z(n41809) );
  XOR U41612 ( .A(n41811), .B(n41808), .Z(n41810) );
  XOR U41613 ( .A(n41812), .B(n41813), .Z(n41800) );
  AND U41614 ( .A(n41814), .B(n41815), .Z(n41813) );
  XOR U41615 ( .A(n41812), .B(n38179), .Z(n41815) );
  XOR U41616 ( .A(n41816), .B(n41817), .Z(n38179) );
  AND U41617 ( .A(n891), .B(n41818), .Z(n41817) );
  XOR U41618 ( .A(n41819), .B(n41816), .Z(n41818) );
  XNOR U41619 ( .A(n38176), .B(n41812), .Z(n41814) );
  XOR U41620 ( .A(n41820), .B(n41821), .Z(n38176) );
  AND U41621 ( .A(n888), .B(n41822), .Z(n41821) );
  XOR U41622 ( .A(n41823), .B(n41820), .Z(n41822) );
  XOR U41623 ( .A(n41824), .B(n41825), .Z(n41812) );
  AND U41624 ( .A(n41826), .B(n41827), .Z(n41825) );
  XOR U41625 ( .A(n41824), .B(n38191), .Z(n41827) );
  XOR U41626 ( .A(n41828), .B(n41829), .Z(n38191) );
  AND U41627 ( .A(n891), .B(n41830), .Z(n41829) );
  XOR U41628 ( .A(n41831), .B(n41828), .Z(n41830) );
  XNOR U41629 ( .A(n38188), .B(n41824), .Z(n41826) );
  XOR U41630 ( .A(n41832), .B(n41833), .Z(n38188) );
  AND U41631 ( .A(n888), .B(n41834), .Z(n41833) );
  XOR U41632 ( .A(n41835), .B(n41832), .Z(n41834) );
  XOR U41633 ( .A(n41836), .B(n41837), .Z(n41824) );
  AND U41634 ( .A(n41838), .B(n41839), .Z(n41837) );
  XOR U41635 ( .A(n41836), .B(n38203), .Z(n41839) );
  XOR U41636 ( .A(n41840), .B(n41841), .Z(n38203) );
  AND U41637 ( .A(n891), .B(n41842), .Z(n41841) );
  XOR U41638 ( .A(n41843), .B(n41840), .Z(n41842) );
  XNOR U41639 ( .A(n38200), .B(n41836), .Z(n41838) );
  XOR U41640 ( .A(n41844), .B(n41845), .Z(n38200) );
  AND U41641 ( .A(n888), .B(n41846), .Z(n41845) );
  XOR U41642 ( .A(n41847), .B(n41844), .Z(n41846) );
  XOR U41643 ( .A(n41848), .B(n41849), .Z(n41836) );
  AND U41644 ( .A(n41850), .B(n41851), .Z(n41849) );
  XOR U41645 ( .A(n41848), .B(n38215), .Z(n41851) );
  XOR U41646 ( .A(n41852), .B(n41853), .Z(n38215) );
  AND U41647 ( .A(n891), .B(n41854), .Z(n41853) );
  XOR U41648 ( .A(n41855), .B(n41852), .Z(n41854) );
  XNOR U41649 ( .A(n38212), .B(n41848), .Z(n41850) );
  XOR U41650 ( .A(n41856), .B(n41857), .Z(n38212) );
  AND U41651 ( .A(n888), .B(n41858), .Z(n41857) );
  XOR U41652 ( .A(n41859), .B(n41856), .Z(n41858) );
  XOR U41653 ( .A(n41860), .B(n41861), .Z(n41848) );
  AND U41654 ( .A(n41862), .B(n41863), .Z(n41861) );
  XOR U41655 ( .A(n41860), .B(n38227), .Z(n41863) );
  XOR U41656 ( .A(n41864), .B(n41865), .Z(n38227) );
  AND U41657 ( .A(n891), .B(n41866), .Z(n41865) );
  XOR U41658 ( .A(n41867), .B(n41864), .Z(n41866) );
  XNOR U41659 ( .A(n38224), .B(n41860), .Z(n41862) );
  XOR U41660 ( .A(n41868), .B(n41869), .Z(n38224) );
  AND U41661 ( .A(n888), .B(n41870), .Z(n41869) );
  XOR U41662 ( .A(n41871), .B(n41868), .Z(n41870) );
  XOR U41663 ( .A(n41872), .B(n41873), .Z(n41860) );
  AND U41664 ( .A(n41874), .B(n41875), .Z(n41873) );
  XOR U41665 ( .A(n41872), .B(n38239), .Z(n41875) );
  XOR U41666 ( .A(n41876), .B(n41877), .Z(n38239) );
  AND U41667 ( .A(n891), .B(n41878), .Z(n41877) );
  XOR U41668 ( .A(n41879), .B(n41876), .Z(n41878) );
  XNOR U41669 ( .A(n38236), .B(n41872), .Z(n41874) );
  XOR U41670 ( .A(n41880), .B(n41881), .Z(n38236) );
  AND U41671 ( .A(n888), .B(n41882), .Z(n41881) );
  XOR U41672 ( .A(n41883), .B(n41880), .Z(n41882) );
  XOR U41673 ( .A(n41884), .B(n41885), .Z(n41872) );
  AND U41674 ( .A(n41886), .B(n41887), .Z(n41885) );
  XOR U41675 ( .A(n41884), .B(n38251), .Z(n41887) );
  XOR U41676 ( .A(n41888), .B(n41889), .Z(n38251) );
  AND U41677 ( .A(n891), .B(n41890), .Z(n41889) );
  XOR U41678 ( .A(n41891), .B(n41888), .Z(n41890) );
  XNOR U41679 ( .A(n38248), .B(n41884), .Z(n41886) );
  XOR U41680 ( .A(n41892), .B(n41893), .Z(n38248) );
  AND U41681 ( .A(n888), .B(n41894), .Z(n41893) );
  XOR U41682 ( .A(n41895), .B(n41892), .Z(n41894) );
  XOR U41683 ( .A(n41896), .B(n41897), .Z(n41884) );
  AND U41684 ( .A(n41898), .B(n41899), .Z(n41897) );
  XOR U41685 ( .A(n41896), .B(n38263), .Z(n41899) );
  XOR U41686 ( .A(n41900), .B(n41901), .Z(n38263) );
  AND U41687 ( .A(n891), .B(n41902), .Z(n41901) );
  XOR U41688 ( .A(n41903), .B(n41900), .Z(n41902) );
  XNOR U41689 ( .A(n38260), .B(n41896), .Z(n41898) );
  XOR U41690 ( .A(n41904), .B(n41905), .Z(n38260) );
  AND U41691 ( .A(n888), .B(n41906), .Z(n41905) );
  XOR U41692 ( .A(n41907), .B(n41904), .Z(n41906) );
  XOR U41693 ( .A(n41908), .B(n41909), .Z(n41896) );
  AND U41694 ( .A(n41910), .B(n41911), .Z(n41909) );
  XOR U41695 ( .A(n41908), .B(n38275), .Z(n41911) );
  XOR U41696 ( .A(n41912), .B(n41913), .Z(n38275) );
  AND U41697 ( .A(n891), .B(n41914), .Z(n41913) );
  XOR U41698 ( .A(n41915), .B(n41912), .Z(n41914) );
  XNOR U41699 ( .A(n38272), .B(n41908), .Z(n41910) );
  XOR U41700 ( .A(n41916), .B(n41917), .Z(n38272) );
  AND U41701 ( .A(n888), .B(n41918), .Z(n41917) );
  XOR U41702 ( .A(n41919), .B(n41916), .Z(n41918) );
  XOR U41703 ( .A(n41920), .B(n41921), .Z(n41908) );
  AND U41704 ( .A(n41922), .B(n41923), .Z(n41921) );
  XOR U41705 ( .A(n41920), .B(n38287), .Z(n41923) );
  XOR U41706 ( .A(n41924), .B(n41925), .Z(n38287) );
  AND U41707 ( .A(n891), .B(n41926), .Z(n41925) );
  XOR U41708 ( .A(n41927), .B(n41924), .Z(n41926) );
  XNOR U41709 ( .A(n38284), .B(n41920), .Z(n41922) );
  XOR U41710 ( .A(n41928), .B(n41929), .Z(n38284) );
  AND U41711 ( .A(n888), .B(n41930), .Z(n41929) );
  XOR U41712 ( .A(n41931), .B(n41928), .Z(n41930) );
  XOR U41713 ( .A(n41932), .B(n41933), .Z(n41920) );
  AND U41714 ( .A(n41934), .B(n41935), .Z(n41933) );
  XOR U41715 ( .A(n41932), .B(n38299), .Z(n41935) );
  XOR U41716 ( .A(n41936), .B(n41937), .Z(n38299) );
  AND U41717 ( .A(n891), .B(n41938), .Z(n41937) );
  XOR U41718 ( .A(n41939), .B(n41936), .Z(n41938) );
  XNOR U41719 ( .A(n38296), .B(n41932), .Z(n41934) );
  XOR U41720 ( .A(n41940), .B(n41941), .Z(n38296) );
  AND U41721 ( .A(n888), .B(n41942), .Z(n41941) );
  XOR U41722 ( .A(n41943), .B(n41940), .Z(n41942) );
  XOR U41723 ( .A(n41944), .B(n41945), .Z(n41932) );
  AND U41724 ( .A(n41946), .B(n41947), .Z(n41945) );
  XOR U41725 ( .A(n41944), .B(n38311), .Z(n41947) );
  XOR U41726 ( .A(n41948), .B(n41949), .Z(n38311) );
  AND U41727 ( .A(n891), .B(n41950), .Z(n41949) );
  XOR U41728 ( .A(n41951), .B(n41948), .Z(n41950) );
  XNOR U41729 ( .A(n38308), .B(n41944), .Z(n41946) );
  XOR U41730 ( .A(n41952), .B(n41953), .Z(n38308) );
  AND U41731 ( .A(n888), .B(n41954), .Z(n41953) );
  XOR U41732 ( .A(n41955), .B(n41952), .Z(n41954) );
  XOR U41733 ( .A(n41956), .B(n41957), .Z(n41944) );
  AND U41734 ( .A(n41958), .B(n41959), .Z(n41957) );
  XOR U41735 ( .A(n41956), .B(n38323), .Z(n41959) );
  XOR U41736 ( .A(n41960), .B(n41961), .Z(n38323) );
  AND U41737 ( .A(n891), .B(n41962), .Z(n41961) );
  XOR U41738 ( .A(n41963), .B(n41960), .Z(n41962) );
  XNOR U41739 ( .A(n38320), .B(n41956), .Z(n41958) );
  XOR U41740 ( .A(n41964), .B(n41965), .Z(n38320) );
  AND U41741 ( .A(n888), .B(n41966), .Z(n41965) );
  XOR U41742 ( .A(n41967), .B(n41964), .Z(n41966) );
  XOR U41743 ( .A(n41968), .B(n41969), .Z(n41956) );
  AND U41744 ( .A(n41970), .B(n41971), .Z(n41969) );
  XNOR U41745 ( .A(n41972), .B(n38336), .Z(n41971) );
  XOR U41746 ( .A(n41973), .B(n41974), .Z(n38336) );
  AND U41747 ( .A(n891), .B(n41975), .Z(n41974) );
  XOR U41748 ( .A(n41973), .B(n41976), .Z(n41975) );
  XNOR U41749 ( .A(n38333), .B(n41968), .Z(n41970) );
  XOR U41750 ( .A(n41977), .B(n41978), .Z(n38333) );
  AND U41751 ( .A(n888), .B(n41979), .Z(n41978) );
  XOR U41752 ( .A(n41977), .B(n41980), .Z(n41979) );
  IV U41753 ( .A(n41972), .Z(n41968) );
  AND U41754 ( .A(n41604), .B(n41607), .Z(n41972) );
  XNOR U41755 ( .A(n41981), .B(n41982), .Z(n41607) );
  AND U41756 ( .A(n891), .B(n41983), .Z(n41982) );
  XNOR U41757 ( .A(n41984), .B(n41981), .Z(n41983) );
  XOR U41758 ( .A(n41985), .B(n41986), .Z(n891) );
  AND U41759 ( .A(n41987), .B(n41988), .Z(n41986) );
  XOR U41760 ( .A(n41985), .B(n41615), .Z(n41988) );
  XNOR U41761 ( .A(n41989), .B(n41990), .Z(n41615) );
  AND U41762 ( .A(n41991), .B(n603), .Z(n41990) );
  AND U41763 ( .A(n41989), .B(n41992), .Z(n41991) );
  XNOR U41764 ( .A(n41612), .B(n41985), .Z(n41987) );
  XOR U41765 ( .A(n41993), .B(n41994), .Z(n41612) );
  AND U41766 ( .A(n41995), .B(n601), .Z(n41994) );
  NOR U41767 ( .A(n41993), .B(n41996), .Z(n41995) );
  XOR U41768 ( .A(n41997), .B(n41998), .Z(n41985) );
  AND U41769 ( .A(n41999), .B(n42000), .Z(n41998) );
  XOR U41770 ( .A(n41997), .B(n41627), .Z(n42000) );
  XOR U41771 ( .A(n42001), .B(n42002), .Z(n41627) );
  AND U41772 ( .A(n603), .B(n42003), .Z(n42002) );
  XOR U41773 ( .A(n42004), .B(n42001), .Z(n42003) );
  XNOR U41774 ( .A(n41624), .B(n41997), .Z(n41999) );
  XOR U41775 ( .A(n42005), .B(n42006), .Z(n41624) );
  AND U41776 ( .A(n601), .B(n42007), .Z(n42006) );
  XOR U41777 ( .A(n42008), .B(n42005), .Z(n42007) );
  XOR U41778 ( .A(n42009), .B(n42010), .Z(n41997) );
  AND U41779 ( .A(n42011), .B(n42012), .Z(n42010) );
  XOR U41780 ( .A(n42009), .B(n41639), .Z(n42012) );
  XOR U41781 ( .A(n42013), .B(n42014), .Z(n41639) );
  AND U41782 ( .A(n603), .B(n42015), .Z(n42014) );
  XOR U41783 ( .A(n42016), .B(n42013), .Z(n42015) );
  XNOR U41784 ( .A(n41636), .B(n42009), .Z(n42011) );
  XOR U41785 ( .A(n42017), .B(n42018), .Z(n41636) );
  AND U41786 ( .A(n601), .B(n42019), .Z(n42018) );
  XOR U41787 ( .A(n42020), .B(n42017), .Z(n42019) );
  XOR U41788 ( .A(n42021), .B(n42022), .Z(n42009) );
  AND U41789 ( .A(n42023), .B(n42024), .Z(n42022) );
  XOR U41790 ( .A(n42021), .B(n41651), .Z(n42024) );
  XOR U41791 ( .A(n42025), .B(n42026), .Z(n41651) );
  AND U41792 ( .A(n603), .B(n42027), .Z(n42026) );
  XOR U41793 ( .A(n42028), .B(n42025), .Z(n42027) );
  XNOR U41794 ( .A(n41648), .B(n42021), .Z(n42023) );
  XOR U41795 ( .A(n42029), .B(n42030), .Z(n41648) );
  AND U41796 ( .A(n601), .B(n42031), .Z(n42030) );
  XOR U41797 ( .A(n42032), .B(n42029), .Z(n42031) );
  XOR U41798 ( .A(n42033), .B(n42034), .Z(n42021) );
  AND U41799 ( .A(n42035), .B(n42036), .Z(n42034) );
  XOR U41800 ( .A(n42033), .B(n41663), .Z(n42036) );
  XOR U41801 ( .A(n42037), .B(n42038), .Z(n41663) );
  AND U41802 ( .A(n603), .B(n42039), .Z(n42038) );
  XOR U41803 ( .A(n42040), .B(n42037), .Z(n42039) );
  XNOR U41804 ( .A(n41660), .B(n42033), .Z(n42035) );
  XOR U41805 ( .A(n42041), .B(n42042), .Z(n41660) );
  AND U41806 ( .A(n601), .B(n42043), .Z(n42042) );
  XOR U41807 ( .A(n42044), .B(n42041), .Z(n42043) );
  XOR U41808 ( .A(n42045), .B(n42046), .Z(n42033) );
  AND U41809 ( .A(n42047), .B(n42048), .Z(n42046) );
  XOR U41810 ( .A(n42045), .B(n41675), .Z(n42048) );
  XOR U41811 ( .A(n42049), .B(n42050), .Z(n41675) );
  AND U41812 ( .A(n603), .B(n42051), .Z(n42050) );
  XOR U41813 ( .A(n42052), .B(n42049), .Z(n42051) );
  XNOR U41814 ( .A(n41672), .B(n42045), .Z(n42047) );
  XOR U41815 ( .A(n42053), .B(n42054), .Z(n41672) );
  AND U41816 ( .A(n601), .B(n42055), .Z(n42054) );
  XOR U41817 ( .A(n42056), .B(n42053), .Z(n42055) );
  XOR U41818 ( .A(n42057), .B(n42058), .Z(n42045) );
  AND U41819 ( .A(n42059), .B(n42060), .Z(n42058) );
  XOR U41820 ( .A(n42057), .B(n41687), .Z(n42060) );
  XOR U41821 ( .A(n42061), .B(n42062), .Z(n41687) );
  AND U41822 ( .A(n603), .B(n42063), .Z(n42062) );
  XOR U41823 ( .A(n42064), .B(n42061), .Z(n42063) );
  XNOR U41824 ( .A(n41684), .B(n42057), .Z(n42059) );
  XOR U41825 ( .A(n42065), .B(n42066), .Z(n41684) );
  AND U41826 ( .A(n601), .B(n42067), .Z(n42066) );
  XOR U41827 ( .A(n42068), .B(n42065), .Z(n42067) );
  XOR U41828 ( .A(n42069), .B(n42070), .Z(n42057) );
  AND U41829 ( .A(n42071), .B(n42072), .Z(n42070) );
  XOR U41830 ( .A(n42069), .B(n41699), .Z(n42072) );
  XOR U41831 ( .A(n42073), .B(n42074), .Z(n41699) );
  AND U41832 ( .A(n603), .B(n42075), .Z(n42074) );
  XOR U41833 ( .A(n42076), .B(n42073), .Z(n42075) );
  XNOR U41834 ( .A(n41696), .B(n42069), .Z(n42071) );
  XOR U41835 ( .A(n42077), .B(n42078), .Z(n41696) );
  AND U41836 ( .A(n601), .B(n42079), .Z(n42078) );
  XOR U41837 ( .A(n42080), .B(n42077), .Z(n42079) );
  XOR U41838 ( .A(n42081), .B(n42082), .Z(n42069) );
  AND U41839 ( .A(n42083), .B(n42084), .Z(n42082) );
  XOR U41840 ( .A(n42081), .B(n41711), .Z(n42084) );
  XOR U41841 ( .A(n42085), .B(n42086), .Z(n41711) );
  AND U41842 ( .A(n603), .B(n42087), .Z(n42086) );
  XOR U41843 ( .A(n42088), .B(n42085), .Z(n42087) );
  XNOR U41844 ( .A(n41708), .B(n42081), .Z(n42083) );
  XOR U41845 ( .A(n42089), .B(n42090), .Z(n41708) );
  AND U41846 ( .A(n601), .B(n42091), .Z(n42090) );
  XOR U41847 ( .A(n42092), .B(n42089), .Z(n42091) );
  XOR U41848 ( .A(n42093), .B(n42094), .Z(n42081) );
  AND U41849 ( .A(n42095), .B(n42096), .Z(n42094) );
  XOR U41850 ( .A(n42093), .B(n41723), .Z(n42096) );
  XOR U41851 ( .A(n42097), .B(n42098), .Z(n41723) );
  AND U41852 ( .A(n603), .B(n42099), .Z(n42098) );
  XOR U41853 ( .A(n42100), .B(n42097), .Z(n42099) );
  XNOR U41854 ( .A(n41720), .B(n42093), .Z(n42095) );
  XOR U41855 ( .A(n42101), .B(n42102), .Z(n41720) );
  AND U41856 ( .A(n601), .B(n42103), .Z(n42102) );
  XOR U41857 ( .A(n42104), .B(n42101), .Z(n42103) );
  XOR U41858 ( .A(n42105), .B(n42106), .Z(n42093) );
  AND U41859 ( .A(n42107), .B(n42108), .Z(n42106) );
  XOR U41860 ( .A(n42105), .B(n41735), .Z(n42108) );
  XOR U41861 ( .A(n42109), .B(n42110), .Z(n41735) );
  AND U41862 ( .A(n603), .B(n42111), .Z(n42110) );
  XOR U41863 ( .A(n42112), .B(n42109), .Z(n42111) );
  XNOR U41864 ( .A(n41732), .B(n42105), .Z(n42107) );
  XOR U41865 ( .A(n42113), .B(n42114), .Z(n41732) );
  AND U41866 ( .A(n601), .B(n42115), .Z(n42114) );
  XOR U41867 ( .A(n42116), .B(n42113), .Z(n42115) );
  XOR U41868 ( .A(n42117), .B(n42118), .Z(n42105) );
  AND U41869 ( .A(n42119), .B(n42120), .Z(n42118) );
  XOR U41870 ( .A(n42117), .B(n41747), .Z(n42120) );
  XOR U41871 ( .A(n42121), .B(n42122), .Z(n41747) );
  AND U41872 ( .A(n603), .B(n42123), .Z(n42122) );
  XOR U41873 ( .A(n42124), .B(n42121), .Z(n42123) );
  XNOR U41874 ( .A(n41744), .B(n42117), .Z(n42119) );
  XOR U41875 ( .A(n42125), .B(n42126), .Z(n41744) );
  AND U41876 ( .A(n601), .B(n42127), .Z(n42126) );
  XOR U41877 ( .A(n42128), .B(n42125), .Z(n42127) );
  XOR U41878 ( .A(n42129), .B(n42130), .Z(n42117) );
  AND U41879 ( .A(n42131), .B(n42132), .Z(n42130) );
  XOR U41880 ( .A(n42129), .B(n41759), .Z(n42132) );
  XOR U41881 ( .A(n42133), .B(n42134), .Z(n41759) );
  AND U41882 ( .A(n603), .B(n42135), .Z(n42134) );
  XOR U41883 ( .A(n42136), .B(n42133), .Z(n42135) );
  XNOR U41884 ( .A(n41756), .B(n42129), .Z(n42131) );
  XOR U41885 ( .A(n42137), .B(n42138), .Z(n41756) );
  AND U41886 ( .A(n601), .B(n42139), .Z(n42138) );
  XOR U41887 ( .A(n42140), .B(n42137), .Z(n42139) );
  XOR U41888 ( .A(n42141), .B(n42142), .Z(n42129) );
  AND U41889 ( .A(n42143), .B(n42144), .Z(n42142) );
  XOR U41890 ( .A(n42141), .B(n41771), .Z(n42144) );
  XOR U41891 ( .A(n42145), .B(n42146), .Z(n41771) );
  AND U41892 ( .A(n603), .B(n42147), .Z(n42146) );
  XOR U41893 ( .A(n42148), .B(n42145), .Z(n42147) );
  XNOR U41894 ( .A(n41768), .B(n42141), .Z(n42143) );
  XOR U41895 ( .A(n42149), .B(n42150), .Z(n41768) );
  AND U41896 ( .A(n601), .B(n42151), .Z(n42150) );
  XOR U41897 ( .A(n42152), .B(n42149), .Z(n42151) );
  XOR U41898 ( .A(n42153), .B(n42154), .Z(n42141) );
  AND U41899 ( .A(n42155), .B(n42156), .Z(n42154) );
  XOR U41900 ( .A(n42153), .B(n41783), .Z(n42156) );
  XOR U41901 ( .A(n42157), .B(n42158), .Z(n41783) );
  AND U41902 ( .A(n603), .B(n42159), .Z(n42158) );
  XOR U41903 ( .A(n42160), .B(n42157), .Z(n42159) );
  XNOR U41904 ( .A(n41780), .B(n42153), .Z(n42155) );
  XOR U41905 ( .A(n42161), .B(n42162), .Z(n41780) );
  AND U41906 ( .A(n601), .B(n42163), .Z(n42162) );
  XOR U41907 ( .A(n42164), .B(n42161), .Z(n42163) );
  XOR U41908 ( .A(n42165), .B(n42166), .Z(n42153) );
  AND U41909 ( .A(n42167), .B(n42168), .Z(n42166) );
  XOR U41910 ( .A(n42165), .B(n41795), .Z(n42168) );
  XOR U41911 ( .A(n42169), .B(n42170), .Z(n41795) );
  AND U41912 ( .A(n603), .B(n42171), .Z(n42170) );
  XOR U41913 ( .A(n42172), .B(n42169), .Z(n42171) );
  XNOR U41914 ( .A(n41792), .B(n42165), .Z(n42167) );
  XOR U41915 ( .A(n42173), .B(n42174), .Z(n41792) );
  AND U41916 ( .A(n601), .B(n42175), .Z(n42174) );
  XOR U41917 ( .A(n42176), .B(n42173), .Z(n42175) );
  XOR U41918 ( .A(n42177), .B(n42178), .Z(n42165) );
  AND U41919 ( .A(n42179), .B(n42180), .Z(n42178) );
  XOR U41920 ( .A(n42177), .B(n41807), .Z(n42180) );
  XOR U41921 ( .A(n42181), .B(n42182), .Z(n41807) );
  AND U41922 ( .A(n603), .B(n42183), .Z(n42182) );
  XOR U41923 ( .A(n42184), .B(n42181), .Z(n42183) );
  XNOR U41924 ( .A(n41804), .B(n42177), .Z(n42179) );
  XOR U41925 ( .A(n42185), .B(n42186), .Z(n41804) );
  AND U41926 ( .A(n601), .B(n42187), .Z(n42186) );
  XOR U41927 ( .A(n42188), .B(n42185), .Z(n42187) );
  XOR U41928 ( .A(n42189), .B(n42190), .Z(n42177) );
  AND U41929 ( .A(n42191), .B(n42192), .Z(n42190) );
  XOR U41930 ( .A(n42189), .B(n41819), .Z(n42192) );
  XOR U41931 ( .A(n42193), .B(n42194), .Z(n41819) );
  AND U41932 ( .A(n603), .B(n42195), .Z(n42194) );
  XOR U41933 ( .A(n42196), .B(n42193), .Z(n42195) );
  XNOR U41934 ( .A(n41816), .B(n42189), .Z(n42191) );
  XOR U41935 ( .A(n42197), .B(n42198), .Z(n41816) );
  AND U41936 ( .A(n601), .B(n42199), .Z(n42198) );
  XOR U41937 ( .A(n42200), .B(n42197), .Z(n42199) );
  XOR U41938 ( .A(n42201), .B(n42202), .Z(n42189) );
  AND U41939 ( .A(n42203), .B(n42204), .Z(n42202) );
  XOR U41940 ( .A(n42201), .B(n41831), .Z(n42204) );
  XOR U41941 ( .A(n42205), .B(n42206), .Z(n41831) );
  AND U41942 ( .A(n603), .B(n42207), .Z(n42206) );
  XOR U41943 ( .A(n42208), .B(n42205), .Z(n42207) );
  XNOR U41944 ( .A(n41828), .B(n42201), .Z(n42203) );
  XOR U41945 ( .A(n42209), .B(n42210), .Z(n41828) );
  AND U41946 ( .A(n601), .B(n42211), .Z(n42210) );
  XOR U41947 ( .A(n42212), .B(n42209), .Z(n42211) );
  XOR U41948 ( .A(n42213), .B(n42214), .Z(n42201) );
  AND U41949 ( .A(n42215), .B(n42216), .Z(n42214) );
  XOR U41950 ( .A(n42213), .B(n41843), .Z(n42216) );
  XOR U41951 ( .A(n42217), .B(n42218), .Z(n41843) );
  AND U41952 ( .A(n603), .B(n42219), .Z(n42218) );
  XOR U41953 ( .A(n42220), .B(n42217), .Z(n42219) );
  XNOR U41954 ( .A(n41840), .B(n42213), .Z(n42215) );
  XOR U41955 ( .A(n42221), .B(n42222), .Z(n41840) );
  AND U41956 ( .A(n601), .B(n42223), .Z(n42222) );
  XOR U41957 ( .A(n42224), .B(n42221), .Z(n42223) );
  XOR U41958 ( .A(n42225), .B(n42226), .Z(n42213) );
  AND U41959 ( .A(n42227), .B(n42228), .Z(n42226) );
  XOR U41960 ( .A(n42225), .B(n41855), .Z(n42228) );
  XOR U41961 ( .A(n42229), .B(n42230), .Z(n41855) );
  AND U41962 ( .A(n603), .B(n42231), .Z(n42230) );
  XOR U41963 ( .A(n42232), .B(n42229), .Z(n42231) );
  XNOR U41964 ( .A(n41852), .B(n42225), .Z(n42227) );
  XOR U41965 ( .A(n42233), .B(n42234), .Z(n41852) );
  AND U41966 ( .A(n601), .B(n42235), .Z(n42234) );
  XOR U41967 ( .A(n42236), .B(n42233), .Z(n42235) );
  XOR U41968 ( .A(n42237), .B(n42238), .Z(n42225) );
  AND U41969 ( .A(n42239), .B(n42240), .Z(n42238) );
  XOR U41970 ( .A(n42237), .B(n41867), .Z(n42240) );
  XOR U41971 ( .A(n42241), .B(n42242), .Z(n41867) );
  AND U41972 ( .A(n603), .B(n42243), .Z(n42242) );
  XOR U41973 ( .A(n42244), .B(n42241), .Z(n42243) );
  XNOR U41974 ( .A(n41864), .B(n42237), .Z(n42239) );
  XOR U41975 ( .A(n42245), .B(n42246), .Z(n41864) );
  AND U41976 ( .A(n601), .B(n42247), .Z(n42246) );
  XOR U41977 ( .A(n42248), .B(n42245), .Z(n42247) );
  XOR U41978 ( .A(n42249), .B(n42250), .Z(n42237) );
  AND U41979 ( .A(n42251), .B(n42252), .Z(n42250) );
  XOR U41980 ( .A(n42249), .B(n41879), .Z(n42252) );
  XOR U41981 ( .A(n42253), .B(n42254), .Z(n41879) );
  AND U41982 ( .A(n603), .B(n42255), .Z(n42254) );
  XOR U41983 ( .A(n42256), .B(n42253), .Z(n42255) );
  XNOR U41984 ( .A(n41876), .B(n42249), .Z(n42251) );
  XOR U41985 ( .A(n42257), .B(n42258), .Z(n41876) );
  AND U41986 ( .A(n601), .B(n42259), .Z(n42258) );
  XOR U41987 ( .A(n42260), .B(n42257), .Z(n42259) );
  XOR U41988 ( .A(n42261), .B(n42262), .Z(n42249) );
  AND U41989 ( .A(n42263), .B(n42264), .Z(n42262) );
  XOR U41990 ( .A(n42261), .B(n41891), .Z(n42264) );
  XOR U41991 ( .A(n42265), .B(n42266), .Z(n41891) );
  AND U41992 ( .A(n603), .B(n42267), .Z(n42266) );
  XOR U41993 ( .A(n42268), .B(n42265), .Z(n42267) );
  XNOR U41994 ( .A(n41888), .B(n42261), .Z(n42263) );
  XOR U41995 ( .A(n42269), .B(n42270), .Z(n41888) );
  AND U41996 ( .A(n601), .B(n42271), .Z(n42270) );
  XOR U41997 ( .A(n42272), .B(n42269), .Z(n42271) );
  XOR U41998 ( .A(n42273), .B(n42274), .Z(n42261) );
  AND U41999 ( .A(n42275), .B(n42276), .Z(n42274) );
  XOR U42000 ( .A(n42273), .B(n41903), .Z(n42276) );
  XOR U42001 ( .A(n42277), .B(n42278), .Z(n41903) );
  AND U42002 ( .A(n603), .B(n42279), .Z(n42278) );
  XOR U42003 ( .A(n42280), .B(n42277), .Z(n42279) );
  XNOR U42004 ( .A(n41900), .B(n42273), .Z(n42275) );
  XOR U42005 ( .A(n42281), .B(n42282), .Z(n41900) );
  AND U42006 ( .A(n601), .B(n42283), .Z(n42282) );
  XOR U42007 ( .A(n42284), .B(n42281), .Z(n42283) );
  XOR U42008 ( .A(n42285), .B(n42286), .Z(n42273) );
  AND U42009 ( .A(n42287), .B(n42288), .Z(n42286) );
  XOR U42010 ( .A(n42285), .B(n41915), .Z(n42288) );
  XOR U42011 ( .A(n42289), .B(n42290), .Z(n41915) );
  AND U42012 ( .A(n603), .B(n42291), .Z(n42290) );
  XOR U42013 ( .A(n42292), .B(n42289), .Z(n42291) );
  XNOR U42014 ( .A(n41912), .B(n42285), .Z(n42287) );
  XOR U42015 ( .A(n42293), .B(n42294), .Z(n41912) );
  AND U42016 ( .A(n601), .B(n42295), .Z(n42294) );
  XOR U42017 ( .A(n42296), .B(n42293), .Z(n42295) );
  XOR U42018 ( .A(n42297), .B(n42298), .Z(n42285) );
  AND U42019 ( .A(n42299), .B(n42300), .Z(n42298) );
  XOR U42020 ( .A(n42297), .B(n41927), .Z(n42300) );
  XOR U42021 ( .A(n42301), .B(n42302), .Z(n41927) );
  AND U42022 ( .A(n603), .B(n42303), .Z(n42302) );
  XOR U42023 ( .A(n42304), .B(n42301), .Z(n42303) );
  XNOR U42024 ( .A(n41924), .B(n42297), .Z(n42299) );
  XOR U42025 ( .A(n42305), .B(n42306), .Z(n41924) );
  AND U42026 ( .A(n601), .B(n42307), .Z(n42306) );
  XOR U42027 ( .A(n42308), .B(n42305), .Z(n42307) );
  XOR U42028 ( .A(n42309), .B(n42310), .Z(n42297) );
  AND U42029 ( .A(n42311), .B(n42312), .Z(n42310) );
  XOR U42030 ( .A(n42309), .B(n41939), .Z(n42312) );
  XOR U42031 ( .A(n42313), .B(n42314), .Z(n41939) );
  AND U42032 ( .A(n603), .B(n42315), .Z(n42314) );
  XOR U42033 ( .A(n42316), .B(n42313), .Z(n42315) );
  XNOR U42034 ( .A(n41936), .B(n42309), .Z(n42311) );
  XOR U42035 ( .A(n42317), .B(n42318), .Z(n41936) );
  AND U42036 ( .A(n601), .B(n42319), .Z(n42318) );
  XOR U42037 ( .A(n42320), .B(n42317), .Z(n42319) );
  XOR U42038 ( .A(n42321), .B(n42322), .Z(n42309) );
  AND U42039 ( .A(n42323), .B(n42324), .Z(n42322) );
  XOR U42040 ( .A(n42321), .B(n41951), .Z(n42324) );
  XOR U42041 ( .A(n42325), .B(n42326), .Z(n41951) );
  AND U42042 ( .A(n603), .B(n42327), .Z(n42326) );
  XOR U42043 ( .A(n42328), .B(n42325), .Z(n42327) );
  XNOR U42044 ( .A(n41948), .B(n42321), .Z(n42323) );
  XOR U42045 ( .A(n42329), .B(n42330), .Z(n41948) );
  AND U42046 ( .A(n601), .B(n42331), .Z(n42330) );
  XOR U42047 ( .A(n42332), .B(n42329), .Z(n42331) );
  XOR U42048 ( .A(n42333), .B(n42334), .Z(n42321) );
  AND U42049 ( .A(n42335), .B(n42336), .Z(n42334) );
  XOR U42050 ( .A(n42333), .B(n41963), .Z(n42336) );
  XOR U42051 ( .A(n42337), .B(n42338), .Z(n41963) );
  AND U42052 ( .A(n603), .B(n42339), .Z(n42338) );
  XOR U42053 ( .A(n42340), .B(n42337), .Z(n42339) );
  XNOR U42054 ( .A(n41960), .B(n42333), .Z(n42335) );
  XOR U42055 ( .A(n42341), .B(n42342), .Z(n41960) );
  AND U42056 ( .A(n601), .B(n42343), .Z(n42342) );
  XOR U42057 ( .A(n42344), .B(n42341), .Z(n42343) );
  XOR U42058 ( .A(n42345), .B(n42346), .Z(n42333) );
  AND U42059 ( .A(n42347), .B(n42348), .Z(n42346) );
  XNOR U42060 ( .A(n42349), .B(n41976), .Z(n42348) );
  XOR U42061 ( .A(n42350), .B(n42351), .Z(n41976) );
  AND U42062 ( .A(n603), .B(n42352), .Z(n42351) );
  XOR U42063 ( .A(n42350), .B(n42353), .Z(n42352) );
  XNOR U42064 ( .A(n41973), .B(n42345), .Z(n42347) );
  XOR U42065 ( .A(n42354), .B(n42355), .Z(n41973) );
  AND U42066 ( .A(n601), .B(n42356), .Z(n42355) );
  XOR U42067 ( .A(n42354), .B(n42357), .Z(n42356) );
  IV U42068 ( .A(n42349), .Z(n42345) );
  AND U42069 ( .A(n41981), .B(n41984), .Z(n42349) );
  XNOR U42070 ( .A(n42358), .B(n42359), .Z(n41984) );
  AND U42071 ( .A(n603), .B(n42360), .Z(n42359) );
  XNOR U42072 ( .A(n42361), .B(n42358), .Z(n42360) );
  XOR U42073 ( .A(n42362), .B(n42363), .Z(n603) );
  AND U42074 ( .A(n42364), .B(n42365), .Z(n42363) );
  XOR U42075 ( .A(n41992), .B(n42362), .Z(n42365) );
  IV U42076 ( .A(n42366), .Z(n41992) );
  AND U42077 ( .A(p_input[2559]), .B(p_input[2527]), .Z(n42366) );
  XOR U42078 ( .A(n42362), .B(n41989), .Z(n42364) );
  AND U42079 ( .A(p_input[2463]), .B(p_input[2495]), .Z(n41989) );
  XOR U42080 ( .A(n42367), .B(n42368), .Z(n42362) );
  AND U42081 ( .A(n42369), .B(n42370), .Z(n42368) );
  XOR U42082 ( .A(n42367), .B(n42004), .Z(n42370) );
  XNOR U42083 ( .A(p_input[2526]), .B(n42371), .Z(n42004) );
  AND U42084 ( .A(n779), .B(n42372), .Z(n42371) );
  XOR U42085 ( .A(p_input[2558]), .B(p_input[2526]), .Z(n42372) );
  XNOR U42086 ( .A(n42001), .B(n42367), .Z(n42369) );
  XOR U42087 ( .A(n42373), .B(n42374), .Z(n42001) );
  AND U42088 ( .A(n777), .B(n42375), .Z(n42374) );
  XOR U42089 ( .A(p_input[2494]), .B(p_input[2462]), .Z(n42375) );
  XOR U42090 ( .A(n42376), .B(n42377), .Z(n42367) );
  AND U42091 ( .A(n42378), .B(n42379), .Z(n42377) );
  XOR U42092 ( .A(n42376), .B(n42016), .Z(n42379) );
  XNOR U42093 ( .A(p_input[2525]), .B(n42380), .Z(n42016) );
  AND U42094 ( .A(n779), .B(n42381), .Z(n42380) );
  XOR U42095 ( .A(p_input[2557]), .B(p_input[2525]), .Z(n42381) );
  XNOR U42096 ( .A(n42013), .B(n42376), .Z(n42378) );
  XOR U42097 ( .A(n42382), .B(n42383), .Z(n42013) );
  AND U42098 ( .A(n777), .B(n42384), .Z(n42383) );
  XOR U42099 ( .A(p_input[2493]), .B(p_input[2461]), .Z(n42384) );
  XOR U42100 ( .A(n42385), .B(n42386), .Z(n42376) );
  AND U42101 ( .A(n42387), .B(n42388), .Z(n42386) );
  XOR U42102 ( .A(n42385), .B(n42028), .Z(n42388) );
  XNOR U42103 ( .A(p_input[2524]), .B(n42389), .Z(n42028) );
  AND U42104 ( .A(n779), .B(n42390), .Z(n42389) );
  XOR U42105 ( .A(p_input[2556]), .B(p_input[2524]), .Z(n42390) );
  XNOR U42106 ( .A(n42025), .B(n42385), .Z(n42387) );
  XOR U42107 ( .A(n42391), .B(n42392), .Z(n42025) );
  AND U42108 ( .A(n777), .B(n42393), .Z(n42392) );
  XOR U42109 ( .A(p_input[2492]), .B(p_input[2460]), .Z(n42393) );
  XOR U42110 ( .A(n42394), .B(n42395), .Z(n42385) );
  AND U42111 ( .A(n42396), .B(n42397), .Z(n42395) );
  XOR U42112 ( .A(n42394), .B(n42040), .Z(n42397) );
  XNOR U42113 ( .A(p_input[2523]), .B(n42398), .Z(n42040) );
  AND U42114 ( .A(n779), .B(n42399), .Z(n42398) );
  XOR U42115 ( .A(p_input[2555]), .B(p_input[2523]), .Z(n42399) );
  XNOR U42116 ( .A(n42037), .B(n42394), .Z(n42396) );
  XOR U42117 ( .A(n42400), .B(n42401), .Z(n42037) );
  AND U42118 ( .A(n777), .B(n42402), .Z(n42401) );
  XOR U42119 ( .A(p_input[2491]), .B(p_input[2459]), .Z(n42402) );
  XOR U42120 ( .A(n42403), .B(n42404), .Z(n42394) );
  AND U42121 ( .A(n42405), .B(n42406), .Z(n42404) );
  XOR U42122 ( .A(n42403), .B(n42052), .Z(n42406) );
  XNOR U42123 ( .A(p_input[2522]), .B(n42407), .Z(n42052) );
  AND U42124 ( .A(n779), .B(n42408), .Z(n42407) );
  XOR U42125 ( .A(p_input[2554]), .B(p_input[2522]), .Z(n42408) );
  XNOR U42126 ( .A(n42049), .B(n42403), .Z(n42405) );
  XOR U42127 ( .A(n42409), .B(n42410), .Z(n42049) );
  AND U42128 ( .A(n777), .B(n42411), .Z(n42410) );
  XOR U42129 ( .A(p_input[2490]), .B(p_input[2458]), .Z(n42411) );
  XOR U42130 ( .A(n42412), .B(n42413), .Z(n42403) );
  AND U42131 ( .A(n42414), .B(n42415), .Z(n42413) );
  XOR U42132 ( .A(n42412), .B(n42064), .Z(n42415) );
  XNOR U42133 ( .A(p_input[2521]), .B(n42416), .Z(n42064) );
  AND U42134 ( .A(n779), .B(n42417), .Z(n42416) );
  XOR U42135 ( .A(p_input[2553]), .B(p_input[2521]), .Z(n42417) );
  XNOR U42136 ( .A(n42061), .B(n42412), .Z(n42414) );
  XOR U42137 ( .A(n42418), .B(n42419), .Z(n42061) );
  AND U42138 ( .A(n777), .B(n42420), .Z(n42419) );
  XOR U42139 ( .A(p_input[2489]), .B(p_input[2457]), .Z(n42420) );
  XOR U42140 ( .A(n42421), .B(n42422), .Z(n42412) );
  AND U42141 ( .A(n42423), .B(n42424), .Z(n42422) );
  XOR U42142 ( .A(n42421), .B(n42076), .Z(n42424) );
  XNOR U42143 ( .A(p_input[2520]), .B(n42425), .Z(n42076) );
  AND U42144 ( .A(n779), .B(n42426), .Z(n42425) );
  XOR U42145 ( .A(p_input[2552]), .B(p_input[2520]), .Z(n42426) );
  XNOR U42146 ( .A(n42073), .B(n42421), .Z(n42423) );
  XOR U42147 ( .A(n42427), .B(n42428), .Z(n42073) );
  AND U42148 ( .A(n777), .B(n42429), .Z(n42428) );
  XOR U42149 ( .A(p_input[2488]), .B(p_input[2456]), .Z(n42429) );
  XOR U42150 ( .A(n42430), .B(n42431), .Z(n42421) );
  AND U42151 ( .A(n42432), .B(n42433), .Z(n42431) );
  XOR U42152 ( .A(n42430), .B(n42088), .Z(n42433) );
  XNOR U42153 ( .A(p_input[2519]), .B(n42434), .Z(n42088) );
  AND U42154 ( .A(n779), .B(n42435), .Z(n42434) );
  XOR U42155 ( .A(p_input[2551]), .B(p_input[2519]), .Z(n42435) );
  XNOR U42156 ( .A(n42085), .B(n42430), .Z(n42432) );
  XOR U42157 ( .A(n42436), .B(n42437), .Z(n42085) );
  AND U42158 ( .A(n777), .B(n42438), .Z(n42437) );
  XOR U42159 ( .A(p_input[2487]), .B(p_input[2455]), .Z(n42438) );
  XOR U42160 ( .A(n42439), .B(n42440), .Z(n42430) );
  AND U42161 ( .A(n42441), .B(n42442), .Z(n42440) );
  XOR U42162 ( .A(n42439), .B(n42100), .Z(n42442) );
  XNOR U42163 ( .A(p_input[2518]), .B(n42443), .Z(n42100) );
  AND U42164 ( .A(n779), .B(n42444), .Z(n42443) );
  XOR U42165 ( .A(p_input[2550]), .B(p_input[2518]), .Z(n42444) );
  XNOR U42166 ( .A(n42097), .B(n42439), .Z(n42441) );
  XOR U42167 ( .A(n42445), .B(n42446), .Z(n42097) );
  AND U42168 ( .A(n777), .B(n42447), .Z(n42446) );
  XOR U42169 ( .A(p_input[2486]), .B(p_input[2454]), .Z(n42447) );
  XOR U42170 ( .A(n42448), .B(n42449), .Z(n42439) );
  AND U42171 ( .A(n42450), .B(n42451), .Z(n42449) );
  XOR U42172 ( .A(n42448), .B(n42112), .Z(n42451) );
  XNOR U42173 ( .A(p_input[2517]), .B(n42452), .Z(n42112) );
  AND U42174 ( .A(n779), .B(n42453), .Z(n42452) );
  XOR U42175 ( .A(p_input[2549]), .B(p_input[2517]), .Z(n42453) );
  XNOR U42176 ( .A(n42109), .B(n42448), .Z(n42450) );
  XOR U42177 ( .A(n42454), .B(n42455), .Z(n42109) );
  AND U42178 ( .A(n777), .B(n42456), .Z(n42455) );
  XOR U42179 ( .A(p_input[2485]), .B(p_input[2453]), .Z(n42456) );
  XOR U42180 ( .A(n42457), .B(n42458), .Z(n42448) );
  AND U42181 ( .A(n42459), .B(n42460), .Z(n42458) );
  XOR U42182 ( .A(n42457), .B(n42124), .Z(n42460) );
  XNOR U42183 ( .A(p_input[2516]), .B(n42461), .Z(n42124) );
  AND U42184 ( .A(n779), .B(n42462), .Z(n42461) );
  XOR U42185 ( .A(p_input[2548]), .B(p_input[2516]), .Z(n42462) );
  XNOR U42186 ( .A(n42121), .B(n42457), .Z(n42459) );
  XOR U42187 ( .A(n42463), .B(n42464), .Z(n42121) );
  AND U42188 ( .A(n777), .B(n42465), .Z(n42464) );
  XOR U42189 ( .A(p_input[2484]), .B(p_input[2452]), .Z(n42465) );
  XOR U42190 ( .A(n42466), .B(n42467), .Z(n42457) );
  AND U42191 ( .A(n42468), .B(n42469), .Z(n42467) );
  XOR U42192 ( .A(n42466), .B(n42136), .Z(n42469) );
  XNOR U42193 ( .A(p_input[2515]), .B(n42470), .Z(n42136) );
  AND U42194 ( .A(n779), .B(n42471), .Z(n42470) );
  XOR U42195 ( .A(p_input[2547]), .B(p_input[2515]), .Z(n42471) );
  XNOR U42196 ( .A(n42133), .B(n42466), .Z(n42468) );
  XOR U42197 ( .A(n42472), .B(n42473), .Z(n42133) );
  AND U42198 ( .A(n777), .B(n42474), .Z(n42473) );
  XOR U42199 ( .A(p_input[2483]), .B(p_input[2451]), .Z(n42474) );
  XOR U42200 ( .A(n42475), .B(n42476), .Z(n42466) );
  AND U42201 ( .A(n42477), .B(n42478), .Z(n42476) );
  XOR U42202 ( .A(n42475), .B(n42148), .Z(n42478) );
  XNOR U42203 ( .A(p_input[2514]), .B(n42479), .Z(n42148) );
  AND U42204 ( .A(n779), .B(n42480), .Z(n42479) );
  XOR U42205 ( .A(p_input[2546]), .B(p_input[2514]), .Z(n42480) );
  XNOR U42206 ( .A(n42145), .B(n42475), .Z(n42477) );
  XOR U42207 ( .A(n42481), .B(n42482), .Z(n42145) );
  AND U42208 ( .A(n777), .B(n42483), .Z(n42482) );
  XOR U42209 ( .A(p_input[2482]), .B(p_input[2450]), .Z(n42483) );
  XOR U42210 ( .A(n42484), .B(n42485), .Z(n42475) );
  AND U42211 ( .A(n42486), .B(n42487), .Z(n42485) );
  XOR U42212 ( .A(n42484), .B(n42160), .Z(n42487) );
  XNOR U42213 ( .A(p_input[2513]), .B(n42488), .Z(n42160) );
  AND U42214 ( .A(n779), .B(n42489), .Z(n42488) );
  XOR U42215 ( .A(p_input[2545]), .B(p_input[2513]), .Z(n42489) );
  XNOR U42216 ( .A(n42157), .B(n42484), .Z(n42486) );
  XOR U42217 ( .A(n42490), .B(n42491), .Z(n42157) );
  AND U42218 ( .A(n777), .B(n42492), .Z(n42491) );
  XOR U42219 ( .A(p_input[2481]), .B(p_input[2449]), .Z(n42492) );
  XOR U42220 ( .A(n42493), .B(n42494), .Z(n42484) );
  AND U42221 ( .A(n42495), .B(n42496), .Z(n42494) );
  XOR U42222 ( .A(n42493), .B(n42172), .Z(n42496) );
  XNOR U42223 ( .A(p_input[2512]), .B(n42497), .Z(n42172) );
  AND U42224 ( .A(n779), .B(n42498), .Z(n42497) );
  XOR U42225 ( .A(p_input[2544]), .B(p_input[2512]), .Z(n42498) );
  XNOR U42226 ( .A(n42169), .B(n42493), .Z(n42495) );
  XOR U42227 ( .A(n42499), .B(n42500), .Z(n42169) );
  AND U42228 ( .A(n777), .B(n42501), .Z(n42500) );
  XOR U42229 ( .A(p_input[2480]), .B(p_input[2448]), .Z(n42501) );
  XOR U42230 ( .A(n42502), .B(n42503), .Z(n42493) );
  AND U42231 ( .A(n42504), .B(n42505), .Z(n42503) );
  XOR U42232 ( .A(n42502), .B(n42184), .Z(n42505) );
  XNOR U42233 ( .A(p_input[2511]), .B(n42506), .Z(n42184) );
  AND U42234 ( .A(n779), .B(n42507), .Z(n42506) );
  XOR U42235 ( .A(p_input[2543]), .B(p_input[2511]), .Z(n42507) );
  XNOR U42236 ( .A(n42181), .B(n42502), .Z(n42504) );
  XOR U42237 ( .A(n42508), .B(n42509), .Z(n42181) );
  AND U42238 ( .A(n777), .B(n42510), .Z(n42509) );
  XOR U42239 ( .A(p_input[2479]), .B(p_input[2447]), .Z(n42510) );
  XOR U42240 ( .A(n42511), .B(n42512), .Z(n42502) );
  AND U42241 ( .A(n42513), .B(n42514), .Z(n42512) );
  XOR U42242 ( .A(n42511), .B(n42196), .Z(n42514) );
  XNOR U42243 ( .A(p_input[2510]), .B(n42515), .Z(n42196) );
  AND U42244 ( .A(n779), .B(n42516), .Z(n42515) );
  XOR U42245 ( .A(p_input[2542]), .B(p_input[2510]), .Z(n42516) );
  XNOR U42246 ( .A(n42193), .B(n42511), .Z(n42513) );
  XOR U42247 ( .A(n42517), .B(n42518), .Z(n42193) );
  AND U42248 ( .A(n777), .B(n42519), .Z(n42518) );
  XOR U42249 ( .A(p_input[2478]), .B(p_input[2446]), .Z(n42519) );
  XOR U42250 ( .A(n42520), .B(n42521), .Z(n42511) );
  AND U42251 ( .A(n42522), .B(n42523), .Z(n42521) );
  XOR U42252 ( .A(n42520), .B(n42208), .Z(n42523) );
  XNOR U42253 ( .A(p_input[2509]), .B(n42524), .Z(n42208) );
  AND U42254 ( .A(n779), .B(n42525), .Z(n42524) );
  XOR U42255 ( .A(p_input[2541]), .B(p_input[2509]), .Z(n42525) );
  XNOR U42256 ( .A(n42205), .B(n42520), .Z(n42522) );
  XOR U42257 ( .A(n42526), .B(n42527), .Z(n42205) );
  AND U42258 ( .A(n777), .B(n42528), .Z(n42527) );
  XOR U42259 ( .A(p_input[2477]), .B(p_input[2445]), .Z(n42528) );
  XOR U42260 ( .A(n42529), .B(n42530), .Z(n42520) );
  AND U42261 ( .A(n42531), .B(n42532), .Z(n42530) );
  XOR U42262 ( .A(n42529), .B(n42220), .Z(n42532) );
  XNOR U42263 ( .A(p_input[2508]), .B(n42533), .Z(n42220) );
  AND U42264 ( .A(n779), .B(n42534), .Z(n42533) );
  XOR U42265 ( .A(p_input[2540]), .B(p_input[2508]), .Z(n42534) );
  XNOR U42266 ( .A(n42217), .B(n42529), .Z(n42531) );
  XOR U42267 ( .A(n42535), .B(n42536), .Z(n42217) );
  AND U42268 ( .A(n777), .B(n42537), .Z(n42536) );
  XOR U42269 ( .A(p_input[2476]), .B(p_input[2444]), .Z(n42537) );
  XOR U42270 ( .A(n42538), .B(n42539), .Z(n42529) );
  AND U42271 ( .A(n42540), .B(n42541), .Z(n42539) );
  XOR U42272 ( .A(n42538), .B(n42232), .Z(n42541) );
  XNOR U42273 ( .A(p_input[2507]), .B(n42542), .Z(n42232) );
  AND U42274 ( .A(n779), .B(n42543), .Z(n42542) );
  XOR U42275 ( .A(p_input[2539]), .B(p_input[2507]), .Z(n42543) );
  XNOR U42276 ( .A(n42229), .B(n42538), .Z(n42540) );
  XOR U42277 ( .A(n42544), .B(n42545), .Z(n42229) );
  AND U42278 ( .A(n777), .B(n42546), .Z(n42545) );
  XOR U42279 ( .A(p_input[2475]), .B(p_input[2443]), .Z(n42546) );
  XOR U42280 ( .A(n42547), .B(n42548), .Z(n42538) );
  AND U42281 ( .A(n42549), .B(n42550), .Z(n42548) );
  XOR U42282 ( .A(n42547), .B(n42244), .Z(n42550) );
  XNOR U42283 ( .A(p_input[2506]), .B(n42551), .Z(n42244) );
  AND U42284 ( .A(n779), .B(n42552), .Z(n42551) );
  XOR U42285 ( .A(p_input[2538]), .B(p_input[2506]), .Z(n42552) );
  XNOR U42286 ( .A(n42241), .B(n42547), .Z(n42549) );
  XOR U42287 ( .A(n42553), .B(n42554), .Z(n42241) );
  AND U42288 ( .A(n777), .B(n42555), .Z(n42554) );
  XOR U42289 ( .A(p_input[2474]), .B(p_input[2442]), .Z(n42555) );
  XOR U42290 ( .A(n42556), .B(n42557), .Z(n42547) );
  AND U42291 ( .A(n42558), .B(n42559), .Z(n42557) );
  XOR U42292 ( .A(n42556), .B(n42256), .Z(n42559) );
  XNOR U42293 ( .A(p_input[2505]), .B(n42560), .Z(n42256) );
  AND U42294 ( .A(n779), .B(n42561), .Z(n42560) );
  XOR U42295 ( .A(p_input[2537]), .B(p_input[2505]), .Z(n42561) );
  XNOR U42296 ( .A(n42253), .B(n42556), .Z(n42558) );
  XOR U42297 ( .A(n42562), .B(n42563), .Z(n42253) );
  AND U42298 ( .A(n777), .B(n42564), .Z(n42563) );
  XOR U42299 ( .A(p_input[2473]), .B(p_input[2441]), .Z(n42564) );
  XOR U42300 ( .A(n42565), .B(n42566), .Z(n42556) );
  AND U42301 ( .A(n42567), .B(n42568), .Z(n42566) );
  XOR U42302 ( .A(n42565), .B(n42268), .Z(n42568) );
  XNOR U42303 ( .A(p_input[2504]), .B(n42569), .Z(n42268) );
  AND U42304 ( .A(n779), .B(n42570), .Z(n42569) );
  XOR U42305 ( .A(p_input[2536]), .B(p_input[2504]), .Z(n42570) );
  XNOR U42306 ( .A(n42265), .B(n42565), .Z(n42567) );
  XOR U42307 ( .A(n42571), .B(n42572), .Z(n42265) );
  AND U42308 ( .A(n777), .B(n42573), .Z(n42572) );
  XOR U42309 ( .A(p_input[2472]), .B(p_input[2440]), .Z(n42573) );
  XOR U42310 ( .A(n42574), .B(n42575), .Z(n42565) );
  AND U42311 ( .A(n42576), .B(n42577), .Z(n42575) );
  XOR U42312 ( .A(n42574), .B(n42280), .Z(n42577) );
  XNOR U42313 ( .A(p_input[2503]), .B(n42578), .Z(n42280) );
  AND U42314 ( .A(n779), .B(n42579), .Z(n42578) );
  XOR U42315 ( .A(p_input[2535]), .B(p_input[2503]), .Z(n42579) );
  XNOR U42316 ( .A(n42277), .B(n42574), .Z(n42576) );
  XOR U42317 ( .A(n42580), .B(n42581), .Z(n42277) );
  AND U42318 ( .A(n777), .B(n42582), .Z(n42581) );
  XOR U42319 ( .A(p_input[2471]), .B(p_input[2439]), .Z(n42582) );
  XOR U42320 ( .A(n42583), .B(n42584), .Z(n42574) );
  AND U42321 ( .A(n42585), .B(n42586), .Z(n42584) );
  XOR U42322 ( .A(n42583), .B(n42292), .Z(n42586) );
  XNOR U42323 ( .A(p_input[2502]), .B(n42587), .Z(n42292) );
  AND U42324 ( .A(n779), .B(n42588), .Z(n42587) );
  XOR U42325 ( .A(p_input[2534]), .B(p_input[2502]), .Z(n42588) );
  XNOR U42326 ( .A(n42289), .B(n42583), .Z(n42585) );
  XOR U42327 ( .A(n42589), .B(n42590), .Z(n42289) );
  AND U42328 ( .A(n777), .B(n42591), .Z(n42590) );
  XOR U42329 ( .A(p_input[2470]), .B(p_input[2438]), .Z(n42591) );
  XOR U42330 ( .A(n42592), .B(n42593), .Z(n42583) );
  AND U42331 ( .A(n42594), .B(n42595), .Z(n42593) );
  XOR U42332 ( .A(n42592), .B(n42304), .Z(n42595) );
  XNOR U42333 ( .A(p_input[2501]), .B(n42596), .Z(n42304) );
  AND U42334 ( .A(n779), .B(n42597), .Z(n42596) );
  XOR U42335 ( .A(p_input[2533]), .B(p_input[2501]), .Z(n42597) );
  XNOR U42336 ( .A(n42301), .B(n42592), .Z(n42594) );
  XOR U42337 ( .A(n42598), .B(n42599), .Z(n42301) );
  AND U42338 ( .A(n777), .B(n42600), .Z(n42599) );
  XOR U42339 ( .A(p_input[2469]), .B(p_input[2437]), .Z(n42600) );
  XOR U42340 ( .A(n42601), .B(n42602), .Z(n42592) );
  AND U42341 ( .A(n42603), .B(n42604), .Z(n42602) );
  XOR U42342 ( .A(n42601), .B(n42316), .Z(n42604) );
  XNOR U42343 ( .A(p_input[2500]), .B(n42605), .Z(n42316) );
  AND U42344 ( .A(n779), .B(n42606), .Z(n42605) );
  XOR U42345 ( .A(p_input[2532]), .B(p_input[2500]), .Z(n42606) );
  XNOR U42346 ( .A(n42313), .B(n42601), .Z(n42603) );
  XOR U42347 ( .A(n42607), .B(n42608), .Z(n42313) );
  AND U42348 ( .A(n777), .B(n42609), .Z(n42608) );
  XOR U42349 ( .A(p_input[2468]), .B(p_input[2436]), .Z(n42609) );
  XOR U42350 ( .A(n42610), .B(n42611), .Z(n42601) );
  AND U42351 ( .A(n42612), .B(n42613), .Z(n42611) );
  XOR U42352 ( .A(n42610), .B(n42328), .Z(n42613) );
  XNOR U42353 ( .A(p_input[2499]), .B(n42614), .Z(n42328) );
  AND U42354 ( .A(n779), .B(n42615), .Z(n42614) );
  XOR U42355 ( .A(p_input[2531]), .B(p_input[2499]), .Z(n42615) );
  XNOR U42356 ( .A(n42325), .B(n42610), .Z(n42612) );
  XOR U42357 ( .A(n42616), .B(n42617), .Z(n42325) );
  AND U42358 ( .A(n777), .B(n42618), .Z(n42617) );
  XOR U42359 ( .A(p_input[2467]), .B(p_input[2435]), .Z(n42618) );
  XOR U42360 ( .A(n42619), .B(n42620), .Z(n42610) );
  AND U42361 ( .A(n42621), .B(n42622), .Z(n42620) );
  XOR U42362 ( .A(n42619), .B(n42340), .Z(n42622) );
  XNOR U42363 ( .A(p_input[2498]), .B(n42623), .Z(n42340) );
  AND U42364 ( .A(n779), .B(n42624), .Z(n42623) );
  XOR U42365 ( .A(p_input[2530]), .B(p_input[2498]), .Z(n42624) );
  XNOR U42366 ( .A(n42337), .B(n42619), .Z(n42621) );
  XOR U42367 ( .A(n42625), .B(n42626), .Z(n42337) );
  AND U42368 ( .A(n777), .B(n42627), .Z(n42626) );
  XOR U42369 ( .A(p_input[2466]), .B(p_input[2434]), .Z(n42627) );
  XOR U42370 ( .A(n42628), .B(n42629), .Z(n42619) );
  AND U42371 ( .A(n42630), .B(n42631), .Z(n42629) );
  XNOR U42372 ( .A(n42632), .B(n42353), .Z(n42631) );
  XNOR U42373 ( .A(p_input[2497]), .B(n42633), .Z(n42353) );
  AND U42374 ( .A(n779), .B(n42634), .Z(n42633) );
  XNOR U42375 ( .A(p_input[2529]), .B(n42635), .Z(n42634) );
  IV U42376 ( .A(p_input[2497]), .Z(n42635) );
  XNOR U42377 ( .A(n42350), .B(n42628), .Z(n42630) );
  XNOR U42378 ( .A(p_input[2433]), .B(n42636), .Z(n42350) );
  AND U42379 ( .A(n777), .B(n42637), .Z(n42636) );
  XOR U42380 ( .A(p_input[2465]), .B(p_input[2433]), .Z(n42637) );
  IV U42381 ( .A(n42632), .Z(n42628) );
  AND U42382 ( .A(n42358), .B(n42361), .Z(n42632) );
  XOR U42383 ( .A(p_input[2496]), .B(n42638), .Z(n42361) );
  AND U42384 ( .A(n779), .B(n42639), .Z(n42638) );
  XOR U42385 ( .A(p_input[2528]), .B(p_input[2496]), .Z(n42639) );
  XOR U42386 ( .A(n42640), .B(n42641), .Z(n779) );
  AND U42387 ( .A(n42642), .B(n42643), .Z(n42641) );
  XNOR U42388 ( .A(p_input[2559]), .B(n42640), .Z(n42643) );
  XOR U42389 ( .A(n42640), .B(p_input[2527]), .Z(n42642) );
  XOR U42390 ( .A(n42644), .B(n42645), .Z(n42640) );
  AND U42391 ( .A(n42646), .B(n42647), .Z(n42645) );
  XNOR U42392 ( .A(p_input[2558]), .B(n42644), .Z(n42647) );
  XOR U42393 ( .A(n42644), .B(p_input[2526]), .Z(n42646) );
  XOR U42394 ( .A(n42648), .B(n42649), .Z(n42644) );
  AND U42395 ( .A(n42650), .B(n42651), .Z(n42649) );
  XNOR U42396 ( .A(p_input[2557]), .B(n42648), .Z(n42651) );
  XOR U42397 ( .A(n42648), .B(p_input[2525]), .Z(n42650) );
  XOR U42398 ( .A(n42652), .B(n42653), .Z(n42648) );
  AND U42399 ( .A(n42654), .B(n42655), .Z(n42653) );
  XNOR U42400 ( .A(p_input[2556]), .B(n42652), .Z(n42655) );
  XOR U42401 ( .A(n42652), .B(p_input[2524]), .Z(n42654) );
  XOR U42402 ( .A(n42656), .B(n42657), .Z(n42652) );
  AND U42403 ( .A(n42658), .B(n42659), .Z(n42657) );
  XNOR U42404 ( .A(p_input[2555]), .B(n42656), .Z(n42659) );
  XOR U42405 ( .A(n42656), .B(p_input[2523]), .Z(n42658) );
  XOR U42406 ( .A(n42660), .B(n42661), .Z(n42656) );
  AND U42407 ( .A(n42662), .B(n42663), .Z(n42661) );
  XNOR U42408 ( .A(p_input[2554]), .B(n42660), .Z(n42663) );
  XOR U42409 ( .A(n42660), .B(p_input[2522]), .Z(n42662) );
  XOR U42410 ( .A(n42664), .B(n42665), .Z(n42660) );
  AND U42411 ( .A(n42666), .B(n42667), .Z(n42665) );
  XNOR U42412 ( .A(p_input[2553]), .B(n42664), .Z(n42667) );
  XOR U42413 ( .A(n42664), .B(p_input[2521]), .Z(n42666) );
  XOR U42414 ( .A(n42668), .B(n42669), .Z(n42664) );
  AND U42415 ( .A(n42670), .B(n42671), .Z(n42669) );
  XNOR U42416 ( .A(p_input[2552]), .B(n42668), .Z(n42671) );
  XOR U42417 ( .A(n42668), .B(p_input[2520]), .Z(n42670) );
  XOR U42418 ( .A(n42672), .B(n42673), .Z(n42668) );
  AND U42419 ( .A(n42674), .B(n42675), .Z(n42673) );
  XNOR U42420 ( .A(p_input[2551]), .B(n42672), .Z(n42675) );
  XOR U42421 ( .A(n42672), .B(p_input[2519]), .Z(n42674) );
  XOR U42422 ( .A(n42676), .B(n42677), .Z(n42672) );
  AND U42423 ( .A(n42678), .B(n42679), .Z(n42677) );
  XNOR U42424 ( .A(p_input[2550]), .B(n42676), .Z(n42679) );
  XOR U42425 ( .A(n42676), .B(p_input[2518]), .Z(n42678) );
  XOR U42426 ( .A(n42680), .B(n42681), .Z(n42676) );
  AND U42427 ( .A(n42682), .B(n42683), .Z(n42681) );
  XNOR U42428 ( .A(p_input[2549]), .B(n42680), .Z(n42683) );
  XOR U42429 ( .A(n42680), .B(p_input[2517]), .Z(n42682) );
  XOR U42430 ( .A(n42684), .B(n42685), .Z(n42680) );
  AND U42431 ( .A(n42686), .B(n42687), .Z(n42685) );
  XNOR U42432 ( .A(p_input[2548]), .B(n42684), .Z(n42687) );
  XOR U42433 ( .A(n42684), .B(p_input[2516]), .Z(n42686) );
  XOR U42434 ( .A(n42688), .B(n42689), .Z(n42684) );
  AND U42435 ( .A(n42690), .B(n42691), .Z(n42689) );
  XNOR U42436 ( .A(p_input[2547]), .B(n42688), .Z(n42691) );
  XOR U42437 ( .A(n42688), .B(p_input[2515]), .Z(n42690) );
  XOR U42438 ( .A(n42692), .B(n42693), .Z(n42688) );
  AND U42439 ( .A(n42694), .B(n42695), .Z(n42693) );
  XNOR U42440 ( .A(p_input[2546]), .B(n42692), .Z(n42695) );
  XOR U42441 ( .A(n42692), .B(p_input[2514]), .Z(n42694) );
  XOR U42442 ( .A(n42696), .B(n42697), .Z(n42692) );
  AND U42443 ( .A(n42698), .B(n42699), .Z(n42697) );
  XNOR U42444 ( .A(p_input[2545]), .B(n42696), .Z(n42699) );
  XOR U42445 ( .A(n42696), .B(p_input[2513]), .Z(n42698) );
  XOR U42446 ( .A(n42700), .B(n42701), .Z(n42696) );
  AND U42447 ( .A(n42702), .B(n42703), .Z(n42701) );
  XNOR U42448 ( .A(p_input[2544]), .B(n42700), .Z(n42703) );
  XOR U42449 ( .A(n42700), .B(p_input[2512]), .Z(n42702) );
  XOR U42450 ( .A(n42704), .B(n42705), .Z(n42700) );
  AND U42451 ( .A(n42706), .B(n42707), .Z(n42705) );
  XNOR U42452 ( .A(p_input[2543]), .B(n42704), .Z(n42707) );
  XOR U42453 ( .A(n42704), .B(p_input[2511]), .Z(n42706) );
  XOR U42454 ( .A(n42708), .B(n42709), .Z(n42704) );
  AND U42455 ( .A(n42710), .B(n42711), .Z(n42709) );
  XNOR U42456 ( .A(p_input[2542]), .B(n42708), .Z(n42711) );
  XOR U42457 ( .A(n42708), .B(p_input[2510]), .Z(n42710) );
  XOR U42458 ( .A(n42712), .B(n42713), .Z(n42708) );
  AND U42459 ( .A(n42714), .B(n42715), .Z(n42713) );
  XNOR U42460 ( .A(p_input[2541]), .B(n42712), .Z(n42715) );
  XOR U42461 ( .A(n42712), .B(p_input[2509]), .Z(n42714) );
  XOR U42462 ( .A(n42716), .B(n42717), .Z(n42712) );
  AND U42463 ( .A(n42718), .B(n42719), .Z(n42717) );
  XNOR U42464 ( .A(p_input[2540]), .B(n42716), .Z(n42719) );
  XOR U42465 ( .A(n42716), .B(p_input[2508]), .Z(n42718) );
  XOR U42466 ( .A(n42720), .B(n42721), .Z(n42716) );
  AND U42467 ( .A(n42722), .B(n42723), .Z(n42721) );
  XNOR U42468 ( .A(p_input[2539]), .B(n42720), .Z(n42723) );
  XOR U42469 ( .A(n42720), .B(p_input[2507]), .Z(n42722) );
  XOR U42470 ( .A(n42724), .B(n42725), .Z(n42720) );
  AND U42471 ( .A(n42726), .B(n42727), .Z(n42725) );
  XNOR U42472 ( .A(p_input[2538]), .B(n42724), .Z(n42727) );
  XOR U42473 ( .A(n42724), .B(p_input[2506]), .Z(n42726) );
  XOR U42474 ( .A(n42728), .B(n42729), .Z(n42724) );
  AND U42475 ( .A(n42730), .B(n42731), .Z(n42729) );
  XNOR U42476 ( .A(p_input[2537]), .B(n42728), .Z(n42731) );
  XOR U42477 ( .A(n42728), .B(p_input[2505]), .Z(n42730) );
  XOR U42478 ( .A(n42732), .B(n42733), .Z(n42728) );
  AND U42479 ( .A(n42734), .B(n42735), .Z(n42733) );
  XNOR U42480 ( .A(p_input[2536]), .B(n42732), .Z(n42735) );
  XOR U42481 ( .A(n42732), .B(p_input[2504]), .Z(n42734) );
  XOR U42482 ( .A(n42736), .B(n42737), .Z(n42732) );
  AND U42483 ( .A(n42738), .B(n42739), .Z(n42737) );
  XNOR U42484 ( .A(p_input[2535]), .B(n42736), .Z(n42739) );
  XOR U42485 ( .A(n42736), .B(p_input[2503]), .Z(n42738) );
  XOR U42486 ( .A(n42740), .B(n42741), .Z(n42736) );
  AND U42487 ( .A(n42742), .B(n42743), .Z(n42741) );
  XNOR U42488 ( .A(p_input[2534]), .B(n42740), .Z(n42743) );
  XOR U42489 ( .A(n42740), .B(p_input[2502]), .Z(n42742) );
  XOR U42490 ( .A(n42744), .B(n42745), .Z(n42740) );
  AND U42491 ( .A(n42746), .B(n42747), .Z(n42745) );
  XNOR U42492 ( .A(p_input[2533]), .B(n42744), .Z(n42747) );
  XOR U42493 ( .A(n42744), .B(p_input[2501]), .Z(n42746) );
  XOR U42494 ( .A(n42748), .B(n42749), .Z(n42744) );
  AND U42495 ( .A(n42750), .B(n42751), .Z(n42749) );
  XNOR U42496 ( .A(p_input[2532]), .B(n42748), .Z(n42751) );
  XOR U42497 ( .A(n42748), .B(p_input[2500]), .Z(n42750) );
  XOR U42498 ( .A(n42752), .B(n42753), .Z(n42748) );
  AND U42499 ( .A(n42754), .B(n42755), .Z(n42753) );
  XNOR U42500 ( .A(p_input[2531]), .B(n42752), .Z(n42755) );
  XOR U42501 ( .A(n42752), .B(p_input[2499]), .Z(n42754) );
  XOR U42502 ( .A(n42756), .B(n42757), .Z(n42752) );
  AND U42503 ( .A(n42758), .B(n42759), .Z(n42757) );
  XNOR U42504 ( .A(p_input[2530]), .B(n42756), .Z(n42759) );
  XOR U42505 ( .A(n42756), .B(p_input[2498]), .Z(n42758) );
  XNOR U42506 ( .A(n42760), .B(n42761), .Z(n42756) );
  AND U42507 ( .A(n42762), .B(n42763), .Z(n42761) );
  XOR U42508 ( .A(p_input[2529]), .B(n42760), .Z(n42763) );
  XNOR U42509 ( .A(p_input[2497]), .B(n42760), .Z(n42762) );
  AND U42510 ( .A(p_input[2528]), .B(n42764), .Z(n42760) );
  IV U42511 ( .A(p_input[2496]), .Z(n42764) );
  XNOR U42512 ( .A(p_input[2432]), .B(n42765), .Z(n42358) );
  AND U42513 ( .A(n777), .B(n42766), .Z(n42765) );
  XOR U42514 ( .A(p_input[2464]), .B(p_input[2432]), .Z(n42766) );
  XOR U42515 ( .A(n42767), .B(n42768), .Z(n777) );
  AND U42516 ( .A(n42769), .B(n42770), .Z(n42768) );
  XNOR U42517 ( .A(p_input[2495]), .B(n42767), .Z(n42770) );
  XOR U42518 ( .A(n42767), .B(p_input[2463]), .Z(n42769) );
  XOR U42519 ( .A(n42771), .B(n42772), .Z(n42767) );
  AND U42520 ( .A(n42773), .B(n42774), .Z(n42772) );
  XNOR U42521 ( .A(p_input[2494]), .B(n42771), .Z(n42774) );
  XNOR U42522 ( .A(n42771), .B(n42373), .Z(n42773) );
  IV U42523 ( .A(p_input[2462]), .Z(n42373) );
  XOR U42524 ( .A(n42775), .B(n42776), .Z(n42771) );
  AND U42525 ( .A(n42777), .B(n42778), .Z(n42776) );
  XNOR U42526 ( .A(p_input[2493]), .B(n42775), .Z(n42778) );
  XNOR U42527 ( .A(n42775), .B(n42382), .Z(n42777) );
  IV U42528 ( .A(p_input[2461]), .Z(n42382) );
  XOR U42529 ( .A(n42779), .B(n42780), .Z(n42775) );
  AND U42530 ( .A(n42781), .B(n42782), .Z(n42780) );
  XNOR U42531 ( .A(p_input[2492]), .B(n42779), .Z(n42782) );
  XNOR U42532 ( .A(n42779), .B(n42391), .Z(n42781) );
  IV U42533 ( .A(p_input[2460]), .Z(n42391) );
  XOR U42534 ( .A(n42783), .B(n42784), .Z(n42779) );
  AND U42535 ( .A(n42785), .B(n42786), .Z(n42784) );
  XNOR U42536 ( .A(p_input[2491]), .B(n42783), .Z(n42786) );
  XNOR U42537 ( .A(n42783), .B(n42400), .Z(n42785) );
  IV U42538 ( .A(p_input[2459]), .Z(n42400) );
  XOR U42539 ( .A(n42787), .B(n42788), .Z(n42783) );
  AND U42540 ( .A(n42789), .B(n42790), .Z(n42788) );
  XNOR U42541 ( .A(p_input[2490]), .B(n42787), .Z(n42790) );
  XNOR U42542 ( .A(n42787), .B(n42409), .Z(n42789) );
  IV U42543 ( .A(p_input[2458]), .Z(n42409) );
  XOR U42544 ( .A(n42791), .B(n42792), .Z(n42787) );
  AND U42545 ( .A(n42793), .B(n42794), .Z(n42792) );
  XNOR U42546 ( .A(p_input[2489]), .B(n42791), .Z(n42794) );
  XNOR U42547 ( .A(n42791), .B(n42418), .Z(n42793) );
  IV U42548 ( .A(p_input[2457]), .Z(n42418) );
  XOR U42549 ( .A(n42795), .B(n42796), .Z(n42791) );
  AND U42550 ( .A(n42797), .B(n42798), .Z(n42796) );
  XNOR U42551 ( .A(p_input[2488]), .B(n42795), .Z(n42798) );
  XNOR U42552 ( .A(n42795), .B(n42427), .Z(n42797) );
  IV U42553 ( .A(p_input[2456]), .Z(n42427) );
  XOR U42554 ( .A(n42799), .B(n42800), .Z(n42795) );
  AND U42555 ( .A(n42801), .B(n42802), .Z(n42800) );
  XNOR U42556 ( .A(p_input[2487]), .B(n42799), .Z(n42802) );
  XNOR U42557 ( .A(n42799), .B(n42436), .Z(n42801) );
  IV U42558 ( .A(p_input[2455]), .Z(n42436) );
  XOR U42559 ( .A(n42803), .B(n42804), .Z(n42799) );
  AND U42560 ( .A(n42805), .B(n42806), .Z(n42804) );
  XNOR U42561 ( .A(p_input[2486]), .B(n42803), .Z(n42806) );
  XNOR U42562 ( .A(n42803), .B(n42445), .Z(n42805) );
  IV U42563 ( .A(p_input[2454]), .Z(n42445) );
  XOR U42564 ( .A(n42807), .B(n42808), .Z(n42803) );
  AND U42565 ( .A(n42809), .B(n42810), .Z(n42808) );
  XNOR U42566 ( .A(p_input[2485]), .B(n42807), .Z(n42810) );
  XNOR U42567 ( .A(n42807), .B(n42454), .Z(n42809) );
  IV U42568 ( .A(p_input[2453]), .Z(n42454) );
  XOR U42569 ( .A(n42811), .B(n42812), .Z(n42807) );
  AND U42570 ( .A(n42813), .B(n42814), .Z(n42812) );
  XNOR U42571 ( .A(p_input[2484]), .B(n42811), .Z(n42814) );
  XNOR U42572 ( .A(n42811), .B(n42463), .Z(n42813) );
  IV U42573 ( .A(p_input[2452]), .Z(n42463) );
  XOR U42574 ( .A(n42815), .B(n42816), .Z(n42811) );
  AND U42575 ( .A(n42817), .B(n42818), .Z(n42816) );
  XNOR U42576 ( .A(p_input[2483]), .B(n42815), .Z(n42818) );
  XNOR U42577 ( .A(n42815), .B(n42472), .Z(n42817) );
  IV U42578 ( .A(p_input[2451]), .Z(n42472) );
  XOR U42579 ( .A(n42819), .B(n42820), .Z(n42815) );
  AND U42580 ( .A(n42821), .B(n42822), .Z(n42820) );
  XNOR U42581 ( .A(p_input[2482]), .B(n42819), .Z(n42822) );
  XNOR U42582 ( .A(n42819), .B(n42481), .Z(n42821) );
  IV U42583 ( .A(p_input[2450]), .Z(n42481) );
  XOR U42584 ( .A(n42823), .B(n42824), .Z(n42819) );
  AND U42585 ( .A(n42825), .B(n42826), .Z(n42824) );
  XNOR U42586 ( .A(p_input[2481]), .B(n42823), .Z(n42826) );
  XNOR U42587 ( .A(n42823), .B(n42490), .Z(n42825) );
  IV U42588 ( .A(p_input[2449]), .Z(n42490) );
  XOR U42589 ( .A(n42827), .B(n42828), .Z(n42823) );
  AND U42590 ( .A(n42829), .B(n42830), .Z(n42828) );
  XNOR U42591 ( .A(p_input[2480]), .B(n42827), .Z(n42830) );
  XNOR U42592 ( .A(n42827), .B(n42499), .Z(n42829) );
  IV U42593 ( .A(p_input[2448]), .Z(n42499) );
  XOR U42594 ( .A(n42831), .B(n42832), .Z(n42827) );
  AND U42595 ( .A(n42833), .B(n42834), .Z(n42832) );
  XNOR U42596 ( .A(p_input[2479]), .B(n42831), .Z(n42834) );
  XNOR U42597 ( .A(n42831), .B(n42508), .Z(n42833) );
  IV U42598 ( .A(p_input[2447]), .Z(n42508) );
  XOR U42599 ( .A(n42835), .B(n42836), .Z(n42831) );
  AND U42600 ( .A(n42837), .B(n42838), .Z(n42836) );
  XNOR U42601 ( .A(p_input[2478]), .B(n42835), .Z(n42838) );
  XNOR U42602 ( .A(n42835), .B(n42517), .Z(n42837) );
  IV U42603 ( .A(p_input[2446]), .Z(n42517) );
  XOR U42604 ( .A(n42839), .B(n42840), .Z(n42835) );
  AND U42605 ( .A(n42841), .B(n42842), .Z(n42840) );
  XNOR U42606 ( .A(p_input[2477]), .B(n42839), .Z(n42842) );
  XNOR U42607 ( .A(n42839), .B(n42526), .Z(n42841) );
  IV U42608 ( .A(p_input[2445]), .Z(n42526) );
  XOR U42609 ( .A(n42843), .B(n42844), .Z(n42839) );
  AND U42610 ( .A(n42845), .B(n42846), .Z(n42844) );
  XNOR U42611 ( .A(p_input[2476]), .B(n42843), .Z(n42846) );
  XNOR U42612 ( .A(n42843), .B(n42535), .Z(n42845) );
  IV U42613 ( .A(p_input[2444]), .Z(n42535) );
  XOR U42614 ( .A(n42847), .B(n42848), .Z(n42843) );
  AND U42615 ( .A(n42849), .B(n42850), .Z(n42848) );
  XNOR U42616 ( .A(p_input[2475]), .B(n42847), .Z(n42850) );
  XNOR U42617 ( .A(n42847), .B(n42544), .Z(n42849) );
  IV U42618 ( .A(p_input[2443]), .Z(n42544) );
  XOR U42619 ( .A(n42851), .B(n42852), .Z(n42847) );
  AND U42620 ( .A(n42853), .B(n42854), .Z(n42852) );
  XNOR U42621 ( .A(p_input[2474]), .B(n42851), .Z(n42854) );
  XNOR U42622 ( .A(n42851), .B(n42553), .Z(n42853) );
  IV U42623 ( .A(p_input[2442]), .Z(n42553) );
  XOR U42624 ( .A(n42855), .B(n42856), .Z(n42851) );
  AND U42625 ( .A(n42857), .B(n42858), .Z(n42856) );
  XNOR U42626 ( .A(p_input[2473]), .B(n42855), .Z(n42858) );
  XNOR U42627 ( .A(n42855), .B(n42562), .Z(n42857) );
  IV U42628 ( .A(p_input[2441]), .Z(n42562) );
  XOR U42629 ( .A(n42859), .B(n42860), .Z(n42855) );
  AND U42630 ( .A(n42861), .B(n42862), .Z(n42860) );
  XNOR U42631 ( .A(p_input[2472]), .B(n42859), .Z(n42862) );
  XNOR U42632 ( .A(n42859), .B(n42571), .Z(n42861) );
  IV U42633 ( .A(p_input[2440]), .Z(n42571) );
  XOR U42634 ( .A(n42863), .B(n42864), .Z(n42859) );
  AND U42635 ( .A(n42865), .B(n42866), .Z(n42864) );
  XNOR U42636 ( .A(p_input[2471]), .B(n42863), .Z(n42866) );
  XNOR U42637 ( .A(n42863), .B(n42580), .Z(n42865) );
  IV U42638 ( .A(p_input[2439]), .Z(n42580) );
  XOR U42639 ( .A(n42867), .B(n42868), .Z(n42863) );
  AND U42640 ( .A(n42869), .B(n42870), .Z(n42868) );
  XNOR U42641 ( .A(p_input[2470]), .B(n42867), .Z(n42870) );
  XNOR U42642 ( .A(n42867), .B(n42589), .Z(n42869) );
  IV U42643 ( .A(p_input[2438]), .Z(n42589) );
  XOR U42644 ( .A(n42871), .B(n42872), .Z(n42867) );
  AND U42645 ( .A(n42873), .B(n42874), .Z(n42872) );
  XNOR U42646 ( .A(p_input[2469]), .B(n42871), .Z(n42874) );
  XNOR U42647 ( .A(n42871), .B(n42598), .Z(n42873) );
  IV U42648 ( .A(p_input[2437]), .Z(n42598) );
  XOR U42649 ( .A(n42875), .B(n42876), .Z(n42871) );
  AND U42650 ( .A(n42877), .B(n42878), .Z(n42876) );
  XNOR U42651 ( .A(p_input[2468]), .B(n42875), .Z(n42878) );
  XNOR U42652 ( .A(n42875), .B(n42607), .Z(n42877) );
  IV U42653 ( .A(p_input[2436]), .Z(n42607) );
  XOR U42654 ( .A(n42879), .B(n42880), .Z(n42875) );
  AND U42655 ( .A(n42881), .B(n42882), .Z(n42880) );
  XNOR U42656 ( .A(p_input[2467]), .B(n42879), .Z(n42882) );
  XNOR U42657 ( .A(n42879), .B(n42616), .Z(n42881) );
  IV U42658 ( .A(p_input[2435]), .Z(n42616) );
  XOR U42659 ( .A(n42883), .B(n42884), .Z(n42879) );
  AND U42660 ( .A(n42885), .B(n42886), .Z(n42884) );
  XNOR U42661 ( .A(p_input[2466]), .B(n42883), .Z(n42886) );
  XNOR U42662 ( .A(n42883), .B(n42625), .Z(n42885) );
  IV U42663 ( .A(p_input[2434]), .Z(n42625) );
  XNOR U42664 ( .A(n42887), .B(n42888), .Z(n42883) );
  AND U42665 ( .A(n42889), .B(n42890), .Z(n42888) );
  XOR U42666 ( .A(p_input[2465]), .B(n42887), .Z(n42890) );
  XNOR U42667 ( .A(p_input[2433]), .B(n42887), .Z(n42889) );
  AND U42668 ( .A(p_input[2464]), .B(n42891), .Z(n42887) );
  IV U42669 ( .A(p_input[2432]), .Z(n42891) );
  XOR U42670 ( .A(n42892), .B(n42893), .Z(n41981) );
  AND U42671 ( .A(n601), .B(n42894), .Z(n42893) );
  XNOR U42672 ( .A(n42895), .B(n42892), .Z(n42894) );
  XOR U42673 ( .A(n42896), .B(n42897), .Z(n601) );
  AND U42674 ( .A(n42898), .B(n42899), .Z(n42897) );
  XNOR U42675 ( .A(n41996), .B(n42896), .Z(n42899) );
  AND U42676 ( .A(p_input[2431]), .B(p_input[2399]), .Z(n41996) );
  XNOR U42677 ( .A(n42896), .B(n41993), .Z(n42898) );
  IV U42678 ( .A(n42900), .Z(n41993) );
  AND U42679 ( .A(p_input[2335]), .B(p_input[2367]), .Z(n42900) );
  XOR U42680 ( .A(n42901), .B(n42902), .Z(n42896) );
  AND U42681 ( .A(n42903), .B(n42904), .Z(n42902) );
  XOR U42682 ( .A(n42901), .B(n42008), .Z(n42904) );
  XNOR U42683 ( .A(p_input[2398]), .B(n42905), .Z(n42008) );
  AND U42684 ( .A(n783), .B(n42906), .Z(n42905) );
  XOR U42685 ( .A(p_input[2430]), .B(p_input[2398]), .Z(n42906) );
  XNOR U42686 ( .A(n42005), .B(n42901), .Z(n42903) );
  XOR U42687 ( .A(n42907), .B(n42908), .Z(n42005) );
  AND U42688 ( .A(n780), .B(n42909), .Z(n42908) );
  XOR U42689 ( .A(p_input[2366]), .B(p_input[2334]), .Z(n42909) );
  XOR U42690 ( .A(n42910), .B(n42911), .Z(n42901) );
  AND U42691 ( .A(n42912), .B(n42913), .Z(n42911) );
  XOR U42692 ( .A(n42910), .B(n42020), .Z(n42913) );
  XNOR U42693 ( .A(p_input[2397]), .B(n42914), .Z(n42020) );
  AND U42694 ( .A(n783), .B(n42915), .Z(n42914) );
  XOR U42695 ( .A(p_input[2429]), .B(p_input[2397]), .Z(n42915) );
  XNOR U42696 ( .A(n42017), .B(n42910), .Z(n42912) );
  XOR U42697 ( .A(n42916), .B(n42917), .Z(n42017) );
  AND U42698 ( .A(n780), .B(n42918), .Z(n42917) );
  XOR U42699 ( .A(p_input[2365]), .B(p_input[2333]), .Z(n42918) );
  XOR U42700 ( .A(n42919), .B(n42920), .Z(n42910) );
  AND U42701 ( .A(n42921), .B(n42922), .Z(n42920) );
  XOR U42702 ( .A(n42919), .B(n42032), .Z(n42922) );
  XNOR U42703 ( .A(p_input[2396]), .B(n42923), .Z(n42032) );
  AND U42704 ( .A(n783), .B(n42924), .Z(n42923) );
  XOR U42705 ( .A(p_input[2428]), .B(p_input[2396]), .Z(n42924) );
  XNOR U42706 ( .A(n42029), .B(n42919), .Z(n42921) );
  XOR U42707 ( .A(n42925), .B(n42926), .Z(n42029) );
  AND U42708 ( .A(n780), .B(n42927), .Z(n42926) );
  XOR U42709 ( .A(p_input[2364]), .B(p_input[2332]), .Z(n42927) );
  XOR U42710 ( .A(n42928), .B(n42929), .Z(n42919) );
  AND U42711 ( .A(n42930), .B(n42931), .Z(n42929) );
  XOR U42712 ( .A(n42928), .B(n42044), .Z(n42931) );
  XNOR U42713 ( .A(p_input[2395]), .B(n42932), .Z(n42044) );
  AND U42714 ( .A(n783), .B(n42933), .Z(n42932) );
  XOR U42715 ( .A(p_input[2427]), .B(p_input[2395]), .Z(n42933) );
  XNOR U42716 ( .A(n42041), .B(n42928), .Z(n42930) );
  XOR U42717 ( .A(n42934), .B(n42935), .Z(n42041) );
  AND U42718 ( .A(n780), .B(n42936), .Z(n42935) );
  XOR U42719 ( .A(p_input[2363]), .B(p_input[2331]), .Z(n42936) );
  XOR U42720 ( .A(n42937), .B(n42938), .Z(n42928) );
  AND U42721 ( .A(n42939), .B(n42940), .Z(n42938) );
  XOR U42722 ( .A(n42937), .B(n42056), .Z(n42940) );
  XNOR U42723 ( .A(p_input[2394]), .B(n42941), .Z(n42056) );
  AND U42724 ( .A(n783), .B(n42942), .Z(n42941) );
  XOR U42725 ( .A(p_input[2426]), .B(p_input[2394]), .Z(n42942) );
  XNOR U42726 ( .A(n42053), .B(n42937), .Z(n42939) );
  XOR U42727 ( .A(n42943), .B(n42944), .Z(n42053) );
  AND U42728 ( .A(n780), .B(n42945), .Z(n42944) );
  XOR U42729 ( .A(p_input[2362]), .B(p_input[2330]), .Z(n42945) );
  XOR U42730 ( .A(n42946), .B(n42947), .Z(n42937) );
  AND U42731 ( .A(n42948), .B(n42949), .Z(n42947) );
  XOR U42732 ( .A(n42946), .B(n42068), .Z(n42949) );
  XNOR U42733 ( .A(p_input[2393]), .B(n42950), .Z(n42068) );
  AND U42734 ( .A(n783), .B(n42951), .Z(n42950) );
  XOR U42735 ( .A(p_input[2425]), .B(p_input[2393]), .Z(n42951) );
  XNOR U42736 ( .A(n42065), .B(n42946), .Z(n42948) );
  XOR U42737 ( .A(n42952), .B(n42953), .Z(n42065) );
  AND U42738 ( .A(n780), .B(n42954), .Z(n42953) );
  XOR U42739 ( .A(p_input[2361]), .B(p_input[2329]), .Z(n42954) );
  XOR U42740 ( .A(n42955), .B(n42956), .Z(n42946) );
  AND U42741 ( .A(n42957), .B(n42958), .Z(n42956) );
  XOR U42742 ( .A(n42955), .B(n42080), .Z(n42958) );
  XNOR U42743 ( .A(p_input[2392]), .B(n42959), .Z(n42080) );
  AND U42744 ( .A(n783), .B(n42960), .Z(n42959) );
  XOR U42745 ( .A(p_input[2424]), .B(p_input[2392]), .Z(n42960) );
  XNOR U42746 ( .A(n42077), .B(n42955), .Z(n42957) );
  XOR U42747 ( .A(n42961), .B(n42962), .Z(n42077) );
  AND U42748 ( .A(n780), .B(n42963), .Z(n42962) );
  XOR U42749 ( .A(p_input[2360]), .B(p_input[2328]), .Z(n42963) );
  XOR U42750 ( .A(n42964), .B(n42965), .Z(n42955) );
  AND U42751 ( .A(n42966), .B(n42967), .Z(n42965) );
  XOR U42752 ( .A(n42964), .B(n42092), .Z(n42967) );
  XNOR U42753 ( .A(p_input[2391]), .B(n42968), .Z(n42092) );
  AND U42754 ( .A(n783), .B(n42969), .Z(n42968) );
  XOR U42755 ( .A(p_input[2423]), .B(p_input[2391]), .Z(n42969) );
  XNOR U42756 ( .A(n42089), .B(n42964), .Z(n42966) );
  XOR U42757 ( .A(n42970), .B(n42971), .Z(n42089) );
  AND U42758 ( .A(n780), .B(n42972), .Z(n42971) );
  XOR U42759 ( .A(p_input[2359]), .B(p_input[2327]), .Z(n42972) );
  XOR U42760 ( .A(n42973), .B(n42974), .Z(n42964) );
  AND U42761 ( .A(n42975), .B(n42976), .Z(n42974) );
  XOR U42762 ( .A(n42973), .B(n42104), .Z(n42976) );
  XNOR U42763 ( .A(p_input[2390]), .B(n42977), .Z(n42104) );
  AND U42764 ( .A(n783), .B(n42978), .Z(n42977) );
  XOR U42765 ( .A(p_input[2422]), .B(p_input[2390]), .Z(n42978) );
  XNOR U42766 ( .A(n42101), .B(n42973), .Z(n42975) );
  XOR U42767 ( .A(n42979), .B(n42980), .Z(n42101) );
  AND U42768 ( .A(n780), .B(n42981), .Z(n42980) );
  XOR U42769 ( .A(p_input[2358]), .B(p_input[2326]), .Z(n42981) );
  XOR U42770 ( .A(n42982), .B(n42983), .Z(n42973) );
  AND U42771 ( .A(n42984), .B(n42985), .Z(n42983) );
  XOR U42772 ( .A(n42982), .B(n42116), .Z(n42985) );
  XNOR U42773 ( .A(p_input[2389]), .B(n42986), .Z(n42116) );
  AND U42774 ( .A(n783), .B(n42987), .Z(n42986) );
  XOR U42775 ( .A(p_input[2421]), .B(p_input[2389]), .Z(n42987) );
  XNOR U42776 ( .A(n42113), .B(n42982), .Z(n42984) );
  XOR U42777 ( .A(n42988), .B(n42989), .Z(n42113) );
  AND U42778 ( .A(n780), .B(n42990), .Z(n42989) );
  XOR U42779 ( .A(p_input[2357]), .B(p_input[2325]), .Z(n42990) );
  XOR U42780 ( .A(n42991), .B(n42992), .Z(n42982) );
  AND U42781 ( .A(n42993), .B(n42994), .Z(n42992) );
  XOR U42782 ( .A(n42991), .B(n42128), .Z(n42994) );
  XNOR U42783 ( .A(p_input[2388]), .B(n42995), .Z(n42128) );
  AND U42784 ( .A(n783), .B(n42996), .Z(n42995) );
  XOR U42785 ( .A(p_input[2420]), .B(p_input[2388]), .Z(n42996) );
  XNOR U42786 ( .A(n42125), .B(n42991), .Z(n42993) );
  XOR U42787 ( .A(n42997), .B(n42998), .Z(n42125) );
  AND U42788 ( .A(n780), .B(n42999), .Z(n42998) );
  XOR U42789 ( .A(p_input[2356]), .B(p_input[2324]), .Z(n42999) );
  XOR U42790 ( .A(n43000), .B(n43001), .Z(n42991) );
  AND U42791 ( .A(n43002), .B(n43003), .Z(n43001) );
  XOR U42792 ( .A(n43000), .B(n42140), .Z(n43003) );
  XNOR U42793 ( .A(p_input[2387]), .B(n43004), .Z(n42140) );
  AND U42794 ( .A(n783), .B(n43005), .Z(n43004) );
  XOR U42795 ( .A(p_input[2419]), .B(p_input[2387]), .Z(n43005) );
  XNOR U42796 ( .A(n42137), .B(n43000), .Z(n43002) );
  XOR U42797 ( .A(n43006), .B(n43007), .Z(n42137) );
  AND U42798 ( .A(n780), .B(n43008), .Z(n43007) );
  XOR U42799 ( .A(p_input[2355]), .B(p_input[2323]), .Z(n43008) );
  XOR U42800 ( .A(n43009), .B(n43010), .Z(n43000) );
  AND U42801 ( .A(n43011), .B(n43012), .Z(n43010) );
  XOR U42802 ( .A(n43009), .B(n42152), .Z(n43012) );
  XNOR U42803 ( .A(p_input[2386]), .B(n43013), .Z(n42152) );
  AND U42804 ( .A(n783), .B(n43014), .Z(n43013) );
  XOR U42805 ( .A(p_input[2418]), .B(p_input[2386]), .Z(n43014) );
  XNOR U42806 ( .A(n42149), .B(n43009), .Z(n43011) );
  XOR U42807 ( .A(n43015), .B(n43016), .Z(n42149) );
  AND U42808 ( .A(n780), .B(n43017), .Z(n43016) );
  XOR U42809 ( .A(p_input[2354]), .B(p_input[2322]), .Z(n43017) );
  XOR U42810 ( .A(n43018), .B(n43019), .Z(n43009) );
  AND U42811 ( .A(n43020), .B(n43021), .Z(n43019) );
  XOR U42812 ( .A(n43018), .B(n42164), .Z(n43021) );
  XNOR U42813 ( .A(p_input[2385]), .B(n43022), .Z(n42164) );
  AND U42814 ( .A(n783), .B(n43023), .Z(n43022) );
  XOR U42815 ( .A(p_input[2417]), .B(p_input[2385]), .Z(n43023) );
  XNOR U42816 ( .A(n42161), .B(n43018), .Z(n43020) );
  XOR U42817 ( .A(n43024), .B(n43025), .Z(n42161) );
  AND U42818 ( .A(n780), .B(n43026), .Z(n43025) );
  XOR U42819 ( .A(p_input[2353]), .B(p_input[2321]), .Z(n43026) );
  XOR U42820 ( .A(n43027), .B(n43028), .Z(n43018) );
  AND U42821 ( .A(n43029), .B(n43030), .Z(n43028) );
  XOR U42822 ( .A(n43027), .B(n42176), .Z(n43030) );
  XNOR U42823 ( .A(p_input[2384]), .B(n43031), .Z(n42176) );
  AND U42824 ( .A(n783), .B(n43032), .Z(n43031) );
  XOR U42825 ( .A(p_input[2416]), .B(p_input[2384]), .Z(n43032) );
  XNOR U42826 ( .A(n42173), .B(n43027), .Z(n43029) );
  XOR U42827 ( .A(n43033), .B(n43034), .Z(n42173) );
  AND U42828 ( .A(n780), .B(n43035), .Z(n43034) );
  XOR U42829 ( .A(p_input[2352]), .B(p_input[2320]), .Z(n43035) );
  XOR U42830 ( .A(n43036), .B(n43037), .Z(n43027) );
  AND U42831 ( .A(n43038), .B(n43039), .Z(n43037) );
  XOR U42832 ( .A(n43036), .B(n42188), .Z(n43039) );
  XNOR U42833 ( .A(p_input[2383]), .B(n43040), .Z(n42188) );
  AND U42834 ( .A(n783), .B(n43041), .Z(n43040) );
  XOR U42835 ( .A(p_input[2415]), .B(p_input[2383]), .Z(n43041) );
  XNOR U42836 ( .A(n42185), .B(n43036), .Z(n43038) );
  XOR U42837 ( .A(n43042), .B(n43043), .Z(n42185) );
  AND U42838 ( .A(n780), .B(n43044), .Z(n43043) );
  XOR U42839 ( .A(p_input[2351]), .B(p_input[2319]), .Z(n43044) );
  XOR U42840 ( .A(n43045), .B(n43046), .Z(n43036) );
  AND U42841 ( .A(n43047), .B(n43048), .Z(n43046) );
  XOR U42842 ( .A(n43045), .B(n42200), .Z(n43048) );
  XNOR U42843 ( .A(p_input[2382]), .B(n43049), .Z(n42200) );
  AND U42844 ( .A(n783), .B(n43050), .Z(n43049) );
  XOR U42845 ( .A(p_input[2414]), .B(p_input[2382]), .Z(n43050) );
  XNOR U42846 ( .A(n42197), .B(n43045), .Z(n43047) );
  XOR U42847 ( .A(n43051), .B(n43052), .Z(n42197) );
  AND U42848 ( .A(n780), .B(n43053), .Z(n43052) );
  XOR U42849 ( .A(p_input[2350]), .B(p_input[2318]), .Z(n43053) );
  XOR U42850 ( .A(n43054), .B(n43055), .Z(n43045) );
  AND U42851 ( .A(n43056), .B(n43057), .Z(n43055) );
  XOR U42852 ( .A(n43054), .B(n42212), .Z(n43057) );
  XNOR U42853 ( .A(p_input[2381]), .B(n43058), .Z(n42212) );
  AND U42854 ( .A(n783), .B(n43059), .Z(n43058) );
  XOR U42855 ( .A(p_input[2413]), .B(p_input[2381]), .Z(n43059) );
  XNOR U42856 ( .A(n42209), .B(n43054), .Z(n43056) );
  XOR U42857 ( .A(n43060), .B(n43061), .Z(n42209) );
  AND U42858 ( .A(n780), .B(n43062), .Z(n43061) );
  XOR U42859 ( .A(p_input[2349]), .B(p_input[2317]), .Z(n43062) );
  XOR U42860 ( .A(n43063), .B(n43064), .Z(n43054) );
  AND U42861 ( .A(n43065), .B(n43066), .Z(n43064) );
  XOR U42862 ( .A(n43063), .B(n42224), .Z(n43066) );
  XNOR U42863 ( .A(p_input[2380]), .B(n43067), .Z(n42224) );
  AND U42864 ( .A(n783), .B(n43068), .Z(n43067) );
  XOR U42865 ( .A(p_input[2412]), .B(p_input[2380]), .Z(n43068) );
  XNOR U42866 ( .A(n42221), .B(n43063), .Z(n43065) );
  XOR U42867 ( .A(n43069), .B(n43070), .Z(n42221) );
  AND U42868 ( .A(n780), .B(n43071), .Z(n43070) );
  XOR U42869 ( .A(p_input[2348]), .B(p_input[2316]), .Z(n43071) );
  XOR U42870 ( .A(n43072), .B(n43073), .Z(n43063) );
  AND U42871 ( .A(n43074), .B(n43075), .Z(n43073) );
  XOR U42872 ( .A(n43072), .B(n42236), .Z(n43075) );
  XNOR U42873 ( .A(p_input[2379]), .B(n43076), .Z(n42236) );
  AND U42874 ( .A(n783), .B(n43077), .Z(n43076) );
  XOR U42875 ( .A(p_input[2411]), .B(p_input[2379]), .Z(n43077) );
  XNOR U42876 ( .A(n42233), .B(n43072), .Z(n43074) );
  XOR U42877 ( .A(n43078), .B(n43079), .Z(n42233) );
  AND U42878 ( .A(n780), .B(n43080), .Z(n43079) );
  XOR U42879 ( .A(p_input[2347]), .B(p_input[2315]), .Z(n43080) );
  XOR U42880 ( .A(n43081), .B(n43082), .Z(n43072) );
  AND U42881 ( .A(n43083), .B(n43084), .Z(n43082) );
  XOR U42882 ( .A(n43081), .B(n42248), .Z(n43084) );
  XNOR U42883 ( .A(p_input[2378]), .B(n43085), .Z(n42248) );
  AND U42884 ( .A(n783), .B(n43086), .Z(n43085) );
  XOR U42885 ( .A(p_input[2410]), .B(p_input[2378]), .Z(n43086) );
  XNOR U42886 ( .A(n42245), .B(n43081), .Z(n43083) );
  XOR U42887 ( .A(n43087), .B(n43088), .Z(n42245) );
  AND U42888 ( .A(n780), .B(n43089), .Z(n43088) );
  XOR U42889 ( .A(p_input[2346]), .B(p_input[2314]), .Z(n43089) );
  XOR U42890 ( .A(n43090), .B(n43091), .Z(n43081) );
  AND U42891 ( .A(n43092), .B(n43093), .Z(n43091) );
  XOR U42892 ( .A(n43090), .B(n42260), .Z(n43093) );
  XNOR U42893 ( .A(p_input[2377]), .B(n43094), .Z(n42260) );
  AND U42894 ( .A(n783), .B(n43095), .Z(n43094) );
  XOR U42895 ( .A(p_input[2409]), .B(p_input[2377]), .Z(n43095) );
  XNOR U42896 ( .A(n42257), .B(n43090), .Z(n43092) );
  XOR U42897 ( .A(n43096), .B(n43097), .Z(n42257) );
  AND U42898 ( .A(n780), .B(n43098), .Z(n43097) );
  XOR U42899 ( .A(p_input[2345]), .B(p_input[2313]), .Z(n43098) );
  XOR U42900 ( .A(n43099), .B(n43100), .Z(n43090) );
  AND U42901 ( .A(n43101), .B(n43102), .Z(n43100) );
  XOR U42902 ( .A(n43099), .B(n42272), .Z(n43102) );
  XNOR U42903 ( .A(p_input[2376]), .B(n43103), .Z(n42272) );
  AND U42904 ( .A(n783), .B(n43104), .Z(n43103) );
  XOR U42905 ( .A(p_input[2408]), .B(p_input[2376]), .Z(n43104) );
  XNOR U42906 ( .A(n42269), .B(n43099), .Z(n43101) );
  XOR U42907 ( .A(n43105), .B(n43106), .Z(n42269) );
  AND U42908 ( .A(n780), .B(n43107), .Z(n43106) );
  XOR U42909 ( .A(p_input[2344]), .B(p_input[2312]), .Z(n43107) );
  XOR U42910 ( .A(n43108), .B(n43109), .Z(n43099) );
  AND U42911 ( .A(n43110), .B(n43111), .Z(n43109) );
  XOR U42912 ( .A(n43108), .B(n42284), .Z(n43111) );
  XNOR U42913 ( .A(p_input[2375]), .B(n43112), .Z(n42284) );
  AND U42914 ( .A(n783), .B(n43113), .Z(n43112) );
  XOR U42915 ( .A(p_input[2407]), .B(p_input[2375]), .Z(n43113) );
  XNOR U42916 ( .A(n42281), .B(n43108), .Z(n43110) );
  XOR U42917 ( .A(n43114), .B(n43115), .Z(n42281) );
  AND U42918 ( .A(n780), .B(n43116), .Z(n43115) );
  XOR U42919 ( .A(p_input[2343]), .B(p_input[2311]), .Z(n43116) );
  XOR U42920 ( .A(n43117), .B(n43118), .Z(n43108) );
  AND U42921 ( .A(n43119), .B(n43120), .Z(n43118) );
  XOR U42922 ( .A(n43117), .B(n42296), .Z(n43120) );
  XNOR U42923 ( .A(p_input[2374]), .B(n43121), .Z(n42296) );
  AND U42924 ( .A(n783), .B(n43122), .Z(n43121) );
  XOR U42925 ( .A(p_input[2406]), .B(p_input[2374]), .Z(n43122) );
  XNOR U42926 ( .A(n42293), .B(n43117), .Z(n43119) );
  XOR U42927 ( .A(n43123), .B(n43124), .Z(n42293) );
  AND U42928 ( .A(n780), .B(n43125), .Z(n43124) );
  XOR U42929 ( .A(p_input[2342]), .B(p_input[2310]), .Z(n43125) );
  XOR U42930 ( .A(n43126), .B(n43127), .Z(n43117) );
  AND U42931 ( .A(n43128), .B(n43129), .Z(n43127) );
  XOR U42932 ( .A(n43126), .B(n42308), .Z(n43129) );
  XNOR U42933 ( .A(p_input[2373]), .B(n43130), .Z(n42308) );
  AND U42934 ( .A(n783), .B(n43131), .Z(n43130) );
  XOR U42935 ( .A(p_input[2405]), .B(p_input[2373]), .Z(n43131) );
  XNOR U42936 ( .A(n42305), .B(n43126), .Z(n43128) );
  XOR U42937 ( .A(n43132), .B(n43133), .Z(n42305) );
  AND U42938 ( .A(n780), .B(n43134), .Z(n43133) );
  XOR U42939 ( .A(p_input[2341]), .B(p_input[2309]), .Z(n43134) );
  XOR U42940 ( .A(n43135), .B(n43136), .Z(n43126) );
  AND U42941 ( .A(n43137), .B(n43138), .Z(n43136) );
  XOR U42942 ( .A(n43135), .B(n42320), .Z(n43138) );
  XNOR U42943 ( .A(p_input[2372]), .B(n43139), .Z(n42320) );
  AND U42944 ( .A(n783), .B(n43140), .Z(n43139) );
  XOR U42945 ( .A(p_input[2404]), .B(p_input[2372]), .Z(n43140) );
  XNOR U42946 ( .A(n42317), .B(n43135), .Z(n43137) );
  XOR U42947 ( .A(n43141), .B(n43142), .Z(n42317) );
  AND U42948 ( .A(n780), .B(n43143), .Z(n43142) );
  XOR U42949 ( .A(p_input[2340]), .B(p_input[2308]), .Z(n43143) );
  XOR U42950 ( .A(n43144), .B(n43145), .Z(n43135) );
  AND U42951 ( .A(n43146), .B(n43147), .Z(n43145) );
  XOR U42952 ( .A(n43144), .B(n42332), .Z(n43147) );
  XNOR U42953 ( .A(p_input[2371]), .B(n43148), .Z(n42332) );
  AND U42954 ( .A(n783), .B(n43149), .Z(n43148) );
  XOR U42955 ( .A(p_input[2403]), .B(p_input[2371]), .Z(n43149) );
  XNOR U42956 ( .A(n42329), .B(n43144), .Z(n43146) );
  XOR U42957 ( .A(n43150), .B(n43151), .Z(n42329) );
  AND U42958 ( .A(n780), .B(n43152), .Z(n43151) );
  XOR U42959 ( .A(p_input[2339]), .B(p_input[2307]), .Z(n43152) );
  XOR U42960 ( .A(n43153), .B(n43154), .Z(n43144) );
  AND U42961 ( .A(n43155), .B(n43156), .Z(n43154) );
  XOR U42962 ( .A(n43153), .B(n42344), .Z(n43156) );
  XNOR U42963 ( .A(p_input[2370]), .B(n43157), .Z(n42344) );
  AND U42964 ( .A(n783), .B(n43158), .Z(n43157) );
  XOR U42965 ( .A(p_input[2402]), .B(p_input[2370]), .Z(n43158) );
  XNOR U42966 ( .A(n42341), .B(n43153), .Z(n43155) );
  XOR U42967 ( .A(n43159), .B(n43160), .Z(n42341) );
  AND U42968 ( .A(n780), .B(n43161), .Z(n43160) );
  XOR U42969 ( .A(p_input[2338]), .B(p_input[2306]), .Z(n43161) );
  XOR U42970 ( .A(n43162), .B(n43163), .Z(n43153) );
  AND U42971 ( .A(n43164), .B(n43165), .Z(n43163) );
  XNOR U42972 ( .A(n43166), .B(n42357), .Z(n43165) );
  XNOR U42973 ( .A(p_input[2369]), .B(n43167), .Z(n42357) );
  AND U42974 ( .A(n783), .B(n43168), .Z(n43167) );
  XNOR U42975 ( .A(p_input[2401]), .B(n43169), .Z(n43168) );
  IV U42976 ( .A(p_input[2369]), .Z(n43169) );
  XNOR U42977 ( .A(n42354), .B(n43162), .Z(n43164) );
  XNOR U42978 ( .A(p_input[2305]), .B(n43170), .Z(n42354) );
  AND U42979 ( .A(n780), .B(n43171), .Z(n43170) );
  XOR U42980 ( .A(p_input[2337]), .B(p_input[2305]), .Z(n43171) );
  IV U42981 ( .A(n43166), .Z(n43162) );
  AND U42982 ( .A(n42892), .B(n42895), .Z(n43166) );
  XOR U42983 ( .A(p_input[2368]), .B(n43172), .Z(n42895) );
  AND U42984 ( .A(n783), .B(n43173), .Z(n43172) );
  XOR U42985 ( .A(p_input[2400]), .B(p_input[2368]), .Z(n43173) );
  XOR U42986 ( .A(n43174), .B(n43175), .Z(n783) );
  AND U42987 ( .A(n43176), .B(n43177), .Z(n43175) );
  XNOR U42988 ( .A(p_input[2431]), .B(n43174), .Z(n43177) );
  XOR U42989 ( .A(n43174), .B(p_input[2399]), .Z(n43176) );
  XOR U42990 ( .A(n43178), .B(n43179), .Z(n43174) );
  AND U42991 ( .A(n43180), .B(n43181), .Z(n43179) );
  XNOR U42992 ( .A(p_input[2430]), .B(n43178), .Z(n43181) );
  XOR U42993 ( .A(n43178), .B(p_input[2398]), .Z(n43180) );
  XOR U42994 ( .A(n43182), .B(n43183), .Z(n43178) );
  AND U42995 ( .A(n43184), .B(n43185), .Z(n43183) );
  XNOR U42996 ( .A(p_input[2429]), .B(n43182), .Z(n43185) );
  XOR U42997 ( .A(n43182), .B(p_input[2397]), .Z(n43184) );
  XOR U42998 ( .A(n43186), .B(n43187), .Z(n43182) );
  AND U42999 ( .A(n43188), .B(n43189), .Z(n43187) );
  XNOR U43000 ( .A(p_input[2428]), .B(n43186), .Z(n43189) );
  XOR U43001 ( .A(n43186), .B(p_input[2396]), .Z(n43188) );
  XOR U43002 ( .A(n43190), .B(n43191), .Z(n43186) );
  AND U43003 ( .A(n43192), .B(n43193), .Z(n43191) );
  XNOR U43004 ( .A(p_input[2427]), .B(n43190), .Z(n43193) );
  XOR U43005 ( .A(n43190), .B(p_input[2395]), .Z(n43192) );
  XOR U43006 ( .A(n43194), .B(n43195), .Z(n43190) );
  AND U43007 ( .A(n43196), .B(n43197), .Z(n43195) );
  XNOR U43008 ( .A(p_input[2426]), .B(n43194), .Z(n43197) );
  XOR U43009 ( .A(n43194), .B(p_input[2394]), .Z(n43196) );
  XOR U43010 ( .A(n43198), .B(n43199), .Z(n43194) );
  AND U43011 ( .A(n43200), .B(n43201), .Z(n43199) );
  XNOR U43012 ( .A(p_input[2425]), .B(n43198), .Z(n43201) );
  XOR U43013 ( .A(n43198), .B(p_input[2393]), .Z(n43200) );
  XOR U43014 ( .A(n43202), .B(n43203), .Z(n43198) );
  AND U43015 ( .A(n43204), .B(n43205), .Z(n43203) );
  XNOR U43016 ( .A(p_input[2424]), .B(n43202), .Z(n43205) );
  XOR U43017 ( .A(n43202), .B(p_input[2392]), .Z(n43204) );
  XOR U43018 ( .A(n43206), .B(n43207), .Z(n43202) );
  AND U43019 ( .A(n43208), .B(n43209), .Z(n43207) );
  XNOR U43020 ( .A(p_input[2423]), .B(n43206), .Z(n43209) );
  XOR U43021 ( .A(n43206), .B(p_input[2391]), .Z(n43208) );
  XOR U43022 ( .A(n43210), .B(n43211), .Z(n43206) );
  AND U43023 ( .A(n43212), .B(n43213), .Z(n43211) );
  XNOR U43024 ( .A(p_input[2422]), .B(n43210), .Z(n43213) );
  XOR U43025 ( .A(n43210), .B(p_input[2390]), .Z(n43212) );
  XOR U43026 ( .A(n43214), .B(n43215), .Z(n43210) );
  AND U43027 ( .A(n43216), .B(n43217), .Z(n43215) );
  XNOR U43028 ( .A(p_input[2421]), .B(n43214), .Z(n43217) );
  XOR U43029 ( .A(n43214), .B(p_input[2389]), .Z(n43216) );
  XOR U43030 ( .A(n43218), .B(n43219), .Z(n43214) );
  AND U43031 ( .A(n43220), .B(n43221), .Z(n43219) );
  XNOR U43032 ( .A(p_input[2420]), .B(n43218), .Z(n43221) );
  XOR U43033 ( .A(n43218), .B(p_input[2388]), .Z(n43220) );
  XOR U43034 ( .A(n43222), .B(n43223), .Z(n43218) );
  AND U43035 ( .A(n43224), .B(n43225), .Z(n43223) );
  XNOR U43036 ( .A(p_input[2419]), .B(n43222), .Z(n43225) );
  XOR U43037 ( .A(n43222), .B(p_input[2387]), .Z(n43224) );
  XOR U43038 ( .A(n43226), .B(n43227), .Z(n43222) );
  AND U43039 ( .A(n43228), .B(n43229), .Z(n43227) );
  XNOR U43040 ( .A(p_input[2418]), .B(n43226), .Z(n43229) );
  XOR U43041 ( .A(n43226), .B(p_input[2386]), .Z(n43228) );
  XOR U43042 ( .A(n43230), .B(n43231), .Z(n43226) );
  AND U43043 ( .A(n43232), .B(n43233), .Z(n43231) );
  XNOR U43044 ( .A(p_input[2417]), .B(n43230), .Z(n43233) );
  XOR U43045 ( .A(n43230), .B(p_input[2385]), .Z(n43232) );
  XOR U43046 ( .A(n43234), .B(n43235), .Z(n43230) );
  AND U43047 ( .A(n43236), .B(n43237), .Z(n43235) );
  XNOR U43048 ( .A(p_input[2416]), .B(n43234), .Z(n43237) );
  XOR U43049 ( .A(n43234), .B(p_input[2384]), .Z(n43236) );
  XOR U43050 ( .A(n43238), .B(n43239), .Z(n43234) );
  AND U43051 ( .A(n43240), .B(n43241), .Z(n43239) );
  XNOR U43052 ( .A(p_input[2415]), .B(n43238), .Z(n43241) );
  XOR U43053 ( .A(n43238), .B(p_input[2383]), .Z(n43240) );
  XOR U43054 ( .A(n43242), .B(n43243), .Z(n43238) );
  AND U43055 ( .A(n43244), .B(n43245), .Z(n43243) );
  XNOR U43056 ( .A(p_input[2414]), .B(n43242), .Z(n43245) );
  XOR U43057 ( .A(n43242), .B(p_input[2382]), .Z(n43244) );
  XOR U43058 ( .A(n43246), .B(n43247), .Z(n43242) );
  AND U43059 ( .A(n43248), .B(n43249), .Z(n43247) );
  XNOR U43060 ( .A(p_input[2413]), .B(n43246), .Z(n43249) );
  XOR U43061 ( .A(n43246), .B(p_input[2381]), .Z(n43248) );
  XOR U43062 ( .A(n43250), .B(n43251), .Z(n43246) );
  AND U43063 ( .A(n43252), .B(n43253), .Z(n43251) );
  XNOR U43064 ( .A(p_input[2412]), .B(n43250), .Z(n43253) );
  XOR U43065 ( .A(n43250), .B(p_input[2380]), .Z(n43252) );
  XOR U43066 ( .A(n43254), .B(n43255), .Z(n43250) );
  AND U43067 ( .A(n43256), .B(n43257), .Z(n43255) );
  XNOR U43068 ( .A(p_input[2411]), .B(n43254), .Z(n43257) );
  XOR U43069 ( .A(n43254), .B(p_input[2379]), .Z(n43256) );
  XOR U43070 ( .A(n43258), .B(n43259), .Z(n43254) );
  AND U43071 ( .A(n43260), .B(n43261), .Z(n43259) );
  XNOR U43072 ( .A(p_input[2410]), .B(n43258), .Z(n43261) );
  XOR U43073 ( .A(n43258), .B(p_input[2378]), .Z(n43260) );
  XOR U43074 ( .A(n43262), .B(n43263), .Z(n43258) );
  AND U43075 ( .A(n43264), .B(n43265), .Z(n43263) );
  XNOR U43076 ( .A(p_input[2409]), .B(n43262), .Z(n43265) );
  XOR U43077 ( .A(n43262), .B(p_input[2377]), .Z(n43264) );
  XOR U43078 ( .A(n43266), .B(n43267), .Z(n43262) );
  AND U43079 ( .A(n43268), .B(n43269), .Z(n43267) );
  XNOR U43080 ( .A(p_input[2408]), .B(n43266), .Z(n43269) );
  XOR U43081 ( .A(n43266), .B(p_input[2376]), .Z(n43268) );
  XOR U43082 ( .A(n43270), .B(n43271), .Z(n43266) );
  AND U43083 ( .A(n43272), .B(n43273), .Z(n43271) );
  XNOR U43084 ( .A(p_input[2407]), .B(n43270), .Z(n43273) );
  XOR U43085 ( .A(n43270), .B(p_input[2375]), .Z(n43272) );
  XOR U43086 ( .A(n43274), .B(n43275), .Z(n43270) );
  AND U43087 ( .A(n43276), .B(n43277), .Z(n43275) );
  XNOR U43088 ( .A(p_input[2406]), .B(n43274), .Z(n43277) );
  XOR U43089 ( .A(n43274), .B(p_input[2374]), .Z(n43276) );
  XOR U43090 ( .A(n43278), .B(n43279), .Z(n43274) );
  AND U43091 ( .A(n43280), .B(n43281), .Z(n43279) );
  XNOR U43092 ( .A(p_input[2405]), .B(n43278), .Z(n43281) );
  XOR U43093 ( .A(n43278), .B(p_input[2373]), .Z(n43280) );
  XOR U43094 ( .A(n43282), .B(n43283), .Z(n43278) );
  AND U43095 ( .A(n43284), .B(n43285), .Z(n43283) );
  XNOR U43096 ( .A(p_input[2404]), .B(n43282), .Z(n43285) );
  XOR U43097 ( .A(n43282), .B(p_input[2372]), .Z(n43284) );
  XOR U43098 ( .A(n43286), .B(n43287), .Z(n43282) );
  AND U43099 ( .A(n43288), .B(n43289), .Z(n43287) );
  XNOR U43100 ( .A(p_input[2403]), .B(n43286), .Z(n43289) );
  XOR U43101 ( .A(n43286), .B(p_input[2371]), .Z(n43288) );
  XOR U43102 ( .A(n43290), .B(n43291), .Z(n43286) );
  AND U43103 ( .A(n43292), .B(n43293), .Z(n43291) );
  XNOR U43104 ( .A(p_input[2402]), .B(n43290), .Z(n43293) );
  XOR U43105 ( .A(n43290), .B(p_input[2370]), .Z(n43292) );
  XNOR U43106 ( .A(n43294), .B(n43295), .Z(n43290) );
  AND U43107 ( .A(n43296), .B(n43297), .Z(n43295) );
  XOR U43108 ( .A(p_input[2401]), .B(n43294), .Z(n43297) );
  XNOR U43109 ( .A(p_input[2369]), .B(n43294), .Z(n43296) );
  AND U43110 ( .A(p_input[2400]), .B(n43298), .Z(n43294) );
  IV U43111 ( .A(p_input[2368]), .Z(n43298) );
  XNOR U43112 ( .A(p_input[2304]), .B(n43299), .Z(n42892) );
  AND U43113 ( .A(n780), .B(n43300), .Z(n43299) );
  XOR U43114 ( .A(p_input[2336]), .B(p_input[2304]), .Z(n43300) );
  XOR U43115 ( .A(n43301), .B(n43302), .Z(n780) );
  AND U43116 ( .A(n43303), .B(n43304), .Z(n43302) );
  XNOR U43117 ( .A(p_input[2367]), .B(n43301), .Z(n43304) );
  XOR U43118 ( .A(n43301), .B(p_input[2335]), .Z(n43303) );
  XOR U43119 ( .A(n43305), .B(n43306), .Z(n43301) );
  AND U43120 ( .A(n43307), .B(n43308), .Z(n43306) );
  XNOR U43121 ( .A(p_input[2366]), .B(n43305), .Z(n43308) );
  XNOR U43122 ( .A(n43305), .B(n42907), .Z(n43307) );
  IV U43123 ( .A(p_input[2334]), .Z(n42907) );
  XOR U43124 ( .A(n43309), .B(n43310), .Z(n43305) );
  AND U43125 ( .A(n43311), .B(n43312), .Z(n43310) );
  XNOR U43126 ( .A(p_input[2365]), .B(n43309), .Z(n43312) );
  XNOR U43127 ( .A(n43309), .B(n42916), .Z(n43311) );
  IV U43128 ( .A(p_input[2333]), .Z(n42916) );
  XOR U43129 ( .A(n43313), .B(n43314), .Z(n43309) );
  AND U43130 ( .A(n43315), .B(n43316), .Z(n43314) );
  XNOR U43131 ( .A(p_input[2364]), .B(n43313), .Z(n43316) );
  XNOR U43132 ( .A(n43313), .B(n42925), .Z(n43315) );
  IV U43133 ( .A(p_input[2332]), .Z(n42925) );
  XOR U43134 ( .A(n43317), .B(n43318), .Z(n43313) );
  AND U43135 ( .A(n43319), .B(n43320), .Z(n43318) );
  XNOR U43136 ( .A(p_input[2363]), .B(n43317), .Z(n43320) );
  XNOR U43137 ( .A(n43317), .B(n42934), .Z(n43319) );
  IV U43138 ( .A(p_input[2331]), .Z(n42934) );
  XOR U43139 ( .A(n43321), .B(n43322), .Z(n43317) );
  AND U43140 ( .A(n43323), .B(n43324), .Z(n43322) );
  XNOR U43141 ( .A(p_input[2362]), .B(n43321), .Z(n43324) );
  XNOR U43142 ( .A(n43321), .B(n42943), .Z(n43323) );
  IV U43143 ( .A(p_input[2330]), .Z(n42943) );
  XOR U43144 ( .A(n43325), .B(n43326), .Z(n43321) );
  AND U43145 ( .A(n43327), .B(n43328), .Z(n43326) );
  XNOR U43146 ( .A(p_input[2361]), .B(n43325), .Z(n43328) );
  XNOR U43147 ( .A(n43325), .B(n42952), .Z(n43327) );
  IV U43148 ( .A(p_input[2329]), .Z(n42952) );
  XOR U43149 ( .A(n43329), .B(n43330), .Z(n43325) );
  AND U43150 ( .A(n43331), .B(n43332), .Z(n43330) );
  XNOR U43151 ( .A(p_input[2360]), .B(n43329), .Z(n43332) );
  XNOR U43152 ( .A(n43329), .B(n42961), .Z(n43331) );
  IV U43153 ( .A(p_input[2328]), .Z(n42961) );
  XOR U43154 ( .A(n43333), .B(n43334), .Z(n43329) );
  AND U43155 ( .A(n43335), .B(n43336), .Z(n43334) );
  XNOR U43156 ( .A(p_input[2359]), .B(n43333), .Z(n43336) );
  XNOR U43157 ( .A(n43333), .B(n42970), .Z(n43335) );
  IV U43158 ( .A(p_input[2327]), .Z(n42970) );
  XOR U43159 ( .A(n43337), .B(n43338), .Z(n43333) );
  AND U43160 ( .A(n43339), .B(n43340), .Z(n43338) );
  XNOR U43161 ( .A(p_input[2358]), .B(n43337), .Z(n43340) );
  XNOR U43162 ( .A(n43337), .B(n42979), .Z(n43339) );
  IV U43163 ( .A(p_input[2326]), .Z(n42979) );
  XOR U43164 ( .A(n43341), .B(n43342), .Z(n43337) );
  AND U43165 ( .A(n43343), .B(n43344), .Z(n43342) );
  XNOR U43166 ( .A(p_input[2357]), .B(n43341), .Z(n43344) );
  XNOR U43167 ( .A(n43341), .B(n42988), .Z(n43343) );
  IV U43168 ( .A(p_input[2325]), .Z(n42988) );
  XOR U43169 ( .A(n43345), .B(n43346), .Z(n43341) );
  AND U43170 ( .A(n43347), .B(n43348), .Z(n43346) );
  XNOR U43171 ( .A(p_input[2356]), .B(n43345), .Z(n43348) );
  XNOR U43172 ( .A(n43345), .B(n42997), .Z(n43347) );
  IV U43173 ( .A(p_input[2324]), .Z(n42997) );
  XOR U43174 ( .A(n43349), .B(n43350), .Z(n43345) );
  AND U43175 ( .A(n43351), .B(n43352), .Z(n43350) );
  XNOR U43176 ( .A(p_input[2355]), .B(n43349), .Z(n43352) );
  XNOR U43177 ( .A(n43349), .B(n43006), .Z(n43351) );
  IV U43178 ( .A(p_input[2323]), .Z(n43006) );
  XOR U43179 ( .A(n43353), .B(n43354), .Z(n43349) );
  AND U43180 ( .A(n43355), .B(n43356), .Z(n43354) );
  XNOR U43181 ( .A(p_input[2354]), .B(n43353), .Z(n43356) );
  XNOR U43182 ( .A(n43353), .B(n43015), .Z(n43355) );
  IV U43183 ( .A(p_input[2322]), .Z(n43015) );
  XOR U43184 ( .A(n43357), .B(n43358), .Z(n43353) );
  AND U43185 ( .A(n43359), .B(n43360), .Z(n43358) );
  XNOR U43186 ( .A(p_input[2353]), .B(n43357), .Z(n43360) );
  XNOR U43187 ( .A(n43357), .B(n43024), .Z(n43359) );
  IV U43188 ( .A(p_input[2321]), .Z(n43024) );
  XOR U43189 ( .A(n43361), .B(n43362), .Z(n43357) );
  AND U43190 ( .A(n43363), .B(n43364), .Z(n43362) );
  XNOR U43191 ( .A(p_input[2352]), .B(n43361), .Z(n43364) );
  XNOR U43192 ( .A(n43361), .B(n43033), .Z(n43363) );
  IV U43193 ( .A(p_input[2320]), .Z(n43033) );
  XOR U43194 ( .A(n43365), .B(n43366), .Z(n43361) );
  AND U43195 ( .A(n43367), .B(n43368), .Z(n43366) );
  XNOR U43196 ( .A(p_input[2351]), .B(n43365), .Z(n43368) );
  XNOR U43197 ( .A(n43365), .B(n43042), .Z(n43367) );
  IV U43198 ( .A(p_input[2319]), .Z(n43042) );
  XOR U43199 ( .A(n43369), .B(n43370), .Z(n43365) );
  AND U43200 ( .A(n43371), .B(n43372), .Z(n43370) );
  XNOR U43201 ( .A(p_input[2350]), .B(n43369), .Z(n43372) );
  XNOR U43202 ( .A(n43369), .B(n43051), .Z(n43371) );
  IV U43203 ( .A(p_input[2318]), .Z(n43051) );
  XOR U43204 ( .A(n43373), .B(n43374), .Z(n43369) );
  AND U43205 ( .A(n43375), .B(n43376), .Z(n43374) );
  XNOR U43206 ( .A(p_input[2349]), .B(n43373), .Z(n43376) );
  XNOR U43207 ( .A(n43373), .B(n43060), .Z(n43375) );
  IV U43208 ( .A(p_input[2317]), .Z(n43060) );
  XOR U43209 ( .A(n43377), .B(n43378), .Z(n43373) );
  AND U43210 ( .A(n43379), .B(n43380), .Z(n43378) );
  XNOR U43211 ( .A(p_input[2348]), .B(n43377), .Z(n43380) );
  XNOR U43212 ( .A(n43377), .B(n43069), .Z(n43379) );
  IV U43213 ( .A(p_input[2316]), .Z(n43069) );
  XOR U43214 ( .A(n43381), .B(n43382), .Z(n43377) );
  AND U43215 ( .A(n43383), .B(n43384), .Z(n43382) );
  XNOR U43216 ( .A(p_input[2347]), .B(n43381), .Z(n43384) );
  XNOR U43217 ( .A(n43381), .B(n43078), .Z(n43383) );
  IV U43218 ( .A(p_input[2315]), .Z(n43078) );
  XOR U43219 ( .A(n43385), .B(n43386), .Z(n43381) );
  AND U43220 ( .A(n43387), .B(n43388), .Z(n43386) );
  XNOR U43221 ( .A(p_input[2346]), .B(n43385), .Z(n43388) );
  XNOR U43222 ( .A(n43385), .B(n43087), .Z(n43387) );
  IV U43223 ( .A(p_input[2314]), .Z(n43087) );
  XOR U43224 ( .A(n43389), .B(n43390), .Z(n43385) );
  AND U43225 ( .A(n43391), .B(n43392), .Z(n43390) );
  XNOR U43226 ( .A(p_input[2345]), .B(n43389), .Z(n43392) );
  XNOR U43227 ( .A(n43389), .B(n43096), .Z(n43391) );
  IV U43228 ( .A(p_input[2313]), .Z(n43096) );
  XOR U43229 ( .A(n43393), .B(n43394), .Z(n43389) );
  AND U43230 ( .A(n43395), .B(n43396), .Z(n43394) );
  XNOR U43231 ( .A(p_input[2344]), .B(n43393), .Z(n43396) );
  XNOR U43232 ( .A(n43393), .B(n43105), .Z(n43395) );
  IV U43233 ( .A(p_input[2312]), .Z(n43105) );
  XOR U43234 ( .A(n43397), .B(n43398), .Z(n43393) );
  AND U43235 ( .A(n43399), .B(n43400), .Z(n43398) );
  XNOR U43236 ( .A(p_input[2343]), .B(n43397), .Z(n43400) );
  XNOR U43237 ( .A(n43397), .B(n43114), .Z(n43399) );
  IV U43238 ( .A(p_input[2311]), .Z(n43114) );
  XOR U43239 ( .A(n43401), .B(n43402), .Z(n43397) );
  AND U43240 ( .A(n43403), .B(n43404), .Z(n43402) );
  XNOR U43241 ( .A(p_input[2342]), .B(n43401), .Z(n43404) );
  XNOR U43242 ( .A(n43401), .B(n43123), .Z(n43403) );
  IV U43243 ( .A(p_input[2310]), .Z(n43123) );
  XOR U43244 ( .A(n43405), .B(n43406), .Z(n43401) );
  AND U43245 ( .A(n43407), .B(n43408), .Z(n43406) );
  XNOR U43246 ( .A(p_input[2341]), .B(n43405), .Z(n43408) );
  XNOR U43247 ( .A(n43405), .B(n43132), .Z(n43407) );
  IV U43248 ( .A(p_input[2309]), .Z(n43132) );
  XOR U43249 ( .A(n43409), .B(n43410), .Z(n43405) );
  AND U43250 ( .A(n43411), .B(n43412), .Z(n43410) );
  XNOR U43251 ( .A(p_input[2340]), .B(n43409), .Z(n43412) );
  XNOR U43252 ( .A(n43409), .B(n43141), .Z(n43411) );
  IV U43253 ( .A(p_input[2308]), .Z(n43141) );
  XOR U43254 ( .A(n43413), .B(n43414), .Z(n43409) );
  AND U43255 ( .A(n43415), .B(n43416), .Z(n43414) );
  XNOR U43256 ( .A(p_input[2339]), .B(n43413), .Z(n43416) );
  XNOR U43257 ( .A(n43413), .B(n43150), .Z(n43415) );
  IV U43258 ( .A(p_input[2307]), .Z(n43150) );
  XOR U43259 ( .A(n43417), .B(n43418), .Z(n43413) );
  AND U43260 ( .A(n43419), .B(n43420), .Z(n43418) );
  XNOR U43261 ( .A(p_input[2338]), .B(n43417), .Z(n43420) );
  XNOR U43262 ( .A(n43417), .B(n43159), .Z(n43419) );
  IV U43263 ( .A(p_input[2306]), .Z(n43159) );
  XNOR U43264 ( .A(n43421), .B(n43422), .Z(n43417) );
  AND U43265 ( .A(n43423), .B(n43424), .Z(n43422) );
  XOR U43266 ( .A(p_input[2337]), .B(n43421), .Z(n43424) );
  XNOR U43267 ( .A(p_input[2305]), .B(n43421), .Z(n43423) );
  AND U43268 ( .A(p_input[2336]), .B(n43425), .Z(n43421) );
  IV U43269 ( .A(p_input[2304]), .Z(n43425) );
  XOR U43270 ( .A(n43426), .B(n43427), .Z(n41604) );
  AND U43271 ( .A(n888), .B(n43428), .Z(n43427) );
  XNOR U43272 ( .A(n43429), .B(n43426), .Z(n43428) );
  XOR U43273 ( .A(n43430), .B(n43431), .Z(n888) );
  AND U43274 ( .A(n43432), .B(n43433), .Z(n43431) );
  XOR U43275 ( .A(n43430), .B(n41619), .Z(n43433) );
  XNOR U43276 ( .A(n43434), .B(n43435), .Z(n41619) );
  AND U43277 ( .A(n43436), .B(n607), .Z(n43435) );
  AND U43278 ( .A(n43434), .B(n43437), .Z(n43436) );
  XNOR U43279 ( .A(n41616), .B(n43430), .Z(n43432) );
  XOR U43280 ( .A(n43438), .B(n43439), .Z(n41616) );
  AND U43281 ( .A(n43440), .B(n604), .Z(n43439) );
  NOR U43282 ( .A(n43438), .B(n43441), .Z(n43440) );
  XOR U43283 ( .A(n43442), .B(n43443), .Z(n43430) );
  AND U43284 ( .A(n43444), .B(n43445), .Z(n43443) );
  XOR U43285 ( .A(n43442), .B(n41631), .Z(n43445) );
  XOR U43286 ( .A(n43446), .B(n43447), .Z(n41631) );
  AND U43287 ( .A(n607), .B(n43448), .Z(n43447) );
  XOR U43288 ( .A(n43449), .B(n43446), .Z(n43448) );
  XNOR U43289 ( .A(n41628), .B(n43442), .Z(n43444) );
  XOR U43290 ( .A(n43450), .B(n43451), .Z(n41628) );
  AND U43291 ( .A(n604), .B(n43452), .Z(n43451) );
  XOR U43292 ( .A(n43453), .B(n43450), .Z(n43452) );
  XOR U43293 ( .A(n43454), .B(n43455), .Z(n43442) );
  AND U43294 ( .A(n43456), .B(n43457), .Z(n43455) );
  XOR U43295 ( .A(n43454), .B(n41643), .Z(n43457) );
  XOR U43296 ( .A(n43458), .B(n43459), .Z(n41643) );
  AND U43297 ( .A(n607), .B(n43460), .Z(n43459) );
  XOR U43298 ( .A(n43461), .B(n43458), .Z(n43460) );
  XNOR U43299 ( .A(n41640), .B(n43454), .Z(n43456) );
  XOR U43300 ( .A(n43462), .B(n43463), .Z(n41640) );
  AND U43301 ( .A(n604), .B(n43464), .Z(n43463) );
  XOR U43302 ( .A(n43465), .B(n43462), .Z(n43464) );
  XOR U43303 ( .A(n43466), .B(n43467), .Z(n43454) );
  AND U43304 ( .A(n43468), .B(n43469), .Z(n43467) );
  XOR U43305 ( .A(n43466), .B(n41655), .Z(n43469) );
  XOR U43306 ( .A(n43470), .B(n43471), .Z(n41655) );
  AND U43307 ( .A(n607), .B(n43472), .Z(n43471) );
  XOR U43308 ( .A(n43473), .B(n43470), .Z(n43472) );
  XNOR U43309 ( .A(n41652), .B(n43466), .Z(n43468) );
  XOR U43310 ( .A(n43474), .B(n43475), .Z(n41652) );
  AND U43311 ( .A(n604), .B(n43476), .Z(n43475) );
  XOR U43312 ( .A(n43477), .B(n43474), .Z(n43476) );
  XOR U43313 ( .A(n43478), .B(n43479), .Z(n43466) );
  AND U43314 ( .A(n43480), .B(n43481), .Z(n43479) );
  XOR U43315 ( .A(n43478), .B(n41667), .Z(n43481) );
  XOR U43316 ( .A(n43482), .B(n43483), .Z(n41667) );
  AND U43317 ( .A(n607), .B(n43484), .Z(n43483) );
  XOR U43318 ( .A(n43485), .B(n43482), .Z(n43484) );
  XNOR U43319 ( .A(n41664), .B(n43478), .Z(n43480) );
  XOR U43320 ( .A(n43486), .B(n43487), .Z(n41664) );
  AND U43321 ( .A(n604), .B(n43488), .Z(n43487) );
  XOR U43322 ( .A(n43489), .B(n43486), .Z(n43488) );
  XOR U43323 ( .A(n43490), .B(n43491), .Z(n43478) );
  AND U43324 ( .A(n43492), .B(n43493), .Z(n43491) );
  XOR U43325 ( .A(n43490), .B(n41679), .Z(n43493) );
  XOR U43326 ( .A(n43494), .B(n43495), .Z(n41679) );
  AND U43327 ( .A(n607), .B(n43496), .Z(n43495) );
  XOR U43328 ( .A(n43497), .B(n43494), .Z(n43496) );
  XNOR U43329 ( .A(n41676), .B(n43490), .Z(n43492) );
  XOR U43330 ( .A(n43498), .B(n43499), .Z(n41676) );
  AND U43331 ( .A(n604), .B(n43500), .Z(n43499) );
  XOR U43332 ( .A(n43501), .B(n43498), .Z(n43500) );
  XOR U43333 ( .A(n43502), .B(n43503), .Z(n43490) );
  AND U43334 ( .A(n43504), .B(n43505), .Z(n43503) );
  XOR U43335 ( .A(n43502), .B(n41691), .Z(n43505) );
  XOR U43336 ( .A(n43506), .B(n43507), .Z(n41691) );
  AND U43337 ( .A(n607), .B(n43508), .Z(n43507) );
  XOR U43338 ( .A(n43509), .B(n43506), .Z(n43508) );
  XNOR U43339 ( .A(n41688), .B(n43502), .Z(n43504) );
  XOR U43340 ( .A(n43510), .B(n43511), .Z(n41688) );
  AND U43341 ( .A(n604), .B(n43512), .Z(n43511) );
  XOR U43342 ( .A(n43513), .B(n43510), .Z(n43512) );
  XOR U43343 ( .A(n43514), .B(n43515), .Z(n43502) );
  AND U43344 ( .A(n43516), .B(n43517), .Z(n43515) );
  XOR U43345 ( .A(n43514), .B(n41703), .Z(n43517) );
  XOR U43346 ( .A(n43518), .B(n43519), .Z(n41703) );
  AND U43347 ( .A(n607), .B(n43520), .Z(n43519) );
  XOR U43348 ( .A(n43521), .B(n43518), .Z(n43520) );
  XNOR U43349 ( .A(n41700), .B(n43514), .Z(n43516) );
  XOR U43350 ( .A(n43522), .B(n43523), .Z(n41700) );
  AND U43351 ( .A(n604), .B(n43524), .Z(n43523) );
  XOR U43352 ( .A(n43525), .B(n43522), .Z(n43524) );
  XOR U43353 ( .A(n43526), .B(n43527), .Z(n43514) );
  AND U43354 ( .A(n43528), .B(n43529), .Z(n43527) );
  XOR U43355 ( .A(n43526), .B(n41715), .Z(n43529) );
  XOR U43356 ( .A(n43530), .B(n43531), .Z(n41715) );
  AND U43357 ( .A(n607), .B(n43532), .Z(n43531) );
  XOR U43358 ( .A(n43533), .B(n43530), .Z(n43532) );
  XNOR U43359 ( .A(n41712), .B(n43526), .Z(n43528) );
  XOR U43360 ( .A(n43534), .B(n43535), .Z(n41712) );
  AND U43361 ( .A(n604), .B(n43536), .Z(n43535) );
  XOR U43362 ( .A(n43537), .B(n43534), .Z(n43536) );
  XOR U43363 ( .A(n43538), .B(n43539), .Z(n43526) );
  AND U43364 ( .A(n43540), .B(n43541), .Z(n43539) );
  XOR U43365 ( .A(n43538), .B(n41727), .Z(n43541) );
  XOR U43366 ( .A(n43542), .B(n43543), .Z(n41727) );
  AND U43367 ( .A(n607), .B(n43544), .Z(n43543) );
  XOR U43368 ( .A(n43545), .B(n43542), .Z(n43544) );
  XNOR U43369 ( .A(n41724), .B(n43538), .Z(n43540) );
  XOR U43370 ( .A(n43546), .B(n43547), .Z(n41724) );
  AND U43371 ( .A(n604), .B(n43548), .Z(n43547) );
  XOR U43372 ( .A(n43549), .B(n43546), .Z(n43548) );
  XOR U43373 ( .A(n43550), .B(n43551), .Z(n43538) );
  AND U43374 ( .A(n43552), .B(n43553), .Z(n43551) );
  XOR U43375 ( .A(n43550), .B(n41739), .Z(n43553) );
  XOR U43376 ( .A(n43554), .B(n43555), .Z(n41739) );
  AND U43377 ( .A(n607), .B(n43556), .Z(n43555) );
  XOR U43378 ( .A(n43557), .B(n43554), .Z(n43556) );
  XNOR U43379 ( .A(n41736), .B(n43550), .Z(n43552) );
  XOR U43380 ( .A(n43558), .B(n43559), .Z(n41736) );
  AND U43381 ( .A(n604), .B(n43560), .Z(n43559) );
  XOR U43382 ( .A(n43561), .B(n43558), .Z(n43560) );
  XOR U43383 ( .A(n43562), .B(n43563), .Z(n43550) );
  AND U43384 ( .A(n43564), .B(n43565), .Z(n43563) );
  XOR U43385 ( .A(n43562), .B(n41751), .Z(n43565) );
  XOR U43386 ( .A(n43566), .B(n43567), .Z(n41751) );
  AND U43387 ( .A(n607), .B(n43568), .Z(n43567) );
  XOR U43388 ( .A(n43569), .B(n43566), .Z(n43568) );
  XNOR U43389 ( .A(n41748), .B(n43562), .Z(n43564) );
  XOR U43390 ( .A(n43570), .B(n43571), .Z(n41748) );
  AND U43391 ( .A(n604), .B(n43572), .Z(n43571) );
  XOR U43392 ( .A(n43573), .B(n43570), .Z(n43572) );
  XOR U43393 ( .A(n43574), .B(n43575), .Z(n43562) );
  AND U43394 ( .A(n43576), .B(n43577), .Z(n43575) );
  XOR U43395 ( .A(n43574), .B(n41763), .Z(n43577) );
  XOR U43396 ( .A(n43578), .B(n43579), .Z(n41763) );
  AND U43397 ( .A(n607), .B(n43580), .Z(n43579) );
  XOR U43398 ( .A(n43581), .B(n43578), .Z(n43580) );
  XNOR U43399 ( .A(n41760), .B(n43574), .Z(n43576) );
  XOR U43400 ( .A(n43582), .B(n43583), .Z(n41760) );
  AND U43401 ( .A(n604), .B(n43584), .Z(n43583) );
  XOR U43402 ( .A(n43585), .B(n43582), .Z(n43584) );
  XOR U43403 ( .A(n43586), .B(n43587), .Z(n43574) );
  AND U43404 ( .A(n43588), .B(n43589), .Z(n43587) );
  XOR U43405 ( .A(n43586), .B(n41775), .Z(n43589) );
  XOR U43406 ( .A(n43590), .B(n43591), .Z(n41775) );
  AND U43407 ( .A(n607), .B(n43592), .Z(n43591) );
  XOR U43408 ( .A(n43593), .B(n43590), .Z(n43592) );
  XNOR U43409 ( .A(n41772), .B(n43586), .Z(n43588) );
  XOR U43410 ( .A(n43594), .B(n43595), .Z(n41772) );
  AND U43411 ( .A(n604), .B(n43596), .Z(n43595) );
  XOR U43412 ( .A(n43597), .B(n43594), .Z(n43596) );
  XOR U43413 ( .A(n43598), .B(n43599), .Z(n43586) );
  AND U43414 ( .A(n43600), .B(n43601), .Z(n43599) );
  XOR U43415 ( .A(n43598), .B(n41787), .Z(n43601) );
  XOR U43416 ( .A(n43602), .B(n43603), .Z(n41787) );
  AND U43417 ( .A(n607), .B(n43604), .Z(n43603) );
  XOR U43418 ( .A(n43605), .B(n43602), .Z(n43604) );
  XNOR U43419 ( .A(n41784), .B(n43598), .Z(n43600) );
  XOR U43420 ( .A(n43606), .B(n43607), .Z(n41784) );
  AND U43421 ( .A(n604), .B(n43608), .Z(n43607) );
  XOR U43422 ( .A(n43609), .B(n43606), .Z(n43608) );
  XOR U43423 ( .A(n43610), .B(n43611), .Z(n43598) );
  AND U43424 ( .A(n43612), .B(n43613), .Z(n43611) );
  XOR U43425 ( .A(n43610), .B(n41799), .Z(n43613) );
  XOR U43426 ( .A(n43614), .B(n43615), .Z(n41799) );
  AND U43427 ( .A(n607), .B(n43616), .Z(n43615) );
  XOR U43428 ( .A(n43617), .B(n43614), .Z(n43616) );
  XNOR U43429 ( .A(n41796), .B(n43610), .Z(n43612) );
  XOR U43430 ( .A(n43618), .B(n43619), .Z(n41796) );
  AND U43431 ( .A(n604), .B(n43620), .Z(n43619) );
  XOR U43432 ( .A(n43621), .B(n43618), .Z(n43620) );
  XOR U43433 ( .A(n43622), .B(n43623), .Z(n43610) );
  AND U43434 ( .A(n43624), .B(n43625), .Z(n43623) );
  XOR U43435 ( .A(n43622), .B(n41811), .Z(n43625) );
  XOR U43436 ( .A(n43626), .B(n43627), .Z(n41811) );
  AND U43437 ( .A(n607), .B(n43628), .Z(n43627) );
  XOR U43438 ( .A(n43629), .B(n43626), .Z(n43628) );
  XNOR U43439 ( .A(n41808), .B(n43622), .Z(n43624) );
  XOR U43440 ( .A(n43630), .B(n43631), .Z(n41808) );
  AND U43441 ( .A(n604), .B(n43632), .Z(n43631) );
  XOR U43442 ( .A(n43633), .B(n43630), .Z(n43632) );
  XOR U43443 ( .A(n43634), .B(n43635), .Z(n43622) );
  AND U43444 ( .A(n43636), .B(n43637), .Z(n43635) );
  XOR U43445 ( .A(n43634), .B(n41823), .Z(n43637) );
  XOR U43446 ( .A(n43638), .B(n43639), .Z(n41823) );
  AND U43447 ( .A(n607), .B(n43640), .Z(n43639) );
  XOR U43448 ( .A(n43641), .B(n43638), .Z(n43640) );
  XNOR U43449 ( .A(n41820), .B(n43634), .Z(n43636) );
  XOR U43450 ( .A(n43642), .B(n43643), .Z(n41820) );
  AND U43451 ( .A(n604), .B(n43644), .Z(n43643) );
  XOR U43452 ( .A(n43645), .B(n43642), .Z(n43644) );
  XOR U43453 ( .A(n43646), .B(n43647), .Z(n43634) );
  AND U43454 ( .A(n43648), .B(n43649), .Z(n43647) );
  XOR U43455 ( .A(n43646), .B(n41835), .Z(n43649) );
  XOR U43456 ( .A(n43650), .B(n43651), .Z(n41835) );
  AND U43457 ( .A(n607), .B(n43652), .Z(n43651) );
  XOR U43458 ( .A(n43653), .B(n43650), .Z(n43652) );
  XNOR U43459 ( .A(n41832), .B(n43646), .Z(n43648) );
  XOR U43460 ( .A(n43654), .B(n43655), .Z(n41832) );
  AND U43461 ( .A(n604), .B(n43656), .Z(n43655) );
  XOR U43462 ( .A(n43657), .B(n43654), .Z(n43656) );
  XOR U43463 ( .A(n43658), .B(n43659), .Z(n43646) );
  AND U43464 ( .A(n43660), .B(n43661), .Z(n43659) );
  XOR U43465 ( .A(n43658), .B(n41847), .Z(n43661) );
  XOR U43466 ( .A(n43662), .B(n43663), .Z(n41847) );
  AND U43467 ( .A(n607), .B(n43664), .Z(n43663) );
  XOR U43468 ( .A(n43665), .B(n43662), .Z(n43664) );
  XNOR U43469 ( .A(n41844), .B(n43658), .Z(n43660) );
  XOR U43470 ( .A(n43666), .B(n43667), .Z(n41844) );
  AND U43471 ( .A(n604), .B(n43668), .Z(n43667) );
  XOR U43472 ( .A(n43669), .B(n43666), .Z(n43668) );
  XOR U43473 ( .A(n43670), .B(n43671), .Z(n43658) );
  AND U43474 ( .A(n43672), .B(n43673), .Z(n43671) );
  XOR U43475 ( .A(n43670), .B(n41859), .Z(n43673) );
  XOR U43476 ( .A(n43674), .B(n43675), .Z(n41859) );
  AND U43477 ( .A(n607), .B(n43676), .Z(n43675) );
  XOR U43478 ( .A(n43677), .B(n43674), .Z(n43676) );
  XNOR U43479 ( .A(n41856), .B(n43670), .Z(n43672) );
  XOR U43480 ( .A(n43678), .B(n43679), .Z(n41856) );
  AND U43481 ( .A(n604), .B(n43680), .Z(n43679) );
  XOR U43482 ( .A(n43681), .B(n43678), .Z(n43680) );
  XOR U43483 ( .A(n43682), .B(n43683), .Z(n43670) );
  AND U43484 ( .A(n43684), .B(n43685), .Z(n43683) );
  XOR U43485 ( .A(n43682), .B(n41871), .Z(n43685) );
  XOR U43486 ( .A(n43686), .B(n43687), .Z(n41871) );
  AND U43487 ( .A(n607), .B(n43688), .Z(n43687) );
  XOR U43488 ( .A(n43689), .B(n43686), .Z(n43688) );
  XNOR U43489 ( .A(n41868), .B(n43682), .Z(n43684) );
  XOR U43490 ( .A(n43690), .B(n43691), .Z(n41868) );
  AND U43491 ( .A(n604), .B(n43692), .Z(n43691) );
  XOR U43492 ( .A(n43693), .B(n43690), .Z(n43692) );
  XOR U43493 ( .A(n43694), .B(n43695), .Z(n43682) );
  AND U43494 ( .A(n43696), .B(n43697), .Z(n43695) );
  XOR U43495 ( .A(n43694), .B(n41883), .Z(n43697) );
  XOR U43496 ( .A(n43698), .B(n43699), .Z(n41883) );
  AND U43497 ( .A(n607), .B(n43700), .Z(n43699) );
  XOR U43498 ( .A(n43701), .B(n43698), .Z(n43700) );
  XNOR U43499 ( .A(n41880), .B(n43694), .Z(n43696) );
  XOR U43500 ( .A(n43702), .B(n43703), .Z(n41880) );
  AND U43501 ( .A(n604), .B(n43704), .Z(n43703) );
  XOR U43502 ( .A(n43705), .B(n43702), .Z(n43704) );
  XOR U43503 ( .A(n43706), .B(n43707), .Z(n43694) );
  AND U43504 ( .A(n43708), .B(n43709), .Z(n43707) );
  XOR U43505 ( .A(n43706), .B(n41895), .Z(n43709) );
  XOR U43506 ( .A(n43710), .B(n43711), .Z(n41895) );
  AND U43507 ( .A(n607), .B(n43712), .Z(n43711) );
  XOR U43508 ( .A(n43713), .B(n43710), .Z(n43712) );
  XNOR U43509 ( .A(n41892), .B(n43706), .Z(n43708) );
  XOR U43510 ( .A(n43714), .B(n43715), .Z(n41892) );
  AND U43511 ( .A(n604), .B(n43716), .Z(n43715) );
  XOR U43512 ( .A(n43717), .B(n43714), .Z(n43716) );
  XOR U43513 ( .A(n43718), .B(n43719), .Z(n43706) );
  AND U43514 ( .A(n43720), .B(n43721), .Z(n43719) );
  XOR U43515 ( .A(n43718), .B(n41907), .Z(n43721) );
  XOR U43516 ( .A(n43722), .B(n43723), .Z(n41907) );
  AND U43517 ( .A(n607), .B(n43724), .Z(n43723) );
  XOR U43518 ( .A(n43725), .B(n43722), .Z(n43724) );
  XNOR U43519 ( .A(n41904), .B(n43718), .Z(n43720) );
  XOR U43520 ( .A(n43726), .B(n43727), .Z(n41904) );
  AND U43521 ( .A(n604), .B(n43728), .Z(n43727) );
  XOR U43522 ( .A(n43729), .B(n43726), .Z(n43728) );
  XOR U43523 ( .A(n43730), .B(n43731), .Z(n43718) );
  AND U43524 ( .A(n43732), .B(n43733), .Z(n43731) );
  XOR U43525 ( .A(n43730), .B(n41919), .Z(n43733) );
  XOR U43526 ( .A(n43734), .B(n43735), .Z(n41919) );
  AND U43527 ( .A(n607), .B(n43736), .Z(n43735) );
  XOR U43528 ( .A(n43737), .B(n43734), .Z(n43736) );
  XNOR U43529 ( .A(n41916), .B(n43730), .Z(n43732) );
  XOR U43530 ( .A(n43738), .B(n43739), .Z(n41916) );
  AND U43531 ( .A(n604), .B(n43740), .Z(n43739) );
  XOR U43532 ( .A(n43741), .B(n43738), .Z(n43740) );
  XOR U43533 ( .A(n43742), .B(n43743), .Z(n43730) );
  AND U43534 ( .A(n43744), .B(n43745), .Z(n43743) );
  XOR U43535 ( .A(n43742), .B(n41931), .Z(n43745) );
  XOR U43536 ( .A(n43746), .B(n43747), .Z(n41931) );
  AND U43537 ( .A(n607), .B(n43748), .Z(n43747) );
  XOR U43538 ( .A(n43749), .B(n43746), .Z(n43748) );
  XNOR U43539 ( .A(n41928), .B(n43742), .Z(n43744) );
  XOR U43540 ( .A(n43750), .B(n43751), .Z(n41928) );
  AND U43541 ( .A(n604), .B(n43752), .Z(n43751) );
  XOR U43542 ( .A(n43753), .B(n43750), .Z(n43752) );
  XOR U43543 ( .A(n43754), .B(n43755), .Z(n43742) );
  AND U43544 ( .A(n43756), .B(n43757), .Z(n43755) );
  XOR U43545 ( .A(n43754), .B(n41943), .Z(n43757) );
  XOR U43546 ( .A(n43758), .B(n43759), .Z(n41943) );
  AND U43547 ( .A(n607), .B(n43760), .Z(n43759) );
  XOR U43548 ( .A(n43761), .B(n43758), .Z(n43760) );
  XNOR U43549 ( .A(n41940), .B(n43754), .Z(n43756) );
  XOR U43550 ( .A(n43762), .B(n43763), .Z(n41940) );
  AND U43551 ( .A(n604), .B(n43764), .Z(n43763) );
  XOR U43552 ( .A(n43765), .B(n43762), .Z(n43764) );
  XOR U43553 ( .A(n43766), .B(n43767), .Z(n43754) );
  AND U43554 ( .A(n43768), .B(n43769), .Z(n43767) );
  XOR U43555 ( .A(n43766), .B(n41955), .Z(n43769) );
  XOR U43556 ( .A(n43770), .B(n43771), .Z(n41955) );
  AND U43557 ( .A(n607), .B(n43772), .Z(n43771) );
  XOR U43558 ( .A(n43773), .B(n43770), .Z(n43772) );
  XNOR U43559 ( .A(n41952), .B(n43766), .Z(n43768) );
  XOR U43560 ( .A(n43774), .B(n43775), .Z(n41952) );
  AND U43561 ( .A(n604), .B(n43776), .Z(n43775) );
  XOR U43562 ( .A(n43777), .B(n43774), .Z(n43776) );
  XOR U43563 ( .A(n43778), .B(n43779), .Z(n43766) );
  AND U43564 ( .A(n43780), .B(n43781), .Z(n43779) );
  XOR U43565 ( .A(n43778), .B(n41967), .Z(n43781) );
  XOR U43566 ( .A(n43782), .B(n43783), .Z(n41967) );
  AND U43567 ( .A(n607), .B(n43784), .Z(n43783) );
  XOR U43568 ( .A(n43785), .B(n43782), .Z(n43784) );
  XNOR U43569 ( .A(n41964), .B(n43778), .Z(n43780) );
  XOR U43570 ( .A(n43786), .B(n43787), .Z(n41964) );
  AND U43571 ( .A(n604), .B(n43788), .Z(n43787) );
  XOR U43572 ( .A(n43789), .B(n43786), .Z(n43788) );
  XOR U43573 ( .A(n43790), .B(n43791), .Z(n43778) );
  AND U43574 ( .A(n43792), .B(n43793), .Z(n43791) );
  XNOR U43575 ( .A(n43794), .B(n41980), .Z(n43793) );
  XOR U43576 ( .A(n43795), .B(n43796), .Z(n41980) );
  AND U43577 ( .A(n607), .B(n43797), .Z(n43796) );
  XOR U43578 ( .A(n43795), .B(n43798), .Z(n43797) );
  XNOR U43579 ( .A(n41977), .B(n43790), .Z(n43792) );
  XOR U43580 ( .A(n43799), .B(n43800), .Z(n41977) );
  AND U43581 ( .A(n604), .B(n43801), .Z(n43800) );
  XOR U43582 ( .A(n43799), .B(n43802), .Z(n43801) );
  IV U43583 ( .A(n43794), .Z(n43790) );
  AND U43584 ( .A(n43426), .B(n43429), .Z(n43794) );
  XNOR U43585 ( .A(n43803), .B(n43804), .Z(n43429) );
  AND U43586 ( .A(n607), .B(n43805), .Z(n43804) );
  XNOR U43587 ( .A(n43806), .B(n43803), .Z(n43805) );
  XOR U43588 ( .A(n43807), .B(n43808), .Z(n607) );
  AND U43589 ( .A(n43809), .B(n43810), .Z(n43808) );
  XOR U43590 ( .A(n43437), .B(n43807), .Z(n43810) );
  IV U43591 ( .A(n43811), .Z(n43437) );
  AND U43592 ( .A(p_input[2303]), .B(p_input[2271]), .Z(n43811) );
  XOR U43593 ( .A(n43807), .B(n43434), .Z(n43809) );
  AND U43594 ( .A(p_input[2207]), .B(p_input[2239]), .Z(n43434) );
  XOR U43595 ( .A(n43812), .B(n43813), .Z(n43807) );
  AND U43596 ( .A(n43814), .B(n43815), .Z(n43813) );
  XOR U43597 ( .A(n43812), .B(n43449), .Z(n43815) );
  XNOR U43598 ( .A(p_input[2270]), .B(n43816), .Z(n43449) );
  AND U43599 ( .A(n791), .B(n43817), .Z(n43816) );
  XOR U43600 ( .A(p_input[2302]), .B(p_input[2270]), .Z(n43817) );
  XNOR U43601 ( .A(n43446), .B(n43812), .Z(n43814) );
  XOR U43602 ( .A(n43818), .B(n43819), .Z(n43446) );
  AND U43603 ( .A(n789), .B(n43820), .Z(n43819) );
  XOR U43604 ( .A(p_input[2238]), .B(p_input[2206]), .Z(n43820) );
  XOR U43605 ( .A(n43821), .B(n43822), .Z(n43812) );
  AND U43606 ( .A(n43823), .B(n43824), .Z(n43822) );
  XOR U43607 ( .A(n43821), .B(n43461), .Z(n43824) );
  XNOR U43608 ( .A(p_input[2269]), .B(n43825), .Z(n43461) );
  AND U43609 ( .A(n791), .B(n43826), .Z(n43825) );
  XOR U43610 ( .A(p_input[2301]), .B(p_input[2269]), .Z(n43826) );
  XNOR U43611 ( .A(n43458), .B(n43821), .Z(n43823) );
  XOR U43612 ( .A(n43827), .B(n43828), .Z(n43458) );
  AND U43613 ( .A(n789), .B(n43829), .Z(n43828) );
  XOR U43614 ( .A(p_input[2237]), .B(p_input[2205]), .Z(n43829) );
  XOR U43615 ( .A(n43830), .B(n43831), .Z(n43821) );
  AND U43616 ( .A(n43832), .B(n43833), .Z(n43831) );
  XOR U43617 ( .A(n43830), .B(n43473), .Z(n43833) );
  XNOR U43618 ( .A(p_input[2268]), .B(n43834), .Z(n43473) );
  AND U43619 ( .A(n791), .B(n43835), .Z(n43834) );
  XOR U43620 ( .A(p_input[2300]), .B(p_input[2268]), .Z(n43835) );
  XNOR U43621 ( .A(n43470), .B(n43830), .Z(n43832) );
  XOR U43622 ( .A(n43836), .B(n43837), .Z(n43470) );
  AND U43623 ( .A(n789), .B(n43838), .Z(n43837) );
  XOR U43624 ( .A(p_input[2236]), .B(p_input[2204]), .Z(n43838) );
  XOR U43625 ( .A(n43839), .B(n43840), .Z(n43830) );
  AND U43626 ( .A(n43841), .B(n43842), .Z(n43840) );
  XOR U43627 ( .A(n43839), .B(n43485), .Z(n43842) );
  XNOR U43628 ( .A(p_input[2267]), .B(n43843), .Z(n43485) );
  AND U43629 ( .A(n791), .B(n43844), .Z(n43843) );
  XOR U43630 ( .A(p_input[2299]), .B(p_input[2267]), .Z(n43844) );
  XNOR U43631 ( .A(n43482), .B(n43839), .Z(n43841) );
  XOR U43632 ( .A(n43845), .B(n43846), .Z(n43482) );
  AND U43633 ( .A(n789), .B(n43847), .Z(n43846) );
  XOR U43634 ( .A(p_input[2235]), .B(p_input[2203]), .Z(n43847) );
  XOR U43635 ( .A(n43848), .B(n43849), .Z(n43839) );
  AND U43636 ( .A(n43850), .B(n43851), .Z(n43849) );
  XOR U43637 ( .A(n43848), .B(n43497), .Z(n43851) );
  XNOR U43638 ( .A(p_input[2266]), .B(n43852), .Z(n43497) );
  AND U43639 ( .A(n791), .B(n43853), .Z(n43852) );
  XOR U43640 ( .A(p_input[2298]), .B(p_input[2266]), .Z(n43853) );
  XNOR U43641 ( .A(n43494), .B(n43848), .Z(n43850) );
  XOR U43642 ( .A(n43854), .B(n43855), .Z(n43494) );
  AND U43643 ( .A(n789), .B(n43856), .Z(n43855) );
  XOR U43644 ( .A(p_input[2234]), .B(p_input[2202]), .Z(n43856) );
  XOR U43645 ( .A(n43857), .B(n43858), .Z(n43848) );
  AND U43646 ( .A(n43859), .B(n43860), .Z(n43858) );
  XOR U43647 ( .A(n43857), .B(n43509), .Z(n43860) );
  XNOR U43648 ( .A(p_input[2265]), .B(n43861), .Z(n43509) );
  AND U43649 ( .A(n791), .B(n43862), .Z(n43861) );
  XOR U43650 ( .A(p_input[2297]), .B(p_input[2265]), .Z(n43862) );
  XNOR U43651 ( .A(n43506), .B(n43857), .Z(n43859) );
  XOR U43652 ( .A(n43863), .B(n43864), .Z(n43506) );
  AND U43653 ( .A(n789), .B(n43865), .Z(n43864) );
  XOR U43654 ( .A(p_input[2233]), .B(p_input[2201]), .Z(n43865) );
  XOR U43655 ( .A(n43866), .B(n43867), .Z(n43857) );
  AND U43656 ( .A(n43868), .B(n43869), .Z(n43867) );
  XOR U43657 ( .A(n43866), .B(n43521), .Z(n43869) );
  XNOR U43658 ( .A(p_input[2264]), .B(n43870), .Z(n43521) );
  AND U43659 ( .A(n791), .B(n43871), .Z(n43870) );
  XOR U43660 ( .A(p_input[2296]), .B(p_input[2264]), .Z(n43871) );
  XNOR U43661 ( .A(n43518), .B(n43866), .Z(n43868) );
  XOR U43662 ( .A(n43872), .B(n43873), .Z(n43518) );
  AND U43663 ( .A(n789), .B(n43874), .Z(n43873) );
  XOR U43664 ( .A(p_input[2232]), .B(p_input[2200]), .Z(n43874) );
  XOR U43665 ( .A(n43875), .B(n43876), .Z(n43866) );
  AND U43666 ( .A(n43877), .B(n43878), .Z(n43876) );
  XOR U43667 ( .A(n43875), .B(n43533), .Z(n43878) );
  XNOR U43668 ( .A(p_input[2263]), .B(n43879), .Z(n43533) );
  AND U43669 ( .A(n791), .B(n43880), .Z(n43879) );
  XOR U43670 ( .A(p_input[2295]), .B(p_input[2263]), .Z(n43880) );
  XNOR U43671 ( .A(n43530), .B(n43875), .Z(n43877) );
  XOR U43672 ( .A(n43881), .B(n43882), .Z(n43530) );
  AND U43673 ( .A(n789), .B(n43883), .Z(n43882) );
  XOR U43674 ( .A(p_input[2231]), .B(p_input[2199]), .Z(n43883) );
  XOR U43675 ( .A(n43884), .B(n43885), .Z(n43875) );
  AND U43676 ( .A(n43886), .B(n43887), .Z(n43885) );
  XOR U43677 ( .A(n43884), .B(n43545), .Z(n43887) );
  XNOR U43678 ( .A(p_input[2262]), .B(n43888), .Z(n43545) );
  AND U43679 ( .A(n791), .B(n43889), .Z(n43888) );
  XOR U43680 ( .A(p_input[2294]), .B(p_input[2262]), .Z(n43889) );
  XNOR U43681 ( .A(n43542), .B(n43884), .Z(n43886) );
  XOR U43682 ( .A(n43890), .B(n43891), .Z(n43542) );
  AND U43683 ( .A(n789), .B(n43892), .Z(n43891) );
  XOR U43684 ( .A(p_input[2230]), .B(p_input[2198]), .Z(n43892) );
  XOR U43685 ( .A(n43893), .B(n43894), .Z(n43884) );
  AND U43686 ( .A(n43895), .B(n43896), .Z(n43894) );
  XOR U43687 ( .A(n43893), .B(n43557), .Z(n43896) );
  XNOR U43688 ( .A(p_input[2261]), .B(n43897), .Z(n43557) );
  AND U43689 ( .A(n791), .B(n43898), .Z(n43897) );
  XOR U43690 ( .A(p_input[2293]), .B(p_input[2261]), .Z(n43898) );
  XNOR U43691 ( .A(n43554), .B(n43893), .Z(n43895) );
  XOR U43692 ( .A(n43899), .B(n43900), .Z(n43554) );
  AND U43693 ( .A(n789), .B(n43901), .Z(n43900) );
  XOR U43694 ( .A(p_input[2229]), .B(p_input[2197]), .Z(n43901) );
  XOR U43695 ( .A(n43902), .B(n43903), .Z(n43893) );
  AND U43696 ( .A(n43904), .B(n43905), .Z(n43903) );
  XOR U43697 ( .A(n43902), .B(n43569), .Z(n43905) );
  XNOR U43698 ( .A(p_input[2260]), .B(n43906), .Z(n43569) );
  AND U43699 ( .A(n791), .B(n43907), .Z(n43906) );
  XOR U43700 ( .A(p_input[2292]), .B(p_input[2260]), .Z(n43907) );
  XNOR U43701 ( .A(n43566), .B(n43902), .Z(n43904) );
  XOR U43702 ( .A(n43908), .B(n43909), .Z(n43566) );
  AND U43703 ( .A(n789), .B(n43910), .Z(n43909) );
  XOR U43704 ( .A(p_input[2228]), .B(p_input[2196]), .Z(n43910) );
  XOR U43705 ( .A(n43911), .B(n43912), .Z(n43902) );
  AND U43706 ( .A(n43913), .B(n43914), .Z(n43912) );
  XOR U43707 ( .A(n43911), .B(n43581), .Z(n43914) );
  XNOR U43708 ( .A(p_input[2259]), .B(n43915), .Z(n43581) );
  AND U43709 ( .A(n791), .B(n43916), .Z(n43915) );
  XOR U43710 ( .A(p_input[2291]), .B(p_input[2259]), .Z(n43916) );
  XNOR U43711 ( .A(n43578), .B(n43911), .Z(n43913) );
  XOR U43712 ( .A(n43917), .B(n43918), .Z(n43578) );
  AND U43713 ( .A(n789), .B(n43919), .Z(n43918) );
  XOR U43714 ( .A(p_input[2227]), .B(p_input[2195]), .Z(n43919) );
  XOR U43715 ( .A(n43920), .B(n43921), .Z(n43911) );
  AND U43716 ( .A(n43922), .B(n43923), .Z(n43921) );
  XOR U43717 ( .A(n43920), .B(n43593), .Z(n43923) );
  XNOR U43718 ( .A(p_input[2258]), .B(n43924), .Z(n43593) );
  AND U43719 ( .A(n791), .B(n43925), .Z(n43924) );
  XOR U43720 ( .A(p_input[2290]), .B(p_input[2258]), .Z(n43925) );
  XNOR U43721 ( .A(n43590), .B(n43920), .Z(n43922) );
  XOR U43722 ( .A(n43926), .B(n43927), .Z(n43590) );
  AND U43723 ( .A(n789), .B(n43928), .Z(n43927) );
  XOR U43724 ( .A(p_input[2226]), .B(p_input[2194]), .Z(n43928) );
  XOR U43725 ( .A(n43929), .B(n43930), .Z(n43920) );
  AND U43726 ( .A(n43931), .B(n43932), .Z(n43930) );
  XOR U43727 ( .A(n43929), .B(n43605), .Z(n43932) );
  XNOR U43728 ( .A(p_input[2257]), .B(n43933), .Z(n43605) );
  AND U43729 ( .A(n791), .B(n43934), .Z(n43933) );
  XOR U43730 ( .A(p_input[2289]), .B(p_input[2257]), .Z(n43934) );
  XNOR U43731 ( .A(n43602), .B(n43929), .Z(n43931) );
  XOR U43732 ( .A(n43935), .B(n43936), .Z(n43602) );
  AND U43733 ( .A(n789), .B(n43937), .Z(n43936) );
  XOR U43734 ( .A(p_input[2225]), .B(p_input[2193]), .Z(n43937) );
  XOR U43735 ( .A(n43938), .B(n43939), .Z(n43929) );
  AND U43736 ( .A(n43940), .B(n43941), .Z(n43939) );
  XOR U43737 ( .A(n43938), .B(n43617), .Z(n43941) );
  XNOR U43738 ( .A(p_input[2256]), .B(n43942), .Z(n43617) );
  AND U43739 ( .A(n791), .B(n43943), .Z(n43942) );
  XOR U43740 ( .A(p_input[2288]), .B(p_input[2256]), .Z(n43943) );
  XNOR U43741 ( .A(n43614), .B(n43938), .Z(n43940) );
  XOR U43742 ( .A(n43944), .B(n43945), .Z(n43614) );
  AND U43743 ( .A(n789), .B(n43946), .Z(n43945) );
  XOR U43744 ( .A(p_input[2224]), .B(p_input[2192]), .Z(n43946) );
  XOR U43745 ( .A(n43947), .B(n43948), .Z(n43938) );
  AND U43746 ( .A(n43949), .B(n43950), .Z(n43948) );
  XOR U43747 ( .A(n43947), .B(n43629), .Z(n43950) );
  XNOR U43748 ( .A(p_input[2255]), .B(n43951), .Z(n43629) );
  AND U43749 ( .A(n791), .B(n43952), .Z(n43951) );
  XOR U43750 ( .A(p_input[2287]), .B(p_input[2255]), .Z(n43952) );
  XNOR U43751 ( .A(n43626), .B(n43947), .Z(n43949) );
  XOR U43752 ( .A(n43953), .B(n43954), .Z(n43626) );
  AND U43753 ( .A(n789), .B(n43955), .Z(n43954) );
  XOR U43754 ( .A(p_input[2223]), .B(p_input[2191]), .Z(n43955) );
  XOR U43755 ( .A(n43956), .B(n43957), .Z(n43947) );
  AND U43756 ( .A(n43958), .B(n43959), .Z(n43957) );
  XOR U43757 ( .A(n43956), .B(n43641), .Z(n43959) );
  XNOR U43758 ( .A(p_input[2254]), .B(n43960), .Z(n43641) );
  AND U43759 ( .A(n791), .B(n43961), .Z(n43960) );
  XOR U43760 ( .A(p_input[2286]), .B(p_input[2254]), .Z(n43961) );
  XNOR U43761 ( .A(n43638), .B(n43956), .Z(n43958) );
  XOR U43762 ( .A(n43962), .B(n43963), .Z(n43638) );
  AND U43763 ( .A(n789), .B(n43964), .Z(n43963) );
  XOR U43764 ( .A(p_input[2222]), .B(p_input[2190]), .Z(n43964) );
  XOR U43765 ( .A(n43965), .B(n43966), .Z(n43956) );
  AND U43766 ( .A(n43967), .B(n43968), .Z(n43966) );
  XOR U43767 ( .A(n43965), .B(n43653), .Z(n43968) );
  XNOR U43768 ( .A(p_input[2253]), .B(n43969), .Z(n43653) );
  AND U43769 ( .A(n791), .B(n43970), .Z(n43969) );
  XOR U43770 ( .A(p_input[2285]), .B(p_input[2253]), .Z(n43970) );
  XNOR U43771 ( .A(n43650), .B(n43965), .Z(n43967) );
  XOR U43772 ( .A(n43971), .B(n43972), .Z(n43650) );
  AND U43773 ( .A(n789), .B(n43973), .Z(n43972) );
  XOR U43774 ( .A(p_input[2221]), .B(p_input[2189]), .Z(n43973) );
  XOR U43775 ( .A(n43974), .B(n43975), .Z(n43965) );
  AND U43776 ( .A(n43976), .B(n43977), .Z(n43975) );
  XOR U43777 ( .A(n43974), .B(n43665), .Z(n43977) );
  XNOR U43778 ( .A(p_input[2252]), .B(n43978), .Z(n43665) );
  AND U43779 ( .A(n791), .B(n43979), .Z(n43978) );
  XOR U43780 ( .A(p_input[2284]), .B(p_input[2252]), .Z(n43979) );
  XNOR U43781 ( .A(n43662), .B(n43974), .Z(n43976) );
  XOR U43782 ( .A(n43980), .B(n43981), .Z(n43662) );
  AND U43783 ( .A(n789), .B(n43982), .Z(n43981) );
  XOR U43784 ( .A(p_input[2220]), .B(p_input[2188]), .Z(n43982) );
  XOR U43785 ( .A(n43983), .B(n43984), .Z(n43974) );
  AND U43786 ( .A(n43985), .B(n43986), .Z(n43984) );
  XOR U43787 ( .A(n43983), .B(n43677), .Z(n43986) );
  XNOR U43788 ( .A(p_input[2251]), .B(n43987), .Z(n43677) );
  AND U43789 ( .A(n791), .B(n43988), .Z(n43987) );
  XOR U43790 ( .A(p_input[2283]), .B(p_input[2251]), .Z(n43988) );
  XNOR U43791 ( .A(n43674), .B(n43983), .Z(n43985) );
  XOR U43792 ( .A(n43989), .B(n43990), .Z(n43674) );
  AND U43793 ( .A(n789), .B(n43991), .Z(n43990) );
  XOR U43794 ( .A(p_input[2219]), .B(p_input[2187]), .Z(n43991) );
  XOR U43795 ( .A(n43992), .B(n43993), .Z(n43983) );
  AND U43796 ( .A(n43994), .B(n43995), .Z(n43993) );
  XOR U43797 ( .A(n43992), .B(n43689), .Z(n43995) );
  XNOR U43798 ( .A(p_input[2250]), .B(n43996), .Z(n43689) );
  AND U43799 ( .A(n791), .B(n43997), .Z(n43996) );
  XOR U43800 ( .A(p_input[2282]), .B(p_input[2250]), .Z(n43997) );
  XNOR U43801 ( .A(n43686), .B(n43992), .Z(n43994) );
  XOR U43802 ( .A(n43998), .B(n43999), .Z(n43686) );
  AND U43803 ( .A(n789), .B(n44000), .Z(n43999) );
  XOR U43804 ( .A(p_input[2218]), .B(p_input[2186]), .Z(n44000) );
  XOR U43805 ( .A(n44001), .B(n44002), .Z(n43992) );
  AND U43806 ( .A(n44003), .B(n44004), .Z(n44002) );
  XOR U43807 ( .A(n44001), .B(n43701), .Z(n44004) );
  XNOR U43808 ( .A(p_input[2249]), .B(n44005), .Z(n43701) );
  AND U43809 ( .A(n791), .B(n44006), .Z(n44005) );
  XOR U43810 ( .A(p_input[2281]), .B(p_input[2249]), .Z(n44006) );
  XNOR U43811 ( .A(n43698), .B(n44001), .Z(n44003) );
  XOR U43812 ( .A(n44007), .B(n44008), .Z(n43698) );
  AND U43813 ( .A(n789), .B(n44009), .Z(n44008) );
  XOR U43814 ( .A(p_input[2217]), .B(p_input[2185]), .Z(n44009) );
  XOR U43815 ( .A(n44010), .B(n44011), .Z(n44001) );
  AND U43816 ( .A(n44012), .B(n44013), .Z(n44011) );
  XOR U43817 ( .A(n44010), .B(n43713), .Z(n44013) );
  XNOR U43818 ( .A(p_input[2248]), .B(n44014), .Z(n43713) );
  AND U43819 ( .A(n791), .B(n44015), .Z(n44014) );
  XOR U43820 ( .A(p_input[2280]), .B(p_input[2248]), .Z(n44015) );
  XNOR U43821 ( .A(n43710), .B(n44010), .Z(n44012) );
  XOR U43822 ( .A(n44016), .B(n44017), .Z(n43710) );
  AND U43823 ( .A(n789), .B(n44018), .Z(n44017) );
  XOR U43824 ( .A(p_input[2216]), .B(p_input[2184]), .Z(n44018) );
  XOR U43825 ( .A(n44019), .B(n44020), .Z(n44010) );
  AND U43826 ( .A(n44021), .B(n44022), .Z(n44020) );
  XOR U43827 ( .A(n44019), .B(n43725), .Z(n44022) );
  XNOR U43828 ( .A(p_input[2247]), .B(n44023), .Z(n43725) );
  AND U43829 ( .A(n791), .B(n44024), .Z(n44023) );
  XOR U43830 ( .A(p_input[2279]), .B(p_input[2247]), .Z(n44024) );
  XNOR U43831 ( .A(n43722), .B(n44019), .Z(n44021) );
  XOR U43832 ( .A(n44025), .B(n44026), .Z(n43722) );
  AND U43833 ( .A(n789), .B(n44027), .Z(n44026) );
  XOR U43834 ( .A(p_input[2215]), .B(p_input[2183]), .Z(n44027) );
  XOR U43835 ( .A(n44028), .B(n44029), .Z(n44019) );
  AND U43836 ( .A(n44030), .B(n44031), .Z(n44029) );
  XOR U43837 ( .A(n44028), .B(n43737), .Z(n44031) );
  XNOR U43838 ( .A(p_input[2246]), .B(n44032), .Z(n43737) );
  AND U43839 ( .A(n791), .B(n44033), .Z(n44032) );
  XOR U43840 ( .A(p_input[2278]), .B(p_input[2246]), .Z(n44033) );
  XNOR U43841 ( .A(n43734), .B(n44028), .Z(n44030) );
  XOR U43842 ( .A(n44034), .B(n44035), .Z(n43734) );
  AND U43843 ( .A(n789), .B(n44036), .Z(n44035) );
  XOR U43844 ( .A(p_input[2214]), .B(p_input[2182]), .Z(n44036) );
  XOR U43845 ( .A(n44037), .B(n44038), .Z(n44028) );
  AND U43846 ( .A(n44039), .B(n44040), .Z(n44038) );
  XOR U43847 ( .A(n44037), .B(n43749), .Z(n44040) );
  XNOR U43848 ( .A(p_input[2245]), .B(n44041), .Z(n43749) );
  AND U43849 ( .A(n791), .B(n44042), .Z(n44041) );
  XOR U43850 ( .A(p_input[2277]), .B(p_input[2245]), .Z(n44042) );
  XNOR U43851 ( .A(n43746), .B(n44037), .Z(n44039) );
  XOR U43852 ( .A(n44043), .B(n44044), .Z(n43746) );
  AND U43853 ( .A(n789), .B(n44045), .Z(n44044) );
  XOR U43854 ( .A(p_input[2213]), .B(p_input[2181]), .Z(n44045) );
  XOR U43855 ( .A(n44046), .B(n44047), .Z(n44037) );
  AND U43856 ( .A(n44048), .B(n44049), .Z(n44047) );
  XOR U43857 ( .A(n44046), .B(n43761), .Z(n44049) );
  XNOR U43858 ( .A(p_input[2244]), .B(n44050), .Z(n43761) );
  AND U43859 ( .A(n791), .B(n44051), .Z(n44050) );
  XOR U43860 ( .A(p_input[2276]), .B(p_input[2244]), .Z(n44051) );
  XNOR U43861 ( .A(n43758), .B(n44046), .Z(n44048) );
  XOR U43862 ( .A(n44052), .B(n44053), .Z(n43758) );
  AND U43863 ( .A(n789), .B(n44054), .Z(n44053) );
  XOR U43864 ( .A(p_input[2212]), .B(p_input[2180]), .Z(n44054) );
  XOR U43865 ( .A(n44055), .B(n44056), .Z(n44046) );
  AND U43866 ( .A(n44057), .B(n44058), .Z(n44056) );
  XOR U43867 ( .A(n44055), .B(n43773), .Z(n44058) );
  XNOR U43868 ( .A(p_input[2243]), .B(n44059), .Z(n43773) );
  AND U43869 ( .A(n791), .B(n44060), .Z(n44059) );
  XOR U43870 ( .A(p_input[2275]), .B(p_input[2243]), .Z(n44060) );
  XNOR U43871 ( .A(n43770), .B(n44055), .Z(n44057) );
  XOR U43872 ( .A(n44061), .B(n44062), .Z(n43770) );
  AND U43873 ( .A(n789), .B(n44063), .Z(n44062) );
  XOR U43874 ( .A(p_input[2211]), .B(p_input[2179]), .Z(n44063) );
  XOR U43875 ( .A(n44064), .B(n44065), .Z(n44055) );
  AND U43876 ( .A(n44066), .B(n44067), .Z(n44065) );
  XOR U43877 ( .A(n44064), .B(n43785), .Z(n44067) );
  XNOR U43878 ( .A(p_input[2242]), .B(n44068), .Z(n43785) );
  AND U43879 ( .A(n791), .B(n44069), .Z(n44068) );
  XOR U43880 ( .A(p_input[2274]), .B(p_input[2242]), .Z(n44069) );
  XNOR U43881 ( .A(n43782), .B(n44064), .Z(n44066) );
  XOR U43882 ( .A(n44070), .B(n44071), .Z(n43782) );
  AND U43883 ( .A(n789), .B(n44072), .Z(n44071) );
  XOR U43884 ( .A(p_input[2210]), .B(p_input[2178]), .Z(n44072) );
  XOR U43885 ( .A(n44073), .B(n44074), .Z(n44064) );
  AND U43886 ( .A(n44075), .B(n44076), .Z(n44074) );
  XNOR U43887 ( .A(n44077), .B(n43798), .Z(n44076) );
  XNOR U43888 ( .A(p_input[2241]), .B(n44078), .Z(n43798) );
  AND U43889 ( .A(n791), .B(n44079), .Z(n44078) );
  XNOR U43890 ( .A(p_input[2273]), .B(n44080), .Z(n44079) );
  IV U43891 ( .A(p_input[2241]), .Z(n44080) );
  XNOR U43892 ( .A(n43795), .B(n44073), .Z(n44075) );
  XNOR U43893 ( .A(p_input[2177]), .B(n44081), .Z(n43795) );
  AND U43894 ( .A(n789), .B(n44082), .Z(n44081) );
  XOR U43895 ( .A(p_input[2209]), .B(p_input[2177]), .Z(n44082) );
  IV U43896 ( .A(n44077), .Z(n44073) );
  AND U43897 ( .A(n43803), .B(n43806), .Z(n44077) );
  XOR U43898 ( .A(p_input[2240]), .B(n44083), .Z(n43806) );
  AND U43899 ( .A(n791), .B(n44084), .Z(n44083) );
  XOR U43900 ( .A(p_input[2272]), .B(p_input[2240]), .Z(n44084) );
  XOR U43901 ( .A(n44085), .B(n44086), .Z(n791) );
  AND U43902 ( .A(n44087), .B(n44088), .Z(n44086) );
  XNOR U43903 ( .A(p_input[2303]), .B(n44085), .Z(n44088) );
  XOR U43904 ( .A(n44085), .B(p_input[2271]), .Z(n44087) );
  XOR U43905 ( .A(n44089), .B(n44090), .Z(n44085) );
  AND U43906 ( .A(n44091), .B(n44092), .Z(n44090) );
  XNOR U43907 ( .A(p_input[2302]), .B(n44089), .Z(n44092) );
  XOR U43908 ( .A(n44089), .B(p_input[2270]), .Z(n44091) );
  XOR U43909 ( .A(n44093), .B(n44094), .Z(n44089) );
  AND U43910 ( .A(n44095), .B(n44096), .Z(n44094) );
  XNOR U43911 ( .A(p_input[2301]), .B(n44093), .Z(n44096) );
  XOR U43912 ( .A(n44093), .B(p_input[2269]), .Z(n44095) );
  XOR U43913 ( .A(n44097), .B(n44098), .Z(n44093) );
  AND U43914 ( .A(n44099), .B(n44100), .Z(n44098) );
  XNOR U43915 ( .A(p_input[2300]), .B(n44097), .Z(n44100) );
  XOR U43916 ( .A(n44097), .B(p_input[2268]), .Z(n44099) );
  XOR U43917 ( .A(n44101), .B(n44102), .Z(n44097) );
  AND U43918 ( .A(n44103), .B(n44104), .Z(n44102) );
  XNOR U43919 ( .A(p_input[2299]), .B(n44101), .Z(n44104) );
  XOR U43920 ( .A(n44101), .B(p_input[2267]), .Z(n44103) );
  XOR U43921 ( .A(n44105), .B(n44106), .Z(n44101) );
  AND U43922 ( .A(n44107), .B(n44108), .Z(n44106) );
  XNOR U43923 ( .A(p_input[2298]), .B(n44105), .Z(n44108) );
  XOR U43924 ( .A(n44105), .B(p_input[2266]), .Z(n44107) );
  XOR U43925 ( .A(n44109), .B(n44110), .Z(n44105) );
  AND U43926 ( .A(n44111), .B(n44112), .Z(n44110) );
  XNOR U43927 ( .A(p_input[2297]), .B(n44109), .Z(n44112) );
  XOR U43928 ( .A(n44109), .B(p_input[2265]), .Z(n44111) );
  XOR U43929 ( .A(n44113), .B(n44114), .Z(n44109) );
  AND U43930 ( .A(n44115), .B(n44116), .Z(n44114) );
  XNOR U43931 ( .A(p_input[2296]), .B(n44113), .Z(n44116) );
  XOR U43932 ( .A(n44113), .B(p_input[2264]), .Z(n44115) );
  XOR U43933 ( .A(n44117), .B(n44118), .Z(n44113) );
  AND U43934 ( .A(n44119), .B(n44120), .Z(n44118) );
  XNOR U43935 ( .A(p_input[2295]), .B(n44117), .Z(n44120) );
  XOR U43936 ( .A(n44117), .B(p_input[2263]), .Z(n44119) );
  XOR U43937 ( .A(n44121), .B(n44122), .Z(n44117) );
  AND U43938 ( .A(n44123), .B(n44124), .Z(n44122) );
  XNOR U43939 ( .A(p_input[2294]), .B(n44121), .Z(n44124) );
  XOR U43940 ( .A(n44121), .B(p_input[2262]), .Z(n44123) );
  XOR U43941 ( .A(n44125), .B(n44126), .Z(n44121) );
  AND U43942 ( .A(n44127), .B(n44128), .Z(n44126) );
  XNOR U43943 ( .A(p_input[2293]), .B(n44125), .Z(n44128) );
  XOR U43944 ( .A(n44125), .B(p_input[2261]), .Z(n44127) );
  XOR U43945 ( .A(n44129), .B(n44130), .Z(n44125) );
  AND U43946 ( .A(n44131), .B(n44132), .Z(n44130) );
  XNOR U43947 ( .A(p_input[2292]), .B(n44129), .Z(n44132) );
  XOR U43948 ( .A(n44129), .B(p_input[2260]), .Z(n44131) );
  XOR U43949 ( .A(n44133), .B(n44134), .Z(n44129) );
  AND U43950 ( .A(n44135), .B(n44136), .Z(n44134) );
  XNOR U43951 ( .A(p_input[2291]), .B(n44133), .Z(n44136) );
  XOR U43952 ( .A(n44133), .B(p_input[2259]), .Z(n44135) );
  XOR U43953 ( .A(n44137), .B(n44138), .Z(n44133) );
  AND U43954 ( .A(n44139), .B(n44140), .Z(n44138) );
  XNOR U43955 ( .A(p_input[2290]), .B(n44137), .Z(n44140) );
  XOR U43956 ( .A(n44137), .B(p_input[2258]), .Z(n44139) );
  XOR U43957 ( .A(n44141), .B(n44142), .Z(n44137) );
  AND U43958 ( .A(n44143), .B(n44144), .Z(n44142) );
  XNOR U43959 ( .A(p_input[2289]), .B(n44141), .Z(n44144) );
  XOR U43960 ( .A(n44141), .B(p_input[2257]), .Z(n44143) );
  XOR U43961 ( .A(n44145), .B(n44146), .Z(n44141) );
  AND U43962 ( .A(n44147), .B(n44148), .Z(n44146) );
  XNOR U43963 ( .A(p_input[2288]), .B(n44145), .Z(n44148) );
  XOR U43964 ( .A(n44145), .B(p_input[2256]), .Z(n44147) );
  XOR U43965 ( .A(n44149), .B(n44150), .Z(n44145) );
  AND U43966 ( .A(n44151), .B(n44152), .Z(n44150) );
  XNOR U43967 ( .A(p_input[2287]), .B(n44149), .Z(n44152) );
  XOR U43968 ( .A(n44149), .B(p_input[2255]), .Z(n44151) );
  XOR U43969 ( .A(n44153), .B(n44154), .Z(n44149) );
  AND U43970 ( .A(n44155), .B(n44156), .Z(n44154) );
  XNOR U43971 ( .A(p_input[2286]), .B(n44153), .Z(n44156) );
  XOR U43972 ( .A(n44153), .B(p_input[2254]), .Z(n44155) );
  XOR U43973 ( .A(n44157), .B(n44158), .Z(n44153) );
  AND U43974 ( .A(n44159), .B(n44160), .Z(n44158) );
  XNOR U43975 ( .A(p_input[2285]), .B(n44157), .Z(n44160) );
  XOR U43976 ( .A(n44157), .B(p_input[2253]), .Z(n44159) );
  XOR U43977 ( .A(n44161), .B(n44162), .Z(n44157) );
  AND U43978 ( .A(n44163), .B(n44164), .Z(n44162) );
  XNOR U43979 ( .A(p_input[2284]), .B(n44161), .Z(n44164) );
  XOR U43980 ( .A(n44161), .B(p_input[2252]), .Z(n44163) );
  XOR U43981 ( .A(n44165), .B(n44166), .Z(n44161) );
  AND U43982 ( .A(n44167), .B(n44168), .Z(n44166) );
  XNOR U43983 ( .A(p_input[2283]), .B(n44165), .Z(n44168) );
  XOR U43984 ( .A(n44165), .B(p_input[2251]), .Z(n44167) );
  XOR U43985 ( .A(n44169), .B(n44170), .Z(n44165) );
  AND U43986 ( .A(n44171), .B(n44172), .Z(n44170) );
  XNOR U43987 ( .A(p_input[2282]), .B(n44169), .Z(n44172) );
  XOR U43988 ( .A(n44169), .B(p_input[2250]), .Z(n44171) );
  XOR U43989 ( .A(n44173), .B(n44174), .Z(n44169) );
  AND U43990 ( .A(n44175), .B(n44176), .Z(n44174) );
  XNOR U43991 ( .A(p_input[2281]), .B(n44173), .Z(n44176) );
  XOR U43992 ( .A(n44173), .B(p_input[2249]), .Z(n44175) );
  XOR U43993 ( .A(n44177), .B(n44178), .Z(n44173) );
  AND U43994 ( .A(n44179), .B(n44180), .Z(n44178) );
  XNOR U43995 ( .A(p_input[2280]), .B(n44177), .Z(n44180) );
  XOR U43996 ( .A(n44177), .B(p_input[2248]), .Z(n44179) );
  XOR U43997 ( .A(n44181), .B(n44182), .Z(n44177) );
  AND U43998 ( .A(n44183), .B(n44184), .Z(n44182) );
  XNOR U43999 ( .A(p_input[2279]), .B(n44181), .Z(n44184) );
  XOR U44000 ( .A(n44181), .B(p_input[2247]), .Z(n44183) );
  XOR U44001 ( .A(n44185), .B(n44186), .Z(n44181) );
  AND U44002 ( .A(n44187), .B(n44188), .Z(n44186) );
  XNOR U44003 ( .A(p_input[2278]), .B(n44185), .Z(n44188) );
  XOR U44004 ( .A(n44185), .B(p_input[2246]), .Z(n44187) );
  XOR U44005 ( .A(n44189), .B(n44190), .Z(n44185) );
  AND U44006 ( .A(n44191), .B(n44192), .Z(n44190) );
  XNOR U44007 ( .A(p_input[2277]), .B(n44189), .Z(n44192) );
  XOR U44008 ( .A(n44189), .B(p_input[2245]), .Z(n44191) );
  XOR U44009 ( .A(n44193), .B(n44194), .Z(n44189) );
  AND U44010 ( .A(n44195), .B(n44196), .Z(n44194) );
  XNOR U44011 ( .A(p_input[2276]), .B(n44193), .Z(n44196) );
  XOR U44012 ( .A(n44193), .B(p_input[2244]), .Z(n44195) );
  XOR U44013 ( .A(n44197), .B(n44198), .Z(n44193) );
  AND U44014 ( .A(n44199), .B(n44200), .Z(n44198) );
  XNOR U44015 ( .A(p_input[2275]), .B(n44197), .Z(n44200) );
  XOR U44016 ( .A(n44197), .B(p_input[2243]), .Z(n44199) );
  XOR U44017 ( .A(n44201), .B(n44202), .Z(n44197) );
  AND U44018 ( .A(n44203), .B(n44204), .Z(n44202) );
  XNOR U44019 ( .A(p_input[2274]), .B(n44201), .Z(n44204) );
  XOR U44020 ( .A(n44201), .B(p_input[2242]), .Z(n44203) );
  XNOR U44021 ( .A(n44205), .B(n44206), .Z(n44201) );
  AND U44022 ( .A(n44207), .B(n44208), .Z(n44206) );
  XOR U44023 ( .A(p_input[2273]), .B(n44205), .Z(n44208) );
  XNOR U44024 ( .A(p_input[2241]), .B(n44205), .Z(n44207) );
  AND U44025 ( .A(p_input[2272]), .B(n44209), .Z(n44205) );
  IV U44026 ( .A(p_input[2240]), .Z(n44209) );
  XNOR U44027 ( .A(p_input[2176]), .B(n44210), .Z(n43803) );
  AND U44028 ( .A(n789), .B(n44211), .Z(n44210) );
  XOR U44029 ( .A(p_input[2208]), .B(p_input[2176]), .Z(n44211) );
  XOR U44030 ( .A(n44212), .B(n44213), .Z(n789) );
  AND U44031 ( .A(n44214), .B(n44215), .Z(n44213) );
  XNOR U44032 ( .A(p_input[2239]), .B(n44212), .Z(n44215) );
  XOR U44033 ( .A(n44212), .B(p_input[2207]), .Z(n44214) );
  XOR U44034 ( .A(n44216), .B(n44217), .Z(n44212) );
  AND U44035 ( .A(n44218), .B(n44219), .Z(n44217) );
  XNOR U44036 ( .A(p_input[2238]), .B(n44216), .Z(n44219) );
  XNOR U44037 ( .A(n44216), .B(n43818), .Z(n44218) );
  IV U44038 ( .A(p_input[2206]), .Z(n43818) );
  XOR U44039 ( .A(n44220), .B(n44221), .Z(n44216) );
  AND U44040 ( .A(n44222), .B(n44223), .Z(n44221) );
  XNOR U44041 ( .A(p_input[2237]), .B(n44220), .Z(n44223) );
  XNOR U44042 ( .A(n44220), .B(n43827), .Z(n44222) );
  IV U44043 ( .A(p_input[2205]), .Z(n43827) );
  XOR U44044 ( .A(n44224), .B(n44225), .Z(n44220) );
  AND U44045 ( .A(n44226), .B(n44227), .Z(n44225) );
  XNOR U44046 ( .A(p_input[2236]), .B(n44224), .Z(n44227) );
  XNOR U44047 ( .A(n44224), .B(n43836), .Z(n44226) );
  IV U44048 ( .A(p_input[2204]), .Z(n43836) );
  XOR U44049 ( .A(n44228), .B(n44229), .Z(n44224) );
  AND U44050 ( .A(n44230), .B(n44231), .Z(n44229) );
  XNOR U44051 ( .A(p_input[2235]), .B(n44228), .Z(n44231) );
  XNOR U44052 ( .A(n44228), .B(n43845), .Z(n44230) );
  IV U44053 ( .A(p_input[2203]), .Z(n43845) );
  XOR U44054 ( .A(n44232), .B(n44233), .Z(n44228) );
  AND U44055 ( .A(n44234), .B(n44235), .Z(n44233) );
  XNOR U44056 ( .A(p_input[2234]), .B(n44232), .Z(n44235) );
  XNOR U44057 ( .A(n44232), .B(n43854), .Z(n44234) );
  IV U44058 ( .A(p_input[2202]), .Z(n43854) );
  XOR U44059 ( .A(n44236), .B(n44237), .Z(n44232) );
  AND U44060 ( .A(n44238), .B(n44239), .Z(n44237) );
  XNOR U44061 ( .A(p_input[2233]), .B(n44236), .Z(n44239) );
  XNOR U44062 ( .A(n44236), .B(n43863), .Z(n44238) );
  IV U44063 ( .A(p_input[2201]), .Z(n43863) );
  XOR U44064 ( .A(n44240), .B(n44241), .Z(n44236) );
  AND U44065 ( .A(n44242), .B(n44243), .Z(n44241) );
  XNOR U44066 ( .A(p_input[2232]), .B(n44240), .Z(n44243) );
  XNOR U44067 ( .A(n44240), .B(n43872), .Z(n44242) );
  IV U44068 ( .A(p_input[2200]), .Z(n43872) );
  XOR U44069 ( .A(n44244), .B(n44245), .Z(n44240) );
  AND U44070 ( .A(n44246), .B(n44247), .Z(n44245) );
  XNOR U44071 ( .A(p_input[2231]), .B(n44244), .Z(n44247) );
  XNOR U44072 ( .A(n44244), .B(n43881), .Z(n44246) );
  IV U44073 ( .A(p_input[2199]), .Z(n43881) );
  XOR U44074 ( .A(n44248), .B(n44249), .Z(n44244) );
  AND U44075 ( .A(n44250), .B(n44251), .Z(n44249) );
  XNOR U44076 ( .A(p_input[2230]), .B(n44248), .Z(n44251) );
  XNOR U44077 ( .A(n44248), .B(n43890), .Z(n44250) );
  IV U44078 ( .A(p_input[2198]), .Z(n43890) );
  XOR U44079 ( .A(n44252), .B(n44253), .Z(n44248) );
  AND U44080 ( .A(n44254), .B(n44255), .Z(n44253) );
  XNOR U44081 ( .A(p_input[2229]), .B(n44252), .Z(n44255) );
  XNOR U44082 ( .A(n44252), .B(n43899), .Z(n44254) );
  IV U44083 ( .A(p_input[2197]), .Z(n43899) );
  XOR U44084 ( .A(n44256), .B(n44257), .Z(n44252) );
  AND U44085 ( .A(n44258), .B(n44259), .Z(n44257) );
  XNOR U44086 ( .A(p_input[2228]), .B(n44256), .Z(n44259) );
  XNOR U44087 ( .A(n44256), .B(n43908), .Z(n44258) );
  IV U44088 ( .A(p_input[2196]), .Z(n43908) );
  XOR U44089 ( .A(n44260), .B(n44261), .Z(n44256) );
  AND U44090 ( .A(n44262), .B(n44263), .Z(n44261) );
  XNOR U44091 ( .A(p_input[2227]), .B(n44260), .Z(n44263) );
  XNOR U44092 ( .A(n44260), .B(n43917), .Z(n44262) );
  IV U44093 ( .A(p_input[2195]), .Z(n43917) );
  XOR U44094 ( .A(n44264), .B(n44265), .Z(n44260) );
  AND U44095 ( .A(n44266), .B(n44267), .Z(n44265) );
  XNOR U44096 ( .A(p_input[2226]), .B(n44264), .Z(n44267) );
  XNOR U44097 ( .A(n44264), .B(n43926), .Z(n44266) );
  IV U44098 ( .A(p_input[2194]), .Z(n43926) );
  XOR U44099 ( .A(n44268), .B(n44269), .Z(n44264) );
  AND U44100 ( .A(n44270), .B(n44271), .Z(n44269) );
  XNOR U44101 ( .A(p_input[2225]), .B(n44268), .Z(n44271) );
  XNOR U44102 ( .A(n44268), .B(n43935), .Z(n44270) );
  IV U44103 ( .A(p_input[2193]), .Z(n43935) );
  XOR U44104 ( .A(n44272), .B(n44273), .Z(n44268) );
  AND U44105 ( .A(n44274), .B(n44275), .Z(n44273) );
  XNOR U44106 ( .A(p_input[2224]), .B(n44272), .Z(n44275) );
  XNOR U44107 ( .A(n44272), .B(n43944), .Z(n44274) );
  IV U44108 ( .A(p_input[2192]), .Z(n43944) );
  XOR U44109 ( .A(n44276), .B(n44277), .Z(n44272) );
  AND U44110 ( .A(n44278), .B(n44279), .Z(n44277) );
  XNOR U44111 ( .A(p_input[2223]), .B(n44276), .Z(n44279) );
  XNOR U44112 ( .A(n44276), .B(n43953), .Z(n44278) );
  IV U44113 ( .A(p_input[2191]), .Z(n43953) );
  XOR U44114 ( .A(n44280), .B(n44281), .Z(n44276) );
  AND U44115 ( .A(n44282), .B(n44283), .Z(n44281) );
  XNOR U44116 ( .A(p_input[2222]), .B(n44280), .Z(n44283) );
  XNOR U44117 ( .A(n44280), .B(n43962), .Z(n44282) );
  IV U44118 ( .A(p_input[2190]), .Z(n43962) );
  XOR U44119 ( .A(n44284), .B(n44285), .Z(n44280) );
  AND U44120 ( .A(n44286), .B(n44287), .Z(n44285) );
  XNOR U44121 ( .A(p_input[2221]), .B(n44284), .Z(n44287) );
  XNOR U44122 ( .A(n44284), .B(n43971), .Z(n44286) );
  IV U44123 ( .A(p_input[2189]), .Z(n43971) );
  XOR U44124 ( .A(n44288), .B(n44289), .Z(n44284) );
  AND U44125 ( .A(n44290), .B(n44291), .Z(n44289) );
  XNOR U44126 ( .A(p_input[2220]), .B(n44288), .Z(n44291) );
  XNOR U44127 ( .A(n44288), .B(n43980), .Z(n44290) );
  IV U44128 ( .A(p_input[2188]), .Z(n43980) );
  XOR U44129 ( .A(n44292), .B(n44293), .Z(n44288) );
  AND U44130 ( .A(n44294), .B(n44295), .Z(n44293) );
  XNOR U44131 ( .A(p_input[2219]), .B(n44292), .Z(n44295) );
  XNOR U44132 ( .A(n44292), .B(n43989), .Z(n44294) );
  IV U44133 ( .A(p_input[2187]), .Z(n43989) );
  XOR U44134 ( .A(n44296), .B(n44297), .Z(n44292) );
  AND U44135 ( .A(n44298), .B(n44299), .Z(n44297) );
  XNOR U44136 ( .A(p_input[2218]), .B(n44296), .Z(n44299) );
  XNOR U44137 ( .A(n44296), .B(n43998), .Z(n44298) );
  IV U44138 ( .A(p_input[2186]), .Z(n43998) );
  XOR U44139 ( .A(n44300), .B(n44301), .Z(n44296) );
  AND U44140 ( .A(n44302), .B(n44303), .Z(n44301) );
  XNOR U44141 ( .A(p_input[2217]), .B(n44300), .Z(n44303) );
  XNOR U44142 ( .A(n44300), .B(n44007), .Z(n44302) );
  IV U44143 ( .A(p_input[2185]), .Z(n44007) );
  XOR U44144 ( .A(n44304), .B(n44305), .Z(n44300) );
  AND U44145 ( .A(n44306), .B(n44307), .Z(n44305) );
  XNOR U44146 ( .A(p_input[2216]), .B(n44304), .Z(n44307) );
  XNOR U44147 ( .A(n44304), .B(n44016), .Z(n44306) );
  IV U44148 ( .A(p_input[2184]), .Z(n44016) );
  XOR U44149 ( .A(n44308), .B(n44309), .Z(n44304) );
  AND U44150 ( .A(n44310), .B(n44311), .Z(n44309) );
  XNOR U44151 ( .A(p_input[2215]), .B(n44308), .Z(n44311) );
  XNOR U44152 ( .A(n44308), .B(n44025), .Z(n44310) );
  IV U44153 ( .A(p_input[2183]), .Z(n44025) );
  XOR U44154 ( .A(n44312), .B(n44313), .Z(n44308) );
  AND U44155 ( .A(n44314), .B(n44315), .Z(n44313) );
  XNOR U44156 ( .A(p_input[2214]), .B(n44312), .Z(n44315) );
  XNOR U44157 ( .A(n44312), .B(n44034), .Z(n44314) );
  IV U44158 ( .A(p_input[2182]), .Z(n44034) );
  XOR U44159 ( .A(n44316), .B(n44317), .Z(n44312) );
  AND U44160 ( .A(n44318), .B(n44319), .Z(n44317) );
  XNOR U44161 ( .A(p_input[2213]), .B(n44316), .Z(n44319) );
  XNOR U44162 ( .A(n44316), .B(n44043), .Z(n44318) );
  IV U44163 ( .A(p_input[2181]), .Z(n44043) );
  XOR U44164 ( .A(n44320), .B(n44321), .Z(n44316) );
  AND U44165 ( .A(n44322), .B(n44323), .Z(n44321) );
  XNOR U44166 ( .A(p_input[2212]), .B(n44320), .Z(n44323) );
  XNOR U44167 ( .A(n44320), .B(n44052), .Z(n44322) );
  IV U44168 ( .A(p_input[2180]), .Z(n44052) );
  XOR U44169 ( .A(n44324), .B(n44325), .Z(n44320) );
  AND U44170 ( .A(n44326), .B(n44327), .Z(n44325) );
  XNOR U44171 ( .A(p_input[2211]), .B(n44324), .Z(n44327) );
  XNOR U44172 ( .A(n44324), .B(n44061), .Z(n44326) );
  IV U44173 ( .A(p_input[2179]), .Z(n44061) );
  XOR U44174 ( .A(n44328), .B(n44329), .Z(n44324) );
  AND U44175 ( .A(n44330), .B(n44331), .Z(n44329) );
  XNOR U44176 ( .A(p_input[2210]), .B(n44328), .Z(n44331) );
  XNOR U44177 ( .A(n44328), .B(n44070), .Z(n44330) );
  IV U44178 ( .A(p_input[2178]), .Z(n44070) );
  XNOR U44179 ( .A(n44332), .B(n44333), .Z(n44328) );
  AND U44180 ( .A(n44334), .B(n44335), .Z(n44333) );
  XOR U44181 ( .A(p_input[2209]), .B(n44332), .Z(n44335) );
  XNOR U44182 ( .A(p_input[2177]), .B(n44332), .Z(n44334) );
  AND U44183 ( .A(p_input[2208]), .B(n44336), .Z(n44332) );
  IV U44184 ( .A(p_input[2176]), .Z(n44336) );
  XOR U44185 ( .A(n44337), .B(n44338), .Z(n43426) );
  AND U44186 ( .A(n604), .B(n44339), .Z(n44338) );
  XNOR U44187 ( .A(n44340), .B(n44337), .Z(n44339) );
  XOR U44188 ( .A(n44341), .B(n44342), .Z(n604) );
  AND U44189 ( .A(n44343), .B(n44344), .Z(n44342) );
  XNOR U44190 ( .A(n43441), .B(n44341), .Z(n44344) );
  AND U44191 ( .A(p_input[2175]), .B(p_input[2143]), .Z(n43441) );
  XNOR U44192 ( .A(n44341), .B(n43438), .Z(n44343) );
  IV U44193 ( .A(n44345), .Z(n43438) );
  AND U44194 ( .A(p_input[2079]), .B(p_input[2111]), .Z(n44345) );
  XOR U44195 ( .A(n44346), .B(n44347), .Z(n44341) );
  AND U44196 ( .A(n44348), .B(n44349), .Z(n44347) );
  XOR U44197 ( .A(n44346), .B(n43453), .Z(n44349) );
  XNOR U44198 ( .A(p_input[2142]), .B(n44350), .Z(n43453) );
  AND U44199 ( .A(n795), .B(n44351), .Z(n44350) );
  XOR U44200 ( .A(p_input[2174]), .B(p_input[2142]), .Z(n44351) );
  XNOR U44201 ( .A(n43450), .B(n44346), .Z(n44348) );
  XOR U44202 ( .A(n44352), .B(n44353), .Z(n43450) );
  AND U44203 ( .A(n792), .B(n44354), .Z(n44353) );
  XOR U44204 ( .A(p_input[2110]), .B(p_input[2078]), .Z(n44354) );
  XOR U44205 ( .A(n44355), .B(n44356), .Z(n44346) );
  AND U44206 ( .A(n44357), .B(n44358), .Z(n44356) );
  XOR U44207 ( .A(n44355), .B(n43465), .Z(n44358) );
  XNOR U44208 ( .A(p_input[2141]), .B(n44359), .Z(n43465) );
  AND U44209 ( .A(n795), .B(n44360), .Z(n44359) );
  XOR U44210 ( .A(p_input[2173]), .B(p_input[2141]), .Z(n44360) );
  XNOR U44211 ( .A(n43462), .B(n44355), .Z(n44357) );
  XOR U44212 ( .A(n44361), .B(n44362), .Z(n43462) );
  AND U44213 ( .A(n792), .B(n44363), .Z(n44362) );
  XOR U44214 ( .A(p_input[2109]), .B(p_input[2077]), .Z(n44363) );
  XOR U44215 ( .A(n44364), .B(n44365), .Z(n44355) );
  AND U44216 ( .A(n44366), .B(n44367), .Z(n44365) );
  XOR U44217 ( .A(n44364), .B(n43477), .Z(n44367) );
  XNOR U44218 ( .A(p_input[2140]), .B(n44368), .Z(n43477) );
  AND U44219 ( .A(n795), .B(n44369), .Z(n44368) );
  XOR U44220 ( .A(p_input[2172]), .B(p_input[2140]), .Z(n44369) );
  XNOR U44221 ( .A(n43474), .B(n44364), .Z(n44366) );
  XOR U44222 ( .A(n44370), .B(n44371), .Z(n43474) );
  AND U44223 ( .A(n792), .B(n44372), .Z(n44371) );
  XOR U44224 ( .A(p_input[2108]), .B(p_input[2076]), .Z(n44372) );
  XOR U44225 ( .A(n44373), .B(n44374), .Z(n44364) );
  AND U44226 ( .A(n44375), .B(n44376), .Z(n44374) );
  XOR U44227 ( .A(n44373), .B(n43489), .Z(n44376) );
  XNOR U44228 ( .A(p_input[2139]), .B(n44377), .Z(n43489) );
  AND U44229 ( .A(n795), .B(n44378), .Z(n44377) );
  XOR U44230 ( .A(p_input[2171]), .B(p_input[2139]), .Z(n44378) );
  XNOR U44231 ( .A(n43486), .B(n44373), .Z(n44375) );
  XOR U44232 ( .A(n44379), .B(n44380), .Z(n43486) );
  AND U44233 ( .A(n792), .B(n44381), .Z(n44380) );
  XOR U44234 ( .A(p_input[2107]), .B(p_input[2075]), .Z(n44381) );
  XOR U44235 ( .A(n44382), .B(n44383), .Z(n44373) );
  AND U44236 ( .A(n44384), .B(n44385), .Z(n44383) );
  XOR U44237 ( .A(n44382), .B(n43501), .Z(n44385) );
  XNOR U44238 ( .A(p_input[2138]), .B(n44386), .Z(n43501) );
  AND U44239 ( .A(n795), .B(n44387), .Z(n44386) );
  XOR U44240 ( .A(p_input[2170]), .B(p_input[2138]), .Z(n44387) );
  XNOR U44241 ( .A(n43498), .B(n44382), .Z(n44384) );
  XOR U44242 ( .A(n44388), .B(n44389), .Z(n43498) );
  AND U44243 ( .A(n792), .B(n44390), .Z(n44389) );
  XOR U44244 ( .A(p_input[2106]), .B(p_input[2074]), .Z(n44390) );
  XOR U44245 ( .A(n44391), .B(n44392), .Z(n44382) );
  AND U44246 ( .A(n44393), .B(n44394), .Z(n44392) );
  XOR U44247 ( .A(n44391), .B(n43513), .Z(n44394) );
  XNOR U44248 ( .A(p_input[2137]), .B(n44395), .Z(n43513) );
  AND U44249 ( .A(n795), .B(n44396), .Z(n44395) );
  XOR U44250 ( .A(p_input[2169]), .B(p_input[2137]), .Z(n44396) );
  XNOR U44251 ( .A(n43510), .B(n44391), .Z(n44393) );
  XOR U44252 ( .A(n44397), .B(n44398), .Z(n43510) );
  AND U44253 ( .A(n792), .B(n44399), .Z(n44398) );
  XOR U44254 ( .A(p_input[2105]), .B(p_input[2073]), .Z(n44399) );
  XOR U44255 ( .A(n44400), .B(n44401), .Z(n44391) );
  AND U44256 ( .A(n44402), .B(n44403), .Z(n44401) );
  XOR U44257 ( .A(n44400), .B(n43525), .Z(n44403) );
  XNOR U44258 ( .A(p_input[2136]), .B(n44404), .Z(n43525) );
  AND U44259 ( .A(n795), .B(n44405), .Z(n44404) );
  XOR U44260 ( .A(p_input[2168]), .B(p_input[2136]), .Z(n44405) );
  XNOR U44261 ( .A(n43522), .B(n44400), .Z(n44402) );
  XOR U44262 ( .A(n44406), .B(n44407), .Z(n43522) );
  AND U44263 ( .A(n792), .B(n44408), .Z(n44407) );
  XOR U44264 ( .A(p_input[2104]), .B(p_input[2072]), .Z(n44408) );
  XOR U44265 ( .A(n44409), .B(n44410), .Z(n44400) );
  AND U44266 ( .A(n44411), .B(n44412), .Z(n44410) );
  XOR U44267 ( .A(n44409), .B(n43537), .Z(n44412) );
  XNOR U44268 ( .A(p_input[2135]), .B(n44413), .Z(n43537) );
  AND U44269 ( .A(n795), .B(n44414), .Z(n44413) );
  XOR U44270 ( .A(p_input[2167]), .B(p_input[2135]), .Z(n44414) );
  XNOR U44271 ( .A(n43534), .B(n44409), .Z(n44411) );
  XOR U44272 ( .A(n44415), .B(n44416), .Z(n43534) );
  AND U44273 ( .A(n792), .B(n44417), .Z(n44416) );
  XOR U44274 ( .A(p_input[2103]), .B(p_input[2071]), .Z(n44417) );
  XOR U44275 ( .A(n44418), .B(n44419), .Z(n44409) );
  AND U44276 ( .A(n44420), .B(n44421), .Z(n44419) );
  XOR U44277 ( .A(n44418), .B(n43549), .Z(n44421) );
  XNOR U44278 ( .A(p_input[2134]), .B(n44422), .Z(n43549) );
  AND U44279 ( .A(n795), .B(n44423), .Z(n44422) );
  XOR U44280 ( .A(p_input[2166]), .B(p_input[2134]), .Z(n44423) );
  XNOR U44281 ( .A(n43546), .B(n44418), .Z(n44420) );
  XOR U44282 ( .A(n44424), .B(n44425), .Z(n43546) );
  AND U44283 ( .A(n792), .B(n44426), .Z(n44425) );
  XOR U44284 ( .A(p_input[2102]), .B(p_input[2070]), .Z(n44426) );
  XOR U44285 ( .A(n44427), .B(n44428), .Z(n44418) );
  AND U44286 ( .A(n44429), .B(n44430), .Z(n44428) );
  XOR U44287 ( .A(n44427), .B(n43561), .Z(n44430) );
  XNOR U44288 ( .A(p_input[2133]), .B(n44431), .Z(n43561) );
  AND U44289 ( .A(n795), .B(n44432), .Z(n44431) );
  XOR U44290 ( .A(p_input[2165]), .B(p_input[2133]), .Z(n44432) );
  XNOR U44291 ( .A(n43558), .B(n44427), .Z(n44429) );
  XOR U44292 ( .A(n44433), .B(n44434), .Z(n43558) );
  AND U44293 ( .A(n792), .B(n44435), .Z(n44434) );
  XOR U44294 ( .A(p_input[2101]), .B(p_input[2069]), .Z(n44435) );
  XOR U44295 ( .A(n44436), .B(n44437), .Z(n44427) );
  AND U44296 ( .A(n44438), .B(n44439), .Z(n44437) );
  XOR U44297 ( .A(n44436), .B(n43573), .Z(n44439) );
  XNOR U44298 ( .A(p_input[2132]), .B(n44440), .Z(n43573) );
  AND U44299 ( .A(n795), .B(n44441), .Z(n44440) );
  XOR U44300 ( .A(p_input[2164]), .B(p_input[2132]), .Z(n44441) );
  XNOR U44301 ( .A(n43570), .B(n44436), .Z(n44438) );
  XOR U44302 ( .A(n44442), .B(n44443), .Z(n43570) );
  AND U44303 ( .A(n792), .B(n44444), .Z(n44443) );
  XOR U44304 ( .A(p_input[2100]), .B(p_input[2068]), .Z(n44444) );
  XOR U44305 ( .A(n44445), .B(n44446), .Z(n44436) );
  AND U44306 ( .A(n44447), .B(n44448), .Z(n44446) );
  XOR U44307 ( .A(n44445), .B(n43585), .Z(n44448) );
  XNOR U44308 ( .A(p_input[2131]), .B(n44449), .Z(n43585) );
  AND U44309 ( .A(n795), .B(n44450), .Z(n44449) );
  XOR U44310 ( .A(p_input[2163]), .B(p_input[2131]), .Z(n44450) );
  XNOR U44311 ( .A(n43582), .B(n44445), .Z(n44447) );
  XOR U44312 ( .A(n44451), .B(n44452), .Z(n43582) );
  AND U44313 ( .A(n792), .B(n44453), .Z(n44452) );
  XOR U44314 ( .A(p_input[2099]), .B(p_input[2067]), .Z(n44453) );
  XOR U44315 ( .A(n44454), .B(n44455), .Z(n44445) );
  AND U44316 ( .A(n44456), .B(n44457), .Z(n44455) );
  XOR U44317 ( .A(n44454), .B(n43597), .Z(n44457) );
  XNOR U44318 ( .A(p_input[2130]), .B(n44458), .Z(n43597) );
  AND U44319 ( .A(n795), .B(n44459), .Z(n44458) );
  XOR U44320 ( .A(p_input[2162]), .B(p_input[2130]), .Z(n44459) );
  XNOR U44321 ( .A(n43594), .B(n44454), .Z(n44456) );
  XOR U44322 ( .A(n44460), .B(n44461), .Z(n43594) );
  AND U44323 ( .A(n792), .B(n44462), .Z(n44461) );
  XOR U44324 ( .A(p_input[2098]), .B(p_input[2066]), .Z(n44462) );
  XOR U44325 ( .A(n44463), .B(n44464), .Z(n44454) );
  AND U44326 ( .A(n44465), .B(n44466), .Z(n44464) );
  XOR U44327 ( .A(n44463), .B(n43609), .Z(n44466) );
  XNOR U44328 ( .A(p_input[2129]), .B(n44467), .Z(n43609) );
  AND U44329 ( .A(n795), .B(n44468), .Z(n44467) );
  XOR U44330 ( .A(p_input[2161]), .B(p_input[2129]), .Z(n44468) );
  XNOR U44331 ( .A(n43606), .B(n44463), .Z(n44465) );
  XOR U44332 ( .A(n44469), .B(n44470), .Z(n43606) );
  AND U44333 ( .A(n792), .B(n44471), .Z(n44470) );
  XOR U44334 ( .A(p_input[2097]), .B(p_input[2065]), .Z(n44471) );
  XOR U44335 ( .A(n44472), .B(n44473), .Z(n44463) );
  AND U44336 ( .A(n44474), .B(n44475), .Z(n44473) );
  XOR U44337 ( .A(n44472), .B(n43621), .Z(n44475) );
  XNOR U44338 ( .A(p_input[2128]), .B(n44476), .Z(n43621) );
  AND U44339 ( .A(n795), .B(n44477), .Z(n44476) );
  XOR U44340 ( .A(p_input[2160]), .B(p_input[2128]), .Z(n44477) );
  XNOR U44341 ( .A(n43618), .B(n44472), .Z(n44474) );
  XOR U44342 ( .A(n44478), .B(n44479), .Z(n43618) );
  AND U44343 ( .A(n792), .B(n44480), .Z(n44479) );
  XOR U44344 ( .A(p_input[2096]), .B(p_input[2064]), .Z(n44480) );
  XOR U44345 ( .A(n44481), .B(n44482), .Z(n44472) );
  AND U44346 ( .A(n44483), .B(n44484), .Z(n44482) );
  XOR U44347 ( .A(n44481), .B(n43633), .Z(n44484) );
  XNOR U44348 ( .A(p_input[2127]), .B(n44485), .Z(n43633) );
  AND U44349 ( .A(n795), .B(n44486), .Z(n44485) );
  XOR U44350 ( .A(p_input[2159]), .B(p_input[2127]), .Z(n44486) );
  XNOR U44351 ( .A(n43630), .B(n44481), .Z(n44483) );
  XOR U44352 ( .A(n44487), .B(n44488), .Z(n43630) );
  AND U44353 ( .A(n792), .B(n44489), .Z(n44488) );
  XOR U44354 ( .A(p_input[2095]), .B(p_input[2063]), .Z(n44489) );
  XOR U44355 ( .A(n44490), .B(n44491), .Z(n44481) );
  AND U44356 ( .A(n44492), .B(n44493), .Z(n44491) );
  XOR U44357 ( .A(n44490), .B(n43645), .Z(n44493) );
  XNOR U44358 ( .A(p_input[2126]), .B(n44494), .Z(n43645) );
  AND U44359 ( .A(n795), .B(n44495), .Z(n44494) );
  XOR U44360 ( .A(p_input[2158]), .B(p_input[2126]), .Z(n44495) );
  XNOR U44361 ( .A(n43642), .B(n44490), .Z(n44492) );
  XOR U44362 ( .A(n44496), .B(n44497), .Z(n43642) );
  AND U44363 ( .A(n792), .B(n44498), .Z(n44497) );
  XOR U44364 ( .A(p_input[2094]), .B(p_input[2062]), .Z(n44498) );
  XOR U44365 ( .A(n44499), .B(n44500), .Z(n44490) );
  AND U44366 ( .A(n44501), .B(n44502), .Z(n44500) );
  XOR U44367 ( .A(n44499), .B(n43657), .Z(n44502) );
  XNOR U44368 ( .A(p_input[2125]), .B(n44503), .Z(n43657) );
  AND U44369 ( .A(n795), .B(n44504), .Z(n44503) );
  XOR U44370 ( .A(p_input[2157]), .B(p_input[2125]), .Z(n44504) );
  XNOR U44371 ( .A(n43654), .B(n44499), .Z(n44501) );
  XOR U44372 ( .A(n44505), .B(n44506), .Z(n43654) );
  AND U44373 ( .A(n792), .B(n44507), .Z(n44506) );
  XOR U44374 ( .A(p_input[2093]), .B(p_input[2061]), .Z(n44507) );
  XOR U44375 ( .A(n44508), .B(n44509), .Z(n44499) );
  AND U44376 ( .A(n44510), .B(n44511), .Z(n44509) );
  XOR U44377 ( .A(n44508), .B(n43669), .Z(n44511) );
  XNOR U44378 ( .A(p_input[2124]), .B(n44512), .Z(n43669) );
  AND U44379 ( .A(n795), .B(n44513), .Z(n44512) );
  XOR U44380 ( .A(p_input[2156]), .B(p_input[2124]), .Z(n44513) );
  XNOR U44381 ( .A(n43666), .B(n44508), .Z(n44510) );
  XOR U44382 ( .A(n44514), .B(n44515), .Z(n43666) );
  AND U44383 ( .A(n792), .B(n44516), .Z(n44515) );
  XOR U44384 ( .A(p_input[2092]), .B(p_input[2060]), .Z(n44516) );
  XOR U44385 ( .A(n44517), .B(n44518), .Z(n44508) );
  AND U44386 ( .A(n44519), .B(n44520), .Z(n44518) );
  XOR U44387 ( .A(n44517), .B(n43681), .Z(n44520) );
  XNOR U44388 ( .A(p_input[2123]), .B(n44521), .Z(n43681) );
  AND U44389 ( .A(n795), .B(n44522), .Z(n44521) );
  XOR U44390 ( .A(p_input[2155]), .B(p_input[2123]), .Z(n44522) );
  XNOR U44391 ( .A(n43678), .B(n44517), .Z(n44519) );
  XOR U44392 ( .A(n44523), .B(n44524), .Z(n43678) );
  AND U44393 ( .A(n792), .B(n44525), .Z(n44524) );
  XOR U44394 ( .A(p_input[2091]), .B(p_input[2059]), .Z(n44525) );
  XOR U44395 ( .A(n44526), .B(n44527), .Z(n44517) );
  AND U44396 ( .A(n44528), .B(n44529), .Z(n44527) );
  XOR U44397 ( .A(n44526), .B(n43693), .Z(n44529) );
  XNOR U44398 ( .A(p_input[2122]), .B(n44530), .Z(n43693) );
  AND U44399 ( .A(n795), .B(n44531), .Z(n44530) );
  XOR U44400 ( .A(p_input[2154]), .B(p_input[2122]), .Z(n44531) );
  XNOR U44401 ( .A(n43690), .B(n44526), .Z(n44528) );
  XOR U44402 ( .A(n44532), .B(n44533), .Z(n43690) );
  AND U44403 ( .A(n792), .B(n44534), .Z(n44533) );
  XOR U44404 ( .A(p_input[2090]), .B(p_input[2058]), .Z(n44534) );
  XOR U44405 ( .A(n44535), .B(n44536), .Z(n44526) );
  AND U44406 ( .A(n44537), .B(n44538), .Z(n44536) );
  XOR U44407 ( .A(n44535), .B(n43705), .Z(n44538) );
  XNOR U44408 ( .A(p_input[2121]), .B(n44539), .Z(n43705) );
  AND U44409 ( .A(n795), .B(n44540), .Z(n44539) );
  XOR U44410 ( .A(p_input[2153]), .B(p_input[2121]), .Z(n44540) );
  XNOR U44411 ( .A(n43702), .B(n44535), .Z(n44537) );
  XOR U44412 ( .A(n44541), .B(n44542), .Z(n43702) );
  AND U44413 ( .A(n792), .B(n44543), .Z(n44542) );
  XOR U44414 ( .A(p_input[2089]), .B(p_input[2057]), .Z(n44543) );
  XOR U44415 ( .A(n44544), .B(n44545), .Z(n44535) );
  AND U44416 ( .A(n44546), .B(n44547), .Z(n44545) );
  XOR U44417 ( .A(n44544), .B(n43717), .Z(n44547) );
  XNOR U44418 ( .A(p_input[2120]), .B(n44548), .Z(n43717) );
  AND U44419 ( .A(n795), .B(n44549), .Z(n44548) );
  XOR U44420 ( .A(p_input[2152]), .B(p_input[2120]), .Z(n44549) );
  XNOR U44421 ( .A(n43714), .B(n44544), .Z(n44546) );
  XOR U44422 ( .A(n44550), .B(n44551), .Z(n43714) );
  AND U44423 ( .A(n792), .B(n44552), .Z(n44551) );
  XOR U44424 ( .A(p_input[2088]), .B(p_input[2056]), .Z(n44552) );
  XOR U44425 ( .A(n44553), .B(n44554), .Z(n44544) );
  AND U44426 ( .A(n44555), .B(n44556), .Z(n44554) );
  XOR U44427 ( .A(n44553), .B(n43729), .Z(n44556) );
  XNOR U44428 ( .A(p_input[2119]), .B(n44557), .Z(n43729) );
  AND U44429 ( .A(n795), .B(n44558), .Z(n44557) );
  XOR U44430 ( .A(p_input[2151]), .B(p_input[2119]), .Z(n44558) );
  XNOR U44431 ( .A(n43726), .B(n44553), .Z(n44555) );
  XOR U44432 ( .A(n44559), .B(n44560), .Z(n43726) );
  AND U44433 ( .A(n792), .B(n44561), .Z(n44560) );
  XOR U44434 ( .A(p_input[2087]), .B(p_input[2055]), .Z(n44561) );
  XOR U44435 ( .A(n44562), .B(n44563), .Z(n44553) );
  AND U44436 ( .A(n44564), .B(n44565), .Z(n44563) );
  XOR U44437 ( .A(n44562), .B(n43741), .Z(n44565) );
  XNOR U44438 ( .A(p_input[2118]), .B(n44566), .Z(n43741) );
  AND U44439 ( .A(n795), .B(n44567), .Z(n44566) );
  XOR U44440 ( .A(p_input[2150]), .B(p_input[2118]), .Z(n44567) );
  XNOR U44441 ( .A(n43738), .B(n44562), .Z(n44564) );
  XOR U44442 ( .A(n44568), .B(n44569), .Z(n43738) );
  AND U44443 ( .A(n792), .B(n44570), .Z(n44569) );
  XOR U44444 ( .A(p_input[2086]), .B(p_input[2054]), .Z(n44570) );
  XOR U44445 ( .A(n44571), .B(n44572), .Z(n44562) );
  AND U44446 ( .A(n44573), .B(n44574), .Z(n44572) );
  XOR U44447 ( .A(n44571), .B(n43753), .Z(n44574) );
  XNOR U44448 ( .A(p_input[2117]), .B(n44575), .Z(n43753) );
  AND U44449 ( .A(n795), .B(n44576), .Z(n44575) );
  XOR U44450 ( .A(p_input[2149]), .B(p_input[2117]), .Z(n44576) );
  XNOR U44451 ( .A(n43750), .B(n44571), .Z(n44573) );
  XOR U44452 ( .A(n44577), .B(n44578), .Z(n43750) );
  AND U44453 ( .A(n792), .B(n44579), .Z(n44578) );
  XOR U44454 ( .A(p_input[2085]), .B(p_input[2053]), .Z(n44579) );
  XOR U44455 ( .A(n44580), .B(n44581), .Z(n44571) );
  AND U44456 ( .A(n44582), .B(n44583), .Z(n44581) );
  XOR U44457 ( .A(n44580), .B(n43765), .Z(n44583) );
  XNOR U44458 ( .A(p_input[2116]), .B(n44584), .Z(n43765) );
  AND U44459 ( .A(n795), .B(n44585), .Z(n44584) );
  XOR U44460 ( .A(p_input[2148]), .B(p_input[2116]), .Z(n44585) );
  XNOR U44461 ( .A(n43762), .B(n44580), .Z(n44582) );
  XOR U44462 ( .A(n44586), .B(n44587), .Z(n43762) );
  AND U44463 ( .A(n792), .B(n44588), .Z(n44587) );
  XOR U44464 ( .A(p_input[2084]), .B(p_input[2052]), .Z(n44588) );
  XOR U44465 ( .A(n44589), .B(n44590), .Z(n44580) );
  AND U44466 ( .A(n44591), .B(n44592), .Z(n44590) );
  XOR U44467 ( .A(n44589), .B(n43777), .Z(n44592) );
  XNOR U44468 ( .A(p_input[2115]), .B(n44593), .Z(n43777) );
  AND U44469 ( .A(n795), .B(n44594), .Z(n44593) );
  XOR U44470 ( .A(p_input[2147]), .B(p_input[2115]), .Z(n44594) );
  XNOR U44471 ( .A(n43774), .B(n44589), .Z(n44591) );
  XOR U44472 ( .A(n44595), .B(n44596), .Z(n43774) );
  AND U44473 ( .A(n792), .B(n44597), .Z(n44596) );
  XOR U44474 ( .A(p_input[2083]), .B(p_input[2051]), .Z(n44597) );
  XOR U44475 ( .A(n44598), .B(n44599), .Z(n44589) );
  AND U44476 ( .A(n44600), .B(n44601), .Z(n44599) );
  XOR U44477 ( .A(n44598), .B(n43789), .Z(n44601) );
  XNOR U44478 ( .A(p_input[2114]), .B(n44602), .Z(n43789) );
  AND U44479 ( .A(n795), .B(n44603), .Z(n44602) );
  XOR U44480 ( .A(p_input[2146]), .B(p_input[2114]), .Z(n44603) );
  XNOR U44481 ( .A(n43786), .B(n44598), .Z(n44600) );
  XOR U44482 ( .A(n44604), .B(n44605), .Z(n43786) );
  AND U44483 ( .A(n792), .B(n44606), .Z(n44605) );
  XOR U44484 ( .A(p_input[2082]), .B(p_input[2050]), .Z(n44606) );
  XOR U44485 ( .A(n44607), .B(n44608), .Z(n44598) );
  AND U44486 ( .A(n44609), .B(n44610), .Z(n44608) );
  XNOR U44487 ( .A(n44611), .B(n43802), .Z(n44610) );
  XNOR U44488 ( .A(p_input[2113]), .B(n44612), .Z(n43802) );
  AND U44489 ( .A(n795), .B(n44613), .Z(n44612) );
  XNOR U44490 ( .A(p_input[2145]), .B(n44614), .Z(n44613) );
  IV U44491 ( .A(p_input[2113]), .Z(n44614) );
  XNOR U44492 ( .A(n43799), .B(n44607), .Z(n44609) );
  XNOR U44493 ( .A(p_input[2049]), .B(n44615), .Z(n43799) );
  AND U44494 ( .A(n792), .B(n44616), .Z(n44615) );
  XOR U44495 ( .A(p_input[2081]), .B(p_input[2049]), .Z(n44616) );
  IV U44496 ( .A(n44611), .Z(n44607) );
  AND U44497 ( .A(n44337), .B(n44340), .Z(n44611) );
  XOR U44498 ( .A(p_input[2112]), .B(n44617), .Z(n44340) );
  AND U44499 ( .A(n795), .B(n44618), .Z(n44617) );
  XOR U44500 ( .A(p_input[2144]), .B(p_input[2112]), .Z(n44618) );
  XOR U44501 ( .A(n44619), .B(n44620), .Z(n795) );
  AND U44502 ( .A(n44621), .B(n44622), .Z(n44620) );
  XNOR U44503 ( .A(p_input[2175]), .B(n44619), .Z(n44622) );
  XOR U44504 ( .A(n44619), .B(p_input[2143]), .Z(n44621) );
  XOR U44505 ( .A(n44623), .B(n44624), .Z(n44619) );
  AND U44506 ( .A(n44625), .B(n44626), .Z(n44624) );
  XNOR U44507 ( .A(p_input[2174]), .B(n44623), .Z(n44626) );
  XOR U44508 ( .A(n44623), .B(p_input[2142]), .Z(n44625) );
  XOR U44509 ( .A(n44627), .B(n44628), .Z(n44623) );
  AND U44510 ( .A(n44629), .B(n44630), .Z(n44628) );
  XNOR U44511 ( .A(p_input[2173]), .B(n44627), .Z(n44630) );
  XOR U44512 ( .A(n44627), .B(p_input[2141]), .Z(n44629) );
  XOR U44513 ( .A(n44631), .B(n44632), .Z(n44627) );
  AND U44514 ( .A(n44633), .B(n44634), .Z(n44632) );
  XNOR U44515 ( .A(p_input[2172]), .B(n44631), .Z(n44634) );
  XOR U44516 ( .A(n44631), .B(p_input[2140]), .Z(n44633) );
  XOR U44517 ( .A(n44635), .B(n44636), .Z(n44631) );
  AND U44518 ( .A(n44637), .B(n44638), .Z(n44636) );
  XNOR U44519 ( .A(p_input[2171]), .B(n44635), .Z(n44638) );
  XOR U44520 ( .A(n44635), .B(p_input[2139]), .Z(n44637) );
  XOR U44521 ( .A(n44639), .B(n44640), .Z(n44635) );
  AND U44522 ( .A(n44641), .B(n44642), .Z(n44640) );
  XNOR U44523 ( .A(p_input[2170]), .B(n44639), .Z(n44642) );
  XOR U44524 ( .A(n44639), .B(p_input[2138]), .Z(n44641) );
  XOR U44525 ( .A(n44643), .B(n44644), .Z(n44639) );
  AND U44526 ( .A(n44645), .B(n44646), .Z(n44644) );
  XNOR U44527 ( .A(p_input[2169]), .B(n44643), .Z(n44646) );
  XOR U44528 ( .A(n44643), .B(p_input[2137]), .Z(n44645) );
  XOR U44529 ( .A(n44647), .B(n44648), .Z(n44643) );
  AND U44530 ( .A(n44649), .B(n44650), .Z(n44648) );
  XNOR U44531 ( .A(p_input[2168]), .B(n44647), .Z(n44650) );
  XOR U44532 ( .A(n44647), .B(p_input[2136]), .Z(n44649) );
  XOR U44533 ( .A(n44651), .B(n44652), .Z(n44647) );
  AND U44534 ( .A(n44653), .B(n44654), .Z(n44652) );
  XNOR U44535 ( .A(p_input[2167]), .B(n44651), .Z(n44654) );
  XOR U44536 ( .A(n44651), .B(p_input[2135]), .Z(n44653) );
  XOR U44537 ( .A(n44655), .B(n44656), .Z(n44651) );
  AND U44538 ( .A(n44657), .B(n44658), .Z(n44656) );
  XNOR U44539 ( .A(p_input[2166]), .B(n44655), .Z(n44658) );
  XOR U44540 ( .A(n44655), .B(p_input[2134]), .Z(n44657) );
  XOR U44541 ( .A(n44659), .B(n44660), .Z(n44655) );
  AND U44542 ( .A(n44661), .B(n44662), .Z(n44660) );
  XNOR U44543 ( .A(p_input[2165]), .B(n44659), .Z(n44662) );
  XOR U44544 ( .A(n44659), .B(p_input[2133]), .Z(n44661) );
  XOR U44545 ( .A(n44663), .B(n44664), .Z(n44659) );
  AND U44546 ( .A(n44665), .B(n44666), .Z(n44664) );
  XNOR U44547 ( .A(p_input[2164]), .B(n44663), .Z(n44666) );
  XOR U44548 ( .A(n44663), .B(p_input[2132]), .Z(n44665) );
  XOR U44549 ( .A(n44667), .B(n44668), .Z(n44663) );
  AND U44550 ( .A(n44669), .B(n44670), .Z(n44668) );
  XNOR U44551 ( .A(p_input[2163]), .B(n44667), .Z(n44670) );
  XOR U44552 ( .A(n44667), .B(p_input[2131]), .Z(n44669) );
  XOR U44553 ( .A(n44671), .B(n44672), .Z(n44667) );
  AND U44554 ( .A(n44673), .B(n44674), .Z(n44672) );
  XNOR U44555 ( .A(p_input[2162]), .B(n44671), .Z(n44674) );
  XOR U44556 ( .A(n44671), .B(p_input[2130]), .Z(n44673) );
  XOR U44557 ( .A(n44675), .B(n44676), .Z(n44671) );
  AND U44558 ( .A(n44677), .B(n44678), .Z(n44676) );
  XNOR U44559 ( .A(p_input[2161]), .B(n44675), .Z(n44678) );
  XOR U44560 ( .A(n44675), .B(p_input[2129]), .Z(n44677) );
  XOR U44561 ( .A(n44679), .B(n44680), .Z(n44675) );
  AND U44562 ( .A(n44681), .B(n44682), .Z(n44680) );
  XNOR U44563 ( .A(p_input[2160]), .B(n44679), .Z(n44682) );
  XOR U44564 ( .A(n44679), .B(p_input[2128]), .Z(n44681) );
  XOR U44565 ( .A(n44683), .B(n44684), .Z(n44679) );
  AND U44566 ( .A(n44685), .B(n44686), .Z(n44684) );
  XNOR U44567 ( .A(p_input[2159]), .B(n44683), .Z(n44686) );
  XOR U44568 ( .A(n44683), .B(p_input[2127]), .Z(n44685) );
  XOR U44569 ( .A(n44687), .B(n44688), .Z(n44683) );
  AND U44570 ( .A(n44689), .B(n44690), .Z(n44688) );
  XNOR U44571 ( .A(p_input[2158]), .B(n44687), .Z(n44690) );
  XOR U44572 ( .A(n44687), .B(p_input[2126]), .Z(n44689) );
  XOR U44573 ( .A(n44691), .B(n44692), .Z(n44687) );
  AND U44574 ( .A(n44693), .B(n44694), .Z(n44692) );
  XNOR U44575 ( .A(p_input[2157]), .B(n44691), .Z(n44694) );
  XOR U44576 ( .A(n44691), .B(p_input[2125]), .Z(n44693) );
  XOR U44577 ( .A(n44695), .B(n44696), .Z(n44691) );
  AND U44578 ( .A(n44697), .B(n44698), .Z(n44696) );
  XNOR U44579 ( .A(p_input[2156]), .B(n44695), .Z(n44698) );
  XOR U44580 ( .A(n44695), .B(p_input[2124]), .Z(n44697) );
  XOR U44581 ( .A(n44699), .B(n44700), .Z(n44695) );
  AND U44582 ( .A(n44701), .B(n44702), .Z(n44700) );
  XNOR U44583 ( .A(p_input[2155]), .B(n44699), .Z(n44702) );
  XOR U44584 ( .A(n44699), .B(p_input[2123]), .Z(n44701) );
  XOR U44585 ( .A(n44703), .B(n44704), .Z(n44699) );
  AND U44586 ( .A(n44705), .B(n44706), .Z(n44704) );
  XNOR U44587 ( .A(p_input[2154]), .B(n44703), .Z(n44706) );
  XOR U44588 ( .A(n44703), .B(p_input[2122]), .Z(n44705) );
  XOR U44589 ( .A(n44707), .B(n44708), .Z(n44703) );
  AND U44590 ( .A(n44709), .B(n44710), .Z(n44708) );
  XNOR U44591 ( .A(p_input[2153]), .B(n44707), .Z(n44710) );
  XOR U44592 ( .A(n44707), .B(p_input[2121]), .Z(n44709) );
  XOR U44593 ( .A(n44711), .B(n44712), .Z(n44707) );
  AND U44594 ( .A(n44713), .B(n44714), .Z(n44712) );
  XNOR U44595 ( .A(p_input[2152]), .B(n44711), .Z(n44714) );
  XOR U44596 ( .A(n44711), .B(p_input[2120]), .Z(n44713) );
  XOR U44597 ( .A(n44715), .B(n44716), .Z(n44711) );
  AND U44598 ( .A(n44717), .B(n44718), .Z(n44716) );
  XNOR U44599 ( .A(p_input[2151]), .B(n44715), .Z(n44718) );
  XOR U44600 ( .A(n44715), .B(p_input[2119]), .Z(n44717) );
  XOR U44601 ( .A(n44719), .B(n44720), .Z(n44715) );
  AND U44602 ( .A(n44721), .B(n44722), .Z(n44720) );
  XNOR U44603 ( .A(p_input[2150]), .B(n44719), .Z(n44722) );
  XOR U44604 ( .A(n44719), .B(p_input[2118]), .Z(n44721) );
  XOR U44605 ( .A(n44723), .B(n44724), .Z(n44719) );
  AND U44606 ( .A(n44725), .B(n44726), .Z(n44724) );
  XNOR U44607 ( .A(p_input[2149]), .B(n44723), .Z(n44726) );
  XOR U44608 ( .A(n44723), .B(p_input[2117]), .Z(n44725) );
  XOR U44609 ( .A(n44727), .B(n44728), .Z(n44723) );
  AND U44610 ( .A(n44729), .B(n44730), .Z(n44728) );
  XNOR U44611 ( .A(p_input[2148]), .B(n44727), .Z(n44730) );
  XOR U44612 ( .A(n44727), .B(p_input[2116]), .Z(n44729) );
  XOR U44613 ( .A(n44731), .B(n44732), .Z(n44727) );
  AND U44614 ( .A(n44733), .B(n44734), .Z(n44732) );
  XNOR U44615 ( .A(p_input[2147]), .B(n44731), .Z(n44734) );
  XOR U44616 ( .A(n44731), .B(p_input[2115]), .Z(n44733) );
  XOR U44617 ( .A(n44735), .B(n44736), .Z(n44731) );
  AND U44618 ( .A(n44737), .B(n44738), .Z(n44736) );
  XNOR U44619 ( .A(p_input[2146]), .B(n44735), .Z(n44738) );
  XOR U44620 ( .A(n44735), .B(p_input[2114]), .Z(n44737) );
  XNOR U44621 ( .A(n44739), .B(n44740), .Z(n44735) );
  AND U44622 ( .A(n44741), .B(n44742), .Z(n44740) );
  XOR U44623 ( .A(p_input[2145]), .B(n44739), .Z(n44742) );
  XNOR U44624 ( .A(p_input[2113]), .B(n44739), .Z(n44741) );
  AND U44625 ( .A(p_input[2144]), .B(n44743), .Z(n44739) );
  IV U44626 ( .A(p_input[2112]), .Z(n44743) );
  XNOR U44627 ( .A(p_input[2048]), .B(n44744), .Z(n44337) );
  AND U44628 ( .A(n792), .B(n44745), .Z(n44744) );
  XOR U44629 ( .A(p_input[2080]), .B(p_input[2048]), .Z(n44745) );
  XOR U44630 ( .A(n44746), .B(n44747), .Z(n792) );
  AND U44631 ( .A(n44748), .B(n44749), .Z(n44747) );
  XNOR U44632 ( .A(p_input[2111]), .B(n44746), .Z(n44749) );
  XOR U44633 ( .A(n44746), .B(p_input[2079]), .Z(n44748) );
  XOR U44634 ( .A(n44750), .B(n44751), .Z(n44746) );
  AND U44635 ( .A(n44752), .B(n44753), .Z(n44751) );
  XNOR U44636 ( .A(p_input[2110]), .B(n44750), .Z(n44753) );
  XNOR U44637 ( .A(n44750), .B(n44352), .Z(n44752) );
  IV U44638 ( .A(p_input[2078]), .Z(n44352) );
  XOR U44639 ( .A(n44754), .B(n44755), .Z(n44750) );
  AND U44640 ( .A(n44756), .B(n44757), .Z(n44755) );
  XNOR U44641 ( .A(p_input[2109]), .B(n44754), .Z(n44757) );
  XNOR U44642 ( .A(n44754), .B(n44361), .Z(n44756) );
  IV U44643 ( .A(p_input[2077]), .Z(n44361) );
  XOR U44644 ( .A(n44758), .B(n44759), .Z(n44754) );
  AND U44645 ( .A(n44760), .B(n44761), .Z(n44759) );
  XNOR U44646 ( .A(p_input[2108]), .B(n44758), .Z(n44761) );
  XNOR U44647 ( .A(n44758), .B(n44370), .Z(n44760) );
  IV U44648 ( .A(p_input[2076]), .Z(n44370) );
  XOR U44649 ( .A(n44762), .B(n44763), .Z(n44758) );
  AND U44650 ( .A(n44764), .B(n44765), .Z(n44763) );
  XNOR U44651 ( .A(p_input[2107]), .B(n44762), .Z(n44765) );
  XNOR U44652 ( .A(n44762), .B(n44379), .Z(n44764) );
  IV U44653 ( .A(p_input[2075]), .Z(n44379) );
  XOR U44654 ( .A(n44766), .B(n44767), .Z(n44762) );
  AND U44655 ( .A(n44768), .B(n44769), .Z(n44767) );
  XNOR U44656 ( .A(p_input[2106]), .B(n44766), .Z(n44769) );
  XNOR U44657 ( .A(n44766), .B(n44388), .Z(n44768) );
  IV U44658 ( .A(p_input[2074]), .Z(n44388) );
  XOR U44659 ( .A(n44770), .B(n44771), .Z(n44766) );
  AND U44660 ( .A(n44772), .B(n44773), .Z(n44771) );
  XNOR U44661 ( .A(p_input[2105]), .B(n44770), .Z(n44773) );
  XNOR U44662 ( .A(n44770), .B(n44397), .Z(n44772) );
  IV U44663 ( .A(p_input[2073]), .Z(n44397) );
  XOR U44664 ( .A(n44774), .B(n44775), .Z(n44770) );
  AND U44665 ( .A(n44776), .B(n44777), .Z(n44775) );
  XNOR U44666 ( .A(p_input[2104]), .B(n44774), .Z(n44777) );
  XNOR U44667 ( .A(n44774), .B(n44406), .Z(n44776) );
  IV U44668 ( .A(p_input[2072]), .Z(n44406) );
  XOR U44669 ( .A(n44778), .B(n44779), .Z(n44774) );
  AND U44670 ( .A(n44780), .B(n44781), .Z(n44779) );
  XNOR U44671 ( .A(p_input[2103]), .B(n44778), .Z(n44781) );
  XNOR U44672 ( .A(n44778), .B(n44415), .Z(n44780) );
  IV U44673 ( .A(p_input[2071]), .Z(n44415) );
  XOR U44674 ( .A(n44782), .B(n44783), .Z(n44778) );
  AND U44675 ( .A(n44784), .B(n44785), .Z(n44783) );
  XNOR U44676 ( .A(p_input[2102]), .B(n44782), .Z(n44785) );
  XNOR U44677 ( .A(n44782), .B(n44424), .Z(n44784) );
  IV U44678 ( .A(p_input[2070]), .Z(n44424) );
  XOR U44679 ( .A(n44786), .B(n44787), .Z(n44782) );
  AND U44680 ( .A(n44788), .B(n44789), .Z(n44787) );
  XNOR U44681 ( .A(p_input[2101]), .B(n44786), .Z(n44789) );
  XNOR U44682 ( .A(n44786), .B(n44433), .Z(n44788) );
  IV U44683 ( .A(p_input[2069]), .Z(n44433) );
  XOR U44684 ( .A(n44790), .B(n44791), .Z(n44786) );
  AND U44685 ( .A(n44792), .B(n44793), .Z(n44791) );
  XNOR U44686 ( .A(p_input[2100]), .B(n44790), .Z(n44793) );
  XNOR U44687 ( .A(n44790), .B(n44442), .Z(n44792) );
  IV U44688 ( .A(p_input[2068]), .Z(n44442) );
  XOR U44689 ( .A(n44794), .B(n44795), .Z(n44790) );
  AND U44690 ( .A(n44796), .B(n44797), .Z(n44795) );
  XNOR U44691 ( .A(p_input[2099]), .B(n44794), .Z(n44797) );
  XNOR U44692 ( .A(n44794), .B(n44451), .Z(n44796) );
  IV U44693 ( .A(p_input[2067]), .Z(n44451) );
  XOR U44694 ( .A(n44798), .B(n44799), .Z(n44794) );
  AND U44695 ( .A(n44800), .B(n44801), .Z(n44799) );
  XNOR U44696 ( .A(p_input[2098]), .B(n44798), .Z(n44801) );
  XNOR U44697 ( .A(n44798), .B(n44460), .Z(n44800) );
  IV U44698 ( .A(p_input[2066]), .Z(n44460) );
  XOR U44699 ( .A(n44802), .B(n44803), .Z(n44798) );
  AND U44700 ( .A(n44804), .B(n44805), .Z(n44803) );
  XNOR U44701 ( .A(p_input[2097]), .B(n44802), .Z(n44805) );
  XNOR U44702 ( .A(n44802), .B(n44469), .Z(n44804) );
  IV U44703 ( .A(p_input[2065]), .Z(n44469) );
  XOR U44704 ( .A(n44806), .B(n44807), .Z(n44802) );
  AND U44705 ( .A(n44808), .B(n44809), .Z(n44807) );
  XNOR U44706 ( .A(p_input[2096]), .B(n44806), .Z(n44809) );
  XNOR U44707 ( .A(n44806), .B(n44478), .Z(n44808) );
  IV U44708 ( .A(p_input[2064]), .Z(n44478) );
  XOR U44709 ( .A(n44810), .B(n44811), .Z(n44806) );
  AND U44710 ( .A(n44812), .B(n44813), .Z(n44811) );
  XNOR U44711 ( .A(p_input[2095]), .B(n44810), .Z(n44813) );
  XNOR U44712 ( .A(n44810), .B(n44487), .Z(n44812) );
  IV U44713 ( .A(p_input[2063]), .Z(n44487) );
  XOR U44714 ( .A(n44814), .B(n44815), .Z(n44810) );
  AND U44715 ( .A(n44816), .B(n44817), .Z(n44815) );
  XNOR U44716 ( .A(p_input[2094]), .B(n44814), .Z(n44817) );
  XNOR U44717 ( .A(n44814), .B(n44496), .Z(n44816) );
  IV U44718 ( .A(p_input[2062]), .Z(n44496) );
  XOR U44719 ( .A(n44818), .B(n44819), .Z(n44814) );
  AND U44720 ( .A(n44820), .B(n44821), .Z(n44819) );
  XNOR U44721 ( .A(p_input[2093]), .B(n44818), .Z(n44821) );
  XNOR U44722 ( .A(n44818), .B(n44505), .Z(n44820) );
  IV U44723 ( .A(p_input[2061]), .Z(n44505) );
  XOR U44724 ( .A(n44822), .B(n44823), .Z(n44818) );
  AND U44725 ( .A(n44824), .B(n44825), .Z(n44823) );
  XNOR U44726 ( .A(p_input[2092]), .B(n44822), .Z(n44825) );
  XNOR U44727 ( .A(n44822), .B(n44514), .Z(n44824) );
  IV U44728 ( .A(p_input[2060]), .Z(n44514) );
  XOR U44729 ( .A(n44826), .B(n44827), .Z(n44822) );
  AND U44730 ( .A(n44828), .B(n44829), .Z(n44827) );
  XNOR U44731 ( .A(p_input[2091]), .B(n44826), .Z(n44829) );
  XNOR U44732 ( .A(n44826), .B(n44523), .Z(n44828) );
  IV U44733 ( .A(p_input[2059]), .Z(n44523) );
  XOR U44734 ( .A(n44830), .B(n44831), .Z(n44826) );
  AND U44735 ( .A(n44832), .B(n44833), .Z(n44831) );
  XNOR U44736 ( .A(p_input[2090]), .B(n44830), .Z(n44833) );
  XNOR U44737 ( .A(n44830), .B(n44532), .Z(n44832) );
  IV U44738 ( .A(p_input[2058]), .Z(n44532) );
  XOR U44739 ( .A(n44834), .B(n44835), .Z(n44830) );
  AND U44740 ( .A(n44836), .B(n44837), .Z(n44835) );
  XNOR U44741 ( .A(p_input[2089]), .B(n44834), .Z(n44837) );
  XNOR U44742 ( .A(n44834), .B(n44541), .Z(n44836) );
  IV U44743 ( .A(p_input[2057]), .Z(n44541) );
  XOR U44744 ( .A(n44838), .B(n44839), .Z(n44834) );
  AND U44745 ( .A(n44840), .B(n44841), .Z(n44839) );
  XNOR U44746 ( .A(p_input[2088]), .B(n44838), .Z(n44841) );
  XNOR U44747 ( .A(n44838), .B(n44550), .Z(n44840) );
  IV U44748 ( .A(p_input[2056]), .Z(n44550) );
  XOR U44749 ( .A(n44842), .B(n44843), .Z(n44838) );
  AND U44750 ( .A(n44844), .B(n44845), .Z(n44843) );
  XNOR U44751 ( .A(p_input[2087]), .B(n44842), .Z(n44845) );
  XNOR U44752 ( .A(n44842), .B(n44559), .Z(n44844) );
  IV U44753 ( .A(p_input[2055]), .Z(n44559) );
  XOR U44754 ( .A(n44846), .B(n44847), .Z(n44842) );
  AND U44755 ( .A(n44848), .B(n44849), .Z(n44847) );
  XNOR U44756 ( .A(p_input[2086]), .B(n44846), .Z(n44849) );
  XNOR U44757 ( .A(n44846), .B(n44568), .Z(n44848) );
  IV U44758 ( .A(p_input[2054]), .Z(n44568) );
  XOR U44759 ( .A(n44850), .B(n44851), .Z(n44846) );
  AND U44760 ( .A(n44852), .B(n44853), .Z(n44851) );
  XNOR U44761 ( .A(p_input[2085]), .B(n44850), .Z(n44853) );
  XNOR U44762 ( .A(n44850), .B(n44577), .Z(n44852) );
  IV U44763 ( .A(p_input[2053]), .Z(n44577) );
  XOR U44764 ( .A(n44854), .B(n44855), .Z(n44850) );
  AND U44765 ( .A(n44856), .B(n44857), .Z(n44855) );
  XNOR U44766 ( .A(p_input[2084]), .B(n44854), .Z(n44857) );
  XNOR U44767 ( .A(n44854), .B(n44586), .Z(n44856) );
  IV U44768 ( .A(p_input[2052]), .Z(n44586) );
  XOR U44769 ( .A(n44858), .B(n44859), .Z(n44854) );
  AND U44770 ( .A(n44860), .B(n44861), .Z(n44859) );
  XNOR U44771 ( .A(p_input[2083]), .B(n44858), .Z(n44861) );
  XNOR U44772 ( .A(n44858), .B(n44595), .Z(n44860) );
  IV U44773 ( .A(p_input[2051]), .Z(n44595) );
  XOR U44774 ( .A(n44862), .B(n44863), .Z(n44858) );
  AND U44775 ( .A(n44864), .B(n44865), .Z(n44863) );
  XNOR U44776 ( .A(p_input[2082]), .B(n44862), .Z(n44865) );
  XNOR U44777 ( .A(n44862), .B(n44604), .Z(n44864) );
  IV U44778 ( .A(p_input[2050]), .Z(n44604) );
  XNOR U44779 ( .A(n44866), .B(n44867), .Z(n44862) );
  AND U44780 ( .A(n44868), .B(n44869), .Z(n44867) );
  XOR U44781 ( .A(p_input[2081]), .B(n44866), .Z(n44869) );
  XNOR U44782 ( .A(p_input[2049]), .B(n44866), .Z(n44868) );
  AND U44783 ( .A(p_input[2080]), .B(n44870), .Z(n44866) );
  IV U44784 ( .A(p_input[2048]), .Z(n44870) );
  XOR U44785 ( .A(n44871), .B(n44872), .Z(n30295) );
  AND U44786 ( .A(n1128), .B(n44873), .Z(n44872) );
  XNOR U44787 ( .A(n44874), .B(n44871), .Z(n44873) );
  XOR U44788 ( .A(n44875), .B(n44876), .Z(n1128) );
  AND U44789 ( .A(n44877), .B(n44878), .Z(n44876) );
  XOR U44790 ( .A(n44875), .B(n30310), .Z(n44878) );
  XOR U44791 ( .A(n44879), .B(n44880), .Z(n30310) );
  AND U44792 ( .A(n1103), .B(n44881), .Z(n44880) );
  XOR U44793 ( .A(n44882), .B(n44879), .Z(n44881) );
  XNOR U44794 ( .A(n30307), .B(n44875), .Z(n44877) );
  XOR U44795 ( .A(n44883), .B(n44884), .Z(n30307) );
  AND U44796 ( .A(n1100), .B(n44885), .Z(n44884) );
  XOR U44797 ( .A(n44886), .B(n44883), .Z(n44885) );
  XOR U44798 ( .A(n44887), .B(n44888), .Z(n44875) );
  AND U44799 ( .A(n44889), .B(n44890), .Z(n44888) );
  XOR U44800 ( .A(n44887), .B(n30322), .Z(n44890) );
  XOR U44801 ( .A(n44891), .B(n44892), .Z(n30322) );
  AND U44802 ( .A(n1103), .B(n44893), .Z(n44892) );
  XOR U44803 ( .A(n44894), .B(n44891), .Z(n44893) );
  XNOR U44804 ( .A(n30319), .B(n44887), .Z(n44889) );
  XOR U44805 ( .A(n44895), .B(n44896), .Z(n30319) );
  AND U44806 ( .A(n1100), .B(n44897), .Z(n44896) );
  XOR U44807 ( .A(n44898), .B(n44895), .Z(n44897) );
  XOR U44808 ( .A(n44899), .B(n44900), .Z(n44887) );
  AND U44809 ( .A(n44901), .B(n44902), .Z(n44900) );
  XOR U44810 ( .A(n44899), .B(n30334), .Z(n44902) );
  XOR U44811 ( .A(n44903), .B(n44904), .Z(n30334) );
  AND U44812 ( .A(n1103), .B(n44905), .Z(n44904) );
  XOR U44813 ( .A(n44906), .B(n44903), .Z(n44905) );
  XNOR U44814 ( .A(n30331), .B(n44899), .Z(n44901) );
  XOR U44815 ( .A(n44907), .B(n44908), .Z(n30331) );
  AND U44816 ( .A(n1100), .B(n44909), .Z(n44908) );
  XOR U44817 ( .A(n44910), .B(n44907), .Z(n44909) );
  XOR U44818 ( .A(n44911), .B(n44912), .Z(n44899) );
  AND U44819 ( .A(n44913), .B(n44914), .Z(n44912) );
  XOR U44820 ( .A(n44911), .B(n30346), .Z(n44914) );
  XOR U44821 ( .A(n44915), .B(n44916), .Z(n30346) );
  AND U44822 ( .A(n1103), .B(n44917), .Z(n44916) );
  XOR U44823 ( .A(n44918), .B(n44915), .Z(n44917) );
  XNOR U44824 ( .A(n30343), .B(n44911), .Z(n44913) );
  XOR U44825 ( .A(n44919), .B(n44920), .Z(n30343) );
  AND U44826 ( .A(n1100), .B(n44921), .Z(n44920) );
  XOR U44827 ( .A(n44922), .B(n44919), .Z(n44921) );
  XOR U44828 ( .A(n44923), .B(n44924), .Z(n44911) );
  AND U44829 ( .A(n44925), .B(n44926), .Z(n44924) );
  XOR U44830 ( .A(n44923), .B(n30358), .Z(n44926) );
  XOR U44831 ( .A(n44927), .B(n44928), .Z(n30358) );
  AND U44832 ( .A(n1103), .B(n44929), .Z(n44928) );
  XOR U44833 ( .A(n44930), .B(n44927), .Z(n44929) );
  XNOR U44834 ( .A(n30355), .B(n44923), .Z(n44925) );
  XOR U44835 ( .A(n44931), .B(n44932), .Z(n30355) );
  AND U44836 ( .A(n1100), .B(n44933), .Z(n44932) );
  XOR U44837 ( .A(n44934), .B(n44931), .Z(n44933) );
  XOR U44838 ( .A(n44935), .B(n44936), .Z(n44923) );
  AND U44839 ( .A(n44937), .B(n44938), .Z(n44936) );
  XOR U44840 ( .A(n44935), .B(n30370), .Z(n44938) );
  XOR U44841 ( .A(n44939), .B(n44940), .Z(n30370) );
  AND U44842 ( .A(n1103), .B(n44941), .Z(n44940) );
  XOR U44843 ( .A(n44942), .B(n44939), .Z(n44941) );
  XNOR U44844 ( .A(n30367), .B(n44935), .Z(n44937) );
  XOR U44845 ( .A(n44943), .B(n44944), .Z(n30367) );
  AND U44846 ( .A(n1100), .B(n44945), .Z(n44944) );
  XOR U44847 ( .A(n44946), .B(n44943), .Z(n44945) );
  XOR U44848 ( .A(n44947), .B(n44948), .Z(n44935) );
  AND U44849 ( .A(n44949), .B(n44950), .Z(n44948) );
  XOR U44850 ( .A(n44947), .B(n30382), .Z(n44950) );
  XOR U44851 ( .A(n44951), .B(n44952), .Z(n30382) );
  AND U44852 ( .A(n1103), .B(n44953), .Z(n44952) );
  XOR U44853 ( .A(n44954), .B(n44951), .Z(n44953) );
  XNOR U44854 ( .A(n30379), .B(n44947), .Z(n44949) );
  XOR U44855 ( .A(n44955), .B(n44956), .Z(n30379) );
  AND U44856 ( .A(n1100), .B(n44957), .Z(n44956) );
  XOR U44857 ( .A(n44958), .B(n44955), .Z(n44957) );
  XOR U44858 ( .A(n44959), .B(n44960), .Z(n44947) );
  AND U44859 ( .A(n44961), .B(n44962), .Z(n44960) );
  XOR U44860 ( .A(n44959), .B(n30394), .Z(n44962) );
  XOR U44861 ( .A(n44963), .B(n44964), .Z(n30394) );
  AND U44862 ( .A(n1103), .B(n44965), .Z(n44964) );
  XOR U44863 ( .A(n44966), .B(n44963), .Z(n44965) );
  XNOR U44864 ( .A(n30391), .B(n44959), .Z(n44961) );
  XOR U44865 ( .A(n44967), .B(n44968), .Z(n30391) );
  AND U44866 ( .A(n1100), .B(n44969), .Z(n44968) );
  XOR U44867 ( .A(n44970), .B(n44967), .Z(n44969) );
  XOR U44868 ( .A(n44971), .B(n44972), .Z(n44959) );
  AND U44869 ( .A(n44973), .B(n44974), .Z(n44972) );
  XOR U44870 ( .A(n44971), .B(n30406), .Z(n44974) );
  XOR U44871 ( .A(n44975), .B(n44976), .Z(n30406) );
  AND U44872 ( .A(n1103), .B(n44977), .Z(n44976) );
  XOR U44873 ( .A(n44978), .B(n44975), .Z(n44977) );
  XNOR U44874 ( .A(n30403), .B(n44971), .Z(n44973) );
  XOR U44875 ( .A(n44979), .B(n44980), .Z(n30403) );
  AND U44876 ( .A(n1100), .B(n44981), .Z(n44980) );
  XOR U44877 ( .A(n44982), .B(n44979), .Z(n44981) );
  XOR U44878 ( .A(n44983), .B(n44984), .Z(n44971) );
  AND U44879 ( .A(n44985), .B(n44986), .Z(n44984) );
  XOR U44880 ( .A(n44983), .B(n30418), .Z(n44986) );
  XOR U44881 ( .A(n44987), .B(n44988), .Z(n30418) );
  AND U44882 ( .A(n1103), .B(n44989), .Z(n44988) );
  XOR U44883 ( .A(n44990), .B(n44987), .Z(n44989) );
  XNOR U44884 ( .A(n30415), .B(n44983), .Z(n44985) );
  XOR U44885 ( .A(n44991), .B(n44992), .Z(n30415) );
  AND U44886 ( .A(n1100), .B(n44993), .Z(n44992) );
  XOR U44887 ( .A(n44994), .B(n44991), .Z(n44993) );
  XOR U44888 ( .A(n44995), .B(n44996), .Z(n44983) );
  AND U44889 ( .A(n44997), .B(n44998), .Z(n44996) );
  XOR U44890 ( .A(n44995), .B(n30430), .Z(n44998) );
  XOR U44891 ( .A(n44999), .B(n45000), .Z(n30430) );
  AND U44892 ( .A(n1103), .B(n45001), .Z(n45000) );
  XOR U44893 ( .A(n45002), .B(n44999), .Z(n45001) );
  XNOR U44894 ( .A(n30427), .B(n44995), .Z(n44997) );
  XOR U44895 ( .A(n45003), .B(n45004), .Z(n30427) );
  AND U44896 ( .A(n1100), .B(n45005), .Z(n45004) );
  XOR U44897 ( .A(n45006), .B(n45003), .Z(n45005) );
  XOR U44898 ( .A(n45007), .B(n45008), .Z(n44995) );
  AND U44899 ( .A(n45009), .B(n45010), .Z(n45008) );
  XOR U44900 ( .A(n45007), .B(n30442), .Z(n45010) );
  XOR U44901 ( .A(n45011), .B(n45012), .Z(n30442) );
  AND U44902 ( .A(n1103), .B(n45013), .Z(n45012) );
  XOR U44903 ( .A(n45014), .B(n45011), .Z(n45013) );
  XNOR U44904 ( .A(n30439), .B(n45007), .Z(n45009) );
  XOR U44905 ( .A(n45015), .B(n45016), .Z(n30439) );
  AND U44906 ( .A(n1100), .B(n45017), .Z(n45016) );
  XOR U44907 ( .A(n45018), .B(n45015), .Z(n45017) );
  XOR U44908 ( .A(n45019), .B(n45020), .Z(n45007) );
  AND U44909 ( .A(n45021), .B(n45022), .Z(n45020) );
  XOR U44910 ( .A(n45019), .B(n30454), .Z(n45022) );
  XOR U44911 ( .A(n45023), .B(n45024), .Z(n30454) );
  AND U44912 ( .A(n1103), .B(n45025), .Z(n45024) );
  XOR U44913 ( .A(n45026), .B(n45023), .Z(n45025) );
  XNOR U44914 ( .A(n30451), .B(n45019), .Z(n45021) );
  XOR U44915 ( .A(n45027), .B(n45028), .Z(n30451) );
  AND U44916 ( .A(n1100), .B(n45029), .Z(n45028) );
  XOR U44917 ( .A(n45030), .B(n45027), .Z(n45029) );
  XOR U44918 ( .A(n45031), .B(n45032), .Z(n45019) );
  AND U44919 ( .A(n45033), .B(n45034), .Z(n45032) );
  XOR U44920 ( .A(n45031), .B(n30466), .Z(n45034) );
  XOR U44921 ( .A(n45035), .B(n45036), .Z(n30466) );
  AND U44922 ( .A(n1103), .B(n45037), .Z(n45036) );
  XOR U44923 ( .A(n45038), .B(n45035), .Z(n45037) );
  XNOR U44924 ( .A(n30463), .B(n45031), .Z(n45033) );
  XOR U44925 ( .A(n45039), .B(n45040), .Z(n30463) );
  AND U44926 ( .A(n1100), .B(n45041), .Z(n45040) );
  XOR U44927 ( .A(n45042), .B(n45039), .Z(n45041) );
  XOR U44928 ( .A(n45043), .B(n45044), .Z(n45031) );
  AND U44929 ( .A(n45045), .B(n45046), .Z(n45044) );
  XOR U44930 ( .A(n45043), .B(n30478), .Z(n45046) );
  XOR U44931 ( .A(n45047), .B(n45048), .Z(n30478) );
  AND U44932 ( .A(n1103), .B(n45049), .Z(n45048) );
  XOR U44933 ( .A(n45050), .B(n45047), .Z(n45049) );
  XNOR U44934 ( .A(n30475), .B(n45043), .Z(n45045) );
  XOR U44935 ( .A(n45051), .B(n45052), .Z(n30475) );
  AND U44936 ( .A(n1100), .B(n45053), .Z(n45052) );
  XOR U44937 ( .A(n45054), .B(n45051), .Z(n45053) );
  XOR U44938 ( .A(n45055), .B(n45056), .Z(n45043) );
  AND U44939 ( .A(n45057), .B(n45058), .Z(n45056) );
  XOR U44940 ( .A(n45055), .B(n30490), .Z(n45058) );
  XOR U44941 ( .A(n45059), .B(n45060), .Z(n30490) );
  AND U44942 ( .A(n1103), .B(n45061), .Z(n45060) );
  XOR U44943 ( .A(n45062), .B(n45059), .Z(n45061) );
  XNOR U44944 ( .A(n30487), .B(n45055), .Z(n45057) );
  XOR U44945 ( .A(n45063), .B(n45064), .Z(n30487) );
  AND U44946 ( .A(n1100), .B(n45065), .Z(n45064) );
  XOR U44947 ( .A(n45066), .B(n45063), .Z(n45065) );
  XOR U44948 ( .A(n45067), .B(n45068), .Z(n45055) );
  AND U44949 ( .A(n45069), .B(n45070), .Z(n45068) );
  XOR U44950 ( .A(n45067), .B(n30502), .Z(n45070) );
  XOR U44951 ( .A(n45071), .B(n45072), .Z(n30502) );
  AND U44952 ( .A(n1103), .B(n45073), .Z(n45072) );
  XOR U44953 ( .A(n45074), .B(n45071), .Z(n45073) );
  XNOR U44954 ( .A(n30499), .B(n45067), .Z(n45069) );
  XOR U44955 ( .A(n45075), .B(n45076), .Z(n30499) );
  AND U44956 ( .A(n1100), .B(n45077), .Z(n45076) );
  XOR U44957 ( .A(n45078), .B(n45075), .Z(n45077) );
  XOR U44958 ( .A(n45079), .B(n45080), .Z(n45067) );
  AND U44959 ( .A(n45081), .B(n45082), .Z(n45080) );
  XOR U44960 ( .A(n45079), .B(n30514), .Z(n45082) );
  XOR U44961 ( .A(n45083), .B(n45084), .Z(n30514) );
  AND U44962 ( .A(n1103), .B(n45085), .Z(n45084) );
  XOR U44963 ( .A(n45086), .B(n45083), .Z(n45085) );
  XNOR U44964 ( .A(n30511), .B(n45079), .Z(n45081) );
  XOR U44965 ( .A(n45087), .B(n45088), .Z(n30511) );
  AND U44966 ( .A(n1100), .B(n45089), .Z(n45088) );
  XOR U44967 ( .A(n45090), .B(n45087), .Z(n45089) );
  XOR U44968 ( .A(n45091), .B(n45092), .Z(n45079) );
  AND U44969 ( .A(n45093), .B(n45094), .Z(n45092) );
  XOR U44970 ( .A(n45091), .B(n30526), .Z(n45094) );
  XOR U44971 ( .A(n45095), .B(n45096), .Z(n30526) );
  AND U44972 ( .A(n1103), .B(n45097), .Z(n45096) );
  XOR U44973 ( .A(n45098), .B(n45095), .Z(n45097) );
  XNOR U44974 ( .A(n30523), .B(n45091), .Z(n45093) );
  XOR U44975 ( .A(n45099), .B(n45100), .Z(n30523) );
  AND U44976 ( .A(n1100), .B(n45101), .Z(n45100) );
  XOR U44977 ( .A(n45102), .B(n45099), .Z(n45101) );
  XOR U44978 ( .A(n45103), .B(n45104), .Z(n45091) );
  AND U44979 ( .A(n45105), .B(n45106), .Z(n45104) );
  XOR U44980 ( .A(n45103), .B(n30538), .Z(n45106) );
  XOR U44981 ( .A(n45107), .B(n45108), .Z(n30538) );
  AND U44982 ( .A(n1103), .B(n45109), .Z(n45108) );
  XOR U44983 ( .A(n45110), .B(n45107), .Z(n45109) );
  XNOR U44984 ( .A(n30535), .B(n45103), .Z(n45105) );
  XOR U44985 ( .A(n45111), .B(n45112), .Z(n30535) );
  AND U44986 ( .A(n1100), .B(n45113), .Z(n45112) );
  XOR U44987 ( .A(n45114), .B(n45111), .Z(n45113) );
  XOR U44988 ( .A(n45115), .B(n45116), .Z(n45103) );
  AND U44989 ( .A(n45117), .B(n45118), .Z(n45116) );
  XOR U44990 ( .A(n45115), .B(n30550), .Z(n45118) );
  XOR U44991 ( .A(n45119), .B(n45120), .Z(n30550) );
  AND U44992 ( .A(n1103), .B(n45121), .Z(n45120) );
  XOR U44993 ( .A(n45122), .B(n45119), .Z(n45121) );
  XNOR U44994 ( .A(n30547), .B(n45115), .Z(n45117) );
  XOR U44995 ( .A(n45123), .B(n45124), .Z(n30547) );
  AND U44996 ( .A(n1100), .B(n45125), .Z(n45124) );
  XOR U44997 ( .A(n45126), .B(n45123), .Z(n45125) );
  XOR U44998 ( .A(n45127), .B(n45128), .Z(n45115) );
  AND U44999 ( .A(n45129), .B(n45130), .Z(n45128) );
  XOR U45000 ( .A(n45127), .B(n30562), .Z(n45130) );
  XOR U45001 ( .A(n45131), .B(n45132), .Z(n30562) );
  AND U45002 ( .A(n1103), .B(n45133), .Z(n45132) );
  XOR U45003 ( .A(n45134), .B(n45131), .Z(n45133) );
  XNOR U45004 ( .A(n30559), .B(n45127), .Z(n45129) );
  XOR U45005 ( .A(n45135), .B(n45136), .Z(n30559) );
  AND U45006 ( .A(n1100), .B(n45137), .Z(n45136) );
  XOR U45007 ( .A(n45138), .B(n45135), .Z(n45137) );
  XOR U45008 ( .A(n45139), .B(n45140), .Z(n45127) );
  AND U45009 ( .A(n45141), .B(n45142), .Z(n45140) );
  XOR U45010 ( .A(n45139), .B(n30574), .Z(n45142) );
  XOR U45011 ( .A(n45143), .B(n45144), .Z(n30574) );
  AND U45012 ( .A(n1103), .B(n45145), .Z(n45144) );
  XOR U45013 ( .A(n45146), .B(n45143), .Z(n45145) );
  XNOR U45014 ( .A(n30571), .B(n45139), .Z(n45141) );
  XOR U45015 ( .A(n45147), .B(n45148), .Z(n30571) );
  AND U45016 ( .A(n1100), .B(n45149), .Z(n45148) );
  XOR U45017 ( .A(n45150), .B(n45147), .Z(n45149) );
  XOR U45018 ( .A(n45151), .B(n45152), .Z(n45139) );
  AND U45019 ( .A(n45153), .B(n45154), .Z(n45152) );
  XOR U45020 ( .A(n45151), .B(n30586), .Z(n45154) );
  XOR U45021 ( .A(n45155), .B(n45156), .Z(n30586) );
  AND U45022 ( .A(n1103), .B(n45157), .Z(n45156) );
  XOR U45023 ( .A(n45158), .B(n45155), .Z(n45157) );
  XNOR U45024 ( .A(n30583), .B(n45151), .Z(n45153) );
  XOR U45025 ( .A(n45159), .B(n45160), .Z(n30583) );
  AND U45026 ( .A(n1100), .B(n45161), .Z(n45160) );
  XOR U45027 ( .A(n45162), .B(n45159), .Z(n45161) );
  XOR U45028 ( .A(n45163), .B(n45164), .Z(n45151) );
  AND U45029 ( .A(n45165), .B(n45166), .Z(n45164) );
  XOR U45030 ( .A(n45163), .B(n30598), .Z(n45166) );
  XOR U45031 ( .A(n45167), .B(n45168), .Z(n30598) );
  AND U45032 ( .A(n1103), .B(n45169), .Z(n45168) );
  XOR U45033 ( .A(n45170), .B(n45167), .Z(n45169) );
  XNOR U45034 ( .A(n30595), .B(n45163), .Z(n45165) );
  XOR U45035 ( .A(n45171), .B(n45172), .Z(n30595) );
  AND U45036 ( .A(n1100), .B(n45173), .Z(n45172) );
  XOR U45037 ( .A(n45174), .B(n45171), .Z(n45173) );
  XOR U45038 ( .A(n45175), .B(n45176), .Z(n45163) );
  AND U45039 ( .A(n45177), .B(n45178), .Z(n45176) );
  XOR U45040 ( .A(n45175), .B(n30610), .Z(n45178) );
  XOR U45041 ( .A(n45179), .B(n45180), .Z(n30610) );
  AND U45042 ( .A(n1103), .B(n45181), .Z(n45180) );
  XOR U45043 ( .A(n45182), .B(n45179), .Z(n45181) );
  XNOR U45044 ( .A(n30607), .B(n45175), .Z(n45177) );
  XOR U45045 ( .A(n45183), .B(n45184), .Z(n30607) );
  AND U45046 ( .A(n1100), .B(n45185), .Z(n45184) );
  XOR U45047 ( .A(n45186), .B(n45183), .Z(n45185) );
  XOR U45048 ( .A(n45187), .B(n45188), .Z(n45175) );
  AND U45049 ( .A(n45189), .B(n45190), .Z(n45188) );
  XOR U45050 ( .A(n45187), .B(n30622), .Z(n45190) );
  XOR U45051 ( .A(n45191), .B(n45192), .Z(n30622) );
  AND U45052 ( .A(n1103), .B(n45193), .Z(n45192) );
  XOR U45053 ( .A(n45194), .B(n45191), .Z(n45193) );
  XNOR U45054 ( .A(n30619), .B(n45187), .Z(n45189) );
  XOR U45055 ( .A(n45195), .B(n45196), .Z(n30619) );
  AND U45056 ( .A(n1100), .B(n45197), .Z(n45196) );
  XOR U45057 ( .A(n45198), .B(n45195), .Z(n45197) );
  XOR U45058 ( .A(n45199), .B(n45200), .Z(n45187) );
  AND U45059 ( .A(n45201), .B(n45202), .Z(n45200) );
  XOR U45060 ( .A(n45199), .B(n30634), .Z(n45202) );
  XOR U45061 ( .A(n45203), .B(n45204), .Z(n30634) );
  AND U45062 ( .A(n1103), .B(n45205), .Z(n45204) );
  XOR U45063 ( .A(n45206), .B(n45203), .Z(n45205) );
  XNOR U45064 ( .A(n30631), .B(n45199), .Z(n45201) );
  XOR U45065 ( .A(n45207), .B(n45208), .Z(n30631) );
  AND U45066 ( .A(n1100), .B(n45209), .Z(n45208) );
  XOR U45067 ( .A(n45210), .B(n45207), .Z(n45209) );
  XOR U45068 ( .A(n45211), .B(n45212), .Z(n45199) );
  AND U45069 ( .A(n45213), .B(n45214), .Z(n45212) );
  XOR U45070 ( .A(n45211), .B(n30646), .Z(n45214) );
  XOR U45071 ( .A(n45215), .B(n45216), .Z(n30646) );
  AND U45072 ( .A(n1103), .B(n45217), .Z(n45216) );
  XOR U45073 ( .A(n45218), .B(n45215), .Z(n45217) );
  XNOR U45074 ( .A(n30643), .B(n45211), .Z(n45213) );
  XOR U45075 ( .A(n45219), .B(n45220), .Z(n30643) );
  AND U45076 ( .A(n1100), .B(n45221), .Z(n45220) );
  XOR U45077 ( .A(n45222), .B(n45219), .Z(n45221) );
  XOR U45078 ( .A(n45223), .B(n45224), .Z(n45211) );
  AND U45079 ( .A(n45225), .B(n45226), .Z(n45224) );
  XOR U45080 ( .A(n45223), .B(n30658), .Z(n45226) );
  XOR U45081 ( .A(n45227), .B(n45228), .Z(n30658) );
  AND U45082 ( .A(n1103), .B(n45229), .Z(n45228) );
  XOR U45083 ( .A(n45230), .B(n45227), .Z(n45229) );
  XNOR U45084 ( .A(n30655), .B(n45223), .Z(n45225) );
  XOR U45085 ( .A(n45231), .B(n45232), .Z(n30655) );
  AND U45086 ( .A(n1100), .B(n45233), .Z(n45232) );
  XOR U45087 ( .A(n45234), .B(n45231), .Z(n45233) );
  XOR U45088 ( .A(n45235), .B(n45236), .Z(n45223) );
  AND U45089 ( .A(n45237), .B(n45238), .Z(n45236) );
  XNOR U45090 ( .A(n45239), .B(n30671), .Z(n45238) );
  XOR U45091 ( .A(n45240), .B(n45241), .Z(n30671) );
  AND U45092 ( .A(n1103), .B(n45242), .Z(n45241) );
  XOR U45093 ( .A(n45240), .B(n45243), .Z(n45242) );
  XNOR U45094 ( .A(n30668), .B(n45235), .Z(n45237) );
  XOR U45095 ( .A(n45244), .B(n45245), .Z(n30668) );
  AND U45096 ( .A(n1100), .B(n45246), .Z(n45245) );
  XOR U45097 ( .A(n45244), .B(n45247), .Z(n45246) );
  IV U45098 ( .A(n45239), .Z(n45235) );
  AND U45099 ( .A(n44871), .B(n44874), .Z(n45239) );
  XNOR U45100 ( .A(n45248), .B(n45249), .Z(n44874) );
  AND U45101 ( .A(n1103), .B(n45250), .Z(n45249) );
  XNOR U45102 ( .A(n45251), .B(n45248), .Z(n45250) );
  XOR U45103 ( .A(n45252), .B(n45253), .Z(n1103) );
  AND U45104 ( .A(n45254), .B(n45255), .Z(n45253) );
  XOR U45105 ( .A(n45252), .B(n44882), .Z(n45255) );
  XOR U45106 ( .A(n45256), .B(n45257), .Z(n44882) );
  AND U45107 ( .A(n1039), .B(n45258), .Z(n45257) );
  XOR U45108 ( .A(n45259), .B(n45256), .Z(n45258) );
  XNOR U45109 ( .A(n44879), .B(n45252), .Z(n45254) );
  XOR U45110 ( .A(n45260), .B(n45261), .Z(n44879) );
  AND U45111 ( .A(n1037), .B(n45262), .Z(n45261) );
  XOR U45112 ( .A(n45263), .B(n45260), .Z(n45262) );
  XOR U45113 ( .A(n45264), .B(n45265), .Z(n45252) );
  AND U45114 ( .A(n45266), .B(n45267), .Z(n45265) );
  XOR U45115 ( .A(n45264), .B(n44894), .Z(n45267) );
  XOR U45116 ( .A(n45268), .B(n45269), .Z(n44894) );
  AND U45117 ( .A(n1039), .B(n45270), .Z(n45269) );
  XOR U45118 ( .A(n45271), .B(n45268), .Z(n45270) );
  XNOR U45119 ( .A(n44891), .B(n45264), .Z(n45266) );
  XOR U45120 ( .A(n45272), .B(n45273), .Z(n44891) );
  AND U45121 ( .A(n1037), .B(n45274), .Z(n45273) );
  XOR U45122 ( .A(n45275), .B(n45272), .Z(n45274) );
  XOR U45123 ( .A(n45276), .B(n45277), .Z(n45264) );
  AND U45124 ( .A(n45278), .B(n45279), .Z(n45277) );
  XOR U45125 ( .A(n45276), .B(n44906), .Z(n45279) );
  XOR U45126 ( .A(n45280), .B(n45281), .Z(n44906) );
  AND U45127 ( .A(n1039), .B(n45282), .Z(n45281) );
  XOR U45128 ( .A(n45283), .B(n45280), .Z(n45282) );
  XNOR U45129 ( .A(n44903), .B(n45276), .Z(n45278) );
  XOR U45130 ( .A(n45284), .B(n45285), .Z(n44903) );
  AND U45131 ( .A(n1037), .B(n45286), .Z(n45285) );
  XOR U45132 ( .A(n45287), .B(n45284), .Z(n45286) );
  XOR U45133 ( .A(n45288), .B(n45289), .Z(n45276) );
  AND U45134 ( .A(n45290), .B(n45291), .Z(n45289) );
  XOR U45135 ( .A(n45288), .B(n44918), .Z(n45291) );
  XOR U45136 ( .A(n45292), .B(n45293), .Z(n44918) );
  AND U45137 ( .A(n1039), .B(n45294), .Z(n45293) );
  XOR U45138 ( .A(n45295), .B(n45292), .Z(n45294) );
  XNOR U45139 ( .A(n44915), .B(n45288), .Z(n45290) );
  XOR U45140 ( .A(n45296), .B(n45297), .Z(n44915) );
  AND U45141 ( .A(n1037), .B(n45298), .Z(n45297) );
  XOR U45142 ( .A(n45299), .B(n45296), .Z(n45298) );
  XOR U45143 ( .A(n45300), .B(n45301), .Z(n45288) );
  AND U45144 ( .A(n45302), .B(n45303), .Z(n45301) );
  XOR U45145 ( .A(n45300), .B(n44930), .Z(n45303) );
  XOR U45146 ( .A(n45304), .B(n45305), .Z(n44930) );
  AND U45147 ( .A(n1039), .B(n45306), .Z(n45305) );
  XOR U45148 ( .A(n45307), .B(n45304), .Z(n45306) );
  XNOR U45149 ( .A(n44927), .B(n45300), .Z(n45302) );
  XOR U45150 ( .A(n45308), .B(n45309), .Z(n44927) );
  AND U45151 ( .A(n1037), .B(n45310), .Z(n45309) );
  XOR U45152 ( .A(n45311), .B(n45308), .Z(n45310) );
  XOR U45153 ( .A(n45312), .B(n45313), .Z(n45300) );
  AND U45154 ( .A(n45314), .B(n45315), .Z(n45313) );
  XOR U45155 ( .A(n45312), .B(n44942), .Z(n45315) );
  XOR U45156 ( .A(n45316), .B(n45317), .Z(n44942) );
  AND U45157 ( .A(n1039), .B(n45318), .Z(n45317) );
  XOR U45158 ( .A(n45319), .B(n45316), .Z(n45318) );
  XNOR U45159 ( .A(n44939), .B(n45312), .Z(n45314) );
  XOR U45160 ( .A(n45320), .B(n45321), .Z(n44939) );
  AND U45161 ( .A(n1037), .B(n45322), .Z(n45321) );
  XOR U45162 ( .A(n45323), .B(n45320), .Z(n45322) );
  XOR U45163 ( .A(n45324), .B(n45325), .Z(n45312) );
  AND U45164 ( .A(n45326), .B(n45327), .Z(n45325) );
  XOR U45165 ( .A(n45324), .B(n44954), .Z(n45327) );
  XOR U45166 ( .A(n45328), .B(n45329), .Z(n44954) );
  AND U45167 ( .A(n1039), .B(n45330), .Z(n45329) );
  XOR U45168 ( .A(n45331), .B(n45328), .Z(n45330) );
  XNOR U45169 ( .A(n44951), .B(n45324), .Z(n45326) );
  XOR U45170 ( .A(n45332), .B(n45333), .Z(n44951) );
  AND U45171 ( .A(n1037), .B(n45334), .Z(n45333) );
  XOR U45172 ( .A(n45335), .B(n45332), .Z(n45334) );
  XOR U45173 ( .A(n45336), .B(n45337), .Z(n45324) );
  AND U45174 ( .A(n45338), .B(n45339), .Z(n45337) );
  XOR U45175 ( .A(n45336), .B(n44966), .Z(n45339) );
  XOR U45176 ( .A(n45340), .B(n45341), .Z(n44966) );
  AND U45177 ( .A(n1039), .B(n45342), .Z(n45341) );
  XOR U45178 ( .A(n45343), .B(n45340), .Z(n45342) );
  XNOR U45179 ( .A(n44963), .B(n45336), .Z(n45338) );
  XOR U45180 ( .A(n45344), .B(n45345), .Z(n44963) );
  AND U45181 ( .A(n1037), .B(n45346), .Z(n45345) );
  XOR U45182 ( .A(n45347), .B(n45344), .Z(n45346) );
  XOR U45183 ( .A(n45348), .B(n45349), .Z(n45336) );
  AND U45184 ( .A(n45350), .B(n45351), .Z(n45349) );
  XOR U45185 ( .A(n45348), .B(n44978), .Z(n45351) );
  XOR U45186 ( .A(n45352), .B(n45353), .Z(n44978) );
  AND U45187 ( .A(n1039), .B(n45354), .Z(n45353) );
  XOR U45188 ( .A(n45355), .B(n45352), .Z(n45354) );
  XNOR U45189 ( .A(n44975), .B(n45348), .Z(n45350) );
  XOR U45190 ( .A(n45356), .B(n45357), .Z(n44975) );
  AND U45191 ( .A(n1037), .B(n45358), .Z(n45357) );
  XOR U45192 ( .A(n45359), .B(n45356), .Z(n45358) );
  XOR U45193 ( .A(n45360), .B(n45361), .Z(n45348) );
  AND U45194 ( .A(n45362), .B(n45363), .Z(n45361) );
  XOR U45195 ( .A(n45360), .B(n44990), .Z(n45363) );
  XOR U45196 ( .A(n45364), .B(n45365), .Z(n44990) );
  AND U45197 ( .A(n1039), .B(n45366), .Z(n45365) );
  XOR U45198 ( .A(n45367), .B(n45364), .Z(n45366) );
  XNOR U45199 ( .A(n44987), .B(n45360), .Z(n45362) );
  XOR U45200 ( .A(n45368), .B(n45369), .Z(n44987) );
  AND U45201 ( .A(n1037), .B(n45370), .Z(n45369) );
  XOR U45202 ( .A(n45371), .B(n45368), .Z(n45370) );
  XOR U45203 ( .A(n45372), .B(n45373), .Z(n45360) );
  AND U45204 ( .A(n45374), .B(n45375), .Z(n45373) );
  XOR U45205 ( .A(n45372), .B(n45002), .Z(n45375) );
  XOR U45206 ( .A(n45376), .B(n45377), .Z(n45002) );
  AND U45207 ( .A(n1039), .B(n45378), .Z(n45377) );
  XOR U45208 ( .A(n45379), .B(n45376), .Z(n45378) );
  XNOR U45209 ( .A(n44999), .B(n45372), .Z(n45374) );
  XOR U45210 ( .A(n45380), .B(n45381), .Z(n44999) );
  AND U45211 ( .A(n1037), .B(n45382), .Z(n45381) );
  XOR U45212 ( .A(n45383), .B(n45380), .Z(n45382) );
  XOR U45213 ( .A(n45384), .B(n45385), .Z(n45372) );
  AND U45214 ( .A(n45386), .B(n45387), .Z(n45385) );
  XOR U45215 ( .A(n45384), .B(n45014), .Z(n45387) );
  XOR U45216 ( .A(n45388), .B(n45389), .Z(n45014) );
  AND U45217 ( .A(n1039), .B(n45390), .Z(n45389) );
  XOR U45218 ( .A(n45391), .B(n45388), .Z(n45390) );
  XNOR U45219 ( .A(n45011), .B(n45384), .Z(n45386) );
  XOR U45220 ( .A(n45392), .B(n45393), .Z(n45011) );
  AND U45221 ( .A(n1037), .B(n45394), .Z(n45393) );
  XOR U45222 ( .A(n45395), .B(n45392), .Z(n45394) );
  XOR U45223 ( .A(n45396), .B(n45397), .Z(n45384) );
  AND U45224 ( .A(n45398), .B(n45399), .Z(n45397) );
  XOR U45225 ( .A(n45396), .B(n45026), .Z(n45399) );
  XOR U45226 ( .A(n45400), .B(n45401), .Z(n45026) );
  AND U45227 ( .A(n1039), .B(n45402), .Z(n45401) );
  XOR U45228 ( .A(n45403), .B(n45400), .Z(n45402) );
  XNOR U45229 ( .A(n45023), .B(n45396), .Z(n45398) );
  XOR U45230 ( .A(n45404), .B(n45405), .Z(n45023) );
  AND U45231 ( .A(n1037), .B(n45406), .Z(n45405) );
  XOR U45232 ( .A(n45407), .B(n45404), .Z(n45406) );
  XOR U45233 ( .A(n45408), .B(n45409), .Z(n45396) );
  AND U45234 ( .A(n45410), .B(n45411), .Z(n45409) );
  XOR U45235 ( .A(n45408), .B(n45038), .Z(n45411) );
  XOR U45236 ( .A(n45412), .B(n45413), .Z(n45038) );
  AND U45237 ( .A(n1039), .B(n45414), .Z(n45413) );
  XOR U45238 ( .A(n45415), .B(n45412), .Z(n45414) );
  XNOR U45239 ( .A(n45035), .B(n45408), .Z(n45410) );
  XOR U45240 ( .A(n45416), .B(n45417), .Z(n45035) );
  AND U45241 ( .A(n1037), .B(n45418), .Z(n45417) );
  XOR U45242 ( .A(n45419), .B(n45416), .Z(n45418) );
  XOR U45243 ( .A(n45420), .B(n45421), .Z(n45408) );
  AND U45244 ( .A(n45422), .B(n45423), .Z(n45421) );
  XOR U45245 ( .A(n45420), .B(n45050), .Z(n45423) );
  XOR U45246 ( .A(n45424), .B(n45425), .Z(n45050) );
  AND U45247 ( .A(n1039), .B(n45426), .Z(n45425) );
  XOR U45248 ( .A(n45427), .B(n45424), .Z(n45426) );
  XNOR U45249 ( .A(n45047), .B(n45420), .Z(n45422) );
  XOR U45250 ( .A(n45428), .B(n45429), .Z(n45047) );
  AND U45251 ( .A(n1037), .B(n45430), .Z(n45429) );
  XOR U45252 ( .A(n45431), .B(n45428), .Z(n45430) );
  XOR U45253 ( .A(n45432), .B(n45433), .Z(n45420) );
  AND U45254 ( .A(n45434), .B(n45435), .Z(n45433) );
  XOR U45255 ( .A(n45432), .B(n45062), .Z(n45435) );
  XOR U45256 ( .A(n45436), .B(n45437), .Z(n45062) );
  AND U45257 ( .A(n1039), .B(n45438), .Z(n45437) );
  XOR U45258 ( .A(n45439), .B(n45436), .Z(n45438) );
  XNOR U45259 ( .A(n45059), .B(n45432), .Z(n45434) );
  XOR U45260 ( .A(n45440), .B(n45441), .Z(n45059) );
  AND U45261 ( .A(n1037), .B(n45442), .Z(n45441) );
  XOR U45262 ( .A(n45443), .B(n45440), .Z(n45442) );
  XOR U45263 ( .A(n45444), .B(n45445), .Z(n45432) );
  AND U45264 ( .A(n45446), .B(n45447), .Z(n45445) );
  XOR U45265 ( .A(n45444), .B(n45074), .Z(n45447) );
  XOR U45266 ( .A(n45448), .B(n45449), .Z(n45074) );
  AND U45267 ( .A(n1039), .B(n45450), .Z(n45449) );
  XOR U45268 ( .A(n45451), .B(n45448), .Z(n45450) );
  XNOR U45269 ( .A(n45071), .B(n45444), .Z(n45446) );
  XOR U45270 ( .A(n45452), .B(n45453), .Z(n45071) );
  AND U45271 ( .A(n1037), .B(n45454), .Z(n45453) );
  XOR U45272 ( .A(n45455), .B(n45452), .Z(n45454) );
  XOR U45273 ( .A(n45456), .B(n45457), .Z(n45444) );
  AND U45274 ( .A(n45458), .B(n45459), .Z(n45457) );
  XOR U45275 ( .A(n45456), .B(n45086), .Z(n45459) );
  XOR U45276 ( .A(n45460), .B(n45461), .Z(n45086) );
  AND U45277 ( .A(n1039), .B(n45462), .Z(n45461) );
  XOR U45278 ( .A(n45463), .B(n45460), .Z(n45462) );
  XNOR U45279 ( .A(n45083), .B(n45456), .Z(n45458) );
  XOR U45280 ( .A(n45464), .B(n45465), .Z(n45083) );
  AND U45281 ( .A(n1037), .B(n45466), .Z(n45465) );
  XOR U45282 ( .A(n45467), .B(n45464), .Z(n45466) );
  XOR U45283 ( .A(n45468), .B(n45469), .Z(n45456) );
  AND U45284 ( .A(n45470), .B(n45471), .Z(n45469) );
  XOR U45285 ( .A(n45468), .B(n45098), .Z(n45471) );
  XOR U45286 ( .A(n45472), .B(n45473), .Z(n45098) );
  AND U45287 ( .A(n1039), .B(n45474), .Z(n45473) );
  XOR U45288 ( .A(n45475), .B(n45472), .Z(n45474) );
  XNOR U45289 ( .A(n45095), .B(n45468), .Z(n45470) );
  XOR U45290 ( .A(n45476), .B(n45477), .Z(n45095) );
  AND U45291 ( .A(n1037), .B(n45478), .Z(n45477) );
  XOR U45292 ( .A(n45479), .B(n45476), .Z(n45478) );
  XOR U45293 ( .A(n45480), .B(n45481), .Z(n45468) );
  AND U45294 ( .A(n45482), .B(n45483), .Z(n45481) );
  XOR U45295 ( .A(n45480), .B(n45110), .Z(n45483) );
  XOR U45296 ( .A(n45484), .B(n45485), .Z(n45110) );
  AND U45297 ( .A(n1039), .B(n45486), .Z(n45485) );
  XOR U45298 ( .A(n45487), .B(n45484), .Z(n45486) );
  XNOR U45299 ( .A(n45107), .B(n45480), .Z(n45482) );
  XOR U45300 ( .A(n45488), .B(n45489), .Z(n45107) );
  AND U45301 ( .A(n1037), .B(n45490), .Z(n45489) );
  XOR U45302 ( .A(n45491), .B(n45488), .Z(n45490) );
  XOR U45303 ( .A(n45492), .B(n45493), .Z(n45480) );
  AND U45304 ( .A(n45494), .B(n45495), .Z(n45493) );
  XOR U45305 ( .A(n45492), .B(n45122), .Z(n45495) );
  XOR U45306 ( .A(n45496), .B(n45497), .Z(n45122) );
  AND U45307 ( .A(n1039), .B(n45498), .Z(n45497) );
  XOR U45308 ( .A(n45499), .B(n45496), .Z(n45498) );
  XNOR U45309 ( .A(n45119), .B(n45492), .Z(n45494) );
  XOR U45310 ( .A(n45500), .B(n45501), .Z(n45119) );
  AND U45311 ( .A(n1037), .B(n45502), .Z(n45501) );
  XOR U45312 ( .A(n45503), .B(n45500), .Z(n45502) );
  XOR U45313 ( .A(n45504), .B(n45505), .Z(n45492) );
  AND U45314 ( .A(n45506), .B(n45507), .Z(n45505) );
  XOR U45315 ( .A(n45504), .B(n45134), .Z(n45507) );
  XOR U45316 ( .A(n45508), .B(n45509), .Z(n45134) );
  AND U45317 ( .A(n1039), .B(n45510), .Z(n45509) );
  XOR U45318 ( .A(n45511), .B(n45508), .Z(n45510) );
  XNOR U45319 ( .A(n45131), .B(n45504), .Z(n45506) );
  XOR U45320 ( .A(n45512), .B(n45513), .Z(n45131) );
  AND U45321 ( .A(n1037), .B(n45514), .Z(n45513) );
  XOR U45322 ( .A(n45515), .B(n45512), .Z(n45514) );
  XOR U45323 ( .A(n45516), .B(n45517), .Z(n45504) );
  AND U45324 ( .A(n45518), .B(n45519), .Z(n45517) );
  XOR U45325 ( .A(n45516), .B(n45146), .Z(n45519) );
  XOR U45326 ( .A(n45520), .B(n45521), .Z(n45146) );
  AND U45327 ( .A(n1039), .B(n45522), .Z(n45521) );
  XOR U45328 ( .A(n45523), .B(n45520), .Z(n45522) );
  XNOR U45329 ( .A(n45143), .B(n45516), .Z(n45518) );
  XOR U45330 ( .A(n45524), .B(n45525), .Z(n45143) );
  AND U45331 ( .A(n1037), .B(n45526), .Z(n45525) );
  XOR U45332 ( .A(n45527), .B(n45524), .Z(n45526) );
  XOR U45333 ( .A(n45528), .B(n45529), .Z(n45516) );
  AND U45334 ( .A(n45530), .B(n45531), .Z(n45529) );
  XOR U45335 ( .A(n45528), .B(n45158), .Z(n45531) );
  XOR U45336 ( .A(n45532), .B(n45533), .Z(n45158) );
  AND U45337 ( .A(n1039), .B(n45534), .Z(n45533) );
  XOR U45338 ( .A(n45535), .B(n45532), .Z(n45534) );
  XNOR U45339 ( .A(n45155), .B(n45528), .Z(n45530) );
  XOR U45340 ( .A(n45536), .B(n45537), .Z(n45155) );
  AND U45341 ( .A(n1037), .B(n45538), .Z(n45537) );
  XOR U45342 ( .A(n45539), .B(n45536), .Z(n45538) );
  XOR U45343 ( .A(n45540), .B(n45541), .Z(n45528) );
  AND U45344 ( .A(n45542), .B(n45543), .Z(n45541) );
  XOR U45345 ( .A(n45540), .B(n45170), .Z(n45543) );
  XOR U45346 ( .A(n45544), .B(n45545), .Z(n45170) );
  AND U45347 ( .A(n1039), .B(n45546), .Z(n45545) );
  XOR U45348 ( .A(n45547), .B(n45544), .Z(n45546) );
  XNOR U45349 ( .A(n45167), .B(n45540), .Z(n45542) );
  XOR U45350 ( .A(n45548), .B(n45549), .Z(n45167) );
  AND U45351 ( .A(n1037), .B(n45550), .Z(n45549) );
  XOR U45352 ( .A(n45551), .B(n45548), .Z(n45550) );
  XOR U45353 ( .A(n45552), .B(n45553), .Z(n45540) );
  AND U45354 ( .A(n45554), .B(n45555), .Z(n45553) );
  XOR U45355 ( .A(n45552), .B(n45182), .Z(n45555) );
  XOR U45356 ( .A(n45556), .B(n45557), .Z(n45182) );
  AND U45357 ( .A(n1039), .B(n45558), .Z(n45557) );
  XOR U45358 ( .A(n45559), .B(n45556), .Z(n45558) );
  XNOR U45359 ( .A(n45179), .B(n45552), .Z(n45554) );
  XOR U45360 ( .A(n45560), .B(n45561), .Z(n45179) );
  AND U45361 ( .A(n1037), .B(n45562), .Z(n45561) );
  XOR U45362 ( .A(n45563), .B(n45560), .Z(n45562) );
  XOR U45363 ( .A(n45564), .B(n45565), .Z(n45552) );
  AND U45364 ( .A(n45566), .B(n45567), .Z(n45565) );
  XOR U45365 ( .A(n45564), .B(n45194), .Z(n45567) );
  XOR U45366 ( .A(n45568), .B(n45569), .Z(n45194) );
  AND U45367 ( .A(n1039), .B(n45570), .Z(n45569) );
  XOR U45368 ( .A(n45571), .B(n45568), .Z(n45570) );
  XNOR U45369 ( .A(n45191), .B(n45564), .Z(n45566) );
  XOR U45370 ( .A(n45572), .B(n45573), .Z(n45191) );
  AND U45371 ( .A(n1037), .B(n45574), .Z(n45573) );
  XOR U45372 ( .A(n45575), .B(n45572), .Z(n45574) );
  XOR U45373 ( .A(n45576), .B(n45577), .Z(n45564) );
  AND U45374 ( .A(n45578), .B(n45579), .Z(n45577) );
  XOR U45375 ( .A(n45576), .B(n45206), .Z(n45579) );
  XOR U45376 ( .A(n45580), .B(n45581), .Z(n45206) );
  AND U45377 ( .A(n1039), .B(n45582), .Z(n45581) );
  XOR U45378 ( .A(n45583), .B(n45580), .Z(n45582) );
  XNOR U45379 ( .A(n45203), .B(n45576), .Z(n45578) );
  XOR U45380 ( .A(n45584), .B(n45585), .Z(n45203) );
  AND U45381 ( .A(n1037), .B(n45586), .Z(n45585) );
  XOR U45382 ( .A(n45587), .B(n45584), .Z(n45586) );
  XOR U45383 ( .A(n45588), .B(n45589), .Z(n45576) );
  AND U45384 ( .A(n45590), .B(n45591), .Z(n45589) );
  XOR U45385 ( .A(n45588), .B(n45218), .Z(n45591) );
  XOR U45386 ( .A(n45592), .B(n45593), .Z(n45218) );
  AND U45387 ( .A(n1039), .B(n45594), .Z(n45593) );
  XOR U45388 ( .A(n45595), .B(n45592), .Z(n45594) );
  XNOR U45389 ( .A(n45215), .B(n45588), .Z(n45590) );
  XOR U45390 ( .A(n45596), .B(n45597), .Z(n45215) );
  AND U45391 ( .A(n1037), .B(n45598), .Z(n45597) );
  XOR U45392 ( .A(n45599), .B(n45596), .Z(n45598) );
  XOR U45393 ( .A(n45600), .B(n45601), .Z(n45588) );
  AND U45394 ( .A(n45602), .B(n45603), .Z(n45601) );
  XOR U45395 ( .A(n45600), .B(n45230), .Z(n45603) );
  XOR U45396 ( .A(n45604), .B(n45605), .Z(n45230) );
  AND U45397 ( .A(n1039), .B(n45606), .Z(n45605) );
  XOR U45398 ( .A(n45607), .B(n45604), .Z(n45606) );
  XNOR U45399 ( .A(n45227), .B(n45600), .Z(n45602) );
  XOR U45400 ( .A(n45608), .B(n45609), .Z(n45227) );
  AND U45401 ( .A(n1037), .B(n45610), .Z(n45609) );
  XOR U45402 ( .A(n45611), .B(n45608), .Z(n45610) );
  XOR U45403 ( .A(n45612), .B(n45613), .Z(n45600) );
  AND U45404 ( .A(n45614), .B(n45615), .Z(n45613) );
  XNOR U45405 ( .A(n45616), .B(n45243), .Z(n45615) );
  XOR U45406 ( .A(n45617), .B(n45618), .Z(n45243) );
  AND U45407 ( .A(n1039), .B(n45619), .Z(n45618) );
  XOR U45408 ( .A(n45617), .B(n45620), .Z(n45619) );
  XNOR U45409 ( .A(n45240), .B(n45612), .Z(n45614) );
  XOR U45410 ( .A(n45621), .B(n45622), .Z(n45240) );
  AND U45411 ( .A(n1037), .B(n45623), .Z(n45622) );
  XOR U45412 ( .A(n45621), .B(n45624), .Z(n45623) );
  IV U45413 ( .A(n45616), .Z(n45612) );
  AND U45414 ( .A(n45248), .B(n45251), .Z(n45616) );
  XNOR U45415 ( .A(n45625), .B(n45626), .Z(n45251) );
  AND U45416 ( .A(n1039), .B(n45627), .Z(n45626) );
  XNOR U45417 ( .A(n45628), .B(n45625), .Z(n45627) );
  XOR U45418 ( .A(n45629), .B(n45630), .Z(n1039) );
  AND U45419 ( .A(n45631), .B(n45632), .Z(n45630) );
  XOR U45420 ( .A(n45629), .B(n45259), .Z(n45632) );
  XOR U45421 ( .A(n45633), .B(n45634), .Z(n45259) );
  AND U45422 ( .A(n903), .B(n45635), .Z(n45634) );
  XOR U45423 ( .A(n45636), .B(n45633), .Z(n45635) );
  XNOR U45424 ( .A(n45256), .B(n45629), .Z(n45631) );
  XOR U45425 ( .A(n45637), .B(n45638), .Z(n45256) );
  AND U45426 ( .A(n901), .B(n45639), .Z(n45638) );
  XOR U45427 ( .A(n45640), .B(n45637), .Z(n45639) );
  XOR U45428 ( .A(n45641), .B(n45642), .Z(n45629) );
  AND U45429 ( .A(n45643), .B(n45644), .Z(n45642) );
  XOR U45430 ( .A(n45641), .B(n45271), .Z(n45644) );
  XOR U45431 ( .A(n45645), .B(n45646), .Z(n45271) );
  AND U45432 ( .A(n903), .B(n45647), .Z(n45646) );
  XOR U45433 ( .A(n45648), .B(n45645), .Z(n45647) );
  XNOR U45434 ( .A(n45268), .B(n45641), .Z(n45643) );
  XOR U45435 ( .A(n45649), .B(n45650), .Z(n45268) );
  AND U45436 ( .A(n901), .B(n45651), .Z(n45650) );
  XOR U45437 ( .A(n45652), .B(n45649), .Z(n45651) );
  XOR U45438 ( .A(n45653), .B(n45654), .Z(n45641) );
  AND U45439 ( .A(n45655), .B(n45656), .Z(n45654) );
  XOR U45440 ( .A(n45653), .B(n45283), .Z(n45656) );
  XOR U45441 ( .A(n45657), .B(n45658), .Z(n45283) );
  AND U45442 ( .A(n903), .B(n45659), .Z(n45658) );
  XOR U45443 ( .A(n45660), .B(n45657), .Z(n45659) );
  XNOR U45444 ( .A(n45280), .B(n45653), .Z(n45655) );
  XOR U45445 ( .A(n45661), .B(n45662), .Z(n45280) );
  AND U45446 ( .A(n901), .B(n45663), .Z(n45662) );
  XOR U45447 ( .A(n45664), .B(n45661), .Z(n45663) );
  XOR U45448 ( .A(n45665), .B(n45666), .Z(n45653) );
  AND U45449 ( .A(n45667), .B(n45668), .Z(n45666) );
  XOR U45450 ( .A(n45665), .B(n45295), .Z(n45668) );
  XOR U45451 ( .A(n45669), .B(n45670), .Z(n45295) );
  AND U45452 ( .A(n903), .B(n45671), .Z(n45670) );
  XOR U45453 ( .A(n45672), .B(n45669), .Z(n45671) );
  XNOR U45454 ( .A(n45292), .B(n45665), .Z(n45667) );
  XOR U45455 ( .A(n45673), .B(n45674), .Z(n45292) );
  AND U45456 ( .A(n901), .B(n45675), .Z(n45674) );
  XOR U45457 ( .A(n45676), .B(n45673), .Z(n45675) );
  XOR U45458 ( .A(n45677), .B(n45678), .Z(n45665) );
  AND U45459 ( .A(n45679), .B(n45680), .Z(n45678) );
  XOR U45460 ( .A(n45677), .B(n45307), .Z(n45680) );
  XOR U45461 ( .A(n45681), .B(n45682), .Z(n45307) );
  AND U45462 ( .A(n903), .B(n45683), .Z(n45682) );
  XOR U45463 ( .A(n45684), .B(n45681), .Z(n45683) );
  XNOR U45464 ( .A(n45304), .B(n45677), .Z(n45679) );
  XOR U45465 ( .A(n45685), .B(n45686), .Z(n45304) );
  AND U45466 ( .A(n901), .B(n45687), .Z(n45686) );
  XOR U45467 ( .A(n45688), .B(n45685), .Z(n45687) );
  XOR U45468 ( .A(n45689), .B(n45690), .Z(n45677) );
  AND U45469 ( .A(n45691), .B(n45692), .Z(n45690) );
  XOR U45470 ( .A(n45689), .B(n45319), .Z(n45692) );
  XOR U45471 ( .A(n45693), .B(n45694), .Z(n45319) );
  AND U45472 ( .A(n903), .B(n45695), .Z(n45694) );
  XOR U45473 ( .A(n45696), .B(n45693), .Z(n45695) );
  XNOR U45474 ( .A(n45316), .B(n45689), .Z(n45691) );
  XOR U45475 ( .A(n45697), .B(n45698), .Z(n45316) );
  AND U45476 ( .A(n901), .B(n45699), .Z(n45698) );
  XOR U45477 ( .A(n45700), .B(n45697), .Z(n45699) );
  XOR U45478 ( .A(n45701), .B(n45702), .Z(n45689) );
  AND U45479 ( .A(n45703), .B(n45704), .Z(n45702) );
  XOR U45480 ( .A(n45701), .B(n45331), .Z(n45704) );
  XOR U45481 ( .A(n45705), .B(n45706), .Z(n45331) );
  AND U45482 ( .A(n903), .B(n45707), .Z(n45706) );
  XOR U45483 ( .A(n45708), .B(n45705), .Z(n45707) );
  XNOR U45484 ( .A(n45328), .B(n45701), .Z(n45703) );
  XOR U45485 ( .A(n45709), .B(n45710), .Z(n45328) );
  AND U45486 ( .A(n901), .B(n45711), .Z(n45710) );
  XOR U45487 ( .A(n45712), .B(n45709), .Z(n45711) );
  XOR U45488 ( .A(n45713), .B(n45714), .Z(n45701) );
  AND U45489 ( .A(n45715), .B(n45716), .Z(n45714) );
  XOR U45490 ( .A(n45713), .B(n45343), .Z(n45716) );
  XOR U45491 ( .A(n45717), .B(n45718), .Z(n45343) );
  AND U45492 ( .A(n903), .B(n45719), .Z(n45718) );
  XOR U45493 ( .A(n45720), .B(n45717), .Z(n45719) );
  XNOR U45494 ( .A(n45340), .B(n45713), .Z(n45715) );
  XOR U45495 ( .A(n45721), .B(n45722), .Z(n45340) );
  AND U45496 ( .A(n901), .B(n45723), .Z(n45722) );
  XOR U45497 ( .A(n45724), .B(n45721), .Z(n45723) );
  XOR U45498 ( .A(n45725), .B(n45726), .Z(n45713) );
  AND U45499 ( .A(n45727), .B(n45728), .Z(n45726) );
  XOR U45500 ( .A(n45725), .B(n45355), .Z(n45728) );
  XOR U45501 ( .A(n45729), .B(n45730), .Z(n45355) );
  AND U45502 ( .A(n903), .B(n45731), .Z(n45730) );
  XOR U45503 ( .A(n45732), .B(n45729), .Z(n45731) );
  XNOR U45504 ( .A(n45352), .B(n45725), .Z(n45727) );
  XOR U45505 ( .A(n45733), .B(n45734), .Z(n45352) );
  AND U45506 ( .A(n901), .B(n45735), .Z(n45734) );
  XOR U45507 ( .A(n45736), .B(n45733), .Z(n45735) );
  XOR U45508 ( .A(n45737), .B(n45738), .Z(n45725) );
  AND U45509 ( .A(n45739), .B(n45740), .Z(n45738) );
  XOR U45510 ( .A(n45737), .B(n45367), .Z(n45740) );
  XOR U45511 ( .A(n45741), .B(n45742), .Z(n45367) );
  AND U45512 ( .A(n903), .B(n45743), .Z(n45742) );
  XOR U45513 ( .A(n45744), .B(n45741), .Z(n45743) );
  XNOR U45514 ( .A(n45364), .B(n45737), .Z(n45739) );
  XOR U45515 ( .A(n45745), .B(n45746), .Z(n45364) );
  AND U45516 ( .A(n901), .B(n45747), .Z(n45746) );
  XOR U45517 ( .A(n45748), .B(n45745), .Z(n45747) );
  XOR U45518 ( .A(n45749), .B(n45750), .Z(n45737) );
  AND U45519 ( .A(n45751), .B(n45752), .Z(n45750) );
  XOR U45520 ( .A(n45749), .B(n45379), .Z(n45752) );
  XOR U45521 ( .A(n45753), .B(n45754), .Z(n45379) );
  AND U45522 ( .A(n903), .B(n45755), .Z(n45754) );
  XOR U45523 ( .A(n45756), .B(n45753), .Z(n45755) );
  XNOR U45524 ( .A(n45376), .B(n45749), .Z(n45751) );
  XOR U45525 ( .A(n45757), .B(n45758), .Z(n45376) );
  AND U45526 ( .A(n901), .B(n45759), .Z(n45758) );
  XOR U45527 ( .A(n45760), .B(n45757), .Z(n45759) );
  XOR U45528 ( .A(n45761), .B(n45762), .Z(n45749) );
  AND U45529 ( .A(n45763), .B(n45764), .Z(n45762) );
  XOR U45530 ( .A(n45761), .B(n45391), .Z(n45764) );
  XOR U45531 ( .A(n45765), .B(n45766), .Z(n45391) );
  AND U45532 ( .A(n903), .B(n45767), .Z(n45766) );
  XOR U45533 ( .A(n45768), .B(n45765), .Z(n45767) );
  XNOR U45534 ( .A(n45388), .B(n45761), .Z(n45763) );
  XOR U45535 ( .A(n45769), .B(n45770), .Z(n45388) );
  AND U45536 ( .A(n901), .B(n45771), .Z(n45770) );
  XOR U45537 ( .A(n45772), .B(n45769), .Z(n45771) );
  XOR U45538 ( .A(n45773), .B(n45774), .Z(n45761) );
  AND U45539 ( .A(n45775), .B(n45776), .Z(n45774) );
  XOR U45540 ( .A(n45773), .B(n45403), .Z(n45776) );
  XOR U45541 ( .A(n45777), .B(n45778), .Z(n45403) );
  AND U45542 ( .A(n903), .B(n45779), .Z(n45778) );
  XOR U45543 ( .A(n45780), .B(n45777), .Z(n45779) );
  XNOR U45544 ( .A(n45400), .B(n45773), .Z(n45775) );
  XOR U45545 ( .A(n45781), .B(n45782), .Z(n45400) );
  AND U45546 ( .A(n901), .B(n45783), .Z(n45782) );
  XOR U45547 ( .A(n45784), .B(n45781), .Z(n45783) );
  XOR U45548 ( .A(n45785), .B(n45786), .Z(n45773) );
  AND U45549 ( .A(n45787), .B(n45788), .Z(n45786) );
  XOR U45550 ( .A(n45785), .B(n45415), .Z(n45788) );
  XOR U45551 ( .A(n45789), .B(n45790), .Z(n45415) );
  AND U45552 ( .A(n903), .B(n45791), .Z(n45790) );
  XOR U45553 ( .A(n45792), .B(n45789), .Z(n45791) );
  XNOR U45554 ( .A(n45412), .B(n45785), .Z(n45787) );
  XOR U45555 ( .A(n45793), .B(n45794), .Z(n45412) );
  AND U45556 ( .A(n901), .B(n45795), .Z(n45794) );
  XOR U45557 ( .A(n45796), .B(n45793), .Z(n45795) );
  XOR U45558 ( .A(n45797), .B(n45798), .Z(n45785) );
  AND U45559 ( .A(n45799), .B(n45800), .Z(n45798) );
  XOR U45560 ( .A(n45797), .B(n45427), .Z(n45800) );
  XOR U45561 ( .A(n45801), .B(n45802), .Z(n45427) );
  AND U45562 ( .A(n903), .B(n45803), .Z(n45802) );
  XOR U45563 ( .A(n45804), .B(n45801), .Z(n45803) );
  XNOR U45564 ( .A(n45424), .B(n45797), .Z(n45799) );
  XOR U45565 ( .A(n45805), .B(n45806), .Z(n45424) );
  AND U45566 ( .A(n901), .B(n45807), .Z(n45806) );
  XOR U45567 ( .A(n45808), .B(n45805), .Z(n45807) );
  XOR U45568 ( .A(n45809), .B(n45810), .Z(n45797) );
  AND U45569 ( .A(n45811), .B(n45812), .Z(n45810) );
  XOR U45570 ( .A(n45809), .B(n45439), .Z(n45812) );
  XOR U45571 ( .A(n45813), .B(n45814), .Z(n45439) );
  AND U45572 ( .A(n903), .B(n45815), .Z(n45814) );
  XOR U45573 ( .A(n45816), .B(n45813), .Z(n45815) );
  XNOR U45574 ( .A(n45436), .B(n45809), .Z(n45811) );
  XOR U45575 ( .A(n45817), .B(n45818), .Z(n45436) );
  AND U45576 ( .A(n901), .B(n45819), .Z(n45818) );
  XOR U45577 ( .A(n45820), .B(n45817), .Z(n45819) );
  XOR U45578 ( .A(n45821), .B(n45822), .Z(n45809) );
  AND U45579 ( .A(n45823), .B(n45824), .Z(n45822) );
  XOR U45580 ( .A(n45821), .B(n45451), .Z(n45824) );
  XOR U45581 ( .A(n45825), .B(n45826), .Z(n45451) );
  AND U45582 ( .A(n903), .B(n45827), .Z(n45826) );
  XOR U45583 ( .A(n45828), .B(n45825), .Z(n45827) );
  XNOR U45584 ( .A(n45448), .B(n45821), .Z(n45823) );
  XOR U45585 ( .A(n45829), .B(n45830), .Z(n45448) );
  AND U45586 ( .A(n901), .B(n45831), .Z(n45830) );
  XOR U45587 ( .A(n45832), .B(n45829), .Z(n45831) );
  XOR U45588 ( .A(n45833), .B(n45834), .Z(n45821) );
  AND U45589 ( .A(n45835), .B(n45836), .Z(n45834) );
  XOR U45590 ( .A(n45833), .B(n45463), .Z(n45836) );
  XOR U45591 ( .A(n45837), .B(n45838), .Z(n45463) );
  AND U45592 ( .A(n903), .B(n45839), .Z(n45838) );
  XOR U45593 ( .A(n45840), .B(n45837), .Z(n45839) );
  XNOR U45594 ( .A(n45460), .B(n45833), .Z(n45835) );
  XOR U45595 ( .A(n45841), .B(n45842), .Z(n45460) );
  AND U45596 ( .A(n901), .B(n45843), .Z(n45842) );
  XOR U45597 ( .A(n45844), .B(n45841), .Z(n45843) );
  XOR U45598 ( .A(n45845), .B(n45846), .Z(n45833) );
  AND U45599 ( .A(n45847), .B(n45848), .Z(n45846) );
  XOR U45600 ( .A(n45845), .B(n45475), .Z(n45848) );
  XOR U45601 ( .A(n45849), .B(n45850), .Z(n45475) );
  AND U45602 ( .A(n903), .B(n45851), .Z(n45850) );
  XOR U45603 ( .A(n45852), .B(n45849), .Z(n45851) );
  XNOR U45604 ( .A(n45472), .B(n45845), .Z(n45847) );
  XOR U45605 ( .A(n45853), .B(n45854), .Z(n45472) );
  AND U45606 ( .A(n901), .B(n45855), .Z(n45854) );
  XOR U45607 ( .A(n45856), .B(n45853), .Z(n45855) );
  XOR U45608 ( .A(n45857), .B(n45858), .Z(n45845) );
  AND U45609 ( .A(n45859), .B(n45860), .Z(n45858) );
  XOR U45610 ( .A(n45857), .B(n45487), .Z(n45860) );
  XOR U45611 ( .A(n45861), .B(n45862), .Z(n45487) );
  AND U45612 ( .A(n903), .B(n45863), .Z(n45862) );
  XOR U45613 ( .A(n45864), .B(n45861), .Z(n45863) );
  XNOR U45614 ( .A(n45484), .B(n45857), .Z(n45859) );
  XOR U45615 ( .A(n45865), .B(n45866), .Z(n45484) );
  AND U45616 ( .A(n901), .B(n45867), .Z(n45866) );
  XOR U45617 ( .A(n45868), .B(n45865), .Z(n45867) );
  XOR U45618 ( .A(n45869), .B(n45870), .Z(n45857) );
  AND U45619 ( .A(n45871), .B(n45872), .Z(n45870) );
  XOR U45620 ( .A(n45869), .B(n45499), .Z(n45872) );
  XOR U45621 ( .A(n45873), .B(n45874), .Z(n45499) );
  AND U45622 ( .A(n903), .B(n45875), .Z(n45874) );
  XOR U45623 ( .A(n45876), .B(n45873), .Z(n45875) );
  XNOR U45624 ( .A(n45496), .B(n45869), .Z(n45871) );
  XOR U45625 ( .A(n45877), .B(n45878), .Z(n45496) );
  AND U45626 ( .A(n901), .B(n45879), .Z(n45878) );
  XOR U45627 ( .A(n45880), .B(n45877), .Z(n45879) );
  XOR U45628 ( .A(n45881), .B(n45882), .Z(n45869) );
  AND U45629 ( .A(n45883), .B(n45884), .Z(n45882) );
  XOR U45630 ( .A(n45881), .B(n45511), .Z(n45884) );
  XOR U45631 ( .A(n45885), .B(n45886), .Z(n45511) );
  AND U45632 ( .A(n903), .B(n45887), .Z(n45886) );
  XOR U45633 ( .A(n45888), .B(n45885), .Z(n45887) );
  XNOR U45634 ( .A(n45508), .B(n45881), .Z(n45883) );
  XOR U45635 ( .A(n45889), .B(n45890), .Z(n45508) );
  AND U45636 ( .A(n901), .B(n45891), .Z(n45890) );
  XOR U45637 ( .A(n45892), .B(n45889), .Z(n45891) );
  XOR U45638 ( .A(n45893), .B(n45894), .Z(n45881) );
  AND U45639 ( .A(n45895), .B(n45896), .Z(n45894) );
  XOR U45640 ( .A(n45893), .B(n45523), .Z(n45896) );
  XOR U45641 ( .A(n45897), .B(n45898), .Z(n45523) );
  AND U45642 ( .A(n903), .B(n45899), .Z(n45898) );
  XOR U45643 ( .A(n45900), .B(n45897), .Z(n45899) );
  XNOR U45644 ( .A(n45520), .B(n45893), .Z(n45895) );
  XOR U45645 ( .A(n45901), .B(n45902), .Z(n45520) );
  AND U45646 ( .A(n901), .B(n45903), .Z(n45902) );
  XOR U45647 ( .A(n45904), .B(n45901), .Z(n45903) );
  XOR U45648 ( .A(n45905), .B(n45906), .Z(n45893) );
  AND U45649 ( .A(n45907), .B(n45908), .Z(n45906) );
  XOR U45650 ( .A(n45905), .B(n45535), .Z(n45908) );
  XOR U45651 ( .A(n45909), .B(n45910), .Z(n45535) );
  AND U45652 ( .A(n903), .B(n45911), .Z(n45910) );
  XOR U45653 ( .A(n45912), .B(n45909), .Z(n45911) );
  XNOR U45654 ( .A(n45532), .B(n45905), .Z(n45907) );
  XOR U45655 ( .A(n45913), .B(n45914), .Z(n45532) );
  AND U45656 ( .A(n901), .B(n45915), .Z(n45914) );
  XOR U45657 ( .A(n45916), .B(n45913), .Z(n45915) );
  XOR U45658 ( .A(n45917), .B(n45918), .Z(n45905) );
  AND U45659 ( .A(n45919), .B(n45920), .Z(n45918) );
  XOR U45660 ( .A(n45917), .B(n45547), .Z(n45920) );
  XOR U45661 ( .A(n45921), .B(n45922), .Z(n45547) );
  AND U45662 ( .A(n903), .B(n45923), .Z(n45922) );
  XOR U45663 ( .A(n45924), .B(n45921), .Z(n45923) );
  XNOR U45664 ( .A(n45544), .B(n45917), .Z(n45919) );
  XOR U45665 ( .A(n45925), .B(n45926), .Z(n45544) );
  AND U45666 ( .A(n901), .B(n45927), .Z(n45926) );
  XOR U45667 ( .A(n45928), .B(n45925), .Z(n45927) );
  XOR U45668 ( .A(n45929), .B(n45930), .Z(n45917) );
  AND U45669 ( .A(n45931), .B(n45932), .Z(n45930) );
  XOR U45670 ( .A(n45929), .B(n45559), .Z(n45932) );
  XOR U45671 ( .A(n45933), .B(n45934), .Z(n45559) );
  AND U45672 ( .A(n903), .B(n45935), .Z(n45934) );
  XOR U45673 ( .A(n45936), .B(n45933), .Z(n45935) );
  XNOR U45674 ( .A(n45556), .B(n45929), .Z(n45931) );
  XOR U45675 ( .A(n45937), .B(n45938), .Z(n45556) );
  AND U45676 ( .A(n901), .B(n45939), .Z(n45938) );
  XOR U45677 ( .A(n45940), .B(n45937), .Z(n45939) );
  XOR U45678 ( .A(n45941), .B(n45942), .Z(n45929) );
  AND U45679 ( .A(n45943), .B(n45944), .Z(n45942) );
  XOR U45680 ( .A(n45941), .B(n45571), .Z(n45944) );
  XOR U45681 ( .A(n45945), .B(n45946), .Z(n45571) );
  AND U45682 ( .A(n903), .B(n45947), .Z(n45946) );
  XOR U45683 ( .A(n45948), .B(n45945), .Z(n45947) );
  XNOR U45684 ( .A(n45568), .B(n45941), .Z(n45943) );
  XOR U45685 ( .A(n45949), .B(n45950), .Z(n45568) );
  AND U45686 ( .A(n901), .B(n45951), .Z(n45950) );
  XOR U45687 ( .A(n45952), .B(n45949), .Z(n45951) );
  XOR U45688 ( .A(n45953), .B(n45954), .Z(n45941) );
  AND U45689 ( .A(n45955), .B(n45956), .Z(n45954) );
  XOR U45690 ( .A(n45953), .B(n45583), .Z(n45956) );
  XOR U45691 ( .A(n45957), .B(n45958), .Z(n45583) );
  AND U45692 ( .A(n903), .B(n45959), .Z(n45958) );
  XOR U45693 ( .A(n45960), .B(n45957), .Z(n45959) );
  XNOR U45694 ( .A(n45580), .B(n45953), .Z(n45955) );
  XOR U45695 ( .A(n45961), .B(n45962), .Z(n45580) );
  AND U45696 ( .A(n901), .B(n45963), .Z(n45962) );
  XOR U45697 ( .A(n45964), .B(n45961), .Z(n45963) );
  XOR U45698 ( .A(n45965), .B(n45966), .Z(n45953) );
  AND U45699 ( .A(n45967), .B(n45968), .Z(n45966) );
  XOR U45700 ( .A(n45965), .B(n45595), .Z(n45968) );
  XOR U45701 ( .A(n45969), .B(n45970), .Z(n45595) );
  AND U45702 ( .A(n903), .B(n45971), .Z(n45970) );
  XOR U45703 ( .A(n45972), .B(n45969), .Z(n45971) );
  XNOR U45704 ( .A(n45592), .B(n45965), .Z(n45967) );
  XOR U45705 ( .A(n45973), .B(n45974), .Z(n45592) );
  AND U45706 ( .A(n901), .B(n45975), .Z(n45974) );
  XOR U45707 ( .A(n45976), .B(n45973), .Z(n45975) );
  XOR U45708 ( .A(n45977), .B(n45978), .Z(n45965) );
  AND U45709 ( .A(n45979), .B(n45980), .Z(n45978) );
  XOR U45710 ( .A(n45977), .B(n45607), .Z(n45980) );
  XOR U45711 ( .A(n45981), .B(n45982), .Z(n45607) );
  AND U45712 ( .A(n903), .B(n45983), .Z(n45982) );
  XOR U45713 ( .A(n45984), .B(n45981), .Z(n45983) );
  XNOR U45714 ( .A(n45604), .B(n45977), .Z(n45979) );
  XOR U45715 ( .A(n45985), .B(n45986), .Z(n45604) );
  AND U45716 ( .A(n901), .B(n45987), .Z(n45986) );
  XOR U45717 ( .A(n45988), .B(n45985), .Z(n45987) );
  XOR U45718 ( .A(n45989), .B(n45990), .Z(n45977) );
  AND U45719 ( .A(n45991), .B(n45992), .Z(n45990) );
  XNOR U45720 ( .A(n45993), .B(n45620), .Z(n45992) );
  XOR U45721 ( .A(n45994), .B(n45995), .Z(n45620) );
  AND U45722 ( .A(n903), .B(n45996), .Z(n45995) );
  XOR U45723 ( .A(n45994), .B(n45997), .Z(n45996) );
  XNOR U45724 ( .A(n45617), .B(n45989), .Z(n45991) );
  XOR U45725 ( .A(n45998), .B(n45999), .Z(n45617) );
  AND U45726 ( .A(n901), .B(n46000), .Z(n45999) );
  XOR U45727 ( .A(n45998), .B(n46001), .Z(n46000) );
  IV U45728 ( .A(n45993), .Z(n45989) );
  AND U45729 ( .A(n45625), .B(n45628), .Z(n45993) );
  XNOR U45730 ( .A(n46002), .B(n46003), .Z(n45628) );
  AND U45731 ( .A(n903), .B(n46004), .Z(n46003) );
  XNOR U45732 ( .A(n46005), .B(n46002), .Z(n46004) );
  XOR U45733 ( .A(n46006), .B(n46007), .Z(n903) );
  AND U45734 ( .A(n46008), .B(n46009), .Z(n46007) );
  XOR U45735 ( .A(n46006), .B(n45636), .Z(n46009) );
  XNOR U45736 ( .A(n46010), .B(n46011), .Z(n45636) );
  AND U45737 ( .A(n46012), .B(n623), .Z(n46011) );
  AND U45738 ( .A(n46010), .B(n46013), .Z(n46012) );
  XNOR U45739 ( .A(n45633), .B(n46006), .Z(n46008) );
  XOR U45740 ( .A(n46014), .B(n46015), .Z(n45633) );
  AND U45741 ( .A(n46016), .B(n621), .Z(n46015) );
  NOR U45742 ( .A(n46014), .B(n46017), .Z(n46016) );
  XOR U45743 ( .A(n46018), .B(n46019), .Z(n46006) );
  AND U45744 ( .A(n46020), .B(n46021), .Z(n46019) );
  XOR U45745 ( .A(n46018), .B(n45648), .Z(n46021) );
  XOR U45746 ( .A(n46022), .B(n46023), .Z(n45648) );
  AND U45747 ( .A(n623), .B(n46024), .Z(n46023) );
  XOR U45748 ( .A(n46025), .B(n46022), .Z(n46024) );
  XNOR U45749 ( .A(n45645), .B(n46018), .Z(n46020) );
  XOR U45750 ( .A(n46026), .B(n46027), .Z(n45645) );
  AND U45751 ( .A(n621), .B(n46028), .Z(n46027) );
  XOR U45752 ( .A(n46029), .B(n46026), .Z(n46028) );
  XOR U45753 ( .A(n46030), .B(n46031), .Z(n46018) );
  AND U45754 ( .A(n46032), .B(n46033), .Z(n46031) );
  XOR U45755 ( .A(n46030), .B(n45660), .Z(n46033) );
  XOR U45756 ( .A(n46034), .B(n46035), .Z(n45660) );
  AND U45757 ( .A(n623), .B(n46036), .Z(n46035) );
  XOR U45758 ( .A(n46037), .B(n46034), .Z(n46036) );
  XNOR U45759 ( .A(n45657), .B(n46030), .Z(n46032) );
  XOR U45760 ( .A(n46038), .B(n46039), .Z(n45657) );
  AND U45761 ( .A(n621), .B(n46040), .Z(n46039) );
  XOR U45762 ( .A(n46041), .B(n46038), .Z(n46040) );
  XOR U45763 ( .A(n46042), .B(n46043), .Z(n46030) );
  AND U45764 ( .A(n46044), .B(n46045), .Z(n46043) );
  XOR U45765 ( .A(n46042), .B(n45672), .Z(n46045) );
  XOR U45766 ( .A(n46046), .B(n46047), .Z(n45672) );
  AND U45767 ( .A(n623), .B(n46048), .Z(n46047) );
  XOR U45768 ( .A(n46049), .B(n46046), .Z(n46048) );
  XNOR U45769 ( .A(n45669), .B(n46042), .Z(n46044) );
  XOR U45770 ( .A(n46050), .B(n46051), .Z(n45669) );
  AND U45771 ( .A(n621), .B(n46052), .Z(n46051) );
  XOR U45772 ( .A(n46053), .B(n46050), .Z(n46052) );
  XOR U45773 ( .A(n46054), .B(n46055), .Z(n46042) );
  AND U45774 ( .A(n46056), .B(n46057), .Z(n46055) );
  XOR U45775 ( .A(n46054), .B(n45684), .Z(n46057) );
  XOR U45776 ( .A(n46058), .B(n46059), .Z(n45684) );
  AND U45777 ( .A(n623), .B(n46060), .Z(n46059) );
  XOR U45778 ( .A(n46061), .B(n46058), .Z(n46060) );
  XNOR U45779 ( .A(n45681), .B(n46054), .Z(n46056) );
  XOR U45780 ( .A(n46062), .B(n46063), .Z(n45681) );
  AND U45781 ( .A(n621), .B(n46064), .Z(n46063) );
  XOR U45782 ( .A(n46065), .B(n46062), .Z(n46064) );
  XOR U45783 ( .A(n46066), .B(n46067), .Z(n46054) );
  AND U45784 ( .A(n46068), .B(n46069), .Z(n46067) );
  XOR U45785 ( .A(n46066), .B(n45696), .Z(n46069) );
  XOR U45786 ( .A(n46070), .B(n46071), .Z(n45696) );
  AND U45787 ( .A(n623), .B(n46072), .Z(n46071) );
  XOR U45788 ( .A(n46073), .B(n46070), .Z(n46072) );
  XNOR U45789 ( .A(n45693), .B(n46066), .Z(n46068) );
  XOR U45790 ( .A(n46074), .B(n46075), .Z(n45693) );
  AND U45791 ( .A(n621), .B(n46076), .Z(n46075) );
  XOR U45792 ( .A(n46077), .B(n46074), .Z(n46076) );
  XOR U45793 ( .A(n46078), .B(n46079), .Z(n46066) );
  AND U45794 ( .A(n46080), .B(n46081), .Z(n46079) );
  XOR U45795 ( .A(n46078), .B(n45708), .Z(n46081) );
  XOR U45796 ( .A(n46082), .B(n46083), .Z(n45708) );
  AND U45797 ( .A(n623), .B(n46084), .Z(n46083) );
  XOR U45798 ( .A(n46085), .B(n46082), .Z(n46084) );
  XNOR U45799 ( .A(n45705), .B(n46078), .Z(n46080) );
  XOR U45800 ( .A(n46086), .B(n46087), .Z(n45705) );
  AND U45801 ( .A(n621), .B(n46088), .Z(n46087) );
  XOR U45802 ( .A(n46089), .B(n46086), .Z(n46088) );
  XOR U45803 ( .A(n46090), .B(n46091), .Z(n46078) );
  AND U45804 ( .A(n46092), .B(n46093), .Z(n46091) );
  XOR U45805 ( .A(n46090), .B(n45720), .Z(n46093) );
  XOR U45806 ( .A(n46094), .B(n46095), .Z(n45720) );
  AND U45807 ( .A(n623), .B(n46096), .Z(n46095) );
  XOR U45808 ( .A(n46097), .B(n46094), .Z(n46096) );
  XNOR U45809 ( .A(n45717), .B(n46090), .Z(n46092) );
  XOR U45810 ( .A(n46098), .B(n46099), .Z(n45717) );
  AND U45811 ( .A(n621), .B(n46100), .Z(n46099) );
  XOR U45812 ( .A(n46101), .B(n46098), .Z(n46100) );
  XOR U45813 ( .A(n46102), .B(n46103), .Z(n46090) );
  AND U45814 ( .A(n46104), .B(n46105), .Z(n46103) );
  XOR U45815 ( .A(n46102), .B(n45732), .Z(n46105) );
  XOR U45816 ( .A(n46106), .B(n46107), .Z(n45732) );
  AND U45817 ( .A(n623), .B(n46108), .Z(n46107) );
  XOR U45818 ( .A(n46109), .B(n46106), .Z(n46108) );
  XNOR U45819 ( .A(n45729), .B(n46102), .Z(n46104) );
  XOR U45820 ( .A(n46110), .B(n46111), .Z(n45729) );
  AND U45821 ( .A(n621), .B(n46112), .Z(n46111) );
  XOR U45822 ( .A(n46113), .B(n46110), .Z(n46112) );
  XOR U45823 ( .A(n46114), .B(n46115), .Z(n46102) );
  AND U45824 ( .A(n46116), .B(n46117), .Z(n46115) );
  XOR U45825 ( .A(n46114), .B(n45744), .Z(n46117) );
  XOR U45826 ( .A(n46118), .B(n46119), .Z(n45744) );
  AND U45827 ( .A(n623), .B(n46120), .Z(n46119) );
  XOR U45828 ( .A(n46121), .B(n46118), .Z(n46120) );
  XNOR U45829 ( .A(n45741), .B(n46114), .Z(n46116) );
  XOR U45830 ( .A(n46122), .B(n46123), .Z(n45741) );
  AND U45831 ( .A(n621), .B(n46124), .Z(n46123) );
  XOR U45832 ( .A(n46125), .B(n46122), .Z(n46124) );
  XOR U45833 ( .A(n46126), .B(n46127), .Z(n46114) );
  AND U45834 ( .A(n46128), .B(n46129), .Z(n46127) );
  XOR U45835 ( .A(n46126), .B(n45756), .Z(n46129) );
  XOR U45836 ( .A(n46130), .B(n46131), .Z(n45756) );
  AND U45837 ( .A(n623), .B(n46132), .Z(n46131) );
  XOR U45838 ( .A(n46133), .B(n46130), .Z(n46132) );
  XNOR U45839 ( .A(n45753), .B(n46126), .Z(n46128) );
  XOR U45840 ( .A(n46134), .B(n46135), .Z(n45753) );
  AND U45841 ( .A(n621), .B(n46136), .Z(n46135) );
  XOR U45842 ( .A(n46137), .B(n46134), .Z(n46136) );
  XOR U45843 ( .A(n46138), .B(n46139), .Z(n46126) );
  AND U45844 ( .A(n46140), .B(n46141), .Z(n46139) );
  XOR U45845 ( .A(n46138), .B(n45768), .Z(n46141) );
  XOR U45846 ( .A(n46142), .B(n46143), .Z(n45768) );
  AND U45847 ( .A(n623), .B(n46144), .Z(n46143) );
  XOR U45848 ( .A(n46145), .B(n46142), .Z(n46144) );
  XNOR U45849 ( .A(n45765), .B(n46138), .Z(n46140) );
  XOR U45850 ( .A(n46146), .B(n46147), .Z(n45765) );
  AND U45851 ( .A(n621), .B(n46148), .Z(n46147) );
  XOR U45852 ( .A(n46149), .B(n46146), .Z(n46148) );
  XOR U45853 ( .A(n46150), .B(n46151), .Z(n46138) );
  AND U45854 ( .A(n46152), .B(n46153), .Z(n46151) );
  XOR U45855 ( .A(n46150), .B(n45780), .Z(n46153) );
  XOR U45856 ( .A(n46154), .B(n46155), .Z(n45780) );
  AND U45857 ( .A(n623), .B(n46156), .Z(n46155) );
  XOR U45858 ( .A(n46157), .B(n46154), .Z(n46156) );
  XNOR U45859 ( .A(n45777), .B(n46150), .Z(n46152) );
  XOR U45860 ( .A(n46158), .B(n46159), .Z(n45777) );
  AND U45861 ( .A(n621), .B(n46160), .Z(n46159) );
  XOR U45862 ( .A(n46161), .B(n46158), .Z(n46160) );
  XOR U45863 ( .A(n46162), .B(n46163), .Z(n46150) );
  AND U45864 ( .A(n46164), .B(n46165), .Z(n46163) );
  XOR U45865 ( .A(n46162), .B(n45792), .Z(n46165) );
  XOR U45866 ( .A(n46166), .B(n46167), .Z(n45792) );
  AND U45867 ( .A(n623), .B(n46168), .Z(n46167) );
  XOR U45868 ( .A(n46169), .B(n46166), .Z(n46168) );
  XNOR U45869 ( .A(n45789), .B(n46162), .Z(n46164) );
  XOR U45870 ( .A(n46170), .B(n46171), .Z(n45789) );
  AND U45871 ( .A(n621), .B(n46172), .Z(n46171) );
  XOR U45872 ( .A(n46173), .B(n46170), .Z(n46172) );
  XOR U45873 ( .A(n46174), .B(n46175), .Z(n46162) );
  AND U45874 ( .A(n46176), .B(n46177), .Z(n46175) );
  XOR U45875 ( .A(n46174), .B(n45804), .Z(n46177) );
  XOR U45876 ( .A(n46178), .B(n46179), .Z(n45804) );
  AND U45877 ( .A(n623), .B(n46180), .Z(n46179) );
  XOR U45878 ( .A(n46181), .B(n46178), .Z(n46180) );
  XNOR U45879 ( .A(n45801), .B(n46174), .Z(n46176) );
  XOR U45880 ( .A(n46182), .B(n46183), .Z(n45801) );
  AND U45881 ( .A(n621), .B(n46184), .Z(n46183) );
  XOR U45882 ( .A(n46185), .B(n46182), .Z(n46184) );
  XOR U45883 ( .A(n46186), .B(n46187), .Z(n46174) );
  AND U45884 ( .A(n46188), .B(n46189), .Z(n46187) );
  XOR U45885 ( .A(n46186), .B(n45816), .Z(n46189) );
  XOR U45886 ( .A(n46190), .B(n46191), .Z(n45816) );
  AND U45887 ( .A(n623), .B(n46192), .Z(n46191) );
  XOR U45888 ( .A(n46193), .B(n46190), .Z(n46192) );
  XNOR U45889 ( .A(n45813), .B(n46186), .Z(n46188) );
  XOR U45890 ( .A(n46194), .B(n46195), .Z(n45813) );
  AND U45891 ( .A(n621), .B(n46196), .Z(n46195) );
  XOR U45892 ( .A(n46197), .B(n46194), .Z(n46196) );
  XOR U45893 ( .A(n46198), .B(n46199), .Z(n46186) );
  AND U45894 ( .A(n46200), .B(n46201), .Z(n46199) );
  XOR U45895 ( .A(n46198), .B(n45828), .Z(n46201) );
  XOR U45896 ( .A(n46202), .B(n46203), .Z(n45828) );
  AND U45897 ( .A(n623), .B(n46204), .Z(n46203) );
  XOR U45898 ( .A(n46205), .B(n46202), .Z(n46204) );
  XNOR U45899 ( .A(n45825), .B(n46198), .Z(n46200) );
  XOR U45900 ( .A(n46206), .B(n46207), .Z(n45825) );
  AND U45901 ( .A(n621), .B(n46208), .Z(n46207) );
  XOR U45902 ( .A(n46209), .B(n46206), .Z(n46208) );
  XOR U45903 ( .A(n46210), .B(n46211), .Z(n46198) );
  AND U45904 ( .A(n46212), .B(n46213), .Z(n46211) );
  XOR U45905 ( .A(n46210), .B(n45840), .Z(n46213) );
  XOR U45906 ( .A(n46214), .B(n46215), .Z(n45840) );
  AND U45907 ( .A(n623), .B(n46216), .Z(n46215) );
  XOR U45908 ( .A(n46217), .B(n46214), .Z(n46216) );
  XNOR U45909 ( .A(n45837), .B(n46210), .Z(n46212) );
  XOR U45910 ( .A(n46218), .B(n46219), .Z(n45837) );
  AND U45911 ( .A(n621), .B(n46220), .Z(n46219) );
  XOR U45912 ( .A(n46221), .B(n46218), .Z(n46220) );
  XOR U45913 ( .A(n46222), .B(n46223), .Z(n46210) );
  AND U45914 ( .A(n46224), .B(n46225), .Z(n46223) );
  XOR U45915 ( .A(n46222), .B(n45852), .Z(n46225) );
  XOR U45916 ( .A(n46226), .B(n46227), .Z(n45852) );
  AND U45917 ( .A(n623), .B(n46228), .Z(n46227) );
  XOR U45918 ( .A(n46229), .B(n46226), .Z(n46228) );
  XNOR U45919 ( .A(n45849), .B(n46222), .Z(n46224) );
  XOR U45920 ( .A(n46230), .B(n46231), .Z(n45849) );
  AND U45921 ( .A(n621), .B(n46232), .Z(n46231) );
  XOR U45922 ( .A(n46233), .B(n46230), .Z(n46232) );
  XOR U45923 ( .A(n46234), .B(n46235), .Z(n46222) );
  AND U45924 ( .A(n46236), .B(n46237), .Z(n46235) );
  XOR U45925 ( .A(n46234), .B(n45864), .Z(n46237) );
  XOR U45926 ( .A(n46238), .B(n46239), .Z(n45864) );
  AND U45927 ( .A(n623), .B(n46240), .Z(n46239) );
  XOR U45928 ( .A(n46241), .B(n46238), .Z(n46240) );
  XNOR U45929 ( .A(n45861), .B(n46234), .Z(n46236) );
  XOR U45930 ( .A(n46242), .B(n46243), .Z(n45861) );
  AND U45931 ( .A(n621), .B(n46244), .Z(n46243) );
  XOR U45932 ( .A(n46245), .B(n46242), .Z(n46244) );
  XOR U45933 ( .A(n46246), .B(n46247), .Z(n46234) );
  AND U45934 ( .A(n46248), .B(n46249), .Z(n46247) );
  XOR U45935 ( .A(n46246), .B(n45876), .Z(n46249) );
  XOR U45936 ( .A(n46250), .B(n46251), .Z(n45876) );
  AND U45937 ( .A(n623), .B(n46252), .Z(n46251) );
  XOR U45938 ( .A(n46253), .B(n46250), .Z(n46252) );
  XNOR U45939 ( .A(n45873), .B(n46246), .Z(n46248) );
  XOR U45940 ( .A(n46254), .B(n46255), .Z(n45873) );
  AND U45941 ( .A(n621), .B(n46256), .Z(n46255) );
  XOR U45942 ( .A(n46257), .B(n46254), .Z(n46256) );
  XOR U45943 ( .A(n46258), .B(n46259), .Z(n46246) );
  AND U45944 ( .A(n46260), .B(n46261), .Z(n46259) );
  XOR U45945 ( .A(n46258), .B(n45888), .Z(n46261) );
  XOR U45946 ( .A(n46262), .B(n46263), .Z(n45888) );
  AND U45947 ( .A(n623), .B(n46264), .Z(n46263) );
  XOR U45948 ( .A(n46265), .B(n46262), .Z(n46264) );
  XNOR U45949 ( .A(n45885), .B(n46258), .Z(n46260) );
  XOR U45950 ( .A(n46266), .B(n46267), .Z(n45885) );
  AND U45951 ( .A(n621), .B(n46268), .Z(n46267) );
  XOR U45952 ( .A(n46269), .B(n46266), .Z(n46268) );
  XOR U45953 ( .A(n46270), .B(n46271), .Z(n46258) );
  AND U45954 ( .A(n46272), .B(n46273), .Z(n46271) );
  XOR U45955 ( .A(n46270), .B(n45900), .Z(n46273) );
  XOR U45956 ( .A(n46274), .B(n46275), .Z(n45900) );
  AND U45957 ( .A(n623), .B(n46276), .Z(n46275) );
  XOR U45958 ( .A(n46277), .B(n46274), .Z(n46276) );
  XNOR U45959 ( .A(n45897), .B(n46270), .Z(n46272) );
  XOR U45960 ( .A(n46278), .B(n46279), .Z(n45897) );
  AND U45961 ( .A(n621), .B(n46280), .Z(n46279) );
  XOR U45962 ( .A(n46281), .B(n46278), .Z(n46280) );
  XOR U45963 ( .A(n46282), .B(n46283), .Z(n46270) );
  AND U45964 ( .A(n46284), .B(n46285), .Z(n46283) );
  XOR U45965 ( .A(n46282), .B(n45912), .Z(n46285) );
  XOR U45966 ( .A(n46286), .B(n46287), .Z(n45912) );
  AND U45967 ( .A(n623), .B(n46288), .Z(n46287) );
  XOR U45968 ( .A(n46289), .B(n46286), .Z(n46288) );
  XNOR U45969 ( .A(n45909), .B(n46282), .Z(n46284) );
  XOR U45970 ( .A(n46290), .B(n46291), .Z(n45909) );
  AND U45971 ( .A(n621), .B(n46292), .Z(n46291) );
  XOR U45972 ( .A(n46293), .B(n46290), .Z(n46292) );
  XOR U45973 ( .A(n46294), .B(n46295), .Z(n46282) );
  AND U45974 ( .A(n46296), .B(n46297), .Z(n46295) );
  XOR U45975 ( .A(n46294), .B(n45924), .Z(n46297) );
  XOR U45976 ( .A(n46298), .B(n46299), .Z(n45924) );
  AND U45977 ( .A(n623), .B(n46300), .Z(n46299) );
  XOR U45978 ( .A(n46301), .B(n46298), .Z(n46300) );
  XNOR U45979 ( .A(n45921), .B(n46294), .Z(n46296) );
  XOR U45980 ( .A(n46302), .B(n46303), .Z(n45921) );
  AND U45981 ( .A(n621), .B(n46304), .Z(n46303) );
  XOR U45982 ( .A(n46305), .B(n46302), .Z(n46304) );
  XOR U45983 ( .A(n46306), .B(n46307), .Z(n46294) );
  AND U45984 ( .A(n46308), .B(n46309), .Z(n46307) );
  XOR U45985 ( .A(n46306), .B(n45936), .Z(n46309) );
  XOR U45986 ( .A(n46310), .B(n46311), .Z(n45936) );
  AND U45987 ( .A(n623), .B(n46312), .Z(n46311) );
  XOR U45988 ( .A(n46313), .B(n46310), .Z(n46312) );
  XNOR U45989 ( .A(n45933), .B(n46306), .Z(n46308) );
  XOR U45990 ( .A(n46314), .B(n46315), .Z(n45933) );
  AND U45991 ( .A(n621), .B(n46316), .Z(n46315) );
  XOR U45992 ( .A(n46317), .B(n46314), .Z(n46316) );
  XOR U45993 ( .A(n46318), .B(n46319), .Z(n46306) );
  AND U45994 ( .A(n46320), .B(n46321), .Z(n46319) );
  XOR U45995 ( .A(n46318), .B(n45948), .Z(n46321) );
  XOR U45996 ( .A(n46322), .B(n46323), .Z(n45948) );
  AND U45997 ( .A(n623), .B(n46324), .Z(n46323) );
  XOR U45998 ( .A(n46325), .B(n46322), .Z(n46324) );
  XNOR U45999 ( .A(n45945), .B(n46318), .Z(n46320) );
  XOR U46000 ( .A(n46326), .B(n46327), .Z(n45945) );
  AND U46001 ( .A(n621), .B(n46328), .Z(n46327) );
  XOR U46002 ( .A(n46329), .B(n46326), .Z(n46328) );
  XOR U46003 ( .A(n46330), .B(n46331), .Z(n46318) );
  AND U46004 ( .A(n46332), .B(n46333), .Z(n46331) );
  XOR U46005 ( .A(n46330), .B(n45960), .Z(n46333) );
  XOR U46006 ( .A(n46334), .B(n46335), .Z(n45960) );
  AND U46007 ( .A(n623), .B(n46336), .Z(n46335) );
  XOR U46008 ( .A(n46337), .B(n46334), .Z(n46336) );
  XNOR U46009 ( .A(n45957), .B(n46330), .Z(n46332) );
  XOR U46010 ( .A(n46338), .B(n46339), .Z(n45957) );
  AND U46011 ( .A(n621), .B(n46340), .Z(n46339) );
  XOR U46012 ( .A(n46341), .B(n46338), .Z(n46340) );
  XOR U46013 ( .A(n46342), .B(n46343), .Z(n46330) );
  AND U46014 ( .A(n46344), .B(n46345), .Z(n46343) );
  XOR U46015 ( .A(n46342), .B(n45972), .Z(n46345) );
  XOR U46016 ( .A(n46346), .B(n46347), .Z(n45972) );
  AND U46017 ( .A(n623), .B(n46348), .Z(n46347) );
  XOR U46018 ( .A(n46349), .B(n46346), .Z(n46348) );
  XNOR U46019 ( .A(n45969), .B(n46342), .Z(n46344) );
  XOR U46020 ( .A(n46350), .B(n46351), .Z(n45969) );
  AND U46021 ( .A(n621), .B(n46352), .Z(n46351) );
  XOR U46022 ( .A(n46353), .B(n46350), .Z(n46352) );
  XOR U46023 ( .A(n46354), .B(n46355), .Z(n46342) );
  AND U46024 ( .A(n46356), .B(n46357), .Z(n46355) );
  XOR U46025 ( .A(n46354), .B(n45984), .Z(n46357) );
  XOR U46026 ( .A(n46358), .B(n46359), .Z(n45984) );
  AND U46027 ( .A(n623), .B(n46360), .Z(n46359) );
  XOR U46028 ( .A(n46361), .B(n46358), .Z(n46360) );
  XNOR U46029 ( .A(n45981), .B(n46354), .Z(n46356) );
  XOR U46030 ( .A(n46362), .B(n46363), .Z(n45981) );
  AND U46031 ( .A(n621), .B(n46364), .Z(n46363) );
  XOR U46032 ( .A(n46365), .B(n46362), .Z(n46364) );
  XOR U46033 ( .A(n46366), .B(n46367), .Z(n46354) );
  AND U46034 ( .A(n46368), .B(n46369), .Z(n46367) );
  XNOR U46035 ( .A(n46370), .B(n45997), .Z(n46369) );
  XOR U46036 ( .A(n46371), .B(n46372), .Z(n45997) );
  AND U46037 ( .A(n623), .B(n46373), .Z(n46372) );
  XOR U46038 ( .A(n46371), .B(n46374), .Z(n46373) );
  XNOR U46039 ( .A(n45994), .B(n46366), .Z(n46368) );
  XOR U46040 ( .A(n46375), .B(n46376), .Z(n45994) );
  AND U46041 ( .A(n621), .B(n46377), .Z(n46376) );
  XOR U46042 ( .A(n46375), .B(n46378), .Z(n46377) );
  IV U46043 ( .A(n46370), .Z(n46366) );
  AND U46044 ( .A(n46002), .B(n46005), .Z(n46370) );
  XNOR U46045 ( .A(n46379), .B(n46380), .Z(n46005) );
  AND U46046 ( .A(n623), .B(n46381), .Z(n46380) );
  XNOR U46047 ( .A(n46382), .B(n46379), .Z(n46381) );
  XOR U46048 ( .A(n46383), .B(n46384), .Z(n623) );
  AND U46049 ( .A(n46385), .B(n46386), .Z(n46384) );
  XOR U46050 ( .A(n46013), .B(n46383), .Z(n46386) );
  IV U46051 ( .A(n46387), .Z(n46013) );
  AND U46052 ( .A(p_input[2047]), .B(p_input[2015]), .Z(n46387) );
  XOR U46053 ( .A(n46383), .B(n46010), .Z(n46385) );
  AND U46054 ( .A(p_input[1951]), .B(p_input[1983]), .Z(n46010) );
  XOR U46055 ( .A(n46388), .B(n46389), .Z(n46383) );
  AND U46056 ( .A(n46390), .B(n46391), .Z(n46389) );
  XOR U46057 ( .A(n46388), .B(n46025), .Z(n46391) );
  XNOR U46058 ( .A(p_input[2014]), .B(n46392), .Z(n46025) );
  AND U46059 ( .A(n939), .B(n46393), .Z(n46392) );
  XOR U46060 ( .A(p_input[2046]), .B(p_input[2014]), .Z(n46393) );
  XNOR U46061 ( .A(n46022), .B(n46388), .Z(n46390) );
  XOR U46062 ( .A(n46394), .B(n46395), .Z(n46022) );
  AND U46063 ( .A(n937), .B(n46396), .Z(n46395) );
  XOR U46064 ( .A(p_input[1982]), .B(p_input[1950]), .Z(n46396) );
  XOR U46065 ( .A(n46397), .B(n46398), .Z(n46388) );
  AND U46066 ( .A(n46399), .B(n46400), .Z(n46398) );
  XOR U46067 ( .A(n46397), .B(n46037), .Z(n46400) );
  XNOR U46068 ( .A(p_input[2013]), .B(n46401), .Z(n46037) );
  AND U46069 ( .A(n939), .B(n46402), .Z(n46401) );
  XOR U46070 ( .A(p_input[2045]), .B(p_input[2013]), .Z(n46402) );
  XNOR U46071 ( .A(n46034), .B(n46397), .Z(n46399) );
  XOR U46072 ( .A(n46403), .B(n46404), .Z(n46034) );
  AND U46073 ( .A(n937), .B(n46405), .Z(n46404) );
  XOR U46074 ( .A(p_input[1981]), .B(p_input[1949]), .Z(n46405) );
  XOR U46075 ( .A(n46406), .B(n46407), .Z(n46397) );
  AND U46076 ( .A(n46408), .B(n46409), .Z(n46407) );
  XOR U46077 ( .A(n46406), .B(n46049), .Z(n46409) );
  XNOR U46078 ( .A(p_input[2012]), .B(n46410), .Z(n46049) );
  AND U46079 ( .A(n939), .B(n46411), .Z(n46410) );
  XOR U46080 ( .A(p_input[2044]), .B(p_input[2012]), .Z(n46411) );
  XNOR U46081 ( .A(n46046), .B(n46406), .Z(n46408) );
  XOR U46082 ( .A(n46412), .B(n46413), .Z(n46046) );
  AND U46083 ( .A(n937), .B(n46414), .Z(n46413) );
  XOR U46084 ( .A(p_input[1980]), .B(p_input[1948]), .Z(n46414) );
  XOR U46085 ( .A(n46415), .B(n46416), .Z(n46406) );
  AND U46086 ( .A(n46417), .B(n46418), .Z(n46416) );
  XOR U46087 ( .A(n46415), .B(n46061), .Z(n46418) );
  XNOR U46088 ( .A(p_input[2011]), .B(n46419), .Z(n46061) );
  AND U46089 ( .A(n939), .B(n46420), .Z(n46419) );
  XOR U46090 ( .A(p_input[2043]), .B(p_input[2011]), .Z(n46420) );
  XNOR U46091 ( .A(n46058), .B(n46415), .Z(n46417) );
  XOR U46092 ( .A(n46421), .B(n46422), .Z(n46058) );
  AND U46093 ( .A(n937), .B(n46423), .Z(n46422) );
  XOR U46094 ( .A(p_input[1979]), .B(p_input[1947]), .Z(n46423) );
  XOR U46095 ( .A(n46424), .B(n46425), .Z(n46415) );
  AND U46096 ( .A(n46426), .B(n46427), .Z(n46425) );
  XOR U46097 ( .A(n46424), .B(n46073), .Z(n46427) );
  XNOR U46098 ( .A(p_input[2010]), .B(n46428), .Z(n46073) );
  AND U46099 ( .A(n939), .B(n46429), .Z(n46428) );
  XOR U46100 ( .A(p_input[2042]), .B(p_input[2010]), .Z(n46429) );
  XNOR U46101 ( .A(n46070), .B(n46424), .Z(n46426) );
  XOR U46102 ( .A(n46430), .B(n46431), .Z(n46070) );
  AND U46103 ( .A(n937), .B(n46432), .Z(n46431) );
  XOR U46104 ( .A(p_input[1978]), .B(p_input[1946]), .Z(n46432) );
  XOR U46105 ( .A(n46433), .B(n46434), .Z(n46424) );
  AND U46106 ( .A(n46435), .B(n46436), .Z(n46434) );
  XOR U46107 ( .A(n46433), .B(n46085), .Z(n46436) );
  XNOR U46108 ( .A(p_input[2009]), .B(n46437), .Z(n46085) );
  AND U46109 ( .A(n939), .B(n46438), .Z(n46437) );
  XOR U46110 ( .A(p_input[2041]), .B(p_input[2009]), .Z(n46438) );
  XNOR U46111 ( .A(n46082), .B(n46433), .Z(n46435) );
  XOR U46112 ( .A(n46439), .B(n46440), .Z(n46082) );
  AND U46113 ( .A(n937), .B(n46441), .Z(n46440) );
  XOR U46114 ( .A(p_input[1977]), .B(p_input[1945]), .Z(n46441) );
  XOR U46115 ( .A(n46442), .B(n46443), .Z(n46433) );
  AND U46116 ( .A(n46444), .B(n46445), .Z(n46443) );
  XOR U46117 ( .A(n46442), .B(n46097), .Z(n46445) );
  XNOR U46118 ( .A(p_input[2008]), .B(n46446), .Z(n46097) );
  AND U46119 ( .A(n939), .B(n46447), .Z(n46446) );
  XOR U46120 ( .A(p_input[2040]), .B(p_input[2008]), .Z(n46447) );
  XNOR U46121 ( .A(n46094), .B(n46442), .Z(n46444) );
  XOR U46122 ( .A(n46448), .B(n46449), .Z(n46094) );
  AND U46123 ( .A(n937), .B(n46450), .Z(n46449) );
  XOR U46124 ( .A(p_input[1976]), .B(p_input[1944]), .Z(n46450) );
  XOR U46125 ( .A(n46451), .B(n46452), .Z(n46442) );
  AND U46126 ( .A(n46453), .B(n46454), .Z(n46452) );
  XOR U46127 ( .A(n46451), .B(n46109), .Z(n46454) );
  XNOR U46128 ( .A(p_input[2007]), .B(n46455), .Z(n46109) );
  AND U46129 ( .A(n939), .B(n46456), .Z(n46455) );
  XOR U46130 ( .A(p_input[2039]), .B(p_input[2007]), .Z(n46456) );
  XNOR U46131 ( .A(n46106), .B(n46451), .Z(n46453) );
  XOR U46132 ( .A(n46457), .B(n46458), .Z(n46106) );
  AND U46133 ( .A(n937), .B(n46459), .Z(n46458) );
  XOR U46134 ( .A(p_input[1975]), .B(p_input[1943]), .Z(n46459) );
  XOR U46135 ( .A(n46460), .B(n46461), .Z(n46451) );
  AND U46136 ( .A(n46462), .B(n46463), .Z(n46461) );
  XOR U46137 ( .A(n46460), .B(n46121), .Z(n46463) );
  XNOR U46138 ( .A(p_input[2006]), .B(n46464), .Z(n46121) );
  AND U46139 ( .A(n939), .B(n46465), .Z(n46464) );
  XOR U46140 ( .A(p_input[2038]), .B(p_input[2006]), .Z(n46465) );
  XNOR U46141 ( .A(n46118), .B(n46460), .Z(n46462) );
  XOR U46142 ( .A(n46466), .B(n46467), .Z(n46118) );
  AND U46143 ( .A(n937), .B(n46468), .Z(n46467) );
  XOR U46144 ( .A(p_input[1974]), .B(p_input[1942]), .Z(n46468) );
  XOR U46145 ( .A(n46469), .B(n46470), .Z(n46460) );
  AND U46146 ( .A(n46471), .B(n46472), .Z(n46470) );
  XOR U46147 ( .A(n46469), .B(n46133), .Z(n46472) );
  XNOR U46148 ( .A(p_input[2005]), .B(n46473), .Z(n46133) );
  AND U46149 ( .A(n939), .B(n46474), .Z(n46473) );
  XOR U46150 ( .A(p_input[2037]), .B(p_input[2005]), .Z(n46474) );
  XNOR U46151 ( .A(n46130), .B(n46469), .Z(n46471) );
  XOR U46152 ( .A(n46475), .B(n46476), .Z(n46130) );
  AND U46153 ( .A(n937), .B(n46477), .Z(n46476) );
  XOR U46154 ( .A(p_input[1973]), .B(p_input[1941]), .Z(n46477) );
  XOR U46155 ( .A(n46478), .B(n46479), .Z(n46469) );
  AND U46156 ( .A(n46480), .B(n46481), .Z(n46479) );
  XOR U46157 ( .A(n46478), .B(n46145), .Z(n46481) );
  XNOR U46158 ( .A(p_input[2004]), .B(n46482), .Z(n46145) );
  AND U46159 ( .A(n939), .B(n46483), .Z(n46482) );
  XOR U46160 ( .A(p_input[2036]), .B(p_input[2004]), .Z(n46483) );
  XNOR U46161 ( .A(n46142), .B(n46478), .Z(n46480) );
  XOR U46162 ( .A(n46484), .B(n46485), .Z(n46142) );
  AND U46163 ( .A(n937), .B(n46486), .Z(n46485) );
  XOR U46164 ( .A(p_input[1972]), .B(p_input[1940]), .Z(n46486) );
  XOR U46165 ( .A(n46487), .B(n46488), .Z(n46478) );
  AND U46166 ( .A(n46489), .B(n46490), .Z(n46488) );
  XOR U46167 ( .A(n46487), .B(n46157), .Z(n46490) );
  XNOR U46168 ( .A(p_input[2003]), .B(n46491), .Z(n46157) );
  AND U46169 ( .A(n939), .B(n46492), .Z(n46491) );
  XOR U46170 ( .A(p_input[2035]), .B(p_input[2003]), .Z(n46492) );
  XNOR U46171 ( .A(n46154), .B(n46487), .Z(n46489) );
  XOR U46172 ( .A(n46493), .B(n46494), .Z(n46154) );
  AND U46173 ( .A(n937), .B(n46495), .Z(n46494) );
  XOR U46174 ( .A(p_input[1971]), .B(p_input[1939]), .Z(n46495) );
  XOR U46175 ( .A(n46496), .B(n46497), .Z(n46487) );
  AND U46176 ( .A(n46498), .B(n46499), .Z(n46497) );
  XOR U46177 ( .A(n46496), .B(n46169), .Z(n46499) );
  XNOR U46178 ( .A(p_input[2002]), .B(n46500), .Z(n46169) );
  AND U46179 ( .A(n939), .B(n46501), .Z(n46500) );
  XOR U46180 ( .A(p_input[2034]), .B(p_input[2002]), .Z(n46501) );
  XNOR U46181 ( .A(n46166), .B(n46496), .Z(n46498) );
  XOR U46182 ( .A(n46502), .B(n46503), .Z(n46166) );
  AND U46183 ( .A(n937), .B(n46504), .Z(n46503) );
  XOR U46184 ( .A(p_input[1970]), .B(p_input[1938]), .Z(n46504) );
  XOR U46185 ( .A(n46505), .B(n46506), .Z(n46496) );
  AND U46186 ( .A(n46507), .B(n46508), .Z(n46506) );
  XOR U46187 ( .A(n46505), .B(n46181), .Z(n46508) );
  XNOR U46188 ( .A(p_input[2001]), .B(n46509), .Z(n46181) );
  AND U46189 ( .A(n939), .B(n46510), .Z(n46509) );
  XOR U46190 ( .A(p_input[2033]), .B(p_input[2001]), .Z(n46510) );
  XNOR U46191 ( .A(n46178), .B(n46505), .Z(n46507) );
  XOR U46192 ( .A(n46511), .B(n46512), .Z(n46178) );
  AND U46193 ( .A(n937), .B(n46513), .Z(n46512) );
  XOR U46194 ( .A(p_input[1969]), .B(p_input[1937]), .Z(n46513) );
  XOR U46195 ( .A(n46514), .B(n46515), .Z(n46505) );
  AND U46196 ( .A(n46516), .B(n46517), .Z(n46515) );
  XOR U46197 ( .A(n46514), .B(n46193), .Z(n46517) );
  XNOR U46198 ( .A(p_input[2000]), .B(n46518), .Z(n46193) );
  AND U46199 ( .A(n939), .B(n46519), .Z(n46518) );
  XOR U46200 ( .A(p_input[2032]), .B(p_input[2000]), .Z(n46519) );
  XNOR U46201 ( .A(n46190), .B(n46514), .Z(n46516) );
  XOR U46202 ( .A(n46520), .B(n46521), .Z(n46190) );
  AND U46203 ( .A(n937), .B(n46522), .Z(n46521) );
  XOR U46204 ( .A(p_input[1968]), .B(p_input[1936]), .Z(n46522) );
  XOR U46205 ( .A(n46523), .B(n46524), .Z(n46514) );
  AND U46206 ( .A(n46525), .B(n46526), .Z(n46524) );
  XOR U46207 ( .A(n46523), .B(n46205), .Z(n46526) );
  XNOR U46208 ( .A(p_input[1999]), .B(n46527), .Z(n46205) );
  AND U46209 ( .A(n939), .B(n46528), .Z(n46527) );
  XOR U46210 ( .A(p_input[2031]), .B(p_input[1999]), .Z(n46528) );
  XNOR U46211 ( .A(n46202), .B(n46523), .Z(n46525) );
  XOR U46212 ( .A(n46529), .B(n46530), .Z(n46202) );
  AND U46213 ( .A(n937), .B(n46531), .Z(n46530) );
  XOR U46214 ( .A(p_input[1967]), .B(p_input[1935]), .Z(n46531) );
  XOR U46215 ( .A(n46532), .B(n46533), .Z(n46523) );
  AND U46216 ( .A(n46534), .B(n46535), .Z(n46533) );
  XOR U46217 ( .A(n46532), .B(n46217), .Z(n46535) );
  XNOR U46218 ( .A(p_input[1998]), .B(n46536), .Z(n46217) );
  AND U46219 ( .A(n939), .B(n46537), .Z(n46536) );
  XOR U46220 ( .A(p_input[2030]), .B(p_input[1998]), .Z(n46537) );
  XNOR U46221 ( .A(n46214), .B(n46532), .Z(n46534) );
  XOR U46222 ( .A(n46538), .B(n46539), .Z(n46214) );
  AND U46223 ( .A(n937), .B(n46540), .Z(n46539) );
  XOR U46224 ( .A(p_input[1966]), .B(p_input[1934]), .Z(n46540) );
  XOR U46225 ( .A(n46541), .B(n46542), .Z(n46532) );
  AND U46226 ( .A(n46543), .B(n46544), .Z(n46542) );
  XOR U46227 ( .A(n46541), .B(n46229), .Z(n46544) );
  XNOR U46228 ( .A(p_input[1997]), .B(n46545), .Z(n46229) );
  AND U46229 ( .A(n939), .B(n46546), .Z(n46545) );
  XOR U46230 ( .A(p_input[2029]), .B(p_input[1997]), .Z(n46546) );
  XNOR U46231 ( .A(n46226), .B(n46541), .Z(n46543) );
  XOR U46232 ( .A(n46547), .B(n46548), .Z(n46226) );
  AND U46233 ( .A(n937), .B(n46549), .Z(n46548) );
  XOR U46234 ( .A(p_input[1965]), .B(p_input[1933]), .Z(n46549) );
  XOR U46235 ( .A(n46550), .B(n46551), .Z(n46541) );
  AND U46236 ( .A(n46552), .B(n46553), .Z(n46551) );
  XOR U46237 ( .A(n46550), .B(n46241), .Z(n46553) );
  XNOR U46238 ( .A(p_input[1996]), .B(n46554), .Z(n46241) );
  AND U46239 ( .A(n939), .B(n46555), .Z(n46554) );
  XOR U46240 ( .A(p_input[2028]), .B(p_input[1996]), .Z(n46555) );
  XNOR U46241 ( .A(n46238), .B(n46550), .Z(n46552) );
  XOR U46242 ( .A(n46556), .B(n46557), .Z(n46238) );
  AND U46243 ( .A(n937), .B(n46558), .Z(n46557) );
  XOR U46244 ( .A(p_input[1964]), .B(p_input[1932]), .Z(n46558) );
  XOR U46245 ( .A(n46559), .B(n46560), .Z(n46550) );
  AND U46246 ( .A(n46561), .B(n46562), .Z(n46560) );
  XOR U46247 ( .A(n46559), .B(n46253), .Z(n46562) );
  XNOR U46248 ( .A(p_input[1995]), .B(n46563), .Z(n46253) );
  AND U46249 ( .A(n939), .B(n46564), .Z(n46563) );
  XOR U46250 ( .A(p_input[2027]), .B(p_input[1995]), .Z(n46564) );
  XNOR U46251 ( .A(n46250), .B(n46559), .Z(n46561) );
  XOR U46252 ( .A(n46565), .B(n46566), .Z(n46250) );
  AND U46253 ( .A(n937), .B(n46567), .Z(n46566) );
  XOR U46254 ( .A(p_input[1963]), .B(p_input[1931]), .Z(n46567) );
  XOR U46255 ( .A(n46568), .B(n46569), .Z(n46559) );
  AND U46256 ( .A(n46570), .B(n46571), .Z(n46569) );
  XOR U46257 ( .A(n46568), .B(n46265), .Z(n46571) );
  XNOR U46258 ( .A(p_input[1994]), .B(n46572), .Z(n46265) );
  AND U46259 ( .A(n939), .B(n46573), .Z(n46572) );
  XOR U46260 ( .A(p_input[2026]), .B(p_input[1994]), .Z(n46573) );
  XNOR U46261 ( .A(n46262), .B(n46568), .Z(n46570) );
  XOR U46262 ( .A(n46574), .B(n46575), .Z(n46262) );
  AND U46263 ( .A(n937), .B(n46576), .Z(n46575) );
  XOR U46264 ( .A(p_input[1962]), .B(p_input[1930]), .Z(n46576) );
  XOR U46265 ( .A(n46577), .B(n46578), .Z(n46568) );
  AND U46266 ( .A(n46579), .B(n46580), .Z(n46578) );
  XOR U46267 ( .A(n46577), .B(n46277), .Z(n46580) );
  XNOR U46268 ( .A(p_input[1993]), .B(n46581), .Z(n46277) );
  AND U46269 ( .A(n939), .B(n46582), .Z(n46581) );
  XOR U46270 ( .A(p_input[2025]), .B(p_input[1993]), .Z(n46582) );
  XNOR U46271 ( .A(n46274), .B(n46577), .Z(n46579) );
  XOR U46272 ( .A(n46583), .B(n46584), .Z(n46274) );
  AND U46273 ( .A(n937), .B(n46585), .Z(n46584) );
  XOR U46274 ( .A(p_input[1961]), .B(p_input[1929]), .Z(n46585) );
  XOR U46275 ( .A(n46586), .B(n46587), .Z(n46577) );
  AND U46276 ( .A(n46588), .B(n46589), .Z(n46587) );
  XOR U46277 ( .A(n46586), .B(n46289), .Z(n46589) );
  XNOR U46278 ( .A(p_input[1992]), .B(n46590), .Z(n46289) );
  AND U46279 ( .A(n939), .B(n46591), .Z(n46590) );
  XOR U46280 ( .A(p_input[2024]), .B(p_input[1992]), .Z(n46591) );
  XNOR U46281 ( .A(n46286), .B(n46586), .Z(n46588) );
  XOR U46282 ( .A(n46592), .B(n46593), .Z(n46286) );
  AND U46283 ( .A(n937), .B(n46594), .Z(n46593) );
  XOR U46284 ( .A(p_input[1960]), .B(p_input[1928]), .Z(n46594) );
  XOR U46285 ( .A(n46595), .B(n46596), .Z(n46586) );
  AND U46286 ( .A(n46597), .B(n46598), .Z(n46596) );
  XOR U46287 ( .A(n46595), .B(n46301), .Z(n46598) );
  XNOR U46288 ( .A(p_input[1991]), .B(n46599), .Z(n46301) );
  AND U46289 ( .A(n939), .B(n46600), .Z(n46599) );
  XOR U46290 ( .A(p_input[2023]), .B(p_input[1991]), .Z(n46600) );
  XNOR U46291 ( .A(n46298), .B(n46595), .Z(n46597) );
  XOR U46292 ( .A(n46601), .B(n46602), .Z(n46298) );
  AND U46293 ( .A(n937), .B(n46603), .Z(n46602) );
  XOR U46294 ( .A(p_input[1959]), .B(p_input[1927]), .Z(n46603) );
  XOR U46295 ( .A(n46604), .B(n46605), .Z(n46595) );
  AND U46296 ( .A(n46606), .B(n46607), .Z(n46605) );
  XOR U46297 ( .A(n46604), .B(n46313), .Z(n46607) );
  XNOR U46298 ( .A(p_input[1990]), .B(n46608), .Z(n46313) );
  AND U46299 ( .A(n939), .B(n46609), .Z(n46608) );
  XOR U46300 ( .A(p_input[2022]), .B(p_input[1990]), .Z(n46609) );
  XNOR U46301 ( .A(n46310), .B(n46604), .Z(n46606) );
  XOR U46302 ( .A(n46610), .B(n46611), .Z(n46310) );
  AND U46303 ( .A(n937), .B(n46612), .Z(n46611) );
  XOR U46304 ( .A(p_input[1958]), .B(p_input[1926]), .Z(n46612) );
  XOR U46305 ( .A(n46613), .B(n46614), .Z(n46604) );
  AND U46306 ( .A(n46615), .B(n46616), .Z(n46614) );
  XOR U46307 ( .A(n46613), .B(n46325), .Z(n46616) );
  XNOR U46308 ( .A(p_input[1989]), .B(n46617), .Z(n46325) );
  AND U46309 ( .A(n939), .B(n46618), .Z(n46617) );
  XOR U46310 ( .A(p_input[2021]), .B(p_input[1989]), .Z(n46618) );
  XNOR U46311 ( .A(n46322), .B(n46613), .Z(n46615) );
  XOR U46312 ( .A(n46619), .B(n46620), .Z(n46322) );
  AND U46313 ( .A(n937), .B(n46621), .Z(n46620) );
  XOR U46314 ( .A(p_input[1957]), .B(p_input[1925]), .Z(n46621) );
  XOR U46315 ( .A(n46622), .B(n46623), .Z(n46613) );
  AND U46316 ( .A(n46624), .B(n46625), .Z(n46623) );
  XOR U46317 ( .A(n46622), .B(n46337), .Z(n46625) );
  XNOR U46318 ( .A(p_input[1988]), .B(n46626), .Z(n46337) );
  AND U46319 ( .A(n939), .B(n46627), .Z(n46626) );
  XOR U46320 ( .A(p_input[2020]), .B(p_input[1988]), .Z(n46627) );
  XNOR U46321 ( .A(n46334), .B(n46622), .Z(n46624) );
  XOR U46322 ( .A(n46628), .B(n46629), .Z(n46334) );
  AND U46323 ( .A(n937), .B(n46630), .Z(n46629) );
  XOR U46324 ( .A(p_input[1956]), .B(p_input[1924]), .Z(n46630) );
  XOR U46325 ( .A(n46631), .B(n46632), .Z(n46622) );
  AND U46326 ( .A(n46633), .B(n46634), .Z(n46632) );
  XOR U46327 ( .A(n46631), .B(n46349), .Z(n46634) );
  XNOR U46328 ( .A(p_input[1987]), .B(n46635), .Z(n46349) );
  AND U46329 ( .A(n939), .B(n46636), .Z(n46635) );
  XOR U46330 ( .A(p_input[2019]), .B(p_input[1987]), .Z(n46636) );
  XNOR U46331 ( .A(n46346), .B(n46631), .Z(n46633) );
  XOR U46332 ( .A(n46637), .B(n46638), .Z(n46346) );
  AND U46333 ( .A(n937), .B(n46639), .Z(n46638) );
  XOR U46334 ( .A(p_input[1955]), .B(p_input[1923]), .Z(n46639) );
  XOR U46335 ( .A(n46640), .B(n46641), .Z(n46631) );
  AND U46336 ( .A(n46642), .B(n46643), .Z(n46641) );
  XOR U46337 ( .A(n46640), .B(n46361), .Z(n46643) );
  XNOR U46338 ( .A(p_input[1986]), .B(n46644), .Z(n46361) );
  AND U46339 ( .A(n939), .B(n46645), .Z(n46644) );
  XOR U46340 ( .A(p_input[2018]), .B(p_input[1986]), .Z(n46645) );
  XNOR U46341 ( .A(n46358), .B(n46640), .Z(n46642) );
  XOR U46342 ( .A(n46646), .B(n46647), .Z(n46358) );
  AND U46343 ( .A(n937), .B(n46648), .Z(n46647) );
  XOR U46344 ( .A(p_input[1954]), .B(p_input[1922]), .Z(n46648) );
  XOR U46345 ( .A(n46649), .B(n46650), .Z(n46640) );
  AND U46346 ( .A(n46651), .B(n46652), .Z(n46650) );
  XNOR U46347 ( .A(n46653), .B(n46374), .Z(n46652) );
  XNOR U46348 ( .A(p_input[1985]), .B(n46654), .Z(n46374) );
  AND U46349 ( .A(n939), .B(n46655), .Z(n46654) );
  XNOR U46350 ( .A(p_input[2017]), .B(n46656), .Z(n46655) );
  IV U46351 ( .A(p_input[1985]), .Z(n46656) );
  XNOR U46352 ( .A(n46371), .B(n46649), .Z(n46651) );
  XNOR U46353 ( .A(p_input[1921]), .B(n46657), .Z(n46371) );
  AND U46354 ( .A(n937), .B(n46658), .Z(n46657) );
  XOR U46355 ( .A(p_input[1953]), .B(p_input[1921]), .Z(n46658) );
  IV U46356 ( .A(n46653), .Z(n46649) );
  AND U46357 ( .A(n46379), .B(n46382), .Z(n46653) );
  XOR U46358 ( .A(p_input[1984]), .B(n46659), .Z(n46382) );
  AND U46359 ( .A(n939), .B(n46660), .Z(n46659) );
  XOR U46360 ( .A(p_input[2016]), .B(p_input[1984]), .Z(n46660) );
  XOR U46361 ( .A(n46661), .B(n46662), .Z(n939) );
  AND U46362 ( .A(n46663), .B(n46664), .Z(n46662) );
  XNOR U46363 ( .A(p_input[2047]), .B(n46661), .Z(n46664) );
  XOR U46364 ( .A(n46661), .B(p_input[2015]), .Z(n46663) );
  XOR U46365 ( .A(n46665), .B(n46666), .Z(n46661) );
  AND U46366 ( .A(n46667), .B(n46668), .Z(n46666) );
  XNOR U46367 ( .A(p_input[2046]), .B(n46665), .Z(n46668) );
  XOR U46368 ( .A(n46665), .B(p_input[2014]), .Z(n46667) );
  XOR U46369 ( .A(n46669), .B(n46670), .Z(n46665) );
  AND U46370 ( .A(n46671), .B(n46672), .Z(n46670) );
  XNOR U46371 ( .A(p_input[2045]), .B(n46669), .Z(n46672) );
  XOR U46372 ( .A(n46669), .B(p_input[2013]), .Z(n46671) );
  XOR U46373 ( .A(n46673), .B(n46674), .Z(n46669) );
  AND U46374 ( .A(n46675), .B(n46676), .Z(n46674) );
  XNOR U46375 ( .A(p_input[2044]), .B(n46673), .Z(n46676) );
  XOR U46376 ( .A(n46673), .B(p_input[2012]), .Z(n46675) );
  XOR U46377 ( .A(n46677), .B(n46678), .Z(n46673) );
  AND U46378 ( .A(n46679), .B(n46680), .Z(n46678) );
  XNOR U46379 ( .A(p_input[2043]), .B(n46677), .Z(n46680) );
  XOR U46380 ( .A(n46677), .B(p_input[2011]), .Z(n46679) );
  XOR U46381 ( .A(n46681), .B(n46682), .Z(n46677) );
  AND U46382 ( .A(n46683), .B(n46684), .Z(n46682) );
  XNOR U46383 ( .A(p_input[2042]), .B(n46681), .Z(n46684) );
  XOR U46384 ( .A(n46681), .B(p_input[2010]), .Z(n46683) );
  XOR U46385 ( .A(n46685), .B(n46686), .Z(n46681) );
  AND U46386 ( .A(n46687), .B(n46688), .Z(n46686) );
  XNOR U46387 ( .A(p_input[2041]), .B(n46685), .Z(n46688) );
  XOR U46388 ( .A(n46685), .B(p_input[2009]), .Z(n46687) );
  XOR U46389 ( .A(n46689), .B(n46690), .Z(n46685) );
  AND U46390 ( .A(n46691), .B(n46692), .Z(n46690) );
  XNOR U46391 ( .A(p_input[2040]), .B(n46689), .Z(n46692) );
  XOR U46392 ( .A(n46689), .B(p_input[2008]), .Z(n46691) );
  XOR U46393 ( .A(n46693), .B(n46694), .Z(n46689) );
  AND U46394 ( .A(n46695), .B(n46696), .Z(n46694) );
  XNOR U46395 ( .A(p_input[2039]), .B(n46693), .Z(n46696) );
  XOR U46396 ( .A(n46693), .B(p_input[2007]), .Z(n46695) );
  XOR U46397 ( .A(n46697), .B(n46698), .Z(n46693) );
  AND U46398 ( .A(n46699), .B(n46700), .Z(n46698) );
  XNOR U46399 ( .A(p_input[2038]), .B(n46697), .Z(n46700) );
  XOR U46400 ( .A(n46697), .B(p_input[2006]), .Z(n46699) );
  XOR U46401 ( .A(n46701), .B(n46702), .Z(n46697) );
  AND U46402 ( .A(n46703), .B(n46704), .Z(n46702) );
  XNOR U46403 ( .A(p_input[2037]), .B(n46701), .Z(n46704) );
  XOR U46404 ( .A(n46701), .B(p_input[2005]), .Z(n46703) );
  XOR U46405 ( .A(n46705), .B(n46706), .Z(n46701) );
  AND U46406 ( .A(n46707), .B(n46708), .Z(n46706) );
  XNOR U46407 ( .A(p_input[2036]), .B(n46705), .Z(n46708) );
  XOR U46408 ( .A(n46705), .B(p_input[2004]), .Z(n46707) );
  XOR U46409 ( .A(n46709), .B(n46710), .Z(n46705) );
  AND U46410 ( .A(n46711), .B(n46712), .Z(n46710) );
  XNOR U46411 ( .A(p_input[2035]), .B(n46709), .Z(n46712) );
  XOR U46412 ( .A(n46709), .B(p_input[2003]), .Z(n46711) );
  XOR U46413 ( .A(n46713), .B(n46714), .Z(n46709) );
  AND U46414 ( .A(n46715), .B(n46716), .Z(n46714) );
  XNOR U46415 ( .A(p_input[2034]), .B(n46713), .Z(n46716) );
  XOR U46416 ( .A(n46713), .B(p_input[2002]), .Z(n46715) );
  XOR U46417 ( .A(n46717), .B(n46718), .Z(n46713) );
  AND U46418 ( .A(n46719), .B(n46720), .Z(n46718) );
  XNOR U46419 ( .A(p_input[2033]), .B(n46717), .Z(n46720) );
  XOR U46420 ( .A(n46717), .B(p_input[2001]), .Z(n46719) );
  XOR U46421 ( .A(n46721), .B(n46722), .Z(n46717) );
  AND U46422 ( .A(n46723), .B(n46724), .Z(n46722) );
  XNOR U46423 ( .A(p_input[2032]), .B(n46721), .Z(n46724) );
  XOR U46424 ( .A(n46721), .B(p_input[2000]), .Z(n46723) );
  XOR U46425 ( .A(n46725), .B(n46726), .Z(n46721) );
  AND U46426 ( .A(n46727), .B(n46728), .Z(n46726) );
  XNOR U46427 ( .A(p_input[2031]), .B(n46725), .Z(n46728) );
  XOR U46428 ( .A(n46725), .B(p_input[1999]), .Z(n46727) );
  XOR U46429 ( .A(n46729), .B(n46730), .Z(n46725) );
  AND U46430 ( .A(n46731), .B(n46732), .Z(n46730) );
  XNOR U46431 ( .A(p_input[2030]), .B(n46729), .Z(n46732) );
  XOR U46432 ( .A(n46729), .B(p_input[1998]), .Z(n46731) );
  XOR U46433 ( .A(n46733), .B(n46734), .Z(n46729) );
  AND U46434 ( .A(n46735), .B(n46736), .Z(n46734) );
  XNOR U46435 ( .A(p_input[2029]), .B(n46733), .Z(n46736) );
  XOR U46436 ( .A(n46733), .B(p_input[1997]), .Z(n46735) );
  XOR U46437 ( .A(n46737), .B(n46738), .Z(n46733) );
  AND U46438 ( .A(n46739), .B(n46740), .Z(n46738) );
  XNOR U46439 ( .A(p_input[2028]), .B(n46737), .Z(n46740) );
  XOR U46440 ( .A(n46737), .B(p_input[1996]), .Z(n46739) );
  XOR U46441 ( .A(n46741), .B(n46742), .Z(n46737) );
  AND U46442 ( .A(n46743), .B(n46744), .Z(n46742) );
  XNOR U46443 ( .A(p_input[2027]), .B(n46741), .Z(n46744) );
  XOR U46444 ( .A(n46741), .B(p_input[1995]), .Z(n46743) );
  XOR U46445 ( .A(n46745), .B(n46746), .Z(n46741) );
  AND U46446 ( .A(n46747), .B(n46748), .Z(n46746) );
  XNOR U46447 ( .A(p_input[2026]), .B(n46745), .Z(n46748) );
  XOR U46448 ( .A(n46745), .B(p_input[1994]), .Z(n46747) );
  XOR U46449 ( .A(n46749), .B(n46750), .Z(n46745) );
  AND U46450 ( .A(n46751), .B(n46752), .Z(n46750) );
  XNOR U46451 ( .A(p_input[2025]), .B(n46749), .Z(n46752) );
  XOR U46452 ( .A(n46749), .B(p_input[1993]), .Z(n46751) );
  XOR U46453 ( .A(n46753), .B(n46754), .Z(n46749) );
  AND U46454 ( .A(n46755), .B(n46756), .Z(n46754) );
  XNOR U46455 ( .A(p_input[2024]), .B(n46753), .Z(n46756) );
  XOR U46456 ( .A(n46753), .B(p_input[1992]), .Z(n46755) );
  XOR U46457 ( .A(n46757), .B(n46758), .Z(n46753) );
  AND U46458 ( .A(n46759), .B(n46760), .Z(n46758) );
  XNOR U46459 ( .A(p_input[2023]), .B(n46757), .Z(n46760) );
  XOR U46460 ( .A(n46757), .B(p_input[1991]), .Z(n46759) );
  XOR U46461 ( .A(n46761), .B(n46762), .Z(n46757) );
  AND U46462 ( .A(n46763), .B(n46764), .Z(n46762) );
  XNOR U46463 ( .A(p_input[2022]), .B(n46761), .Z(n46764) );
  XOR U46464 ( .A(n46761), .B(p_input[1990]), .Z(n46763) );
  XOR U46465 ( .A(n46765), .B(n46766), .Z(n46761) );
  AND U46466 ( .A(n46767), .B(n46768), .Z(n46766) );
  XNOR U46467 ( .A(p_input[2021]), .B(n46765), .Z(n46768) );
  XOR U46468 ( .A(n46765), .B(p_input[1989]), .Z(n46767) );
  XOR U46469 ( .A(n46769), .B(n46770), .Z(n46765) );
  AND U46470 ( .A(n46771), .B(n46772), .Z(n46770) );
  XNOR U46471 ( .A(p_input[2020]), .B(n46769), .Z(n46772) );
  XOR U46472 ( .A(n46769), .B(p_input[1988]), .Z(n46771) );
  XOR U46473 ( .A(n46773), .B(n46774), .Z(n46769) );
  AND U46474 ( .A(n46775), .B(n46776), .Z(n46774) );
  XNOR U46475 ( .A(p_input[2019]), .B(n46773), .Z(n46776) );
  XOR U46476 ( .A(n46773), .B(p_input[1987]), .Z(n46775) );
  XOR U46477 ( .A(n46777), .B(n46778), .Z(n46773) );
  AND U46478 ( .A(n46779), .B(n46780), .Z(n46778) );
  XNOR U46479 ( .A(p_input[2018]), .B(n46777), .Z(n46780) );
  XOR U46480 ( .A(n46777), .B(p_input[1986]), .Z(n46779) );
  XNOR U46481 ( .A(n46781), .B(n46782), .Z(n46777) );
  AND U46482 ( .A(n46783), .B(n46784), .Z(n46782) );
  XOR U46483 ( .A(p_input[2017]), .B(n46781), .Z(n46784) );
  XNOR U46484 ( .A(p_input[1985]), .B(n46781), .Z(n46783) );
  AND U46485 ( .A(p_input[2016]), .B(n46785), .Z(n46781) );
  IV U46486 ( .A(p_input[1984]), .Z(n46785) );
  XNOR U46487 ( .A(p_input[1920]), .B(n46786), .Z(n46379) );
  AND U46488 ( .A(n937), .B(n46787), .Z(n46786) );
  XOR U46489 ( .A(p_input[1952]), .B(p_input[1920]), .Z(n46787) );
  XOR U46490 ( .A(n46788), .B(n46789), .Z(n937) );
  AND U46491 ( .A(n46790), .B(n46791), .Z(n46789) );
  XNOR U46492 ( .A(p_input[1983]), .B(n46788), .Z(n46791) );
  XOR U46493 ( .A(n46788), .B(p_input[1951]), .Z(n46790) );
  XOR U46494 ( .A(n46792), .B(n46793), .Z(n46788) );
  AND U46495 ( .A(n46794), .B(n46795), .Z(n46793) );
  XNOR U46496 ( .A(p_input[1982]), .B(n46792), .Z(n46795) );
  XNOR U46497 ( .A(n46792), .B(n46394), .Z(n46794) );
  IV U46498 ( .A(p_input[1950]), .Z(n46394) );
  XOR U46499 ( .A(n46796), .B(n46797), .Z(n46792) );
  AND U46500 ( .A(n46798), .B(n46799), .Z(n46797) );
  XNOR U46501 ( .A(p_input[1981]), .B(n46796), .Z(n46799) );
  XNOR U46502 ( .A(n46796), .B(n46403), .Z(n46798) );
  IV U46503 ( .A(p_input[1949]), .Z(n46403) );
  XOR U46504 ( .A(n46800), .B(n46801), .Z(n46796) );
  AND U46505 ( .A(n46802), .B(n46803), .Z(n46801) );
  XNOR U46506 ( .A(p_input[1980]), .B(n46800), .Z(n46803) );
  XNOR U46507 ( .A(n46800), .B(n46412), .Z(n46802) );
  IV U46508 ( .A(p_input[1948]), .Z(n46412) );
  XOR U46509 ( .A(n46804), .B(n46805), .Z(n46800) );
  AND U46510 ( .A(n46806), .B(n46807), .Z(n46805) );
  XNOR U46511 ( .A(p_input[1979]), .B(n46804), .Z(n46807) );
  XNOR U46512 ( .A(n46804), .B(n46421), .Z(n46806) );
  IV U46513 ( .A(p_input[1947]), .Z(n46421) );
  XOR U46514 ( .A(n46808), .B(n46809), .Z(n46804) );
  AND U46515 ( .A(n46810), .B(n46811), .Z(n46809) );
  XNOR U46516 ( .A(p_input[1978]), .B(n46808), .Z(n46811) );
  XNOR U46517 ( .A(n46808), .B(n46430), .Z(n46810) );
  IV U46518 ( .A(p_input[1946]), .Z(n46430) );
  XOR U46519 ( .A(n46812), .B(n46813), .Z(n46808) );
  AND U46520 ( .A(n46814), .B(n46815), .Z(n46813) );
  XNOR U46521 ( .A(p_input[1977]), .B(n46812), .Z(n46815) );
  XNOR U46522 ( .A(n46812), .B(n46439), .Z(n46814) );
  IV U46523 ( .A(p_input[1945]), .Z(n46439) );
  XOR U46524 ( .A(n46816), .B(n46817), .Z(n46812) );
  AND U46525 ( .A(n46818), .B(n46819), .Z(n46817) );
  XNOR U46526 ( .A(p_input[1976]), .B(n46816), .Z(n46819) );
  XNOR U46527 ( .A(n46816), .B(n46448), .Z(n46818) );
  IV U46528 ( .A(p_input[1944]), .Z(n46448) );
  XOR U46529 ( .A(n46820), .B(n46821), .Z(n46816) );
  AND U46530 ( .A(n46822), .B(n46823), .Z(n46821) );
  XNOR U46531 ( .A(p_input[1975]), .B(n46820), .Z(n46823) );
  XNOR U46532 ( .A(n46820), .B(n46457), .Z(n46822) );
  IV U46533 ( .A(p_input[1943]), .Z(n46457) );
  XOR U46534 ( .A(n46824), .B(n46825), .Z(n46820) );
  AND U46535 ( .A(n46826), .B(n46827), .Z(n46825) );
  XNOR U46536 ( .A(p_input[1974]), .B(n46824), .Z(n46827) );
  XNOR U46537 ( .A(n46824), .B(n46466), .Z(n46826) );
  IV U46538 ( .A(p_input[1942]), .Z(n46466) );
  XOR U46539 ( .A(n46828), .B(n46829), .Z(n46824) );
  AND U46540 ( .A(n46830), .B(n46831), .Z(n46829) );
  XNOR U46541 ( .A(p_input[1973]), .B(n46828), .Z(n46831) );
  XNOR U46542 ( .A(n46828), .B(n46475), .Z(n46830) );
  IV U46543 ( .A(p_input[1941]), .Z(n46475) );
  XOR U46544 ( .A(n46832), .B(n46833), .Z(n46828) );
  AND U46545 ( .A(n46834), .B(n46835), .Z(n46833) );
  XNOR U46546 ( .A(p_input[1972]), .B(n46832), .Z(n46835) );
  XNOR U46547 ( .A(n46832), .B(n46484), .Z(n46834) );
  IV U46548 ( .A(p_input[1940]), .Z(n46484) );
  XOR U46549 ( .A(n46836), .B(n46837), .Z(n46832) );
  AND U46550 ( .A(n46838), .B(n46839), .Z(n46837) );
  XNOR U46551 ( .A(p_input[1971]), .B(n46836), .Z(n46839) );
  XNOR U46552 ( .A(n46836), .B(n46493), .Z(n46838) );
  IV U46553 ( .A(p_input[1939]), .Z(n46493) );
  XOR U46554 ( .A(n46840), .B(n46841), .Z(n46836) );
  AND U46555 ( .A(n46842), .B(n46843), .Z(n46841) );
  XNOR U46556 ( .A(p_input[1970]), .B(n46840), .Z(n46843) );
  XNOR U46557 ( .A(n46840), .B(n46502), .Z(n46842) );
  IV U46558 ( .A(p_input[1938]), .Z(n46502) );
  XOR U46559 ( .A(n46844), .B(n46845), .Z(n46840) );
  AND U46560 ( .A(n46846), .B(n46847), .Z(n46845) );
  XNOR U46561 ( .A(p_input[1969]), .B(n46844), .Z(n46847) );
  XNOR U46562 ( .A(n46844), .B(n46511), .Z(n46846) );
  IV U46563 ( .A(p_input[1937]), .Z(n46511) );
  XOR U46564 ( .A(n46848), .B(n46849), .Z(n46844) );
  AND U46565 ( .A(n46850), .B(n46851), .Z(n46849) );
  XNOR U46566 ( .A(p_input[1968]), .B(n46848), .Z(n46851) );
  XNOR U46567 ( .A(n46848), .B(n46520), .Z(n46850) );
  IV U46568 ( .A(p_input[1936]), .Z(n46520) );
  XOR U46569 ( .A(n46852), .B(n46853), .Z(n46848) );
  AND U46570 ( .A(n46854), .B(n46855), .Z(n46853) );
  XNOR U46571 ( .A(p_input[1967]), .B(n46852), .Z(n46855) );
  XNOR U46572 ( .A(n46852), .B(n46529), .Z(n46854) );
  IV U46573 ( .A(p_input[1935]), .Z(n46529) );
  XOR U46574 ( .A(n46856), .B(n46857), .Z(n46852) );
  AND U46575 ( .A(n46858), .B(n46859), .Z(n46857) );
  XNOR U46576 ( .A(p_input[1966]), .B(n46856), .Z(n46859) );
  XNOR U46577 ( .A(n46856), .B(n46538), .Z(n46858) );
  IV U46578 ( .A(p_input[1934]), .Z(n46538) );
  XOR U46579 ( .A(n46860), .B(n46861), .Z(n46856) );
  AND U46580 ( .A(n46862), .B(n46863), .Z(n46861) );
  XNOR U46581 ( .A(p_input[1965]), .B(n46860), .Z(n46863) );
  XNOR U46582 ( .A(n46860), .B(n46547), .Z(n46862) );
  IV U46583 ( .A(p_input[1933]), .Z(n46547) );
  XOR U46584 ( .A(n46864), .B(n46865), .Z(n46860) );
  AND U46585 ( .A(n46866), .B(n46867), .Z(n46865) );
  XNOR U46586 ( .A(p_input[1964]), .B(n46864), .Z(n46867) );
  XNOR U46587 ( .A(n46864), .B(n46556), .Z(n46866) );
  IV U46588 ( .A(p_input[1932]), .Z(n46556) );
  XOR U46589 ( .A(n46868), .B(n46869), .Z(n46864) );
  AND U46590 ( .A(n46870), .B(n46871), .Z(n46869) );
  XNOR U46591 ( .A(p_input[1963]), .B(n46868), .Z(n46871) );
  XNOR U46592 ( .A(n46868), .B(n46565), .Z(n46870) );
  IV U46593 ( .A(p_input[1931]), .Z(n46565) );
  XOR U46594 ( .A(n46872), .B(n46873), .Z(n46868) );
  AND U46595 ( .A(n46874), .B(n46875), .Z(n46873) );
  XNOR U46596 ( .A(p_input[1962]), .B(n46872), .Z(n46875) );
  XNOR U46597 ( .A(n46872), .B(n46574), .Z(n46874) );
  IV U46598 ( .A(p_input[1930]), .Z(n46574) );
  XOR U46599 ( .A(n46876), .B(n46877), .Z(n46872) );
  AND U46600 ( .A(n46878), .B(n46879), .Z(n46877) );
  XNOR U46601 ( .A(p_input[1961]), .B(n46876), .Z(n46879) );
  XNOR U46602 ( .A(n46876), .B(n46583), .Z(n46878) );
  IV U46603 ( .A(p_input[1929]), .Z(n46583) );
  XOR U46604 ( .A(n46880), .B(n46881), .Z(n46876) );
  AND U46605 ( .A(n46882), .B(n46883), .Z(n46881) );
  XNOR U46606 ( .A(p_input[1960]), .B(n46880), .Z(n46883) );
  XNOR U46607 ( .A(n46880), .B(n46592), .Z(n46882) );
  IV U46608 ( .A(p_input[1928]), .Z(n46592) );
  XOR U46609 ( .A(n46884), .B(n46885), .Z(n46880) );
  AND U46610 ( .A(n46886), .B(n46887), .Z(n46885) );
  XNOR U46611 ( .A(p_input[1959]), .B(n46884), .Z(n46887) );
  XNOR U46612 ( .A(n46884), .B(n46601), .Z(n46886) );
  IV U46613 ( .A(p_input[1927]), .Z(n46601) );
  XOR U46614 ( .A(n46888), .B(n46889), .Z(n46884) );
  AND U46615 ( .A(n46890), .B(n46891), .Z(n46889) );
  XNOR U46616 ( .A(p_input[1958]), .B(n46888), .Z(n46891) );
  XNOR U46617 ( .A(n46888), .B(n46610), .Z(n46890) );
  IV U46618 ( .A(p_input[1926]), .Z(n46610) );
  XOR U46619 ( .A(n46892), .B(n46893), .Z(n46888) );
  AND U46620 ( .A(n46894), .B(n46895), .Z(n46893) );
  XNOR U46621 ( .A(p_input[1957]), .B(n46892), .Z(n46895) );
  XNOR U46622 ( .A(n46892), .B(n46619), .Z(n46894) );
  IV U46623 ( .A(p_input[1925]), .Z(n46619) );
  XOR U46624 ( .A(n46896), .B(n46897), .Z(n46892) );
  AND U46625 ( .A(n46898), .B(n46899), .Z(n46897) );
  XNOR U46626 ( .A(p_input[1956]), .B(n46896), .Z(n46899) );
  XNOR U46627 ( .A(n46896), .B(n46628), .Z(n46898) );
  IV U46628 ( .A(p_input[1924]), .Z(n46628) );
  XOR U46629 ( .A(n46900), .B(n46901), .Z(n46896) );
  AND U46630 ( .A(n46902), .B(n46903), .Z(n46901) );
  XNOR U46631 ( .A(p_input[1955]), .B(n46900), .Z(n46903) );
  XNOR U46632 ( .A(n46900), .B(n46637), .Z(n46902) );
  IV U46633 ( .A(p_input[1923]), .Z(n46637) );
  XOR U46634 ( .A(n46904), .B(n46905), .Z(n46900) );
  AND U46635 ( .A(n46906), .B(n46907), .Z(n46905) );
  XNOR U46636 ( .A(p_input[1954]), .B(n46904), .Z(n46907) );
  XNOR U46637 ( .A(n46904), .B(n46646), .Z(n46906) );
  IV U46638 ( .A(p_input[1922]), .Z(n46646) );
  XNOR U46639 ( .A(n46908), .B(n46909), .Z(n46904) );
  AND U46640 ( .A(n46910), .B(n46911), .Z(n46909) );
  XOR U46641 ( .A(p_input[1953]), .B(n46908), .Z(n46911) );
  XNOR U46642 ( .A(p_input[1921]), .B(n46908), .Z(n46910) );
  AND U46643 ( .A(p_input[1952]), .B(n46912), .Z(n46908) );
  IV U46644 ( .A(p_input[1920]), .Z(n46912) );
  XOR U46645 ( .A(n46913), .B(n46914), .Z(n46002) );
  AND U46646 ( .A(n621), .B(n46915), .Z(n46914) );
  XNOR U46647 ( .A(n46916), .B(n46913), .Z(n46915) );
  XOR U46648 ( .A(n46917), .B(n46918), .Z(n621) );
  AND U46649 ( .A(n46919), .B(n46920), .Z(n46918) );
  XNOR U46650 ( .A(n46017), .B(n46917), .Z(n46920) );
  AND U46651 ( .A(p_input[1919]), .B(p_input[1887]), .Z(n46017) );
  XNOR U46652 ( .A(n46917), .B(n46014), .Z(n46919) );
  IV U46653 ( .A(n46921), .Z(n46014) );
  AND U46654 ( .A(p_input[1823]), .B(p_input[1855]), .Z(n46921) );
  XOR U46655 ( .A(n46922), .B(n46923), .Z(n46917) );
  AND U46656 ( .A(n46924), .B(n46925), .Z(n46923) );
  XOR U46657 ( .A(n46922), .B(n46029), .Z(n46925) );
  XNOR U46658 ( .A(p_input[1886]), .B(n46926), .Z(n46029) );
  AND U46659 ( .A(n943), .B(n46927), .Z(n46926) );
  XOR U46660 ( .A(p_input[1918]), .B(p_input[1886]), .Z(n46927) );
  XNOR U46661 ( .A(n46026), .B(n46922), .Z(n46924) );
  XOR U46662 ( .A(n46928), .B(n46929), .Z(n46026) );
  AND U46663 ( .A(n940), .B(n46930), .Z(n46929) );
  XOR U46664 ( .A(p_input[1854]), .B(p_input[1822]), .Z(n46930) );
  XOR U46665 ( .A(n46931), .B(n46932), .Z(n46922) );
  AND U46666 ( .A(n46933), .B(n46934), .Z(n46932) );
  XOR U46667 ( .A(n46931), .B(n46041), .Z(n46934) );
  XNOR U46668 ( .A(p_input[1885]), .B(n46935), .Z(n46041) );
  AND U46669 ( .A(n943), .B(n46936), .Z(n46935) );
  XOR U46670 ( .A(p_input[1917]), .B(p_input[1885]), .Z(n46936) );
  XNOR U46671 ( .A(n46038), .B(n46931), .Z(n46933) );
  XOR U46672 ( .A(n46937), .B(n46938), .Z(n46038) );
  AND U46673 ( .A(n940), .B(n46939), .Z(n46938) );
  XOR U46674 ( .A(p_input[1853]), .B(p_input[1821]), .Z(n46939) );
  XOR U46675 ( .A(n46940), .B(n46941), .Z(n46931) );
  AND U46676 ( .A(n46942), .B(n46943), .Z(n46941) );
  XOR U46677 ( .A(n46940), .B(n46053), .Z(n46943) );
  XNOR U46678 ( .A(p_input[1884]), .B(n46944), .Z(n46053) );
  AND U46679 ( .A(n943), .B(n46945), .Z(n46944) );
  XOR U46680 ( .A(p_input[1916]), .B(p_input[1884]), .Z(n46945) );
  XNOR U46681 ( .A(n46050), .B(n46940), .Z(n46942) );
  XOR U46682 ( .A(n46946), .B(n46947), .Z(n46050) );
  AND U46683 ( .A(n940), .B(n46948), .Z(n46947) );
  XOR U46684 ( .A(p_input[1852]), .B(p_input[1820]), .Z(n46948) );
  XOR U46685 ( .A(n46949), .B(n46950), .Z(n46940) );
  AND U46686 ( .A(n46951), .B(n46952), .Z(n46950) );
  XOR U46687 ( .A(n46949), .B(n46065), .Z(n46952) );
  XNOR U46688 ( .A(p_input[1883]), .B(n46953), .Z(n46065) );
  AND U46689 ( .A(n943), .B(n46954), .Z(n46953) );
  XOR U46690 ( .A(p_input[1915]), .B(p_input[1883]), .Z(n46954) );
  XNOR U46691 ( .A(n46062), .B(n46949), .Z(n46951) );
  XOR U46692 ( .A(n46955), .B(n46956), .Z(n46062) );
  AND U46693 ( .A(n940), .B(n46957), .Z(n46956) );
  XOR U46694 ( .A(p_input[1851]), .B(p_input[1819]), .Z(n46957) );
  XOR U46695 ( .A(n46958), .B(n46959), .Z(n46949) );
  AND U46696 ( .A(n46960), .B(n46961), .Z(n46959) );
  XOR U46697 ( .A(n46958), .B(n46077), .Z(n46961) );
  XNOR U46698 ( .A(p_input[1882]), .B(n46962), .Z(n46077) );
  AND U46699 ( .A(n943), .B(n46963), .Z(n46962) );
  XOR U46700 ( .A(p_input[1914]), .B(p_input[1882]), .Z(n46963) );
  XNOR U46701 ( .A(n46074), .B(n46958), .Z(n46960) );
  XOR U46702 ( .A(n46964), .B(n46965), .Z(n46074) );
  AND U46703 ( .A(n940), .B(n46966), .Z(n46965) );
  XOR U46704 ( .A(p_input[1850]), .B(p_input[1818]), .Z(n46966) );
  XOR U46705 ( .A(n46967), .B(n46968), .Z(n46958) );
  AND U46706 ( .A(n46969), .B(n46970), .Z(n46968) );
  XOR U46707 ( .A(n46967), .B(n46089), .Z(n46970) );
  XNOR U46708 ( .A(p_input[1881]), .B(n46971), .Z(n46089) );
  AND U46709 ( .A(n943), .B(n46972), .Z(n46971) );
  XOR U46710 ( .A(p_input[1913]), .B(p_input[1881]), .Z(n46972) );
  XNOR U46711 ( .A(n46086), .B(n46967), .Z(n46969) );
  XOR U46712 ( .A(n46973), .B(n46974), .Z(n46086) );
  AND U46713 ( .A(n940), .B(n46975), .Z(n46974) );
  XOR U46714 ( .A(p_input[1849]), .B(p_input[1817]), .Z(n46975) );
  XOR U46715 ( .A(n46976), .B(n46977), .Z(n46967) );
  AND U46716 ( .A(n46978), .B(n46979), .Z(n46977) );
  XOR U46717 ( .A(n46976), .B(n46101), .Z(n46979) );
  XNOR U46718 ( .A(p_input[1880]), .B(n46980), .Z(n46101) );
  AND U46719 ( .A(n943), .B(n46981), .Z(n46980) );
  XOR U46720 ( .A(p_input[1912]), .B(p_input[1880]), .Z(n46981) );
  XNOR U46721 ( .A(n46098), .B(n46976), .Z(n46978) );
  XOR U46722 ( .A(n46982), .B(n46983), .Z(n46098) );
  AND U46723 ( .A(n940), .B(n46984), .Z(n46983) );
  XOR U46724 ( .A(p_input[1848]), .B(p_input[1816]), .Z(n46984) );
  XOR U46725 ( .A(n46985), .B(n46986), .Z(n46976) );
  AND U46726 ( .A(n46987), .B(n46988), .Z(n46986) );
  XOR U46727 ( .A(n46985), .B(n46113), .Z(n46988) );
  XNOR U46728 ( .A(p_input[1879]), .B(n46989), .Z(n46113) );
  AND U46729 ( .A(n943), .B(n46990), .Z(n46989) );
  XOR U46730 ( .A(p_input[1911]), .B(p_input[1879]), .Z(n46990) );
  XNOR U46731 ( .A(n46110), .B(n46985), .Z(n46987) );
  XOR U46732 ( .A(n46991), .B(n46992), .Z(n46110) );
  AND U46733 ( .A(n940), .B(n46993), .Z(n46992) );
  XOR U46734 ( .A(p_input[1847]), .B(p_input[1815]), .Z(n46993) );
  XOR U46735 ( .A(n46994), .B(n46995), .Z(n46985) );
  AND U46736 ( .A(n46996), .B(n46997), .Z(n46995) );
  XOR U46737 ( .A(n46994), .B(n46125), .Z(n46997) );
  XNOR U46738 ( .A(p_input[1878]), .B(n46998), .Z(n46125) );
  AND U46739 ( .A(n943), .B(n46999), .Z(n46998) );
  XOR U46740 ( .A(p_input[1910]), .B(p_input[1878]), .Z(n46999) );
  XNOR U46741 ( .A(n46122), .B(n46994), .Z(n46996) );
  XOR U46742 ( .A(n47000), .B(n47001), .Z(n46122) );
  AND U46743 ( .A(n940), .B(n47002), .Z(n47001) );
  XOR U46744 ( .A(p_input[1846]), .B(p_input[1814]), .Z(n47002) );
  XOR U46745 ( .A(n47003), .B(n47004), .Z(n46994) );
  AND U46746 ( .A(n47005), .B(n47006), .Z(n47004) );
  XOR U46747 ( .A(n47003), .B(n46137), .Z(n47006) );
  XNOR U46748 ( .A(p_input[1877]), .B(n47007), .Z(n46137) );
  AND U46749 ( .A(n943), .B(n47008), .Z(n47007) );
  XOR U46750 ( .A(p_input[1909]), .B(p_input[1877]), .Z(n47008) );
  XNOR U46751 ( .A(n46134), .B(n47003), .Z(n47005) );
  XOR U46752 ( .A(n47009), .B(n47010), .Z(n46134) );
  AND U46753 ( .A(n940), .B(n47011), .Z(n47010) );
  XOR U46754 ( .A(p_input[1845]), .B(p_input[1813]), .Z(n47011) );
  XOR U46755 ( .A(n47012), .B(n47013), .Z(n47003) );
  AND U46756 ( .A(n47014), .B(n47015), .Z(n47013) );
  XOR U46757 ( .A(n47012), .B(n46149), .Z(n47015) );
  XNOR U46758 ( .A(p_input[1876]), .B(n47016), .Z(n46149) );
  AND U46759 ( .A(n943), .B(n47017), .Z(n47016) );
  XOR U46760 ( .A(p_input[1908]), .B(p_input[1876]), .Z(n47017) );
  XNOR U46761 ( .A(n46146), .B(n47012), .Z(n47014) );
  XOR U46762 ( .A(n47018), .B(n47019), .Z(n46146) );
  AND U46763 ( .A(n940), .B(n47020), .Z(n47019) );
  XOR U46764 ( .A(p_input[1844]), .B(p_input[1812]), .Z(n47020) );
  XOR U46765 ( .A(n47021), .B(n47022), .Z(n47012) );
  AND U46766 ( .A(n47023), .B(n47024), .Z(n47022) );
  XOR U46767 ( .A(n47021), .B(n46161), .Z(n47024) );
  XNOR U46768 ( .A(p_input[1875]), .B(n47025), .Z(n46161) );
  AND U46769 ( .A(n943), .B(n47026), .Z(n47025) );
  XOR U46770 ( .A(p_input[1907]), .B(p_input[1875]), .Z(n47026) );
  XNOR U46771 ( .A(n46158), .B(n47021), .Z(n47023) );
  XOR U46772 ( .A(n47027), .B(n47028), .Z(n46158) );
  AND U46773 ( .A(n940), .B(n47029), .Z(n47028) );
  XOR U46774 ( .A(p_input[1843]), .B(p_input[1811]), .Z(n47029) );
  XOR U46775 ( .A(n47030), .B(n47031), .Z(n47021) );
  AND U46776 ( .A(n47032), .B(n47033), .Z(n47031) );
  XOR U46777 ( .A(n47030), .B(n46173), .Z(n47033) );
  XNOR U46778 ( .A(p_input[1874]), .B(n47034), .Z(n46173) );
  AND U46779 ( .A(n943), .B(n47035), .Z(n47034) );
  XOR U46780 ( .A(p_input[1906]), .B(p_input[1874]), .Z(n47035) );
  XNOR U46781 ( .A(n46170), .B(n47030), .Z(n47032) );
  XOR U46782 ( .A(n47036), .B(n47037), .Z(n46170) );
  AND U46783 ( .A(n940), .B(n47038), .Z(n47037) );
  XOR U46784 ( .A(p_input[1842]), .B(p_input[1810]), .Z(n47038) );
  XOR U46785 ( .A(n47039), .B(n47040), .Z(n47030) );
  AND U46786 ( .A(n47041), .B(n47042), .Z(n47040) );
  XOR U46787 ( .A(n47039), .B(n46185), .Z(n47042) );
  XNOR U46788 ( .A(p_input[1873]), .B(n47043), .Z(n46185) );
  AND U46789 ( .A(n943), .B(n47044), .Z(n47043) );
  XOR U46790 ( .A(p_input[1905]), .B(p_input[1873]), .Z(n47044) );
  XNOR U46791 ( .A(n46182), .B(n47039), .Z(n47041) );
  XOR U46792 ( .A(n47045), .B(n47046), .Z(n46182) );
  AND U46793 ( .A(n940), .B(n47047), .Z(n47046) );
  XOR U46794 ( .A(p_input[1841]), .B(p_input[1809]), .Z(n47047) );
  XOR U46795 ( .A(n47048), .B(n47049), .Z(n47039) );
  AND U46796 ( .A(n47050), .B(n47051), .Z(n47049) );
  XOR U46797 ( .A(n47048), .B(n46197), .Z(n47051) );
  XNOR U46798 ( .A(p_input[1872]), .B(n47052), .Z(n46197) );
  AND U46799 ( .A(n943), .B(n47053), .Z(n47052) );
  XOR U46800 ( .A(p_input[1904]), .B(p_input[1872]), .Z(n47053) );
  XNOR U46801 ( .A(n46194), .B(n47048), .Z(n47050) );
  XOR U46802 ( .A(n47054), .B(n47055), .Z(n46194) );
  AND U46803 ( .A(n940), .B(n47056), .Z(n47055) );
  XOR U46804 ( .A(p_input[1840]), .B(p_input[1808]), .Z(n47056) );
  XOR U46805 ( .A(n47057), .B(n47058), .Z(n47048) );
  AND U46806 ( .A(n47059), .B(n47060), .Z(n47058) );
  XOR U46807 ( .A(n47057), .B(n46209), .Z(n47060) );
  XNOR U46808 ( .A(p_input[1871]), .B(n47061), .Z(n46209) );
  AND U46809 ( .A(n943), .B(n47062), .Z(n47061) );
  XOR U46810 ( .A(p_input[1903]), .B(p_input[1871]), .Z(n47062) );
  XNOR U46811 ( .A(n46206), .B(n47057), .Z(n47059) );
  XOR U46812 ( .A(n47063), .B(n47064), .Z(n46206) );
  AND U46813 ( .A(n940), .B(n47065), .Z(n47064) );
  XOR U46814 ( .A(p_input[1839]), .B(p_input[1807]), .Z(n47065) );
  XOR U46815 ( .A(n47066), .B(n47067), .Z(n47057) );
  AND U46816 ( .A(n47068), .B(n47069), .Z(n47067) );
  XOR U46817 ( .A(n47066), .B(n46221), .Z(n47069) );
  XNOR U46818 ( .A(p_input[1870]), .B(n47070), .Z(n46221) );
  AND U46819 ( .A(n943), .B(n47071), .Z(n47070) );
  XOR U46820 ( .A(p_input[1902]), .B(p_input[1870]), .Z(n47071) );
  XNOR U46821 ( .A(n46218), .B(n47066), .Z(n47068) );
  XOR U46822 ( .A(n47072), .B(n47073), .Z(n46218) );
  AND U46823 ( .A(n940), .B(n47074), .Z(n47073) );
  XOR U46824 ( .A(p_input[1838]), .B(p_input[1806]), .Z(n47074) );
  XOR U46825 ( .A(n47075), .B(n47076), .Z(n47066) );
  AND U46826 ( .A(n47077), .B(n47078), .Z(n47076) );
  XOR U46827 ( .A(n47075), .B(n46233), .Z(n47078) );
  XNOR U46828 ( .A(p_input[1869]), .B(n47079), .Z(n46233) );
  AND U46829 ( .A(n943), .B(n47080), .Z(n47079) );
  XOR U46830 ( .A(p_input[1901]), .B(p_input[1869]), .Z(n47080) );
  XNOR U46831 ( .A(n46230), .B(n47075), .Z(n47077) );
  XOR U46832 ( .A(n47081), .B(n47082), .Z(n46230) );
  AND U46833 ( .A(n940), .B(n47083), .Z(n47082) );
  XOR U46834 ( .A(p_input[1837]), .B(p_input[1805]), .Z(n47083) );
  XOR U46835 ( .A(n47084), .B(n47085), .Z(n47075) );
  AND U46836 ( .A(n47086), .B(n47087), .Z(n47085) );
  XOR U46837 ( .A(n47084), .B(n46245), .Z(n47087) );
  XNOR U46838 ( .A(p_input[1868]), .B(n47088), .Z(n46245) );
  AND U46839 ( .A(n943), .B(n47089), .Z(n47088) );
  XOR U46840 ( .A(p_input[1900]), .B(p_input[1868]), .Z(n47089) );
  XNOR U46841 ( .A(n46242), .B(n47084), .Z(n47086) );
  XOR U46842 ( .A(n47090), .B(n47091), .Z(n46242) );
  AND U46843 ( .A(n940), .B(n47092), .Z(n47091) );
  XOR U46844 ( .A(p_input[1836]), .B(p_input[1804]), .Z(n47092) );
  XOR U46845 ( .A(n47093), .B(n47094), .Z(n47084) );
  AND U46846 ( .A(n47095), .B(n47096), .Z(n47094) );
  XOR U46847 ( .A(n47093), .B(n46257), .Z(n47096) );
  XNOR U46848 ( .A(p_input[1867]), .B(n47097), .Z(n46257) );
  AND U46849 ( .A(n943), .B(n47098), .Z(n47097) );
  XOR U46850 ( .A(p_input[1899]), .B(p_input[1867]), .Z(n47098) );
  XNOR U46851 ( .A(n46254), .B(n47093), .Z(n47095) );
  XOR U46852 ( .A(n47099), .B(n47100), .Z(n46254) );
  AND U46853 ( .A(n940), .B(n47101), .Z(n47100) );
  XOR U46854 ( .A(p_input[1835]), .B(p_input[1803]), .Z(n47101) );
  XOR U46855 ( .A(n47102), .B(n47103), .Z(n47093) );
  AND U46856 ( .A(n47104), .B(n47105), .Z(n47103) );
  XOR U46857 ( .A(n47102), .B(n46269), .Z(n47105) );
  XNOR U46858 ( .A(p_input[1866]), .B(n47106), .Z(n46269) );
  AND U46859 ( .A(n943), .B(n47107), .Z(n47106) );
  XOR U46860 ( .A(p_input[1898]), .B(p_input[1866]), .Z(n47107) );
  XNOR U46861 ( .A(n46266), .B(n47102), .Z(n47104) );
  XOR U46862 ( .A(n47108), .B(n47109), .Z(n46266) );
  AND U46863 ( .A(n940), .B(n47110), .Z(n47109) );
  XOR U46864 ( .A(p_input[1834]), .B(p_input[1802]), .Z(n47110) );
  XOR U46865 ( .A(n47111), .B(n47112), .Z(n47102) );
  AND U46866 ( .A(n47113), .B(n47114), .Z(n47112) );
  XOR U46867 ( .A(n47111), .B(n46281), .Z(n47114) );
  XNOR U46868 ( .A(p_input[1865]), .B(n47115), .Z(n46281) );
  AND U46869 ( .A(n943), .B(n47116), .Z(n47115) );
  XOR U46870 ( .A(p_input[1897]), .B(p_input[1865]), .Z(n47116) );
  XNOR U46871 ( .A(n46278), .B(n47111), .Z(n47113) );
  XOR U46872 ( .A(n47117), .B(n47118), .Z(n46278) );
  AND U46873 ( .A(n940), .B(n47119), .Z(n47118) );
  XOR U46874 ( .A(p_input[1833]), .B(p_input[1801]), .Z(n47119) );
  XOR U46875 ( .A(n47120), .B(n47121), .Z(n47111) );
  AND U46876 ( .A(n47122), .B(n47123), .Z(n47121) );
  XOR U46877 ( .A(n47120), .B(n46293), .Z(n47123) );
  XNOR U46878 ( .A(p_input[1864]), .B(n47124), .Z(n46293) );
  AND U46879 ( .A(n943), .B(n47125), .Z(n47124) );
  XOR U46880 ( .A(p_input[1896]), .B(p_input[1864]), .Z(n47125) );
  XNOR U46881 ( .A(n46290), .B(n47120), .Z(n47122) );
  XOR U46882 ( .A(n47126), .B(n47127), .Z(n46290) );
  AND U46883 ( .A(n940), .B(n47128), .Z(n47127) );
  XOR U46884 ( .A(p_input[1832]), .B(p_input[1800]), .Z(n47128) );
  XOR U46885 ( .A(n47129), .B(n47130), .Z(n47120) );
  AND U46886 ( .A(n47131), .B(n47132), .Z(n47130) );
  XOR U46887 ( .A(n47129), .B(n46305), .Z(n47132) );
  XNOR U46888 ( .A(p_input[1863]), .B(n47133), .Z(n46305) );
  AND U46889 ( .A(n943), .B(n47134), .Z(n47133) );
  XOR U46890 ( .A(p_input[1895]), .B(p_input[1863]), .Z(n47134) );
  XNOR U46891 ( .A(n46302), .B(n47129), .Z(n47131) );
  XOR U46892 ( .A(n47135), .B(n47136), .Z(n46302) );
  AND U46893 ( .A(n940), .B(n47137), .Z(n47136) );
  XOR U46894 ( .A(p_input[1831]), .B(p_input[1799]), .Z(n47137) );
  XOR U46895 ( .A(n47138), .B(n47139), .Z(n47129) );
  AND U46896 ( .A(n47140), .B(n47141), .Z(n47139) );
  XOR U46897 ( .A(n47138), .B(n46317), .Z(n47141) );
  XNOR U46898 ( .A(p_input[1862]), .B(n47142), .Z(n46317) );
  AND U46899 ( .A(n943), .B(n47143), .Z(n47142) );
  XOR U46900 ( .A(p_input[1894]), .B(p_input[1862]), .Z(n47143) );
  XNOR U46901 ( .A(n46314), .B(n47138), .Z(n47140) );
  XOR U46902 ( .A(n47144), .B(n47145), .Z(n46314) );
  AND U46903 ( .A(n940), .B(n47146), .Z(n47145) );
  XOR U46904 ( .A(p_input[1830]), .B(p_input[1798]), .Z(n47146) );
  XOR U46905 ( .A(n47147), .B(n47148), .Z(n47138) );
  AND U46906 ( .A(n47149), .B(n47150), .Z(n47148) );
  XOR U46907 ( .A(n47147), .B(n46329), .Z(n47150) );
  XNOR U46908 ( .A(p_input[1861]), .B(n47151), .Z(n46329) );
  AND U46909 ( .A(n943), .B(n47152), .Z(n47151) );
  XOR U46910 ( .A(p_input[1893]), .B(p_input[1861]), .Z(n47152) );
  XNOR U46911 ( .A(n46326), .B(n47147), .Z(n47149) );
  XOR U46912 ( .A(n47153), .B(n47154), .Z(n46326) );
  AND U46913 ( .A(n940), .B(n47155), .Z(n47154) );
  XOR U46914 ( .A(p_input[1829]), .B(p_input[1797]), .Z(n47155) );
  XOR U46915 ( .A(n47156), .B(n47157), .Z(n47147) );
  AND U46916 ( .A(n47158), .B(n47159), .Z(n47157) );
  XOR U46917 ( .A(n47156), .B(n46341), .Z(n47159) );
  XNOR U46918 ( .A(p_input[1860]), .B(n47160), .Z(n46341) );
  AND U46919 ( .A(n943), .B(n47161), .Z(n47160) );
  XOR U46920 ( .A(p_input[1892]), .B(p_input[1860]), .Z(n47161) );
  XNOR U46921 ( .A(n46338), .B(n47156), .Z(n47158) );
  XOR U46922 ( .A(n47162), .B(n47163), .Z(n46338) );
  AND U46923 ( .A(n940), .B(n47164), .Z(n47163) );
  XOR U46924 ( .A(p_input[1828]), .B(p_input[1796]), .Z(n47164) );
  XOR U46925 ( .A(n47165), .B(n47166), .Z(n47156) );
  AND U46926 ( .A(n47167), .B(n47168), .Z(n47166) );
  XOR U46927 ( .A(n47165), .B(n46353), .Z(n47168) );
  XNOR U46928 ( .A(p_input[1859]), .B(n47169), .Z(n46353) );
  AND U46929 ( .A(n943), .B(n47170), .Z(n47169) );
  XOR U46930 ( .A(p_input[1891]), .B(p_input[1859]), .Z(n47170) );
  XNOR U46931 ( .A(n46350), .B(n47165), .Z(n47167) );
  XOR U46932 ( .A(n47171), .B(n47172), .Z(n46350) );
  AND U46933 ( .A(n940), .B(n47173), .Z(n47172) );
  XOR U46934 ( .A(p_input[1827]), .B(p_input[1795]), .Z(n47173) );
  XOR U46935 ( .A(n47174), .B(n47175), .Z(n47165) );
  AND U46936 ( .A(n47176), .B(n47177), .Z(n47175) );
  XOR U46937 ( .A(n47174), .B(n46365), .Z(n47177) );
  XNOR U46938 ( .A(p_input[1858]), .B(n47178), .Z(n46365) );
  AND U46939 ( .A(n943), .B(n47179), .Z(n47178) );
  XOR U46940 ( .A(p_input[1890]), .B(p_input[1858]), .Z(n47179) );
  XNOR U46941 ( .A(n46362), .B(n47174), .Z(n47176) );
  XOR U46942 ( .A(n47180), .B(n47181), .Z(n46362) );
  AND U46943 ( .A(n940), .B(n47182), .Z(n47181) );
  XOR U46944 ( .A(p_input[1826]), .B(p_input[1794]), .Z(n47182) );
  XOR U46945 ( .A(n47183), .B(n47184), .Z(n47174) );
  AND U46946 ( .A(n47185), .B(n47186), .Z(n47184) );
  XNOR U46947 ( .A(n47187), .B(n46378), .Z(n47186) );
  XNOR U46948 ( .A(p_input[1857]), .B(n47188), .Z(n46378) );
  AND U46949 ( .A(n943), .B(n47189), .Z(n47188) );
  XNOR U46950 ( .A(p_input[1889]), .B(n47190), .Z(n47189) );
  IV U46951 ( .A(p_input[1857]), .Z(n47190) );
  XNOR U46952 ( .A(n46375), .B(n47183), .Z(n47185) );
  XNOR U46953 ( .A(p_input[1793]), .B(n47191), .Z(n46375) );
  AND U46954 ( .A(n940), .B(n47192), .Z(n47191) );
  XOR U46955 ( .A(p_input[1825]), .B(p_input[1793]), .Z(n47192) );
  IV U46956 ( .A(n47187), .Z(n47183) );
  AND U46957 ( .A(n46913), .B(n46916), .Z(n47187) );
  XOR U46958 ( .A(p_input[1856]), .B(n47193), .Z(n46916) );
  AND U46959 ( .A(n943), .B(n47194), .Z(n47193) );
  XOR U46960 ( .A(p_input[1888]), .B(p_input[1856]), .Z(n47194) );
  XOR U46961 ( .A(n47195), .B(n47196), .Z(n943) );
  AND U46962 ( .A(n47197), .B(n47198), .Z(n47196) );
  XNOR U46963 ( .A(p_input[1919]), .B(n47195), .Z(n47198) );
  XOR U46964 ( .A(n47195), .B(p_input[1887]), .Z(n47197) );
  XOR U46965 ( .A(n47199), .B(n47200), .Z(n47195) );
  AND U46966 ( .A(n47201), .B(n47202), .Z(n47200) );
  XNOR U46967 ( .A(p_input[1918]), .B(n47199), .Z(n47202) );
  XOR U46968 ( .A(n47199), .B(p_input[1886]), .Z(n47201) );
  XOR U46969 ( .A(n47203), .B(n47204), .Z(n47199) );
  AND U46970 ( .A(n47205), .B(n47206), .Z(n47204) );
  XNOR U46971 ( .A(p_input[1917]), .B(n47203), .Z(n47206) );
  XOR U46972 ( .A(n47203), .B(p_input[1885]), .Z(n47205) );
  XOR U46973 ( .A(n47207), .B(n47208), .Z(n47203) );
  AND U46974 ( .A(n47209), .B(n47210), .Z(n47208) );
  XNOR U46975 ( .A(p_input[1916]), .B(n47207), .Z(n47210) );
  XOR U46976 ( .A(n47207), .B(p_input[1884]), .Z(n47209) );
  XOR U46977 ( .A(n47211), .B(n47212), .Z(n47207) );
  AND U46978 ( .A(n47213), .B(n47214), .Z(n47212) );
  XNOR U46979 ( .A(p_input[1915]), .B(n47211), .Z(n47214) );
  XOR U46980 ( .A(n47211), .B(p_input[1883]), .Z(n47213) );
  XOR U46981 ( .A(n47215), .B(n47216), .Z(n47211) );
  AND U46982 ( .A(n47217), .B(n47218), .Z(n47216) );
  XNOR U46983 ( .A(p_input[1914]), .B(n47215), .Z(n47218) );
  XOR U46984 ( .A(n47215), .B(p_input[1882]), .Z(n47217) );
  XOR U46985 ( .A(n47219), .B(n47220), .Z(n47215) );
  AND U46986 ( .A(n47221), .B(n47222), .Z(n47220) );
  XNOR U46987 ( .A(p_input[1913]), .B(n47219), .Z(n47222) );
  XOR U46988 ( .A(n47219), .B(p_input[1881]), .Z(n47221) );
  XOR U46989 ( .A(n47223), .B(n47224), .Z(n47219) );
  AND U46990 ( .A(n47225), .B(n47226), .Z(n47224) );
  XNOR U46991 ( .A(p_input[1912]), .B(n47223), .Z(n47226) );
  XOR U46992 ( .A(n47223), .B(p_input[1880]), .Z(n47225) );
  XOR U46993 ( .A(n47227), .B(n47228), .Z(n47223) );
  AND U46994 ( .A(n47229), .B(n47230), .Z(n47228) );
  XNOR U46995 ( .A(p_input[1911]), .B(n47227), .Z(n47230) );
  XOR U46996 ( .A(n47227), .B(p_input[1879]), .Z(n47229) );
  XOR U46997 ( .A(n47231), .B(n47232), .Z(n47227) );
  AND U46998 ( .A(n47233), .B(n47234), .Z(n47232) );
  XNOR U46999 ( .A(p_input[1910]), .B(n47231), .Z(n47234) );
  XOR U47000 ( .A(n47231), .B(p_input[1878]), .Z(n47233) );
  XOR U47001 ( .A(n47235), .B(n47236), .Z(n47231) );
  AND U47002 ( .A(n47237), .B(n47238), .Z(n47236) );
  XNOR U47003 ( .A(p_input[1909]), .B(n47235), .Z(n47238) );
  XOR U47004 ( .A(n47235), .B(p_input[1877]), .Z(n47237) );
  XOR U47005 ( .A(n47239), .B(n47240), .Z(n47235) );
  AND U47006 ( .A(n47241), .B(n47242), .Z(n47240) );
  XNOR U47007 ( .A(p_input[1908]), .B(n47239), .Z(n47242) );
  XOR U47008 ( .A(n47239), .B(p_input[1876]), .Z(n47241) );
  XOR U47009 ( .A(n47243), .B(n47244), .Z(n47239) );
  AND U47010 ( .A(n47245), .B(n47246), .Z(n47244) );
  XNOR U47011 ( .A(p_input[1907]), .B(n47243), .Z(n47246) );
  XOR U47012 ( .A(n47243), .B(p_input[1875]), .Z(n47245) );
  XOR U47013 ( .A(n47247), .B(n47248), .Z(n47243) );
  AND U47014 ( .A(n47249), .B(n47250), .Z(n47248) );
  XNOR U47015 ( .A(p_input[1906]), .B(n47247), .Z(n47250) );
  XOR U47016 ( .A(n47247), .B(p_input[1874]), .Z(n47249) );
  XOR U47017 ( .A(n47251), .B(n47252), .Z(n47247) );
  AND U47018 ( .A(n47253), .B(n47254), .Z(n47252) );
  XNOR U47019 ( .A(p_input[1905]), .B(n47251), .Z(n47254) );
  XOR U47020 ( .A(n47251), .B(p_input[1873]), .Z(n47253) );
  XOR U47021 ( .A(n47255), .B(n47256), .Z(n47251) );
  AND U47022 ( .A(n47257), .B(n47258), .Z(n47256) );
  XNOR U47023 ( .A(p_input[1904]), .B(n47255), .Z(n47258) );
  XOR U47024 ( .A(n47255), .B(p_input[1872]), .Z(n47257) );
  XOR U47025 ( .A(n47259), .B(n47260), .Z(n47255) );
  AND U47026 ( .A(n47261), .B(n47262), .Z(n47260) );
  XNOR U47027 ( .A(p_input[1903]), .B(n47259), .Z(n47262) );
  XOR U47028 ( .A(n47259), .B(p_input[1871]), .Z(n47261) );
  XOR U47029 ( .A(n47263), .B(n47264), .Z(n47259) );
  AND U47030 ( .A(n47265), .B(n47266), .Z(n47264) );
  XNOR U47031 ( .A(p_input[1902]), .B(n47263), .Z(n47266) );
  XOR U47032 ( .A(n47263), .B(p_input[1870]), .Z(n47265) );
  XOR U47033 ( .A(n47267), .B(n47268), .Z(n47263) );
  AND U47034 ( .A(n47269), .B(n47270), .Z(n47268) );
  XNOR U47035 ( .A(p_input[1901]), .B(n47267), .Z(n47270) );
  XOR U47036 ( .A(n47267), .B(p_input[1869]), .Z(n47269) );
  XOR U47037 ( .A(n47271), .B(n47272), .Z(n47267) );
  AND U47038 ( .A(n47273), .B(n47274), .Z(n47272) );
  XNOR U47039 ( .A(p_input[1900]), .B(n47271), .Z(n47274) );
  XOR U47040 ( .A(n47271), .B(p_input[1868]), .Z(n47273) );
  XOR U47041 ( .A(n47275), .B(n47276), .Z(n47271) );
  AND U47042 ( .A(n47277), .B(n47278), .Z(n47276) );
  XNOR U47043 ( .A(p_input[1899]), .B(n47275), .Z(n47278) );
  XOR U47044 ( .A(n47275), .B(p_input[1867]), .Z(n47277) );
  XOR U47045 ( .A(n47279), .B(n47280), .Z(n47275) );
  AND U47046 ( .A(n47281), .B(n47282), .Z(n47280) );
  XNOR U47047 ( .A(p_input[1898]), .B(n47279), .Z(n47282) );
  XOR U47048 ( .A(n47279), .B(p_input[1866]), .Z(n47281) );
  XOR U47049 ( .A(n47283), .B(n47284), .Z(n47279) );
  AND U47050 ( .A(n47285), .B(n47286), .Z(n47284) );
  XNOR U47051 ( .A(p_input[1897]), .B(n47283), .Z(n47286) );
  XOR U47052 ( .A(n47283), .B(p_input[1865]), .Z(n47285) );
  XOR U47053 ( .A(n47287), .B(n47288), .Z(n47283) );
  AND U47054 ( .A(n47289), .B(n47290), .Z(n47288) );
  XNOR U47055 ( .A(p_input[1896]), .B(n47287), .Z(n47290) );
  XOR U47056 ( .A(n47287), .B(p_input[1864]), .Z(n47289) );
  XOR U47057 ( .A(n47291), .B(n47292), .Z(n47287) );
  AND U47058 ( .A(n47293), .B(n47294), .Z(n47292) );
  XNOR U47059 ( .A(p_input[1895]), .B(n47291), .Z(n47294) );
  XOR U47060 ( .A(n47291), .B(p_input[1863]), .Z(n47293) );
  XOR U47061 ( .A(n47295), .B(n47296), .Z(n47291) );
  AND U47062 ( .A(n47297), .B(n47298), .Z(n47296) );
  XNOR U47063 ( .A(p_input[1894]), .B(n47295), .Z(n47298) );
  XOR U47064 ( .A(n47295), .B(p_input[1862]), .Z(n47297) );
  XOR U47065 ( .A(n47299), .B(n47300), .Z(n47295) );
  AND U47066 ( .A(n47301), .B(n47302), .Z(n47300) );
  XNOR U47067 ( .A(p_input[1893]), .B(n47299), .Z(n47302) );
  XOR U47068 ( .A(n47299), .B(p_input[1861]), .Z(n47301) );
  XOR U47069 ( .A(n47303), .B(n47304), .Z(n47299) );
  AND U47070 ( .A(n47305), .B(n47306), .Z(n47304) );
  XNOR U47071 ( .A(p_input[1892]), .B(n47303), .Z(n47306) );
  XOR U47072 ( .A(n47303), .B(p_input[1860]), .Z(n47305) );
  XOR U47073 ( .A(n47307), .B(n47308), .Z(n47303) );
  AND U47074 ( .A(n47309), .B(n47310), .Z(n47308) );
  XNOR U47075 ( .A(p_input[1891]), .B(n47307), .Z(n47310) );
  XOR U47076 ( .A(n47307), .B(p_input[1859]), .Z(n47309) );
  XOR U47077 ( .A(n47311), .B(n47312), .Z(n47307) );
  AND U47078 ( .A(n47313), .B(n47314), .Z(n47312) );
  XNOR U47079 ( .A(p_input[1890]), .B(n47311), .Z(n47314) );
  XOR U47080 ( .A(n47311), .B(p_input[1858]), .Z(n47313) );
  XNOR U47081 ( .A(n47315), .B(n47316), .Z(n47311) );
  AND U47082 ( .A(n47317), .B(n47318), .Z(n47316) );
  XOR U47083 ( .A(p_input[1889]), .B(n47315), .Z(n47318) );
  XNOR U47084 ( .A(p_input[1857]), .B(n47315), .Z(n47317) );
  AND U47085 ( .A(p_input[1888]), .B(n47319), .Z(n47315) );
  IV U47086 ( .A(p_input[1856]), .Z(n47319) );
  XNOR U47087 ( .A(p_input[1792]), .B(n47320), .Z(n46913) );
  AND U47088 ( .A(n940), .B(n47321), .Z(n47320) );
  XOR U47089 ( .A(p_input[1824]), .B(p_input[1792]), .Z(n47321) );
  XOR U47090 ( .A(n47322), .B(n47323), .Z(n940) );
  AND U47091 ( .A(n47324), .B(n47325), .Z(n47323) );
  XNOR U47092 ( .A(p_input[1855]), .B(n47322), .Z(n47325) );
  XOR U47093 ( .A(n47322), .B(p_input[1823]), .Z(n47324) );
  XOR U47094 ( .A(n47326), .B(n47327), .Z(n47322) );
  AND U47095 ( .A(n47328), .B(n47329), .Z(n47327) );
  XNOR U47096 ( .A(p_input[1854]), .B(n47326), .Z(n47329) );
  XNOR U47097 ( .A(n47326), .B(n46928), .Z(n47328) );
  IV U47098 ( .A(p_input[1822]), .Z(n46928) );
  XOR U47099 ( .A(n47330), .B(n47331), .Z(n47326) );
  AND U47100 ( .A(n47332), .B(n47333), .Z(n47331) );
  XNOR U47101 ( .A(p_input[1853]), .B(n47330), .Z(n47333) );
  XNOR U47102 ( .A(n47330), .B(n46937), .Z(n47332) );
  IV U47103 ( .A(p_input[1821]), .Z(n46937) );
  XOR U47104 ( .A(n47334), .B(n47335), .Z(n47330) );
  AND U47105 ( .A(n47336), .B(n47337), .Z(n47335) );
  XNOR U47106 ( .A(p_input[1852]), .B(n47334), .Z(n47337) );
  XNOR U47107 ( .A(n47334), .B(n46946), .Z(n47336) );
  IV U47108 ( .A(p_input[1820]), .Z(n46946) );
  XOR U47109 ( .A(n47338), .B(n47339), .Z(n47334) );
  AND U47110 ( .A(n47340), .B(n47341), .Z(n47339) );
  XNOR U47111 ( .A(p_input[1851]), .B(n47338), .Z(n47341) );
  XNOR U47112 ( .A(n47338), .B(n46955), .Z(n47340) );
  IV U47113 ( .A(p_input[1819]), .Z(n46955) );
  XOR U47114 ( .A(n47342), .B(n47343), .Z(n47338) );
  AND U47115 ( .A(n47344), .B(n47345), .Z(n47343) );
  XNOR U47116 ( .A(p_input[1850]), .B(n47342), .Z(n47345) );
  XNOR U47117 ( .A(n47342), .B(n46964), .Z(n47344) );
  IV U47118 ( .A(p_input[1818]), .Z(n46964) );
  XOR U47119 ( .A(n47346), .B(n47347), .Z(n47342) );
  AND U47120 ( .A(n47348), .B(n47349), .Z(n47347) );
  XNOR U47121 ( .A(p_input[1849]), .B(n47346), .Z(n47349) );
  XNOR U47122 ( .A(n47346), .B(n46973), .Z(n47348) );
  IV U47123 ( .A(p_input[1817]), .Z(n46973) );
  XOR U47124 ( .A(n47350), .B(n47351), .Z(n47346) );
  AND U47125 ( .A(n47352), .B(n47353), .Z(n47351) );
  XNOR U47126 ( .A(p_input[1848]), .B(n47350), .Z(n47353) );
  XNOR U47127 ( .A(n47350), .B(n46982), .Z(n47352) );
  IV U47128 ( .A(p_input[1816]), .Z(n46982) );
  XOR U47129 ( .A(n47354), .B(n47355), .Z(n47350) );
  AND U47130 ( .A(n47356), .B(n47357), .Z(n47355) );
  XNOR U47131 ( .A(p_input[1847]), .B(n47354), .Z(n47357) );
  XNOR U47132 ( .A(n47354), .B(n46991), .Z(n47356) );
  IV U47133 ( .A(p_input[1815]), .Z(n46991) );
  XOR U47134 ( .A(n47358), .B(n47359), .Z(n47354) );
  AND U47135 ( .A(n47360), .B(n47361), .Z(n47359) );
  XNOR U47136 ( .A(p_input[1846]), .B(n47358), .Z(n47361) );
  XNOR U47137 ( .A(n47358), .B(n47000), .Z(n47360) );
  IV U47138 ( .A(p_input[1814]), .Z(n47000) );
  XOR U47139 ( .A(n47362), .B(n47363), .Z(n47358) );
  AND U47140 ( .A(n47364), .B(n47365), .Z(n47363) );
  XNOR U47141 ( .A(p_input[1845]), .B(n47362), .Z(n47365) );
  XNOR U47142 ( .A(n47362), .B(n47009), .Z(n47364) );
  IV U47143 ( .A(p_input[1813]), .Z(n47009) );
  XOR U47144 ( .A(n47366), .B(n47367), .Z(n47362) );
  AND U47145 ( .A(n47368), .B(n47369), .Z(n47367) );
  XNOR U47146 ( .A(p_input[1844]), .B(n47366), .Z(n47369) );
  XNOR U47147 ( .A(n47366), .B(n47018), .Z(n47368) );
  IV U47148 ( .A(p_input[1812]), .Z(n47018) );
  XOR U47149 ( .A(n47370), .B(n47371), .Z(n47366) );
  AND U47150 ( .A(n47372), .B(n47373), .Z(n47371) );
  XNOR U47151 ( .A(p_input[1843]), .B(n47370), .Z(n47373) );
  XNOR U47152 ( .A(n47370), .B(n47027), .Z(n47372) );
  IV U47153 ( .A(p_input[1811]), .Z(n47027) );
  XOR U47154 ( .A(n47374), .B(n47375), .Z(n47370) );
  AND U47155 ( .A(n47376), .B(n47377), .Z(n47375) );
  XNOR U47156 ( .A(p_input[1842]), .B(n47374), .Z(n47377) );
  XNOR U47157 ( .A(n47374), .B(n47036), .Z(n47376) );
  IV U47158 ( .A(p_input[1810]), .Z(n47036) );
  XOR U47159 ( .A(n47378), .B(n47379), .Z(n47374) );
  AND U47160 ( .A(n47380), .B(n47381), .Z(n47379) );
  XNOR U47161 ( .A(p_input[1841]), .B(n47378), .Z(n47381) );
  XNOR U47162 ( .A(n47378), .B(n47045), .Z(n47380) );
  IV U47163 ( .A(p_input[1809]), .Z(n47045) );
  XOR U47164 ( .A(n47382), .B(n47383), .Z(n47378) );
  AND U47165 ( .A(n47384), .B(n47385), .Z(n47383) );
  XNOR U47166 ( .A(p_input[1840]), .B(n47382), .Z(n47385) );
  XNOR U47167 ( .A(n47382), .B(n47054), .Z(n47384) );
  IV U47168 ( .A(p_input[1808]), .Z(n47054) );
  XOR U47169 ( .A(n47386), .B(n47387), .Z(n47382) );
  AND U47170 ( .A(n47388), .B(n47389), .Z(n47387) );
  XNOR U47171 ( .A(p_input[1839]), .B(n47386), .Z(n47389) );
  XNOR U47172 ( .A(n47386), .B(n47063), .Z(n47388) );
  IV U47173 ( .A(p_input[1807]), .Z(n47063) );
  XOR U47174 ( .A(n47390), .B(n47391), .Z(n47386) );
  AND U47175 ( .A(n47392), .B(n47393), .Z(n47391) );
  XNOR U47176 ( .A(p_input[1838]), .B(n47390), .Z(n47393) );
  XNOR U47177 ( .A(n47390), .B(n47072), .Z(n47392) );
  IV U47178 ( .A(p_input[1806]), .Z(n47072) );
  XOR U47179 ( .A(n47394), .B(n47395), .Z(n47390) );
  AND U47180 ( .A(n47396), .B(n47397), .Z(n47395) );
  XNOR U47181 ( .A(p_input[1837]), .B(n47394), .Z(n47397) );
  XNOR U47182 ( .A(n47394), .B(n47081), .Z(n47396) );
  IV U47183 ( .A(p_input[1805]), .Z(n47081) );
  XOR U47184 ( .A(n47398), .B(n47399), .Z(n47394) );
  AND U47185 ( .A(n47400), .B(n47401), .Z(n47399) );
  XNOR U47186 ( .A(p_input[1836]), .B(n47398), .Z(n47401) );
  XNOR U47187 ( .A(n47398), .B(n47090), .Z(n47400) );
  IV U47188 ( .A(p_input[1804]), .Z(n47090) );
  XOR U47189 ( .A(n47402), .B(n47403), .Z(n47398) );
  AND U47190 ( .A(n47404), .B(n47405), .Z(n47403) );
  XNOR U47191 ( .A(p_input[1835]), .B(n47402), .Z(n47405) );
  XNOR U47192 ( .A(n47402), .B(n47099), .Z(n47404) );
  IV U47193 ( .A(p_input[1803]), .Z(n47099) );
  XOR U47194 ( .A(n47406), .B(n47407), .Z(n47402) );
  AND U47195 ( .A(n47408), .B(n47409), .Z(n47407) );
  XNOR U47196 ( .A(p_input[1834]), .B(n47406), .Z(n47409) );
  XNOR U47197 ( .A(n47406), .B(n47108), .Z(n47408) );
  IV U47198 ( .A(p_input[1802]), .Z(n47108) );
  XOR U47199 ( .A(n47410), .B(n47411), .Z(n47406) );
  AND U47200 ( .A(n47412), .B(n47413), .Z(n47411) );
  XNOR U47201 ( .A(p_input[1833]), .B(n47410), .Z(n47413) );
  XNOR U47202 ( .A(n47410), .B(n47117), .Z(n47412) );
  IV U47203 ( .A(p_input[1801]), .Z(n47117) );
  XOR U47204 ( .A(n47414), .B(n47415), .Z(n47410) );
  AND U47205 ( .A(n47416), .B(n47417), .Z(n47415) );
  XNOR U47206 ( .A(p_input[1832]), .B(n47414), .Z(n47417) );
  XNOR U47207 ( .A(n47414), .B(n47126), .Z(n47416) );
  IV U47208 ( .A(p_input[1800]), .Z(n47126) );
  XOR U47209 ( .A(n47418), .B(n47419), .Z(n47414) );
  AND U47210 ( .A(n47420), .B(n47421), .Z(n47419) );
  XNOR U47211 ( .A(p_input[1831]), .B(n47418), .Z(n47421) );
  XNOR U47212 ( .A(n47418), .B(n47135), .Z(n47420) );
  IV U47213 ( .A(p_input[1799]), .Z(n47135) );
  XOR U47214 ( .A(n47422), .B(n47423), .Z(n47418) );
  AND U47215 ( .A(n47424), .B(n47425), .Z(n47423) );
  XNOR U47216 ( .A(p_input[1830]), .B(n47422), .Z(n47425) );
  XNOR U47217 ( .A(n47422), .B(n47144), .Z(n47424) );
  IV U47218 ( .A(p_input[1798]), .Z(n47144) );
  XOR U47219 ( .A(n47426), .B(n47427), .Z(n47422) );
  AND U47220 ( .A(n47428), .B(n47429), .Z(n47427) );
  XNOR U47221 ( .A(p_input[1829]), .B(n47426), .Z(n47429) );
  XNOR U47222 ( .A(n47426), .B(n47153), .Z(n47428) );
  IV U47223 ( .A(p_input[1797]), .Z(n47153) );
  XOR U47224 ( .A(n47430), .B(n47431), .Z(n47426) );
  AND U47225 ( .A(n47432), .B(n47433), .Z(n47431) );
  XNOR U47226 ( .A(p_input[1828]), .B(n47430), .Z(n47433) );
  XNOR U47227 ( .A(n47430), .B(n47162), .Z(n47432) );
  IV U47228 ( .A(p_input[1796]), .Z(n47162) );
  XOR U47229 ( .A(n47434), .B(n47435), .Z(n47430) );
  AND U47230 ( .A(n47436), .B(n47437), .Z(n47435) );
  XNOR U47231 ( .A(p_input[1827]), .B(n47434), .Z(n47437) );
  XNOR U47232 ( .A(n47434), .B(n47171), .Z(n47436) );
  IV U47233 ( .A(p_input[1795]), .Z(n47171) );
  XOR U47234 ( .A(n47438), .B(n47439), .Z(n47434) );
  AND U47235 ( .A(n47440), .B(n47441), .Z(n47439) );
  XNOR U47236 ( .A(p_input[1826]), .B(n47438), .Z(n47441) );
  XNOR U47237 ( .A(n47438), .B(n47180), .Z(n47440) );
  IV U47238 ( .A(p_input[1794]), .Z(n47180) );
  XNOR U47239 ( .A(n47442), .B(n47443), .Z(n47438) );
  AND U47240 ( .A(n47444), .B(n47445), .Z(n47443) );
  XOR U47241 ( .A(p_input[1825]), .B(n47442), .Z(n47445) );
  XNOR U47242 ( .A(p_input[1793]), .B(n47442), .Z(n47444) );
  AND U47243 ( .A(p_input[1824]), .B(n47446), .Z(n47442) );
  IV U47244 ( .A(p_input[1792]), .Z(n47446) );
  XOR U47245 ( .A(n47447), .B(n47448), .Z(n45625) );
  AND U47246 ( .A(n901), .B(n47449), .Z(n47448) );
  XNOR U47247 ( .A(n47450), .B(n47447), .Z(n47449) );
  XOR U47248 ( .A(n47451), .B(n47452), .Z(n901) );
  AND U47249 ( .A(n47453), .B(n47454), .Z(n47452) );
  XOR U47250 ( .A(n47451), .B(n45640), .Z(n47454) );
  XNOR U47251 ( .A(n47455), .B(n47456), .Z(n45640) );
  AND U47252 ( .A(n47457), .B(n627), .Z(n47456) );
  AND U47253 ( .A(n47455), .B(n47458), .Z(n47457) );
  XNOR U47254 ( .A(n45637), .B(n47451), .Z(n47453) );
  XOR U47255 ( .A(n47459), .B(n47460), .Z(n45637) );
  AND U47256 ( .A(n47461), .B(n624), .Z(n47460) );
  NOR U47257 ( .A(n47459), .B(n47462), .Z(n47461) );
  XOR U47258 ( .A(n47463), .B(n47464), .Z(n47451) );
  AND U47259 ( .A(n47465), .B(n47466), .Z(n47464) );
  XOR U47260 ( .A(n47463), .B(n45652), .Z(n47466) );
  XOR U47261 ( .A(n47467), .B(n47468), .Z(n45652) );
  AND U47262 ( .A(n627), .B(n47469), .Z(n47468) );
  XOR U47263 ( .A(n47470), .B(n47467), .Z(n47469) );
  XNOR U47264 ( .A(n45649), .B(n47463), .Z(n47465) );
  XOR U47265 ( .A(n47471), .B(n47472), .Z(n45649) );
  AND U47266 ( .A(n624), .B(n47473), .Z(n47472) );
  XOR U47267 ( .A(n47474), .B(n47471), .Z(n47473) );
  XOR U47268 ( .A(n47475), .B(n47476), .Z(n47463) );
  AND U47269 ( .A(n47477), .B(n47478), .Z(n47476) );
  XOR U47270 ( .A(n47475), .B(n45664), .Z(n47478) );
  XOR U47271 ( .A(n47479), .B(n47480), .Z(n45664) );
  AND U47272 ( .A(n627), .B(n47481), .Z(n47480) );
  XOR U47273 ( .A(n47482), .B(n47479), .Z(n47481) );
  XNOR U47274 ( .A(n45661), .B(n47475), .Z(n47477) );
  XOR U47275 ( .A(n47483), .B(n47484), .Z(n45661) );
  AND U47276 ( .A(n624), .B(n47485), .Z(n47484) );
  XOR U47277 ( .A(n47486), .B(n47483), .Z(n47485) );
  XOR U47278 ( .A(n47487), .B(n47488), .Z(n47475) );
  AND U47279 ( .A(n47489), .B(n47490), .Z(n47488) );
  XOR U47280 ( .A(n47487), .B(n45676), .Z(n47490) );
  XOR U47281 ( .A(n47491), .B(n47492), .Z(n45676) );
  AND U47282 ( .A(n627), .B(n47493), .Z(n47492) );
  XOR U47283 ( .A(n47494), .B(n47491), .Z(n47493) );
  XNOR U47284 ( .A(n45673), .B(n47487), .Z(n47489) );
  XOR U47285 ( .A(n47495), .B(n47496), .Z(n45673) );
  AND U47286 ( .A(n624), .B(n47497), .Z(n47496) );
  XOR U47287 ( .A(n47498), .B(n47495), .Z(n47497) );
  XOR U47288 ( .A(n47499), .B(n47500), .Z(n47487) );
  AND U47289 ( .A(n47501), .B(n47502), .Z(n47500) );
  XOR U47290 ( .A(n47499), .B(n45688), .Z(n47502) );
  XOR U47291 ( .A(n47503), .B(n47504), .Z(n45688) );
  AND U47292 ( .A(n627), .B(n47505), .Z(n47504) );
  XOR U47293 ( .A(n47506), .B(n47503), .Z(n47505) );
  XNOR U47294 ( .A(n45685), .B(n47499), .Z(n47501) );
  XOR U47295 ( .A(n47507), .B(n47508), .Z(n45685) );
  AND U47296 ( .A(n624), .B(n47509), .Z(n47508) );
  XOR U47297 ( .A(n47510), .B(n47507), .Z(n47509) );
  XOR U47298 ( .A(n47511), .B(n47512), .Z(n47499) );
  AND U47299 ( .A(n47513), .B(n47514), .Z(n47512) );
  XOR U47300 ( .A(n47511), .B(n45700), .Z(n47514) );
  XOR U47301 ( .A(n47515), .B(n47516), .Z(n45700) );
  AND U47302 ( .A(n627), .B(n47517), .Z(n47516) );
  XOR U47303 ( .A(n47518), .B(n47515), .Z(n47517) );
  XNOR U47304 ( .A(n45697), .B(n47511), .Z(n47513) );
  XOR U47305 ( .A(n47519), .B(n47520), .Z(n45697) );
  AND U47306 ( .A(n624), .B(n47521), .Z(n47520) );
  XOR U47307 ( .A(n47522), .B(n47519), .Z(n47521) );
  XOR U47308 ( .A(n47523), .B(n47524), .Z(n47511) );
  AND U47309 ( .A(n47525), .B(n47526), .Z(n47524) );
  XOR U47310 ( .A(n47523), .B(n45712), .Z(n47526) );
  XOR U47311 ( .A(n47527), .B(n47528), .Z(n45712) );
  AND U47312 ( .A(n627), .B(n47529), .Z(n47528) );
  XOR U47313 ( .A(n47530), .B(n47527), .Z(n47529) );
  XNOR U47314 ( .A(n45709), .B(n47523), .Z(n47525) );
  XOR U47315 ( .A(n47531), .B(n47532), .Z(n45709) );
  AND U47316 ( .A(n624), .B(n47533), .Z(n47532) );
  XOR U47317 ( .A(n47534), .B(n47531), .Z(n47533) );
  XOR U47318 ( .A(n47535), .B(n47536), .Z(n47523) );
  AND U47319 ( .A(n47537), .B(n47538), .Z(n47536) );
  XOR U47320 ( .A(n47535), .B(n45724), .Z(n47538) );
  XOR U47321 ( .A(n47539), .B(n47540), .Z(n45724) );
  AND U47322 ( .A(n627), .B(n47541), .Z(n47540) );
  XOR U47323 ( .A(n47542), .B(n47539), .Z(n47541) );
  XNOR U47324 ( .A(n45721), .B(n47535), .Z(n47537) );
  XOR U47325 ( .A(n47543), .B(n47544), .Z(n45721) );
  AND U47326 ( .A(n624), .B(n47545), .Z(n47544) );
  XOR U47327 ( .A(n47546), .B(n47543), .Z(n47545) );
  XOR U47328 ( .A(n47547), .B(n47548), .Z(n47535) );
  AND U47329 ( .A(n47549), .B(n47550), .Z(n47548) );
  XOR U47330 ( .A(n47547), .B(n45736), .Z(n47550) );
  XOR U47331 ( .A(n47551), .B(n47552), .Z(n45736) );
  AND U47332 ( .A(n627), .B(n47553), .Z(n47552) );
  XOR U47333 ( .A(n47554), .B(n47551), .Z(n47553) );
  XNOR U47334 ( .A(n45733), .B(n47547), .Z(n47549) );
  XOR U47335 ( .A(n47555), .B(n47556), .Z(n45733) );
  AND U47336 ( .A(n624), .B(n47557), .Z(n47556) );
  XOR U47337 ( .A(n47558), .B(n47555), .Z(n47557) );
  XOR U47338 ( .A(n47559), .B(n47560), .Z(n47547) );
  AND U47339 ( .A(n47561), .B(n47562), .Z(n47560) );
  XOR U47340 ( .A(n47559), .B(n45748), .Z(n47562) );
  XOR U47341 ( .A(n47563), .B(n47564), .Z(n45748) );
  AND U47342 ( .A(n627), .B(n47565), .Z(n47564) );
  XOR U47343 ( .A(n47566), .B(n47563), .Z(n47565) );
  XNOR U47344 ( .A(n45745), .B(n47559), .Z(n47561) );
  XOR U47345 ( .A(n47567), .B(n47568), .Z(n45745) );
  AND U47346 ( .A(n624), .B(n47569), .Z(n47568) );
  XOR U47347 ( .A(n47570), .B(n47567), .Z(n47569) );
  XOR U47348 ( .A(n47571), .B(n47572), .Z(n47559) );
  AND U47349 ( .A(n47573), .B(n47574), .Z(n47572) );
  XOR U47350 ( .A(n47571), .B(n45760), .Z(n47574) );
  XOR U47351 ( .A(n47575), .B(n47576), .Z(n45760) );
  AND U47352 ( .A(n627), .B(n47577), .Z(n47576) );
  XOR U47353 ( .A(n47578), .B(n47575), .Z(n47577) );
  XNOR U47354 ( .A(n45757), .B(n47571), .Z(n47573) );
  XOR U47355 ( .A(n47579), .B(n47580), .Z(n45757) );
  AND U47356 ( .A(n624), .B(n47581), .Z(n47580) );
  XOR U47357 ( .A(n47582), .B(n47579), .Z(n47581) );
  XOR U47358 ( .A(n47583), .B(n47584), .Z(n47571) );
  AND U47359 ( .A(n47585), .B(n47586), .Z(n47584) );
  XOR U47360 ( .A(n47583), .B(n45772), .Z(n47586) );
  XOR U47361 ( .A(n47587), .B(n47588), .Z(n45772) );
  AND U47362 ( .A(n627), .B(n47589), .Z(n47588) );
  XOR U47363 ( .A(n47590), .B(n47587), .Z(n47589) );
  XNOR U47364 ( .A(n45769), .B(n47583), .Z(n47585) );
  XOR U47365 ( .A(n47591), .B(n47592), .Z(n45769) );
  AND U47366 ( .A(n624), .B(n47593), .Z(n47592) );
  XOR U47367 ( .A(n47594), .B(n47591), .Z(n47593) );
  XOR U47368 ( .A(n47595), .B(n47596), .Z(n47583) );
  AND U47369 ( .A(n47597), .B(n47598), .Z(n47596) );
  XOR U47370 ( .A(n47595), .B(n45784), .Z(n47598) );
  XOR U47371 ( .A(n47599), .B(n47600), .Z(n45784) );
  AND U47372 ( .A(n627), .B(n47601), .Z(n47600) );
  XOR U47373 ( .A(n47602), .B(n47599), .Z(n47601) );
  XNOR U47374 ( .A(n45781), .B(n47595), .Z(n47597) );
  XOR U47375 ( .A(n47603), .B(n47604), .Z(n45781) );
  AND U47376 ( .A(n624), .B(n47605), .Z(n47604) );
  XOR U47377 ( .A(n47606), .B(n47603), .Z(n47605) );
  XOR U47378 ( .A(n47607), .B(n47608), .Z(n47595) );
  AND U47379 ( .A(n47609), .B(n47610), .Z(n47608) );
  XOR U47380 ( .A(n47607), .B(n45796), .Z(n47610) );
  XOR U47381 ( .A(n47611), .B(n47612), .Z(n45796) );
  AND U47382 ( .A(n627), .B(n47613), .Z(n47612) );
  XOR U47383 ( .A(n47614), .B(n47611), .Z(n47613) );
  XNOR U47384 ( .A(n45793), .B(n47607), .Z(n47609) );
  XOR U47385 ( .A(n47615), .B(n47616), .Z(n45793) );
  AND U47386 ( .A(n624), .B(n47617), .Z(n47616) );
  XOR U47387 ( .A(n47618), .B(n47615), .Z(n47617) );
  XOR U47388 ( .A(n47619), .B(n47620), .Z(n47607) );
  AND U47389 ( .A(n47621), .B(n47622), .Z(n47620) );
  XOR U47390 ( .A(n47619), .B(n45808), .Z(n47622) );
  XOR U47391 ( .A(n47623), .B(n47624), .Z(n45808) );
  AND U47392 ( .A(n627), .B(n47625), .Z(n47624) );
  XOR U47393 ( .A(n47626), .B(n47623), .Z(n47625) );
  XNOR U47394 ( .A(n45805), .B(n47619), .Z(n47621) );
  XOR U47395 ( .A(n47627), .B(n47628), .Z(n45805) );
  AND U47396 ( .A(n624), .B(n47629), .Z(n47628) );
  XOR U47397 ( .A(n47630), .B(n47627), .Z(n47629) );
  XOR U47398 ( .A(n47631), .B(n47632), .Z(n47619) );
  AND U47399 ( .A(n47633), .B(n47634), .Z(n47632) );
  XOR U47400 ( .A(n47631), .B(n45820), .Z(n47634) );
  XOR U47401 ( .A(n47635), .B(n47636), .Z(n45820) );
  AND U47402 ( .A(n627), .B(n47637), .Z(n47636) );
  XOR U47403 ( .A(n47638), .B(n47635), .Z(n47637) );
  XNOR U47404 ( .A(n45817), .B(n47631), .Z(n47633) );
  XOR U47405 ( .A(n47639), .B(n47640), .Z(n45817) );
  AND U47406 ( .A(n624), .B(n47641), .Z(n47640) );
  XOR U47407 ( .A(n47642), .B(n47639), .Z(n47641) );
  XOR U47408 ( .A(n47643), .B(n47644), .Z(n47631) );
  AND U47409 ( .A(n47645), .B(n47646), .Z(n47644) );
  XOR U47410 ( .A(n47643), .B(n45832), .Z(n47646) );
  XOR U47411 ( .A(n47647), .B(n47648), .Z(n45832) );
  AND U47412 ( .A(n627), .B(n47649), .Z(n47648) );
  XOR U47413 ( .A(n47650), .B(n47647), .Z(n47649) );
  XNOR U47414 ( .A(n45829), .B(n47643), .Z(n47645) );
  XOR U47415 ( .A(n47651), .B(n47652), .Z(n45829) );
  AND U47416 ( .A(n624), .B(n47653), .Z(n47652) );
  XOR U47417 ( .A(n47654), .B(n47651), .Z(n47653) );
  XOR U47418 ( .A(n47655), .B(n47656), .Z(n47643) );
  AND U47419 ( .A(n47657), .B(n47658), .Z(n47656) );
  XOR U47420 ( .A(n47655), .B(n45844), .Z(n47658) );
  XOR U47421 ( .A(n47659), .B(n47660), .Z(n45844) );
  AND U47422 ( .A(n627), .B(n47661), .Z(n47660) );
  XOR U47423 ( .A(n47662), .B(n47659), .Z(n47661) );
  XNOR U47424 ( .A(n45841), .B(n47655), .Z(n47657) );
  XOR U47425 ( .A(n47663), .B(n47664), .Z(n45841) );
  AND U47426 ( .A(n624), .B(n47665), .Z(n47664) );
  XOR U47427 ( .A(n47666), .B(n47663), .Z(n47665) );
  XOR U47428 ( .A(n47667), .B(n47668), .Z(n47655) );
  AND U47429 ( .A(n47669), .B(n47670), .Z(n47668) );
  XOR U47430 ( .A(n47667), .B(n45856), .Z(n47670) );
  XOR U47431 ( .A(n47671), .B(n47672), .Z(n45856) );
  AND U47432 ( .A(n627), .B(n47673), .Z(n47672) );
  XOR U47433 ( .A(n47674), .B(n47671), .Z(n47673) );
  XNOR U47434 ( .A(n45853), .B(n47667), .Z(n47669) );
  XOR U47435 ( .A(n47675), .B(n47676), .Z(n45853) );
  AND U47436 ( .A(n624), .B(n47677), .Z(n47676) );
  XOR U47437 ( .A(n47678), .B(n47675), .Z(n47677) );
  XOR U47438 ( .A(n47679), .B(n47680), .Z(n47667) );
  AND U47439 ( .A(n47681), .B(n47682), .Z(n47680) );
  XOR U47440 ( .A(n47679), .B(n45868), .Z(n47682) );
  XOR U47441 ( .A(n47683), .B(n47684), .Z(n45868) );
  AND U47442 ( .A(n627), .B(n47685), .Z(n47684) );
  XOR U47443 ( .A(n47686), .B(n47683), .Z(n47685) );
  XNOR U47444 ( .A(n45865), .B(n47679), .Z(n47681) );
  XOR U47445 ( .A(n47687), .B(n47688), .Z(n45865) );
  AND U47446 ( .A(n624), .B(n47689), .Z(n47688) );
  XOR U47447 ( .A(n47690), .B(n47687), .Z(n47689) );
  XOR U47448 ( .A(n47691), .B(n47692), .Z(n47679) );
  AND U47449 ( .A(n47693), .B(n47694), .Z(n47692) );
  XOR U47450 ( .A(n47691), .B(n45880), .Z(n47694) );
  XOR U47451 ( .A(n47695), .B(n47696), .Z(n45880) );
  AND U47452 ( .A(n627), .B(n47697), .Z(n47696) );
  XOR U47453 ( .A(n47698), .B(n47695), .Z(n47697) );
  XNOR U47454 ( .A(n45877), .B(n47691), .Z(n47693) );
  XOR U47455 ( .A(n47699), .B(n47700), .Z(n45877) );
  AND U47456 ( .A(n624), .B(n47701), .Z(n47700) );
  XOR U47457 ( .A(n47702), .B(n47699), .Z(n47701) );
  XOR U47458 ( .A(n47703), .B(n47704), .Z(n47691) );
  AND U47459 ( .A(n47705), .B(n47706), .Z(n47704) );
  XOR U47460 ( .A(n47703), .B(n45892), .Z(n47706) );
  XOR U47461 ( .A(n47707), .B(n47708), .Z(n45892) );
  AND U47462 ( .A(n627), .B(n47709), .Z(n47708) );
  XOR U47463 ( .A(n47710), .B(n47707), .Z(n47709) );
  XNOR U47464 ( .A(n45889), .B(n47703), .Z(n47705) );
  XOR U47465 ( .A(n47711), .B(n47712), .Z(n45889) );
  AND U47466 ( .A(n624), .B(n47713), .Z(n47712) );
  XOR U47467 ( .A(n47714), .B(n47711), .Z(n47713) );
  XOR U47468 ( .A(n47715), .B(n47716), .Z(n47703) );
  AND U47469 ( .A(n47717), .B(n47718), .Z(n47716) );
  XOR U47470 ( .A(n47715), .B(n45904), .Z(n47718) );
  XOR U47471 ( .A(n47719), .B(n47720), .Z(n45904) );
  AND U47472 ( .A(n627), .B(n47721), .Z(n47720) );
  XOR U47473 ( .A(n47722), .B(n47719), .Z(n47721) );
  XNOR U47474 ( .A(n45901), .B(n47715), .Z(n47717) );
  XOR U47475 ( .A(n47723), .B(n47724), .Z(n45901) );
  AND U47476 ( .A(n624), .B(n47725), .Z(n47724) );
  XOR U47477 ( .A(n47726), .B(n47723), .Z(n47725) );
  XOR U47478 ( .A(n47727), .B(n47728), .Z(n47715) );
  AND U47479 ( .A(n47729), .B(n47730), .Z(n47728) );
  XOR U47480 ( .A(n47727), .B(n45916), .Z(n47730) );
  XOR U47481 ( .A(n47731), .B(n47732), .Z(n45916) );
  AND U47482 ( .A(n627), .B(n47733), .Z(n47732) );
  XOR U47483 ( .A(n47734), .B(n47731), .Z(n47733) );
  XNOR U47484 ( .A(n45913), .B(n47727), .Z(n47729) );
  XOR U47485 ( .A(n47735), .B(n47736), .Z(n45913) );
  AND U47486 ( .A(n624), .B(n47737), .Z(n47736) );
  XOR U47487 ( .A(n47738), .B(n47735), .Z(n47737) );
  XOR U47488 ( .A(n47739), .B(n47740), .Z(n47727) );
  AND U47489 ( .A(n47741), .B(n47742), .Z(n47740) );
  XOR U47490 ( .A(n47739), .B(n45928), .Z(n47742) );
  XOR U47491 ( .A(n47743), .B(n47744), .Z(n45928) );
  AND U47492 ( .A(n627), .B(n47745), .Z(n47744) );
  XOR U47493 ( .A(n47746), .B(n47743), .Z(n47745) );
  XNOR U47494 ( .A(n45925), .B(n47739), .Z(n47741) );
  XOR U47495 ( .A(n47747), .B(n47748), .Z(n45925) );
  AND U47496 ( .A(n624), .B(n47749), .Z(n47748) );
  XOR U47497 ( .A(n47750), .B(n47747), .Z(n47749) );
  XOR U47498 ( .A(n47751), .B(n47752), .Z(n47739) );
  AND U47499 ( .A(n47753), .B(n47754), .Z(n47752) );
  XOR U47500 ( .A(n47751), .B(n45940), .Z(n47754) );
  XOR U47501 ( .A(n47755), .B(n47756), .Z(n45940) );
  AND U47502 ( .A(n627), .B(n47757), .Z(n47756) );
  XOR U47503 ( .A(n47758), .B(n47755), .Z(n47757) );
  XNOR U47504 ( .A(n45937), .B(n47751), .Z(n47753) );
  XOR U47505 ( .A(n47759), .B(n47760), .Z(n45937) );
  AND U47506 ( .A(n624), .B(n47761), .Z(n47760) );
  XOR U47507 ( .A(n47762), .B(n47759), .Z(n47761) );
  XOR U47508 ( .A(n47763), .B(n47764), .Z(n47751) );
  AND U47509 ( .A(n47765), .B(n47766), .Z(n47764) );
  XOR U47510 ( .A(n47763), .B(n45952), .Z(n47766) );
  XOR U47511 ( .A(n47767), .B(n47768), .Z(n45952) );
  AND U47512 ( .A(n627), .B(n47769), .Z(n47768) );
  XOR U47513 ( .A(n47770), .B(n47767), .Z(n47769) );
  XNOR U47514 ( .A(n45949), .B(n47763), .Z(n47765) );
  XOR U47515 ( .A(n47771), .B(n47772), .Z(n45949) );
  AND U47516 ( .A(n624), .B(n47773), .Z(n47772) );
  XOR U47517 ( .A(n47774), .B(n47771), .Z(n47773) );
  XOR U47518 ( .A(n47775), .B(n47776), .Z(n47763) );
  AND U47519 ( .A(n47777), .B(n47778), .Z(n47776) );
  XOR U47520 ( .A(n47775), .B(n45964), .Z(n47778) );
  XOR U47521 ( .A(n47779), .B(n47780), .Z(n45964) );
  AND U47522 ( .A(n627), .B(n47781), .Z(n47780) );
  XOR U47523 ( .A(n47782), .B(n47779), .Z(n47781) );
  XNOR U47524 ( .A(n45961), .B(n47775), .Z(n47777) );
  XOR U47525 ( .A(n47783), .B(n47784), .Z(n45961) );
  AND U47526 ( .A(n624), .B(n47785), .Z(n47784) );
  XOR U47527 ( .A(n47786), .B(n47783), .Z(n47785) );
  XOR U47528 ( .A(n47787), .B(n47788), .Z(n47775) );
  AND U47529 ( .A(n47789), .B(n47790), .Z(n47788) );
  XOR U47530 ( .A(n47787), .B(n45976), .Z(n47790) );
  XOR U47531 ( .A(n47791), .B(n47792), .Z(n45976) );
  AND U47532 ( .A(n627), .B(n47793), .Z(n47792) );
  XOR U47533 ( .A(n47794), .B(n47791), .Z(n47793) );
  XNOR U47534 ( .A(n45973), .B(n47787), .Z(n47789) );
  XOR U47535 ( .A(n47795), .B(n47796), .Z(n45973) );
  AND U47536 ( .A(n624), .B(n47797), .Z(n47796) );
  XOR U47537 ( .A(n47798), .B(n47795), .Z(n47797) );
  XOR U47538 ( .A(n47799), .B(n47800), .Z(n47787) );
  AND U47539 ( .A(n47801), .B(n47802), .Z(n47800) );
  XOR U47540 ( .A(n47799), .B(n45988), .Z(n47802) );
  XOR U47541 ( .A(n47803), .B(n47804), .Z(n45988) );
  AND U47542 ( .A(n627), .B(n47805), .Z(n47804) );
  XOR U47543 ( .A(n47806), .B(n47803), .Z(n47805) );
  XNOR U47544 ( .A(n45985), .B(n47799), .Z(n47801) );
  XOR U47545 ( .A(n47807), .B(n47808), .Z(n45985) );
  AND U47546 ( .A(n624), .B(n47809), .Z(n47808) );
  XOR U47547 ( .A(n47810), .B(n47807), .Z(n47809) );
  XOR U47548 ( .A(n47811), .B(n47812), .Z(n47799) );
  AND U47549 ( .A(n47813), .B(n47814), .Z(n47812) );
  XNOR U47550 ( .A(n47815), .B(n46001), .Z(n47814) );
  XOR U47551 ( .A(n47816), .B(n47817), .Z(n46001) );
  AND U47552 ( .A(n627), .B(n47818), .Z(n47817) );
  XOR U47553 ( .A(n47816), .B(n47819), .Z(n47818) );
  XNOR U47554 ( .A(n45998), .B(n47811), .Z(n47813) );
  XOR U47555 ( .A(n47820), .B(n47821), .Z(n45998) );
  AND U47556 ( .A(n624), .B(n47822), .Z(n47821) );
  XOR U47557 ( .A(n47820), .B(n47823), .Z(n47822) );
  IV U47558 ( .A(n47815), .Z(n47811) );
  AND U47559 ( .A(n47447), .B(n47450), .Z(n47815) );
  XNOR U47560 ( .A(n47824), .B(n47825), .Z(n47450) );
  AND U47561 ( .A(n627), .B(n47826), .Z(n47825) );
  XNOR U47562 ( .A(n47827), .B(n47824), .Z(n47826) );
  XOR U47563 ( .A(n47828), .B(n47829), .Z(n627) );
  AND U47564 ( .A(n47830), .B(n47831), .Z(n47829) );
  XOR U47565 ( .A(n47458), .B(n47828), .Z(n47831) );
  IV U47566 ( .A(n47832), .Z(n47458) );
  AND U47567 ( .A(p_input[1791]), .B(p_input[1759]), .Z(n47832) );
  XOR U47568 ( .A(n47828), .B(n47455), .Z(n47830) );
  AND U47569 ( .A(p_input[1695]), .B(p_input[1727]), .Z(n47455) );
  XOR U47570 ( .A(n47833), .B(n47834), .Z(n47828) );
  AND U47571 ( .A(n47835), .B(n47836), .Z(n47834) );
  XOR U47572 ( .A(n47833), .B(n47470), .Z(n47836) );
  XNOR U47573 ( .A(p_input[1758]), .B(n47837), .Z(n47470) );
  AND U47574 ( .A(n951), .B(n47838), .Z(n47837) );
  XOR U47575 ( .A(p_input[1790]), .B(p_input[1758]), .Z(n47838) );
  XNOR U47576 ( .A(n47467), .B(n47833), .Z(n47835) );
  XOR U47577 ( .A(n47839), .B(n47840), .Z(n47467) );
  AND U47578 ( .A(n949), .B(n47841), .Z(n47840) );
  XOR U47579 ( .A(p_input[1726]), .B(p_input[1694]), .Z(n47841) );
  XOR U47580 ( .A(n47842), .B(n47843), .Z(n47833) );
  AND U47581 ( .A(n47844), .B(n47845), .Z(n47843) );
  XOR U47582 ( .A(n47842), .B(n47482), .Z(n47845) );
  XNOR U47583 ( .A(p_input[1757]), .B(n47846), .Z(n47482) );
  AND U47584 ( .A(n951), .B(n47847), .Z(n47846) );
  XOR U47585 ( .A(p_input[1789]), .B(p_input[1757]), .Z(n47847) );
  XNOR U47586 ( .A(n47479), .B(n47842), .Z(n47844) );
  XOR U47587 ( .A(n47848), .B(n47849), .Z(n47479) );
  AND U47588 ( .A(n949), .B(n47850), .Z(n47849) );
  XOR U47589 ( .A(p_input[1725]), .B(p_input[1693]), .Z(n47850) );
  XOR U47590 ( .A(n47851), .B(n47852), .Z(n47842) );
  AND U47591 ( .A(n47853), .B(n47854), .Z(n47852) );
  XOR U47592 ( .A(n47851), .B(n47494), .Z(n47854) );
  XNOR U47593 ( .A(p_input[1756]), .B(n47855), .Z(n47494) );
  AND U47594 ( .A(n951), .B(n47856), .Z(n47855) );
  XOR U47595 ( .A(p_input[1788]), .B(p_input[1756]), .Z(n47856) );
  XNOR U47596 ( .A(n47491), .B(n47851), .Z(n47853) );
  XOR U47597 ( .A(n47857), .B(n47858), .Z(n47491) );
  AND U47598 ( .A(n949), .B(n47859), .Z(n47858) );
  XOR U47599 ( .A(p_input[1724]), .B(p_input[1692]), .Z(n47859) );
  XOR U47600 ( .A(n47860), .B(n47861), .Z(n47851) );
  AND U47601 ( .A(n47862), .B(n47863), .Z(n47861) );
  XOR U47602 ( .A(n47860), .B(n47506), .Z(n47863) );
  XNOR U47603 ( .A(p_input[1755]), .B(n47864), .Z(n47506) );
  AND U47604 ( .A(n951), .B(n47865), .Z(n47864) );
  XOR U47605 ( .A(p_input[1787]), .B(p_input[1755]), .Z(n47865) );
  XNOR U47606 ( .A(n47503), .B(n47860), .Z(n47862) );
  XOR U47607 ( .A(n47866), .B(n47867), .Z(n47503) );
  AND U47608 ( .A(n949), .B(n47868), .Z(n47867) );
  XOR U47609 ( .A(p_input[1723]), .B(p_input[1691]), .Z(n47868) );
  XOR U47610 ( .A(n47869), .B(n47870), .Z(n47860) );
  AND U47611 ( .A(n47871), .B(n47872), .Z(n47870) );
  XOR U47612 ( .A(n47869), .B(n47518), .Z(n47872) );
  XNOR U47613 ( .A(p_input[1754]), .B(n47873), .Z(n47518) );
  AND U47614 ( .A(n951), .B(n47874), .Z(n47873) );
  XOR U47615 ( .A(p_input[1786]), .B(p_input[1754]), .Z(n47874) );
  XNOR U47616 ( .A(n47515), .B(n47869), .Z(n47871) );
  XOR U47617 ( .A(n47875), .B(n47876), .Z(n47515) );
  AND U47618 ( .A(n949), .B(n47877), .Z(n47876) );
  XOR U47619 ( .A(p_input[1722]), .B(p_input[1690]), .Z(n47877) );
  XOR U47620 ( .A(n47878), .B(n47879), .Z(n47869) );
  AND U47621 ( .A(n47880), .B(n47881), .Z(n47879) );
  XOR U47622 ( .A(n47878), .B(n47530), .Z(n47881) );
  XNOR U47623 ( .A(p_input[1753]), .B(n47882), .Z(n47530) );
  AND U47624 ( .A(n951), .B(n47883), .Z(n47882) );
  XOR U47625 ( .A(p_input[1785]), .B(p_input[1753]), .Z(n47883) );
  XNOR U47626 ( .A(n47527), .B(n47878), .Z(n47880) );
  XOR U47627 ( .A(n47884), .B(n47885), .Z(n47527) );
  AND U47628 ( .A(n949), .B(n47886), .Z(n47885) );
  XOR U47629 ( .A(p_input[1721]), .B(p_input[1689]), .Z(n47886) );
  XOR U47630 ( .A(n47887), .B(n47888), .Z(n47878) );
  AND U47631 ( .A(n47889), .B(n47890), .Z(n47888) );
  XOR U47632 ( .A(n47887), .B(n47542), .Z(n47890) );
  XNOR U47633 ( .A(p_input[1752]), .B(n47891), .Z(n47542) );
  AND U47634 ( .A(n951), .B(n47892), .Z(n47891) );
  XOR U47635 ( .A(p_input[1784]), .B(p_input[1752]), .Z(n47892) );
  XNOR U47636 ( .A(n47539), .B(n47887), .Z(n47889) );
  XOR U47637 ( .A(n47893), .B(n47894), .Z(n47539) );
  AND U47638 ( .A(n949), .B(n47895), .Z(n47894) );
  XOR U47639 ( .A(p_input[1720]), .B(p_input[1688]), .Z(n47895) );
  XOR U47640 ( .A(n47896), .B(n47897), .Z(n47887) );
  AND U47641 ( .A(n47898), .B(n47899), .Z(n47897) );
  XOR U47642 ( .A(n47896), .B(n47554), .Z(n47899) );
  XNOR U47643 ( .A(p_input[1751]), .B(n47900), .Z(n47554) );
  AND U47644 ( .A(n951), .B(n47901), .Z(n47900) );
  XOR U47645 ( .A(p_input[1783]), .B(p_input[1751]), .Z(n47901) );
  XNOR U47646 ( .A(n47551), .B(n47896), .Z(n47898) );
  XOR U47647 ( .A(n47902), .B(n47903), .Z(n47551) );
  AND U47648 ( .A(n949), .B(n47904), .Z(n47903) );
  XOR U47649 ( .A(p_input[1719]), .B(p_input[1687]), .Z(n47904) );
  XOR U47650 ( .A(n47905), .B(n47906), .Z(n47896) );
  AND U47651 ( .A(n47907), .B(n47908), .Z(n47906) );
  XOR U47652 ( .A(n47905), .B(n47566), .Z(n47908) );
  XNOR U47653 ( .A(p_input[1750]), .B(n47909), .Z(n47566) );
  AND U47654 ( .A(n951), .B(n47910), .Z(n47909) );
  XOR U47655 ( .A(p_input[1782]), .B(p_input[1750]), .Z(n47910) );
  XNOR U47656 ( .A(n47563), .B(n47905), .Z(n47907) );
  XOR U47657 ( .A(n47911), .B(n47912), .Z(n47563) );
  AND U47658 ( .A(n949), .B(n47913), .Z(n47912) );
  XOR U47659 ( .A(p_input[1718]), .B(p_input[1686]), .Z(n47913) );
  XOR U47660 ( .A(n47914), .B(n47915), .Z(n47905) );
  AND U47661 ( .A(n47916), .B(n47917), .Z(n47915) );
  XOR U47662 ( .A(n47914), .B(n47578), .Z(n47917) );
  XNOR U47663 ( .A(p_input[1749]), .B(n47918), .Z(n47578) );
  AND U47664 ( .A(n951), .B(n47919), .Z(n47918) );
  XOR U47665 ( .A(p_input[1781]), .B(p_input[1749]), .Z(n47919) );
  XNOR U47666 ( .A(n47575), .B(n47914), .Z(n47916) );
  XOR U47667 ( .A(n47920), .B(n47921), .Z(n47575) );
  AND U47668 ( .A(n949), .B(n47922), .Z(n47921) );
  XOR U47669 ( .A(p_input[1717]), .B(p_input[1685]), .Z(n47922) );
  XOR U47670 ( .A(n47923), .B(n47924), .Z(n47914) );
  AND U47671 ( .A(n47925), .B(n47926), .Z(n47924) );
  XOR U47672 ( .A(n47923), .B(n47590), .Z(n47926) );
  XNOR U47673 ( .A(p_input[1748]), .B(n47927), .Z(n47590) );
  AND U47674 ( .A(n951), .B(n47928), .Z(n47927) );
  XOR U47675 ( .A(p_input[1780]), .B(p_input[1748]), .Z(n47928) );
  XNOR U47676 ( .A(n47587), .B(n47923), .Z(n47925) );
  XOR U47677 ( .A(n47929), .B(n47930), .Z(n47587) );
  AND U47678 ( .A(n949), .B(n47931), .Z(n47930) );
  XOR U47679 ( .A(p_input[1716]), .B(p_input[1684]), .Z(n47931) );
  XOR U47680 ( .A(n47932), .B(n47933), .Z(n47923) );
  AND U47681 ( .A(n47934), .B(n47935), .Z(n47933) );
  XOR U47682 ( .A(n47932), .B(n47602), .Z(n47935) );
  XNOR U47683 ( .A(p_input[1747]), .B(n47936), .Z(n47602) );
  AND U47684 ( .A(n951), .B(n47937), .Z(n47936) );
  XOR U47685 ( .A(p_input[1779]), .B(p_input[1747]), .Z(n47937) );
  XNOR U47686 ( .A(n47599), .B(n47932), .Z(n47934) );
  XOR U47687 ( .A(n47938), .B(n47939), .Z(n47599) );
  AND U47688 ( .A(n949), .B(n47940), .Z(n47939) );
  XOR U47689 ( .A(p_input[1715]), .B(p_input[1683]), .Z(n47940) );
  XOR U47690 ( .A(n47941), .B(n47942), .Z(n47932) );
  AND U47691 ( .A(n47943), .B(n47944), .Z(n47942) );
  XOR U47692 ( .A(n47941), .B(n47614), .Z(n47944) );
  XNOR U47693 ( .A(p_input[1746]), .B(n47945), .Z(n47614) );
  AND U47694 ( .A(n951), .B(n47946), .Z(n47945) );
  XOR U47695 ( .A(p_input[1778]), .B(p_input[1746]), .Z(n47946) );
  XNOR U47696 ( .A(n47611), .B(n47941), .Z(n47943) );
  XOR U47697 ( .A(n47947), .B(n47948), .Z(n47611) );
  AND U47698 ( .A(n949), .B(n47949), .Z(n47948) );
  XOR U47699 ( .A(p_input[1714]), .B(p_input[1682]), .Z(n47949) );
  XOR U47700 ( .A(n47950), .B(n47951), .Z(n47941) );
  AND U47701 ( .A(n47952), .B(n47953), .Z(n47951) );
  XOR U47702 ( .A(n47950), .B(n47626), .Z(n47953) );
  XNOR U47703 ( .A(p_input[1745]), .B(n47954), .Z(n47626) );
  AND U47704 ( .A(n951), .B(n47955), .Z(n47954) );
  XOR U47705 ( .A(p_input[1777]), .B(p_input[1745]), .Z(n47955) );
  XNOR U47706 ( .A(n47623), .B(n47950), .Z(n47952) );
  XOR U47707 ( .A(n47956), .B(n47957), .Z(n47623) );
  AND U47708 ( .A(n949), .B(n47958), .Z(n47957) );
  XOR U47709 ( .A(p_input[1713]), .B(p_input[1681]), .Z(n47958) );
  XOR U47710 ( .A(n47959), .B(n47960), .Z(n47950) );
  AND U47711 ( .A(n47961), .B(n47962), .Z(n47960) );
  XOR U47712 ( .A(n47959), .B(n47638), .Z(n47962) );
  XNOR U47713 ( .A(p_input[1744]), .B(n47963), .Z(n47638) );
  AND U47714 ( .A(n951), .B(n47964), .Z(n47963) );
  XOR U47715 ( .A(p_input[1776]), .B(p_input[1744]), .Z(n47964) );
  XNOR U47716 ( .A(n47635), .B(n47959), .Z(n47961) );
  XOR U47717 ( .A(n47965), .B(n47966), .Z(n47635) );
  AND U47718 ( .A(n949), .B(n47967), .Z(n47966) );
  XOR U47719 ( .A(p_input[1712]), .B(p_input[1680]), .Z(n47967) );
  XOR U47720 ( .A(n47968), .B(n47969), .Z(n47959) );
  AND U47721 ( .A(n47970), .B(n47971), .Z(n47969) );
  XOR U47722 ( .A(n47968), .B(n47650), .Z(n47971) );
  XNOR U47723 ( .A(p_input[1743]), .B(n47972), .Z(n47650) );
  AND U47724 ( .A(n951), .B(n47973), .Z(n47972) );
  XOR U47725 ( .A(p_input[1775]), .B(p_input[1743]), .Z(n47973) );
  XNOR U47726 ( .A(n47647), .B(n47968), .Z(n47970) );
  XOR U47727 ( .A(n47974), .B(n47975), .Z(n47647) );
  AND U47728 ( .A(n949), .B(n47976), .Z(n47975) );
  XOR U47729 ( .A(p_input[1711]), .B(p_input[1679]), .Z(n47976) );
  XOR U47730 ( .A(n47977), .B(n47978), .Z(n47968) );
  AND U47731 ( .A(n47979), .B(n47980), .Z(n47978) );
  XOR U47732 ( .A(n47977), .B(n47662), .Z(n47980) );
  XNOR U47733 ( .A(p_input[1742]), .B(n47981), .Z(n47662) );
  AND U47734 ( .A(n951), .B(n47982), .Z(n47981) );
  XOR U47735 ( .A(p_input[1774]), .B(p_input[1742]), .Z(n47982) );
  XNOR U47736 ( .A(n47659), .B(n47977), .Z(n47979) );
  XOR U47737 ( .A(n47983), .B(n47984), .Z(n47659) );
  AND U47738 ( .A(n949), .B(n47985), .Z(n47984) );
  XOR U47739 ( .A(p_input[1710]), .B(p_input[1678]), .Z(n47985) );
  XOR U47740 ( .A(n47986), .B(n47987), .Z(n47977) );
  AND U47741 ( .A(n47988), .B(n47989), .Z(n47987) );
  XOR U47742 ( .A(n47986), .B(n47674), .Z(n47989) );
  XNOR U47743 ( .A(p_input[1741]), .B(n47990), .Z(n47674) );
  AND U47744 ( .A(n951), .B(n47991), .Z(n47990) );
  XOR U47745 ( .A(p_input[1773]), .B(p_input[1741]), .Z(n47991) );
  XNOR U47746 ( .A(n47671), .B(n47986), .Z(n47988) );
  XOR U47747 ( .A(n47992), .B(n47993), .Z(n47671) );
  AND U47748 ( .A(n949), .B(n47994), .Z(n47993) );
  XOR U47749 ( .A(p_input[1709]), .B(p_input[1677]), .Z(n47994) );
  XOR U47750 ( .A(n47995), .B(n47996), .Z(n47986) );
  AND U47751 ( .A(n47997), .B(n47998), .Z(n47996) );
  XOR U47752 ( .A(n47995), .B(n47686), .Z(n47998) );
  XNOR U47753 ( .A(p_input[1740]), .B(n47999), .Z(n47686) );
  AND U47754 ( .A(n951), .B(n48000), .Z(n47999) );
  XOR U47755 ( .A(p_input[1772]), .B(p_input[1740]), .Z(n48000) );
  XNOR U47756 ( .A(n47683), .B(n47995), .Z(n47997) );
  XOR U47757 ( .A(n48001), .B(n48002), .Z(n47683) );
  AND U47758 ( .A(n949), .B(n48003), .Z(n48002) );
  XOR U47759 ( .A(p_input[1708]), .B(p_input[1676]), .Z(n48003) );
  XOR U47760 ( .A(n48004), .B(n48005), .Z(n47995) );
  AND U47761 ( .A(n48006), .B(n48007), .Z(n48005) );
  XOR U47762 ( .A(n48004), .B(n47698), .Z(n48007) );
  XNOR U47763 ( .A(p_input[1739]), .B(n48008), .Z(n47698) );
  AND U47764 ( .A(n951), .B(n48009), .Z(n48008) );
  XOR U47765 ( .A(p_input[1771]), .B(p_input[1739]), .Z(n48009) );
  XNOR U47766 ( .A(n47695), .B(n48004), .Z(n48006) );
  XOR U47767 ( .A(n48010), .B(n48011), .Z(n47695) );
  AND U47768 ( .A(n949), .B(n48012), .Z(n48011) );
  XOR U47769 ( .A(p_input[1707]), .B(p_input[1675]), .Z(n48012) );
  XOR U47770 ( .A(n48013), .B(n48014), .Z(n48004) );
  AND U47771 ( .A(n48015), .B(n48016), .Z(n48014) );
  XOR U47772 ( .A(n48013), .B(n47710), .Z(n48016) );
  XNOR U47773 ( .A(p_input[1738]), .B(n48017), .Z(n47710) );
  AND U47774 ( .A(n951), .B(n48018), .Z(n48017) );
  XOR U47775 ( .A(p_input[1770]), .B(p_input[1738]), .Z(n48018) );
  XNOR U47776 ( .A(n47707), .B(n48013), .Z(n48015) );
  XOR U47777 ( .A(n48019), .B(n48020), .Z(n47707) );
  AND U47778 ( .A(n949), .B(n48021), .Z(n48020) );
  XOR U47779 ( .A(p_input[1706]), .B(p_input[1674]), .Z(n48021) );
  XOR U47780 ( .A(n48022), .B(n48023), .Z(n48013) );
  AND U47781 ( .A(n48024), .B(n48025), .Z(n48023) );
  XOR U47782 ( .A(n48022), .B(n47722), .Z(n48025) );
  XNOR U47783 ( .A(p_input[1737]), .B(n48026), .Z(n47722) );
  AND U47784 ( .A(n951), .B(n48027), .Z(n48026) );
  XOR U47785 ( .A(p_input[1769]), .B(p_input[1737]), .Z(n48027) );
  XNOR U47786 ( .A(n47719), .B(n48022), .Z(n48024) );
  XOR U47787 ( .A(n48028), .B(n48029), .Z(n47719) );
  AND U47788 ( .A(n949), .B(n48030), .Z(n48029) );
  XOR U47789 ( .A(p_input[1705]), .B(p_input[1673]), .Z(n48030) );
  XOR U47790 ( .A(n48031), .B(n48032), .Z(n48022) );
  AND U47791 ( .A(n48033), .B(n48034), .Z(n48032) );
  XOR U47792 ( .A(n48031), .B(n47734), .Z(n48034) );
  XNOR U47793 ( .A(p_input[1736]), .B(n48035), .Z(n47734) );
  AND U47794 ( .A(n951), .B(n48036), .Z(n48035) );
  XOR U47795 ( .A(p_input[1768]), .B(p_input[1736]), .Z(n48036) );
  XNOR U47796 ( .A(n47731), .B(n48031), .Z(n48033) );
  XOR U47797 ( .A(n48037), .B(n48038), .Z(n47731) );
  AND U47798 ( .A(n949), .B(n48039), .Z(n48038) );
  XOR U47799 ( .A(p_input[1704]), .B(p_input[1672]), .Z(n48039) );
  XOR U47800 ( .A(n48040), .B(n48041), .Z(n48031) );
  AND U47801 ( .A(n48042), .B(n48043), .Z(n48041) );
  XOR U47802 ( .A(n48040), .B(n47746), .Z(n48043) );
  XNOR U47803 ( .A(p_input[1735]), .B(n48044), .Z(n47746) );
  AND U47804 ( .A(n951), .B(n48045), .Z(n48044) );
  XOR U47805 ( .A(p_input[1767]), .B(p_input[1735]), .Z(n48045) );
  XNOR U47806 ( .A(n47743), .B(n48040), .Z(n48042) );
  XOR U47807 ( .A(n48046), .B(n48047), .Z(n47743) );
  AND U47808 ( .A(n949), .B(n48048), .Z(n48047) );
  XOR U47809 ( .A(p_input[1703]), .B(p_input[1671]), .Z(n48048) );
  XOR U47810 ( .A(n48049), .B(n48050), .Z(n48040) );
  AND U47811 ( .A(n48051), .B(n48052), .Z(n48050) );
  XOR U47812 ( .A(n48049), .B(n47758), .Z(n48052) );
  XNOR U47813 ( .A(p_input[1734]), .B(n48053), .Z(n47758) );
  AND U47814 ( .A(n951), .B(n48054), .Z(n48053) );
  XOR U47815 ( .A(p_input[1766]), .B(p_input[1734]), .Z(n48054) );
  XNOR U47816 ( .A(n47755), .B(n48049), .Z(n48051) );
  XOR U47817 ( .A(n48055), .B(n48056), .Z(n47755) );
  AND U47818 ( .A(n949), .B(n48057), .Z(n48056) );
  XOR U47819 ( .A(p_input[1702]), .B(p_input[1670]), .Z(n48057) );
  XOR U47820 ( .A(n48058), .B(n48059), .Z(n48049) );
  AND U47821 ( .A(n48060), .B(n48061), .Z(n48059) );
  XOR U47822 ( .A(n48058), .B(n47770), .Z(n48061) );
  XNOR U47823 ( .A(p_input[1733]), .B(n48062), .Z(n47770) );
  AND U47824 ( .A(n951), .B(n48063), .Z(n48062) );
  XOR U47825 ( .A(p_input[1765]), .B(p_input[1733]), .Z(n48063) );
  XNOR U47826 ( .A(n47767), .B(n48058), .Z(n48060) );
  XOR U47827 ( .A(n48064), .B(n48065), .Z(n47767) );
  AND U47828 ( .A(n949), .B(n48066), .Z(n48065) );
  XOR U47829 ( .A(p_input[1701]), .B(p_input[1669]), .Z(n48066) );
  XOR U47830 ( .A(n48067), .B(n48068), .Z(n48058) );
  AND U47831 ( .A(n48069), .B(n48070), .Z(n48068) );
  XOR U47832 ( .A(n48067), .B(n47782), .Z(n48070) );
  XNOR U47833 ( .A(p_input[1732]), .B(n48071), .Z(n47782) );
  AND U47834 ( .A(n951), .B(n48072), .Z(n48071) );
  XOR U47835 ( .A(p_input[1764]), .B(p_input[1732]), .Z(n48072) );
  XNOR U47836 ( .A(n47779), .B(n48067), .Z(n48069) );
  XOR U47837 ( .A(n48073), .B(n48074), .Z(n47779) );
  AND U47838 ( .A(n949), .B(n48075), .Z(n48074) );
  XOR U47839 ( .A(p_input[1700]), .B(p_input[1668]), .Z(n48075) );
  XOR U47840 ( .A(n48076), .B(n48077), .Z(n48067) );
  AND U47841 ( .A(n48078), .B(n48079), .Z(n48077) );
  XOR U47842 ( .A(n48076), .B(n47794), .Z(n48079) );
  XNOR U47843 ( .A(p_input[1731]), .B(n48080), .Z(n47794) );
  AND U47844 ( .A(n951), .B(n48081), .Z(n48080) );
  XOR U47845 ( .A(p_input[1763]), .B(p_input[1731]), .Z(n48081) );
  XNOR U47846 ( .A(n47791), .B(n48076), .Z(n48078) );
  XOR U47847 ( .A(n48082), .B(n48083), .Z(n47791) );
  AND U47848 ( .A(n949), .B(n48084), .Z(n48083) );
  XOR U47849 ( .A(p_input[1699]), .B(p_input[1667]), .Z(n48084) );
  XOR U47850 ( .A(n48085), .B(n48086), .Z(n48076) );
  AND U47851 ( .A(n48087), .B(n48088), .Z(n48086) );
  XOR U47852 ( .A(n48085), .B(n47806), .Z(n48088) );
  XNOR U47853 ( .A(p_input[1730]), .B(n48089), .Z(n47806) );
  AND U47854 ( .A(n951), .B(n48090), .Z(n48089) );
  XOR U47855 ( .A(p_input[1762]), .B(p_input[1730]), .Z(n48090) );
  XNOR U47856 ( .A(n47803), .B(n48085), .Z(n48087) );
  XOR U47857 ( .A(n48091), .B(n48092), .Z(n47803) );
  AND U47858 ( .A(n949), .B(n48093), .Z(n48092) );
  XOR U47859 ( .A(p_input[1698]), .B(p_input[1666]), .Z(n48093) );
  XOR U47860 ( .A(n48094), .B(n48095), .Z(n48085) );
  AND U47861 ( .A(n48096), .B(n48097), .Z(n48095) );
  XNOR U47862 ( .A(n48098), .B(n47819), .Z(n48097) );
  XNOR U47863 ( .A(p_input[1729]), .B(n48099), .Z(n47819) );
  AND U47864 ( .A(n951), .B(n48100), .Z(n48099) );
  XNOR U47865 ( .A(p_input[1761]), .B(n48101), .Z(n48100) );
  IV U47866 ( .A(p_input[1729]), .Z(n48101) );
  XNOR U47867 ( .A(n47816), .B(n48094), .Z(n48096) );
  XNOR U47868 ( .A(p_input[1665]), .B(n48102), .Z(n47816) );
  AND U47869 ( .A(n949), .B(n48103), .Z(n48102) );
  XOR U47870 ( .A(p_input[1697]), .B(p_input[1665]), .Z(n48103) );
  IV U47871 ( .A(n48098), .Z(n48094) );
  AND U47872 ( .A(n47824), .B(n47827), .Z(n48098) );
  XOR U47873 ( .A(p_input[1728]), .B(n48104), .Z(n47827) );
  AND U47874 ( .A(n951), .B(n48105), .Z(n48104) );
  XOR U47875 ( .A(p_input[1760]), .B(p_input[1728]), .Z(n48105) );
  XOR U47876 ( .A(n48106), .B(n48107), .Z(n951) );
  AND U47877 ( .A(n48108), .B(n48109), .Z(n48107) );
  XNOR U47878 ( .A(p_input[1791]), .B(n48106), .Z(n48109) );
  XOR U47879 ( .A(n48106), .B(p_input[1759]), .Z(n48108) );
  XOR U47880 ( .A(n48110), .B(n48111), .Z(n48106) );
  AND U47881 ( .A(n48112), .B(n48113), .Z(n48111) );
  XNOR U47882 ( .A(p_input[1790]), .B(n48110), .Z(n48113) );
  XOR U47883 ( .A(n48110), .B(p_input[1758]), .Z(n48112) );
  XOR U47884 ( .A(n48114), .B(n48115), .Z(n48110) );
  AND U47885 ( .A(n48116), .B(n48117), .Z(n48115) );
  XNOR U47886 ( .A(p_input[1789]), .B(n48114), .Z(n48117) );
  XOR U47887 ( .A(n48114), .B(p_input[1757]), .Z(n48116) );
  XOR U47888 ( .A(n48118), .B(n48119), .Z(n48114) );
  AND U47889 ( .A(n48120), .B(n48121), .Z(n48119) );
  XNOR U47890 ( .A(p_input[1788]), .B(n48118), .Z(n48121) );
  XOR U47891 ( .A(n48118), .B(p_input[1756]), .Z(n48120) );
  XOR U47892 ( .A(n48122), .B(n48123), .Z(n48118) );
  AND U47893 ( .A(n48124), .B(n48125), .Z(n48123) );
  XNOR U47894 ( .A(p_input[1787]), .B(n48122), .Z(n48125) );
  XOR U47895 ( .A(n48122), .B(p_input[1755]), .Z(n48124) );
  XOR U47896 ( .A(n48126), .B(n48127), .Z(n48122) );
  AND U47897 ( .A(n48128), .B(n48129), .Z(n48127) );
  XNOR U47898 ( .A(p_input[1786]), .B(n48126), .Z(n48129) );
  XOR U47899 ( .A(n48126), .B(p_input[1754]), .Z(n48128) );
  XOR U47900 ( .A(n48130), .B(n48131), .Z(n48126) );
  AND U47901 ( .A(n48132), .B(n48133), .Z(n48131) );
  XNOR U47902 ( .A(p_input[1785]), .B(n48130), .Z(n48133) );
  XOR U47903 ( .A(n48130), .B(p_input[1753]), .Z(n48132) );
  XOR U47904 ( .A(n48134), .B(n48135), .Z(n48130) );
  AND U47905 ( .A(n48136), .B(n48137), .Z(n48135) );
  XNOR U47906 ( .A(p_input[1784]), .B(n48134), .Z(n48137) );
  XOR U47907 ( .A(n48134), .B(p_input[1752]), .Z(n48136) );
  XOR U47908 ( .A(n48138), .B(n48139), .Z(n48134) );
  AND U47909 ( .A(n48140), .B(n48141), .Z(n48139) );
  XNOR U47910 ( .A(p_input[1783]), .B(n48138), .Z(n48141) );
  XOR U47911 ( .A(n48138), .B(p_input[1751]), .Z(n48140) );
  XOR U47912 ( .A(n48142), .B(n48143), .Z(n48138) );
  AND U47913 ( .A(n48144), .B(n48145), .Z(n48143) );
  XNOR U47914 ( .A(p_input[1782]), .B(n48142), .Z(n48145) );
  XOR U47915 ( .A(n48142), .B(p_input[1750]), .Z(n48144) );
  XOR U47916 ( .A(n48146), .B(n48147), .Z(n48142) );
  AND U47917 ( .A(n48148), .B(n48149), .Z(n48147) );
  XNOR U47918 ( .A(p_input[1781]), .B(n48146), .Z(n48149) );
  XOR U47919 ( .A(n48146), .B(p_input[1749]), .Z(n48148) );
  XOR U47920 ( .A(n48150), .B(n48151), .Z(n48146) );
  AND U47921 ( .A(n48152), .B(n48153), .Z(n48151) );
  XNOR U47922 ( .A(p_input[1780]), .B(n48150), .Z(n48153) );
  XOR U47923 ( .A(n48150), .B(p_input[1748]), .Z(n48152) );
  XOR U47924 ( .A(n48154), .B(n48155), .Z(n48150) );
  AND U47925 ( .A(n48156), .B(n48157), .Z(n48155) );
  XNOR U47926 ( .A(p_input[1779]), .B(n48154), .Z(n48157) );
  XOR U47927 ( .A(n48154), .B(p_input[1747]), .Z(n48156) );
  XOR U47928 ( .A(n48158), .B(n48159), .Z(n48154) );
  AND U47929 ( .A(n48160), .B(n48161), .Z(n48159) );
  XNOR U47930 ( .A(p_input[1778]), .B(n48158), .Z(n48161) );
  XOR U47931 ( .A(n48158), .B(p_input[1746]), .Z(n48160) );
  XOR U47932 ( .A(n48162), .B(n48163), .Z(n48158) );
  AND U47933 ( .A(n48164), .B(n48165), .Z(n48163) );
  XNOR U47934 ( .A(p_input[1777]), .B(n48162), .Z(n48165) );
  XOR U47935 ( .A(n48162), .B(p_input[1745]), .Z(n48164) );
  XOR U47936 ( .A(n48166), .B(n48167), .Z(n48162) );
  AND U47937 ( .A(n48168), .B(n48169), .Z(n48167) );
  XNOR U47938 ( .A(p_input[1776]), .B(n48166), .Z(n48169) );
  XOR U47939 ( .A(n48166), .B(p_input[1744]), .Z(n48168) );
  XOR U47940 ( .A(n48170), .B(n48171), .Z(n48166) );
  AND U47941 ( .A(n48172), .B(n48173), .Z(n48171) );
  XNOR U47942 ( .A(p_input[1775]), .B(n48170), .Z(n48173) );
  XOR U47943 ( .A(n48170), .B(p_input[1743]), .Z(n48172) );
  XOR U47944 ( .A(n48174), .B(n48175), .Z(n48170) );
  AND U47945 ( .A(n48176), .B(n48177), .Z(n48175) );
  XNOR U47946 ( .A(p_input[1774]), .B(n48174), .Z(n48177) );
  XOR U47947 ( .A(n48174), .B(p_input[1742]), .Z(n48176) );
  XOR U47948 ( .A(n48178), .B(n48179), .Z(n48174) );
  AND U47949 ( .A(n48180), .B(n48181), .Z(n48179) );
  XNOR U47950 ( .A(p_input[1773]), .B(n48178), .Z(n48181) );
  XOR U47951 ( .A(n48178), .B(p_input[1741]), .Z(n48180) );
  XOR U47952 ( .A(n48182), .B(n48183), .Z(n48178) );
  AND U47953 ( .A(n48184), .B(n48185), .Z(n48183) );
  XNOR U47954 ( .A(p_input[1772]), .B(n48182), .Z(n48185) );
  XOR U47955 ( .A(n48182), .B(p_input[1740]), .Z(n48184) );
  XOR U47956 ( .A(n48186), .B(n48187), .Z(n48182) );
  AND U47957 ( .A(n48188), .B(n48189), .Z(n48187) );
  XNOR U47958 ( .A(p_input[1771]), .B(n48186), .Z(n48189) );
  XOR U47959 ( .A(n48186), .B(p_input[1739]), .Z(n48188) );
  XOR U47960 ( .A(n48190), .B(n48191), .Z(n48186) );
  AND U47961 ( .A(n48192), .B(n48193), .Z(n48191) );
  XNOR U47962 ( .A(p_input[1770]), .B(n48190), .Z(n48193) );
  XOR U47963 ( .A(n48190), .B(p_input[1738]), .Z(n48192) );
  XOR U47964 ( .A(n48194), .B(n48195), .Z(n48190) );
  AND U47965 ( .A(n48196), .B(n48197), .Z(n48195) );
  XNOR U47966 ( .A(p_input[1769]), .B(n48194), .Z(n48197) );
  XOR U47967 ( .A(n48194), .B(p_input[1737]), .Z(n48196) );
  XOR U47968 ( .A(n48198), .B(n48199), .Z(n48194) );
  AND U47969 ( .A(n48200), .B(n48201), .Z(n48199) );
  XNOR U47970 ( .A(p_input[1768]), .B(n48198), .Z(n48201) );
  XOR U47971 ( .A(n48198), .B(p_input[1736]), .Z(n48200) );
  XOR U47972 ( .A(n48202), .B(n48203), .Z(n48198) );
  AND U47973 ( .A(n48204), .B(n48205), .Z(n48203) );
  XNOR U47974 ( .A(p_input[1767]), .B(n48202), .Z(n48205) );
  XOR U47975 ( .A(n48202), .B(p_input[1735]), .Z(n48204) );
  XOR U47976 ( .A(n48206), .B(n48207), .Z(n48202) );
  AND U47977 ( .A(n48208), .B(n48209), .Z(n48207) );
  XNOR U47978 ( .A(p_input[1766]), .B(n48206), .Z(n48209) );
  XOR U47979 ( .A(n48206), .B(p_input[1734]), .Z(n48208) );
  XOR U47980 ( .A(n48210), .B(n48211), .Z(n48206) );
  AND U47981 ( .A(n48212), .B(n48213), .Z(n48211) );
  XNOR U47982 ( .A(p_input[1765]), .B(n48210), .Z(n48213) );
  XOR U47983 ( .A(n48210), .B(p_input[1733]), .Z(n48212) );
  XOR U47984 ( .A(n48214), .B(n48215), .Z(n48210) );
  AND U47985 ( .A(n48216), .B(n48217), .Z(n48215) );
  XNOR U47986 ( .A(p_input[1764]), .B(n48214), .Z(n48217) );
  XOR U47987 ( .A(n48214), .B(p_input[1732]), .Z(n48216) );
  XOR U47988 ( .A(n48218), .B(n48219), .Z(n48214) );
  AND U47989 ( .A(n48220), .B(n48221), .Z(n48219) );
  XNOR U47990 ( .A(p_input[1763]), .B(n48218), .Z(n48221) );
  XOR U47991 ( .A(n48218), .B(p_input[1731]), .Z(n48220) );
  XOR U47992 ( .A(n48222), .B(n48223), .Z(n48218) );
  AND U47993 ( .A(n48224), .B(n48225), .Z(n48223) );
  XNOR U47994 ( .A(p_input[1762]), .B(n48222), .Z(n48225) );
  XOR U47995 ( .A(n48222), .B(p_input[1730]), .Z(n48224) );
  XNOR U47996 ( .A(n48226), .B(n48227), .Z(n48222) );
  AND U47997 ( .A(n48228), .B(n48229), .Z(n48227) );
  XOR U47998 ( .A(p_input[1761]), .B(n48226), .Z(n48229) );
  XNOR U47999 ( .A(p_input[1729]), .B(n48226), .Z(n48228) );
  AND U48000 ( .A(p_input[1760]), .B(n48230), .Z(n48226) );
  IV U48001 ( .A(p_input[1728]), .Z(n48230) );
  XNOR U48002 ( .A(p_input[1664]), .B(n48231), .Z(n47824) );
  AND U48003 ( .A(n949), .B(n48232), .Z(n48231) );
  XOR U48004 ( .A(p_input[1696]), .B(p_input[1664]), .Z(n48232) );
  XOR U48005 ( .A(n48233), .B(n48234), .Z(n949) );
  AND U48006 ( .A(n48235), .B(n48236), .Z(n48234) );
  XNOR U48007 ( .A(p_input[1727]), .B(n48233), .Z(n48236) );
  XOR U48008 ( .A(n48233), .B(p_input[1695]), .Z(n48235) );
  XOR U48009 ( .A(n48237), .B(n48238), .Z(n48233) );
  AND U48010 ( .A(n48239), .B(n48240), .Z(n48238) );
  XNOR U48011 ( .A(p_input[1726]), .B(n48237), .Z(n48240) );
  XNOR U48012 ( .A(n48237), .B(n47839), .Z(n48239) );
  IV U48013 ( .A(p_input[1694]), .Z(n47839) );
  XOR U48014 ( .A(n48241), .B(n48242), .Z(n48237) );
  AND U48015 ( .A(n48243), .B(n48244), .Z(n48242) );
  XNOR U48016 ( .A(p_input[1725]), .B(n48241), .Z(n48244) );
  XNOR U48017 ( .A(n48241), .B(n47848), .Z(n48243) );
  IV U48018 ( .A(p_input[1693]), .Z(n47848) );
  XOR U48019 ( .A(n48245), .B(n48246), .Z(n48241) );
  AND U48020 ( .A(n48247), .B(n48248), .Z(n48246) );
  XNOR U48021 ( .A(p_input[1724]), .B(n48245), .Z(n48248) );
  XNOR U48022 ( .A(n48245), .B(n47857), .Z(n48247) );
  IV U48023 ( .A(p_input[1692]), .Z(n47857) );
  XOR U48024 ( .A(n48249), .B(n48250), .Z(n48245) );
  AND U48025 ( .A(n48251), .B(n48252), .Z(n48250) );
  XNOR U48026 ( .A(p_input[1723]), .B(n48249), .Z(n48252) );
  XNOR U48027 ( .A(n48249), .B(n47866), .Z(n48251) );
  IV U48028 ( .A(p_input[1691]), .Z(n47866) );
  XOR U48029 ( .A(n48253), .B(n48254), .Z(n48249) );
  AND U48030 ( .A(n48255), .B(n48256), .Z(n48254) );
  XNOR U48031 ( .A(p_input[1722]), .B(n48253), .Z(n48256) );
  XNOR U48032 ( .A(n48253), .B(n47875), .Z(n48255) );
  IV U48033 ( .A(p_input[1690]), .Z(n47875) );
  XOR U48034 ( .A(n48257), .B(n48258), .Z(n48253) );
  AND U48035 ( .A(n48259), .B(n48260), .Z(n48258) );
  XNOR U48036 ( .A(p_input[1721]), .B(n48257), .Z(n48260) );
  XNOR U48037 ( .A(n48257), .B(n47884), .Z(n48259) );
  IV U48038 ( .A(p_input[1689]), .Z(n47884) );
  XOR U48039 ( .A(n48261), .B(n48262), .Z(n48257) );
  AND U48040 ( .A(n48263), .B(n48264), .Z(n48262) );
  XNOR U48041 ( .A(p_input[1720]), .B(n48261), .Z(n48264) );
  XNOR U48042 ( .A(n48261), .B(n47893), .Z(n48263) );
  IV U48043 ( .A(p_input[1688]), .Z(n47893) );
  XOR U48044 ( .A(n48265), .B(n48266), .Z(n48261) );
  AND U48045 ( .A(n48267), .B(n48268), .Z(n48266) );
  XNOR U48046 ( .A(p_input[1719]), .B(n48265), .Z(n48268) );
  XNOR U48047 ( .A(n48265), .B(n47902), .Z(n48267) );
  IV U48048 ( .A(p_input[1687]), .Z(n47902) );
  XOR U48049 ( .A(n48269), .B(n48270), .Z(n48265) );
  AND U48050 ( .A(n48271), .B(n48272), .Z(n48270) );
  XNOR U48051 ( .A(p_input[1718]), .B(n48269), .Z(n48272) );
  XNOR U48052 ( .A(n48269), .B(n47911), .Z(n48271) );
  IV U48053 ( .A(p_input[1686]), .Z(n47911) );
  XOR U48054 ( .A(n48273), .B(n48274), .Z(n48269) );
  AND U48055 ( .A(n48275), .B(n48276), .Z(n48274) );
  XNOR U48056 ( .A(p_input[1717]), .B(n48273), .Z(n48276) );
  XNOR U48057 ( .A(n48273), .B(n47920), .Z(n48275) );
  IV U48058 ( .A(p_input[1685]), .Z(n47920) );
  XOR U48059 ( .A(n48277), .B(n48278), .Z(n48273) );
  AND U48060 ( .A(n48279), .B(n48280), .Z(n48278) );
  XNOR U48061 ( .A(p_input[1716]), .B(n48277), .Z(n48280) );
  XNOR U48062 ( .A(n48277), .B(n47929), .Z(n48279) );
  IV U48063 ( .A(p_input[1684]), .Z(n47929) );
  XOR U48064 ( .A(n48281), .B(n48282), .Z(n48277) );
  AND U48065 ( .A(n48283), .B(n48284), .Z(n48282) );
  XNOR U48066 ( .A(p_input[1715]), .B(n48281), .Z(n48284) );
  XNOR U48067 ( .A(n48281), .B(n47938), .Z(n48283) );
  IV U48068 ( .A(p_input[1683]), .Z(n47938) );
  XOR U48069 ( .A(n48285), .B(n48286), .Z(n48281) );
  AND U48070 ( .A(n48287), .B(n48288), .Z(n48286) );
  XNOR U48071 ( .A(p_input[1714]), .B(n48285), .Z(n48288) );
  XNOR U48072 ( .A(n48285), .B(n47947), .Z(n48287) );
  IV U48073 ( .A(p_input[1682]), .Z(n47947) );
  XOR U48074 ( .A(n48289), .B(n48290), .Z(n48285) );
  AND U48075 ( .A(n48291), .B(n48292), .Z(n48290) );
  XNOR U48076 ( .A(p_input[1713]), .B(n48289), .Z(n48292) );
  XNOR U48077 ( .A(n48289), .B(n47956), .Z(n48291) );
  IV U48078 ( .A(p_input[1681]), .Z(n47956) );
  XOR U48079 ( .A(n48293), .B(n48294), .Z(n48289) );
  AND U48080 ( .A(n48295), .B(n48296), .Z(n48294) );
  XNOR U48081 ( .A(p_input[1712]), .B(n48293), .Z(n48296) );
  XNOR U48082 ( .A(n48293), .B(n47965), .Z(n48295) );
  IV U48083 ( .A(p_input[1680]), .Z(n47965) );
  XOR U48084 ( .A(n48297), .B(n48298), .Z(n48293) );
  AND U48085 ( .A(n48299), .B(n48300), .Z(n48298) );
  XNOR U48086 ( .A(p_input[1711]), .B(n48297), .Z(n48300) );
  XNOR U48087 ( .A(n48297), .B(n47974), .Z(n48299) );
  IV U48088 ( .A(p_input[1679]), .Z(n47974) );
  XOR U48089 ( .A(n48301), .B(n48302), .Z(n48297) );
  AND U48090 ( .A(n48303), .B(n48304), .Z(n48302) );
  XNOR U48091 ( .A(p_input[1710]), .B(n48301), .Z(n48304) );
  XNOR U48092 ( .A(n48301), .B(n47983), .Z(n48303) );
  IV U48093 ( .A(p_input[1678]), .Z(n47983) );
  XOR U48094 ( .A(n48305), .B(n48306), .Z(n48301) );
  AND U48095 ( .A(n48307), .B(n48308), .Z(n48306) );
  XNOR U48096 ( .A(p_input[1709]), .B(n48305), .Z(n48308) );
  XNOR U48097 ( .A(n48305), .B(n47992), .Z(n48307) );
  IV U48098 ( .A(p_input[1677]), .Z(n47992) );
  XOR U48099 ( .A(n48309), .B(n48310), .Z(n48305) );
  AND U48100 ( .A(n48311), .B(n48312), .Z(n48310) );
  XNOR U48101 ( .A(p_input[1708]), .B(n48309), .Z(n48312) );
  XNOR U48102 ( .A(n48309), .B(n48001), .Z(n48311) );
  IV U48103 ( .A(p_input[1676]), .Z(n48001) );
  XOR U48104 ( .A(n48313), .B(n48314), .Z(n48309) );
  AND U48105 ( .A(n48315), .B(n48316), .Z(n48314) );
  XNOR U48106 ( .A(p_input[1707]), .B(n48313), .Z(n48316) );
  XNOR U48107 ( .A(n48313), .B(n48010), .Z(n48315) );
  IV U48108 ( .A(p_input[1675]), .Z(n48010) );
  XOR U48109 ( .A(n48317), .B(n48318), .Z(n48313) );
  AND U48110 ( .A(n48319), .B(n48320), .Z(n48318) );
  XNOR U48111 ( .A(p_input[1706]), .B(n48317), .Z(n48320) );
  XNOR U48112 ( .A(n48317), .B(n48019), .Z(n48319) );
  IV U48113 ( .A(p_input[1674]), .Z(n48019) );
  XOR U48114 ( .A(n48321), .B(n48322), .Z(n48317) );
  AND U48115 ( .A(n48323), .B(n48324), .Z(n48322) );
  XNOR U48116 ( .A(p_input[1705]), .B(n48321), .Z(n48324) );
  XNOR U48117 ( .A(n48321), .B(n48028), .Z(n48323) );
  IV U48118 ( .A(p_input[1673]), .Z(n48028) );
  XOR U48119 ( .A(n48325), .B(n48326), .Z(n48321) );
  AND U48120 ( .A(n48327), .B(n48328), .Z(n48326) );
  XNOR U48121 ( .A(p_input[1704]), .B(n48325), .Z(n48328) );
  XNOR U48122 ( .A(n48325), .B(n48037), .Z(n48327) );
  IV U48123 ( .A(p_input[1672]), .Z(n48037) );
  XOR U48124 ( .A(n48329), .B(n48330), .Z(n48325) );
  AND U48125 ( .A(n48331), .B(n48332), .Z(n48330) );
  XNOR U48126 ( .A(p_input[1703]), .B(n48329), .Z(n48332) );
  XNOR U48127 ( .A(n48329), .B(n48046), .Z(n48331) );
  IV U48128 ( .A(p_input[1671]), .Z(n48046) );
  XOR U48129 ( .A(n48333), .B(n48334), .Z(n48329) );
  AND U48130 ( .A(n48335), .B(n48336), .Z(n48334) );
  XNOR U48131 ( .A(p_input[1702]), .B(n48333), .Z(n48336) );
  XNOR U48132 ( .A(n48333), .B(n48055), .Z(n48335) );
  IV U48133 ( .A(p_input[1670]), .Z(n48055) );
  XOR U48134 ( .A(n48337), .B(n48338), .Z(n48333) );
  AND U48135 ( .A(n48339), .B(n48340), .Z(n48338) );
  XNOR U48136 ( .A(p_input[1701]), .B(n48337), .Z(n48340) );
  XNOR U48137 ( .A(n48337), .B(n48064), .Z(n48339) );
  IV U48138 ( .A(p_input[1669]), .Z(n48064) );
  XOR U48139 ( .A(n48341), .B(n48342), .Z(n48337) );
  AND U48140 ( .A(n48343), .B(n48344), .Z(n48342) );
  XNOR U48141 ( .A(p_input[1700]), .B(n48341), .Z(n48344) );
  XNOR U48142 ( .A(n48341), .B(n48073), .Z(n48343) );
  IV U48143 ( .A(p_input[1668]), .Z(n48073) );
  XOR U48144 ( .A(n48345), .B(n48346), .Z(n48341) );
  AND U48145 ( .A(n48347), .B(n48348), .Z(n48346) );
  XNOR U48146 ( .A(p_input[1699]), .B(n48345), .Z(n48348) );
  XNOR U48147 ( .A(n48345), .B(n48082), .Z(n48347) );
  IV U48148 ( .A(p_input[1667]), .Z(n48082) );
  XOR U48149 ( .A(n48349), .B(n48350), .Z(n48345) );
  AND U48150 ( .A(n48351), .B(n48352), .Z(n48350) );
  XNOR U48151 ( .A(p_input[1698]), .B(n48349), .Z(n48352) );
  XNOR U48152 ( .A(n48349), .B(n48091), .Z(n48351) );
  IV U48153 ( .A(p_input[1666]), .Z(n48091) );
  XNOR U48154 ( .A(n48353), .B(n48354), .Z(n48349) );
  AND U48155 ( .A(n48355), .B(n48356), .Z(n48354) );
  XOR U48156 ( .A(p_input[1697]), .B(n48353), .Z(n48356) );
  XNOR U48157 ( .A(p_input[1665]), .B(n48353), .Z(n48355) );
  AND U48158 ( .A(p_input[1696]), .B(n48357), .Z(n48353) );
  IV U48159 ( .A(p_input[1664]), .Z(n48357) );
  XOR U48160 ( .A(n48358), .B(n48359), .Z(n47447) );
  AND U48161 ( .A(n624), .B(n48360), .Z(n48359) );
  XNOR U48162 ( .A(n48361), .B(n48358), .Z(n48360) );
  XOR U48163 ( .A(n48362), .B(n48363), .Z(n624) );
  AND U48164 ( .A(n48364), .B(n48365), .Z(n48363) );
  XNOR U48165 ( .A(n47462), .B(n48362), .Z(n48365) );
  AND U48166 ( .A(p_input[1663]), .B(p_input[1631]), .Z(n47462) );
  XNOR U48167 ( .A(n48362), .B(n47459), .Z(n48364) );
  IV U48168 ( .A(n48366), .Z(n47459) );
  AND U48169 ( .A(p_input[1567]), .B(p_input[1599]), .Z(n48366) );
  XOR U48170 ( .A(n48367), .B(n48368), .Z(n48362) );
  AND U48171 ( .A(n48369), .B(n48370), .Z(n48368) );
  XOR U48172 ( .A(n48367), .B(n47474), .Z(n48370) );
  XNOR U48173 ( .A(p_input[1630]), .B(n48371), .Z(n47474) );
  AND U48174 ( .A(n955), .B(n48372), .Z(n48371) );
  XOR U48175 ( .A(p_input[1662]), .B(p_input[1630]), .Z(n48372) );
  XNOR U48176 ( .A(n47471), .B(n48367), .Z(n48369) );
  XOR U48177 ( .A(n48373), .B(n48374), .Z(n47471) );
  AND U48178 ( .A(n952), .B(n48375), .Z(n48374) );
  XOR U48179 ( .A(p_input[1598]), .B(p_input[1566]), .Z(n48375) );
  XOR U48180 ( .A(n48376), .B(n48377), .Z(n48367) );
  AND U48181 ( .A(n48378), .B(n48379), .Z(n48377) );
  XOR U48182 ( .A(n48376), .B(n47486), .Z(n48379) );
  XNOR U48183 ( .A(p_input[1629]), .B(n48380), .Z(n47486) );
  AND U48184 ( .A(n955), .B(n48381), .Z(n48380) );
  XOR U48185 ( .A(p_input[1661]), .B(p_input[1629]), .Z(n48381) );
  XNOR U48186 ( .A(n47483), .B(n48376), .Z(n48378) );
  XOR U48187 ( .A(n48382), .B(n48383), .Z(n47483) );
  AND U48188 ( .A(n952), .B(n48384), .Z(n48383) );
  XOR U48189 ( .A(p_input[1597]), .B(p_input[1565]), .Z(n48384) );
  XOR U48190 ( .A(n48385), .B(n48386), .Z(n48376) );
  AND U48191 ( .A(n48387), .B(n48388), .Z(n48386) );
  XOR U48192 ( .A(n48385), .B(n47498), .Z(n48388) );
  XNOR U48193 ( .A(p_input[1628]), .B(n48389), .Z(n47498) );
  AND U48194 ( .A(n955), .B(n48390), .Z(n48389) );
  XOR U48195 ( .A(p_input[1660]), .B(p_input[1628]), .Z(n48390) );
  XNOR U48196 ( .A(n47495), .B(n48385), .Z(n48387) );
  XOR U48197 ( .A(n48391), .B(n48392), .Z(n47495) );
  AND U48198 ( .A(n952), .B(n48393), .Z(n48392) );
  XOR U48199 ( .A(p_input[1596]), .B(p_input[1564]), .Z(n48393) );
  XOR U48200 ( .A(n48394), .B(n48395), .Z(n48385) );
  AND U48201 ( .A(n48396), .B(n48397), .Z(n48395) );
  XOR U48202 ( .A(n48394), .B(n47510), .Z(n48397) );
  XNOR U48203 ( .A(p_input[1627]), .B(n48398), .Z(n47510) );
  AND U48204 ( .A(n955), .B(n48399), .Z(n48398) );
  XOR U48205 ( .A(p_input[1659]), .B(p_input[1627]), .Z(n48399) );
  XNOR U48206 ( .A(n47507), .B(n48394), .Z(n48396) );
  XOR U48207 ( .A(n48400), .B(n48401), .Z(n47507) );
  AND U48208 ( .A(n952), .B(n48402), .Z(n48401) );
  XOR U48209 ( .A(p_input[1595]), .B(p_input[1563]), .Z(n48402) );
  XOR U48210 ( .A(n48403), .B(n48404), .Z(n48394) );
  AND U48211 ( .A(n48405), .B(n48406), .Z(n48404) );
  XOR U48212 ( .A(n48403), .B(n47522), .Z(n48406) );
  XNOR U48213 ( .A(p_input[1626]), .B(n48407), .Z(n47522) );
  AND U48214 ( .A(n955), .B(n48408), .Z(n48407) );
  XOR U48215 ( .A(p_input[1658]), .B(p_input[1626]), .Z(n48408) );
  XNOR U48216 ( .A(n47519), .B(n48403), .Z(n48405) );
  XOR U48217 ( .A(n48409), .B(n48410), .Z(n47519) );
  AND U48218 ( .A(n952), .B(n48411), .Z(n48410) );
  XOR U48219 ( .A(p_input[1594]), .B(p_input[1562]), .Z(n48411) );
  XOR U48220 ( .A(n48412), .B(n48413), .Z(n48403) );
  AND U48221 ( .A(n48414), .B(n48415), .Z(n48413) );
  XOR U48222 ( .A(n48412), .B(n47534), .Z(n48415) );
  XNOR U48223 ( .A(p_input[1625]), .B(n48416), .Z(n47534) );
  AND U48224 ( .A(n955), .B(n48417), .Z(n48416) );
  XOR U48225 ( .A(p_input[1657]), .B(p_input[1625]), .Z(n48417) );
  XNOR U48226 ( .A(n47531), .B(n48412), .Z(n48414) );
  XOR U48227 ( .A(n48418), .B(n48419), .Z(n47531) );
  AND U48228 ( .A(n952), .B(n48420), .Z(n48419) );
  XOR U48229 ( .A(p_input[1593]), .B(p_input[1561]), .Z(n48420) );
  XOR U48230 ( .A(n48421), .B(n48422), .Z(n48412) );
  AND U48231 ( .A(n48423), .B(n48424), .Z(n48422) );
  XOR U48232 ( .A(n48421), .B(n47546), .Z(n48424) );
  XNOR U48233 ( .A(p_input[1624]), .B(n48425), .Z(n47546) );
  AND U48234 ( .A(n955), .B(n48426), .Z(n48425) );
  XOR U48235 ( .A(p_input[1656]), .B(p_input[1624]), .Z(n48426) );
  XNOR U48236 ( .A(n47543), .B(n48421), .Z(n48423) );
  XOR U48237 ( .A(n48427), .B(n48428), .Z(n47543) );
  AND U48238 ( .A(n952), .B(n48429), .Z(n48428) );
  XOR U48239 ( .A(p_input[1592]), .B(p_input[1560]), .Z(n48429) );
  XOR U48240 ( .A(n48430), .B(n48431), .Z(n48421) );
  AND U48241 ( .A(n48432), .B(n48433), .Z(n48431) );
  XOR U48242 ( .A(n48430), .B(n47558), .Z(n48433) );
  XNOR U48243 ( .A(p_input[1623]), .B(n48434), .Z(n47558) );
  AND U48244 ( .A(n955), .B(n48435), .Z(n48434) );
  XOR U48245 ( .A(p_input[1655]), .B(p_input[1623]), .Z(n48435) );
  XNOR U48246 ( .A(n47555), .B(n48430), .Z(n48432) );
  XOR U48247 ( .A(n48436), .B(n48437), .Z(n47555) );
  AND U48248 ( .A(n952), .B(n48438), .Z(n48437) );
  XOR U48249 ( .A(p_input[1591]), .B(p_input[1559]), .Z(n48438) );
  XOR U48250 ( .A(n48439), .B(n48440), .Z(n48430) );
  AND U48251 ( .A(n48441), .B(n48442), .Z(n48440) );
  XOR U48252 ( .A(n48439), .B(n47570), .Z(n48442) );
  XNOR U48253 ( .A(p_input[1622]), .B(n48443), .Z(n47570) );
  AND U48254 ( .A(n955), .B(n48444), .Z(n48443) );
  XOR U48255 ( .A(p_input[1654]), .B(p_input[1622]), .Z(n48444) );
  XNOR U48256 ( .A(n47567), .B(n48439), .Z(n48441) );
  XOR U48257 ( .A(n48445), .B(n48446), .Z(n47567) );
  AND U48258 ( .A(n952), .B(n48447), .Z(n48446) );
  XOR U48259 ( .A(p_input[1590]), .B(p_input[1558]), .Z(n48447) );
  XOR U48260 ( .A(n48448), .B(n48449), .Z(n48439) );
  AND U48261 ( .A(n48450), .B(n48451), .Z(n48449) );
  XOR U48262 ( .A(n48448), .B(n47582), .Z(n48451) );
  XNOR U48263 ( .A(p_input[1621]), .B(n48452), .Z(n47582) );
  AND U48264 ( .A(n955), .B(n48453), .Z(n48452) );
  XOR U48265 ( .A(p_input[1653]), .B(p_input[1621]), .Z(n48453) );
  XNOR U48266 ( .A(n47579), .B(n48448), .Z(n48450) );
  XOR U48267 ( .A(n48454), .B(n48455), .Z(n47579) );
  AND U48268 ( .A(n952), .B(n48456), .Z(n48455) );
  XOR U48269 ( .A(p_input[1589]), .B(p_input[1557]), .Z(n48456) );
  XOR U48270 ( .A(n48457), .B(n48458), .Z(n48448) );
  AND U48271 ( .A(n48459), .B(n48460), .Z(n48458) );
  XOR U48272 ( .A(n48457), .B(n47594), .Z(n48460) );
  XNOR U48273 ( .A(p_input[1620]), .B(n48461), .Z(n47594) );
  AND U48274 ( .A(n955), .B(n48462), .Z(n48461) );
  XOR U48275 ( .A(p_input[1652]), .B(p_input[1620]), .Z(n48462) );
  XNOR U48276 ( .A(n47591), .B(n48457), .Z(n48459) );
  XOR U48277 ( .A(n48463), .B(n48464), .Z(n47591) );
  AND U48278 ( .A(n952), .B(n48465), .Z(n48464) );
  XOR U48279 ( .A(p_input[1588]), .B(p_input[1556]), .Z(n48465) );
  XOR U48280 ( .A(n48466), .B(n48467), .Z(n48457) );
  AND U48281 ( .A(n48468), .B(n48469), .Z(n48467) );
  XOR U48282 ( .A(n48466), .B(n47606), .Z(n48469) );
  XNOR U48283 ( .A(p_input[1619]), .B(n48470), .Z(n47606) );
  AND U48284 ( .A(n955), .B(n48471), .Z(n48470) );
  XOR U48285 ( .A(p_input[1651]), .B(p_input[1619]), .Z(n48471) );
  XNOR U48286 ( .A(n47603), .B(n48466), .Z(n48468) );
  XOR U48287 ( .A(n48472), .B(n48473), .Z(n47603) );
  AND U48288 ( .A(n952), .B(n48474), .Z(n48473) );
  XOR U48289 ( .A(p_input[1587]), .B(p_input[1555]), .Z(n48474) );
  XOR U48290 ( .A(n48475), .B(n48476), .Z(n48466) );
  AND U48291 ( .A(n48477), .B(n48478), .Z(n48476) );
  XOR U48292 ( .A(n48475), .B(n47618), .Z(n48478) );
  XNOR U48293 ( .A(p_input[1618]), .B(n48479), .Z(n47618) );
  AND U48294 ( .A(n955), .B(n48480), .Z(n48479) );
  XOR U48295 ( .A(p_input[1650]), .B(p_input[1618]), .Z(n48480) );
  XNOR U48296 ( .A(n47615), .B(n48475), .Z(n48477) );
  XOR U48297 ( .A(n48481), .B(n48482), .Z(n47615) );
  AND U48298 ( .A(n952), .B(n48483), .Z(n48482) );
  XOR U48299 ( .A(p_input[1586]), .B(p_input[1554]), .Z(n48483) );
  XOR U48300 ( .A(n48484), .B(n48485), .Z(n48475) );
  AND U48301 ( .A(n48486), .B(n48487), .Z(n48485) );
  XOR U48302 ( .A(n48484), .B(n47630), .Z(n48487) );
  XNOR U48303 ( .A(p_input[1617]), .B(n48488), .Z(n47630) );
  AND U48304 ( .A(n955), .B(n48489), .Z(n48488) );
  XOR U48305 ( .A(p_input[1649]), .B(p_input[1617]), .Z(n48489) );
  XNOR U48306 ( .A(n47627), .B(n48484), .Z(n48486) );
  XOR U48307 ( .A(n48490), .B(n48491), .Z(n47627) );
  AND U48308 ( .A(n952), .B(n48492), .Z(n48491) );
  XOR U48309 ( .A(p_input[1585]), .B(p_input[1553]), .Z(n48492) );
  XOR U48310 ( .A(n48493), .B(n48494), .Z(n48484) );
  AND U48311 ( .A(n48495), .B(n48496), .Z(n48494) );
  XOR U48312 ( .A(n48493), .B(n47642), .Z(n48496) );
  XNOR U48313 ( .A(p_input[1616]), .B(n48497), .Z(n47642) );
  AND U48314 ( .A(n955), .B(n48498), .Z(n48497) );
  XOR U48315 ( .A(p_input[1648]), .B(p_input[1616]), .Z(n48498) );
  XNOR U48316 ( .A(n47639), .B(n48493), .Z(n48495) );
  XOR U48317 ( .A(n48499), .B(n48500), .Z(n47639) );
  AND U48318 ( .A(n952), .B(n48501), .Z(n48500) );
  XOR U48319 ( .A(p_input[1584]), .B(p_input[1552]), .Z(n48501) );
  XOR U48320 ( .A(n48502), .B(n48503), .Z(n48493) );
  AND U48321 ( .A(n48504), .B(n48505), .Z(n48503) );
  XOR U48322 ( .A(n48502), .B(n47654), .Z(n48505) );
  XNOR U48323 ( .A(p_input[1615]), .B(n48506), .Z(n47654) );
  AND U48324 ( .A(n955), .B(n48507), .Z(n48506) );
  XOR U48325 ( .A(p_input[1647]), .B(p_input[1615]), .Z(n48507) );
  XNOR U48326 ( .A(n47651), .B(n48502), .Z(n48504) );
  XOR U48327 ( .A(n48508), .B(n48509), .Z(n47651) );
  AND U48328 ( .A(n952), .B(n48510), .Z(n48509) );
  XOR U48329 ( .A(p_input[1583]), .B(p_input[1551]), .Z(n48510) );
  XOR U48330 ( .A(n48511), .B(n48512), .Z(n48502) );
  AND U48331 ( .A(n48513), .B(n48514), .Z(n48512) );
  XOR U48332 ( .A(n48511), .B(n47666), .Z(n48514) );
  XNOR U48333 ( .A(p_input[1614]), .B(n48515), .Z(n47666) );
  AND U48334 ( .A(n955), .B(n48516), .Z(n48515) );
  XOR U48335 ( .A(p_input[1646]), .B(p_input[1614]), .Z(n48516) );
  XNOR U48336 ( .A(n47663), .B(n48511), .Z(n48513) );
  XOR U48337 ( .A(n48517), .B(n48518), .Z(n47663) );
  AND U48338 ( .A(n952), .B(n48519), .Z(n48518) );
  XOR U48339 ( .A(p_input[1582]), .B(p_input[1550]), .Z(n48519) );
  XOR U48340 ( .A(n48520), .B(n48521), .Z(n48511) );
  AND U48341 ( .A(n48522), .B(n48523), .Z(n48521) );
  XOR U48342 ( .A(n48520), .B(n47678), .Z(n48523) );
  XNOR U48343 ( .A(p_input[1613]), .B(n48524), .Z(n47678) );
  AND U48344 ( .A(n955), .B(n48525), .Z(n48524) );
  XOR U48345 ( .A(p_input[1645]), .B(p_input[1613]), .Z(n48525) );
  XNOR U48346 ( .A(n47675), .B(n48520), .Z(n48522) );
  XOR U48347 ( .A(n48526), .B(n48527), .Z(n47675) );
  AND U48348 ( .A(n952), .B(n48528), .Z(n48527) );
  XOR U48349 ( .A(p_input[1581]), .B(p_input[1549]), .Z(n48528) );
  XOR U48350 ( .A(n48529), .B(n48530), .Z(n48520) );
  AND U48351 ( .A(n48531), .B(n48532), .Z(n48530) );
  XOR U48352 ( .A(n48529), .B(n47690), .Z(n48532) );
  XNOR U48353 ( .A(p_input[1612]), .B(n48533), .Z(n47690) );
  AND U48354 ( .A(n955), .B(n48534), .Z(n48533) );
  XOR U48355 ( .A(p_input[1644]), .B(p_input[1612]), .Z(n48534) );
  XNOR U48356 ( .A(n47687), .B(n48529), .Z(n48531) );
  XOR U48357 ( .A(n48535), .B(n48536), .Z(n47687) );
  AND U48358 ( .A(n952), .B(n48537), .Z(n48536) );
  XOR U48359 ( .A(p_input[1580]), .B(p_input[1548]), .Z(n48537) );
  XOR U48360 ( .A(n48538), .B(n48539), .Z(n48529) );
  AND U48361 ( .A(n48540), .B(n48541), .Z(n48539) );
  XOR U48362 ( .A(n48538), .B(n47702), .Z(n48541) );
  XNOR U48363 ( .A(p_input[1611]), .B(n48542), .Z(n47702) );
  AND U48364 ( .A(n955), .B(n48543), .Z(n48542) );
  XOR U48365 ( .A(p_input[1643]), .B(p_input[1611]), .Z(n48543) );
  XNOR U48366 ( .A(n47699), .B(n48538), .Z(n48540) );
  XOR U48367 ( .A(n48544), .B(n48545), .Z(n47699) );
  AND U48368 ( .A(n952), .B(n48546), .Z(n48545) );
  XOR U48369 ( .A(p_input[1579]), .B(p_input[1547]), .Z(n48546) );
  XOR U48370 ( .A(n48547), .B(n48548), .Z(n48538) );
  AND U48371 ( .A(n48549), .B(n48550), .Z(n48548) );
  XOR U48372 ( .A(n48547), .B(n47714), .Z(n48550) );
  XNOR U48373 ( .A(p_input[1610]), .B(n48551), .Z(n47714) );
  AND U48374 ( .A(n955), .B(n48552), .Z(n48551) );
  XOR U48375 ( .A(p_input[1642]), .B(p_input[1610]), .Z(n48552) );
  XNOR U48376 ( .A(n47711), .B(n48547), .Z(n48549) );
  XOR U48377 ( .A(n48553), .B(n48554), .Z(n47711) );
  AND U48378 ( .A(n952), .B(n48555), .Z(n48554) );
  XOR U48379 ( .A(p_input[1578]), .B(p_input[1546]), .Z(n48555) );
  XOR U48380 ( .A(n48556), .B(n48557), .Z(n48547) );
  AND U48381 ( .A(n48558), .B(n48559), .Z(n48557) );
  XOR U48382 ( .A(n48556), .B(n47726), .Z(n48559) );
  XNOR U48383 ( .A(p_input[1609]), .B(n48560), .Z(n47726) );
  AND U48384 ( .A(n955), .B(n48561), .Z(n48560) );
  XOR U48385 ( .A(p_input[1641]), .B(p_input[1609]), .Z(n48561) );
  XNOR U48386 ( .A(n47723), .B(n48556), .Z(n48558) );
  XOR U48387 ( .A(n48562), .B(n48563), .Z(n47723) );
  AND U48388 ( .A(n952), .B(n48564), .Z(n48563) );
  XOR U48389 ( .A(p_input[1577]), .B(p_input[1545]), .Z(n48564) );
  XOR U48390 ( .A(n48565), .B(n48566), .Z(n48556) );
  AND U48391 ( .A(n48567), .B(n48568), .Z(n48566) );
  XOR U48392 ( .A(n48565), .B(n47738), .Z(n48568) );
  XNOR U48393 ( .A(p_input[1608]), .B(n48569), .Z(n47738) );
  AND U48394 ( .A(n955), .B(n48570), .Z(n48569) );
  XOR U48395 ( .A(p_input[1640]), .B(p_input[1608]), .Z(n48570) );
  XNOR U48396 ( .A(n47735), .B(n48565), .Z(n48567) );
  XOR U48397 ( .A(n48571), .B(n48572), .Z(n47735) );
  AND U48398 ( .A(n952), .B(n48573), .Z(n48572) );
  XOR U48399 ( .A(p_input[1576]), .B(p_input[1544]), .Z(n48573) );
  XOR U48400 ( .A(n48574), .B(n48575), .Z(n48565) );
  AND U48401 ( .A(n48576), .B(n48577), .Z(n48575) );
  XOR U48402 ( .A(n48574), .B(n47750), .Z(n48577) );
  XNOR U48403 ( .A(p_input[1607]), .B(n48578), .Z(n47750) );
  AND U48404 ( .A(n955), .B(n48579), .Z(n48578) );
  XOR U48405 ( .A(p_input[1639]), .B(p_input[1607]), .Z(n48579) );
  XNOR U48406 ( .A(n47747), .B(n48574), .Z(n48576) );
  XOR U48407 ( .A(n48580), .B(n48581), .Z(n47747) );
  AND U48408 ( .A(n952), .B(n48582), .Z(n48581) );
  XOR U48409 ( .A(p_input[1575]), .B(p_input[1543]), .Z(n48582) );
  XOR U48410 ( .A(n48583), .B(n48584), .Z(n48574) );
  AND U48411 ( .A(n48585), .B(n48586), .Z(n48584) );
  XOR U48412 ( .A(n48583), .B(n47762), .Z(n48586) );
  XNOR U48413 ( .A(p_input[1606]), .B(n48587), .Z(n47762) );
  AND U48414 ( .A(n955), .B(n48588), .Z(n48587) );
  XOR U48415 ( .A(p_input[1638]), .B(p_input[1606]), .Z(n48588) );
  XNOR U48416 ( .A(n47759), .B(n48583), .Z(n48585) );
  XOR U48417 ( .A(n48589), .B(n48590), .Z(n47759) );
  AND U48418 ( .A(n952), .B(n48591), .Z(n48590) );
  XOR U48419 ( .A(p_input[1574]), .B(p_input[1542]), .Z(n48591) );
  XOR U48420 ( .A(n48592), .B(n48593), .Z(n48583) );
  AND U48421 ( .A(n48594), .B(n48595), .Z(n48593) );
  XOR U48422 ( .A(n48592), .B(n47774), .Z(n48595) );
  XNOR U48423 ( .A(p_input[1605]), .B(n48596), .Z(n47774) );
  AND U48424 ( .A(n955), .B(n48597), .Z(n48596) );
  XOR U48425 ( .A(p_input[1637]), .B(p_input[1605]), .Z(n48597) );
  XNOR U48426 ( .A(n47771), .B(n48592), .Z(n48594) );
  XOR U48427 ( .A(n48598), .B(n48599), .Z(n47771) );
  AND U48428 ( .A(n952), .B(n48600), .Z(n48599) );
  XOR U48429 ( .A(p_input[1573]), .B(p_input[1541]), .Z(n48600) );
  XOR U48430 ( .A(n48601), .B(n48602), .Z(n48592) );
  AND U48431 ( .A(n48603), .B(n48604), .Z(n48602) );
  XOR U48432 ( .A(n48601), .B(n47786), .Z(n48604) );
  XNOR U48433 ( .A(p_input[1604]), .B(n48605), .Z(n47786) );
  AND U48434 ( .A(n955), .B(n48606), .Z(n48605) );
  XOR U48435 ( .A(p_input[1636]), .B(p_input[1604]), .Z(n48606) );
  XNOR U48436 ( .A(n47783), .B(n48601), .Z(n48603) );
  XOR U48437 ( .A(n48607), .B(n48608), .Z(n47783) );
  AND U48438 ( .A(n952), .B(n48609), .Z(n48608) );
  XOR U48439 ( .A(p_input[1572]), .B(p_input[1540]), .Z(n48609) );
  XOR U48440 ( .A(n48610), .B(n48611), .Z(n48601) );
  AND U48441 ( .A(n48612), .B(n48613), .Z(n48611) );
  XOR U48442 ( .A(n48610), .B(n47798), .Z(n48613) );
  XNOR U48443 ( .A(p_input[1603]), .B(n48614), .Z(n47798) );
  AND U48444 ( .A(n955), .B(n48615), .Z(n48614) );
  XOR U48445 ( .A(p_input[1635]), .B(p_input[1603]), .Z(n48615) );
  XNOR U48446 ( .A(n47795), .B(n48610), .Z(n48612) );
  XOR U48447 ( .A(n48616), .B(n48617), .Z(n47795) );
  AND U48448 ( .A(n952), .B(n48618), .Z(n48617) );
  XOR U48449 ( .A(p_input[1571]), .B(p_input[1539]), .Z(n48618) );
  XOR U48450 ( .A(n48619), .B(n48620), .Z(n48610) );
  AND U48451 ( .A(n48621), .B(n48622), .Z(n48620) );
  XOR U48452 ( .A(n48619), .B(n47810), .Z(n48622) );
  XNOR U48453 ( .A(p_input[1602]), .B(n48623), .Z(n47810) );
  AND U48454 ( .A(n955), .B(n48624), .Z(n48623) );
  XOR U48455 ( .A(p_input[1634]), .B(p_input[1602]), .Z(n48624) );
  XNOR U48456 ( .A(n47807), .B(n48619), .Z(n48621) );
  XOR U48457 ( .A(n48625), .B(n48626), .Z(n47807) );
  AND U48458 ( .A(n952), .B(n48627), .Z(n48626) );
  XOR U48459 ( .A(p_input[1570]), .B(p_input[1538]), .Z(n48627) );
  XOR U48460 ( .A(n48628), .B(n48629), .Z(n48619) );
  AND U48461 ( .A(n48630), .B(n48631), .Z(n48629) );
  XNOR U48462 ( .A(n48632), .B(n47823), .Z(n48631) );
  XNOR U48463 ( .A(p_input[1601]), .B(n48633), .Z(n47823) );
  AND U48464 ( .A(n955), .B(n48634), .Z(n48633) );
  XNOR U48465 ( .A(p_input[1633]), .B(n48635), .Z(n48634) );
  IV U48466 ( .A(p_input[1601]), .Z(n48635) );
  XNOR U48467 ( .A(n47820), .B(n48628), .Z(n48630) );
  XNOR U48468 ( .A(p_input[1537]), .B(n48636), .Z(n47820) );
  AND U48469 ( .A(n952), .B(n48637), .Z(n48636) );
  XOR U48470 ( .A(p_input[1569]), .B(p_input[1537]), .Z(n48637) );
  IV U48471 ( .A(n48632), .Z(n48628) );
  AND U48472 ( .A(n48358), .B(n48361), .Z(n48632) );
  XOR U48473 ( .A(p_input[1600]), .B(n48638), .Z(n48361) );
  AND U48474 ( .A(n955), .B(n48639), .Z(n48638) );
  XOR U48475 ( .A(p_input[1632]), .B(p_input[1600]), .Z(n48639) );
  XOR U48476 ( .A(n48640), .B(n48641), .Z(n955) );
  AND U48477 ( .A(n48642), .B(n48643), .Z(n48641) );
  XNOR U48478 ( .A(p_input[1663]), .B(n48640), .Z(n48643) );
  XOR U48479 ( .A(n48640), .B(p_input[1631]), .Z(n48642) );
  XOR U48480 ( .A(n48644), .B(n48645), .Z(n48640) );
  AND U48481 ( .A(n48646), .B(n48647), .Z(n48645) );
  XNOR U48482 ( .A(p_input[1662]), .B(n48644), .Z(n48647) );
  XOR U48483 ( .A(n48644), .B(p_input[1630]), .Z(n48646) );
  XOR U48484 ( .A(n48648), .B(n48649), .Z(n48644) );
  AND U48485 ( .A(n48650), .B(n48651), .Z(n48649) );
  XNOR U48486 ( .A(p_input[1661]), .B(n48648), .Z(n48651) );
  XOR U48487 ( .A(n48648), .B(p_input[1629]), .Z(n48650) );
  XOR U48488 ( .A(n48652), .B(n48653), .Z(n48648) );
  AND U48489 ( .A(n48654), .B(n48655), .Z(n48653) );
  XNOR U48490 ( .A(p_input[1660]), .B(n48652), .Z(n48655) );
  XOR U48491 ( .A(n48652), .B(p_input[1628]), .Z(n48654) );
  XOR U48492 ( .A(n48656), .B(n48657), .Z(n48652) );
  AND U48493 ( .A(n48658), .B(n48659), .Z(n48657) );
  XNOR U48494 ( .A(p_input[1659]), .B(n48656), .Z(n48659) );
  XOR U48495 ( .A(n48656), .B(p_input[1627]), .Z(n48658) );
  XOR U48496 ( .A(n48660), .B(n48661), .Z(n48656) );
  AND U48497 ( .A(n48662), .B(n48663), .Z(n48661) );
  XNOR U48498 ( .A(p_input[1658]), .B(n48660), .Z(n48663) );
  XOR U48499 ( .A(n48660), .B(p_input[1626]), .Z(n48662) );
  XOR U48500 ( .A(n48664), .B(n48665), .Z(n48660) );
  AND U48501 ( .A(n48666), .B(n48667), .Z(n48665) );
  XNOR U48502 ( .A(p_input[1657]), .B(n48664), .Z(n48667) );
  XOR U48503 ( .A(n48664), .B(p_input[1625]), .Z(n48666) );
  XOR U48504 ( .A(n48668), .B(n48669), .Z(n48664) );
  AND U48505 ( .A(n48670), .B(n48671), .Z(n48669) );
  XNOR U48506 ( .A(p_input[1656]), .B(n48668), .Z(n48671) );
  XOR U48507 ( .A(n48668), .B(p_input[1624]), .Z(n48670) );
  XOR U48508 ( .A(n48672), .B(n48673), .Z(n48668) );
  AND U48509 ( .A(n48674), .B(n48675), .Z(n48673) );
  XNOR U48510 ( .A(p_input[1655]), .B(n48672), .Z(n48675) );
  XOR U48511 ( .A(n48672), .B(p_input[1623]), .Z(n48674) );
  XOR U48512 ( .A(n48676), .B(n48677), .Z(n48672) );
  AND U48513 ( .A(n48678), .B(n48679), .Z(n48677) );
  XNOR U48514 ( .A(p_input[1654]), .B(n48676), .Z(n48679) );
  XOR U48515 ( .A(n48676), .B(p_input[1622]), .Z(n48678) );
  XOR U48516 ( .A(n48680), .B(n48681), .Z(n48676) );
  AND U48517 ( .A(n48682), .B(n48683), .Z(n48681) );
  XNOR U48518 ( .A(p_input[1653]), .B(n48680), .Z(n48683) );
  XOR U48519 ( .A(n48680), .B(p_input[1621]), .Z(n48682) );
  XOR U48520 ( .A(n48684), .B(n48685), .Z(n48680) );
  AND U48521 ( .A(n48686), .B(n48687), .Z(n48685) );
  XNOR U48522 ( .A(p_input[1652]), .B(n48684), .Z(n48687) );
  XOR U48523 ( .A(n48684), .B(p_input[1620]), .Z(n48686) );
  XOR U48524 ( .A(n48688), .B(n48689), .Z(n48684) );
  AND U48525 ( .A(n48690), .B(n48691), .Z(n48689) );
  XNOR U48526 ( .A(p_input[1651]), .B(n48688), .Z(n48691) );
  XOR U48527 ( .A(n48688), .B(p_input[1619]), .Z(n48690) );
  XOR U48528 ( .A(n48692), .B(n48693), .Z(n48688) );
  AND U48529 ( .A(n48694), .B(n48695), .Z(n48693) );
  XNOR U48530 ( .A(p_input[1650]), .B(n48692), .Z(n48695) );
  XOR U48531 ( .A(n48692), .B(p_input[1618]), .Z(n48694) );
  XOR U48532 ( .A(n48696), .B(n48697), .Z(n48692) );
  AND U48533 ( .A(n48698), .B(n48699), .Z(n48697) );
  XNOR U48534 ( .A(p_input[1649]), .B(n48696), .Z(n48699) );
  XOR U48535 ( .A(n48696), .B(p_input[1617]), .Z(n48698) );
  XOR U48536 ( .A(n48700), .B(n48701), .Z(n48696) );
  AND U48537 ( .A(n48702), .B(n48703), .Z(n48701) );
  XNOR U48538 ( .A(p_input[1648]), .B(n48700), .Z(n48703) );
  XOR U48539 ( .A(n48700), .B(p_input[1616]), .Z(n48702) );
  XOR U48540 ( .A(n48704), .B(n48705), .Z(n48700) );
  AND U48541 ( .A(n48706), .B(n48707), .Z(n48705) );
  XNOR U48542 ( .A(p_input[1647]), .B(n48704), .Z(n48707) );
  XOR U48543 ( .A(n48704), .B(p_input[1615]), .Z(n48706) );
  XOR U48544 ( .A(n48708), .B(n48709), .Z(n48704) );
  AND U48545 ( .A(n48710), .B(n48711), .Z(n48709) );
  XNOR U48546 ( .A(p_input[1646]), .B(n48708), .Z(n48711) );
  XOR U48547 ( .A(n48708), .B(p_input[1614]), .Z(n48710) );
  XOR U48548 ( .A(n48712), .B(n48713), .Z(n48708) );
  AND U48549 ( .A(n48714), .B(n48715), .Z(n48713) );
  XNOR U48550 ( .A(p_input[1645]), .B(n48712), .Z(n48715) );
  XOR U48551 ( .A(n48712), .B(p_input[1613]), .Z(n48714) );
  XOR U48552 ( .A(n48716), .B(n48717), .Z(n48712) );
  AND U48553 ( .A(n48718), .B(n48719), .Z(n48717) );
  XNOR U48554 ( .A(p_input[1644]), .B(n48716), .Z(n48719) );
  XOR U48555 ( .A(n48716), .B(p_input[1612]), .Z(n48718) );
  XOR U48556 ( .A(n48720), .B(n48721), .Z(n48716) );
  AND U48557 ( .A(n48722), .B(n48723), .Z(n48721) );
  XNOR U48558 ( .A(p_input[1643]), .B(n48720), .Z(n48723) );
  XOR U48559 ( .A(n48720), .B(p_input[1611]), .Z(n48722) );
  XOR U48560 ( .A(n48724), .B(n48725), .Z(n48720) );
  AND U48561 ( .A(n48726), .B(n48727), .Z(n48725) );
  XNOR U48562 ( .A(p_input[1642]), .B(n48724), .Z(n48727) );
  XOR U48563 ( .A(n48724), .B(p_input[1610]), .Z(n48726) );
  XOR U48564 ( .A(n48728), .B(n48729), .Z(n48724) );
  AND U48565 ( .A(n48730), .B(n48731), .Z(n48729) );
  XNOR U48566 ( .A(p_input[1641]), .B(n48728), .Z(n48731) );
  XOR U48567 ( .A(n48728), .B(p_input[1609]), .Z(n48730) );
  XOR U48568 ( .A(n48732), .B(n48733), .Z(n48728) );
  AND U48569 ( .A(n48734), .B(n48735), .Z(n48733) );
  XNOR U48570 ( .A(p_input[1640]), .B(n48732), .Z(n48735) );
  XOR U48571 ( .A(n48732), .B(p_input[1608]), .Z(n48734) );
  XOR U48572 ( .A(n48736), .B(n48737), .Z(n48732) );
  AND U48573 ( .A(n48738), .B(n48739), .Z(n48737) );
  XNOR U48574 ( .A(p_input[1639]), .B(n48736), .Z(n48739) );
  XOR U48575 ( .A(n48736), .B(p_input[1607]), .Z(n48738) );
  XOR U48576 ( .A(n48740), .B(n48741), .Z(n48736) );
  AND U48577 ( .A(n48742), .B(n48743), .Z(n48741) );
  XNOR U48578 ( .A(p_input[1638]), .B(n48740), .Z(n48743) );
  XOR U48579 ( .A(n48740), .B(p_input[1606]), .Z(n48742) );
  XOR U48580 ( .A(n48744), .B(n48745), .Z(n48740) );
  AND U48581 ( .A(n48746), .B(n48747), .Z(n48745) );
  XNOR U48582 ( .A(p_input[1637]), .B(n48744), .Z(n48747) );
  XOR U48583 ( .A(n48744), .B(p_input[1605]), .Z(n48746) );
  XOR U48584 ( .A(n48748), .B(n48749), .Z(n48744) );
  AND U48585 ( .A(n48750), .B(n48751), .Z(n48749) );
  XNOR U48586 ( .A(p_input[1636]), .B(n48748), .Z(n48751) );
  XOR U48587 ( .A(n48748), .B(p_input[1604]), .Z(n48750) );
  XOR U48588 ( .A(n48752), .B(n48753), .Z(n48748) );
  AND U48589 ( .A(n48754), .B(n48755), .Z(n48753) );
  XNOR U48590 ( .A(p_input[1635]), .B(n48752), .Z(n48755) );
  XOR U48591 ( .A(n48752), .B(p_input[1603]), .Z(n48754) );
  XOR U48592 ( .A(n48756), .B(n48757), .Z(n48752) );
  AND U48593 ( .A(n48758), .B(n48759), .Z(n48757) );
  XNOR U48594 ( .A(p_input[1634]), .B(n48756), .Z(n48759) );
  XOR U48595 ( .A(n48756), .B(p_input[1602]), .Z(n48758) );
  XNOR U48596 ( .A(n48760), .B(n48761), .Z(n48756) );
  AND U48597 ( .A(n48762), .B(n48763), .Z(n48761) );
  XOR U48598 ( .A(p_input[1633]), .B(n48760), .Z(n48763) );
  XNOR U48599 ( .A(p_input[1601]), .B(n48760), .Z(n48762) );
  AND U48600 ( .A(p_input[1632]), .B(n48764), .Z(n48760) );
  IV U48601 ( .A(p_input[1600]), .Z(n48764) );
  XNOR U48602 ( .A(p_input[1536]), .B(n48765), .Z(n48358) );
  AND U48603 ( .A(n952), .B(n48766), .Z(n48765) );
  XOR U48604 ( .A(p_input[1568]), .B(p_input[1536]), .Z(n48766) );
  XOR U48605 ( .A(n48767), .B(n48768), .Z(n952) );
  AND U48606 ( .A(n48769), .B(n48770), .Z(n48768) );
  XNOR U48607 ( .A(p_input[1599]), .B(n48767), .Z(n48770) );
  XOR U48608 ( .A(n48767), .B(p_input[1567]), .Z(n48769) );
  XOR U48609 ( .A(n48771), .B(n48772), .Z(n48767) );
  AND U48610 ( .A(n48773), .B(n48774), .Z(n48772) );
  XNOR U48611 ( .A(p_input[1598]), .B(n48771), .Z(n48774) );
  XNOR U48612 ( .A(n48771), .B(n48373), .Z(n48773) );
  IV U48613 ( .A(p_input[1566]), .Z(n48373) );
  XOR U48614 ( .A(n48775), .B(n48776), .Z(n48771) );
  AND U48615 ( .A(n48777), .B(n48778), .Z(n48776) );
  XNOR U48616 ( .A(p_input[1597]), .B(n48775), .Z(n48778) );
  XNOR U48617 ( .A(n48775), .B(n48382), .Z(n48777) );
  IV U48618 ( .A(p_input[1565]), .Z(n48382) );
  XOR U48619 ( .A(n48779), .B(n48780), .Z(n48775) );
  AND U48620 ( .A(n48781), .B(n48782), .Z(n48780) );
  XNOR U48621 ( .A(p_input[1596]), .B(n48779), .Z(n48782) );
  XNOR U48622 ( .A(n48779), .B(n48391), .Z(n48781) );
  IV U48623 ( .A(p_input[1564]), .Z(n48391) );
  XOR U48624 ( .A(n48783), .B(n48784), .Z(n48779) );
  AND U48625 ( .A(n48785), .B(n48786), .Z(n48784) );
  XNOR U48626 ( .A(p_input[1595]), .B(n48783), .Z(n48786) );
  XNOR U48627 ( .A(n48783), .B(n48400), .Z(n48785) );
  IV U48628 ( .A(p_input[1563]), .Z(n48400) );
  XOR U48629 ( .A(n48787), .B(n48788), .Z(n48783) );
  AND U48630 ( .A(n48789), .B(n48790), .Z(n48788) );
  XNOR U48631 ( .A(p_input[1594]), .B(n48787), .Z(n48790) );
  XNOR U48632 ( .A(n48787), .B(n48409), .Z(n48789) );
  IV U48633 ( .A(p_input[1562]), .Z(n48409) );
  XOR U48634 ( .A(n48791), .B(n48792), .Z(n48787) );
  AND U48635 ( .A(n48793), .B(n48794), .Z(n48792) );
  XNOR U48636 ( .A(p_input[1593]), .B(n48791), .Z(n48794) );
  XNOR U48637 ( .A(n48791), .B(n48418), .Z(n48793) );
  IV U48638 ( .A(p_input[1561]), .Z(n48418) );
  XOR U48639 ( .A(n48795), .B(n48796), .Z(n48791) );
  AND U48640 ( .A(n48797), .B(n48798), .Z(n48796) );
  XNOR U48641 ( .A(p_input[1592]), .B(n48795), .Z(n48798) );
  XNOR U48642 ( .A(n48795), .B(n48427), .Z(n48797) );
  IV U48643 ( .A(p_input[1560]), .Z(n48427) );
  XOR U48644 ( .A(n48799), .B(n48800), .Z(n48795) );
  AND U48645 ( .A(n48801), .B(n48802), .Z(n48800) );
  XNOR U48646 ( .A(p_input[1591]), .B(n48799), .Z(n48802) );
  XNOR U48647 ( .A(n48799), .B(n48436), .Z(n48801) );
  IV U48648 ( .A(p_input[1559]), .Z(n48436) );
  XOR U48649 ( .A(n48803), .B(n48804), .Z(n48799) );
  AND U48650 ( .A(n48805), .B(n48806), .Z(n48804) );
  XNOR U48651 ( .A(p_input[1590]), .B(n48803), .Z(n48806) );
  XNOR U48652 ( .A(n48803), .B(n48445), .Z(n48805) );
  IV U48653 ( .A(p_input[1558]), .Z(n48445) );
  XOR U48654 ( .A(n48807), .B(n48808), .Z(n48803) );
  AND U48655 ( .A(n48809), .B(n48810), .Z(n48808) );
  XNOR U48656 ( .A(p_input[1589]), .B(n48807), .Z(n48810) );
  XNOR U48657 ( .A(n48807), .B(n48454), .Z(n48809) );
  IV U48658 ( .A(p_input[1557]), .Z(n48454) );
  XOR U48659 ( .A(n48811), .B(n48812), .Z(n48807) );
  AND U48660 ( .A(n48813), .B(n48814), .Z(n48812) );
  XNOR U48661 ( .A(p_input[1588]), .B(n48811), .Z(n48814) );
  XNOR U48662 ( .A(n48811), .B(n48463), .Z(n48813) );
  IV U48663 ( .A(p_input[1556]), .Z(n48463) );
  XOR U48664 ( .A(n48815), .B(n48816), .Z(n48811) );
  AND U48665 ( .A(n48817), .B(n48818), .Z(n48816) );
  XNOR U48666 ( .A(p_input[1587]), .B(n48815), .Z(n48818) );
  XNOR U48667 ( .A(n48815), .B(n48472), .Z(n48817) );
  IV U48668 ( .A(p_input[1555]), .Z(n48472) );
  XOR U48669 ( .A(n48819), .B(n48820), .Z(n48815) );
  AND U48670 ( .A(n48821), .B(n48822), .Z(n48820) );
  XNOR U48671 ( .A(p_input[1586]), .B(n48819), .Z(n48822) );
  XNOR U48672 ( .A(n48819), .B(n48481), .Z(n48821) );
  IV U48673 ( .A(p_input[1554]), .Z(n48481) );
  XOR U48674 ( .A(n48823), .B(n48824), .Z(n48819) );
  AND U48675 ( .A(n48825), .B(n48826), .Z(n48824) );
  XNOR U48676 ( .A(p_input[1585]), .B(n48823), .Z(n48826) );
  XNOR U48677 ( .A(n48823), .B(n48490), .Z(n48825) );
  IV U48678 ( .A(p_input[1553]), .Z(n48490) );
  XOR U48679 ( .A(n48827), .B(n48828), .Z(n48823) );
  AND U48680 ( .A(n48829), .B(n48830), .Z(n48828) );
  XNOR U48681 ( .A(p_input[1584]), .B(n48827), .Z(n48830) );
  XNOR U48682 ( .A(n48827), .B(n48499), .Z(n48829) );
  IV U48683 ( .A(p_input[1552]), .Z(n48499) );
  XOR U48684 ( .A(n48831), .B(n48832), .Z(n48827) );
  AND U48685 ( .A(n48833), .B(n48834), .Z(n48832) );
  XNOR U48686 ( .A(p_input[1583]), .B(n48831), .Z(n48834) );
  XNOR U48687 ( .A(n48831), .B(n48508), .Z(n48833) );
  IV U48688 ( .A(p_input[1551]), .Z(n48508) );
  XOR U48689 ( .A(n48835), .B(n48836), .Z(n48831) );
  AND U48690 ( .A(n48837), .B(n48838), .Z(n48836) );
  XNOR U48691 ( .A(p_input[1582]), .B(n48835), .Z(n48838) );
  XNOR U48692 ( .A(n48835), .B(n48517), .Z(n48837) );
  IV U48693 ( .A(p_input[1550]), .Z(n48517) );
  XOR U48694 ( .A(n48839), .B(n48840), .Z(n48835) );
  AND U48695 ( .A(n48841), .B(n48842), .Z(n48840) );
  XNOR U48696 ( .A(p_input[1581]), .B(n48839), .Z(n48842) );
  XNOR U48697 ( .A(n48839), .B(n48526), .Z(n48841) );
  IV U48698 ( .A(p_input[1549]), .Z(n48526) );
  XOR U48699 ( .A(n48843), .B(n48844), .Z(n48839) );
  AND U48700 ( .A(n48845), .B(n48846), .Z(n48844) );
  XNOR U48701 ( .A(p_input[1580]), .B(n48843), .Z(n48846) );
  XNOR U48702 ( .A(n48843), .B(n48535), .Z(n48845) );
  IV U48703 ( .A(p_input[1548]), .Z(n48535) );
  XOR U48704 ( .A(n48847), .B(n48848), .Z(n48843) );
  AND U48705 ( .A(n48849), .B(n48850), .Z(n48848) );
  XNOR U48706 ( .A(p_input[1579]), .B(n48847), .Z(n48850) );
  XNOR U48707 ( .A(n48847), .B(n48544), .Z(n48849) );
  IV U48708 ( .A(p_input[1547]), .Z(n48544) );
  XOR U48709 ( .A(n48851), .B(n48852), .Z(n48847) );
  AND U48710 ( .A(n48853), .B(n48854), .Z(n48852) );
  XNOR U48711 ( .A(p_input[1578]), .B(n48851), .Z(n48854) );
  XNOR U48712 ( .A(n48851), .B(n48553), .Z(n48853) );
  IV U48713 ( .A(p_input[1546]), .Z(n48553) );
  XOR U48714 ( .A(n48855), .B(n48856), .Z(n48851) );
  AND U48715 ( .A(n48857), .B(n48858), .Z(n48856) );
  XNOR U48716 ( .A(p_input[1577]), .B(n48855), .Z(n48858) );
  XNOR U48717 ( .A(n48855), .B(n48562), .Z(n48857) );
  IV U48718 ( .A(p_input[1545]), .Z(n48562) );
  XOR U48719 ( .A(n48859), .B(n48860), .Z(n48855) );
  AND U48720 ( .A(n48861), .B(n48862), .Z(n48860) );
  XNOR U48721 ( .A(p_input[1576]), .B(n48859), .Z(n48862) );
  XNOR U48722 ( .A(n48859), .B(n48571), .Z(n48861) );
  IV U48723 ( .A(p_input[1544]), .Z(n48571) );
  XOR U48724 ( .A(n48863), .B(n48864), .Z(n48859) );
  AND U48725 ( .A(n48865), .B(n48866), .Z(n48864) );
  XNOR U48726 ( .A(p_input[1575]), .B(n48863), .Z(n48866) );
  XNOR U48727 ( .A(n48863), .B(n48580), .Z(n48865) );
  IV U48728 ( .A(p_input[1543]), .Z(n48580) );
  XOR U48729 ( .A(n48867), .B(n48868), .Z(n48863) );
  AND U48730 ( .A(n48869), .B(n48870), .Z(n48868) );
  XNOR U48731 ( .A(p_input[1574]), .B(n48867), .Z(n48870) );
  XNOR U48732 ( .A(n48867), .B(n48589), .Z(n48869) );
  IV U48733 ( .A(p_input[1542]), .Z(n48589) );
  XOR U48734 ( .A(n48871), .B(n48872), .Z(n48867) );
  AND U48735 ( .A(n48873), .B(n48874), .Z(n48872) );
  XNOR U48736 ( .A(p_input[1573]), .B(n48871), .Z(n48874) );
  XNOR U48737 ( .A(n48871), .B(n48598), .Z(n48873) );
  IV U48738 ( .A(p_input[1541]), .Z(n48598) );
  XOR U48739 ( .A(n48875), .B(n48876), .Z(n48871) );
  AND U48740 ( .A(n48877), .B(n48878), .Z(n48876) );
  XNOR U48741 ( .A(p_input[1572]), .B(n48875), .Z(n48878) );
  XNOR U48742 ( .A(n48875), .B(n48607), .Z(n48877) );
  IV U48743 ( .A(p_input[1540]), .Z(n48607) );
  XOR U48744 ( .A(n48879), .B(n48880), .Z(n48875) );
  AND U48745 ( .A(n48881), .B(n48882), .Z(n48880) );
  XNOR U48746 ( .A(p_input[1571]), .B(n48879), .Z(n48882) );
  XNOR U48747 ( .A(n48879), .B(n48616), .Z(n48881) );
  IV U48748 ( .A(p_input[1539]), .Z(n48616) );
  XOR U48749 ( .A(n48883), .B(n48884), .Z(n48879) );
  AND U48750 ( .A(n48885), .B(n48886), .Z(n48884) );
  XNOR U48751 ( .A(p_input[1570]), .B(n48883), .Z(n48886) );
  XNOR U48752 ( .A(n48883), .B(n48625), .Z(n48885) );
  IV U48753 ( .A(p_input[1538]), .Z(n48625) );
  XNOR U48754 ( .A(n48887), .B(n48888), .Z(n48883) );
  AND U48755 ( .A(n48889), .B(n48890), .Z(n48888) );
  XOR U48756 ( .A(p_input[1569]), .B(n48887), .Z(n48890) );
  XNOR U48757 ( .A(p_input[1537]), .B(n48887), .Z(n48889) );
  AND U48758 ( .A(p_input[1568]), .B(n48891), .Z(n48887) );
  IV U48759 ( .A(p_input[1536]), .Z(n48891) );
  XOR U48760 ( .A(n48892), .B(n48893), .Z(n45248) );
  AND U48761 ( .A(n1037), .B(n48894), .Z(n48893) );
  XNOR U48762 ( .A(n48895), .B(n48892), .Z(n48894) );
  XOR U48763 ( .A(n48896), .B(n48897), .Z(n1037) );
  AND U48764 ( .A(n48898), .B(n48899), .Z(n48897) );
  XOR U48765 ( .A(n48896), .B(n45263), .Z(n48899) );
  XOR U48766 ( .A(n48900), .B(n48901), .Z(n45263) );
  AND U48767 ( .A(n907), .B(n48902), .Z(n48901) );
  XOR U48768 ( .A(n48903), .B(n48900), .Z(n48902) );
  XNOR U48769 ( .A(n45260), .B(n48896), .Z(n48898) );
  XOR U48770 ( .A(n48904), .B(n48905), .Z(n45260) );
  AND U48771 ( .A(n904), .B(n48906), .Z(n48905) );
  XOR U48772 ( .A(n48907), .B(n48904), .Z(n48906) );
  XOR U48773 ( .A(n48908), .B(n48909), .Z(n48896) );
  AND U48774 ( .A(n48910), .B(n48911), .Z(n48909) );
  XOR U48775 ( .A(n48908), .B(n45275), .Z(n48911) );
  XOR U48776 ( .A(n48912), .B(n48913), .Z(n45275) );
  AND U48777 ( .A(n907), .B(n48914), .Z(n48913) );
  XOR U48778 ( .A(n48915), .B(n48912), .Z(n48914) );
  XNOR U48779 ( .A(n45272), .B(n48908), .Z(n48910) );
  XOR U48780 ( .A(n48916), .B(n48917), .Z(n45272) );
  AND U48781 ( .A(n904), .B(n48918), .Z(n48917) );
  XOR U48782 ( .A(n48919), .B(n48916), .Z(n48918) );
  XOR U48783 ( .A(n48920), .B(n48921), .Z(n48908) );
  AND U48784 ( .A(n48922), .B(n48923), .Z(n48921) );
  XOR U48785 ( .A(n48920), .B(n45287), .Z(n48923) );
  XOR U48786 ( .A(n48924), .B(n48925), .Z(n45287) );
  AND U48787 ( .A(n907), .B(n48926), .Z(n48925) );
  XOR U48788 ( .A(n48927), .B(n48924), .Z(n48926) );
  XNOR U48789 ( .A(n45284), .B(n48920), .Z(n48922) );
  XOR U48790 ( .A(n48928), .B(n48929), .Z(n45284) );
  AND U48791 ( .A(n904), .B(n48930), .Z(n48929) );
  XOR U48792 ( .A(n48931), .B(n48928), .Z(n48930) );
  XOR U48793 ( .A(n48932), .B(n48933), .Z(n48920) );
  AND U48794 ( .A(n48934), .B(n48935), .Z(n48933) );
  XOR U48795 ( .A(n48932), .B(n45299), .Z(n48935) );
  XOR U48796 ( .A(n48936), .B(n48937), .Z(n45299) );
  AND U48797 ( .A(n907), .B(n48938), .Z(n48937) );
  XOR U48798 ( .A(n48939), .B(n48936), .Z(n48938) );
  XNOR U48799 ( .A(n45296), .B(n48932), .Z(n48934) );
  XOR U48800 ( .A(n48940), .B(n48941), .Z(n45296) );
  AND U48801 ( .A(n904), .B(n48942), .Z(n48941) );
  XOR U48802 ( .A(n48943), .B(n48940), .Z(n48942) );
  XOR U48803 ( .A(n48944), .B(n48945), .Z(n48932) );
  AND U48804 ( .A(n48946), .B(n48947), .Z(n48945) );
  XOR U48805 ( .A(n48944), .B(n45311), .Z(n48947) );
  XOR U48806 ( .A(n48948), .B(n48949), .Z(n45311) );
  AND U48807 ( .A(n907), .B(n48950), .Z(n48949) );
  XOR U48808 ( .A(n48951), .B(n48948), .Z(n48950) );
  XNOR U48809 ( .A(n45308), .B(n48944), .Z(n48946) );
  XOR U48810 ( .A(n48952), .B(n48953), .Z(n45308) );
  AND U48811 ( .A(n904), .B(n48954), .Z(n48953) );
  XOR U48812 ( .A(n48955), .B(n48952), .Z(n48954) );
  XOR U48813 ( .A(n48956), .B(n48957), .Z(n48944) );
  AND U48814 ( .A(n48958), .B(n48959), .Z(n48957) );
  XOR U48815 ( .A(n48956), .B(n45323), .Z(n48959) );
  XOR U48816 ( .A(n48960), .B(n48961), .Z(n45323) );
  AND U48817 ( .A(n907), .B(n48962), .Z(n48961) );
  XOR U48818 ( .A(n48963), .B(n48960), .Z(n48962) );
  XNOR U48819 ( .A(n45320), .B(n48956), .Z(n48958) );
  XOR U48820 ( .A(n48964), .B(n48965), .Z(n45320) );
  AND U48821 ( .A(n904), .B(n48966), .Z(n48965) );
  XOR U48822 ( .A(n48967), .B(n48964), .Z(n48966) );
  XOR U48823 ( .A(n48968), .B(n48969), .Z(n48956) );
  AND U48824 ( .A(n48970), .B(n48971), .Z(n48969) );
  XOR U48825 ( .A(n48968), .B(n45335), .Z(n48971) );
  XOR U48826 ( .A(n48972), .B(n48973), .Z(n45335) );
  AND U48827 ( .A(n907), .B(n48974), .Z(n48973) );
  XOR U48828 ( .A(n48975), .B(n48972), .Z(n48974) );
  XNOR U48829 ( .A(n45332), .B(n48968), .Z(n48970) );
  XOR U48830 ( .A(n48976), .B(n48977), .Z(n45332) );
  AND U48831 ( .A(n904), .B(n48978), .Z(n48977) );
  XOR U48832 ( .A(n48979), .B(n48976), .Z(n48978) );
  XOR U48833 ( .A(n48980), .B(n48981), .Z(n48968) );
  AND U48834 ( .A(n48982), .B(n48983), .Z(n48981) );
  XOR U48835 ( .A(n48980), .B(n45347), .Z(n48983) );
  XOR U48836 ( .A(n48984), .B(n48985), .Z(n45347) );
  AND U48837 ( .A(n907), .B(n48986), .Z(n48985) );
  XOR U48838 ( .A(n48987), .B(n48984), .Z(n48986) );
  XNOR U48839 ( .A(n45344), .B(n48980), .Z(n48982) );
  XOR U48840 ( .A(n48988), .B(n48989), .Z(n45344) );
  AND U48841 ( .A(n904), .B(n48990), .Z(n48989) );
  XOR U48842 ( .A(n48991), .B(n48988), .Z(n48990) );
  XOR U48843 ( .A(n48992), .B(n48993), .Z(n48980) );
  AND U48844 ( .A(n48994), .B(n48995), .Z(n48993) );
  XOR U48845 ( .A(n48992), .B(n45359), .Z(n48995) );
  XOR U48846 ( .A(n48996), .B(n48997), .Z(n45359) );
  AND U48847 ( .A(n907), .B(n48998), .Z(n48997) );
  XOR U48848 ( .A(n48999), .B(n48996), .Z(n48998) );
  XNOR U48849 ( .A(n45356), .B(n48992), .Z(n48994) );
  XOR U48850 ( .A(n49000), .B(n49001), .Z(n45356) );
  AND U48851 ( .A(n904), .B(n49002), .Z(n49001) );
  XOR U48852 ( .A(n49003), .B(n49000), .Z(n49002) );
  XOR U48853 ( .A(n49004), .B(n49005), .Z(n48992) );
  AND U48854 ( .A(n49006), .B(n49007), .Z(n49005) );
  XOR U48855 ( .A(n49004), .B(n45371), .Z(n49007) );
  XOR U48856 ( .A(n49008), .B(n49009), .Z(n45371) );
  AND U48857 ( .A(n907), .B(n49010), .Z(n49009) );
  XOR U48858 ( .A(n49011), .B(n49008), .Z(n49010) );
  XNOR U48859 ( .A(n45368), .B(n49004), .Z(n49006) );
  XOR U48860 ( .A(n49012), .B(n49013), .Z(n45368) );
  AND U48861 ( .A(n904), .B(n49014), .Z(n49013) );
  XOR U48862 ( .A(n49015), .B(n49012), .Z(n49014) );
  XOR U48863 ( .A(n49016), .B(n49017), .Z(n49004) );
  AND U48864 ( .A(n49018), .B(n49019), .Z(n49017) );
  XOR U48865 ( .A(n49016), .B(n45383), .Z(n49019) );
  XOR U48866 ( .A(n49020), .B(n49021), .Z(n45383) );
  AND U48867 ( .A(n907), .B(n49022), .Z(n49021) );
  XOR U48868 ( .A(n49023), .B(n49020), .Z(n49022) );
  XNOR U48869 ( .A(n45380), .B(n49016), .Z(n49018) );
  XOR U48870 ( .A(n49024), .B(n49025), .Z(n45380) );
  AND U48871 ( .A(n904), .B(n49026), .Z(n49025) );
  XOR U48872 ( .A(n49027), .B(n49024), .Z(n49026) );
  XOR U48873 ( .A(n49028), .B(n49029), .Z(n49016) );
  AND U48874 ( .A(n49030), .B(n49031), .Z(n49029) );
  XOR U48875 ( .A(n49028), .B(n45395), .Z(n49031) );
  XOR U48876 ( .A(n49032), .B(n49033), .Z(n45395) );
  AND U48877 ( .A(n907), .B(n49034), .Z(n49033) );
  XOR U48878 ( .A(n49035), .B(n49032), .Z(n49034) );
  XNOR U48879 ( .A(n45392), .B(n49028), .Z(n49030) );
  XOR U48880 ( .A(n49036), .B(n49037), .Z(n45392) );
  AND U48881 ( .A(n904), .B(n49038), .Z(n49037) );
  XOR U48882 ( .A(n49039), .B(n49036), .Z(n49038) );
  XOR U48883 ( .A(n49040), .B(n49041), .Z(n49028) );
  AND U48884 ( .A(n49042), .B(n49043), .Z(n49041) );
  XOR U48885 ( .A(n49040), .B(n45407), .Z(n49043) );
  XOR U48886 ( .A(n49044), .B(n49045), .Z(n45407) );
  AND U48887 ( .A(n907), .B(n49046), .Z(n49045) );
  XOR U48888 ( .A(n49047), .B(n49044), .Z(n49046) );
  XNOR U48889 ( .A(n45404), .B(n49040), .Z(n49042) );
  XOR U48890 ( .A(n49048), .B(n49049), .Z(n45404) );
  AND U48891 ( .A(n904), .B(n49050), .Z(n49049) );
  XOR U48892 ( .A(n49051), .B(n49048), .Z(n49050) );
  XOR U48893 ( .A(n49052), .B(n49053), .Z(n49040) );
  AND U48894 ( .A(n49054), .B(n49055), .Z(n49053) );
  XOR U48895 ( .A(n49052), .B(n45419), .Z(n49055) );
  XOR U48896 ( .A(n49056), .B(n49057), .Z(n45419) );
  AND U48897 ( .A(n907), .B(n49058), .Z(n49057) );
  XOR U48898 ( .A(n49059), .B(n49056), .Z(n49058) );
  XNOR U48899 ( .A(n45416), .B(n49052), .Z(n49054) );
  XOR U48900 ( .A(n49060), .B(n49061), .Z(n45416) );
  AND U48901 ( .A(n904), .B(n49062), .Z(n49061) );
  XOR U48902 ( .A(n49063), .B(n49060), .Z(n49062) );
  XOR U48903 ( .A(n49064), .B(n49065), .Z(n49052) );
  AND U48904 ( .A(n49066), .B(n49067), .Z(n49065) );
  XOR U48905 ( .A(n49064), .B(n45431), .Z(n49067) );
  XOR U48906 ( .A(n49068), .B(n49069), .Z(n45431) );
  AND U48907 ( .A(n907), .B(n49070), .Z(n49069) );
  XOR U48908 ( .A(n49071), .B(n49068), .Z(n49070) );
  XNOR U48909 ( .A(n45428), .B(n49064), .Z(n49066) );
  XOR U48910 ( .A(n49072), .B(n49073), .Z(n45428) );
  AND U48911 ( .A(n904), .B(n49074), .Z(n49073) );
  XOR U48912 ( .A(n49075), .B(n49072), .Z(n49074) );
  XOR U48913 ( .A(n49076), .B(n49077), .Z(n49064) );
  AND U48914 ( .A(n49078), .B(n49079), .Z(n49077) );
  XOR U48915 ( .A(n49076), .B(n45443), .Z(n49079) );
  XOR U48916 ( .A(n49080), .B(n49081), .Z(n45443) );
  AND U48917 ( .A(n907), .B(n49082), .Z(n49081) );
  XOR U48918 ( .A(n49083), .B(n49080), .Z(n49082) );
  XNOR U48919 ( .A(n45440), .B(n49076), .Z(n49078) );
  XOR U48920 ( .A(n49084), .B(n49085), .Z(n45440) );
  AND U48921 ( .A(n904), .B(n49086), .Z(n49085) );
  XOR U48922 ( .A(n49087), .B(n49084), .Z(n49086) );
  XOR U48923 ( .A(n49088), .B(n49089), .Z(n49076) );
  AND U48924 ( .A(n49090), .B(n49091), .Z(n49089) );
  XOR U48925 ( .A(n49088), .B(n45455), .Z(n49091) );
  XOR U48926 ( .A(n49092), .B(n49093), .Z(n45455) );
  AND U48927 ( .A(n907), .B(n49094), .Z(n49093) );
  XOR U48928 ( .A(n49095), .B(n49092), .Z(n49094) );
  XNOR U48929 ( .A(n45452), .B(n49088), .Z(n49090) );
  XOR U48930 ( .A(n49096), .B(n49097), .Z(n45452) );
  AND U48931 ( .A(n904), .B(n49098), .Z(n49097) );
  XOR U48932 ( .A(n49099), .B(n49096), .Z(n49098) );
  XOR U48933 ( .A(n49100), .B(n49101), .Z(n49088) );
  AND U48934 ( .A(n49102), .B(n49103), .Z(n49101) );
  XOR U48935 ( .A(n49100), .B(n45467), .Z(n49103) );
  XOR U48936 ( .A(n49104), .B(n49105), .Z(n45467) );
  AND U48937 ( .A(n907), .B(n49106), .Z(n49105) );
  XOR U48938 ( .A(n49107), .B(n49104), .Z(n49106) );
  XNOR U48939 ( .A(n45464), .B(n49100), .Z(n49102) );
  XOR U48940 ( .A(n49108), .B(n49109), .Z(n45464) );
  AND U48941 ( .A(n904), .B(n49110), .Z(n49109) );
  XOR U48942 ( .A(n49111), .B(n49108), .Z(n49110) );
  XOR U48943 ( .A(n49112), .B(n49113), .Z(n49100) );
  AND U48944 ( .A(n49114), .B(n49115), .Z(n49113) );
  XOR U48945 ( .A(n49112), .B(n45479), .Z(n49115) );
  XOR U48946 ( .A(n49116), .B(n49117), .Z(n45479) );
  AND U48947 ( .A(n907), .B(n49118), .Z(n49117) );
  XOR U48948 ( .A(n49119), .B(n49116), .Z(n49118) );
  XNOR U48949 ( .A(n45476), .B(n49112), .Z(n49114) );
  XOR U48950 ( .A(n49120), .B(n49121), .Z(n45476) );
  AND U48951 ( .A(n904), .B(n49122), .Z(n49121) );
  XOR U48952 ( .A(n49123), .B(n49120), .Z(n49122) );
  XOR U48953 ( .A(n49124), .B(n49125), .Z(n49112) );
  AND U48954 ( .A(n49126), .B(n49127), .Z(n49125) );
  XOR U48955 ( .A(n49124), .B(n45491), .Z(n49127) );
  XOR U48956 ( .A(n49128), .B(n49129), .Z(n45491) );
  AND U48957 ( .A(n907), .B(n49130), .Z(n49129) );
  XOR U48958 ( .A(n49131), .B(n49128), .Z(n49130) );
  XNOR U48959 ( .A(n45488), .B(n49124), .Z(n49126) );
  XOR U48960 ( .A(n49132), .B(n49133), .Z(n45488) );
  AND U48961 ( .A(n904), .B(n49134), .Z(n49133) );
  XOR U48962 ( .A(n49135), .B(n49132), .Z(n49134) );
  XOR U48963 ( .A(n49136), .B(n49137), .Z(n49124) );
  AND U48964 ( .A(n49138), .B(n49139), .Z(n49137) );
  XOR U48965 ( .A(n49136), .B(n45503), .Z(n49139) );
  XOR U48966 ( .A(n49140), .B(n49141), .Z(n45503) );
  AND U48967 ( .A(n907), .B(n49142), .Z(n49141) );
  XOR U48968 ( .A(n49143), .B(n49140), .Z(n49142) );
  XNOR U48969 ( .A(n45500), .B(n49136), .Z(n49138) );
  XOR U48970 ( .A(n49144), .B(n49145), .Z(n45500) );
  AND U48971 ( .A(n904), .B(n49146), .Z(n49145) );
  XOR U48972 ( .A(n49147), .B(n49144), .Z(n49146) );
  XOR U48973 ( .A(n49148), .B(n49149), .Z(n49136) );
  AND U48974 ( .A(n49150), .B(n49151), .Z(n49149) );
  XOR U48975 ( .A(n49148), .B(n45515), .Z(n49151) );
  XOR U48976 ( .A(n49152), .B(n49153), .Z(n45515) );
  AND U48977 ( .A(n907), .B(n49154), .Z(n49153) );
  XOR U48978 ( .A(n49155), .B(n49152), .Z(n49154) );
  XNOR U48979 ( .A(n45512), .B(n49148), .Z(n49150) );
  XOR U48980 ( .A(n49156), .B(n49157), .Z(n45512) );
  AND U48981 ( .A(n904), .B(n49158), .Z(n49157) );
  XOR U48982 ( .A(n49159), .B(n49156), .Z(n49158) );
  XOR U48983 ( .A(n49160), .B(n49161), .Z(n49148) );
  AND U48984 ( .A(n49162), .B(n49163), .Z(n49161) );
  XOR U48985 ( .A(n49160), .B(n45527), .Z(n49163) );
  XOR U48986 ( .A(n49164), .B(n49165), .Z(n45527) );
  AND U48987 ( .A(n907), .B(n49166), .Z(n49165) );
  XOR U48988 ( .A(n49167), .B(n49164), .Z(n49166) );
  XNOR U48989 ( .A(n45524), .B(n49160), .Z(n49162) );
  XOR U48990 ( .A(n49168), .B(n49169), .Z(n45524) );
  AND U48991 ( .A(n904), .B(n49170), .Z(n49169) );
  XOR U48992 ( .A(n49171), .B(n49168), .Z(n49170) );
  XOR U48993 ( .A(n49172), .B(n49173), .Z(n49160) );
  AND U48994 ( .A(n49174), .B(n49175), .Z(n49173) );
  XOR U48995 ( .A(n49172), .B(n45539), .Z(n49175) );
  XOR U48996 ( .A(n49176), .B(n49177), .Z(n45539) );
  AND U48997 ( .A(n907), .B(n49178), .Z(n49177) );
  XOR U48998 ( .A(n49179), .B(n49176), .Z(n49178) );
  XNOR U48999 ( .A(n45536), .B(n49172), .Z(n49174) );
  XOR U49000 ( .A(n49180), .B(n49181), .Z(n45536) );
  AND U49001 ( .A(n904), .B(n49182), .Z(n49181) );
  XOR U49002 ( .A(n49183), .B(n49180), .Z(n49182) );
  XOR U49003 ( .A(n49184), .B(n49185), .Z(n49172) );
  AND U49004 ( .A(n49186), .B(n49187), .Z(n49185) );
  XOR U49005 ( .A(n49184), .B(n45551), .Z(n49187) );
  XOR U49006 ( .A(n49188), .B(n49189), .Z(n45551) );
  AND U49007 ( .A(n907), .B(n49190), .Z(n49189) );
  XOR U49008 ( .A(n49191), .B(n49188), .Z(n49190) );
  XNOR U49009 ( .A(n45548), .B(n49184), .Z(n49186) );
  XOR U49010 ( .A(n49192), .B(n49193), .Z(n45548) );
  AND U49011 ( .A(n904), .B(n49194), .Z(n49193) );
  XOR U49012 ( .A(n49195), .B(n49192), .Z(n49194) );
  XOR U49013 ( .A(n49196), .B(n49197), .Z(n49184) );
  AND U49014 ( .A(n49198), .B(n49199), .Z(n49197) );
  XOR U49015 ( .A(n49196), .B(n45563), .Z(n49199) );
  XOR U49016 ( .A(n49200), .B(n49201), .Z(n45563) );
  AND U49017 ( .A(n907), .B(n49202), .Z(n49201) );
  XOR U49018 ( .A(n49203), .B(n49200), .Z(n49202) );
  XNOR U49019 ( .A(n45560), .B(n49196), .Z(n49198) );
  XOR U49020 ( .A(n49204), .B(n49205), .Z(n45560) );
  AND U49021 ( .A(n904), .B(n49206), .Z(n49205) );
  XOR U49022 ( .A(n49207), .B(n49204), .Z(n49206) );
  XOR U49023 ( .A(n49208), .B(n49209), .Z(n49196) );
  AND U49024 ( .A(n49210), .B(n49211), .Z(n49209) );
  XOR U49025 ( .A(n49208), .B(n45575), .Z(n49211) );
  XOR U49026 ( .A(n49212), .B(n49213), .Z(n45575) );
  AND U49027 ( .A(n907), .B(n49214), .Z(n49213) );
  XOR U49028 ( .A(n49215), .B(n49212), .Z(n49214) );
  XNOR U49029 ( .A(n45572), .B(n49208), .Z(n49210) );
  XOR U49030 ( .A(n49216), .B(n49217), .Z(n45572) );
  AND U49031 ( .A(n904), .B(n49218), .Z(n49217) );
  XOR U49032 ( .A(n49219), .B(n49216), .Z(n49218) );
  XOR U49033 ( .A(n49220), .B(n49221), .Z(n49208) );
  AND U49034 ( .A(n49222), .B(n49223), .Z(n49221) );
  XOR U49035 ( .A(n49220), .B(n45587), .Z(n49223) );
  XOR U49036 ( .A(n49224), .B(n49225), .Z(n45587) );
  AND U49037 ( .A(n907), .B(n49226), .Z(n49225) );
  XOR U49038 ( .A(n49227), .B(n49224), .Z(n49226) );
  XNOR U49039 ( .A(n45584), .B(n49220), .Z(n49222) );
  XOR U49040 ( .A(n49228), .B(n49229), .Z(n45584) );
  AND U49041 ( .A(n904), .B(n49230), .Z(n49229) );
  XOR U49042 ( .A(n49231), .B(n49228), .Z(n49230) );
  XOR U49043 ( .A(n49232), .B(n49233), .Z(n49220) );
  AND U49044 ( .A(n49234), .B(n49235), .Z(n49233) );
  XOR U49045 ( .A(n49232), .B(n45599), .Z(n49235) );
  XOR U49046 ( .A(n49236), .B(n49237), .Z(n45599) );
  AND U49047 ( .A(n907), .B(n49238), .Z(n49237) );
  XOR U49048 ( .A(n49239), .B(n49236), .Z(n49238) );
  XNOR U49049 ( .A(n45596), .B(n49232), .Z(n49234) );
  XOR U49050 ( .A(n49240), .B(n49241), .Z(n45596) );
  AND U49051 ( .A(n904), .B(n49242), .Z(n49241) );
  XOR U49052 ( .A(n49243), .B(n49240), .Z(n49242) );
  XOR U49053 ( .A(n49244), .B(n49245), .Z(n49232) );
  AND U49054 ( .A(n49246), .B(n49247), .Z(n49245) );
  XOR U49055 ( .A(n49244), .B(n45611), .Z(n49247) );
  XOR U49056 ( .A(n49248), .B(n49249), .Z(n45611) );
  AND U49057 ( .A(n907), .B(n49250), .Z(n49249) );
  XOR U49058 ( .A(n49251), .B(n49248), .Z(n49250) );
  XNOR U49059 ( .A(n45608), .B(n49244), .Z(n49246) );
  XOR U49060 ( .A(n49252), .B(n49253), .Z(n45608) );
  AND U49061 ( .A(n904), .B(n49254), .Z(n49253) );
  XOR U49062 ( .A(n49255), .B(n49252), .Z(n49254) );
  XOR U49063 ( .A(n49256), .B(n49257), .Z(n49244) );
  AND U49064 ( .A(n49258), .B(n49259), .Z(n49257) );
  XNOR U49065 ( .A(n49260), .B(n45624), .Z(n49259) );
  XOR U49066 ( .A(n49261), .B(n49262), .Z(n45624) );
  AND U49067 ( .A(n907), .B(n49263), .Z(n49262) );
  XOR U49068 ( .A(n49261), .B(n49264), .Z(n49263) );
  XNOR U49069 ( .A(n45621), .B(n49256), .Z(n49258) );
  XOR U49070 ( .A(n49265), .B(n49266), .Z(n45621) );
  AND U49071 ( .A(n904), .B(n49267), .Z(n49266) );
  XOR U49072 ( .A(n49265), .B(n49268), .Z(n49267) );
  IV U49073 ( .A(n49260), .Z(n49256) );
  AND U49074 ( .A(n48892), .B(n48895), .Z(n49260) );
  XNOR U49075 ( .A(n49269), .B(n49270), .Z(n48895) );
  AND U49076 ( .A(n907), .B(n49271), .Z(n49270) );
  XNOR U49077 ( .A(n49272), .B(n49269), .Z(n49271) );
  XOR U49078 ( .A(n49273), .B(n49274), .Z(n907) );
  AND U49079 ( .A(n49275), .B(n49276), .Z(n49274) );
  XOR U49080 ( .A(n49273), .B(n48903), .Z(n49276) );
  XNOR U49081 ( .A(n49277), .B(n49278), .Z(n48903) );
  AND U49082 ( .A(n49279), .B(n635), .Z(n49278) );
  AND U49083 ( .A(n49277), .B(n49280), .Z(n49279) );
  XNOR U49084 ( .A(n48900), .B(n49273), .Z(n49275) );
  XOR U49085 ( .A(n49281), .B(n49282), .Z(n48900) );
  AND U49086 ( .A(n49283), .B(n633), .Z(n49282) );
  NOR U49087 ( .A(n49281), .B(n49284), .Z(n49283) );
  XOR U49088 ( .A(n49285), .B(n49286), .Z(n49273) );
  AND U49089 ( .A(n49287), .B(n49288), .Z(n49286) );
  XOR U49090 ( .A(n49285), .B(n48915), .Z(n49288) );
  XOR U49091 ( .A(n49289), .B(n49290), .Z(n48915) );
  AND U49092 ( .A(n635), .B(n49291), .Z(n49290) );
  XOR U49093 ( .A(n49292), .B(n49289), .Z(n49291) );
  XNOR U49094 ( .A(n48912), .B(n49285), .Z(n49287) );
  XOR U49095 ( .A(n49293), .B(n49294), .Z(n48912) );
  AND U49096 ( .A(n633), .B(n49295), .Z(n49294) );
  XOR U49097 ( .A(n49296), .B(n49293), .Z(n49295) );
  XOR U49098 ( .A(n49297), .B(n49298), .Z(n49285) );
  AND U49099 ( .A(n49299), .B(n49300), .Z(n49298) );
  XOR U49100 ( .A(n49297), .B(n48927), .Z(n49300) );
  XOR U49101 ( .A(n49301), .B(n49302), .Z(n48927) );
  AND U49102 ( .A(n635), .B(n49303), .Z(n49302) );
  XOR U49103 ( .A(n49304), .B(n49301), .Z(n49303) );
  XNOR U49104 ( .A(n48924), .B(n49297), .Z(n49299) );
  XOR U49105 ( .A(n49305), .B(n49306), .Z(n48924) );
  AND U49106 ( .A(n633), .B(n49307), .Z(n49306) );
  XOR U49107 ( .A(n49308), .B(n49305), .Z(n49307) );
  XOR U49108 ( .A(n49309), .B(n49310), .Z(n49297) );
  AND U49109 ( .A(n49311), .B(n49312), .Z(n49310) );
  XOR U49110 ( .A(n49309), .B(n48939), .Z(n49312) );
  XOR U49111 ( .A(n49313), .B(n49314), .Z(n48939) );
  AND U49112 ( .A(n635), .B(n49315), .Z(n49314) );
  XOR U49113 ( .A(n49316), .B(n49313), .Z(n49315) );
  XNOR U49114 ( .A(n48936), .B(n49309), .Z(n49311) );
  XOR U49115 ( .A(n49317), .B(n49318), .Z(n48936) );
  AND U49116 ( .A(n633), .B(n49319), .Z(n49318) );
  XOR U49117 ( .A(n49320), .B(n49317), .Z(n49319) );
  XOR U49118 ( .A(n49321), .B(n49322), .Z(n49309) );
  AND U49119 ( .A(n49323), .B(n49324), .Z(n49322) );
  XOR U49120 ( .A(n49321), .B(n48951), .Z(n49324) );
  XOR U49121 ( .A(n49325), .B(n49326), .Z(n48951) );
  AND U49122 ( .A(n635), .B(n49327), .Z(n49326) );
  XOR U49123 ( .A(n49328), .B(n49325), .Z(n49327) );
  XNOR U49124 ( .A(n48948), .B(n49321), .Z(n49323) );
  XOR U49125 ( .A(n49329), .B(n49330), .Z(n48948) );
  AND U49126 ( .A(n633), .B(n49331), .Z(n49330) );
  XOR U49127 ( .A(n49332), .B(n49329), .Z(n49331) );
  XOR U49128 ( .A(n49333), .B(n49334), .Z(n49321) );
  AND U49129 ( .A(n49335), .B(n49336), .Z(n49334) );
  XOR U49130 ( .A(n49333), .B(n48963), .Z(n49336) );
  XOR U49131 ( .A(n49337), .B(n49338), .Z(n48963) );
  AND U49132 ( .A(n635), .B(n49339), .Z(n49338) );
  XOR U49133 ( .A(n49340), .B(n49337), .Z(n49339) );
  XNOR U49134 ( .A(n48960), .B(n49333), .Z(n49335) );
  XOR U49135 ( .A(n49341), .B(n49342), .Z(n48960) );
  AND U49136 ( .A(n633), .B(n49343), .Z(n49342) );
  XOR U49137 ( .A(n49344), .B(n49341), .Z(n49343) );
  XOR U49138 ( .A(n49345), .B(n49346), .Z(n49333) );
  AND U49139 ( .A(n49347), .B(n49348), .Z(n49346) );
  XOR U49140 ( .A(n49345), .B(n48975), .Z(n49348) );
  XOR U49141 ( .A(n49349), .B(n49350), .Z(n48975) );
  AND U49142 ( .A(n635), .B(n49351), .Z(n49350) );
  XOR U49143 ( .A(n49352), .B(n49349), .Z(n49351) );
  XNOR U49144 ( .A(n48972), .B(n49345), .Z(n49347) );
  XOR U49145 ( .A(n49353), .B(n49354), .Z(n48972) );
  AND U49146 ( .A(n633), .B(n49355), .Z(n49354) );
  XOR U49147 ( .A(n49356), .B(n49353), .Z(n49355) );
  XOR U49148 ( .A(n49357), .B(n49358), .Z(n49345) );
  AND U49149 ( .A(n49359), .B(n49360), .Z(n49358) );
  XOR U49150 ( .A(n49357), .B(n48987), .Z(n49360) );
  XOR U49151 ( .A(n49361), .B(n49362), .Z(n48987) );
  AND U49152 ( .A(n635), .B(n49363), .Z(n49362) );
  XOR U49153 ( .A(n49364), .B(n49361), .Z(n49363) );
  XNOR U49154 ( .A(n48984), .B(n49357), .Z(n49359) );
  XOR U49155 ( .A(n49365), .B(n49366), .Z(n48984) );
  AND U49156 ( .A(n633), .B(n49367), .Z(n49366) );
  XOR U49157 ( .A(n49368), .B(n49365), .Z(n49367) );
  XOR U49158 ( .A(n49369), .B(n49370), .Z(n49357) );
  AND U49159 ( .A(n49371), .B(n49372), .Z(n49370) );
  XOR U49160 ( .A(n49369), .B(n48999), .Z(n49372) );
  XOR U49161 ( .A(n49373), .B(n49374), .Z(n48999) );
  AND U49162 ( .A(n635), .B(n49375), .Z(n49374) );
  XOR U49163 ( .A(n49376), .B(n49373), .Z(n49375) );
  XNOR U49164 ( .A(n48996), .B(n49369), .Z(n49371) );
  XOR U49165 ( .A(n49377), .B(n49378), .Z(n48996) );
  AND U49166 ( .A(n633), .B(n49379), .Z(n49378) );
  XOR U49167 ( .A(n49380), .B(n49377), .Z(n49379) );
  XOR U49168 ( .A(n49381), .B(n49382), .Z(n49369) );
  AND U49169 ( .A(n49383), .B(n49384), .Z(n49382) );
  XOR U49170 ( .A(n49381), .B(n49011), .Z(n49384) );
  XOR U49171 ( .A(n49385), .B(n49386), .Z(n49011) );
  AND U49172 ( .A(n635), .B(n49387), .Z(n49386) );
  XOR U49173 ( .A(n49388), .B(n49385), .Z(n49387) );
  XNOR U49174 ( .A(n49008), .B(n49381), .Z(n49383) );
  XOR U49175 ( .A(n49389), .B(n49390), .Z(n49008) );
  AND U49176 ( .A(n633), .B(n49391), .Z(n49390) );
  XOR U49177 ( .A(n49392), .B(n49389), .Z(n49391) );
  XOR U49178 ( .A(n49393), .B(n49394), .Z(n49381) );
  AND U49179 ( .A(n49395), .B(n49396), .Z(n49394) );
  XOR U49180 ( .A(n49393), .B(n49023), .Z(n49396) );
  XOR U49181 ( .A(n49397), .B(n49398), .Z(n49023) );
  AND U49182 ( .A(n635), .B(n49399), .Z(n49398) );
  XOR U49183 ( .A(n49400), .B(n49397), .Z(n49399) );
  XNOR U49184 ( .A(n49020), .B(n49393), .Z(n49395) );
  XOR U49185 ( .A(n49401), .B(n49402), .Z(n49020) );
  AND U49186 ( .A(n633), .B(n49403), .Z(n49402) );
  XOR U49187 ( .A(n49404), .B(n49401), .Z(n49403) );
  XOR U49188 ( .A(n49405), .B(n49406), .Z(n49393) );
  AND U49189 ( .A(n49407), .B(n49408), .Z(n49406) );
  XOR U49190 ( .A(n49405), .B(n49035), .Z(n49408) );
  XOR U49191 ( .A(n49409), .B(n49410), .Z(n49035) );
  AND U49192 ( .A(n635), .B(n49411), .Z(n49410) );
  XOR U49193 ( .A(n49412), .B(n49409), .Z(n49411) );
  XNOR U49194 ( .A(n49032), .B(n49405), .Z(n49407) );
  XOR U49195 ( .A(n49413), .B(n49414), .Z(n49032) );
  AND U49196 ( .A(n633), .B(n49415), .Z(n49414) );
  XOR U49197 ( .A(n49416), .B(n49413), .Z(n49415) );
  XOR U49198 ( .A(n49417), .B(n49418), .Z(n49405) );
  AND U49199 ( .A(n49419), .B(n49420), .Z(n49418) );
  XOR U49200 ( .A(n49417), .B(n49047), .Z(n49420) );
  XOR U49201 ( .A(n49421), .B(n49422), .Z(n49047) );
  AND U49202 ( .A(n635), .B(n49423), .Z(n49422) );
  XOR U49203 ( .A(n49424), .B(n49421), .Z(n49423) );
  XNOR U49204 ( .A(n49044), .B(n49417), .Z(n49419) );
  XOR U49205 ( .A(n49425), .B(n49426), .Z(n49044) );
  AND U49206 ( .A(n633), .B(n49427), .Z(n49426) );
  XOR U49207 ( .A(n49428), .B(n49425), .Z(n49427) );
  XOR U49208 ( .A(n49429), .B(n49430), .Z(n49417) );
  AND U49209 ( .A(n49431), .B(n49432), .Z(n49430) );
  XOR U49210 ( .A(n49429), .B(n49059), .Z(n49432) );
  XOR U49211 ( .A(n49433), .B(n49434), .Z(n49059) );
  AND U49212 ( .A(n635), .B(n49435), .Z(n49434) );
  XOR U49213 ( .A(n49436), .B(n49433), .Z(n49435) );
  XNOR U49214 ( .A(n49056), .B(n49429), .Z(n49431) );
  XOR U49215 ( .A(n49437), .B(n49438), .Z(n49056) );
  AND U49216 ( .A(n633), .B(n49439), .Z(n49438) );
  XOR U49217 ( .A(n49440), .B(n49437), .Z(n49439) );
  XOR U49218 ( .A(n49441), .B(n49442), .Z(n49429) );
  AND U49219 ( .A(n49443), .B(n49444), .Z(n49442) );
  XOR U49220 ( .A(n49441), .B(n49071), .Z(n49444) );
  XOR U49221 ( .A(n49445), .B(n49446), .Z(n49071) );
  AND U49222 ( .A(n635), .B(n49447), .Z(n49446) );
  XOR U49223 ( .A(n49448), .B(n49445), .Z(n49447) );
  XNOR U49224 ( .A(n49068), .B(n49441), .Z(n49443) );
  XOR U49225 ( .A(n49449), .B(n49450), .Z(n49068) );
  AND U49226 ( .A(n633), .B(n49451), .Z(n49450) );
  XOR U49227 ( .A(n49452), .B(n49449), .Z(n49451) );
  XOR U49228 ( .A(n49453), .B(n49454), .Z(n49441) );
  AND U49229 ( .A(n49455), .B(n49456), .Z(n49454) );
  XOR U49230 ( .A(n49453), .B(n49083), .Z(n49456) );
  XOR U49231 ( .A(n49457), .B(n49458), .Z(n49083) );
  AND U49232 ( .A(n635), .B(n49459), .Z(n49458) );
  XOR U49233 ( .A(n49460), .B(n49457), .Z(n49459) );
  XNOR U49234 ( .A(n49080), .B(n49453), .Z(n49455) );
  XOR U49235 ( .A(n49461), .B(n49462), .Z(n49080) );
  AND U49236 ( .A(n633), .B(n49463), .Z(n49462) );
  XOR U49237 ( .A(n49464), .B(n49461), .Z(n49463) );
  XOR U49238 ( .A(n49465), .B(n49466), .Z(n49453) );
  AND U49239 ( .A(n49467), .B(n49468), .Z(n49466) );
  XOR U49240 ( .A(n49465), .B(n49095), .Z(n49468) );
  XOR U49241 ( .A(n49469), .B(n49470), .Z(n49095) );
  AND U49242 ( .A(n635), .B(n49471), .Z(n49470) );
  XOR U49243 ( .A(n49472), .B(n49469), .Z(n49471) );
  XNOR U49244 ( .A(n49092), .B(n49465), .Z(n49467) );
  XOR U49245 ( .A(n49473), .B(n49474), .Z(n49092) );
  AND U49246 ( .A(n633), .B(n49475), .Z(n49474) );
  XOR U49247 ( .A(n49476), .B(n49473), .Z(n49475) );
  XOR U49248 ( .A(n49477), .B(n49478), .Z(n49465) );
  AND U49249 ( .A(n49479), .B(n49480), .Z(n49478) );
  XOR U49250 ( .A(n49477), .B(n49107), .Z(n49480) );
  XOR U49251 ( .A(n49481), .B(n49482), .Z(n49107) );
  AND U49252 ( .A(n635), .B(n49483), .Z(n49482) );
  XOR U49253 ( .A(n49484), .B(n49481), .Z(n49483) );
  XNOR U49254 ( .A(n49104), .B(n49477), .Z(n49479) );
  XOR U49255 ( .A(n49485), .B(n49486), .Z(n49104) );
  AND U49256 ( .A(n633), .B(n49487), .Z(n49486) );
  XOR U49257 ( .A(n49488), .B(n49485), .Z(n49487) );
  XOR U49258 ( .A(n49489), .B(n49490), .Z(n49477) );
  AND U49259 ( .A(n49491), .B(n49492), .Z(n49490) );
  XOR U49260 ( .A(n49489), .B(n49119), .Z(n49492) );
  XOR U49261 ( .A(n49493), .B(n49494), .Z(n49119) );
  AND U49262 ( .A(n635), .B(n49495), .Z(n49494) );
  XOR U49263 ( .A(n49496), .B(n49493), .Z(n49495) );
  XNOR U49264 ( .A(n49116), .B(n49489), .Z(n49491) );
  XOR U49265 ( .A(n49497), .B(n49498), .Z(n49116) );
  AND U49266 ( .A(n633), .B(n49499), .Z(n49498) );
  XOR U49267 ( .A(n49500), .B(n49497), .Z(n49499) );
  XOR U49268 ( .A(n49501), .B(n49502), .Z(n49489) );
  AND U49269 ( .A(n49503), .B(n49504), .Z(n49502) );
  XOR U49270 ( .A(n49501), .B(n49131), .Z(n49504) );
  XOR U49271 ( .A(n49505), .B(n49506), .Z(n49131) );
  AND U49272 ( .A(n635), .B(n49507), .Z(n49506) );
  XOR U49273 ( .A(n49508), .B(n49505), .Z(n49507) );
  XNOR U49274 ( .A(n49128), .B(n49501), .Z(n49503) );
  XOR U49275 ( .A(n49509), .B(n49510), .Z(n49128) );
  AND U49276 ( .A(n633), .B(n49511), .Z(n49510) );
  XOR U49277 ( .A(n49512), .B(n49509), .Z(n49511) );
  XOR U49278 ( .A(n49513), .B(n49514), .Z(n49501) );
  AND U49279 ( .A(n49515), .B(n49516), .Z(n49514) );
  XOR U49280 ( .A(n49513), .B(n49143), .Z(n49516) );
  XOR U49281 ( .A(n49517), .B(n49518), .Z(n49143) );
  AND U49282 ( .A(n635), .B(n49519), .Z(n49518) );
  XOR U49283 ( .A(n49520), .B(n49517), .Z(n49519) );
  XNOR U49284 ( .A(n49140), .B(n49513), .Z(n49515) );
  XOR U49285 ( .A(n49521), .B(n49522), .Z(n49140) );
  AND U49286 ( .A(n633), .B(n49523), .Z(n49522) );
  XOR U49287 ( .A(n49524), .B(n49521), .Z(n49523) );
  XOR U49288 ( .A(n49525), .B(n49526), .Z(n49513) );
  AND U49289 ( .A(n49527), .B(n49528), .Z(n49526) );
  XOR U49290 ( .A(n49525), .B(n49155), .Z(n49528) );
  XOR U49291 ( .A(n49529), .B(n49530), .Z(n49155) );
  AND U49292 ( .A(n635), .B(n49531), .Z(n49530) );
  XOR U49293 ( .A(n49532), .B(n49529), .Z(n49531) );
  XNOR U49294 ( .A(n49152), .B(n49525), .Z(n49527) );
  XOR U49295 ( .A(n49533), .B(n49534), .Z(n49152) );
  AND U49296 ( .A(n633), .B(n49535), .Z(n49534) );
  XOR U49297 ( .A(n49536), .B(n49533), .Z(n49535) );
  XOR U49298 ( .A(n49537), .B(n49538), .Z(n49525) );
  AND U49299 ( .A(n49539), .B(n49540), .Z(n49538) );
  XOR U49300 ( .A(n49537), .B(n49167), .Z(n49540) );
  XOR U49301 ( .A(n49541), .B(n49542), .Z(n49167) );
  AND U49302 ( .A(n635), .B(n49543), .Z(n49542) );
  XOR U49303 ( .A(n49544), .B(n49541), .Z(n49543) );
  XNOR U49304 ( .A(n49164), .B(n49537), .Z(n49539) );
  XOR U49305 ( .A(n49545), .B(n49546), .Z(n49164) );
  AND U49306 ( .A(n633), .B(n49547), .Z(n49546) );
  XOR U49307 ( .A(n49548), .B(n49545), .Z(n49547) );
  XOR U49308 ( .A(n49549), .B(n49550), .Z(n49537) );
  AND U49309 ( .A(n49551), .B(n49552), .Z(n49550) );
  XOR U49310 ( .A(n49549), .B(n49179), .Z(n49552) );
  XOR U49311 ( .A(n49553), .B(n49554), .Z(n49179) );
  AND U49312 ( .A(n635), .B(n49555), .Z(n49554) );
  XOR U49313 ( .A(n49556), .B(n49553), .Z(n49555) );
  XNOR U49314 ( .A(n49176), .B(n49549), .Z(n49551) );
  XOR U49315 ( .A(n49557), .B(n49558), .Z(n49176) );
  AND U49316 ( .A(n633), .B(n49559), .Z(n49558) );
  XOR U49317 ( .A(n49560), .B(n49557), .Z(n49559) );
  XOR U49318 ( .A(n49561), .B(n49562), .Z(n49549) );
  AND U49319 ( .A(n49563), .B(n49564), .Z(n49562) );
  XOR U49320 ( .A(n49561), .B(n49191), .Z(n49564) );
  XOR U49321 ( .A(n49565), .B(n49566), .Z(n49191) );
  AND U49322 ( .A(n635), .B(n49567), .Z(n49566) );
  XOR U49323 ( .A(n49568), .B(n49565), .Z(n49567) );
  XNOR U49324 ( .A(n49188), .B(n49561), .Z(n49563) );
  XOR U49325 ( .A(n49569), .B(n49570), .Z(n49188) );
  AND U49326 ( .A(n633), .B(n49571), .Z(n49570) );
  XOR U49327 ( .A(n49572), .B(n49569), .Z(n49571) );
  XOR U49328 ( .A(n49573), .B(n49574), .Z(n49561) );
  AND U49329 ( .A(n49575), .B(n49576), .Z(n49574) );
  XOR U49330 ( .A(n49573), .B(n49203), .Z(n49576) );
  XOR U49331 ( .A(n49577), .B(n49578), .Z(n49203) );
  AND U49332 ( .A(n635), .B(n49579), .Z(n49578) );
  XOR U49333 ( .A(n49580), .B(n49577), .Z(n49579) );
  XNOR U49334 ( .A(n49200), .B(n49573), .Z(n49575) );
  XOR U49335 ( .A(n49581), .B(n49582), .Z(n49200) );
  AND U49336 ( .A(n633), .B(n49583), .Z(n49582) );
  XOR U49337 ( .A(n49584), .B(n49581), .Z(n49583) );
  XOR U49338 ( .A(n49585), .B(n49586), .Z(n49573) );
  AND U49339 ( .A(n49587), .B(n49588), .Z(n49586) );
  XOR U49340 ( .A(n49585), .B(n49215), .Z(n49588) );
  XOR U49341 ( .A(n49589), .B(n49590), .Z(n49215) );
  AND U49342 ( .A(n635), .B(n49591), .Z(n49590) );
  XOR U49343 ( .A(n49592), .B(n49589), .Z(n49591) );
  XNOR U49344 ( .A(n49212), .B(n49585), .Z(n49587) );
  XOR U49345 ( .A(n49593), .B(n49594), .Z(n49212) );
  AND U49346 ( .A(n633), .B(n49595), .Z(n49594) );
  XOR U49347 ( .A(n49596), .B(n49593), .Z(n49595) );
  XOR U49348 ( .A(n49597), .B(n49598), .Z(n49585) );
  AND U49349 ( .A(n49599), .B(n49600), .Z(n49598) );
  XOR U49350 ( .A(n49597), .B(n49227), .Z(n49600) );
  XOR U49351 ( .A(n49601), .B(n49602), .Z(n49227) );
  AND U49352 ( .A(n635), .B(n49603), .Z(n49602) );
  XOR U49353 ( .A(n49604), .B(n49601), .Z(n49603) );
  XNOR U49354 ( .A(n49224), .B(n49597), .Z(n49599) );
  XOR U49355 ( .A(n49605), .B(n49606), .Z(n49224) );
  AND U49356 ( .A(n633), .B(n49607), .Z(n49606) );
  XOR U49357 ( .A(n49608), .B(n49605), .Z(n49607) );
  XOR U49358 ( .A(n49609), .B(n49610), .Z(n49597) );
  AND U49359 ( .A(n49611), .B(n49612), .Z(n49610) );
  XOR U49360 ( .A(n49609), .B(n49239), .Z(n49612) );
  XOR U49361 ( .A(n49613), .B(n49614), .Z(n49239) );
  AND U49362 ( .A(n635), .B(n49615), .Z(n49614) );
  XOR U49363 ( .A(n49616), .B(n49613), .Z(n49615) );
  XNOR U49364 ( .A(n49236), .B(n49609), .Z(n49611) );
  XOR U49365 ( .A(n49617), .B(n49618), .Z(n49236) );
  AND U49366 ( .A(n633), .B(n49619), .Z(n49618) );
  XOR U49367 ( .A(n49620), .B(n49617), .Z(n49619) );
  XOR U49368 ( .A(n49621), .B(n49622), .Z(n49609) );
  AND U49369 ( .A(n49623), .B(n49624), .Z(n49622) );
  XOR U49370 ( .A(n49621), .B(n49251), .Z(n49624) );
  XOR U49371 ( .A(n49625), .B(n49626), .Z(n49251) );
  AND U49372 ( .A(n635), .B(n49627), .Z(n49626) );
  XOR U49373 ( .A(n49628), .B(n49625), .Z(n49627) );
  XNOR U49374 ( .A(n49248), .B(n49621), .Z(n49623) );
  XOR U49375 ( .A(n49629), .B(n49630), .Z(n49248) );
  AND U49376 ( .A(n633), .B(n49631), .Z(n49630) );
  XOR U49377 ( .A(n49632), .B(n49629), .Z(n49631) );
  XOR U49378 ( .A(n49633), .B(n49634), .Z(n49621) );
  AND U49379 ( .A(n49635), .B(n49636), .Z(n49634) );
  XNOR U49380 ( .A(n49637), .B(n49264), .Z(n49636) );
  XOR U49381 ( .A(n49638), .B(n49639), .Z(n49264) );
  AND U49382 ( .A(n635), .B(n49640), .Z(n49639) );
  XOR U49383 ( .A(n49638), .B(n49641), .Z(n49640) );
  XNOR U49384 ( .A(n49261), .B(n49633), .Z(n49635) );
  XOR U49385 ( .A(n49642), .B(n49643), .Z(n49261) );
  AND U49386 ( .A(n633), .B(n49644), .Z(n49643) );
  XOR U49387 ( .A(n49642), .B(n49645), .Z(n49644) );
  IV U49388 ( .A(n49637), .Z(n49633) );
  AND U49389 ( .A(n49269), .B(n49272), .Z(n49637) );
  XNOR U49390 ( .A(n49646), .B(n49647), .Z(n49272) );
  AND U49391 ( .A(n635), .B(n49648), .Z(n49647) );
  XNOR U49392 ( .A(n49649), .B(n49646), .Z(n49648) );
  XOR U49393 ( .A(n49650), .B(n49651), .Z(n635) );
  AND U49394 ( .A(n49652), .B(n49653), .Z(n49651) );
  XOR U49395 ( .A(n49280), .B(n49650), .Z(n49653) );
  IV U49396 ( .A(n49654), .Z(n49280) );
  AND U49397 ( .A(p_input[1535]), .B(p_input[1503]), .Z(n49654) );
  XOR U49398 ( .A(n49650), .B(n49277), .Z(n49652) );
  AND U49399 ( .A(p_input[1439]), .B(p_input[1471]), .Z(n49277) );
  XOR U49400 ( .A(n49655), .B(n49656), .Z(n49650) );
  AND U49401 ( .A(n49657), .B(n49658), .Z(n49656) );
  XOR U49402 ( .A(n49655), .B(n49292), .Z(n49658) );
  XNOR U49403 ( .A(p_input[1502]), .B(n49659), .Z(n49292) );
  AND U49404 ( .A(n967), .B(n49660), .Z(n49659) );
  XOR U49405 ( .A(p_input[1534]), .B(p_input[1502]), .Z(n49660) );
  XNOR U49406 ( .A(n49289), .B(n49655), .Z(n49657) );
  XOR U49407 ( .A(n49661), .B(n49662), .Z(n49289) );
  AND U49408 ( .A(n965), .B(n49663), .Z(n49662) );
  XOR U49409 ( .A(p_input[1470]), .B(p_input[1438]), .Z(n49663) );
  XOR U49410 ( .A(n49664), .B(n49665), .Z(n49655) );
  AND U49411 ( .A(n49666), .B(n49667), .Z(n49665) );
  XOR U49412 ( .A(n49664), .B(n49304), .Z(n49667) );
  XNOR U49413 ( .A(p_input[1501]), .B(n49668), .Z(n49304) );
  AND U49414 ( .A(n967), .B(n49669), .Z(n49668) );
  XOR U49415 ( .A(p_input[1533]), .B(p_input[1501]), .Z(n49669) );
  XNOR U49416 ( .A(n49301), .B(n49664), .Z(n49666) );
  XOR U49417 ( .A(n49670), .B(n49671), .Z(n49301) );
  AND U49418 ( .A(n965), .B(n49672), .Z(n49671) );
  XOR U49419 ( .A(p_input[1469]), .B(p_input[1437]), .Z(n49672) );
  XOR U49420 ( .A(n49673), .B(n49674), .Z(n49664) );
  AND U49421 ( .A(n49675), .B(n49676), .Z(n49674) );
  XOR U49422 ( .A(n49673), .B(n49316), .Z(n49676) );
  XNOR U49423 ( .A(p_input[1500]), .B(n49677), .Z(n49316) );
  AND U49424 ( .A(n967), .B(n49678), .Z(n49677) );
  XOR U49425 ( .A(p_input[1532]), .B(p_input[1500]), .Z(n49678) );
  XNOR U49426 ( .A(n49313), .B(n49673), .Z(n49675) );
  XOR U49427 ( .A(n49679), .B(n49680), .Z(n49313) );
  AND U49428 ( .A(n965), .B(n49681), .Z(n49680) );
  XOR U49429 ( .A(p_input[1468]), .B(p_input[1436]), .Z(n49681) );
  XOR U49430 ( .A(n49682), .B(n49683), .Z(n49673) );
  AND U49431 ( .A(n49684), .B(n49685), .Z(n49683) );
  XOR U49432 ( .A(n49682), .B(n49328), .Z(n49685) );
  XNOR U49433 ( .A(p_input[1499]), .B(n49686), .Z(n49328) );
  AND U49434 ( .A(n967), .B(n49687), .Z(n49686) );
  XOR U49435 ( .A(p_input[1531]), .B(p_input[1499]), .Z(n49687) );
  XNOR U49436 ( .A(n49325), .B(n49682), .Z(n49684) );
  XOR U49437 ( .A(n49688), .B(n49689), .Z(n49325) );
  AND U49438 ( .A(n965), .B(n49690), .Z(n49689) );
  XOR U49439 ( .A(p_input[1467]), .B(p_input[1435]), .Z(n49690) );
  XOR U49440 ( .A(n49691), .B(n49692), .Z(n49682) );
  AND U49441 ( .A(n49693), .B(n49694), .Z(n49692) );
  XOR U49442 ( .A(n49691), .B(n49340), .Z(n49694) );
  XNOR U49443 ( .A(p_input[1498]), .B(n49695), .Z(n49340) );
  AND U49444 ( .A(n967), .B(n49696), .Z(n49695) );
  XOR U49445 ( .A(p_input[1530]), .B(p_input[1498]), .Z(n49696) );
  XNOR U49446 ( .A(n49337), .B(n49691), .Z(n49693) );
  XOR U49447 ( .A(n49697), .B(n49698), .Z(n49337) );
  AND U49448 ( .A(n965), .B(n49699), .Z(n49698) );
  XOR U49449 ( .A(p_input[1466]), .B(p_input[1434]), .Z(n49699) );
  XOR U49450 ( .A(n49700), .B(n49701), .Z(n49691) );
  AND U49451 ( .A(n49702), .B(n49703), .Z(n49701) );
  XOR U49452 ( .A(n49700), .B(n49352), .Z(n49703) );
  XNOR U49453 ( .A(p_input[1497]), .B(n49704), .Z(n49352) );
  AND U49454 ( .A(n967), .B(n49705), .Z(n49704) );
  XOR U49455 ( .A(p_input[1529]), .B(p_input[1497]), .Z(n49705) );
  XNOR U49456 ( .A(n49349), .B(n49700), .Z(n49702) );
  XOR U49457 ( .A(n49706), .B(n49707), .Z(n49349) );
  AND U49458 ( .A(n965), .B(n49708), .Z(n49707) );
  XOR U49459 ( .A(p_input[1465]), .B(p_input[1433]), .Z(n49708) );
  XOR U49460 ( .A(n49709), .B(n49710), .Z(n49700) );
  AND U49461 ( .A(n49711), .B(n49712), .Z(n49710) );
  XOR U49462 ( .A(n49709), .B(n49364), .Z(n49712) );
  XNOR U49463 ( .A(p_input[1496]), .B(n49713), .Z(n49364) );
  AND U49464 ( .A(n967), .B(n49714), .Z(n49713) );
  XOR U49465 ( .A(p_input[1528]), .B(p_input[1496]), .Z(n49714) );
  XNOR U49466 ( .A(n49361), .B(n49709), .Z(n49711) );
  XOR U49467 ( .A(n49715), .B(n49716), .Z(n49361) );
  AND U49468 ( .A(n965), .B(n49717), .Z(n49716) );
  XOR U49469 ( .A(p_input[1464]), .B(p_input[1432]), .Z(n49717) );
  XOR U49470 ( .A(n49718), .B(n49719), .Z(n49709) );
  AND U49471 ( .A(n49720), .B(n49721), .Z(n49719) );
  XOR U49472 ( .A(n49718), .B(n49376), .Z(n49721) );
  XNOR U49473 ( .A(p_input[1495]), .B(n49722), .Z(n49376) );
  AND U49474 ( .A(n967), .B(n49723), .Z(n49722) );
  XOR U49475 ( .A(p_input[1527]), .B(p_input[1495]), .Z(n49723) );
  XNOR U49476 ( .A(n49373), .B(n49718), .Z(n49720) );
  XOR U49477 ( .A(n49724), .B(n49725), .Z(n49373) );
  AND U49478 ( .A(n965), .B(n49726), .Z(n49725) );
  XOR U49479 ( .A(p_input[1463]), .B(p_input[1431]), .Z(n49726) );
  XOR U49480 ( .A(n49727), .B(n49728), .Z(n49718) );
  AND U49481 ( .A(n49729), .B(n49730), .Z(n49728) );
  XOR U49482 ( .A(n49727), .B(n49388), .Z(n49730) );
  XNOR U49483 ( .A(p_input[1494]), .B(n49731), .Z(n49388) );
  AND U49484 ( .A(n967), .B(n49732), .Z(n49731) );
  XOR U49485 ( .A(p_input[1526]), .B(p_input[1494]), .Z(n49732) );
  XNOR U49486 ( .A(n49385), .B(n49727), .Z(n49729) );
  XOR U49487 ( .A(n49733), .B(n49734), .Z(n49385) );
  AND U49488 ( .A(n965), .B(n49735), .Z(n49734) );
  XOR U49489 ( .A(p_input[1462]), .B(p_input[1430]), .Z(n49735) );
  XOR U49490 ( .A(n49736), .B(n49737), .Z(n49727) );
  AND U49491 ( .A(n49738), .B(n49739), .Z(n49737) );
  XOR U49492 ( .A(n49736), .B(n49400), .Z(n49739) );
  XNOR U49493 ( .A(p_input[1493]), .B(n49740), .Z(n49400) );
  AND U49494 ( .A(n967), .B(n49741), .Z(n49740) );
  XOR U49495 ( .A(p_input[1525]), .B(p_input[1493]), .Z(n49741) );
  XNOR U49496 ( .A(n49397), .B(n49736), .Z(n49738) );
  XOR U49497 ( .A(n49742), .B(n49743), .Z(n49397) );
  AND U49498 ( .A(n965), .B(n49744), .Z(n49743) );
  XOR U49499 ( .A(p_input[1461]), .B(p_input[1429]), .Z(n49744) );
  XOR U49500 ( .A(n49745), .B(n49746), .Z(n49736) );
  AND U49501 ( .A(n49747), .B(n49748), .Z(n49746) );
  XOR U49502 ( .A(n49745), .B(n49412), .Z(n49748) );
  XNOR U49503 ( .A(p_input[1492]), .B(n49749), .Z(n49412) );
  AND U49504 ( .A(n967), .B(n49750), .Z(n49749) );
  XOR U49505 ( .A(p_input[1524]), .B(p_input[1492]), .Z(n49750) );
  XNOR U49506 ( .A(n49409), .B(n49745), .Z(n49747) );
  XOR U49507 ( .A(n49751), .B(n49752), .Z(n49409) );
  AND U49508 ( .A(n965), .B(n49753), .Z(n49752) );
  XOR U49509 ( .A(p_input[1460]), .B(p_input[1428]), .Z(n49753) );
  XOR U49510 ( .A(n49754), .B(n49755), .Z(n49745) );
  AND U49511 ( .A(n49756), .B(n49757), .Z(n49755) );
  XOR U49512 ( .A(n49754), .B(n49424), .Z(n49757) );
  XNOR U49513 ( .A(p_input[1491]), .B(n49758), .Z(n49424) );
  AND U49514 ( .A(n967), .B(n49759), .Z(n49758) );
  XOR U49515 ( .A(p_input[1523]), .B(p_input[1491]), .Z(n49759) );
  XNOR U49516 ( .A(n49421), .B(n49754), .Z(n49756) );
  XOR U49517 ( .A(n49760), .B(n49761), .Z(n49421) );
  AND U49518 ( .A(n965), .B(n49762), .Z(n49761) );
  XOR U49519 ( .A(p_input[1459]), .B(p_input[1427]), .Z(n49762) );
  XOR U49520 ( .A(n49763), .B(n49764), .Z(n49754) );
  AND U49521 ( .A(n49765), .B(n49766), .Z(n49764) );
  XOR U49522 ( .A(n49763), .B(n49436), .Z(n49766) );
  XNOR U49523 ( .A(p_input[1490]), .B(n49767), .Z(n49436) );
  AND U49524 ( .A(n967), .B(n49768), .Z(n49767) );
  XOR U49525 ( .A(p_input[1522]), .B(p_input[1490]), .Z(n49768) );
  XNOR U49526 ( .A(n49433), .B(n49763), .Z(n49765) );
  XOR U49527 ( .A(n49769), .B(n49770), .Z(n49433) );
  AND U49528 ( .A(n965), .B(n49771), .Z(n49770) );
  XOR U49529 ( .A(p_input[1458]), .B(p_input[1426]), .Z(n49771) );
  XOR U49530 ( .A(n49772), .B(n49773), .Z(n49763) );
  AND U49531 ( .A(n49774), .B(n49775), .Z(n49773) );
  XOR U49532 ( .A(n49772), .B(n49448), .Z(n49775) );
  XNOR U49533 ( .A(p_input[1489]), .B(n49776), .Z(n49448) );
  AND U49534 ( .A(n967), .B(n49777), .Z(n49776) );
  XOR U49535 ( .A(p_input[1521]), .B(p_input[1489]), .Z(n49777) );
  XNOR U49536 ( .A(n49445), .B(n49772), .Z(n49774) );
  XOR U49537 ( .A(n49778), .B(n49779), .Z(n49445) );
  AND U49538 ( .A(n965), .B(n49780), .Z(n49779) );
  XOR U49539 ( .A(p_input[1457]), .B(p_input[1425]), .Z(n49780) );
  XOR U49540 ( .A(n49781), .B(n49782), .Z(n49772) );
  AND U49541 ( .A(n49783), .B(n49784), .Z(n49782) );
  XOR U49542 ( .A(n49781), .B(n49460), .Z(n49784) );
  XNOR U49543 ( .A(p_input[1488]), .B(n49785), .Z(n49460) );
  AND U49544 ( .A(n967), .B(n49786), .Z(n49785) );
  XOR U49545 ( .A(p_input[1520]), .B(p_input[1488]), .Z(n49786) );
  XNOR U49546 ( .A(n49457), .B(n49781), .Z(n49783) );
  XOR U49547 ( .A(n49787), .B(n49788), .Z(n49457) );
  AND U49548 ( .A(n965), .B(n49789), .Z(n49788) );
  XOR U49549 ( .A(p_input[1456]), .B(p_input[1424]), .Z(n49789) );
  XOR U49550 ( .A(n49790), .B(n49791), .Z(n49781) );
  AND U49551 ( .A(n49792), .B(n49793), .Z(n49791) );
  XOR U49552 ( .A(n49790), .B(n49472), .Z(n49793) );
  XNOR U49553 ( .A(p_input[1487]), .B(n49794), .Z(n49472) );
  AND U49554 ( .A(n967), .B(n49795), .Z(n49794) );
  XOR U49555 ( .A(p_input[1519]), .B(p_input[1487]), .Z(n49795) );
  XNOR U49556 ( .A(n49469), .B(n49790), .Z(n49792) );
  XOR U49557 ( .A(n49796), .B(n49797), .Z(n49469) );
  AND U49558 ( .A(n965), .B(n49798), .Z(n49797) );
  XOR U49559 ( .A(p_input[1455]), .B(p_input[1423]), .Z(n49798) );
  XOR U49560 ( .A(n49799), .B(n49800), .Z(n49790) );
  AND U49561 ( .A(n49801), .B(n49802), .Z(n49800) );
  XOR U49562 ( .A(n49799), .B(n49484), .Z(n49802) );
  XNOR U49563 ( .A(p_input[1486]), .B(n49803), .Z(n49484) );
  AND U49564 ( .A(n967), .B(n49804), .Z(n49803) );
  XOR U49565 ( .A(p_input[1518]), .B(p_input[1486]), .Z(n49804) );
  XNOR U49566 ( .A(n49481), .B(n49799), .Z(n49801) );
  XOR U49567 ( .A(n49805), .B(n49806), .Z(n49481) );
  AND U49568 ( .A(n965), .B(n49807), .Z(n49806) );
  XOR U49569 ( .A(p_input[1454]), .B(p_input[1422]), .Z(n49807) );
  XOR U49570 ( .A(n49808), .B(n49809), .Z(n49799) );
  AND U49571 ( .A(n49810), .B(n49811), .Z(n49809) );
  XOR U49572 ( .A(n49808), .B(n49496), .Z(n49811) );
  XNOR U49573 ( .A(p_input[1485]), .B(n49812), .Z(n49496) );
  AND U49574 ( .A(n967), .B(n49813), .Z(n49812) );
  XOR U49575 ( .A(p_input[1517]), .B(p_input[1485]), .Z(n49813) );
  XNOR U49576 ( .A(n49493), .B(n49808), .Z(n49810) );
  XOR U49577 ( .A(n49814), .B(n49815), .Z(n49493) );
  AND U49578 ( .A(n965), .B(n49816), .Z(n49815) );
  XOR U49579 ( .A(p_input[1453]), .B(p_input[1421]), .Z(n49816) );
  XOR U49580 ( .A(n49817), .B(n49818), .Z(n49808) );
  AND U49581 ( .A(n49819), .B(n49820), .Z(n49818) );
  XOR U49582 ( .A(n49817), .B(n49508), .Z(n49820) );
  XNOR U49583 ( .A(p_input[1484]), .B(n49821), .Z(n49508) );
  AND U49584 ( .A(n967), .B(n49822), .Z(n49821) );
  XOR U49585 ( .A(p_input[1516]), .B(p_input[1484]), .Z(n49822) );
  XNOR U49586 ( .A(n49505), .B(n49817), .Z(n49819) );
  XOR U49587 ( .A(n49823), .B(n49824), .Z(n49505) );
  AND U49588 ( .A(n965), .B(n49825), .Z(n49824) );
  XOR U49589 ( .A(p_input[1452]), .B(p_input[1420]), .Z(n49825) );
  XOR U49590 ( .A(n49826), .B(n49827), .Z(n49817) );
  AND U49591 ( .A(n49828), .B(n49829), .Z(n49827) );
  XOR U49592 ( .A(n49826), .B(n49520), .Z(n49829) );
  XNOR U49593 ( .A(p_input[1483]), .B(n49830), .Z(n49520) );
  AND U49594 ( .A(n967), .B(n49831), .Z(n49830) );
  XOR U49595 ( .A(p_input[1515]), .B(p_input[1483]), .Z(n49831) );
  XNOR U49596 ( .A(n49517), .B(n49826), .Z(n49828) );
  XOR U49597 ( .A(n49832), .B(n49833), .Z(n49517) );
  AND U49598 ( .A(n965), .B(n49834), .Z(n49833) );
  XOR U49599 ( .A(p_input[1451]), .B(p_input[1419]), .Z(n49834) );
  XOR U49600 ( .A(n49835), .B(n49836), .Z(n49826) );
  AND U49601 ( .A(n49837), .B(n49838), .Z(n49836) );
  XOR U49602 ( .A(n49835), .B(n49532), .Z(n49838) );
  XNOR U49603 ( .A(p_input[1482]), .B(n49839), .Z(n49532) );
  AND U49604 ( .A(n967), .B(n49840), .Z(n49839) );
  XOR U49605 ( .A(p_input[1514]), .B(p_input[1482]), .Z(n49840) );
  XNOR U49606 ( .A(n49529), .B(n49835), .Z(n49837) );
  XOR U49607 ( .A(n49841), .B(n49842), .Z(n49529) );
  AND U49608 ( .A(n965), .B(n49843), .Z(n49842) );
  XOR U49609 ( .A(p_input[1450]), .B(p_input[1418]), .Z(n49843) );
  XOR U49610 ( .A(n49844), .B(n49845), .Z(n49835) );
  AND U49611 ( .A(n49846), .B(n49847), .Z(n49845) );
  XOR U49612 ( .A(n49844), .B(n49544), .Z(n49847) );
  XNOR U49613 ( .A(p_input[1481]), .B(n49848), .Z(n49544) );
  AND U49614 ( .A(n967), .B(n49849), .Z(n49848) );
  XOR U49615 ( .A(p_input[1513]), .B(p_input[1481]), .Z(n49849) );
  XNOR U49616 ( .A(n49541), .B(n49844), .Z(n49846) );
  XOR U49617 ( .A(n49850), .B(n49851), .Z(n49541) );
  AND U49618 ( .A(n965), .B(n49852), .Z(n49851) );
  XOR U49619 ( .A(p_input[1449]), .B(p_input[1417]), .Z(n49852) );
  XOR U49620 ( .A(n49853), .B(n49854), .Z(n49844) );
  AND U49621 ( .A(n49855), .B(n49856), .Z(n49854) );
  XOR U49622 ( .A(n49853), .B(n49556), .Z(n49856) );
  XNOR U49623 ( .A(p_input[1480]), .B(n49857), .Z(n49556) );
  AND U49624 ( .A(n967), .B(n49858), .Z(n49857) );
  XOR U49625 ( .A(p_input[1512]), .B(p_input[1480]), .Z(n49858) );
  XNOR U49626 ( .A(n49553), .B(n49853), .Z(n49855) );
  XOR U49627 ( .A(n49859), .B(n49860), .Z(n49553) );
  AND U49628 ( .A(n965), .B(n49861), .Z(n49860) );
  XOR U49629 ( .A(p_input[1448]), .B(p_input[1416]), .Z(n49861) );
  XOR U49630 ( .A(n49862), .B(n49863), .Z(n49853) );
  AND U49631 ( .A(n49864), .B(n49865), .Z(n49863) );
  XOR U49632 ( .A(n49862), .B(n49568), .Z(n49865) );
  XNOR U49633 ( .A(p_input[1479]), .B(n49866), .Z(n49568) );
  AND U49634 ( .A(n967), .B(n49867), .Z(n49866) );
  XOR U49635 ( .A(p_input[1511]), .B(p_input[1479]), .Z(n49867) );
  XNOR U49636 ( .A(n49565), .B(n49862), .Z(n49864) );
  XOR U49637 ( .A(n49868), .B(n49869), .Z(n49565) );
  AND U49638 ( .A(n965), .B(n49870), .Z(n49869) );
  XOR U49639 ( .A(p_input[1447]), .B(p_input[1415]), .Z(n49870) );
  XOR U49640 ( .A(n49871), .B(n49872), .Z(n49862) );
  AND U49641 ( .A(n49873), .B(n49874), .Z(n49872) );
  XOR U49642 ( .A(n49871), .B(n49580), .Z(n49874) );
  XNOR U49643 ( .A(p_input[1478]), .B(n49875), .Z(n49580) );
  AND U49644 ( .A(n967), .B(n49876), .Z(n49875) );
  XOR U49645 ( .A(p_input[1510]), .B(p_input[1478]), .Z(n49876) );
  XNOR U49646 ( .A(n49577), .B(n49871), .Z(n49873) );
  XOR U49647 ( .A(n49877), .B(n49878), .Z(n49577) );
  AND U49648 ( .A(n965), .B(n49879), .Z(n49878) );
  XOR U49649 ( .A(p_input[1446]), .B(p_input[1414]), .Z(n49879) );
  XOR U49650 ( .A(n49880), .B(n49881), .Z(n49871) );
  AND U49651 ( .A(n49882), .B(n49883), .Z(n49881) );
  XOR U49652 ( .A(n49880), .B(n49592), .Z(n49883) );
  XNOR U49653 ( .A(p_input[1477]), .B(n49884), .Z(n49592) );
  AND U49654 ( .A(n967), .B(n49885), .Z(n49884) );
  XOR U49655 ( .A(p_input[1509]), .B(p_input[1477]), .Z(n49885) );
  XNOR U49656 ( .A(n49589), .B(n49880), .Z(n49882) );
  XOR U49657 ( .A(n49886), .B(n49887), .Z(n49589) );
  AND U49658 ( .A(n965), .B(n49888), .Z(n49887) );
  XOR U49659 ( .A(p_input[1445]), .B(p_input[1413]), .Z(n49888) );
  XOR U49660 ( .A(n49889), .B(n49890), .Z(n49880) );
  AND U49661 ( .A(n49891), .B(n49892), .Z(n49890) );
  XOR U49662 ( .A(n49889), .B(n49604), .Z(n49892) );
  XNOR U49663 ( .A(p_input[1476]), .B(n49893), .Z(n49604) );
  AND U49664 ( .A(n967), .B(n49894), .Z(n49893) );
  XOR U49665 ( .A(p_input[1508]), .B(p_input[1476]), .Z(n49894) );
  XNOR U49666 ( .A(n49601), .B(n49889), .Z(n49891) );
  XOR U49667 ( .A(n49895), .B(n49896), .Z(n49601) );
  AND U49668 ( .A(n965), .B(n49897), .Z(n49896) );
  XOR U49669 ( .A(p_input[1444]), .B(p_input[1412]), .Z(n49897) );
  XOR U49670 ( .A(n49898), .B(n49899), .Z(n49889) );
  AND U49671 ( .A(n49900), .B(n49901), .Z(n49899) );
  XOR U49672 ( .A(n49898), .B(n49616), .Z(n49901) );
  XNOR U49673 ( .A(p_input[1475]), .B(n49902), .Z(n49616) );
  AND U49674 ( .A(n967), .B(n49903), .Z(n49902) );
  XOR U49675 ( .A(p_input[1507]), .B(p_input[1475]), .Z(n49903) );
  XNOR U49676 ( .A(n49613), .B(n49898), .Z(n49900) );
  XOR U49677 ( .A(n49904), .B(n49905), .Z(n49613) );
  AND U49678 ( .A(n965), .B(n49906), .Z(n49905) );
  XOR U49679 ( .A(p_input[1443]), .B(p_input[1411]), .Z(n49906) );
  XOR U49680 ( .A(n49907), .B(n49908), .Z(n49898) );
  AND U49681 ( .A(n49909), .B(n49910), .Z(n49908) );
  XOR U49682 ( .A(n49907), .B(n49628), .Z(n49910) );
  XNOR U49683 ( .A(p_input[1474]), .B(n49911), .Z(n49628) );
  AND U49684 ( .A(n967), .B(n49912), .Z(n49911) );
  XOR U49685 ( .A(p_input[1506]), .B(p_input[1474]), .Z(n49912) );
  XNOR U49686 ( .A(n49625), .B(n49907), .Z(n49909) );
  XOR U49687 ( .A(n49913), .B(n49914), .Z(n49625) );
  AND U49688 ( .A(n965), .B(n49915), .Z(n49914) );
  XOR U49689 ( .A(p_input[1442]), .B(p_input[1410]), .Z(n49915) );
  XOR U49690 ( .A(n49916), .B(n49917), .Z(n49907) );
  AND U49691 ( .A(n49918), .B(n49919), .Z(n49917) );
  XNOR U49692 ( .A(n49920), .B(n49641), .Z(n49919) );
  XNOR U49693 ( .A(p_input[1473]), .B(n49921), .Z(n49641) );
  AND U49694 ( .A(n967), .B(n49922), .Z(n49921) );
  XNOR U49695 ( .A(p_input[1505]), .B(n49923), .Z(n49922) );
  IV U49696 ( .A(p_input[1473]), .Z(n49923) );
  XNOR U49697 ( .A(n49638), .B(n49916), .Z(n49918) );
  XNOR U49698 ( .A(p_input[1409]), .B(n49924), .Z(n49638) );
  AND U49699 ( .A(n965), .B(n49925), .Z(n49924) );
  XOR U49700 ( .A(p_input[1441]), .B(p_input[1409]), .Z(n49925) );
  IV U49701 ( .A(n49920), .Z(n49916) );
  AND U49702 ( .A(n49646), .B(n49649), .Z(n49920) );
  XOR U49703 ( .A(p_input[1472]), .B(n49926), .Z(n49649) );
  AND U49704 ( .A(n967), .B(n49927), .Z(n49926) );
  XOR U49705 ( .A(p_input[1504]), .B(p_input[1472]), .Z(n49927) );
  XOR U49706 ( .A(n49928), .B(n49929), .Z(n967) );
  AND U49707 ( .A(n49930), .B(n49931), .Z(n49929) );
  XNOR U49708 ( .A(p_input[1535]), .B(n49928), .Z(n49931) );
  XOR U49709 ( .A(n49928), .B(p_input[1503]), .Z(n49930) );
  XOR U49710 ( .A(n49932), .B(n49933), .Z(n49928) );
  AND U49711 ( .A(n49934), .B(n49935), .Z(n49933) );
  XNOR U49712 ( .A(p_input[1534]), .B(n49932), .Z(n49935) );
  XOR U49713 ( .A(n49932), .B(p_input[1502]), .Z(n49934) );
  XOR U49714 ( .A(n49936), .B(n49937), .Z(n49932) );
  AND U49715 ( .A(n49938), .B(n49939), .Z(n49937) );
  XNOR U49716 ( .A(p_input[1533]), .B(n49936), .Z(n49939) );
  XOR U49717 ( .A(n49936), .B(p_input[1501]), .Z(n49938) );
  XOR U49718 ( .A(n49940), .B(n49941), .Z(n49936) );
  AND U49719 ( .A(n49942), .B(n49943), .Z(n49941) );
  XNOR U49720 ( .A(p_input[1532]), .B(n49940), .Z(n49943) );
  XOR U49721 ( .A(n49940), .B(p_input[1500]), .Z(n49942) );
  XOR U49722 ( .A(n49944), .B(n49945), .Z(n49940) );
  AND U49723 ( .A(n49946), .B(n49947), .Z(n49945) );
  XNOR U49724 ( .A(p_input[1531]), .B(n49944), .Z(n49947) );
  XOR U49725 ( .A(n49944), .B(p_input[1499]), .Z(n49946) );
  XOR U49726 ( .A(n49948), .B(n49949), .Z(n49944) );
  AND U49727 ( .A(n49950), .B(n49951), .Z(n49949) );
  XNOR U49728 ( .A(p_input[1530]), .B(n49948), .Z(n49951) );
  XOR U49729 ( .A(n49948), .B(p_input[1498]), .Z(n49950) );
  XOR U49730 ( .A(n49952), .B(n49953), .Z(n49948) );
  AND U49731 ( .A(n49954), .B(n49955), .Z(n49953) );
  XNOR U49732 ( .A(p_input[1529]), .B(n49952), .Z(n49955) );
  XOR U49733 ( .A(n49952), .B(p_input[1497]), .Z(n49954) );
  XOR U49734 ( .A(n49956), .B(n49957), .Z(n49952) );
  AND U49735 ( .A(n49958), .B(n49959), .Z(n49957) );
  XNOR U49736 ( .A(p_input[1528]), .B(n49956), .Z(n49959) );
  XOR U49737 ( .A(n49956), .B(p_input[1496]), .Z(n49958) );
  XOR U49738 ( .A(n49960), .B(n49961), .Z(n49956) );
  AND U49739 ( .A(n49962), .B(n49963), .Z(n49961) );
  XNOR U49740 ( .A(p_input[1527]), .B(n49960), .Z(n49963) );
  XOR U49741 ( .A(n49960), .B(p_input[1495]), .Z(n49962) );
  XOR U49742 ( .A(n49964), .B(n49965), .Z(n49960) );
  AND U49743 ( .A(n49966), .B(n49967), .Z(n49965) );
  XNOR U49744 ( .A(p_input[1526]), .B(n49964), .Z(n49967) );
  XOR U49745 ( .A(n49964), .B(p_input[1494]), .Z(n49966) );
  XOR U49746 ( .A(n49968), .B(n49969), .Z(n49964) );
  AND U49747 ( .A(n49970), .B(n49971), .Z(n49969) );
  XNOR U49748 ( .A(p_input[1525]), .B(n49968), .Z(n49971) );
  XOR U49749 ( .A(n49968), .B(p_input[1493]), .Z(n49970) );
  XOR U49750 ( .A(n49972), .B(n49973), .Z(n49968) );
  AND U49751 ( .A(n49974), .B(n49975), .Z(n49973) );
  XNOR U49752 ( .A(p_input[1524]), .B(n49972), .Z(n49975) );
  XOR U49753 ( .A(n49972), .B(p_input[1492]), .Z(n49974) );
  XOR U49754 ( .A(n49976), .B(n49977), .Z(n49972) );
  AND U49755 ( .A(n49978), .B(n49979), .Z(n49977) );
  XNOR U49756 ( .A(p_input[1523]), .B(n49976), .Z(n49979) );
  XOR U49757 ( .A(n49976), .B(p_input[1491]), .Z(n49978) );
  XOR U49758 ( .A(n49980), .B(n49981), .Z(n49976) );
  AND U49759 ( .A(n49982), .B(n49983), .Z(n49981) );
  XNOR U49760 ( .A(p_input[1522]), .B(n49980), .Z(n49983) );
  XOR U49761 ( .A(n49980), .B(p_input[1490]), .Z(n49982) );
  XOR U49762 ( .A(n49984), .B(n49985), .Z(n49980) );
  AND U49763 ( .A(n49986), .B(n49987), .Z(n49985) );
  XNOR U49764 ( .A(p_input[1521]), .B(n49984), .Z(n49987) );
  XOR U49765 ( .A(n49984), .B(p_input[1489]), .Z(n49986) );
  XOR U49766 ( .A(n49988), .B(n49989), .Z(n49984) );
  AND U49767 ( .A(n49990), .B(n49991), .Z(n49989) );
  XNOR U49768 ( .A(p_input[1520]), .B(n49988), .Z(n49991) );
  XOR U49769 ( .A(n49988), .B(p_input[1488]), .Z(n49990) );
  XOR U49770 ( .A(n49992), .B(n49993), .Z(n49988) );
  AND U49771 ( .A(n49994), .B(n49995), .Z(n49993) );
  XNOR U49772 ( .A(p_input[1519]), .B(n49992), .Z(n49995) );
  XOR U49773 ( .A(n49992), .B(p_input[1487]), .Z(n49994) );
  XOR U49774 ( .A(n49996), .B(n49997), .Z(n49992) );
  AND U49775 ( .A(n49998), .B(n49999), .Z(n49997) );
  XNOR U49776 ( .A(p_input[1518]), .B(n49996), .Z(n49999) );
  XOR U49777 ( .A(n49996), .B(p_input[1486]), .Z(n49998) );
  XOR U49778 ( .A(n50000), .B(n50001), .Z(n49996) );
  AND U49779 ( .A(n50002), .B(n50003), .Z(n50001) );
  XNOR U49780 ( .A(p_input[1517]), .B(n50000), .Z(n50003) );
  XOR U49781 ( .A(n50000), .B(p_input[1485]), .Z(n50002) );
  XOR U49782 ( .A(n50004), .B(n50005), .Z(n50000) );
  AND U49783 ( .A(n50006), .B(n50007), .Z(n50005) );
  XNOR U49784 ( .A(p_input[1516]), .B(n50004), .Z(n50007) );
  XOR U49785 ( .A(n50004), .B(p_input[1484]), .Z(n50006) );
  XOR U49786 ( .A(n50008), .B(n50009), .Z(n50004) );
  AND U49787 ( .A(n50010), .B(n50011), .Z(n50009) );
  XNOR U49788 ( .A(p_input[1515]), .B(n50008), .Z(n50011) );
  XOR U49789 ( .A(n50008), .B(p_input[1483]), .Z(n50010) );
  XOR U49790 ( .A(n50012), .B(n50013), .Z(n50008) );
  AND U49791 ( .A(n50014), .B(n50015), .Z(n50013) );
  XNOR U49792 ( .A(p_input[1514]), .B(n50012), .Z(n50015) );
  XOR U49793 ( .A(n50012), .B(p_input[1482]), .Z(n50014) );
  XOR U49794 ( .A(n50016), .B(n50017), .Z(n50012) );
  AND U49795 ( .A(n50018), .B(n50019), .Z(n50017) );
  XNOR U49796 ( .A(p_input[1513]), .B(n50016), .Z(n50019) );
  XOR U49797 ( .A(n50016), .B(p_input[1481]), .Z(n50018) );
  XOR U49798 ( .A(n50020), .B(n50021), .Z(n50016) );
  AND U49799 ( .A(n50022), .B(n50023), .Z(n50021) );
  XNOR U49800 ( .A(p_input[1512]), .B(n50020), .Z(n50023) );
  XOR U49801 ( .A(n50020), .B(p_input[1480]), .Z(n50022) );
  XOR U49802 ( .A(n50024), .B(n50025), .Z(n50020) );
  AND U49803 ( .A(n50026), .B(n50027), .Z(n50025) );
  XNOR U49804 ( .A(p_input[1511]), .B(n50024), .Z(n50027) );
  XOR U49805 ( .A(n50024), .B(p_input[1479]), .Z(n50026) );
  XOR U49806 ( .A(n50028), .B(n50029), .Z(n50024) );
  AND U49807 ( .A(n50030), .B(n50031), .Z(n50029) );
  XNOR U49808 ( .A(p_input[1510]), .B(n50028), .Z(n50031) );
  XOR U49809 ( .A(n50028), .B(p_input[1478]), .Z(n50030) );
  XOR U49810 ( .A(n50032), .B(n50033), .Z(n50028) );
  AND U49811 ( .A(n50034), .B(n50035), .Z(n50033) );
  XNOR U49812 ( .A(p_input[1509]), .B(n50032), .Z(n50035) );
  XOR U49813 ( .A(n50032), .B(p_input[1477]), .Z(n50034) );
  XOR U49814 ( .A(n50036), .B(n50037), .Z(n50032) );
  AND U49815 ( .A(n50038), .B(n50039), .Z(n50037) );
  XNOR U49816 ( .A(p_input[1508]), .B(n50036), .Z(n50039) );
  XOR U49817 ( .A(n50036), .B(p_input[1476]), .Z(n50038) );
  XOR U49818 ( .A(n50040), .B(n50041), .Z(n50036) );
  AND U49819 ( .A(n50042), .B(n50043), .Z(n50041) );
  XNOR U49820 ( .A(p_input[1507]), .B(n50040), .Z(n50043) );
  XOR U49821 ( .A(n50040), .B(p_input[1475]), .Z(n50042) );
  XOR U49822 ( .A(n50044), .B(n50045), .Z(n50040) );
  AND U49823 ( .A(n50046), .B(n50047), .Z(n50045) );
  XNOR U49824 ( .A(p_input[1506]), .B(n50044), .Z(n50047) );
  XOR U49825 ( .A(n50044), .B(p_input[1474]), .Z(n50046) );
  XNOR U49826 ( .A(n50048), .B(n50049), .Z(n50044) );
  AND U49827 ( .A(n50050), .B(n50051), .Z(n50049) );
  XOR U49828 ( .A(p_input[1505]), .B(n50048), .Z(n50051) );
  XNOR U49829 ( .A(p_input[1473]), .B(n50048), .Z(n50050) );
  AND U49830 ( .A(p_input[1504]), .B(n50052), .Z(n50048) );
  IV U49831 ( .A(p_input[1472]), .Z(n50052) );
  XNOR U49832 ( .A(p_input[1408]), .B(n50053), .Z(n49646) );
  AND U49833 ( .A(n965), .B(n50054), .Z(n50053) );
  XOR U49834 ( .A(p_input[1440]), .B(p_input[1408]), .Z(n50054) );
  XOR U49835 ( .A(n50055), .B(n50056), .Z(n965) );
  AND U49836 ( .A(n50057), .B(n50058), .Z(n50056) );
  XNOR U49837 ( .A(p_input[1471]), .B(n50055), .Z(n50058) );
  XOR U49838 ( .A(n50055), .B(p_input[1439]), .Z(n50057) );
  XOR U49839 ( .A(n50059), .B(n50060), .Z(n50055) );
  AND U49840 ( .A(n50061), .B(n50062), .Z(n50060) );
  XNOR U49841 ( .A(p_input[1470]), .B(n50059), .Z(n50062) );
  XNOR U49842 ( .A(n50059), .B(n49661), .Z(n50061) );
  IV U49843 ( .A(p_input[1438]), .Z(n49661) );
  XOR U49844 ( .A(n50063), .B(n50064), .Z(n50059) );
  AND U49845 ( .A(n50065), .B(n50066), .Z(n50064) );
  XNOR U49846 ( .A(p_input[1469]), .B(n50063), .Z(n50066) );
  XNOR U49847 ( .A(n50063), .B(n49670), .Z(n50065) );
  IV U49848 ( .A(p_input[1437]), .Z(n49670) );
  XOR U49849 ( .A(n50067), .B(n50068), .Z(n50063) );
  AND U49850 ( .A(n50069), .B(n50070), .Z(n50068) );
  XNOR U49851 ( .A(p_input[1468]), .B(n50067), .Z(n50070) );
  XNOR U49852 ( .A(n50067), .B(n49679), .Z(n50069) );
  IV U49853 ( .A(p_input[1436]), .Z(n49679) );
  XOR U49854 ( .A(n50071), .B(n50072), .Z(n50067) );
  AND U49855 ( .A(n50073), .B(n50074), .Z(n50072) );
  XNOR U49856 ( .A(p_input[1467]), .B(n50071), .Z(n50074) );
  XNOR U49857 ( .A(n50071), .B(n49688), .Z(n50073) );
  IV U49858 ( .A(p_input[1435]), .Z(n49688) );
  XOR U49859 ( .A(n50075), .B(n50076), .Z(n50071) );
  AND U49860 ( .A(n50077), .B(n50078), .Z(n50076) );
  XNOR U49861 ( .A(p_input[1466]), .B(n50075), .Z(n50078) );
  XNOR U49862 ( .A(n50075), .B(n49697), .Z(n50077) );
  IV U49863 ( .A(p_input[1434]), .Z(n49697) );
  XOR U49864 ( .A(n50079), .B(n50080), .Z(n50075) );
  AND U49865 ( .A(n50081), .B(n50082), .Z(n50080) );
  XNOR U49866 ( .A(p_input[1465]), .B(n50079), .Z(n50082) );
  XNOR U49867 ( .A(n50079), .B(n49706), .Z(n50081) );
  IV U49868 ( .A(p_input[1433]), .Z(n49706) );
  XOR U49869 ( .A(n50083), .B(n50084), .Z(n50079) );
  AND U49870 ( .A(n50085), .B(n50086), .Z(n50084) );
  XNOR U49871 ( .A(p_input[1464]), .B(n50083), .Z(n50086) );
  XNOR U49872 ( .A(n50083), .B(n49715), .Z(n50085) );
  IV U49873 ( .A(p_input[1432]), .Z(n49715) );
  XOR U49874 ( .A(n50087), .B(n50088), .Z(n50083) );
  AND U49875 ( .A(n50089), .B(n50090), .Z(n50088) );
  XNOR U49876 ( .A(p_input[1463]), .B(n50087), .Z(n50090) );
  XNOR U49877 ( .A(n50087), .B(n49724), .Z(n50089) );
  IV U49878 ( .A(p_input[1431]), .Z(n49724) );
  XOR U49879 ( .A(n50091), .B(n50092), .Z(n50087) );
  AND U49880 ( .A(n50093), .B(n50094), .Z(n50092) );
  XNOR U49881 ( .A(p_input[1462]), .B(n50091), .Z(n50094) );
  XNOR U49882 ( .A(n50091), .B(n49733), .Z(n50093) );
  IV U49883 ( .A(p_input[1430]), .Z(n49733) );
  XOR U49884 ( .A(n50095), .B(n50096), .Z(n50091) );
  AND U49885 ( .A(n50097), .B(n50098), .Z(n50096) );
  XNOR U49886 ( .A(p_input[1461]), .B(n50095), .Z(n50098) );
  XNOR U49887 ( .A(n50095), .B(n49742), .Z(n50097) );
  IV U49888 ( .A(p_input[1429]), .Z(n49742) );
  XOR U49889 ( .A(n50099), .B(n50100), .Z(n50095) );
  AND U49890 ( .A(n50101), .B(n50102), .Z(n50100) );
  XNOR U49891 ( .A(p_input[1460]), .B(n50099), .Z(n50102) );
  XNOR U49892 ( .A(n50099), .B(n49751), .Z(n50101) );
  IV U49893 ( .A(p_input[1428]), .Z(n49751) );
  XOR U49894 ( .A(n50103), .B(n50104), .Z(n50099) );
  AND U49895 ( .A(n50105), .B(n50106), .Z(n50104) );
  XNOR U49896 ( .A(p_input[1459]), .B(n50103), .Z(n50106) );
  XNOR U49897 ( .A(n50103), .B(n49760), .Z(n50105) );
  IV U49898 ( .A(p_input[1427]), .Z(n49760) );
  XOR U49899 ( .A(n50107), .B(n50108), .Z(n50103) );
  AND U49900 ( .A(n50109), .B(n50110), .Z(n50108) );
  XNOR U49901 ( .A(p_input[1458]), .B(n50107), .Z(n50110) );
  XNOR U49902 ( .A(n50107), .B(n49769), .Z(n50109) );
  IV U49903 ( .A(p_input[1426]), .Z(n49769) );
  XOR U49904 ( .A(n50111), .B(n50112), .Z(n50107) );
  AND U49905 ( .A(n50113), .B(n50114), .Z(n50112) );
  XNOR U49906 ( .A(p_input[1457]), .B(n50111), .Z(n50114) );
  XNOR U49907 ( .A(n50111), .B(n49778), .Z(n50113) );
  IV U49908 ( .A(p_input[1425]), .Z(n49778) );
  XOR U49909 ( .A(n50115), .B(n50116), .Z(n50111) );
  AND U49910 ( .A(n50117), .B(n50118), .Z(n50116) );
  XNOR U49911 ( .A(p_input[1456]), .B(n50115), .Z(n50118) );
  XNOR U49912 ( .A(n50115), .B(n49787), .Z(n50117) );
  IV U49913 ( .A(p_input[1424]), .Z(n49787) );
  XOR U49914 ( .A(n50119), .B(n50120), .Z(n50115) );
  AND U49915 ( .A(n50121), .B(n50122), .Z(n50120) );
  XNOR U49916 ( .A(p_input[1455]), .B(n50119), .Z(n50122) );
  XNOR U49917 ( .A(n50119), .B(n49796), .Z(n50121) );
  IV U49918 ( .A(p_input[1423]), .Z(n49796) );
  XOR U49919 ( .A(n50123), .B(n50124), .Z(n50119) );
  AND U49920 ( .A(n50125), .B(n50126), .Z(n50124) );
  XNOR U49921 ( .A(p_input[1454]), .B(n50123), .Z(n50126) );
  XNOR U49922 ( .A(n50123), .B(n49805), .Z(n50125) );
  IV U49923 ( .A(p_input[1422]), .Z(n49805) );
  XOR U49924 ( .A(n50127), .B(n50128), .Z(n50123) );
  AND U49925 ( .A(n50129), .B(n50130), .Z(n50128) );
  XNOR U49926 ( .A(p_input[1453]), .B(n50127), .Z(n50130) );
  XNOR U49927 ( .A(n50127), .B(n49814), .Z(n50129) );
  IV U49928 ( .A(p_input[1421]), .Z(n49814) );
  XOR U49929 ( .A(n50131), .B(n50132), .Z(n50127) );
  AND U49930 ( .A(n50133), .B(n50134), .Z(n50132) );
  XNOR U49931 ( .A(p_input[1452]), .B(n50131), .Z(n50134) );
  XNOR U49932 ( .A(n50131), .B(n49823), .Z(n50133) );
  IV U49933 ( .A(p_input[1420]), .Z(n49823) );
  XOR U49934 ( .A(n50135), .B(n50136), .Z(n50131) );
  AND U49935 ( .A(n50137), .B(n50138), .Z(n50136) );
  XNOR U49936 ( .A(p_input[1451]), .B(n50135), .Z(n50138) );
  XNOR U49937 ( .A(n50135), .B(n49832), .Z(n50137) );
  IV U49938 ( .A(p_input[1419]), .Z(n49832) );
  XOR U49939 ( .A(n50139), .B(n50140), .Z(n50135) );
  AND U49940 ( .A(n50141), .B(n50142), .Z(n50140) );
  XNOR U49941 ( .A(p_input[1450]), .B(n50139), .Z(n50142) );
  XNOR U49942 ( .A(n50139), .B(n49841), .Z(n50141) );
  IV U49943 ( .A(p_input[1418]), .Z(n49841) );
  XOR U49944 ( .A(n50143), .B(n50144), .Z(n50139) );
  AND U49945 ( .A(n50145), .B(n50146), .Z(n50144) );
  XNOR U49946 ( .A(p_input[1449]), .B(n50143), .Z(n50146) );
  XNOR U49947 ( .A(n50143), .B(n49850), .Z(n50145) );
  IV U49948 ( .A(p_input[1417]), .Z(n49850) );
  XOR U49949 ( .A(n50147), .B(n50148), .Z(n50143) );
  AND U49950 ( .A(n50149), .B(n50150), .Z(n50148) );
  XNOR U49951 ( .A(p_input[1448]), .B(n50147), .Z(n50150) );
  XNOR U49952 ( .A(n50147), .B(n49859), .Z(n50149) );
  IV U49953 ( .A(p_input[1416]), .Z(n49859) );
  XOR U49954 ( .A(n50151), .B(n50152), .Z(n50147) );
  AND U49955 ( .A(n50153), .B(n50154), .Z(n50152) );
  XNOR U49956 ( .A(p_input[1447]), .B(n50151), .Z(n50154) );
  XNOR U49957 ( .A(n50151), .B(n49868), .Z(n50153) );
  IV U49958 ( .A(p_input[1415]), .Z(n49868) );
  XOR U49959 ( .A(n50155), .B(n50156), .Z(n50151) );
  AND U49960 ( .A(n50157), .B(n50158), .Z(n50156) );
  XNOR U49961 ( .A(p_input[1446]), .B(n50155), .Z(n50158) );
  XNOR U49962 ( .A(n50155), .B(n49877), .Z(n50157) );
  IV U49963 ( .A(p_input[1414]), .Z(n49877) );
  XOR U49964 ( .A(n50159), .B(n50160), .Z(n50155) );
  AND U49965 ( .A(n50161), .B(n50162), .Z(n50160) );
  XNOR U49966 ( .A(p_input[1445]), .B(n50159), .Z(n50162) );
  XNOR U49967 ( .A(n50159), .B(n49886), .Z(n50161) );
  IV U49968 ( .A(p_input[1413]), .Z(n49886) );
  XOR U49969 ( .A(n50163), .B(n50164), .Z(n50159) );
  AND U49970 ( .A(n50165), .B(n50166), .Z(n50164) );
  XNOR U49971 ( .A(p_input[1444]), .B(n50163), .Z(n50166) );
  XNOR U49972 ( .A(n50163), .B(n49895), .Z(n50165) );
  IV U49973 ( .A(p_input[1412]), .Z(n49895) );
  XOR U49974 ( .A(n50167), .B(n50168), .Z(n50163) );
  AND U49975 ( .A(n50169), .B(n50170), .Z(n50168) );
  XNOR U49976 ( .A(p_input[1443]), .B(n50167), .Z(n50170) );
  XNOR U49977 ( .A(n50167), .B(n49904), .Z(n50169) );
  IV U49978 ( .A(p_input[1411]), .Z(n49904) );
  XOR U49979 ( .A(n50171), .B(n50172), .Z(n50167) );
  AND U49980 ( .A(n50173), .B(n50174), .Z(n50172) );
  XNOR U49981 ( .A(p_input[1442]), .B(n50171), .Z(n50174) );
  XNOR U49982 ( .A(n50171), .B(n49913), .Z(n50173) );
  IV U49983 ( .A(p_input[1410]), .Z(n49913) );
  XNOR U49984 ( .A(n50175), .B(n50176), .Z(n50171) );
  AND U49985 ( .A(n50177), .B(n50178), .Z(n50176) );
  XOR U49986 ( .A(p_input[1441]), .B(n50175), .Z(n50178) );
  XNOR U49987 ( .A(p_input[1409]), .B(n50175), .Z(n50177) );
  AND U49988 ( .A(p_input[1440]), .B(n50179), .Z(n50175) );
  IV U49989 ( .A(p_input[1408]), .Z(n50179) );
  XOR U49990 ( .A(n50180), .B(n50181), .Z(n49269) );
  AND U49991 ( .A(n633), .B(n50182), .Z(n50181) );
  XNOR U49992 ( .A(n50183), .B(n50180), .Z(n50182) );
  XOR U49993 ( .A(n50184), .B(n50185), .Z(n633) );
  AND U49994 ( .A(n50186), .B(n50187), .Z(n50185) );
  XNOR U49995 ( .A(n49284), .B(n50184), .Z(n50187) );
  AND U49996 ( .A(p_input[1407]), .B(p_input[1375]), .Z(n49284) );
  XNOR U49997 ( .A(n50184), .B(n49281), .Z(n50186) );
  IV U49998 ( .A(n50188), .Z(n49281) );
  AND U49999 ( .A(p_input[1311]), .B(p_input[1343]), .Z(n50188) );
  XOR U50000 ( .A(n50189), .B(n50190), .Z(n50184) );
  AND U50001 ( .A(n50191), .B(n50192), .Z(n50190) );
  XOR U50002 ( .A(n50189), .B(n49296), .Z(n50192) );
  XNOR U50003 ( .A(p_input[1374]), .B(n50193), .Z(n49296) );
  AND U50004 ( .A(n971), .B(n50194), .Z(n50193) );
  XOR U50005 ( .A(p_input[1406]), .B(p_input[1374]), .Z(n50194) );
  XNOR U50006 ( .A(n49293), .B(n50189), .Z(n50191) );
  XOR U50007 ( .A(n50195), .B(n50196), .Z(n49293) );
  AND U50008 ( .A(n968), .B(n50197), .Z(n50196) );
  XOR U50009 ( .A(p_input[1342]), .B(p_input[1310]), .Z(n50197) );
  XOR U50010 ( .A(n50198), .B(n50199), .Z(n50189) );
  AND U50011 ( .A(n50200), .B(n50201), .Z(n50199) );
  XOR U50012 ( .A(n50198), .B(n49308), .Z(n50201) );
  XNOR U50013 ( .A(p_input[1373]), .B(n50202), .Z(n49308) );
  AND U50014 ( .A(n971), .B(n50203), .Z(n50202) );
  XOR U50015 ( .A(p_input[1405]), .B(p_input[1373]), .Z(n50203) );
  XNOR U50016 ( .A(n49305), .B(n50198), .Z(n50200) );
  XOR U50017 ( .A(n50204), .B(n50205), .Z(n49305) );
  AND U50018 ( .A(n968), .B(n50206), .Z(n50205) );
  XOR U50019 ( .A(p_input[1341]), .B(p_input[1309]), .Z(n50206) );
  XOR U50020 ( .A(n50207), .B(n50208), .Z(n50198) );
  AND U50021 ( .A(n50209), .B(n50210), .Z(n50208) );
  XOR U50022 ( .A(n50207), .B(n49320), .Z(n50210) );
  XNOR U50023 ( .A(p_input[1372]), .B(n50211), .Z(n49320) );
  AND U50024 ( .A(n971), .B(n50212), .Z(n50211) );
  XOR U50025 ( .A(p_input[1404]), .B(p_input[1372]), .Z(n50212) );
  XNOR U50026 ( .A(n49317), .B(n50207), .Z(n50209) );
  XOR U50027 ( .A(n50213), .B(n50214), .Z(n49317) );
  AND U50028 ( .A(n968), .B(n50215), .Z(n50214) );
  XOR U50029 ( .A(p_input[1340]), .B(p_input[1308]), .Z(n50215) );
  XOR U50030 ( .A(n50216), .B(n50217), .Z(n50207) );
  AND U50031 ( .A(n50218), .B(n50219), .Z(n50217) );
  XOR U50032 ( .A(n50216), .B(n49332), .Z(n50219) );
  XNOR U50033 ( .A(p_input[1371]), .B(n50220), .Z(n49332) );
  AND U50034 ( .A(n971), .B(n50221), .Z(n50220) );
  XOR U50035 ( .A(p_input[1403]), .B(p_input[1371]), .Z(n50221) );
  XNOR U50036 ( .A(n49329), .B(n50216), .Z(n50218) );
  XOR U50037 ( .A(n50222), .B(n50223), .Z(n49329) );
  AND U50038 ( .A(n968), .B(n50224), .Z(n50223) );
  XOR U50039 ( .A(p_input[1339]), .B(p_input[1307]), .Z(n50224) );
  XOR U50040 ( .A(n50225), .B(n50226), .Z(n50216) );
  AND U50041 ( .A(n50227), .B(n50228), .Z(n50226) );
  XOR U50042 ( .A(n50225), .B(n49344), .Z(n50228) );
  XNOR U50043 ( .A(p_input[1370]), .B(n50229), .Z(n49344) );
  AND U50044 ( .A(n971), .B(n50230), .Z(n50229) );
  XOR U50045 ( .A(p_input[1402]), .B(p_input[1370]), .Z(n50230) );
  XNOR U50046 ( .A(n49341), .B(n50225), .Z(n50227) );
  XOR U50047 ( .A(n50231), .B(n50232), .Z(n49341) );
  AND U50048 ( .A(n968), .B(n50233), .Z(n50232) );
  XOR U50049 ( .A(p_input[1338]), .B(p_input[1306]), .Z(n50233) );
  XOR U50050 ( .A(n50234), .B(n50235), .Z(n50225) );
  AND U50051 ( .A(n50236), .B(n50237), .Z(n50235) );
  XOR U50052 ( .A(n50234), .B(n49356), .Z(n50237) );
  XNOR U50053 ( .A(p_input[1369]), .B(n50238), .Z(n49356) );
  AND U50054 ( .A(n971), .B(n50239), .Z(n50238) );
  XOR U50055 ( .A(p_input[1401]), .B(p_input[1369]), .Z(n50239) );
  XNOR U50056 ( .A(n49353), .B(n50234), .Z(n50236) );
  XOR U50057 ( .A(n50240), .B(n50241), .Z(n49353) );
  AND U50058 ( .A(n968), .B(n50242), .Z(n50241) );
  XOR U50059 ( .A(p_input[1337]), .B(p_input[1305]), .Z(n50242) );
  XOR U50060 ( .A(n50243), .B(n50244), .Z(n50234) );
  AND U50061 ( .A(n50245), .B(n50246), .Z(n50244) );
  XOR U50062 ( .A(n50243), .B(n49368), .Z(n50246) );
  XNOR U50063 ( .A(p_input[1368]), .B(n50247), .Z(n49368) );
  AND U50064 ( .A(n971), .B(n50248), .Z(n50247) );
  XOR U50065 ( .A(p_input[1400]), .B(p_input[1368]), .Z(n50248) );
  XNOR U50066 ( .A(n49365), .B(n50243), .Z(n50245) );
  XOR U50067 ( .A(n50249), .B(n50250), .Z(n49365) );
  AND U50068 ( .A(n968), .B(n50251), .Z(n50250) );
  XOR U50069 ( .A(p_input[1336]), .B(p_input[1304]), .Z(n50251) );
  XOR U50070 ( .A(n50252), .B(n50253), .Z(n50243) );
  AND U50071 ( .A(n50254), .B(n50255), .Z(n50253) );
  XOR U50072 ( .A(n50252), .B(n49380), .Z(n50255) );
  XNOR U50073 ( .A(p_input[1367]), .B(n50256), .Z(n49380) );
  AND U50074 ( .A(n971), .B(n50257), .Z(n50256) );
  XOR U50075 ( .A(p_input[1399]), .B(p_input[1367]), .Z(n50257) );
  XNOR U50076 ( .A(n49377), .B(n50252), .Z(n50254) );
  XOR U50077 ( .A(n50258), .B(n50259), .Z(n49377) );
  AND U50078 ( .A(n968), .B(n50260), .Z(n50259) );
  XOR U50079 ( .A(p_input[1335]), .B(p_input[1303]), .Z(n50260) );
  XOR U50080 ( .A(n50261), .B(n50262), .Z(n50252) );
  AND U50081 ( .A(n50263), .B(n50264), .Z(n50262) );
  XOR U50082 ( .A(n50261), .B(n49392), .Z(n50264) );
  XNOR U50083 ( .A(p_input[1366]), .B(n50265), .Z(n49392) );
  AND U50084 ( .A(n971), .B(n50266), .Z(n50265) );
  XOR U50085 ( .A(p_input[1398]), .B(p_input[1366]), .Z(n50266) );
  XNOR U50086 ( .A(n49389), .B(n50261), .Z(n50263) );
  XOR U50087 ( .A(n50267), .B(n50268), .Z(n49389) );
  AND U50088 ( .A(n968), .B(n50269), .Z(n50268) );
  XOR U50089 ( .A(p_input[1334]), .B(p_input[1302]), .Z(n50269) );
  XOR U50090 ( .A(n50270), .B(n50271), .Z(n50261) );
  AND U50091 ( .A(n50272), .B(n50273), .Z(n50271) );
  XOR U50092 ( .A(n50270), .B(n49404), .Z(n50273) );
  XNOR U50093 ( .A(p_input[1365]), .B(n50274), .Z(n49404) );
  AND U50094 ( .A(n971), .B(n50275), .Z(n50274) );
  XOR U50095 ( .A(p_input[1397]), .B(p_input[1365]), .Z(n50275) );
  XNOR U50096 ( .A(n49401), .B(n50270), .Z(n50272) );
  XOR U50097 ( .A(n50276), .B(n50277), .Z(n49401) );
  AND U50098 ( .A(n968), .B(n50278), .Z(n50277) );
  XOR U50099 ( .A(p_input[1333]), .B(p_input[1301]), .Z(n50278) );
  XOR U50100 ( .A(n50279), .B(n50280), .Z(n50270) );
  AND U50101 ( .A(n50281), .B(n50282), .Z(n50280) );
  XOR U50102 ( .A(n50279), .B(n49416), .Z(n50282) );
  XNOR U50103 ( .A(p_input[1364]), .B(n50283), .Z(n49416) );
  AND U50104 ( .A(n971), .B(n50284), .Z(n50283) );
  XOR U50105 ( .A(p_input[1396]), .B(p_input[1364]), .Z(n50284) );
  XNOR U50106 ( .A(n49413), .B(n50279), .Z(n50281) );
  XOR U50107 ( .A(n50285), .B(n50286), .Z(n49413) );
  AND U50108 ( .A(n968), .B(n50287), .Z(n50286) );
  XOR U50109 ( .A(p_input[1332]), .B(p_input[1300]), .Z(n50287) );
  XOR U50110 ( .A(n50288), .B(n50289), .Z(n50279) );
  AND U50111 ( .A(n50290), .B(n50291), .Z(n50289) );
  XOR U50112 ( .A(n50288), .B(n49428), .Z(n50291) );
  XNOR U50113 ( .A(p_input[1363]), .B(n50292), .Z(n49428) );
  AND U50114 ( .A(n971), .B(n50293), .Z(n50292) );
  XOR U50115 ( .A(p_input[1395]), .B(p_input[1363]), .Z(n50293) );
  XNOR U50116 ( .A(n49425), .B(n50288), .Z(n50290) );
  XOR U50117 ( .A(n50294), .B(n50295), .Z(n49425) );
  AND U50118 ( .A(n968), .B(n50296), .Z(n50295) );
  XOR U50119 ( .A(p_input[1331]), .B(p_input[1299]), .Z(n50296) );
  XOR U50120 ( .A(n50297), .B(n50298), .Z(n50288) );
  AND U50121 ( .A(n50299), .B(n50300), .Z(n50298) );
  XOR U50122 ( .A(n50297), .B(n49440), .Z(n50300) );
  XNOR U50123 ( .A(p_input[1362]), .B(n50301), .Z(n49440) );
  AND U50124 ( .A(n971), .B(n50302), .Z(n50301) );
  XOR U50125 ( .A(p_input[1394]), .B(p_input[1362]), .Z(n50302) );
  XNOR U50126 ( .A(n49437), .B(n50297), .Z(n50299) );
  XOR U50127 ( .A(n50303), .B(n50304), .Z(n49437) );
  AND U50128 ( .A(n968), .B(n50305), .Z(n50304) );
  XOR U50129 ( .A(p_input[1330]), .B(p_input[1298]), .Z(n50305) );
  XOR U50130 ( .A(n50306), .B(n50307), .Z(n50297) );
  AND U50131 ( .A(n50308), .B(n50309), .Z(n50307) );
  XOR U50132 ( .A(n50306), .B(n49452), .Z(n50309) );
  XNOR U50133 ( .A(p_input[1361]), .B(n50310), .Z(n49452) );
  AND U50134 ( .A(n971), .B(n50311), .Z(n50310) );
  XOR U50135 ( .A(p_input[1393]), .B(p_input[1361]), .Z(n50311) );
  XNOR U50136 ( .A(n49449), .B(n50306), .Z(n50308) );
  XOR U50137 ( .A(n50312), .B(n50313), .Z(n49449) );
  AND U50138 ( .A(n968), .B(n50314), .Z(n50313) );
  XOR U50139 ( .A(p_input[1329]), .B(p_input[1297]), .Z(n50314) );
  XOR U50140 ( .A(n50315), .B(n50316), .Z(n50306) );
  AND U50141 ( .A(n50317), .B(n50318), .Z(n50316) );
  XOR U50142 ( .A(n50315), .B(n49464), .Z(n50318) );
  XNOR U50143 ( .A(p_input[1360]), .B(n50319), .Z(n49464) );
  AND U50144 ( .A(n971), .B(n50320), .Z(n50319) );
  XOR U50145 ( .A(p_input[1392]), .B(p_input[1360]), .Z(n50320) );
  XNOR U50146 ( .A(n49461), .B(n50315), .Z(n50317) );
  XOR U50147 ( .A(n50321), .B(n50322), .Z(n49461) );
  AND U50148 ( .A(n968), .B(n50323), .Z(n50322) );
  XOR U50149 ( .A(p_input[1328]), .B(p_input[1296]), .Z(n50323) );
  XOR U50150 ( .A(n50324), .B(n50325), .Z(n50315) );
  AND U50151 ( .A(n50326), .B(n50327), .Z(n50325) );
  XOR U50152 ( .A(n50324), .B(n49476), .Z(n50327) );
  XNOR U50153 ( .A(p_input[1359]), .B(n50328), .Z(n49476) );
  AND U50154 ( .A(n971), .B(n50329), .Z(n50328) );
  XOR U50155 ( .A(p_input[1391]), .B(p_input[1359]), .Z(n50329) );
  XNOR U50156 ( .A(n49473), .B(n50324), .Z(n50326) );
  XOR U50157 ( .A(n50330), .B(n50331), .Z(n49473) );
  AND U50158 ( .A(n968), .B(n50332), .Z(n50331) );
  XOR U50159 ( .A(p_input[1327]), .B(p_input[1295]), .Z(n50332) );
  XOR U50160 ( .A(n50333), .B(n50334), .Z(n50324) );
  AND U50161 ( .A(n50335), .B(n50336), .Z(n50334) );
  XOR U50162 ( .A(n50333), .B(n49488), .Z(n50336) );
  XNOR U50163 ( .A(p_input[1358]), .B(n50337), .Z(n49488) );
  AND U50164 ( .A(n971), .B(n50338), .Z(n50337) );
  XOR U50165 ( .A(p_input[1390]), .B(p_input[1358]), .Z(n50338) );
  XNOR U50166 ( .A(n49485), .B(n50333), .Z(n50335) );
  XOR U50167 ( .A(n50339), .B(n50340), .Z(n49485) );
  AND U50168 ( .A(n968), .B(n50341), .Z(n50340) );
  XOR U50169 ( .A(p_input[1326]), .B(p_input[1294]), .Z(n50341) );
  XOR U50170 ( .A(n50342), .B(n50343), .Z(n50333) );
  AND U50171 ( .A(n50344), .B(n50345), .Z(n50343) );
  XOR U50172 ( .A(n50342), .B(n49500), .Z(n50345) );
  XNOR U50173 ( .A(p_input[1357]), .B(n50346), .Z(n49500) );
  AND U50174 ( .A(n971), .B(n50347), .Z(n50346) );
  XOR U50175 ( .A(p_input[1389]), .B(p_input[1357]), .Z(n50347) );
  XNOR U50176 ( .A(n49497), .B(n50342), .Z(n50344) );
  XOR U50177 ( .A(n50348), .B(n50349), .Z(n49497) );
  AND U50178 ( .A(n968), .B(n50350), .Z(n50349) );
  XOR U50179 ( .A(p_input[1325]), .B(p_input[1293]), .Z(n50350) );
  XOR U50180 ( .A(n50351), .B(n50352), .Z(n50342) );
  AND U50181 ( .A(n50353), .B(n50354), .Z(n50352) );
  XOR U50182 ( .A(n50351), .B(n49512), .Z(n50354) );
  XNOR U50183 ( .A(p_input[1356]), .B(n50355), .Z(n49512) );
  AND U50184 ( .A(n971), .B(n50356), .Z(n50355) );
  XOR U50185 ( .A(p_input[1388]), .B(p_input[1356]), .Z(n50356) );
  XNOR U50186 ( .A(n49509), .B(n50351), .Z(n50353) );
  XOR U50187 ( .A(n50357), .B(n50358), .Z(n49509) );
  AND U50188 ( .A(n968), .B(n50359), .Z(n50358) );
  XOR U50189 ( .A(p_input[1324]), .B(p_input[1292]), .Z(n50359) );
  XOR U50190 ( .A(n50360), .B(n50361), .Z(n50351) );
  AND U50191 ( .A(n50362), .B(n50363), .Z(n50361) );
  XOR U50192 ( .A(n50360), .B(n49524), .Z(n50363) );
  XNOR U50193 ( .A(p_input[1355]), .B(n50364), .Z(n49524) );
  AND U50194 ( .A(n971), .B(n50365), .Z(n50364) );
  XOR U50195 ( .A(p_input[1387]), .B(p_input[1355]), .Z(n50365) );
  XNOR U50196 ( .A(n49521), .B(n50360), .Z(n50362) );
  XOR U50197 ( .A(n50366), .B(n50367), .Z(n49521) );
  AND U50198 ( .A(n968), .B(n50368), .Z(n50367) );
  XOR U50199 ( .A(p_input[1323]), .B(p_input[1291]), .Z(n50368) );
  XOR U50200 ( .A(n50369), .B(n50370), .Z(n50360) );
  AND U50201 ( .A(n50371), .B(n50372), .Z(n50370) );
  XOR U50202 ( .A(n50369), .B(n49536), .Z(n50372) );
  XNOR U50203 ( .A(p_input[1354]), .B(n50373), .Z(n49536) );
  AND U50204 ( .A(n971), .B(n50374), .Z(n50373) );
  XOR U50205 ( .A(p_input[1386]), .B(p_input[1354]), .Z(n50374) );
  XNOR U50206 ( .A(n49533), .B(n50369), .Z(n50371) );
  XOR U50207 ( .A(n50375), .B(n50376), .Z(n49533) );
  AND U50208 ( .A(n968), .B(n50377), .Z(n50376) );
  XOR U50209 ( .A(p_input[1322]), .B(p_input[1290]), .Z(n50377) );
  XOR U50210 ( .A(n50378), .B(n50379), .Z(n50369) );
  AND U50211 ( .A(n50380), .B(n50381), .Z(n50379) );
  XOR U50212 ( .A(n50378), .B(n49548), .Z(n50381) );
  XNOR U50213 ( .A(p_input[1353]), .B(n50382), .Z(n49548) );
  AND U50214 ( .A(n971), .B(n50383), .Z(n50382) );
  XOR U50215 ( .A(p_input[1385]), .B(p_input[1353]), .Z(n50383) );
  XNOR U50216 ( .A(n49545), .B(n50378), .Z(n50380) );
  XOR U50217 ( .A(n50384), .B(n50385), .Z(n49545) );
  AND U50218 ( .A(n968), .B(n50386), .Z(n50385) );
  XOR U50219 ( .A(p_input[1321]), .B(p_input[1289]), .Z(n50386) );
  XOR U50220 ( .A(n50387), .B(n50388), .Z(n50378) );
  AND U50221 ( .A(n50389), .B(n50390), .Z(n50388) );
  XOR U50222 ( .A(n50387), .B(n49560), .Z(n50390) );
  XNOR U50223 ( .A(p_input[1352]), .B(n50391), .Z(n49560) );
  AND U50224 ( .A(n971), .B(n50392), .Z(n50391) );
  XOR U50225 ( .A(p_input[1384]), .B(p_input[1352]), .Z(n50392) );
  XNOR U50226 ( .A(n49557), .B(n50387), .Z(n50389) );
  XOR U50227 ( .A(n50393), .B(n50394), .Z(n49557) );
  AND U50228 ( .A(n968), .B(n50395), .Z(n50394) );
  XOR U50229 ( .A(p_input[1320]), .B(p_input[1288]), .Z(n50395) );
  XOR U50230 ( .A(n50396), .B(n50397), .Z(n50387) );
  AND U50231 ( .A(n50398), .B(n50399), .Z(n50397) );
  XOR U50232 ( .A(n50396), .B(n49572), .Z(n50399) );
  XNOR U50233 ( .A(p_input[1351]), .B(n50400), .Z(n49572) );
  AND U50234 ( .A(n971), .B(n50401), .Z(n50400) );
  XOR U50235 ( .A(p_input[1383]), .B(p_input[1351]), .Z(n50401) );
  XNOR U50236 ( .A(n49569), .B(n50396), .Z(n50398) );
  XOR U50237 ( .A(n50402), .B(n50403), .Z(n49569) );
  AND U50238 ( .A(n968), .B(n50404), .Z(n50403) );
  XOR U50239 ( .A(p_input[1319]), .B(p_input[1287]), .Z(n50404) );
  XOR U50240 ( .A(n50405), .B(n50406), .Z(n50396) );
  AND U50241 ( .A(n50407), .B(n50408), .Z(n50406) );
  XOR U50242 ( .A(n50405), .B(n49584), .Z(n50408) );
  XNOR U50243 ( .A(p_input[1350]), .B(n50409), .Z(n49584) );
  AND U50244 ( .A(n971), .B(n50410), .Z(n50409) );
  XOR U50245 ( .A(p_input[1382]), .B(p_input[1350]), .Z(n50410) );
  XNOR U50246 ( .A(n49581), .B(n50405), .Z(n50407) );
  XOR U50247 ( .A(n50411), .B(n50412), .Z(n49581) );
  AND U50248 ( .A(n968), .B(n50413), .Z(n50412) );
  XOR U50249 ( .A(p_input[1318]), .B(p_input[1286]), .Z(n50413) );
  XOR U50250 ( .A(n50414), .B(n50415), .Z(n50405) );
  AND U50251 ( .A(n50416), .B(n50417), .Z(n50415) );
  XOR U50252 ( .A(n50414), .B(n49596), .Z(n50417) );
  XNOR U50253 ( .A(p_input[1349]), .B(n50418), .Z(n49596) );
  AND U50254 ( .A(n971), .B(n50419), .Z(n50418) );
  XOR U50255 ( .A(p_input[1381]), .B(p_input[1349]), .Z(n50419) );
  XNOR U50256 ( .A(n49593), .B(n50414), .Z(n50416) );
  XOR U50257 ( .A(n50420), .B(n50421), .Z(n49593) );
  AND U50258 ( .A(n968), .B(n50422), .Z(n50421) );
  XOR U50259 ( .A(p_input[1317]), .B(p_input[1285]), .Z(n50422) );
  XOR U50260 ( .A(n50423), .B(n50424), .Z(n50414) );
  AND U50261 ( .A(n50425), .B(n50426), .Z(n50424) );
  XOR U50262 ( .A(n50423), .B(n49608), .Z(n50426) );
  XNOR U50263 ( .A(p_input[1348]), .B(n50427), .Z(n49608) );
  AND U50264 ( .A(n971), .B(n50428), .Z(n50427) );
  XOR U50265 ( .A(p_input[1380]), .B(p_input[1348]), .Z(n50428) );
  XNOR U50266 ( .A(n49605), .B(n50423), .Z(n50425) );
  XOR U50267 ( .A(n50429), .B(n50430), .Z(n49605) );
  AND U50268 ( .A(n968), .B(n50431), .Z(n50430) );
  XOR U50269 ( .A(p_input[1316]), .B(p_input[1284]), .Z(n50431) );
  XOR U50270 ( .A(n50432), .B(n50433), .Z(n50423) );
  AND U50271 ( .A(n50434), .B(n50435), .Z(n50433) );
  XOR U50272 ( .A(n50432), .B(n49620), .Z(n50435) );
  XNOR U50273 ( .A(p_input[1347]), .B(n50436), .Z(n49620) );
  AND U50274 ( .A(n971), .B(n50437), .Z(n50436) );
  XOR U50275 ( .A(p_input[1379]), .B(p_input[1347]), .Z(n50437) );
  XNOR U50276 ( .A(n49617), .B(n50432), .Z(n50434) );
  XOR U50277 ( .A(n50438), .B(n50439), .Z(n49617) );
  AND U50278 ( .A(n968), .B(n50440), .Z(n50439) );
  XOR U50279 ( .A(p_input[1315]), .B(p_input[1283]), .Z(n50440) );
  XOR U50280 ( .A(n50441), .B(n50442), .Z(n50432) );
  AND U50281 ( .A(n50443), .B(n50444), .Z(n50442) );
  XOR U50282 ( .A(n50441), .B(n49632), .Z(n50444) );
  XNOR U50283 ( .A(p_input[1346]), .B(n50445), .Z(n49632) );
  AND U50284 ( .A(n971), .B(n50446), .Z(n50445) );
  XOR U50285 ( .A(p_input[1378]), .B(p_input[1346]), .Z(n50446) );
  XNOR U50286 ( .A(n49629), .B(n50441), .Z(n50443) );
  XOR U50287 ( .A(n50447), .B(n50448), .Z(n49629) );
  AND U50288 ( .A(n968), .B(n50449), .Z(n50448) );
  XOR U50289 ( .A(p_input[1314]), .B(p_input[1282]), .Z(n50449) );
  XOR U50290 ( .A(n50450), .B(n50451), .Z(n50441) );
  AND U50291 ( .A(n50452), .B(n50453), .Z(n50451) );
  XNOR U50292 ( .A(n50454), .B(n49645), .Z(n50453) );
  XNOR U50293 ( .A(p_input[1345]), .B(n50455), .Z(n49645) );
  AND U50294 ( .A(n971), .B(n50456), .Z(n50455) );
  XNOR U50295 ( .A(p_input[1377]), .B(n50457), .Z(n50456) );
  IV U50296 ( .A(p_input[1345]), .Z(n50457) );
  XNOR U50297 ( .A(n49642), .B(n50450), .Z(n50452) );
  XNOR U50298 ( .A(p_input[1281]), .B(n50458), .Z(n49642) );
  AND U50299 ( .A(n968), .B(n50459), .Z(n50458) );
  XOR U50300 ( .A(p_input[1313]), .B(p_input[1281]), .Z(n50459) );
  IV U50301 ( .A(n50454), .Z(n50450) );
  AND U50302 ( .A(n50180), .B(n50183), .Z(n50454) );
  XOR U50303 ( .A(p_input[1344]), .B(n50460), .Z(n50183) );
  AND U50304 ( .A(n971), .B(n50461), .Z(n50460) );
  XOR U50305 ( .A(p_input[1376]), .B(p_input[1344]), .Z(n50461) );
  XOR U50306 ( .A(n50462), .B(n50463), .Z(n971) );
  AND U50307 ( .A(n50464), .B(n50465), .Z(n50463) );
  XNOR U50308 ( .A(p_input[1407]), .B(n50462), .Z(n50465) );
  XOR U50309 ( .A(n50462), .B(p_input[1375]), .Z(n50464) );
  XOR U50310 ( .A(n50466), .B(n50467), .Z(n50462) );
  AND U50311 ( .A(n50468), .B(n50469), .Z(n50467) );
  XNOR U50312 ( .A(p_input[1406]), .B(n50466), .Z(n50469) );
  XOR U50313 ( .A(n50466), .B(p_input[1374]), .Z(n50468) );
  XOR U50314 ( .A(n50470), .B(n50471), .Z(n50466) );
  AND U50315 ( .A(n50472), .B(n50473), .Z(n50471) );
  XNOR U50316 ( .A(p_input[1405]), .B(n50470), .Z(n50473) );
  XOR U50317 ( .A(n50470), .B(p_input[1373]), .Z(n50472) );
  XOR U50318 ( .A(n50474), .B(n50475), .Z(n50470) );
  AND U50319 ( .A(n50476), .B(n50477), .Z(n50475) );
  XNOR U50320 ( .A(p_input[1404]), .B(n50474), .Z(n50477) );
  XOR U50321 ( .A(n50474), .B(p_input[1372]), .Z(n50476) );
  XOR U50322 ( .A(n50478), .B(n50479), .Z(n50474) );
  AND U50323 ( .A(n50480), .B(n50481), .Z(n50479) );
  XNOR U50324 ( .A(p_input[1403]), .B(n50478), .Z(n50481) );
  XOR U50325 ( .A(n50478), .B(p_input[1371]), .Z(n50480) );
  XOR U50326 ( .A(n50482), .B(n50483), .Z(n50478) );
  AND U50327 ( .A(n50484), .B(n50485), .Z(n50483) );
  XNOR U50328 ( .A(p_input[1402]), .B(n50482), .Z(n50485) );
  XOR U50329 ( .A(n50482), .B(p_input[1370]), .Z(n50484) );
  XOR U50330 ( .A(n50486), .B(n50487), .Z(n50482) );
  AND U50331 ( .A(n50488), .B(n50489), .Z(n50487) );
  XNOR U50332 ( .A(p_input[1401]), .B(n50486), .Z(n50489) );
  XOR U50333 ( .A(n50486), .B(p_input[1369]), .Z(n50488) );
  XOR U50334 ( .A(n50490), .B(n50491), .Z(n50486) );
  AND U50335 ( .A(n50492), .B(n50493), .Z(n50491) );
  XNOR U50336 ( .A(p_input[1400]), .B(n50490), .Z(n50493) );
  XOR U50337 ( .A(n50490), .B(p_input[1368]), .Z(n50492) );
  XOR U50338 ( .A(n50494), .B(n50495), .Z(n50490) );
  AND U50339 ( .A(n50496), .B(n50497), .Z(n50495) );
  XNOR U50340 ( .A(p_input[1399]), .B(n50494), .Z(n50497) );
  XOR U50341 ( .A(n50494), .B(p_input[1367]), .Z(n50496) );
  XOR U50342 ( .A(n50498), .B(n50499), .Z(n50494) );
  AND U50343 ( .A(n50500), .B(n50501), .Z(n50499) );
  XNOR U50344 ( .A(p_input[1398]), .B(n50498), .Z(n50501) );
  XOR U50345 ( .A(n50498), .B(p_input[1366]), .Z(n50500) );
  XOR U50346 ( .A(n50502), .B(n50503), .Z(n50498) );
  AND U50347 ( .A(n50504), .B(n50505), .Z(n50503) );
  XNOR U50348 ( .A(p_input[1397]), .B(n50502), .Z(n50505) );
  XOR U50349 ( .A(n50502), .B(p_input[1365]), .Z(n50504) );
  XOR U50350 ( .A(n50506), .B(n50507), .Z(n50502) );
  AND U50351 ( .A(n50508), .B(n50509), .Z(n50507) );
  XNOR U50352 ( .A(p_input[1396]), .B(n50506), .Z(n50509) );
  XOR U50353 ( .A(n50506), .B(p_input[1364]), .Z(n50508) );
  XOR U50354 ( .A(n50510), .B(n50511), .Z(n50506) );
  AND U50355 ( .A(n50512), .B(n50513), .Z(n50511) );
  XNOR U50356 ( .A(p_input[1395]), .B(n50510), .Z(n50513) );
  XOR U50357 ( .A(n50510), .B(p_input[1363]), .Z(n50512) );
  XOR U50358 ( .A(n50514), .B(n50515), .Z(n50510) );
  AND U50359 ( .A(n50516), .B(n50517), .Z(n50515) );
  XNOR U50360 ( .A(p_input[1394]), .B(n50514), .Z(n50517) );
  XOR U50361 ( .A(n50514), .B(p_input[1362]), .Z(n50516) );
  XOR U50362 ( .A(n50518), .B(n50519), .Z(n50514) );
  AND U50363 ( .A(n50520), .B(n50521), .Z(n50519) );
  XNOR U50364 ( .A(p_input[1393]), .B(n50518), .Z(n50521) );
  XOR U50365 ( .A(n50518), .B(p_input[1361]), .Z(n50520) );
  XOR U50366 ( .A(n50522), .B(n50523), .Z(n50518) );
  AND U50367 ( .A(n50524), .B(n50525), .Z(n50523) );
  XNOR U50368 ( .A(p_input[1392]), .B(n50522), .Z(n50525) );
  XOR U50369 ( .A(n50522), .B(p_input[1360]), .Z(n50524) );
  XOR U50370 ( .A(n50526), .B(n50527), .Z(n50522) );
  AND U50371 ( .A(n50528), .B(n50529), .Z(n50527) );
  XNOR U50372 ( .A(p_input[1391]), .B(n50526), .Z(n50529) );
  XOR U50373 ( .A(n50526), .B(p_input[1359]), .Z(n50528) );
  XOR U50374 ( .A(n50530), .B(n50531), .Z(n50526) );
  AND U50375 ( .A(n50532), .B(n50533), .Z(n50531) );
  XNOR U50376 ( .A(p_input[1390]), .B(n50530), .Z(n50533) );
  XOR U50377 ( .A(n50530), .B(p_input[1358]), .Z(n50532) );
  XOR U50378 ( .A(n50534), .B(n50535), .Z(n50530) );
  AND U50379 ( .A(n50536), .B(n50537), .Z(n50535) );
  XNOR U50380 ( .A(p_input[1389]), .B(n50534), .Z(n50537) );
  XOR U50381 ( .A(n50534), .B(p_input[1357]), .Z(n50536) );
  XOR U50382 ( .A(n50538), .B(n50539), .Z(n50534) );
  AND U50383 ( .A(n50540), .B(n50541), .Z(n50539) );
  XNOR U50384 ( .A(p_input[1388]), .B(n50538), .Z(n50541) );
  XOR U50385 ( .A(n50538), .B(p_input[1356]), .Z(n50540) );
  XOR U50386 ( .A(n50542), .B(n50543), .Z(n50538) );
  AND U50387 ( .A(n50544), .B(n50545), .Z(n50543) );
  XNOR U50388 ( .A(p_input[1387]), .B(n50542), .Z(n50545) );
  XOR U50389 ( .A(n50542), .B(p_input[1355]), .Z(n50544) );
  XOR U50390 ( .A(n50546), .B(n50547), .Z(n50542) );
  AND U50391 ( .A(n50548), .B(n50549), .Z(n50547) );
  XNOR U50392 ( .A(p_input[1386]), .B(n50546), .Z(n50549) );
  XOR U50393 ( .A(n50546), .B(p_input[1354]), .Z(n50548) );
  XOR U50394 ( .A(n50550), .B(n50551), .Z(n50546) );
  AND U50395 ( .A(n50552), .B(n50553), .Z(n50551) );
  XNOR U50396 ( .A(p_input[1385]), .B(n50550), .Z(n50553) );
  XOR U50397 ( .A(n50550), .B(p_input[1353]), .Z(n50552) );
  XOR U50398 ( .A(n50554), .B(n50555), .Z(n50550) );
  AND U50399 ( .A(n50556), .B(n50557), .Z(n50555) );
  XNOR U50400 ( .A(p_input[1384]), .B(n50554), .Z(n50557) );
  XOR U50401 ( .A(n50554), .B(p_input[1352]), .Z(n50556) );
  XOR U50402 ( .A(n50558), .B(n50559), .Z(n50554) );
  AND U50403 ( .A(n50560), .B(n50561), .Z(n50559) );
  XNOR U50404 ( .A(p_input[1383]), .B(n50558), .Z(n50561) );
  XOR U50405 ( .A(n50558), .B(p_input[1351]), .Z(n50560) );
  XOR U50406 ( .A(n50562), .B(n50563), .Z(n50558) );
  AND U50407 ( .A(n50564), .B(n50565), .Z(n50563) );
  XNOR U50408 ( .A(p_input[1382]), .B(n50562), .Z(n50565) );
  XOR U50409 ( .A(n50562), .B(p_input[1350]), .Z(n50564) );
  XOR U50410 ( .A(n50566), .B(n50567), .Z(n50562) );
  AND U50411 ( .A(n50568), .B(n50569), .Z(n50567) );
  XNOR U50412 ( .A(p_input[1381]), .B(n50566), .Z(n50569) );
  XOR U50413 ( .A(n50566), .B(p_input[1349]), .Z(n50568) );
  XOR U50414 ( .A(n50570), .B(n50571), .Z(n50566) );
  AND U50415 ( .A(n50572), .B(n50573), .Z(n50571) );
  XNOR U50416 ( .A(p_input[1380]), .B(n50570), .Z(n50573) );
  XOR U50417 ( .A(n50570), .B(p_input[1348]), .Z(n50572) );
  XOR U50418 ( .A(n50574), .B(n50575), .Z(n50570) );
  AND U50419 ( .A(n50576), .B(n50577), .Z(n50575) );
  XNOR U50420 ( .A(p_input[1379]), .B(n50574), .Z(n50577) );
  XOR U50421 ( .A(n50574), .B(p_input[1347]), .Z(n50576) );
  XOR U50422 ( .A(n50578), .B(n50579), .Z(n50574) );
  AND U50423 ( .A(n50580), .B(n50581), .Z(n50579) );
  XNOR U50424 ( .A(p_input[1378]), .B(n50578), .Z(n50581) );
  XOR U50425 ( .A(n50578), .B(p_input[1346]), .Z(n50580) );
  XNOR U50426 ( .A(n50582), .B(n50583), .Z(n50578) );
  AND U50427 ( .A(n50584), .B(n50585), .Z(n50583) );
  XOR U50428 ( .A(p_input[1377]), .B(n50582), .Z(n50585) );
  XNOR U50429 ( .A(p_input[1345]), .B(n50582), .Z(n50584) );
  AND U50430 ( .A(p_input[1376]), .B(n50586), .Z(n50582) );
  IV U50431 ( .A(p_input[1344]), .Z(n50586) );
  XNOR U50432 ( .A(p_input[1280]), .B(n50587), .Z(n50180) );
  AND U50433 ( .A(n968), .B(n50588), .Z(n50587) );
  XOR U50434 ( .A(p_input[1312]), .B(p_input[1280]), .Z(n50588) );
  XOR U50435 ( .A(n50589), .B(n50590), .Z(n968) );
  AND U50436 ( .A(n50591), .B(n50592), .Z(n50590) );
  XNOR U50437 ( .A(p_input[1343]), .B(n50589), .Z(n50592) );
  XOR U50438 ( .A(n50589), .B(p_input[1311]), .Z(n50591) );
  XOR U50439 ( .A(n50593), .B(n50594), .Z(n50589) );
  AND U50440 ( .A(n50595), .B(n50596), .Z(n50594) );
  XNOR U50441 ( .A(p_input[1342]), .B(n50593), .Z(n50596) );
  XNOR U50442 ( .A(n50593), .B(n50195), .Z(n50595) );
  IV U50443 ( .A(p_input[1310]), .Z(n50195) );
  XOR U50444 ( .A(n50597), .B(n50598), .Z(n50593) );
  AND U50445 ( .A(n50599), .B(n50600), .Z(n50598) );
  XNOR U50446 ( .A(p_input[1341]), .B(n50597), .Z(n50600) );
  XNOR U50447 ( .A(n50597), .B(n50204), .Z(n50599) );
  IV U50448 ( .A(p_input[1309]), .Z(n50204) );
  XOR U50449 ( .A(n50601), .B(n50602), .Z(n50597) );
  AND U50450 ( .A(n50603), .B(n50604), .Z(n50602) );
  XNOR U50451 ( .A(p_input[1340]), .B(n50601), .Z(n50604) );
  XNOR U50452 ( .A(n50601), .B(n50213), .Z(n50603) );
  IV U50453 ( .A(p_input[1308]), .Z(n50213) );
  XOR U50454 ( .A(n50605), .B(n50606), .Z(n50601) );
  AND U50455 ( .A(n50607), .B(n50608), .Z(n50606) );
  XNOR U50456 ( .A(p_input[1339]), .B(n50605), .Z(n50608) );
  XNOR U50457 ( .A(n50605), .B(n50222), .Z(n50607) );
  IV U50458 ( .A(p_input[1307]), .Z(n50222) );
  XOR U50459 ( .A(n50609), .B(n50610), .Z(n50605) );
  AND U50460 ( .A(n50611), .B(n50612), .Z(n50610) );
  XNOR U50461 ( .A(p_input[1338]), .B(n50609), .Z(n50612) );
  XNOR U50462 ( .A(n50609), .B(n50231), .Z(n50611) );
  IV U50463 ( .A(p_input[1306]), .Z(n50231) );
  XOR U50464 ( .A(n50613), .B(n50614), .Z(n50609) );
  AND U50465 ( .A(n50615), .B(n50616), .Z(n50614) );
  XNOR U50466 ( .A(p_input[1337]), .B(n50613), .Z(n50616) );
  XNOR U50467 ( .A(n50613), .B(n50240), .Z(n50615) );
  IV U50468 ( .A(p_input[1305]), .Z(n50240) );
  XOR U50469 ( .A(n50617), .B(n50618), .Z(n50613) );
  AND U50470 ( .A(n50619), .B(n50620), .Z(n50618) );
  XNOR U50471 ( .A(p_input[1336]), .B(n50617), .Z(n50620) );
  XNOR U50472 ( .A(n50617), .B(n50249), .Z(n50619) );
  IV U50473 ( .A(p_input[1304]), .Z(n50249) );
  XOR U50474 ( .A(n50621), .B(n50622), .Z(n50617) );
  AND U50475 ( .A(n50623), .B(n50624), .Z(n50622) );
  XNOR U50476 ( .A(p_input[1335]), .B(n50621), .Z(n50624) );
  XNOR U50477 ( .A(n50621), .B(n50258), .Z(n50623) );
  IV U50478 ( .A(p_input[1303]), .Z(n50258) );
  XOR U50479 ( .A(n50625), .B(n50626), .Z(n50621) );
  AND U50480 ( .A(n50627), .B(n50628), .Z(n50626) );
  XNOR U50481 ( .A(p_input[1334]), .B(n50625), .Z(n50628) );
  XNOR U50482 ( .A(n50625), .B(n50267), .Z(n50627) );
  IV U50483 ( .A(p_input[1302]), .Z(n50267) );
  XOR U50484 ( .A(n50629), .B(n50630), .Z(n50625) );
  AND U50485 ( .A(n50631), .B(n50632), .Z(n50630) );
  XNOR U50486 ( .A(p_input[1333]), .B(n50629), .Z(n50632) );
  XNOR U50487 ( .A(n50629), .B(n50276), .Z(n50631) );
  IV U50488 ( .A(p_input[1301]), .Z(n50276) );
  XOR U50489 ( .A(n50633), .B(n50634), .Z(n50629) );
  AND U50490 ( .A(n50635), .B(n50636), .Z(n50634) );
  XNOR U50491 ( .A(p_input[1332]), .B(n50633), .Z(n50636) );
  XNOR U50492 ( .A(n50633), .B(n50285), .Z(n50635) );
  IV U50493 ( .A(p_input[1300]), .Z(n50285) );
  XOR U50494 ( .A(n50637), .B(n50638), .Z(n50633) );
  AND U50495 ( .A(n50639), .B(n50640), .Z(n50638) );
  XNOR U50496 ( .A(p_input[1331]), .B(n50637), .Z(n50640) );
  XNOR U50497 ( .A(n50637), .B(n50294), .Z(n50639) );
  IV U50498 ( .A(p_input[1299]), .Z(n50294) );
  XOR U50499 ( .A(n50641), .B(n50642), .Z(n50637) );
  AND U50500 ( .A(n50643), .B(n50644), .Z(n50642) );
  XNOR U50501 ( .A(p_input[1330]), .B(n50641), .Z(n50644) );
  XNOR U50502 ( .A(n50641), .B(n50303), .Z(n50643) );
  IV U50503 ( .A(p_input[1298]), .Z(n50303) );
  XOR U50504 ( .A(n50645), .B(n50646), .Z(n50641) );
  AND U50505 ( .A(n50647), .B(n50648), .Z(n50646) );
  XNOR U50506 ( .A(p_input[1329]), .B(n50645), .Z(n50648) );
  XNOR U50507 ( .A(n50645), .B(n50312), .Z(n50647) );
  IV U50508 ( .A(p_input[1297]), .Z(n50312) );
  XOR U50509 ( .A(n50649), .B(n50650), .Z(n50645) );
  AND U50510 ( .A(n50651), .B(n50652), .Z(n50650) );
  XNOR U50511 ( .A(p_input[1328]), .B(n50649), .Z(n50652) );
  XNOR U50512 ( .A(n50649), .B(n50321), .Z(n50651) );
  IV U50513 ( .A(p_input[1296]), .Z(n50321) );
  XOR U50514 ( .A(n50653), .B(n50654), .Z(n50649) );
  AND U50515 ( .A(n50655), .B(n50656), .Z(n50654) );
  XNOR U50516 ( .A(p_input[1327]), .B(n50653), .Z(n50656) );
  XNOR U50517 ( .A(n50653), .B(n50330), .Z(n50655) );
  IV U50518 ( .A(p_input[1295]), .Z(n50330) );
  XOR U50519 ( .A(n50657), .B(n50658), .Z(n50653) );
  AND U50520 ( .A(n50659), .B(n50660), .Z(n50658) );
  XNOR U50521 ( .A(p_input[1326]), .B(n50657), .Z(n50660) );
  XNOR U50522 ( .A(n50657), .B(n50339), .Z(n50659) );
  IV U50523 ( .A(p_input[1294]), .Z(n50339) );
  XOR U50524 ( .A(n50661), .B(n50662), .Z(n50657) );
  AND U50525 ( .A(n50663), .B(n50664), .Z(n50662) );
  XNOR U50526 ( .A(p_input[1325]), .B(n50661), .Z(n50664) );
  XNOR U50527 ( .A(n50661), .B(n50348), .Z(n50663) );
  IV U50528 ( .A(p_input[1293]), .Z(n50348) );
  XOR U50529 ( .A(n50665), .B(n50666), .Z(n50661) );
  AND U50530 ( .A(n50667), .B(n50668), .Z(n50666) );
  XNOR U50531 ( .A(p_input[1324]), .B(n50665), .Z(n50668) );
  XNOR U50532 ( .A(n50665), .B(n50357), .Z(n50667) );
  IV U50533 ( .A(p_input[1292]), .Z(n50357) );
  XOR U50534 ( .A(n50669), .B(n50670), .Z(n50665) );
  AND U50535 ( .A(n50671), .B(n50672), .Z(n50670) );
  XNOR U50536 ( .A(p_input[1323]), .B(n50669), .Z(n50672) );
  XNOR U50537 ( .A(n50669), .B(n50366), .Z(n50671) );
  IV U50538 ( .A(p_input[1291]), .Z(n50366) );
  XOR U50539 ( .A(n50673), .B(n50674), .Z(n50669) );
  AND U50540 ( .A(n50675), .B(n50676), .Z(n50674) );
  XNOR U50541 ( .A(p_input[1322]), .B(n50673), .Z(n50676) );
  XNOR U50542 ( .A(n50673), .B(n50375), .Z(n50675) );
  IV U50543 ( .A(p_input[1290]), .Z(n50375) );
  XOR U50544 ( .A(n50677), .B(n50678), .Z(n50673) );
  AND U50545 ( .A(n50679), .B(n50680), .Z(n50678) );
  XNOR U50546 ( .A(p_input[1321]), .B(n50677), .Z(n50680) );
  XNOR U50547 ( .A(n50677), .B(n50384), .Z(n50679) );
  IV U50548 ( .A(p_input[1289]), .Z(n50384) );
  XOR U50549 ( .A(n50681), .B(n50682), .Z(n50677) );
  AND U50550 ( .A(n50683), .B(n50684), .Z(n50682) );
  XNOR U50551 ( .A(p_input[1320]), .B(n50681), .Z(n50684) );
  XNOR U50552 ( .A(n50681), .B(n50393), .Z(n50683) );
  IV U50553 ( .A(p_input[1288]), .Z(n50393) );
  XOR U50554 ( .A(n50685), .B(n50686), .Z(n50681) );
  AND U50555 ( .A(n50687), .B(n50688), .Z(n50686) );
  XNOR U50556 ( .A(p_input[1319]), .B(n50685), .Z(n50688) );
  XNOR U50557 ( .A(n50685), .B(n50402), .Z(n50687) );
  IV U50558 ( .A(p_input[1287]), .Z(n50402) );
  XOR U50559 ( .A(n50689), .B(n50690), .Z(n50685) );
  AND U50560 ( .A(n50691), .B(n50692), .Z(n50690) );
  XNOR U50561 ( .A(p_input[1318]), .B(n50689), .Z(n50692) );
  XNOR U50562 ( .A(n50689), .B(n50411), .Z(n50691) );
  IV U50563 ( .A(p_input[1286]), .Z(n50411) );
  XOR U50564 ( .A(n50693), .B(n50694), .Z(n50689) );
  AND U50565 ( .A(n50695), .B(n50696), .Z(n50694) );
  XNOR U50566 ( .A(p_input[1317]), .B(n50693), .Z(n50696) );
  XNOR U50567 ( .A(n50693), .B(n50420), .Z(n50695) );
  IV U50568 ( .A(p_input[1285]), .Z(n50420) );
  XOR U50569 ( .A(n50697), .B(n50698), .Z(n50693) );
  AND U50570 ( .A(n50699), .B(n50700), .Z(n50698) );
  XNOR U50571 ( .A(p_input[1316]), .B(n50697), .Z(n50700) );
  XNOR U50572 ( .A(n50697), .B(n50429), .Z(n50699) );
  IV U50573 ( .A(p_input[1284]), .Z(n50429) );
  XOR U50574 ( .A(n50701), .B(n50702), .Z(n50697) );
  AND U50575 ( .A(n50703), .B(n50704), .Z(n50702) );
  XNOR U50576 ( .A(p_input[1315]), .B(n50701), .Z(n50704) );
  XNOR U50577 ( .A(n50701), .B(n50438), .Z(n50703) );
  IV U50578 ( .A(p_input[1283]), .Z(n50438) );
  XOR U50579 ( .A(n50705), .B(n50706), .Z(n50701) );
  AND U50580 ( .A(n50707), .B(n50708), .Z(n50706) );
  XNOR U50581 ( .A(p_input[1314]), .B(n50705), .Z(n50708) );
  XNOR U50582 ( .A(n50705), .B(n50447), .Z(n50707) );
  IV U50583 ( .A(p_input[1282]), .Z(n50447) );
  XNOR U50584 ( .A(n50709), .B(n50710), .Z(n50705) );
  AND U50585 ( .A(n50711), .B(n50712), .Z(n50710) );
  XOR U50586 ( .A(p_input[1313]), .B(n50709), .Z(n50712) );
  XNOR U50587 ( .A(p_input[1281]), .B(n50709), .Z(n50711) );
  AND U50588 ( .A(p_input[1312]), .B(n50713), .Z(n50709) );
  IV U50589 ( .A(p_input[1280]), .Z(n50713) );
  XOR U50590 ( .A(n50714), .B(n50715), .Z(n48892) );
  AND U50591 ( .A(n904), .B(n50716), .Z(n50715) );
  XNOR U50592 ( .A(n50717), .B(n50714), .Z(n50716) );
  XOR U50593 ( .A(n50718), .B(n50719), .Z(n904) );
  AND U50594 ( .A(n50720), .B(n50721), .Z(n50719) );
  XOR U50595 ( .A(n50718), .B(n48907), .Z(n50721) );
  XNOR U50596 ( .A(n50722), .B(n50723), .Z(n48907) );
  AND U50597 ( .A(n50724), .B(n639), .Z(n50723) );
  AND U50598 ( .A(n50722), .B(n50725), .Z(n50724) );
  XNOR U50599 ( .A(n48904), .B(n50718), .Z(n50720) );
  XOR U50600 ( .A(n50726), .B(n50727), .Z(n48904) );
  AND U50601 ( .A(n50728), .B(n636), .Z(n50727) );
  NOR U50602 ( .A(n50726), .B(n50729), .Z(n50728) );
  XOR U50603 ( .A(n50730), .B(n50731), .Z(n50718) );
  AND U50604 ( .A(n50732), .B(n50733), .Z(n50731) );
  XOR U50605 ( .A(n50730), .B(n48919), .Z(n50733) );
  XOR U50606 ( .A(n50734), .B(n50735), .Z(n48919) );
  AND U50607 ( .A(n639), .B(n50736), .Z(n50735) );
  XOR U50608 ( .A(n50737), .B(n50734), .Z(n50736) );
  XNOR U50609 ( .A(n48916), .B(n50730), .Z(n50732) );
  XOR U50610 ( .A(n50738), .B(n50739), .Z(n48916) );
  AND U50611 ( .A(n636), .B(n50740), .Z(n50739) );
  XOR U50612 ( .A(n50741), .B(n50738), .Z(n50740) );
  XOR U50613 ( .A(n50742), .B(n50743), .Z(n50730) );
  AND U50614 ( .A(n50744), .B(n50745), .Z(n50743) );
  XOR U50615 ( .A(n50742), .B(n48931), .Z(n50745) );
  XOR U50616 ( .A(n50746), .B(n50747), .Z(n48931) );
  AND U50617 ( .A(n639), .B(n50748), .Z(n50747) );
  XOR U50618 ( .A(n50749), .B(n50746), .Z(n50748) );
  XNOR U50619 ( .A(n48928), .B(n50742), .Z(n50744) );
  XOR U50620 ( .A(n50750), .B(n50751), .Z(n48928) );
  AND U50621 ( .A(n636), .B(n50752), .Z(n50751) );
  XOR U50622 ( .A(n50753), .B(n50750), .Z(n50752) );
  XOR U50623 ( .A(n50754), .B(n50755), .Z(n50742) );
  AND U50624 ( .A(n50756), .B(n50757), .Z(n50755) );
  XOR U50625 ( .A(n50754), .B(n48943), .Z(n50757) );
  XOR U50626 ( .A(n50758), .B(n50759), .Z(n48943) );
  AND U50627 ( .A(n639), .B(n50760), .Z(n50759) );
  XOR U50628 ( .A(n50761), .B(n50758), .Z(n50760) );
  XNOR U50629 ( .A(n48940), .B(n50754), .Z(n50756) );
  XOR U50630 ( .A(n50762), .B(n50763), .Z(n48940) );
  AND U50631 ( .A(n636), .B(n50764), .Z(n50763) );
  XOR U50632 ( .A(n50765), .B(n50762), .Z(n50764) );
  XOR U50633 ( .A(n50766), .B(n50767), .Z(n50754) );
  AND U50634 ( .A(n50768), .B(n50769), .Z(n50767) );
  XOR U50635 ( .A(n50766), .B(n48955), .Z(n50769) );
  XOR U50636 ( .A(n50770), .B(n50771), .Z(n48955) );
  AND U50637 ( .A(n639), .B(n50772), .Z(n50771) );
  XOR U50638 ( .A(n50773), .B(n50770), .Z(n50772) );
  XNOR U50639 ( .A(n48952), .B(n50766), .Z(n50768) );
  XOR U50640 ( .A(n50774), .B(n50775), .Z(n48952) );
  AND U50641 ( .A(n636), .B(n50776), .Z(n50775) );
  XOR U50642 ( .A(n50777), .B(n50774), .Z(n50776) );
  XOR U50643 ( .A(n50778), .B(n50779), .Z(n50766) );
  AND U50644 ( .A(n50780), .B(n50781), .Z(n50779) );
  XOR U50645 ( .A(n50778), .B(n48967), .Z(n50781) );
  XOR U50646 ( .A(n50782), .B(n50783), .Z(n48967) );
  AND U50647 ( .A(n639), .B(n50784), .Z(n50783) );
  XOR U50648 ( .A(n50785), .B(n50782), .Z(n50784) );
  XNOR U50649 ( .A(n48964), .B(n50778), .Z(n50780) );
  XOR U50650 ( .A(n50786), .B(n50787), .Z(n48964) );
  AND U50651 ( .A(n636), .B(n50788), .Z(n50787) );
  XOR U50652 ( .A(n50789), .B(n50786), .Z(n50788) );
  XOR U50653 ( .A(n50790), .B(n50791), .Z(n50778) );
  AND U50654 ( .A(n50792), .B(n50793), .Z(n50791) );
  XOR U50655 ( .A(n50790), .B(n48979), .Z(n50793) );
  XOR U50656 ( .A(n50794), .B(n50795), .Z(n48979) );
  AND U50657 ( .A(n639), .B(n50796), .Z(n50795) );
  XOR U50658 ( .A(n50797), .B(n50794), .Z(n50796) );
  XNOR U50659 ( .A(n48976), .B(n50790), .Z(n50792) );
  XOR U50660 ( .A(n50798), .B(n50799), .Z(n48976) );
  AND U50661 ( .A(n636), .B(n50800), .Z(n50799) );
  XOR U50662 ( .A(n50801), .B(n50798), .Z(n50800) );
  XOR U50663 ( .A(n50802), .B(n50803), .Z(n50790) );
  AND U50664 ( .A(n50804), .B(n50805), .Z(n50803) );
  XOR U50665 ( .A(n50802), .B(n48991), .Z(n50805) );
  XOR U50666 ( .A(n50806), .B(n50807), .Z(n48991) );
  AND U50667 ( .A(n639), .B(n50808), .Z(n50807) );
  XOR U50668 ( .A(n50809), .B(n50806), .Z(n50808) );
  XNOR U50669 ( .A(n48988), .B(n50802), .Z(n50804) );
  XOR U50670 ( .A(n50810), .B(n50811), .Z(n48988) );
  AND U50671 ( .A(n636), .B(n50812), .Z(n50811) );
  XOR U50672 ( .A(n50813), .B(n50810), .Z(n50812) );
  XOR U50673 ( .A(n50814), .B(n50815), .Z(n50802) );
  AND U50674 ( .A(n50816), .B(n50817), .Z(n50815) );
  XOR U50675 ( .A(n50814), .B(n49003), .Z(n50817) );
  XOR U50676 ( .A(n50818), .B(n50819), .Z(n49003) );
  AND U50677 ( .A(n639), .B(n50820), .Z(n50819) );
  XOR U50678 ( .A(n50821), .B(n50818), .Z(n50820) );
  XNOR U50679 ( .A(n49000), .B(n50814), .Z(n50816) );
  XOR U50680 ( .A(n50822), .B(n50823), .Z(n49000) );
  AND U50681 ( .A(n636), .B(n50824), .Z(n50823) );
  XOR U50682 ( .A(n50825), .B(n50822), .Z(n50824) );
  XOR U50683 ( .A(n50826), .B(n50827), .Z(n50814) );
  AND U50684 ( .A(n50828), .B(n50829), .Z(n50827) );
  XOR U50685 ( .A(n50826), .B(n49015), .Z(n50829) );
  XOR U50686 ( .A(n50830), .B(n50831), .Z(n49015) );
  AND U50687 ( .A(n639), .B(n50832), .Z(n50831) );
  XOR U50688 ( .A(n50833), .B(n50830), .Z(n50832) );
  XNOR U50689 ( .A(n49012), .B(n50826), .Z(n50828) );
  XOR U50690 ( .A(n50834), .B(n50835), .Z(n49012) );
  AND U50691 ( .A(n636), .B(n50836), .Z(n50835) );
  XOR U50692 ( .A(n50837), .B(n50834), .Z(n50836) );
  XOR U50693 ( .A(n50838), .B(n50839), .Z(n50826) );
  AND U50694 ( .A(n50840), .B(n50841), .Z(n50839) );
  XOR U50695 ( .A(n50838), .B(n49027), .Z(n50841) );
  XOR U50696 ( .A(n50842), .B(n50843), .Z(n49027) );
  AND U50697 ( .A(n639), .B(n50844), .Z(n50843) );
  XOR U50698 ( .A(n50845), .B(n50842), .Z(n50844) );
  XNOR U50699 ( .A(n49024), .B(n50838), .Z(n50840) );
  XOR U50700 ( .A(n50846), .B(n50847), .Z(n49024) );
  AND U50701 ( .A(n636), .B(n50848), .Z(n50847) );
  XOR U50702 ( .A(n50849), .B(n50846), .Z(n50848) );
  XOR U50703 ( .A(n50850), .B(n50851), .Z(n50838) );
  AND U50704 ( .A(n50852), .B(n50853), .Z(n50851) );
  XOR U50705 ( .A(n50850), .B(n49039), .Z(n50853) );
  XOR U50706 ( .A(n50854), .B(n50855), .Z(n49039) );
  AND U50707 ( .A(n639), .B(n50856), .Z(n50855) );
  XOR U50708 ( .A(n50857), .B(n50854), .Z(n50856) );
  XNOR U50709 ( .A(n49036), .B(n50850), .Z(n50852) );
  XOR U50710 ( .A(n50858), .B(n50859), .Z(n49036) );
  AND U50711 ( .A(n636), .B(n50860), .Z(n50859) );
  XOR U50712 ( .A(n50861), .B(n50858), .Z(n50860) );
  XOR U50713 ( .A(n50862), .B(n50863), .Z(n50850) );
  AND U50714 ( .A(n50864), .B(n50865), .Z(n50863) );
  XOR U50715 ( .A(n50862), .B(n49051), .Z(n50865) );
  XOR U50716 ( .A(n50866), .B(n50867), .Z(n49051) );
  AND U50717 ( .A(n639), .B(n50868), .Z(n50867) );
  XOR U50718 ( .A(n50869), .B(n50866), .Z(n50868) );
  XNOR U50719 ( .A(n49048), .B(n50862), .Z(n50864) );
  XOR U50720 ( .A(n50870), .B(n50871), .Z(n49048) );
  AND U50721 ( .A(n636), .B(n50872), .Z(n50871) );
  XOR U50722 ( .A(n50873), .B(n50870), .Z(n50872) );
  XOR U50723 ( .A(n50874), .B(n50875), .Z(n50862) );
  AND U50724 ( .A(n50876), .B(n50877), .Z(n50875) );
  XOR U50725 ( .A(n50874), .B(n49063), .Z(n50877) );
  XOR U50726 ( .A(n50878), .B(n50879), .Z(n49063) );
  AND U50727 ( .A(n639), .B(n50880), .Z(n50879) );
  XOR U50728 ( .A(n50881), .B(n50878), .Z(n50880) );
  XNOR U50729 ( .A(n49060), .B(n50874), .Z(n50876) );
  XOR U50730 ( .A(n50882), .B(n50883), .Z(n49060) );
  AND U50731 ( .A(n636), .B(n50884), .Z(n50883) );
  XOR U50732 ( .A(n50885), .B(n50882), .Z(n50884) );
  XOR U50733 ( .A(n50886), .B(n50887), .Z(n50874) );
  AND U50734 ( .A(n50888), .B(n50889), .Z(n50887) );
  XOR U50735 ( .A(n50886), .B(n49075), .Z(n50889) );
  XOR U50736 ( .A(n50890), .B(n50891), .Z(n49075) );
  AND U50737 ( .A(n639), .B(n50892), .Z(n50891) );
  XOR U50738 ( .A(n50893), .B(n50890), .Z(n50892) );
  XNOR U50739 ( .A(n49072), .B(n50886), .Z(n50888) );
  XOR U50740 ( .A(n50894), .B(n50895), .Z(n49072) );
  AND U50741 ( .A(n636), .B(n50896), .Z(n50895) );
  XOR U50742 ( .A(n50897), .B(n50894), .Z(n50896) );
  XOR U50743 ( .A(n50898), .B(n50899), .Z(n50886) );
  AND U50744 ( .A(n50900), .B(n50901), .Z(n50899) );
  XOR U50745 ( .A(n50898), .B(n49087), .Z(n50901) );
  XOR U50746 ( .A(n50902), .B(n50903), .Z(n49087) );
  AND U50747 ( .A(n639), .B(n50904), .Z(n50903) );
  XOR U50748 ( .A(n50905), .B(n50902), .Z(n50904) );
  XNOR U50749 ( .A(n49084), .B(n50898), .Z(n50900) );
  XOR U50750 ( .A(n50906), .B(n50907), .Z(n49084) );
  AND U50751 ( .A(n636), .B(n50908), .Z(n50907) );
  XOR U50752 ( .A(n50909), .B(n50906), .Z(n50908) );
  XOR U50753 ( .A(n50910), .B(n50911), .Z(n50898) );
  AND U50754 ( .A(n50912), .B(n50913), .Z(n50911) );
  XOR U50755 ( .A(n50910), .B(n49099), .Z(n50913) );
  XOR U50756 ( .A(n50914), .B(n50915), .Z(n49099) );
  AND U50757 ( .A(n639), .B(n50916), .Z(n50915) );
  XOR U50758 ( .A(n50917), .B(n50914), .Z(n50916) );
  XNOR U50759 ( .A(n49096), .B(n50910), .Z(n50912) );
  XOR U50760 ( .A(n50918), .B(n50919), .Z(n49096) );
  AND U50761 ( .A(n636), .B(n50920), .Z(n50919) );
  XOR U50762 ( .A(n50921), .B(n50918), .Z(n50920) );
  XOR U50763 ( .A(n50922), .B(n50923), .Z(n50910) );
  AND U50764 ( .A(n50924), .B(n50925), .Z(n50923) );
  XOR U50765 ( .A(n50922), .B(n49111), .Z(n50925) );
  XOR U50766 ( .A(n50926), .B(n50927), .Z(n49111) );
  AND U50767 ( .A(n639), .B(n50928), .Z(n50927) );
  XOR U50768 ( .A(n50929), .B(n50926), .Z(n50928) );
  XNOR U50769 ( .A(n49108), .B(n50922), .Z(n50924) );
  XOR U50770 ( .A(n50930), .B(n50931), .Z(n49108) );
  AND U50771 ( .A(n636), .B(n50932), .Z(n50931) );
  XOR U50772 ( .A(n50933), .B(n50930), .Z(n50932) );
  XOR U50773 ( .A(n50934), .B(n50935), .Z(n50922) );
  AND U50774 ( .A(n50936), .B(n50937), .Z(n50935) );
  XOR U50775 ( .A(n50934), .B(n49123), .Z(n50937) );
  XOR U50776 ( .A(n50938), .B(n50939), .Z(n49123) );
  AND U50777 ( .A(n639), .B(n50940), .Z(n50939) );
  XOR U50778 ( .A(n50941), .B(n50938), .Z(n50940) );
  XNOR U50779 ( .A(n49120), .B(n50934), .Z(n50936) );
  XOR U50780 ( .A(n50942), .B(n50943), .Z(n49120) );
  AND U50781 ( .A(n636), .B(n50944), .Z(n50943) );
  XOR U50782 ( .A(n50945), .B(n50942), .Z(n50944) );
  XOR U50783 ( .A(n50946), .B(n50947), .Z(n50934) );
  AND U50784 ( .A(n50948), .B(n50949), .Z(n50947) );
  XOR U50785 ( .A(n50946), .B(n49135), .Z(n50949) );
  XOR U50786 ( .A(n50950), .B(n50951), .Z(n49135) );
  AND U50787 ( .A(n639), .B(n50952), .Z(n50951) );
  XOR U50788 ( .A(n50953), .B(n50950), .Z(n50952) );
  XNOR U50789 ( .A(n49132), .B(n50946), .Z(n50948) );
  XOR U50790 ( .A(n50954), .B(n50955), .Z(n49132) );
  AND U50791 ( .A(n636), .B(n50956), .Z(n50955) );
  XOR U50792 ( .A(n50957), .B(n50954), .Z(n50956) );
  XOR U50793 ( .A(n50958), .B(n50959), .Z(n50946) );
  AND U50794 ( .A(n50960), .B(n50961), .Z(n50959) );
  XOR U50795 ( .A(n50958), .B(n49147), .Z(n50961) );
  XOR U50796 ( .A(n50962), .B(n50963), .Z(n49147) );
  AND U50797 ( .A(n639), .B(n50964), .Z(n50963) );
  XOR U50798 ( .A(n50965), .B(n50962), .Z(n50964) );
  XNOR U50799 ( .A(n49144), .B(n50958), .Z(n50960) );
  XOR U50800 ( .A(n50966), .B(n50967), .Z(n49144) );
  AND U50801 ( .A(n636), .B(n50968), .Z(n50967) );
  XOR U50802 ( .A(n50969), .B(n50966), .Z(n50968) );
  XOR U50803 ( .A(n50970), .B(n50971), .Z(n50958) );
  AND U50804 ( .A(n50972), .B(n50973), .Z(n50971) );
  XOR U50805 ( .A(n50970), .B(n49159), .Z(n50973) );
  XOR U50806 ( .A(n50974), .B(n50975), .Z(n49159) );
  AND U50807 ( .A(n639), .B(n50976), .Z(n50975) );
  XOR U50808 ( .A(n50977), .B(n50974), .Z(n50976) );
  XNOR U50809 ( .A(n49156), .B(n50970), .Z(n50972) );
  XOR U50810 ( .A(n50978), .B(n50979), .Z(n49156) );
  AND U50811 ( .A(n636), .B(n50980), .Z(n50979) );
  XOR U50812 ( .A(n50981), .B(n50978), .Z(n50980) );
  XOR U50813 ( .A(n50982), .B(n50983), .Z(n50970) );
  AND U50814 ( .A(n50984), .B(n50985), .Z(n50983) );
  XOR U50815 ( .A(n50982), .B(n49171), .Z(n50985) );
  XOR U50816 ( .A(n50986), .B(n50987), .Z(n49171) );
  AND U50817 ( .A(n639), .B(n50988), .Z(n50987) );
  XOR U50818 ( .A(n50989), .B(n50986), .Z(n50988) );
  XNOR U50819 ( .A(n49168), .B(n50982), .Z(n50984) );
  XOR U50820 ( .A(n50990), .B(n50991), .Z(n49168) );
  AND U50821 ( .A(n636), .B(n50992), .Z(n50991) );
  XOR U50822 ( .A(n50993), .B(n50990), .Z(n50992) );
  XOR U50823 ( .A(n50994), .B(n50995), .Z(n50982) );
  AND U50824 ( .A(n50996), .B(n50997), .Z(n50995) );
  XOR U50825 ( .A(n50994), .B(n49183), .Z(n50997) );
  XOR U50826 ( .A(n50998), .B(n50999), .Z(n49183) );
  AND U50827 ( .A(n639), .B(n51000), .Z(n50999) );
  XOR U50828 ( .A(n51001), .B(n50998), .Z(n51000) );
  XNOR U50829 ( .A(n49180), .B(n50994), .Z(n50996) );
  XOR U50830 ( .A(n51002), .B(n51003), .Z(n49180) );
  AND U50831 ( .A(n636), .B(n51004), .Z(n51003) );
  XOR U50832 ( .A(n51005), .B(n51002), .Z(n51004) );
  XOR U50833 ( .A(n51006), .B(n51007), .Z(n50994) );
  AND U50834 ( .A(n51008), .B(n51009), .Z(n51007) );
  XOR U50835 ( .A(n51006), .B(n49195), .Z(n51009) );
  XOR U50836 ( .A(n51010), .B(n51011), .Z(n49195) );
  AND U50837 ( .A(n639), .B(n51012), .Z(n51011) );
  XOR U50838 ( .A(n51013), .B(n51010), .Z(n51012) );
  XNOR U50839 ( .A(n49192), .B(n51006), .Z(n51008) );
  XOR U50840 ( .A(n51014), .B(n51015), .Z(n49192) );
  AND U50841 ( .A(n636), .B(n51016), .Z(n51015) );
  XOR U50842 ( .A(n51017), .B(n51014), .Z(n51016) );
  XOR U50843 ( .A(n51018), .B(n51019), .Z(n51006) );
  AND U50844 ( .A(n51020), .B(n51021), .Z(n51019) );
  XOR U50845 ( .A(n51018), .B(n49207), .Z(n51021) );
  XOR U50846 ( .A(n51022), .B(n51023), .Z(n49207) );
  AND U50847 ( .A(n639), .B(n51024), .Z(n51023) );
  XOR U50848 ( .A(n51025), .B(n51022), .Z(n51024) );
  XNOR U50849 ( .A(n49204), .B(n51018), .Z(n51020) );
  XOR U50850 ( .A(n51026), .B(n51027), .Z(n49204) );
  AND U50851 ( .A(n636), .B(n51028), .Z(n51027) );
  XOR U50852 ( .A(n51029), .B(n51026), .Z(n51028) );
  XOR U50853 ( .A(n51030), .B(n51031), .Z(n51018) );
  AND U50854 ( .A(n51032), .B(n51033), .Z(n51031) );
  XOR U50855 ( .A(n51030), .B(n49219), .Z(n51033) );
  XOR U50856 ( .A(n51034), .B(n51035), .Z(n49219) );
  AND U50857 ( .A(n639), .B(n51036), .Z(n51035) );
  XOR U50858 ( .A(n51037), .B(n51034), .Z(n51036) );
  XNOR U50859 ( .A(n49216), .B(n51030), .Z(n51032) );
  XOR U50860 ( .A(n51038), .B(n51039), .Z(n49216) );
  AND U50861 ( .A(n636), .B(n51040), .Z(n51039) );
  XOR U50862 ( .A(n51041), .B(n51038), .Z(n51040) );
  XOR U50863 ( .A(n51042), .B(n51043), .Z(n51030) );
  AND U50864 ( .A(n51044), .B(n51045), .Z(n51043) );
  XOR U50865 ( .A(n51042), .B(n49231), .Z(n51045) );
  XOR U50866 ( .A(n51046), .B(n51047), .Z(n49231) );
  AND U50867 ( .A(n639), .B(n51048), .Z(n51047) );
  XOR U50868 ( .A(n51049), .B(n51046), .Z(n51048) );
  XNOR U50869 ( .A(n49228), .B(n51042), .Z(n51044) );
  XOR U50870 ( .A(n51050), .B(n51051), .Z(n49228) );
  AND U50871 ( .A(n636), .B(n51052), .Z(n51051) );
  XOR U50872 ( .A(n51053), .B(n51050), .Z(n51052) );
  XOR U50873 ( .A(n51054), .B(n51055), .Z(n51042) );
  AND U50874 ( .A(n51056), .B(n51057), .Z(n51055) );
  XOR U50875 ( .A(n51054), .B(n49243), .Z(n51057) );
  XOR U50876 ( .A(n51058), .B(n51059), .Z(n49243) );
  AND U50877 ( .A(n639), .B(n51060), .Z(n51059) );
  XOR U50878 ( .A(n51061), .B(n51058), .Z(n51060) );
  XNOR U50879 ( .A(n49240), .B(n51054), .Z(n51056) );
  XOR U50880 ( .A(n51062), .B(n51063), .Z(n49240) );
  AND U50881 ( .A(n636), .B(n51064), .Z(n51063) );
  XOR U50882 ( .A(n51065), .B(n51062), .Z(n51064) );
  XOR U50883 ( .A(n51066), .B(n51067), .Z(n51054) );
  AND U50884 ( .A(n51068), .B(n51069), .Z(n51067) );
  XOR U50885 ( .A(n51066), .B(n49255), .Z(n51069) );
  XOR U50886 ( .A(n51070), .B(n51071), .Z(n49255) );
  AND U50887 ( .A(n639), .B(n51072), .Z(n51071) );
  XOR U50888 ( .A(n51073), .B(n51070), .Z(n51072) );
  XNOR U50889 ( .A(n49252), .B(n51066), .Z(n51068) );
  XOR U50890 ( .A(n51074), .B(n51075), .Z(n49252) );
  AND U50891 ( .A(n636), .B(n51076), .Z(n51075) );
  XOR U50892 ( .A(n51077), .B(n51074), .Z(n51076) );
  XOR U50893 ( .A(n51078), .B(n51079), .Z(n51066) );
  AND U50894 ( .A(n51080), .B(n51081), .Z(n51079) );
  XNOR U50895 ( .A(n51082), .B(n49268), .Z(n51081) );
  XOR U50896 ( .A(n51083), .B(n51084), .Z(n49268) );
  AND U50897 ( .A(n639), .B(n51085), .Z(n51084) );
  XOR U50898 ( .A(n51083), .B(n51086), .Z(n51085) );
  XNOR U50899 ( .A(n49265), .B(n51078), .Z(n51080) );
  XOR U50900 ( .A(n51087), .B(n51088), .Z(n49265) );
  AND U50901 ( .A(n636), .B(n51089), .Z(n51088) );
  XOR U50902 ( .A(n51087), .B(n51090), .Z(n51089) );
  IV U50903 ( .A(n51082), .Z(n51078) );
  AND U50904 ( .A(n50714), .B(n50717), .Z(n51082) );
  XNOR U50905 ( .A(n51091), .B(n51092), .Z(n50717) );
  AND U50906 ( .A(n639), .B(n51093), .Z(n51092) );
  XNOR U50907 ( .A(n51094), .B(n51091), .Z(n51093) );
  XOR U50908 ( .A(n51095), .B(n51096), .Z(n639) );
  AND U50909 ( .A(n51097), .B(n51098), .Z(n51096) );
  XOR U50910 ( .A(n50725), .B(n51095), .Z(n51098) );
  IV U50911 ( .A(n51099), .Z(n50725) );
  AND U50912 ( .A(p_input[1279]), .B(p_input[1247]), .Z(n51099) );
  XOR U50913 ( .A(n51095), .B(n50722), .Z(n51097) );
  AND U50914 ( .A(p_input[1183]), .B(p_input[1215]), .Z(n50722) );
  XOR U50915 ( .A(n51100), .B(n51101), .Z(n51095) );
  AND U50916 ( .A(n51102), .B(n51103), .Z(n51101) );
  XOR U50917 ( .A(n51100), .B(n50737), .Z(n51103) );
  XNOR U50918 ( .A(p_input[1246]), .B(n51104), .Z(n50737) );
  AND U50919 ( .A(n979), .B(n51105), .Z(n51104) );
  XOR U50920 ( .A(p_input[1278]), .B(p_input[1246]), .Z(n51105) );
  XNOR U50921 ( .A(n50734), .B(n51100), .Z(n51102) );
  XOR U50922 ( .A(n51106), .B(n51107), .Z(n50734) );
  AND U50923 ( .A(n977), .B(n51108), .Z(n51107) );
  XOR U50924 ( .A(p_input[1214]), .B(p_input[1182]), .Z(n51108) );
  XOR U50925 ( .A(n51109), .B(n51110), .Z(n51100) );
  AND U50926 ( .A(n51111), .B(n51112), .Z(n51110) );
  XOR U50927 ( .A(n51109), .B(n50749), .Z(n51112) );
  XNOR U50928 ( .A(p_input[1245]), .B(n51113), .Z(n50749) );
  AND U50929 ( .A(n979), .B(n51114), .Z(n51113) );
  XOR U50930 ( .A(p_input[1277]), .B(p_input[1245]), .Z(n51114) );
  XNOR U50931 ( .A(n50746), .B(n51109), .Z(n51111) );
  XOR U50932 ( .A(n51115), .B(n51116), .Z(n50746) );
  AND U50933 ( .A(n977), .B(n51117), .Z(n51116) );
  XOR U50934 ( .A(p_input[1213]), .B(p_input[1181]), .Z(n51117) );
  XOR U50935 ( .A(n51118), .B(n51119), .Z(n51109) );
  AND U50936 ( .A(n51120), .B(n51121), .Z(n51119) );
  XOR U50937 ( .A(n51118), .B(n50761), .Z(n51121) );
  XNOR U50938 ( .A(p_input[1244]), .B(n51122), .Z(n50761) );
  AND U50939 ( .A(n979), .B(n51123), .Z(n51122) );
  XOR U50940 ( .A(p_input[1276]), .B(p_input[1244]), .Z(n51123) );
  XNOR U50941 ( .A(n50758), .B(n51118), .Z(n51120) );
  XOR U50942 ( .A(n51124), .B(n51125), .Z(n50758) );
  AND U50943 ( .A(n977), .B(n51126), .Z(n51125) );
  XOR U50944 ( .A(p_input[1212]), .B(p_input[1180]), .Z(n51126) );
  XOR U50945 ( .A(n51127), .B(n51128), .Z(n51118) );
  AND U50946 ( .A(n51129), .B(n51130), .Z(n51128) );
  XOR U50947 ( .A(n51127), .B(n50773), .Z(n51130) );
  XNOR U50948 ( .A(p_input[1243]), .B(n51131), .Z(n50773) );
  AND U50949 ( .A(n979), .B(n51132), .Z(n51131) );
  XOR U50950 ( .A(p_input[1275]), .B(p_input[1243]), .Z(n51132) );
  XNOR U50951 ( .A(n50770), .B(n51127), .Z(n51129) );
  XOR U50952 ( .A(n51133), .B(n51134), .Z(n50770) );
  AND U50953 ( .A(n977), .B(n51135), .Z(n51134) );
  XOR U50954 ( .A(p_input[1211]), .B(p_input[1179]), .Z(n51135) );
  XOR U50955 ( .A(n51136), .B(n51137), .Z(n51127) );
  AND U50956 ( .A(n51138), .B(n51139), .Z(n51137) );
  XOR U50957 ( .A(n51136), .B(n50785), .Z(n51139) );
  XNOR U50958 ( .A(p_input[1242]), .B(n51140), .Z(n50785) );
  AND U50959 ( .A(n979), .B(n51141), .Z(n51140) );
  XOR U50960 ( .A(p_input[1274]), .B(p_input[1242]), .Z(n51141) );
  XNOR U50961 ( .A(n50782), .B(n51136), .Z(n51138) );
  XOR U50962 ( .A(n51142), .B(n51143), .Z(n50782) );
  AND U50963 ( .A(n977), .B(n51144), .Z(n51143) );
  XOR U50964 ( .A(p_input[1210]), .B(p_input[1178]), .Z(n51144) );
  XOR U50965 ( .A(n51145), .B(n51146), .Z(n51136) );
  AND U50966 ( .A(n51147), .B(n51148), .Z(n51146) );
  XOR U50967 ( .A(n51145), .B(n50797), .Z(n51148) );
  XNOR U50968 ( .A(p_input[1241]), .B(n51149), .Z(n50797) );
  AND U50969 ( .A(n979), .B(n51150), .Z(n51149) );
  XOR U50970 ( .A(p_input[1273]), .B(p_input[1241]), .Z(n51150) );
  XNOR U50971 ( .A(n50794), .B(n51145), .Z(n51147) );
  XOR U50972 ( .A(n51151), .B(n51152), .Z(n50794) );
  AND U50973 ( .A(n977), .B(n51153), .Z(n51152) );
  XOR U50974 ( .A(p_input[1209]), .B(p_input[1177]), .Z(n51153) );
  XOR U50975 ( .A(n51154), .B(n51155), .Z(n51145) );
  AND U50976 ( .A(n51156), .B(n51157), .Z(n51155) );
  XOR U50977 ( .A(n51154), .B(n50809), .Z(n51157) );
  XNOR U50978 ( .A(p_input[1240]), .B(n51158), .Z(n50809) );
  AND U50979 ( .A(n979), .B(n51159), .Z(n51158) );
  XOR U50980 ( .A(p_input[1272]), .B(p_input[1240]), .Z(n51159) );
  XNOR U50981 ( .A(n50806), .B(n51154), .Z(n51156) );
  XOR U50982 ( .A(n51160), .B(n51161), .Z(n50806) );
  AND U50983 ( .A(n977), .B(n51162), .Z(n51161) );
  XOR U50984 ( .A(p_input[1208]), .B(p_input[1176]), .Z(n51162) );
  XOR U50985 ( .A(n51163), .B(n51164), .Z(n51154) );
  AND U50986 ( .A(n51165), .B(n51166), .Z(n51164) );
  XOR U50987 ( .A(n51163), .B(n50821), .Z(n51166) );
  XNOR U50988 ( .A(p_input[1239]), .B(n51167), .Z(n50821) );
  AND U50989 ( .A(n979), .B(n51168), .Z(n51167) );
  XOR U50990 ( .A(p_input[1271]), .B(p_input[1239]), .Z(n51168) );
  XNOR U50991 ( .A(n50818), .B(n51163), .Z(n51165) );
  XOR U50992 ( .A(n51169), .B(n51170), .Z(n50818) );
  AND U50993 ( .A(n977), .B(n51171), .Z(n51170) );
  XOR U50994 ( .A(p_input[1207]), .B(p_input[1175]), .Z(n51171) );
  XOR U50995 ( .A(n51172), .B(n51173), .Z(n51163) );
  AND U50996 ( .A(n51174), .B(n51175), .Z(n51173) );
  XOR U50997 ( .A(n51172), .B(n50833), .Z(n51175) );
  XNOR U50998 ( .A(p_input[1238]), .B(n51176), .Z(n50833) );
  AND U50999 ( .A(n979), .B(n51177), .Z(n51176) );
  XOR U51000 ( .A(p_input[1270]), .B(p_input[1238]), .Z(n51177) );
  XNOR U51001 ( .A(n50830), .B(n51172), .Z(n51174) );
  XOR U51002 ( .A(n51178), .B(n51179), .Z(n50830) );
  AND U51003 ( .A(n977), .B(n51180), .Z(n51179) );
  XOR U51004 ( .A(p_input[1206]), .B(p_input[1174]), .Z(n51180) );
  XOR U51005 ( .A(n51181), .B(n51182), .Z(n51172) );
  AND U51006 ( .A(n51183), .B(n51184), .Z(n51182) );
  XOR U51007 ( .A(n51181), .B(n50845), .Z(n51184) );
  XNOR U51008 ( .A(p_input[1237]), .B(n51185), .Z(n50845) );
  AND U51009 ( .A(n979), .B(n51186), .Z(n51185) );
  XOR U51010 ( .A(p_input[1269]), .B(p_input[1237]), .Z(n51186) );
  XNOR U51011 ( .A(n50842), .B(n51181), .Z(n51183) );
  XOR U51012 ( .A(n51187), .B(n51188), .Z(n50842) );
  AND U51013 ( .A(n977), .B(n51189), .Z(n51188) );
  XOR U51014 ( .A(p_input[1205]), .B(p_input[1173]), .Z(n51189) );
  XOR U51015 ( .A(n51190), .B(n51191), .Z(n51181) );
  AND U51016 ( .A(n51192), .B(n51193), .Z(n51191) );
  XOR U51017 ( .A(n51190), .B(n50857), .Z(n51193) );
  XNOR U51018 ( .A(p_input[1236]), .B(n51194), .Z(n50857) );
  AND U51019 ( .A(n979), .B(n51195), .Z(n51194) );
  XOR U51020 ( .A(p_input[1268]), .B(p_input[1236]), .Z(n51195) );
  XNOR U51021 ( .A(n50854), .B(n51190), .Z(n51192) );
  XOR U51022 ( .A(n51196), .B(n51197), .Z(n50854) );
  AND U51023 ( .A(n977), .B(n51198), .Z(n51197) );
  XOR U51024 ( .A(p_input[1204]), .B(p_input[1172]), .Z(n51198) );
  XOR U51025 ( .A(n51199), .B(n51200), .Z(n51190) );
  AND U51026 ( .A(n51201), .B(n51202), .Z(n51200) );
  XOR U51027 ( .A(n51199), .B(n50869), .Z(n51202) );
  XNOR U51028 ( .A(p_input[1235]), .B(n51203), .Z(n50869) );
  AND U51029 ( .A(n979), .B(n51204), .Z(n51203) );
  XOR U51030 ( .A(p_input[1267]), .B(p_input[1235]), .Z(n51204) );
  XNOR U51031 ( .A(n50866), .B(n51199), .Z(n51201) );
  XOR U51032 ( .A(n51205), .B(n51206), .Z(n50866) );
  AND U51033 ( .A(n977), .B(n51207), .Z(n51206) );
  XOR U51034 ( .A(p_input[1203]), .B(p_input[1171]), .Z(n51207) );
  XOR U51035 ( .A(n51208), .B(n51209), .Z(n51199) );
  AND U51036 ( .A(n51210), .B(n51211), .Z(n51209) );
  XOR U51037 ( .A(n51208), .B(n50881), .Z(n51211) );
  XNOR U51038 ( .A(p_input[1234]), .B(n51212), .Z(n50881) );
  AND U51039 ( .A(n979), .B(n51213), .Z(n51212) );
  XOR U51040 ( .A(p_input[1266]), .B(p_input[1234]), .Z(n51213) );
  XNOR U51041 ( .A(n50878), .B(n51208), .Z(n51210) );
  XOR U51042 ( .A(n51214), .B(n51215), .Z(n50878) );
  AND U51043 ( .A(n977), .B(n51216), .Z(n51215) );
  XOR U51044 ( .A(p_input[1202]), .B(p_input[1170]), .Z(n51216) );
  XOR U51045 ( .A(n51217), .B(n51218), .Z(n51208) );
  AND U51046 ( .A(n51219), .B(n51220), .Z(n51218) );
  XOR U51047 ( .A(n51217), .B(n50893), .Z(n51220) );
  XNOR U51048 ( .A(p_input[1233]), .B(n51221), .Z(n50893) );
  AND U51049 ( .A(n979), .B(n51222), .Z(n51221) );
  XOR U51050 ( .A(p_input[1265]), .B(p_input[1233]), .Z(n51222) );
  XNOR U51051 ( .A(n50890), .B(n51217), .Z(n51219) );
  XOR U51052 ( .A(n51223), .B(n51224), .Z(n50890) );
  AND U51053 ( .A(n977), .B(n51225), .Z(n51224) );
  XOR U51054 ( .A(p_input[1201]), .B(p_input[1169]), .Z(n51225) );
  XOR U51055 ( .A(n51226), .B(n51227), .Z(n51217) );
  AND U51056 ( .A(n51228), .B(n51229), .Z(n51227) );
  XOR U51057 ( .A(n51226), .B(n50905), .Z(n51229) );
  XNOR U51058 ( .A(p_input[1232]), .B(n51230), .Z(n50905) );
  AND U51059 ( .A(n979), .B(n51231), .Z(n51230) );
  XOR U51060 ( .A(p_input[1264]), .B(p_input[1232]), .Z(n51231) );
  XNOR U51061 ( .A(n50902), .B(n51226), .Z(n51228) );
  XOR U51062 ( .A(n51232), .B(n51233), .Z(n50902) );
  AND U51063 ( .A(n977), .B(n51234), .Z(n51233) );
  XOR U51064 ( .A(p_input[1200]), .B(p_input[1168]), .Z(n51234) );
  XOR U51065 ( .A(n51235), .B(n51236), .Z(n51226) );
  AND U51066 ( .A(n51237), .B(n51238), .Z(n51236) );
  XOR U51067 ( .A(n51235), .B(n50917), .Z(n51238) );
  XNOR U51068 ( .A(p_input[1231]), .B(n51239), .Z(n50917) );
  AND U51069 ( .A(n979), .B(n51240), .Z(n51239) );
  XOR U51070 ( .A(p_input[1263]), .B(p_input[1231]), .Z(n51240) );
  XNOR U51071 ( .A(n50914), .B(n51235), .Z(n51237) );
  XOR U51072 ( .A(n51241), .B(n51242), .Z(n50914) );
  AND U51073 ( .A(n977), .B(n51243), .Z(n51242) );
  XOR U51074 ( .A(p_input[1199]), .B(p_input[1167]), .Z(n51243) );
  XOR U51075 ( .A(n51244), .B(n51245), .Z(n51235) );
  AND U51076 ( .A(n51246), .B(n51247), .Z(n51245) );
  XOR U51077 ( .A(n51244), .B(n50929), .Z(n51247) );
  XNOR U51078 ( .A(p_input[1230]), .B(n51248), .Z(n50929) );
  AND U51079 ( .A(n979), .B(n51249), .Z(n51248) );
  XOR U51080 ( .A(p_input[1262]), .B(p_input[1230]), .Z(n51249) );
  XNOR U51081 ( .A(n50926), .B(n51244), .Z(n51246) );
  XOR U51082 ( .A(n51250), .B(n51251), .Z(n50926) );
  AND U51083 ( .A(n977), .B(n51252), .Z(n51251) );
  XOR U51084 ( .A(p_input[1198]), .B(p_input[1166]), .Z(n51252) );
  XOR U51085 ( .A(n51253), .B(n51254), .Z(n51244) );
  AND U51086 ( .A(n51255), .B(n51256), .Z(n51254) );
  XOR U51087 ( .A(n51253), .B(n50941), .Z(n51256) );
  XNOR U51088 ( .A(p_input[1229]), .B(n51257), .Z(n50941) );
  AND U51089 ( .A(n979), .B(n51258), .Z(n51257) );
  XOR U51090 ( .A(p_input[1261]), .B(p_input[1229]), .Z(n51258) );
  XNOR U51091 ( .A(n50938), .B(n51253), .Z(n51255) );
  XOR U51092 ( .A(n51259), .B(n51260), .Z(n50938) );
  AND U51093 ( .A(n977), .B(n51261), .Z(n51260) );
  XOR U51094 ( .A(p_input[1197]), .B(p_input[1165]), .Z(n51261) );
  XOR U51095 ( .A(n51262), .B(n51263), .Z(n51253) );
  AND U51096 ( .A(n51264), .B(n51265), .Z(n51263) );
  XOR U51097 ( .A(n51262), .B(n50953), .Z(n51265) );
  XNOR U51098 ( .A(p_input[1228]), .B(n51266), .Z(n50953) );
  AND U51099 ( .A(n979), .B(n51267), .Z(n51266) );
  XOR U51100 ( .A(p_input[1260]), .B(p_input[1228]), .Z(n51267) );
  XNOR U51101 ( .A(n50950), .B(n51262), .Z(n51264) );
  XOR U51102 ( .A(n51268), .B(n51269), .Z(n50950) );
  AND U51103 ( .A(n977), .B(n51270), .Z(n51269) );
  XOR U51104 ( .A(p_input[1196]), .B(p_input[1164]), .Z(n51270) );
  XOR U51105 ( .A(n51271), .B(n51272), .Z(n51262) );
  AND U51106 ( .A(n51273), .B(n51274), .Z(n51272) );
  XOR U51107 ( .A(n51271), .B(n50965), .Z(n51274) );
  XNOR U51108 ( .A(p_input[1227]), .B(n51275), .Z(n50965) );
  AND U51109 ( .A(n979), .B(n51276), .Z(n51275) );
  XOR U51110 ( .A(p_input[1259]), .B(p_input[1227]), .Z(n51276) );
  XNOR U51111 ( .A(n50962), .B(n51271), .Z(n51273) );
  XOR U51112 ( .A(n51277), .B(n51278), .Z(n50962) );
  AND U51113 ( .A(n977), .B(n51279), .Z(n51278) );
  XOR U51114 ( .A(p_input[1195]), .B(p_input[1163]), .Z(n51279) );
  XOR U51115 ( .A(n51280), .B(n51281), .Z(n51271) );
  AND U51116 ( .A(n51282), .B(n51283), .Z(n51281) );
  XOR U51117 ( .A(n51280), .B(n50977), .Z(n51283) );
  XNOR U51118 ( .A(p_input[1226]), .B(n51284), .Z(n50977) );
  AND U51119 ( .A(n979), .B(n51285), .Z(n51284) );
  XOR U51120 ( .A(p_input[1258]), .B(p_input[1226]), .Z(n51285) );
  XNOR U51121 ( .A(n50974), .B(n51280), .Z(n51282) );
  XOR U51122 ( .A(n51286), .B(n51287), .Z(n50974) );
  AND U51123 ( .A(n977), .B(n51288), .Z(n51287) );
  XOR U51124 ( .A(p_input[1194]), .B(p_input[1162]), .Z(n51288) );
  XOR U51125 ( .A(n51289), .B(n51290), .Z(n51280) );
  AND U51126 ( .A(n51291), .B(n51292), .Z(n51290) );
  XOR U51127 ( .A(n51289), .B(n50989), .Z(n51292) );
  XNOR U51128 ( .A(p_input[1225]), .B(n51293), .Z(n50989) );
  AND U51129 ( .A(n979), .B(n51294), .Z(n51293) );
  XOR U51130 ( .A(p_input[1257]), .B(p_input[1225]), .Z(n51294) );
  XNOR U51131 ( .A(n50986), .B(n51289), .Z(n51291) );
  XOR U51132 ( .A(n51295), .B(n51296), .Z(n50986) );
  AND U51133 ( .A(n977), .B(n51297), .Z(n51296) );
  XOR U51134 ( .A(p_input[1193]), .B(p_input[1161]), .Z(n51297) );
  XOR U51135 ( .A(n51298), .B(n51299), .Z(n51289) );
  AND U51136 ( .A(n51300), .B(n51301), .Z(n51299) );
  XOR U51137 ( .A(n51298), .B(n51001), .Z(n51301) );
  XNOR U51138 ( .A(p_input[1224]), .B(n51302), .Z(n51001) );
  AND U51139 ( .A(n979), .B(n51303), .Z(n51302) );
  XOR U51140 ( .A(p_input[1256]), .B(p_input[1224]), .Z(n51303) );
  XNOR U51141 ( .A(n50998), .B(n51298), .Z(n51300) );
  XOR U51142 ( .A(n51304), .B(n51305), .Z(n50998) );
  AND U51143 ( .A(n977), .B(n51306), .Z(n51305) );
  XOR U51144 ( .A(p_input[1192]), .B(p_input[1160]), .Z(n51306) );
  XOR U51145 ( .A(n51307), .B(n51308), .Z(n51298) );
  AND U51146 ( .A(n51309), .B(n51310), .Z(n51308) );
  XOR U51147 ( .A(n51307), .B(n51013), .Z(n51310) );
  XNOR U51148 ( .A(p_input[1223]), .B(n51311), .Z(n51013) );
  AND U51149 ( .A(n979), .B(n51312), .Z(n51311) );
  XOR U51150 ( .A(p_input[1255]), .B(p_input[1223]), .Z(n51312) );
  XNOR U51151 ( .A(n51010), .B(n51307), .Z(n51309) );
  XOR U51152 ( .A(n51313), .B(n51314), .Z(n51010) );
  AND U51153 ( .A(n977), .B(n51315), .Z(n51314) );
  XOR U51154 ( .A(p_input[1191]), .B(p_input[1159]), .Z(n51315) );
  XOR U51155 ( .A(n51316), .B(n51317), .Z(n51307) );
  AND U51156 ( .A(n51318), .B(n51319), .Z(n51317) );
  XOR U51157 ( .A(n51316), .B(n51025), .Z(n51319) );
  XNOR U51158 ( .A(p_input[1222]), .B(n51320), .Z(n51025) );
  AND U51159 ( .A(n979), .B(n51321), .Z(n51320) );
  XOR U51160 ( .A(p_input[1254]), .B(p_input[1222]), .Z(n51321) );
  XNOR U51161 ( .A(n51022), .B(n51316), .Z(n51318) );
  XOR U51162 ( .A(n51322), .B(n51323), .Z(n51022) );
  AND U51163 ( .A(n977), .B(n51324), .Z(n51323) );
  XOR U51164 ( .A(p_input[1190]), .B(p_input[1158]), .Z(n51324) );
  XOR U51165 ( .A(n51325), .B(n51326), .Z(n51316) );
  AND U51166 ( .A(n51327), .B(n51328), .Z(n51326) );
  XOR U51167 ( .A(n51325), .B(n51037), .Z(n51328) );
  XNOR U51168 ( .A(p_input[1221]), .B(n51329), .Z(n51037) );
  AND U51169 ( .A(n979), .B(n51330), .Z(n51329) );
  XOR U51170 ( .A(p_input[1253]), .B(p_input[1221]), .Z(n51330) );
  XNOR U51171 ( .A(n51034), .B(n51325), .Z(n51327) );
  XOR U51172 ( .A(n51331), .B(n51332), .Z(n51034) );
  AND U51173 ( .A(n977), .B(n51333), .Z(n51332) );
  XOR U51174 ( .A(p_input[1189]), .B(p_input[1157]), .Z(n51333) );
  XOR U51175 ( .A(n51334), .B(n51335), .Z(n51325) );
  AND U51176 ( .A(n51336), .B(n51337), .Z(n51335) );
  XOR U51177 ( .A(n51334), .B(n51049), .Z(n51337) );
  XNOR U51178 ( .A(p_input[1220]), .B(n51338), .Z(n51049) );
  AND U51179 ( .A(n979), .B(n51339), .Z(n51338) );
  XOR U51180 ( .A(p_input[1252]), .B(p_input[1220]), .Z(n51339) );
  XNOR U51181 ( .A(n51046), .B(n51334), .Z(n51336) );
  XOR U51182 ( .A(n51340), .B(n51341), .Z(n51046) );
  AND U51183 ( .A(n977), .B(n51342), .Z(n51341) );
  XOR U51184 ( .A(p_input[1188]), .B(p_input[1156]), .Z(n51342) );
  XOR U51185 ( .A(n51343), .B(n51344), .Z(n51334) );
  AND U51186 ( .A(n51345), .B(n51346), .Z(n51344) );
  XOR U51187 ( .A(n51343), .B(n51061), .Z(n51346) );
  XNOR U51188 ( .A(p_input[1219]), .B(n51347), .Z(n51061) );
  AND U51189 ( .A(n979), .B(n51348), .Z(n51347) );
  XOR U51190 ( .A(p_input[1251]), .B(p_input[1219]), .Z(n51348) );
  XNOR U51191 ( .A(n51058), .B(n51343), .Z(n51345) );
  XOR U51192 ( .A(n51349), .B(n51350), .Z(n51058) );
  AND U51193 ( .A(n977), .B(n51351), .Z(n51350) );
  XOR U51194 ( .A(p_input[1187]), .B(p_input[1155]), .Z(n51351) );
  XOR U51195 ( .A(n51352), .B(n51353), .Z(n51343) );
  AND U51196 ( .A(n51354), .B(n51355), .Z(n51353) );
  XOR U51197 ( .A(n51352), .B(n51073), .Z(n51355) );
  XNOR U51198 ( .A(p_input[1218]), .B(n51356), .Z(n51073) );
  AND U51199 ( .A(n979), .B(n51357), .Z(n51356) );
  XOR U51200 ( .A(p_input[1250]), .B(p_input[1218]), .Z(n51357) );
  XNOR U51201 ( .A(n51070), .B(n51352), .Z(n51354) );
  XOR U51202 ( .A(n51358), .B(n51359), .Z(n51070) );
  AND U51203 ( .A(n977), .B(n51360), .Z(n51359) );
  XOR U51204 ( .A(p_input[1186]), .B(p_input[1154]), .Z(n51360) );
  XOR U51205 ( .A(n51361), .B(n51362), .Z(n51352) );
  AND U51206 ( .A(n51363), .B(n51364), .Z(n51362) );
  XNOR U51207 ( .A(n51365), .B(n51086), .Z(n51364) );
  XNOR U51208 ( .A(p_input[1217]), .B(n51366), .Z(n51086) );
  AND U51209 ( .A(n979), .B(n51367), .Z(n51366) );
  XNOR U51210 ( .A(p_input[1249]), .B(n51368), .Z(n51367) );
  IV U51211 ( .A(p_input[1217]), .Z(n51368) );
  XNOR U51212 ( .A(n51083), .B(n51361), .Z(n51363) );
  XNOR U51213 ( .A(p_input[1153]), .B(n51369), .Z(n51083) );
  AND U51214 ( .A(n977), .B(n51370), .Z(n51369) );
  XOR U51215 ( .A(p_input[1185]), .B(p_input[1153]), .Z(n51370) );
  IV U51216 ( .A(n51365), .Z(n51361) );
  AND U51217 ( .A(n51091), .B(n51094), .Z(n51365) );
  XOR U51218 ( .A(p_input[1216]), .B(n51371), .Z(n51094) );
  AND U51219 ( .A(n979), .B(n51372), .Z(n51371) );
  XOR U51220 ( .A(p_input[1248]), .B(p_input[1216]), .Z(n51372) );
  XOR U51221 ( .A(n51373), .B(n51374), .Z(n979) );
  AND U51222 ( .A(n51375), .B(n51376), .Z(n51374) );
  XNOR U51223 ( .A(p_input[1279]), .B(n51373), .Z(n51376) );
  XOR U51224 ( .A(n51373), .B(p_input[1247]), .Z(n51375) );
  XOR U51225 ( .A(n51377), .B(n51378), .Z(n51373) );
  AND U51226 ( .A(n51379), .B(n51380), .Z(n51378) );
  XNOR U51227 ( .A(p_input[1278]), .B(n51377), .Z(n51380) );
  XOR U51228 ( .A(n51377), .B(p_input[1246]), .Z(n51379) );
  XOR U51229 ( .A(n51381), .B(n51382), .Z(n51377) );
  AND U51230 ( .A(n51383), .B(n51384), .Z(n51382) );
  XNOR U51231 ( .A(p_input[1277]), .B(n51381), .Z(n51384) );
  XOR U51232 ( .A(n51381), .B(p_input[1245]), .Z(n51383) );
  XOR U51233 ( .A(n51385), .B(n51386), .Z(n51381) );
  AND U51234 ( .A(n51387), .B(n51388), .Z(n51386) );
  XNOR U51235 ( .A(p_input[1276]), .B(n51385), .Z(n51388) );
  XOR U51236 ( .A(n51385), .B(p_input[1244]), .Z(n51387) );
  XOR U51237 ( .A(n51389), .B(n51390), .Z(n51385) );
  AND U51238 ( .A(n51391), .B(n51392), .Z(n51390) );
  XNOR U51239 ( .A(p_input[1275]), .B(n51389), .Z(n51392) );
  XOR U51240 ( .A(n51389), .B(p_input[1243]), .Z(n51391) );
  XOR U51241 ( .A(n51393), .B(n51394), .Z(n51389) );
  AND U51242 ( .A(n51395), .B(n51396), .Z(n51394) );
  XNOR U51243 ( .A(p_input[1274]), .B(n51393), .Z(n51396) );
  XOR U51244 ( .A(n51393), .B(p_input[1242]), .Z(n51395) );
  XOR U51245 ( .A(n51397), .B(n51398), .Z(n51393) );
  AND U51246 ( .A(n51399), .B(n51400), .Z(n51398) );
  XNOR U51247 ( .A(p_input[1273]), .B(n51397), .Z(n51400) );
  XOR U51248 ( .A(n51397), .B(p_input[1241]), .Z(n51399) );
  XOR U51249 ( .A(n51401), .B(n51402), .Z(n51397) );
  AND U51250 ( .A(n51403), .B(n51404), .Z(n51402) );
  XNOR U51251 ( .A(p_input[1272]), .B(n51401), .Z(n51404) );
  XOR U51252 ( .A(n51401), .B(p_input[1240]), .Z(n51403) );
  XOR U51253 ( .A(n51405), .B(n51406), .Z(n51401) );
  AND U51254 ( .A(n51407), .B(n51408), .Z(n51406) );
  XNOR U51255 ( .A(p_input[1271]), .B(n51405), .Z(n51408) );
  XOR U51256 ( .A(n51405), .B(p_input[1239]), .Z(n51407) );
  XOR U51257 ( .A(n51409), .B(n51410), .Z(n51405) );
  AND U51258 ( .A(n51411), .B(n51412), .Z(n51410) );
  XNOR U51259 ( .A(p_input[1270]), .B(n51409), .Z(n51412) );
  XOR U51260 ( .A(n51409), .B(p_input[1238]), .Z(n51411) );
  XOR U51261 ( .A(n51413), .B(n51414), .Z(n51409) );
  AND U51262 ( .A(n51415), .B(n51416), .Z(n51414) );
  XNOR U51263 ( .A(p_input[1269]), .B(n51413), .Z(n51416) );
  XOR U51264 ( .A(n51413), .B(p_input[1237]), .Z(n51415) );
  XOR U51265 ( .A(n51417), .B(n51418), .Z(n51413) );
  AND U51266 ( .A(n51419), .B(n51420), .Z(n51418) );
  XNOR U51267 ( .A(p_input[1268]), .B(n51417), .Z(n51420) );
  XOR U51268 ( .A(n51417), .B(p_input[1236]), .Z(n51419) );
  XOR U51269 ( .A(n51421), .B(n51422), .Z(n51417) );
  AND U51270 ( .A(n51423), .B(n51424), .Z(n51422) );
  XNOR U51271 ( .A(p_input[1267]), .B(n51421), .Z(n51424) );
  XOR U51272 ( .A(n51421), .B(p_input[1235]), .Z(n51423) );
  XOR U51273 ( .A(n51425), .B(n51426), .Z(n51421) );
  AND U51274 ( .A(n51427), .B(n51428), .Z(n51426) );
  XNOR U51275 ( .A(p_input[1266]), .B(n51425), .Z(n51428) );
  XOR U51276 ( .A(n51425), .B(p_input[1234]), .Z(n51427) );
  XOR U51277 ( .A(n51429), .B(n51430), .Z(n51425) );
  AND U51278 ( .A(n51431), .B(n51432), .Z(n51430) );
  XNOR U51279 ( .A(p_input[1265]), .B(n51429), .Z(n51432) );
  XOR U51280 ( .A(n51429), .B(p_input[1233]), .Z(n51431) );
  XOR U51281 ( .A(n51433), .B(n51434), .Z(n51429) );
  AND U51282 ( .A(n51435), .B(n51436), .Z(n51434) );
  XNOR U51283 ( .A(p_input[1264]), .B(n51433), .Z(n51436) );
  XOR U51284 ( .A(n51433), .B(p_input[1232]), .Z(n51435) );
  XOR U51285 ( .A(n51437), .B(n51438), .Z(n51433) );
  AND U51286 ( .A(n51439), .B(n51440), .Z(n51438) );
  XNOR U51287 ( .A(p_input[1263]), .B(n51437), .Z(n51440) );
  XOR U51288 ( .A(n51437), .B(p_input[1231]), .Z(n51439) );
  XOR U51289 ( .A(n51441), .B(n51442), .Z(n51437) );
  AND U51290 ( .A(n51443), .B(n51444), .Z(n51442) );
  XNOR U51291 ( .A(p_input[1262]), .B(n51441), .Z(n51444) );
  XOR U51292 ( .A(n51441), .B(p_input[1230]), .Z(n51443) );
  XOR U51293 ( .A(n51445), .B(n51446), .Z(n51441) );
  AND U51294 ( .A(n51447), .B(n51448), .Z(n51446) );
  XNOR U51295 ( .A(p_input[1261]), .B(n51445), .Z(n51448) );
  XOR U51296 ( .A(n51445), .B(p_input[1229]), .Z(n51447) );
  XOR U51297 ( .A(n51449), .B(n51450), .Z(n51445) );
  AND U51298 ( .A(n51451), .B(n51452), .Z(n51450) );
  XNOR U51299 ( .A(p_input[1260]), .B(n51449), .Z(n51452) );
  XOR U51300 ( .A(n51449), .B(p_input[1228]), .Z(n51451) );
  XOR U51301 ( .A(n51453), .B(n51454), .Z(n51449) );
  AND U51302 ( .A(n51455), .B(n51456), .Z(n51454) );
  XNOR U51303 ( .A(p_input[1259]), .B(n51453), .Z(n51456) );
  XOR U51304 ( .A(n51453), .B(p_input[1227]), .Z(n51455) );
  XOR U51305 ( .A(n51457), .B(n51458), .Z(n51453) );
  AND U51306 ( .A(n51459), .B(n51460), .Z(n51458) );
  XNOR U51307 ( .A(p_input[1258]), .B(n51457), .Z(n51460) );
  XOR U51308 ( .A(n51457), .B(p_input[1226]), .Z(n51459) );
  XOR U51309 ( .A(n51461), .B(n51462), .Z(n51457) );
  AND U51310 ( .A(n51463), .B(n51464), .Z(n51462) );
  XNOR U51311 ( .A(p_input[1257]), .B(n51461), .Z(n51464) );
  XOR U51312 ( .A(n51461), .B(p_input[1225]), .Z(n51463) );
  XOR U51313 ( .A(n51465), .B(n51466), .Z(n51461) );
  AND U51314 ( .A(n51467), .B(n51468), .Z(n51466) );
  XNOR U51315 ( .A(p_input[1256]), .B(n51465), .Z(n51468) );
  XOR U51316 ( .A(n51465), .B(p_input[1224]), .Z(n51467) );
  XOR U51317 ( .A(n51469), .B(n51470), .Z(n51465) );
  AND U51318 ( .A(n51471), .B(n51472), .Z(n51470) );
  XNOR U51319 ( .A(p_input[1255]), .B(n51469), .Z(n51472) );
  XOR U51320 ( .A(n51469), .B(p_input[1223]), .Z(n51471) );
  XOR U51321 ( .A(n51473), .B(n51474), .Z(n51469) );
  AND U51322 ( .A(n51475), .B(n51476), .Z(n51474) );
  XNOR U51323 ( .A(p_input[1254]), .B(n51473), .Z(n51476) );
  XOR U51324 ( .A(n51473), .B(p_input[1222]), .Z(n51475) );
  XOR U51325 ( .A(n51477), .B(n51478), .Z(n51473) );
  AND U51326 ( .A(n51479), .B(n51480), .Z(n51478) );
  XNOR U51327 ( .A(p_input[1253]), .B(n51477), .Z(n51480) );
  XOR U51328 ( .A(n51477), .B(p_input[1221]), .Z(n51479) );
  XOR U51329 ( .A(n51481), .B(n51482), .Z(n51477) );
  AND U51330 ( .A(n51483), .B(n51484), .Z(n51482) );
  XNOR U51331 ( .A(p_input[1252]), .B(n51481), .Z(n51484) );
  XOR U51332 ( .A(n51481), .B(p_input[1220]), .Z(n51483) );
  XOR U51333 ( .A(n51485), .B(n51486), .Z(n51481) );
  AND U51334 ( .A(n51487), .B(n51488), .Z(n51486) );
  XNOR U51335 ( .A(p_input[1251]), .B(n51485), .Z(n51488) );
  XOR U51336 ( .A(n51485), .B(p_input[1219]), .Z(n51487) );
  XOR U51337 ( .A(n51489), .B(n51490), .Z(n51485) );
  AND U51338 ( .A(n51491), .B(n51492), .Z(n51490) );
  XNOR U51339 ( .A(p_input[1250]), .B(n51489), .Z(n51492) );
  XOR U51340 ( .A(n51489), .B(p_input[1218]), .Z(n51491) );
  XNOR U51341 ( .A(n51493), .B(n51494), .Z(n51489) );
  AND U51342 ( .A(n51495), .B(n51496), .Z(n51494) );
  XOR U51343 ( .A(p_input[1249]), .B(n51493), .Z(n51496) );
  XNOR U51344 ( .A(p_input[1217]), .B(n51493), .Z(n51495) );
  AND U51345 ( .A(p_input[1248]), .B(n51497), .Z(n51493) );
  IV U51346 ( .A(p_input[1216]), .Z(n51497) );
  XNOR U51347 ( .A(p_input[1152]), .B(n51498), .Z(n51091) );
  AND U51348 ( .A(n977), .B(n51499), .Z(n51498) );
  XOR U51349 ( .A(p_input[1184]), .B(p_input[1152]), .Z(n51499) );
  XOR U51350 ( .A(n51500), .B(n51501), .Z(n977) );
  AND U51351 ( .A(n51502), .B(n51503), .Z(n51501) );
  XNOR U51352 ( .A(p_input[1215]), .B(n51500), .Z(n51503) );
  XOR U51353 ( .A(n51500), .B(p_input[1183]), .Z(n51502) );
  XOR U51354 ( .A(n51504), .B(n51505), .Z(n51500) );
  AND U51355 ( .A(n51506), .B(n51507), .Z(n51505) );
  XNOR U51356 ( .A(p_input[1214]), .B(n51504), .Z(n51507) );
  XNOR U51357 ( .A(n51504), .B(n51106), .Z(n51506) );
  IV U51358 ( .A(p_input[1182]), .Z(n51106) );
  XOR U51359 ( .A(n51508), .B(n51509), .Z(n51504) );
  AND U51360 ( .A(n51510), .B(n51511), .Z(n51509) );
  XNOR U51361 ( .A(p_input[1213]), .B(n51508), .Z(n51511) );
  XNOR U51362 ( .A(n51508), .B(n51115), .Z(n51510) );
  IV U51363 ( .A(p_input[1181]), .Z(n51115) );
  XOR U51364 ( .A(n51512), .B(n51513), .Z(n51508) );
  AND U51365 ( .A(n51514), .B(n51515), .Z(n51513) );
  XNOR U51366 ( .A(p_input[1212]), .B(n51512), .Z(n51515) );
  XNOR U51367 ( .A(n51512), .B(n51124), .Z(n51514) );
  IV U51368 ( .A(p_input[1180]), .Z(n51124) );
  XOR U51369 ( .A(n51516), .B(n51517), .Z(n51512) );
  AND U51370 ( .A(n51518), .B(n51519), .Z(n51517) );
  XNOR U51371 ( .A(p_input[1211]), .B(n51516), .Z(n51519) );
  XNOR U51372 ( .A(n51516), .B(n51133), .Z(n51518) );
  IV U51373 ( .A(p_input[1179]), .Z(n51133) );
  XOR U51374 ( .A(n51520), .B(n51521), .Z(n51516) );
  AND U51375 ( .A(n51522), .B(n51523), .Z(n51521) );
  XNOR U51376 ( .A(p_input[1210]), .B(n51520), .Z(n51523) );
  XNOR U51377 ( .A(n51520), .B(n51142), .Z(n51522) );
  IV U51378 ( .A(p_input[1178]), .Z(n51142) );
  XOR U51379 ( .A(n51524), .B(n51525), .Z(n51520) );
  AND U51380 ( .A(n51526), .B(n51527), .Z(n51525) );
  XNOR U51381 ( .A(p_input[1209]), .B(n51524), .Z(n51527) );
  XNOR U51382 ( .A(n51524), .B(n51151), .Z(n51526) );
  IV U51383 ( .A(p_input[1177]), .Z(n51151) );
  XOR U51384 ( .A(n51528), .B(n51529), .Z(n51524) );
  AND U51385 ( .A(n51530), .B(n51531), .Z(n51529) );
  XNOR U51386 ( .A(p_input[1208]), .B(n51528), .Z(n51531) );
  XNOR U51387 ( .A(n51528), .B(n51160), .Z(n51530) );
  IV U51388 ( .A(p_input[1176]), .Z(n51160) );
  XOR U51389 ( .A(n51532), .B(n51533), .Z(n51528) );
  AND U51390 ( .A(n51534), .B(n51535), .Z(n51533) );
  XNOR U51391 ( .A(p_input[1207]), .B(n51532), .Z(n51535) );
  XNOR U51392 ( .A(n51532), .B(n51169), .Z(n51534) );
  IV U51393 ( .A(p_input[1175]), .Z(n51169) );
  XOR U51394 ( .A(n51536), .B(n51537), .Z(n51532) );
  AND U51395 ( .A(n51538), .B(n51539), .Z(n51537) );
  XNOR U51396 ( .A(p_input[1206]), .B(n51536), .Z(n51539) );
  XNOR U51397 ( .A(n51536), .B(n51178), .Z(n51538) );
  IV U51398 ( .A(p_input[1174]), .Z(n51178) );
  XOR U51399 ( .A(n51540), .B(n51541), .Z(n51536) );
  AND U51400 ( .A(n51542), .B(n51543), .Z(n51541) );
  XNOR U51401 ( .A(p_input[1205]), .B(n51540), .Z(n51543) );
  XNOR U51402 ( .A(n51540), .B(n51187), .Z(n51542) );
  IV U51403 ( .A(p_input[1173]), .Z(n51187) );
  XOR U51404 ( .A(n51544), .B(n51545), .Z(n51540) );
  AND U51405 ( .A(n51546), .B(n51547), .Z(n51545) );
  XNOR U51406 ( .A(p_input[1204]), .B(n51544), .Z(n51547) );
  XNOR U51407 ( .A(n51544), .B(n51196), .Z(n51546) );
  IV U51408 ( .A(p_input[1172]), .Z(n51196) );
  XOR U51409 ( .A(n51548), .B(n51549), .Z(n51544) );
  AND U51410 ( .A(n51550), .B(n51551), .Z(n51549) );
  XNOR U51411 ( .A(p_input[1203]), .B(n51548), .Z(n51551) );
  XNOR U51412 ( .A(n51548), .B(n51205), .Z(n51550) );
  IV U51413 ( .A(p_input[1171]), .Z(n51205) );
  XOR U51414 ( .A(n51552), .B(n51553), .Z(n51548) );
  AND U51415 ( .A(n51554), .B(n51555), .Z(n51553) );
  XNOR U51416 ( .A(p_input[1202]), .B(n51552), .Z(n51555) );
  XNOR U51417 ( .A(n51552), .B(n51214), .Z(n51554) );
  IV U51418 ( .A(p_input[1170]), .Z(n51214) );
  XOR U51419 ( .A(n51556), .B(n51557), .Z(n51552) );
  AND U51420 ( .A(n51558), .B(n51559), .Z(n51557) );
  XNOR U51421 ( .A(p_input[1201]), .B(n51556), .Z(n51559) );
  XNOR U51422 ( .A(n51556), .B(n51223), .Z(n51558) );
  IV U51423 ( .A(p_input[1169]), .Z(n51223) );
  XOR U51424 ( .A(n51560), .B(n51561), .Z(n51556) );
  AND U51425 ( .A(n51562), .B(n51563), .Z(n51561) );
  XNOR U51426 ( .A(p_input[1200]), .B(n51560), .Z(n51563) );
  XNOR U51427 ( .A(n51560), .B(n51232), .Z(n51562) );
  IV U51428 ( .A(p_input[1168]), .Z(n51232) );
  XOR U51429 ( .A(n51564), .B(n51565), .Z(n51560) );
  AND U51430 ( .A(n51566), .B(n51567), .Z(n51565) );
  XNOR U51431 ( .A(p_input[1199]), .B(n51564), .Z(n51567) );
  XNOR U51432 ( .A(n51564), .B(n51241), .Z(n51566) );
  IV U51433 ( .A(p_input[1167]), .Z(n51241) );
  XOR U51434 ( .A(n51568), .B(n51569), .Z(n51564) );
  AND U51435 ( .A(n51570), .B(n51571), .Z(n51569) );
  XNOR U51436 ( .A(p_input[1198]), .B(n51568), .Z(n51571) );
  XNOR U51437 ( .A(n51568), .B(n51250), .Z(n51570) );
  IV U51438 ( .A(p_input[1166]), .Z(n51250) );
  XOR U51439 ( .A(n51572), .B(n51573), .Z(n51568) );
  AND U51440 ( .A(n51574), .B(n51575), .Z(n51573) );
  XNOR U51441 ( .A(p_input[1197]), .B(n51572), .Z(n51575) );
  XNOR U51442 ( .A(n51572), .B(n51259), .Z(n51574) );
  IV U51443 ( .A(p_input[1165]), .Z(n51259) );
  XOR U51444 ( .A(n51576), .B(n51577), .Z(n51572) );
  AND U51445 ( .A(n51578), .B(n51579), .Z(n51577) );
  XNOR U51446 ( .A(p_input[1196]), .B(n51576), .Z(n51579) );
  XNOR U51447 ( .A(n51576), .B(n51268), .Z(n51578) );
  IV U51448 ( .A(p_input[1164]), .Z(n51268) );
  XOR U51449 ( .A(n51580), .B(n51581), .Z(n51576) );
  AND U51450 ( .A(n51582), .B(n51583), .Z(n51581) );
  XNOR U51451 ( .A(p_input[1195]), .B(n51580), .Z(n51583) );
  XNOR U51452 ( .A(n51580), .B(n51277), .Z(n51582) );
  IV U51453 ( .A(p_input[1163]), .Z(n51277) );
  XOR U51454 ( .A(n51584), .B(n51585), .Z(n51580) );
  AND U51455 ( .A(n51586), .B(n51587), .Z(n51585) );
  XNOR U51456 ( .A(p_input[1194]), .B(n51584), .Z(n51587) );
  XNOR U51457 ( .A(n51584), .B(n51286), .Z(n51586) );
  IV U51458 ( .A(p_input[1162]), .Z(n51286) );
  XOR U51459 ( .A(n51588), .B(n51589), .Z(n51584) );
  AND U51460 ( .A(n51590), .B(n51591), .Z(n51589) );
  XNOR U51461 ( .A(p_input[1193]), .B(n51588), .Z(n51591) );
  XNOR U51462 ( .A(n51588), .B(n51295), .Z(n51590) );
  IV U51463 ( .A(p_input[1161]), .Z(n51295) );
  XOR U51464 ( .A(n51592), .B(n51593), .Z(n51588) );
  AND U51465 ( .A(n51594), .B(n51595), .Z(n51593) );
  XNOR U51466 ( .A(p_input[1192]), .B(n51592), .Z(n51595) );
  XNOR U51467 ( .A(n51592), .B(n51304), .Z(n51594) );
  IV U51468 ( .A(p_input[1160]), .Z(n51304) );
  XOR U51469 ( .A(n51596), .B(n51597), .Z(n51592) );
  AND U51470 ( .A(n51598), .B(n51599), .Z(n51597) );
  XNOR U51471 ( .A(p_input[1191]), .B(n51596), .Z(n51599) );
  XNOR U51472 ( .A(n51596), .B(n51313), .Z(n51598) );
  IV U51473 ( .A(p_input[1159]), .Z(n51313) );
  XOR U51474 ( .A(n51600), .B(n51601), .Z(n51596) );
  AND U51475 ( .A(n51602), .B(n51603), .Z(n51601) );
  XNOR U51476 ( .A(p_input[1190]), .B(n51600), .Z(n51603) );
  XNOR U51477 ( .A(n51600), .B(n51322), .Z(n51602) );
  IV U51478 ( .A(p_input[1158]), .Z(n51322) );
  XOR U51479 ( .A(n51604), .B(n51605), .Z(n51600) );
  AND U51480 ( .A(n51606), .B(n51607), .Z(n51605) );
  XNOR U51481 ( .A(p_input[1189]), .B(n51604), .Z(n51607) );
  XNOR U51482 ( .A(n51604), .B(n51331), .Z(n51606) );
  IV U51483 ( .A(p_input[1157]), .Z(n51331) );
  XOR U51484 ( .A(n51608), .B(n51609), .Z(n51604) );
  AND U51485 ( .A(n51610), .B(n51611), .Z(n51609) );
  XNOR U51486 ( .A(p_input[1188]), .B(n51608), .Z(n51611) );
  XNOR U51487 ( .A(n51608), .B(n51340), .Z(n51610) );
  IV U51488 ( .A(p_input[1156]), .Z(n51340) );
  XOR U51489 ( .A(n51612), .B(n51613), .Z(n51608) );
  AND U51490 ( .A(n51614), .B(n51615), .Z(n51613) );
  XNOR U51491 ( .A(p_input[1187]), .B(n51612), .Z(n51615) );
  XNOR U51492 ( .A(n51612), .B(n51349), .Z(n51614) );
  IV U51493 ( .A(p_input[1155]), .Z(n51349) );
  XOR U51494 ( .A(n51616), .B(n51617), .Z(n51612) );
  AND U51495 ( .A(n51618), .B(n51619), .Z(n51617) );
  XNOR U51496 ( .A(p_input[1186]), .B(n51616), .Z(n51619) );
  XNOR U51497 ( .A(n51616), .B(n51358), .Z(n51618) );
  IV U51498 ( .A(p_input[1154]), .Z(n51358) );
  XNOR U51499 ( .A(n51620), .B(n51621), .Z(n51616) );
  AND U51500 ( .A(n51622), .B(n51623), .Z(n51621) );
  XOR U51501 ( .A(p_input[1185]), .B(n51620), .Z(n51623) );
  XNOR U51502 ( .A(p_input[1153]), .B(n51620), .Z(n51622) );
  AND U51503 ( .A(p_input[1184]), .B(n51624), .Z(n51620) );
  IV U51504 ( .A(p_input[1152]), .Z(n51624) );
  XOR U51505 ( .A(n51625), .B(n51626), .Z(n50714) );
  AND U51506 ( .A(n636), .B(n51627), .Z(n51626) );
  XNOR U51507 ( .A(n51628), .B(n51625), .Z(n51627) );
  XOR U51508 ( .A(n51629), .B(n51630), .Z(n636) );
  AND U51509 ( .A(n51631), .B(n51632), .Z(n51630) );
  XNOR U51510 ( .A(n50729), .B(n51629), .Z(n51632) );
  AND U51511 ( .A(p_input[1151]), .B(p_input[1119]), .Z(n50729) );
  XNOR U51512 ( .A(n51629), .B(n50726), .Z(n51631) );
  IV U51513 ( .A(n51633), .Z(n50726) );
  AND U51514 ( .A(p_input[1055]), .B(p_input[1087]), .Z(n51633) );
  XOR U51515 ( .A(n51634), .B(n51635), .Z(n51629) );
  AND U51516 ( .A(n51636), .B(n51637), .Z(n51635) );
  XOR U51517 ( .A(n51634), .B(n50741), .Z(n51637) );
  XNOR U51518 ( .A(p_input[1118]), .B(n51638), .Z(n50741) );
  AND U51519 ( .A(n983), .B(n51639), .Z(n51638) );
  XOR U51520 ( .A(p_input[1150]), .B(p_input[1118]), .Z(n51639) );
  XNOR U51521 ( .A(n50738), .B(n51634), .Z(n51636) );
  XOR U51522 ( .A(n51640), .B(n51641), .Z(n50738) );
  AND U51523 ( .A(n980), .B(n51642), .Z(n51641) );
  XOR U51524 ( .A(p_input[1086]), .B(p_input[1054]), .Z(n51642) );
  XOR U51525 ( .A(n51643), .B(n51644), .Z(n51634) );
  AND U51526 ( .A(n51645), .B(n51646), .Z(n51644) );
  XOR U51527 ( .A(n51643), .B(n50753), .Z(n51646) );
  XNOR U51528 ( .A(p_input[1117]), .B(n51647), .Z(n50753) );
  AND U51529 ( .A(n983), .B(n51648), .Z(n51647) );
  XOR U51530 ( .A(p_input[1149]), .B(p_input[1117]), .Z(n51648) );
  XNOR U51531 ( .A(n50750), .B(n51643), .Z(n51645) );
  XOR U51532 ( .A(n51649), .B(n51650), .Z(n50750) );
  AND U51533 ( .A(n980), .B(n51651), .Z(n51650) );
  XOR U51534 ( .A(p_input[1085]), .B(p_input[1053]), .Z(n51651) );
  XOR U51535 ( .A(n51652), .B(n51653), .Z(n51643) );
  AND U51536 ( .A(n51654), .B(n51655), .Z(n51653) );
  XOR U51537 ( .A(n51652), .B(n50765), .Z(n51655) );
  XNOR U51538 ( .A(p_input[1116]), .B(n51656), .Z(n50765) );
  AND U51539 ( .A(n983), .B(n51657), .Z(n51656) );
  XOR U51540 ( .A(p_input[1148]), .B(p_input[1116]), .Z(n51657) );
  XNOR U51541 ( .A(n50762), .B(n51652), .Z(n51654) );
  XOR U51542 ( .A(n51658), .B(n51659), .Z(n50762) );
  AND U51543 ( .A(n980), .B(n51660), .Z(n51659) );
  XOR U51544 ( .A(p_input[1084]), .B(p_input[1052]), .Z(n51660) );
  XOR U51545 ( .A(n51661), .B(n51662), .Z(n51652) );
  AND U51546 ( .A(n51663), .B(n51664), .Z(n51662) );
  XOR U51547 ( .A(n51661), .B(n50777), .Z(n51664) );
  XNOR U51548 ( .A(p_input[1115]), .B(n51665), .Z(n50777) );
  AND U51549 ( .A(n983), .B(n51666), .Z(n51665) );
  XOR U51550 ( .A(p_input[1147]), .B(p_input[1115]), .Z(n51666) );
  XNOR U51551 ( .A(n50774), .B(n51661), .Z(n51663) );
  XOR U51552 ( .A(n51667), .B(n51668), .Z(n50774) );
  AND U51553 ( .A(n980), .B(n51669), .Z(n51668) );
  XOR U51554 ( .A(p_input[1083]), .B(p_input[1051]), .Z(n51669) );
  XOR U51555 ( .A(n51670), .B(n51671), .Z(n51661) );
  AND U51556 ( .A(n51672), .B(n51673), .Z(n51671) );
  XOR U51557 ( .A(n51670), .B(n50789), .Z(n51673) );
  XNOR U51558 ( .A(p_input[1114]), .B(n51674), .Z(n50789) );
  AND U51559 ( .A(n983), .B(n51675), .Z(n51674) );
  XOR U51560 ( .A(p_input[1146]), .B(p_input[1114]), .Z(n51675) );
  XNOR U51561 ( .A(n50786), .B(n51670), .Z(n51672) );
  XOR U51562 ( .A(n51676), .B(n51677), .Z(n50786) );
  AND U51563 ( .A(n980), .B(n51678), .Z(n51677) );
  XOR U51564 ( .A(p_input[1082]), .B(p_input[1050]), .Z(n51678) );
  XOR U51565 ( .A(n51679), .B(n51680), .Z(n51670) );
  AND U51566 ( .A(n51681), .B(n51682), .Z(n51680) );
  XOR U51567 ( .A(n51679), .B(n50801), .Z(n51682) );
  XNOR U51568 ( .A(p_input[1113]), .B(n51683), .Z(n50801) );
  AND U51569 ( .A(n983), .B(n51684), .Z(n51683) );
  XOR U51570 ( .A(p_input[1145]), .B(p_input[1113]), .Z(n51684) );
  XNOR U51571 ( .A(n50798), .B(n51679), .Z(n51681) );
  XOR U51572 ( .A(n51685), .B(n51686), .Z(n50798) );
  AND U51573 ( .A(n980), .B(n51687), .Z(n51686) );
  XOR U51574 ( .A(p_input[1081]), .B(p_input[1049]), .Z(n51687) );
  XOR U51575 ( .A(n51688), .B(n51689), .Z(n51679) );
  AND U51576 ( .A(n51690), .B(n51691), .Z(n51689) );
  XOR U51577 ( .A(n51688), .B(n50813), .Z(n51691) );
  XNOR U51578 ( .A(p_input[1112]), .B(n51692), .Z(n50813) );
  AND U51579 ( .A(n983), .B(n51693), .Z(n51692) );
  XOR U51580 ( .A(p_input[1144]), .B(p_input[1112]), .Z(n51693) );
  XNOR U51581 ( .A(n50810), .B(n51688), .Z(n51690) );
  XOR U51582 ( .A(n51694), .B(n51695), .Z(n50810) );
  AND U51583 ( .A(n980), .B(n51696), .Z(n51695) );
  XOR U51584 ( .A(p_input[1080]), .B(p_input[1048]), .Z(n51696) );
  XOR U51585 ( .A(n51697), .B(n51698), .Z(n51688) );
  AND U51586 ( .A(n51699), .B(n51700), .Z(n51698) );
  XOR U51587 ( .A(n51697), .B(n50825), .Z(n51700) );
  XNOR U51588 ( .A(p_input[1111]), .B(n51701), .Z(n50825) );
  AND U51589 ( .A(n983), .B(n51702), .Z(n51701) );
  XOR U51590 ( .A(p_input[1143]), .B(p_input[1111]), .Z(n51702) );
  XNOR U51591 ( .A(n50822), .B(n51697), .Z(n51699) );
  XOR U51592 ( .A(n51703), .B(n51704), .Z(n50822) );
  AND U51593 ( .A(n980), .B(n51705), .Z(n51704) );
  XOR U51594 ( .A(p_input[1079]), .B(p_input[1047]), .Z(n51705) );
  XOR U51595 ( .A(n51706), .B(n51707), .Z(n51697) );
  AND U51596 ( .A(n51708), .B(n51709), .Z(n51707) );
  XOR U51597 ( .A(n51706), .B(n50837), .Z(n51709) );
  XNOR U51598 ( .A(p_input[1110]), .B(n51710), .Z(n50837) );
  AND U51599 ( .A(n983), .B(n51711), .Z(n51710) );
  XOR U51600 ( .A(p_input[1142]), .B(p_input[1110]), .Z(n51711) );
  XNOR U51601 ( .A(n50834), .B(n51706), .Z(n51708) );
  XOR U51602 ( .A(n51712), .B(n51713), .Z(n50834) );
  AND U51603 ( .A(n980), .B(n51714), .Z(n51713) );
  XOR U51604 ( .A(p_input[1078]), .B(p_input[1046]), .Z(n51714) );
  XOR U51605 ( .A(n51715), .B(n51716), .Z(n51706) );
  AND U51606 ( .A(n51717), .B(n51718), .Z(n51716) );
  XOR U51607 ( .A(n51715), .B(n50849), .Z(n51718) );
  XNOR U51608 ( .A(p_input[1109]), .B(n51719), .Z(n50849) );
  AND U51609 ( .A(n983), .B(n51720), .Z(n51719) );
  XOR U51610 ( .A(p_input[1141]), .B(p_input[1109]), .Z(n51720) );
  XNOR U51611 ( .A(n50846), .B(n51715), .Z(n51717) );
  XOR U51612 ( .A(n51721), .B(n51722), .Z(n50846) );
  AND U51613 ( .A(n980), .B(n51723), .Z(n51722) );
  XOR U51614 ( .A(p_input[1077]), .B(p_input[1045]), .Z(n51723) );
  XOR U51615 ( .A(n51724), .B(n51725), .Z(n51715) );
  AND U51616 ( .A(n51726), .B(n51727), .Z(n51725) );
  XOR U51617 ( .A(n51724), .B(n50861), .Z(n51727) );
  XNOR U51618 ( .A(p_input[1108]), .B(n51728), .Z(n50861) );
  AND U51619 ( .A(n983), .B(n51729), .Z(n51728) );
  XOR U51620 ( .A(p_input[1140]), .B(p_input[1108]), .Z(n51729) );
  XNOR U51621 ( .A(n50858), .B(n51724), .Z(n51726) );
  XOR U51622 ( .A(n51730), .B(n51731), .Z(n50858) );
  AND U51623 ( .A(n980), .B(n51732), .Z(n51731) );
  XOR U51624 ( .A(p_input[1076]), .B(p_input[1044]), .Z(n51732) );
  XOR U51625 ( .A(n51733), .B(n51734), .Z(n51724) );
  AND U51626 ( .A(n51735), .B(n51736), .Z(n51734) );
  XOR U51627 ( .A(n51733), .B(n50873), .Z(n51736) );
  XNOR U51628 ( .A(p_input[1107]), .B(n51737), .Z(n50873) );
  AND U51629 ( .A(n983), .B(n51738), .Z(n51737) );
  XOR U51630 ( .A(p_input[1139]), .B(p_input[1107]), .Z(n51738) );
  XNOR U51631 ( .A(n50870), .B(n51733), .Z(n51735) );
  XOR U51632 ( .A(n51739), .B(n51740), .Z(n50870) );
  AND U51633 ( .A(n980), .B(n51741), .Z(n51740) );
  XOR U51634 ( .A(p_input[1075]), .B(p_input[1043]), .Z(n51741) );
  XOR U51635 ( .A(n51742), .B(n51743), .Z(n51733) );
  AND U51636 ( .A(n51744), .B(n51745), .Z(n51743) );
  XOR U51637 ( .A(n51742), .B(n50885), .Z(n51745) );
  XNOR U51638 ( .A(p_input[1106]), .B(n51746), .Z(n50885) );
  AND U51639 ( .A(n983), .B(n51747), .Z(n51746) );
  XOR U51640 ( .A(p_input[1138]), .B(p_input[1106]), .Z(n51747) );
  XNOR U51641 ( .A(n50882), .B(n51742), .Z(n51744) );
  XOR U51642 ( .A(n51748), .B(n51749), .Z(n50882) );
  AND U51643 ( .A(n980), .B(n51750), .Z(n51749) );
  XOR U51644 ( .A(p_input[1074]), .B(p_input[1042]), .Z(n51750) );
  XOR U51645 ( .A(n51751), .B(n51752), .Z(n51742) );
  AND U51646 ( .A(n51753), .B(n51754), .Z(n51752) );
  XOR U51647 ( .A(n51751), .B(n50897), .Z(n51754) );
  XNOR U51648 ( .A(p_input[1105]), .B(n51755), .Z(n50897) );
  AND U51649 ( .A(n983), .B(n51756), .Z(n51755) );
  XOR U51650 ( .A(p_input[1137]), .B(p_input[1105]), .Z(n51756) );
  XNOR U51651 ( .A(n50894), .B(n51751), .Z(n51753) );
  XOR U51652 ( .A(n51757), .B(n51758), .Z(n50894) );
  AND U51653 ( .A(n980), .B(n51759), .Z(n51758) );
  XOR U51654 ( .A(p_input[1073]), .B(p_input[1041]), .Z(n51759) );
  XOR U51655 ( .A(n51760), .B(n51761), .Z(n51751) );
  AND U51656 ( .A(n51762), .B(n51763), .Z(n51761) );
  XOR U51657 ( .A(n51760), .B(n50909), .Z(n51763) );
  XNOR U51658 ( .A(p_input[1104]), .B(n51764), .Z(n50909) );
  AND U51659 ( .A(n983), .B(n51765), .Z(n51764) );
  XOR U51660 ( .A(p_input[1136]), .B(p_input[1104]), .Z(n51765) );
  XNOR U51661 ( .A(n50906), .B(n51760), .Z(n51762) );
  XOR U51662 ( .A(n51766), .B(n51767), .Z(n50906) );
  AND U51663 ( .A(n980), .B(n51768), .Z(n51767) );
  XOR U51664 ( .A(p_input[1072]), .B(p_input[1040]), .Z(n51768) );
  XOR U51665 ( .A(n51769), .B(n51770), .Z(n51760) );
  AND U51666 ( .A(n51771), .B(n51772), .Z(n51770) );
  XOR U51667 ( .A(n51769), .B(n50921), .Z(n51772) );
  XNOR U51668 ( .A(p_input[1103]), .B(n51773), .Z(n50921) );
  AND U51669 ( .A(n983), .B(n51774), .Z(n51773) );
  XOR U51670 ( .A(p_input[1135]), .B(p_input[1103]), .Z(n51774) );
  XNOR U51671 ( .A(n50918), .B(n51769), .Z(n51771) );
  XOR U51672 ( .A(n51775), .B(n51776), .Z(n50918) );
  AND U51673 ( .A(n980), .B(n51777), .Z(n51776) );
  XOR U51674 ( .A(p_input[1071]), .B(p_input[1039]), .Z(n51777) );
  XOR U51675 ( .A(n51778), .B(n51779), .Z(n51769) );
  AND U51676 ( .A(n51780), .B(n51781), .Z(n51779) );
  XOR U51677 ( .A(n51778), .B(n50933), .Z(n51781) );
  XNOR U51678 ( .A(p_input[1102]), .B(n51782), .Z(n50933) );
  AND U51679 ( .A(n983), .B(n51783), .Z(n51782) );
  XOR U51680 ( .A(p_input[1134]), .B(p_input[1102]), .Z(n51783) );
  XNOR U51681 ( .A(n50930), .B(n51778), .Z(n51780) );
  XOR U51682 ( .A(n51784), .B(n51785), .Z(n50930) );
  AND U51683 ( .A(n980), .B(n51786), .Z(n51785) );
  XOR U51684 ( .A(p_input[1070]), .B(p_input[1038]), .Z(n51786) );
  XOR U51685 ( .A(n51787), .B(n51788), .Z(n51778) );
  AND U51686 ( .A(n51789), .B(n51790), .Z(n51788) );
  XOR U51687 ( .A(n51787), .B(n50945), .Z(n51790) );
  XNOR U51688 ( .A(p_input[1101]), .B(n51791), .Z(n50945) );
  AND U51689 ( .A(n983), .B(n51792), .Z(n51791) );
  XOR U51690 ( .A(p_input[1133]), .B(p_input[1101]), .Z(n51792) );
  XNOR U51691 ( .A(n50942), .B(n51787), .Z(n51789) );
  XOR U51692 ( .A(n51793), .B(n51794), .Z(n50942) );
  AND U51693 ( .A(n980), .B(n51795), .Z(n51794) );
  XOR U51694 ( .A(p_input[1069]), .B(p_input[1037]), .Z(n51795) );
  XOR U51695 ( .A(n51796), .B(n51797), .Z(n51787) );
  AND U51696 ( .A(n51798), .B(n51799), .Z(n51797) );
  XOR U51697 ( .A(n51796), .B(n50957), .Z(n51799) );
  XNOR U51698 ( .A(p_input[1100]), .B(n51800), .Z(n50957) );
  AND U51699 ( .A(n983), .B(n51801), .Z(n51800) );
  XOR U51700 ( .A(p_input[1132]), .B(p_input[1100]), .Z(n51801) );
  XNOR U51701 ( .A(n50954), .B(n51796), .Z(n51798) );
  XOR U51702 ( .A(n51802), .B(n51803), .Z(n50954) );
  AND U51703 ( .A(n980), .B(n51804), .Z(n51803) );
  XOR U51704 ( .A(p_input[1068]), .B(p_input[1036]), .Z(n51804) );
  XOR U51705 ( .A(n51805), .B(n51806), .Z(n51796) );
  AND U51706 ( .A(n51807), .B(n51808), .Z(n51806) );
  XOR U51707 ( .A(n51805), .B(n50969), .Z(n51808) );
  XNOR U51708 ( .A(p_input[1099]), .B(n51809), .Z(n50969) );
  AND U51709 ( .A(n983), .B(n51810), .Z(n51809) );
  XOR U51710 ( .A(p_input[1131]), .B(p_input[1099]), .Z(n51810) );
  XNOR U51711 ( .A(n50966), .B(n51805), .Z(n51807) );
  XOR U51712 ( .A(n51811), .B(n51812), .Z(n50966) );
  AND U51713 ( .A(n980), .B(n51813), .Z(n51812) );
  XOR U51714 ( .A(p_input[1067]), .B(p_input[1035]), .Z(n51813) );
  XOR U51715 ( .A(n51814), .B(n51815), .Z(n51805) );
  AND U51716 ( .A(n51816), .B(n51817), .Z(n51815) );
  XOR U51717 ( .A(n51814), .B(n50981), .Z(n51817) );
  XNOR U51718 ( .A(p_input[1098]), .B(n51818), .Z(n50981) );
  AND U51719 ( .A(n983), .B(n51819), .Z(n51818) );
  XOR U51720 ( .A(p_input[1130]), .B(p_input[1098]), .Z(n51819) );
  XNOR U51721 ( .A(n50978), .B(n51814), .Z(n51816) );
  XOR U51722 ( .A(n51820), .B(n51821), .Z(n50978) );
  AND U51723 ( .A(n980), .B(n51822), .Z(n51821) );
  XOR U51724 ( .A(p_input[1066]), .B(p_input[1034]), .Z(n51822) );
  XOR U51725 ( .A(n51823), .B(n51824), .Z(n51814) );
  AND U51726 ( .A(n51825), .B(n51826), .Z(n51824) );
  XOR U51727 ( .A(n51823), .B(n50993), .Z(n51826) );
  XNOR U51728 ( .A(p_input[1097]), .B(n51827), .Z(n50993) );
  AND U51729 ( .A(n983), .B(n51828), .Z(n51827) );
  XOR U51730 ( .A(p_input[1129]), .B(p_input[1097]), .Z(n51828) );
  XNOR U51731 ( .A(n50990), .B(n51823), .Z(n51825) );
  XOR U51732 ( .A(n51829), .B(n51830), .Z(n50990) );
  AND U51733 ( .A(n980), .B(n51831), .Z(n51830) );
  XOR U51734 ( .A(p_input[1065]), .B(p_input[1033]), .Z(n51831) );
  XOR U51735 ( .A(n51832), .B(n51833), .Z(n51823) );
  AND U51736 ( .A(n51834), .B(n51835), .Z(n51833) );
  XOR U51737 ( .A(n51832), .B(n51005), .Z(n51835) );
  XNOR U51738 ( .A(p_input[1096]), .B(n51836), .Z(n51005) );
  AND U51739 ( .A(n983), .B(n51837), .Z(n51836) );
  XOR U51740 ( .A(p_input[1128]), .B(p_input[1096]), .Z(n51837) );
  XNOR U51741 ( .A(n51002), .B(n51832), .Z(n51834) );
  XOR U51742 ( .A(n51838), .B(n51839), .Z(n51002) );
  AND U51743 ( .A(n980), .B(n51840), .Z(n51839) );
  XOR U51744 ( .A(p_input[1064]), .B(p_input[1032]), .Z(n51840) );
  XOR U51745 ( .A(n51841), .B(n51842), .Z(n51832) );
  AND U51746 ( .A(n51843), .B(n51844), .Z(n51842) );
  XOR U51747 ( .A(n51841), .B(n51017), .Z(n51844) );
  XNOR U51748 ( .A(p_input[1095]), .B(n51845), .Z(n51017) );
  AND U51749 ( .A(n983), .B(n51846), .Z(n51845) );
  XOR U51750 ( .A(p_input[1127]), .B(p_input[1095]), .Z(n51846) );
  XNOR U51751 ( .A(n51014), .B(n51841), .Z(n51843) );
  XOR U51752 ( .A(n51847), .B(n51848), .Z(n51014) );
  AND U51753 ( .A(n980), .B(n51849), .Z(n51848) );
  XOR U51754 ( .A(p_input[1063]), .B(p_input[1031]), .Z(n51849) );
  XOR U51755 ( .A(n51850), .B(n51851), .Z(n51841) );
  AND U51756 ( .A(n51852), .B(n51853), .Z(n51851) );
  XOR U51757 ( .A(n51850), .B(n51029), .Z(n51853) );
  XNOR U51758 ( .A(p_input[1094]), .B(n51854), .Z(n51029) );
  AND U51759 ( .A(n983), .B(n51855), .Z(n51854) );
  XOR U51760 ( .A(p_input[1126]), .B(p_input[1094]), .Z(n51855) );
  XNOR U51761 ( .A(n51026), .B(n51850), .Z(n51852) );
  XOR U51762 ( .A(n51856), .B(n51857), .Z(n51026) );
  AND U51763 ( .A(n980), .B(n51858), .Z(n51857) );
  XOR U51764 ( .A(p_input[1062]), .B(p_input[1030]), .Z(n51858) );
  XOR U51765 ( .A(n51859), .B(n51860), .Z(n51850) );
  AND U51766 ( .A(n51861), .B(n51862), .Z(n51860) );
  XOR U51767 ( .A(n51859), .B(n51041), .Z(n51862) );
  XNOR U51768 ( .A(p_input[1093]), .B(n51863), .Z(n51041) );
  AND U51769 ( .A(n983), .B(n51864), .Z(n51863) );
  XOR U51770 ( .A(p_input[1125]), .B(p_input[1093]), .Z(n51864) );
  XNOR U51771 ( .A(n51038), .B(n51859), .Z(n51861) );
  XOR U51772 ( .A(n51865), .B(n51866), .Z(n51038) );
  AND U51773 ( .A(n980), .B(n51867), .Z(n51866) );
  XOR U51774 ( .A(p_input[1061]), .B(p_input[1029]), .Z(n51867) );
  XOR U51775 ( .A(n51868), .B(n51869), .Z(n51859) );
  AND U51776 ( .A(n51870), .B(n51871), .Z(n51869) );
  XOR U51777 ( .A(n51868), .B(n51053), .Z(n51871) );
  XNOR U51778 ( .A(p_input[1092]), .B(n51872), .Z(n51053) );
  AND U51779 ( .A(n983), .B(n51873), .Z(n51872) );
  XOR U51780 ( .A(p_input[1124]), .B(p_input[1092]), .Z(n51873) );
  XNOR U51781 ( .A(n51050), .B(n51868), .Z(n51870) );
  XOR U51782 ( .A(n51874), .B(n51875), .Z(n51050) );
  AND U51783 ( .A(n980), .B(n51876), .Z(n51875) );
  XOR U51784 ( .A(p_input[1060]), .B(p_input[1028]), .Z(n51876) );
  XOR U51785 ( .A(n51877), .B(n51878), .Z(n51868) );
  AND U51786 ( .A(n51879), .B(n51880), .Z(n51878) );
  XOR U51787 ( .A(n51877), .B(n51065), .Z(n51880) );
  XNOR U51788 ( .A(p_input[1091]), .B(n51881), .Z(n51065) );
  AND U51789 ( .A(n983), .B(n51882), .Z(n51881) );
  XOR U51790 ( .A(p_input[1123]), .B(p_input[1091]), .Z(n51882) );
  XNOR U51791 ( .A(n51062), .B(n51877), .Z(n51879) );
  XOR U51792 ( .A(n51883), .B(n51884), .Z(n51062) );
  AND U51793 ( .A(n980), .B(n51885), .Z(n51884) );
  XOR U51794 ( .A(p_input[1059]), .B(p_input[1027]), .Z(n51885) );
  XOR U51795 ( .A(n51886), .B(n51887), .Z(n51877) );
  AND U51796 ( .A(n51888), .B(n51889), .Z(n51887) );
  XOR U51797 ( .A(n51886), .B(n51077), .Z(n51889) );
  XNOR U51798 ( .A(p_input[1090]), .B(n51890), .Z(n51077) );
  AND U51799 ( .A(n983), .B(n51891), .Z(n51890) );
  XOR U51800 ( .A(p_input[1122]), .B(p_input[1090]), .Z(n51891) );
  XNOR U51801 ( .A(n51074), .B(n51886), .Z(n51888) );
  XOR U51802 ( .A(n51892), .B(n51893), .Z(n51074) );
  AND U51803 ( .A(n980), .B(n51894), .Z(n51893) );
  XOR U51804 ( .A(p_input[1058]), .B(p_input[1026]), .Z(n51894) );
  XOR U51805 ( .A(n51895), .B(n51896), .Z(n51886) );
  AND U51806 ( .A(n51897), .B(n51898), .Z(n51896) );
  XNOR U51807 ( .A(n51899), .B(n51090), .Z(n51898) );
  XNOR U51808 ( .A(p_input[1089]), .B(n51900), .Z(n51090) );
  AND U51809 ( .A(n983), .B(n51901), .Z(n51900) );
  XNOR U51810 ( .A(p_input[1121]), .B(n51902), .Z(n51901) );
  IV U51811 ( .A(p_input[1089]), .Z(n51902) );
  XNOR U51812 ( .A(n51087), .B(n51895), .Z(n51897) );
  XNOR U51813 ( .A(p_input[1025]), .B(n51903), .Z(n51087) );
  AND U51814 ( .A(n980), .B(n51904), .Z(n51903) );
  XOR U51815 ( .A(p_input[1057]), .B(p_input[1025]), .Z(n51904) );
  IV U51816 ( .A(n51899), .Z(n51895) );
  AND U51817 ( .A(n51625), .B(n51628), .Z(n51899) );
  XOR U51818 ( .A(p_input[1088]), .B(n51905), .Z(n51628) );
  AND U51819 ( .A(n983), .B(n51906), .Z(n51905) );
  XOR U51820 ( .A(p_input[1120]), .B(p_input[1088]), .Z(n51906) );
  XOR U51821 ( .A(n51907), .B(n51908), .Z(n983) );
  AND U51822 ( .A(n51909), .B(n51910), .Z(n51908) );
  XNOR U51823 ( .A(p_input[1151]), .B(n51907), .Z(n51910) );
  XOR U51824 ( .A(n51907), .B(p_input[1119]), .Z(n51909) );
  XOR U51825 ( .A(n51911), .B(n51912), .Z(n51907) );
  AND U51826 ( .A(n51913), .B(n51914), .Z(n51912) );
  XNOR U51827 ( .A(p_input[1150]), .B(n51911), .Z(n51914) );
  XOR U51828 ( .A(n51911), .B(p_input[1118]), .Z(n51913) );
  XOR U51829 ( .A(n51915), .B(n51916), .Z(n51911) );
  AND U51830 ( .A(n51917), .B(n51918), .Z(n51916) );
  XNOR U51831 ( .A(p_input[1149]), .B(n51915), .Z(n51918) );
  XOR U51832 ( .A(n51915), .B(p_input[1117]), .Z(n51917) );
  XOR U51833 ( .A(n51919), .B(n51920), .Z(n51915) );
  AND U51834 ( .A(n51921), .B(n51922), .Z(n51920) );
  XNOR U51835 ( .A(p_input[1148]), .B(n51919), .Z(n51922) );
  XOR U51836 ( .A(n51919), .B(p_input[1116]), .Z(n51921) );
  XOR U51837 ( .A(n51923), .B(n51924), .Z(n51919) );
  AND U51838 ( .A(n51925), .B(n51926), .Z(n51924) );
  XNOR U51839 ( .A(p_input[1147]), .B(n51923), .Z(n51926) );
  XOR U51840 ( .A(n51923), .B(p_input[1115]), .Z(n51925) );
  XOR U51841 ( .A(n51927), .B(n51928), .Z(n51923) );
  AND U51842 ( .A(n51929), .B(n51930), .Z(n51928) );
  XNOR U51843 ( .A(p_input[1146]), .B(n51927), .Z(n51930) );
  XOR U51844 ( .A(n51927), .B(p_input[1114]), .Z(n51929) );
  XOR U51845 ( .A(n51931), .B(n51932), .Z(n51927) );
  AND U51846 ( .A(n51933), .B(n51934), .Z(n51932) );
  XNOR U51847 ( .A(p_input[1145]), .B(n51931), .Z(n51934) );
  XOR U51848 ( .A(n51931), .B(p_input[1113]), .Z(n51933) );
  XOR U51849 ( .A(n51935), .B(n51936), .Z(n51931) );
  AND U51850 ( .A(n51937), .B(n51938), .Z(n51936) );
  XNOR U51851 ( .A(p_input[1144]), .B(n51935), .Z(n51938) );
  XOR U51852 ( .A(n51935), .B(p_input[1112]), .Z(n51937) );
  XOR U51853 ( .A(n51939), .B(n51940), .Z(n51935) );
  AND U51854 ( .A(n51941), .B(n51942), .Z(n51940) );
  XNOR U51855 ( .A(p_input[1143]), .B(n51939), .Z(n51942) );
  XOR U51856 ( .A(n51939), .B(p_input[1111]), .Z(n51941) );
  XOR U51857 ( .A(n51943), .B(n51944), .Z(n51939) );
  AND U51858 ( .A(n51945), .B(n51946), .Z(n51944) );
  XNOR U51859 ( .A(p_input[1142]), .B(n51943), .Z(n51946) );
  XOR U51860 ( .A(n51943), .B(p_input[1110]), .Z(n51945) );
  XOR U51861 ( .A(n51947), .B(n51948), .Z(n51943) );
  AND U51862 ( .A(n51949), .B(n51950), .Z(n51948) );
  XNOR U51863 ( .A(p_input[1141]), .B(n51947), .Z(n51950) );
  XOR U51864 ( .A(n51947), .B(p_input[1109]), .Z(n51949) );
  XOR U51865 ( .A(n51951), .B(n51952), .Z(n51947) );
  AND U51866 ( .A(n51953), .B(n51954), .Z(n51952) );
  XNOR U51867 ( .A(p_input[1140]), .B(n51951), .Z(n51954) );
  XOR U51868 ( .A(n51951), .B(p_input[1108]), .Z(n51953) );
  XOR U51869 ( .A(n51955), .B(n51956), .Z(n51951) );
  AND U51870 ( .A(n51957), .B(n51958), .Z(n51956) );
  XNOR U51871 ( .A(p_input[1139]), .B(n51955), .Z(n51958) );
  XOR U51872 ( .A(n51955), .B(p_input[1107]), .Z(n51957) );
  XOR U51873 ( .A(n51959), .B(n51960), .Z(n51955) );
  AND U51874 ( .A(n51961), .B(n51962), .Z(n51960) );
  XNOR U51875 ( .A(p_input[1138]), .B(n51959), .Z(n51962) );
  XOR U51876 ( .A(n51959), .B(p_input[1106]), .Z(n51961) );
  XOR U51877 ( .A(n51963), .B(n51964), .Z(n51959) );
  AND U51878 ( .A(n51965), .B(n51966), .Z(n51964) );
  XNOR U51879 ( .A(p_input[1137]), .B(n51963), .Z(n51966) );
  XOR U51880 ( .A(n51963), .B(p_input[1105]), .Z(n51965) );
  XOR U51881 ( .A(n51967), .B(n51968), .Z(n51963) );
  AND U51882 ( .A(n51969), .B(n51970), .Z(n51968) );
  XNOR U51883 ( .A(p_input[1136]), .B(n51967), .Z(n51970) );
  XOR U51884 ( .A(n51967), .B(p_input[1104]), .Z(n51969) );
  XOR U51885 ( .A(n51971), .B(n51972), .Z(n51967) );
  AND U51886 ( .A(n51973), .B(n51974), .Z(n51972) );
  XNOR U51887 ( .A(p_input[1135]), .B(n51971), .Z(n51974) );
  XOR U51888 ( .A(n51971), .B(p_input[1103]), .Z(n51973) );
  XOR U51889 ( .A(n51975), .B(n51976), .Z(n51971) );
  AND U51890 ( .A(n51977), .B(n51978), .Z(n51976) );
  XNOR U51891 ( .A(p_input[1134]), .B(n51975), .Z(n51978) );
  XOR U51892 ( .A(n51975), .B(p_input[1102]), .Z(n51977) );
  XOR U51893 ( .A(n51979), .B(n51980), .Z(n51975) );
  AND U51894 ( .A(n51981), .B(n51982), .Z(n51980) );
  XNOR U51895 ( .A(p_input[1133]), .B(n51979), .Z(n51982) );
  XOR U51896 ( .A(n51979), .B(p_input[1101]), .Z(n51981) );
  XOR U51897 ( .A(n51983), .B(n51984), .Z(n51979) );
  AND U51898 ( .A(n51985), .B(n51986), .Z(n51984) );
  XNOR U51899 ( .A(p_input[1132]), .B(n51983), .Z(n51986) );
  XOR U51900 ( .A(n51983), .B(p_input[1100]), .Z(n51985) );
  XOR U51901 ( .A(n51987), .B(n51988), .Z(n51983) );
  AND U51902 ( .A(n51989), .B(n51990), .Z(n51988) );
  XNOR U51903 ( .A(p_input[1131]), .B(n51987), .Z(n51990) );
  XOR U51904 ( .A(n51987), .B(p_input[1099]), .Z(n51989) );
  XOR U51905 ( .A(n51991), .B(n51992), .Z(n51987) );
  AND U51906 ( .A(n51993), .B(n51994), .Z(n51992) );
  XNOR U51907 ( .A(p_input[1130]), .B(n51991), .Z(n51994) );
  XOR U51908 ( .A(n51991), .B(p_input[1098]), .Z(n51993) );
  XOR U51909 ( .A(n51995), .B(n51996), .Z(n51991) );
  AND U51910 ( .A(n51997), .B(n51998), .Z(n51996) );
  XNOR U51911 ( .A(p_input[1129]), .B(n51995), .Z(n51998) );
  XOR U51912 ( .A(n51995), .B(p_input[1097]), .Z(n51997) );
  XOR U51913 ( .A(n51999), .B(n52000), .Z(n51995) );
  AND U51914 ( .A(n52001), .B(n52002), .Z(n52000) );
  XNOR U51915 ( .A(p_input[1128]), .B(n51999), .Z(n52002) );
  XOR U51916 ( .A(n51999), .B(p_input[1096]), .Z(n52001) );
  XOR U51917 ( .A(n52003), .B(n52004), .Z(n51999) );
  AND U51918 ( .A(n52005), .B(n52006), .Z(n52004) );
  XNOR U51919 ( .A(p_input[1127]), .B(n52003), .Z(n52006) );
  XOR U51920 ( .A(n52003), .B(p_input[1095]), .Z(n52005) );
  XOR U51921 ( .A(n52007), .B(n52008), .Z(n52003) );
  AND U51922 ( .A(n52009), .B(n52010), .Z(n52008) );
  XNOR U51923 ( .A(p_input[1126]), .B(n52007), .Z(n52010) );
  XOR U51924 ( .A(n52007), .B(p_input[1094]), .Z(n52009) );
  XOR U51925 ( .A(n52011), .B(n52012), .Z(n52007) );
  AND U51926 ( .A(n52013), .B(n52014), .Z(n52012) );
  XNOR U51927 ( .A(p_input[1125]), .B(n52011), .Z(n52014) );
  XOR U51928 ( .A(n52011), .B(p_input[1093]), .Z(n52013) );
  XOR U51929 ( .A(n52015), .B(n52016), .Z(n52011) );
  AND U51930 ( .A(n52017), .B(n52018), .Z(n52016) );
  XNOR U51931 ( .A(p_input[1124]), .B(n52015), .Z(n52018) );
  XOR U51932 ( .A(n52015), .B(p_input[1092]), .Z(n52017) );
  XOR U51933 ( .A(n52019), .B(n52020), .Z(n52015) );
  AND U51934 ( .A(n52021), .B(n52022), .Z(n52020) );
  XNOR U51935 ( .A(p_input[1123]), .B(n52019), .Z(n52022) );
  XOR U51936 ( .A(n52019), .B(p_input[1091]), .Z(n52021) );
  XOR U51937 ( .A(n52023), .B(n52024), .Z(n52019) );
  AND U51938 ( .A(n52025), .B(n52026), .Z(n52024) );
  XNOR U51939 ( .A(p_input[1122]), .B(n52023), .Z(n52026) );
  XOR U51940 ( .A(n52023), .B(p_input[1090]), .Z(n52025) );
  XNOR U51941 ( .A(n52027), .B(n52028), .Z(n52023) );
  AND U51942 ( .A(n52029), .B(n52030), .Z(n52028) );
  XOR U51943 ( .A(p_input[1121]), .B(n52027), .Z(n52030) );
  XNOR U51944 ( .A(p_input[1089]), .B(n52027), .Z(n52029) );
  AND U51945 ( .A(p_input[1120]), .B(n52031), .Z(n52027) );
  IV U51946 ( .A(p_input[1088]), .Z(n52031) );
  XNOR U51947 ( .A(p_input[1024]), .B(n52032), .Z(n51625) );
  AND U51948 ( .A(n980), .B(n52033), .Z(n52032) );
  XOR U51949 ( .A(p_input[1056]), .B(p_input[1024]), .Z(n52033) );
  XOR U51950 ( .A(n52034), .B(n52035), .Z(n980) );
  AND U51951 ( .A(n52036), .B(n52037), .Z(n52035) );
  XNOR U51952 ( .A(p_input[1087]), .B(n52034), .Z(n52037) );
  XOR U51953 ( .A(n52034), .B(p_input[1055]), .Z(n52036) );
  XOR U51954 ( .A(n52038), .B(n52039), .Z(n52034) );
  AND U51955 ( .A(n52040), .B(n52041), .Z(n52039) );
  XNOR U51956 ( .A(p_input[1086]), .B(n52038), .Z(n52041) );
  XNOR U51957 ( .A(n52038), .B(n51640), .Z(n52040) );
  IV U51958 ( .A(p_input[1054]), .Z(n51640) );
  XOR U51959 ( .A(n52042), .B(n52043), .Z(n52038) );
  AND U51960 ( .A(n52044), .B(n52045), .Z(n52043) );
  XNOR U51961 ( .A(p_input[1085]), .B(n52042), .Z(n52045) );
  XNOR U51962 ( .A(n52042), .B(n51649), .Z(n52044) );
  IV U51963 ( .A(p_input[1053]), .Z(n51649) );
  XOR U51964 ( .A(n52046), .B(n52047), .Z(n52042) );
  AND U51965 ( .A(n52048), .B(n52049), .Z(n52047) );
  XNOR U51966 ( .A(p_input[1084]), .B(n52046), .Z(n52049) );
  XNOR U51967 ( .A(n52046), .B(n51658), .Z(n52048) );
  IV U51968 ( .A(p_input[1052]), .Z(n51658) );
  XOR U51969 ( .A(n52050), .B(n52051), .Z(n52046) );
  AND U51970 ( .A(n52052), .B(n52053), .Z(n52051) );
  XNOR U51971 ( .A(p_input[1083]), .B(n52050), .Z(n52053) );
  XNOR U51972 ( .A(n52050), .B(n51667), .Z(n52052) );
  IV U51973 ( .A(p_input[1051]), .Z(n51667) );
  XOR U51974 ( .A(n52054), .B(n52055), .Z(n52050) );
  AND U51975 ( .A(n52056), .B(n52057), .Z(n52055) );
  XNOR U51976 ( .A(p_input[1082]), .B(n52054), .Z(n52057) );
  XNOR U51977 ( .A(n52054), .B(n51676), .Z(n52056) );
  IV U51978 ( .A(p_input[1050]), .Z(n51676) );
  XOR U51979 ( .A(n52058), .B(n52059), .Z(n52054) );
  AND U51980 ( .A(n52060), .B(n52061), .Z(n52059) );
  XNOR U51981 ( .A(p_input[1081]), .B(n52058), .Z(n52061) );
  XNOR U51982 ( .A(n52058), .B(n51685), .Z(n52060) );
  IV U51983 ( .A(p_input[1049]), .Z(n51685) );
  XOR U51984 ( .A(n52062), .B(n52063), .Z(n52058) );
  AND U51985 ( .A(n52064), .B(n52065), .Z(n52063) );
  XNOR U51986 ( .A(p_input[1080]), .B(n52062), .Z(n52065) );
  XNOR U51987 ( .A(n52062), .B(n51694), .Z(n52064) );
  IV U51988 ( .A(p_input[1048]), .Z(n51694) );
  XOR U51989 ( .A(n52066), .B(n52067), .Z(n52062) );
  AND U51990 ( .A(n52068), .B(n52069), .Z(n52067) );
  XNOR U51991 ( .A(p_input[1079]), .B(n52066), .Z(n52069) );
  XNOR U51992 ( .A(n52066), .B(n51703), .Z(n52068) );
  IV U51993 ( .A(p_input[1047]), .Z(n51703) );
  XOR U51994 ( .A(n52070), .B(n52071), .Z(n52066) );
  AND U51995 ( .A(n52072), .B(n52073), .Z(n52071) );
  XNOR U51996 ( .A(p_input[1078]), .B(n52070), .Z(n52073) );
  XNOR U51997 ( .A(n52070), .B(n51712), .Z(n52072) );
  IV U51998 ( .A(p_input[1046]), .Z(n51712) );
  XOR U51999 ( .A(n52074), .B(n52075), .Z(n52070) );
  AND U52000 ( .A(n52076), .B(n52077), .Z(n52075) );
  XNOR U52001 ( .A(p_input[1077]), .B(n52074), .Z(n52077) );
  XNOR U52002 ( .A(n52074), .B(n51721), .Z(n52076) );
  IV U52003 ( .A(p_input[1045]), .Z(n51721) );
  XOR U52004 ( .A(n52078), .B(n52079), .Z(n52074) );
  AND U52005 ( .A(n52080), .B(n52081), .Z(n52079) );
  XNOR U52006 ( .A(p_input[1076]), .B(n52078), .Z(n52081) );
  XNOR U52007 ( .A(n52078), .B(n51730), .Z(n52080) );
  IV U52008 ( .A(p_input[1044]), .Z(n51730) );
  XOR U52009 ( .A(n52082), .B(n52083), .Z(n52078) );
  AND U52010 ( .A(n52084), .B(n52085), .Z(n52083) );
  XNOR U52011 ( .A(p_input[1075]), .B(n52082), .Z(n52085) );
  XNOR U52012 ( .A(n52082), .B(n51739), .Z(n52084) );
  IV U52013 ( .A(p_input[1043]), .Z(n51739) );
  XOR U52014 ( .A(n52086), .B(n52087), .Z(n52082) );
  AND U52015 ( .A(n52088), .B(n52089), .Z(n52087) );
  XNOR U52016 ( .A(p_input[1074]), .B(n52086), .Z(n52089) );
  XNOR U52017 ( .A(n52086), .B(n51748), .Z(n52088) );
  IV U52018 ( .A(p_input[1042]), .Z(n51748) );
  XOR U52019 ( .A(n52090), .B(n52091), .Z(n52086) );
  AND U52020 ( .A(n52092), .B(n52093), .Z(n52091) );
  XNOR U52021 ( .A(p_input[1073]), .B(n52090), .Z(n52093) );
  XNOR U52022 ( .A(n52090), .B(n51757), .Z(n52092) );
  IV U52023 ( .A(p_input[1041]), .Z(n51757) );
  XOR U52024 ( .A(n52094), .B(n52095), .Z(n52090) );
  AND U52025 ( .A(n52096), .B(n52097), .Z(n52095) );
  XNOR U52026 ( .A(p_input[1072]), .B(n52094), .Z(n52097) );
  XNOR U52027 ( .A(n52094), .B(n51766), .Z(n52096) );
  IV U52028 ( .A(p_input[1040]), .Z(n51766) );
  XOR U52029 ( .A(n52098), .B(n52099), .Z(n52094) );
  AND U52030 ( .A(n52100), .B(n52101), .Z(n52099) );
  XNOR U52031 ( .A(p_input[1071]), .B(n52098), .Z(n52101) );
  XNOR U52032 ( .A(n52098), .B(n51775), .Z(n52100) );
  IV U52033 ( .A(p_input[1039]), .Z(n51775) );
  XOR U52034 ( .A(n52102), .B(n52103), .Z(n52098) );
  AND U52035 ( .A(n52104), .B(n52105), .Z(n52103) );
  XNOR U52036 ( .A(p_input[1070]), .B(n52102), .Z(n52105) );
  XNOR U52037 ( .A(n52102), .B(n51784), .Z(n52104) );
  IV U52038 ( .A(p_input[1038]), .Z(n51784) );
  XOR U52039 ( .A(n52106), .B(n52107), .Z(n52102) );
  AND U52040 ( .A(n52108), .B(n52109), .Z(n52107) );
  XNOR U52041 ( .A(p_input[1069]), .B(n52106), .Z(n52109) );
  XNOR U52042 ( .A(n52106), .B(n51793), .Z(n52108) );
  IV U52043 ( .A(p_input[1037]), .Z(n51793) );
  XOR U52044 ( .A(n52110), .B(n52111), .Z(n52106) );
  AND U52045 ( .A(n52112), .B(n52113), .Z(n52111) );
  XNOR U52046 ( .A(p_input[1068]), .B(n52110), .Z(n52113) );
  XNOR U52047 ( .A(n52110), .B(n51802), .Z(n52112) );
  IV U52048 ( .A(p_input[1036]), .Z(n51802) );
  XOR U52049 ( .A(n52114), .B(n52115), .Z(n52110) );
  AND U52050 ( .A(n52116), .B(n52117), .Z(n52115) );
  XNOR U52051 ( .A(p_input[1067]), .B(n52114), .Z(n52117) );
  XNOR U52052 ( .A(n52114), .B(n51811), .Z(n52116) );
  IV U52053 ( .A(p_input[1035]), .Z(n51811) );
  XOR U52054 ( .A(n52118), .B(n52119), .Z(n52114) );
  AND U52055 ( .A(n52120), .B(n52121), .Z(n52119) );
  XNOR U52056 ( .A(p_input[1066]), .B(n52118), .Z(n52121) );
  XNOR U52057 ( .A(n52118), .B(n51820), .Z(n52120) );
  IV U52058 ( .A(p_input[1034]), .Z(n51820) );
  XOR U52059 ( .A(n52122), .B(n52123), .Z(n52118) );
  AND U52060 ( .A(n52124), .B(n52125), .Z(n52123) );
  XNOR U52061 ( .A(p_input[1065]), .B(n52122), .Z(n52125) );
  XNOR U52062 ( .A(n52122), .B(n51829), .Z(n52124) );
  IV U52063 ( .A(p_input[1033]), .Z(n51829) );
  XOR U52064 ( .A(n52126), .B(n52127), .Z(n52122) );
  AND U52065 ( .A(n52128), .B(n52129), .Z(n52127) );
  XNOR U52066 ( .A(p_input[1064]), .B(n52126), .Z(n52129) );
  XNOR U52067 ( .A(n52126), .B(n51838), .Z(n52128) );
  IV U52068 ( .A(p_input[1032]), .Z(n51838) );
  XOR U52069 ( .A(n52130), .B(n52131), .Z(n52126) );
  AND U52070 ( .A(n52132), .B(n52133), .Z(n52131) );
  XNOR U52071 ( .A(p_input[1063]), .B(n52130), .Z(n52133) );
  XNOR U52072 ( .A(n52130), .B(n51847), .Z(n52132) );
  IV U52073 ( .A(p_input[1031]), .Z(n51847) );
  XOR U52074 ( .A(n52134), .B(n52135), .Z(n52130) );
  AND U52075 ( .A(n52136), .B(n52137), .Z(n52135) );
  XNOR U52076 ( .A(p_input[1062]), .B(n52134), .Z(n52137) );
  XNOR U52077 ( .A(n52134), .B(n51856), .Z(n52136) );
  IV U52078 ( .A(p_input[1030]), .Z(n51856) );
  XOR U52079 ( .A(n52138), .B(n52139), .Z(n52134) );
  AND U52080 ( .A(n52140), .B(n52141), .Z(n52139) );
  XNOR U52081 ( .A(p_input[1061]), .B(n52138), .Z(n52141) );
  XNOR U52082 ( .A(n52138), .B(n51865), .Z(n52140) );
  IV U52083 ( .A(p_input[1029]), .Z(n51865) );
  XOR U52084 ( .A(n52142), .B(n52143), .Z(n52138) );
  AND U52085 ( .A(n52144), .B(n52145), .Z(n52143) );
  XNOR U52086 ( .A(p_input[1060]), .B(n52142), .Z(n52145) );
  XNOR U52087 ( .A(n52142), .B(n51874), .Z(n52144) );
  IV U52088 ( .A(p_input[1028]), .Z(n51874) );
  XOR U52089 ( .A(n52146), .B(n52147), .Z(n52142) );
  AND U52090 ( .A(n52148), .B(n52149), .Z(n52147) );
  XNOR U52091 ( .A(p_input[1059]), .B(n52146), .Z(n52149) );
  XNOR U52092 ( .A(n52146), .B(n51883), .Z(n52148) );
  IV U52093 ( .A(p_input[1027]), .Z(n51883) );
  XOR U52094 ( .A(n52150), .B(n52151), .Z(n52146) );
  AND U52095 ( .A(n52152), .B(n52153), .Z(n52151) );
  XNOR U52096 ( .A(p_input[1058]), .B(n52150), .Z(n52153) );
  XNOR U52097 ( .A(n52150), .B(n51892), .Z(n52152) );
  IV U52098 ( .A(p_input[1026]), .Z(n51892) );
  XNOR U52099 ( .A(n52154), .B(n52155), .Z(n52150) );
  AND U52100 ( .A(n52156), .B(n52157), .Z(n52155) );
  XOR U52101 ( .A(p_input[1057]), .B(n52154), .Z(n52157) );
  XNOR U52102 ( .A(p_input[1025]), .B(n52154), .Z(n52156) );
  AND U52103 ( .A(p_input[1056]), .B(n52158), .Z(n52154) );
  IV U52104 ( .A(p_input[1024]), .Z(n52158) );
  XOR U52105 ( .A(n52159), .B(n52160), .Z(n44871) );
  AND U52106 ( .A(n1100), .B(n52161), .Z(n52160) );
  XNOR U52107 ( .A(n52162), .B(n52159), .Z(n52161) );
  XOR U52108 ( .A(n52163), .B(n52164), .Z(n1100) );
  AND U52109 ( .A(n52165), .B(n52166), .Z(n52164) );
  XOR U52110 ( .A(n52163), .B(n44886), .Z(n52166) );
  XOR U52111 ( .A(n52167), .B(n52168), .Z(n44886) );
  AND U52112 ( .A(n1043), .B(n52169), .Z(n52168) );
  XOR U52113 ( .A(n52170), .B(n52167), .Z(n52169) );
  XNOR U52114 ( .A(n44883), .B(n52163), .Z(n52165) );
  XOR U52115 ( .A(n52171), .B(n52172), .Z(n44883) );
  AND U52116 ( .A(n1040), .B(n52173), .Z(n52172) );
  XOR U52117 ( .A(n52174), .B(n52171), .Z(n52173) );
  XOR U52118 ( .A(n52175), .B(n52176), .Z(n52163) );
  AND U52119 ( .A(n52177), .B(n52178), .Z(n52176) );
  XOR U52120 ( .A(n52175), .B(n44898), .Z(n52178) );
  XOR U52121 ( .A(n52179), .B(n52180), .Z(n44898) );
  AND U52122 ( .A(n1043), .B(n52181), .Z(n52180) );
  XOR U52123 ( .A(n52182), .B(n52179), .Z(n52181) );
  XNOR U52124 ( .A(n44895), .B(n52175), .Z(n52177) );
  XOR U52125 ( .A(n52183), .B(n52184), .Z(n44895) );
  AND U52126 ( .A(n1040), .B(n52185), .Z(n52184) );
  XOR U52127 ( .A(n52186), .B(n52183), .Z(n52185) );
  XOR U52128 ( .A(n52187), .B(n52188), .Z(n52175) );
  AND U52129 ( .A(n52189), .B(n52190), .Z(n52188) );
  XOR U52130 ( .A(n52187), .B(n44910), .Z(n52190) );
  XOR U52131 ( .A(n52191), .B(n52192), .Z(n44910) );
  AND U52132 ( .A(n1043), .B(n52193), .Z(n52192) );
  XOR U52133 ( .A(n52194), .B(n52191), .Z(n52193) );
  XNOR U52134 ( .A(n44907), .B(n52187), .Z(n52189) );
  XOR U52135 ( .A(n52195), .B(n52196), .Z(n44907) );
  AND U52136 ( .A(n1040), .B(n52197), .Z(n52196) );
  XOR U52137 ( .A(n52198), .B(n52195), .Z(n52197) );
  XOR U52138 ( .A(n52199), .B(n52200), .Z(n52187) );
  AND U52139 ( .A(n52201), .B(n52202), .Z(n52200) );
  XOR U52140 ( .A(n52199), .B(n44922), .Z(n52202) );
  XOR U52141 ( .A(n52203), .B(n52204), .Z(n44922) );
  AND U52142 ( .A(n1043), .B(n52205), .Z(n52204) );
  XOR U52143 ( .A(n52206), .B(n52203), .Z(n52205) );
  XNOR U52144 ( .A(n44919), .B(n52199), .Z(n52201) );
  XOR U52145 ( .A(n52207), .B(n52208), .Z(n44919) );
  AND U52146 ( .A(n1040), .B(n52209), .Z(n52208) );
  XOR U52147 ( .A(n52210), .B(n52207), .Z(n52209) );
  XOR U52148 ( .A(n52211), .B(n52212), .Z(n52199) );
  AND U52149 ( .A(n52213), .B(n52214), .Z(n52212) );
  XOR U52150 ( .A(n52211), .B(n44934), .Z(n52214) );
  XOR U52151 ( .A(n52215), .B(n52216), .Z(n44934) );
  AND U52152 ( .A(n1043), .B(n52217), .Z(n52216) );
  XOR U52153 ( .A(n52218), .B(n52215), .Z(n52217) );
  XNOR U52154 ( .A(n44931), .B(n52211), .Z(n52213) );
  XOR U52155 ( .A(n52219), .B(n52220), .Z(n44931) );
  AND U52156 ( .A(n1040), .B(n52221), .Z(n52220) );
  XOR U52157 ( .A(n52222), .B(n52219), .Z(n52221) );
  XOR U52158 ( .A(n52223), .B(n52224), .Z(n52211) );
  AND U52159 ( .A(n52225), .B(n52226), .Z(n52224) );
  XOR U52160 ( .A(n52223), .B(n44946), .Z(n52226) );
  XOR U52161 ( .A(n52227), .B(n52228), .Z(n44946) );
  AND U52162 ( .A(n1043), .B(n52229), .Z(n52228) );
  XOR U52163 ( .A(n52230), .B(n52227), .Z(n52229) );
  XNOR U52164 ( .A(n44943), .B(n52223), .Z(n52225) );
  XOR U52165 ( .A(n52231), .B(n52232), .Z(n44943) );
  AND U52166 ( .A(n1040), .B(n52233), .Z(n52232) );
  XOR U52167 ( .A(n52234), .B(n52231), .Z(n52233) );
  XOR U52168 ( .A(n52235), .B(n52236), .Z(n52223) );
  AND U52169 ( .A(n52237), .B(n52238), .Z(n52236) );
  XOR U52170 ( .A(n52235), .B(n44958), .Z(n52238) );
  XOR U52171 ( .A(n52239), .B(n52240), .Z(n44958) );
  AND U52172 ( .A(n1043), .B(n52241), .Z(n52240) );
  XOR U52173 ( .A(n52242), .B(n52239), .Z(n52241) );
  XNOR U52174 ( .A(n44955), .B(n52235), .Z(n52237) );
  XOR U52175 ( .A(n52243), .B(n52244), .Z(n44955) );
  AND U52176 ( .A(n1040), .B(n52245), .Z(n52244) );
  XOR U52177 ( .A(n52246), .B(n52243), .Z(n52245) );
  XOR U52178 ( .A(n52247), .B(n52248), .Z(n52235) );
  AND U52179 ( .A(n52249), .B(n52250), .Z(n52248) );
  XOR U52180 ( .A(n52247), .B(n44970), .Z(n52250) );
  XOR U52181 ( .A(n52251), .B(n52252), .Z(n44970) );
  AND U52182 ( .A(n1043), .B(n52253), .Z(n52252) );
  XOR U52183 ( .A(n52254), .B(n52251), .Z(n52253) );
  XNOR U52184 ( .A(n44967), .B(n52247), .Z(n52249) );
  XOR U52185 ( .A(n52255), .B(n52256), .Z(n44967) );
  AND U52186 ( .A(n1040), .B(n52257), .Z(n52256) );
  XOR U52187 ( .A(n52258), .B(n52255), .Z(n52257) );
  XOR U52188 ( .A(n52259), .B(n52260), .Z(n52247) );
  AND U52189 ( .A(n52261), .B(n52262), .Z(n52260) );
  XOR U52190 ( .A(n52259), .B(n44982), .Z(n52262) );
  XOR U52191 ( .A(n52263), .B(n52264), .Z(n44982) );
  AND U52192 ( .A(n1043), .B(n52265), .Z(n52264) );
  XOR U52193 ( .A(n52266), .B(n52263), .Z(n52265) );
  XNOR U52194 ( .A(n44979), .B(n52259), .Z(n52261) );
  XOR U52195 ( .A(n52267), .B(n52268), .Z(n44979) );
  AND U52196 ( .A(n1040), .B(n52269), .Z(n52268) );
  XOR U52197 ( .A(n52270), .B(n52267), .Z(n52269) );
  XOR U52198 ( .A(n52271), .B(n52272), .Z(n52259) );
  AND U52199 ( .A(n52273), .B(n52274), .Z(n52272) );
  XOR U52200 ( .A(n52271), .B(n44994), .Z(n52274) );
  XOR U52201 ( .A(n52275), .B(n52276), .Z(n44994) );
  AND U52202 ( .A(n1043), .B(n52277), .Z(n52276) );
  XOR U52203 ( .A(n52278), .B(n52275), .Z(n52277) );
  XNOR U52204 ( .A(n44991), .B(n52271), .Z(n52273) );
  XOR U52205 ( .A(n52279), .B(n52280), .Z(n44991) );
  AND U52206 ( .A(n1040), .B(n52281), .Z(n52280) );
  XOR U52207 ( .A(n52282), .B(n52279), .Z(n52281) );
  XOR U52208 ( .A(n52283), .B(n52284), .Z(n52271) );
  AND U52209 ( .A(n52285), .B(n52286), .Z(n52284) );
  XOR U52210 ( .A(n52283), .B(n45006), .Z(n52286) );
  XOR U52211 ( .A(n52287), .B(n52288), .Z(n45006) );
  AND U52212 ( .A(n1043), .B(n52289), .Z(n52288) );
  XOR U52213 ( .A(n52290), .B(n52287), .Z(n52289) );
  XNOR U52214 ( .A(n45003), .B(n52283), .Z(n52285) );
  XOR U52215 ( .A(n52291), .B(n52292), .Z(n45003) );
  AND U52216 ( .A(n1040), .B(n52293), .Z(n52292) );
  XOR U52217 ( .A(n52294), .B(n52291), .Z(n52293) );
  XOR U52218 ( .A(n52295), .B(n52296), .Z(n52283) );
  AND U52219 ( .A(n52297), .B(n52298), .Z(n52296) );
  XOR U52220 ( .A(n52295), .B(n45018), .Z(n52298) );
  XOR U52221 ( .A(n52299), .B(n52300), .Z(n45018) );
  AND U52222 ( .A(n1043), .B(n52301), .Z(n52300) );
  XOR U52223 ( .A(n52302), .B(n52299), .Z(n52301) );
  XNOR U52224 ( .A(n45015), .B(n52295), .Z(n52297) );
  XOR U52225 ( .A(n52303), .B(n52304), .Z(n45015) );
  AND U52226 ( .A(n1040), .B(n52305), .Z(n52304) );
  XOR U52227 ( .A(n52306), .B(n52303), .Z(n52305) );
  XOR U52228 ( .A(n52307), .B(n52308), .Z(n52295) );
  AND U52229 ( .A(n52309), .B(n52310), .Z(n52308) );
  XOR U52230 ( .A(n52307), .B(n45030), .Z(n52310) );
  XOR U52231 ( .A(n52311), .B(n52312), .Z(n45030) );
  AND U52232 ( .A(n1043), .B(n52313), .Z(n52312) );
  XOR U52233 ( .A(n52314), .B(n52311), .Z(n52313) );
  XNOR U52234 ( .A(n45027), .B(n52307), .Z(n52309) );
  XOR U52235 ( .A(n52315), .B(n52316), .Z(n45027) );
  AND U52236 ( .A(n1040), .B(n52317), .Z(n52316) );
  XOR U52237 ( .A(n52318), .B(n52315), .Z(n52317) );
  XOR U52238 ( .A(n52319), .B(n52320), .Z(n52307) );
  AND U52239 ( .A(n52321), .B(n52322), .Z(n52320) );
  XOR U52240 ( .A(n52319), .B(n45042), .Z(n52322) );
  XOR U52241 ( .A(n52323), .B(n52324), .Z(n45042) );
  AND U52242 ( .A(n1043), .B(n52325), .Z(n52324) );
  XOR U52243 ( .A(n52326), .B(n52323), .Z(n52325) );
  XNOR U52244 ( .A(n45039), .B(n52319), .Z(n52321) );
  XOR U52245 ( .A(n52327), .B(n52328), .Z(n45039) );
  AND U52246 ( .A(n1040), .B(n52329), .Z(n52328) );
  XOR U52247 ( .A(n52330), .B(n52327), .Z(n52329) );
  XOR U52248 ( .A(n52331), .B(n52332), .Z(n52319) );
  AND U52249 ( .A(n52333), .B(n52334), .Z(n52332) );
  XOR U52250 ( .A(n52331), .B(n45054), .Z(n52334) );
  XOR U52251 ( .A(n52335), .B(n52336), .Z(n45054) );
  AND U52252 ( .A(n1043), .B(n52337), .Z(n52336) );
  XOR U52253 ( .A(n52338), .B(n52335), .Z(n52337) );
  XNOR U52254 ( .A(n45051), .B(n52331), .Z(n52333) );
  XOR U52255 ( .A(n52339), .B(n52340), .Z(n45051) );
  AND U52256 ( .A(n1040), .B(n52341), .Z(n52340) );
  XOR U52257 ( .A(n52342), .B(n52339), .Z(n52341) );
  XOR U52258 ( .A(n52343), .B(n52344), .Z(n52331) );
  AND U52259 ( .A(n52345), .B(n52346), .Z(n52344) );
  XOR U52260 ( .A(n52343), .B(n45066), .Z(n52346) );
  XOR U52261 ( .A(n52347), .B(n52348), .Z(n45066) );
  AND U52262 ( .A(n1043), .B(n52349), .Z(n52348) );
  XOR U52263 ( .A(n52350), .B(n52347), .Z(n52349) );
  XNOR U52264 ( .A(n45063), .B(n52343), .Z(n52345) );
  XOR U52265 ( .A(n52351), .B(n52352), .Z(n45063) );
  AND U52266 ( .A(n1040), .B(n52353), .Z(n52352) );
  XOR U52267 ( .A(n52354), .B(n52351), .Z(n52353) );
  XOR U52268 ( .A(n52355), .B(n52356), .Z(n52343) );
  AND U52269 ( .A(n52357), .B(n52358), .Z(n52356) );
  XOR U52270 ( .A(n52355), .B(n45078), .Z(n52358) );
  XOR U52271 ( .A(n52359), .B(n52360), .Z(n45078) );
  AND U52272 ( .A(n1043), .B(n52361), .Z(n52360) );
  XOR U52273 ( .A(n52362), .B(n52359), .Z(n52361) );
  XNOR U52274 ( .A(n45075), .B(n52355), .Z(n52357) );
  XOR U52275 ( .A(n52363), .B(n52364), .Z(n45075) );
  AND U52276 ( .A(n1040), .B(n52365), .Z(n52364) );
  XOR U52277 ( .A(n52366), .B(n52363), .Z(n52365) );
  XOR U52278 ( .A(n52367), .B(n52368), .Z(n52355) );
  AND U52279 ( .A(n52369), .B(n52370), .Z(n52368) );
  XOR U52280 ( .A(n52367), .B(n45090), .Z(n52370) );
  XOR U52281 ( .A(n52371), .B(n52372), .Z(n45090) );
  AND U52282 ( .A(n1043), .B(n52373), .Z(n52372) );
  XOR U52283 ( .A(n52374), .B(n52371), .Z(n52373) );
  XNOR U52284 ( .A(n45087), .B(n52367), .Z(n52369) );
  XOR U52285 ( .A(n52375), .B(n52376), .Z(n45087) );
  AND U52286 ( .A(n1040), .B(n52377), .Z(n52376) );
  XOR U52287 ( .A(n52378), .B(n52375), .Z(n52377) );
  XOR U52288 ( .A(n52379), .B(n52380), .Z(n52367) );
  AND U52289 ( .A(n52381), .B(n52382), .Z(n52380) );
  XOR U52290 ( .A(n52379), .B(n45102), .Z(n52382) );
  XOR U52291 ( .A(n52383), .B(n52384), .Z(n45102) );
  AND U52292 ( .A(n1043), .B(n52385), .Z(n52384) );
  XOR U52293 ( .A(n52386), .B(n52383), .Z(n52385) );
  XNOR U52294 ( .A(n45099), .B(n52379), .Z(n52381) );
  XOR U52295 ( .A(n52387), .B(n52388), .Z(n45099) );
  AND U52296 ( .A(n1040), .B(n52389), .Z(n52388) );
  XOR U52297 ( .A(n52390), .B(n52387), .Z(n52389) );
  XOR U52298 ( .A(n52391), .B(n52392), .Z(n52379) );
  AND U52299 ( .A(n52393), .B(n52394), .Z(n52392) );
  XOR U52300 ( .A(n52391), .B(n45114), .Z(n52394) );
  XOR U52301 ( .A(n52395), .B(n52396), .Z(n45114) );
  AND U52302 ( .A(n1043), .B(n52397), .Z(n52396) );
  XOR U52303 ( .A(n52398), .B(n52395), .Z(n52397) );
  XNOR U52304 ( .A(n45111), .B(n52391), .Z(n52393) );
  XOR U52305 ( .A(n52399), .B(n52400), .Z(n45111) );
  AND U52306 ( .A(n1040), .B(n52401), .Z(n52400) );
  XOR U52307 ( .A(n52402), .B(n52399), .Z(n52401) );
  XOR U52308 ( .A(n52403), .B(n52404), .Z(n52391) );
  AND U52309 ( .A(n52405), .B(n52406), .Z(n52404) );
  XOR U52310 ( .A(n52403), .B(n45126), .Z(n52406) );
  XOR U52311 ( .A(n52407), .B(n52408), .Z(n45126) );
  AND U52312 ( .A(n1043), .B(n52409), .Z(n52408) );
  XOR U52313 ( .A(n52410), .B(n52407), .Z(n52409) );
  XNOR U52314 ( .A(n45123), .B(n52403), .Z(n52405) );
  XOR U52315 ( .A(n52411), .B(n52412), .Z(n45123) );
  AND U52316 ( .A(n1040), .B(n52413), .Z(n52412) );
  XOR U52317 ( .A(n52414), .B(n52411), .Z(n52413) );
  XOR U52318 ( .A(n52415), .B(n52416), .Z(n52403) );
  AND U52319 ( .A(n52417), .B(n52418), .Z(n52416) );
  XOR U52320 ( .A(n52415), .B(n45138), .Z(n52418) );
  XOR U52321 ( .A(n52419), .B(n52420), .Z(n45138) );
  AND U52322 ( .A(n1043), .B(n52421), .Z(n52420) );
  XOR U52323 ( .A(n52422), .B(n52419), .Z(n52421) );
  XNOR U52324 ( .A(n45135), .B(n52415), .Z(n52417) );
  XOR U52325 ( .A(n52423), .B(n52424), .Z(n45135) );
  AND U52326 ( .A(n1040), .B(n52425), .Z(n52424) );
  XOR U52327 ( .A(n52426), .B(n52423), .Z(n52425) );
  XOR U52328 ( .A(n52427), .B(n52428), .Z(n52415) );
  AND U52329 ( .A(n52429), .B(n52430), .Z(n52428) );
  XOR U52330 ( .A(n52427), .B(n45150), .Z(n52430) );
  XOR U52331 ( .A(n52431), .B(n52432), .Z(n45150) );
  AND U52332 ( .A(n1043), .B(n52433), .Z(n52432) );
  XOR U52333 ( .A(n52434), .B(n52431), .Z(n52433) );
  XNOR U52334 ( .A(n45147), .B(n52427), .Z(n52429) );
  XOR U52335 ( .A(n52435), .B(n52436), .Z(n45147) );
  AND U52336 ( .A(n1040), .B(n52437), .Z(n52436) );
  XOR U52337 ( .A(n52438), .B(n52435), .Z(n52437) );
  XOR U52338 ( .A(n52439), .B(n52440), .Z(n52427) );
  AND U52339 ( .A(n52441), .B(n52442), .Z(n52440) );
  XOR U52340 ( .A(n52439), .B(n45162), .Z(n52442) );
  XOR U52341 ( .A(n52443), .B(n52444), .Z(n45162) );
  AND U52342 ( .A(n1043), .B(n52445), .Z(n52444) );
  XOR U52343 ( .A(n52446), .B(n52443), .Z(n52445) );
  XNOR U52344 ( .A(n45159), .B(n52439), .Z(n52441) );
  XOR U52345 ( .A(n52447), .B(n52448), .Z(n45159) );
  AND U52346 ( .A(n1040), .B(n52449), .Z(n52448) );
  XOR U52347 ( .A(n52450), .B(n52447), .Z(n52449) );
  XOR U52348 ( .A(n52451), .B(n52452), .Z(n52439) );
  AND U52349 ( .A(n52453), .B(n52454), .Z(n52452) );
  XOR U52350 ( .A(n52451), .B(n45174), .Z(n52454) );
  XOR U52351 ( .A(n52455), .B(n52456), .Z(n45174) );
  AND U52352 ( .A(n1043), .B(n52457), .Z(n52456) );
  XOR U52353 ( .A(n52458), .B(n52455), .Z(n52457) );
  XNOR U52354 ( .A(n45171), .B(n52451), .Z(n52453) );
  XOR U52355 ( .A(n52459), .B(n52460), .Z(n45171) );
  AND U52356 ( .A(n1040), .B(n52461), .Z(n52460) );
  XOR U52357 ( .A(n52462), .B(n52459), .Z(n52461) );
  XOR U52358 ( .A(n52463), .B(n52464), .Z(n52451) );
  AND U52359 ( .A(n52465), .B(n52466), .Z(n52464) );
  XOR U52360 ( .A(n52463), .B(n45186), .Z(n52466) );
  XOR U52361 ( .A(n52467), .B(n52468), .Z(n45186) );
  AND U52362 ( .A(n1043), .B(n52469), .Z(n52468) );
  XOR U52363 ( .A(n52470), .B(n52467), .Z(n52469) );
  XNOR U52364 ( .A(n45183), .B(n52463), .Z(n52465) );
  XOR U52365 ( .A(n52471), .B(n52472), .Z(n45183) );
  AND U52366 ( .A(n1040), .B(n52473), .Z(n52472) );
  XOR U52367 ( .A(n52474), .B(n52471), .Z(n52473) );
  XOR U52368 ( .A(n52475), .B(n52476), .Z(n52463) );
  AND U52369 ( .A(n52477), .B(n52478), .Z(n52476) );
  XOR U52370 ( .A(n52475), .B(n45198), .Z(n52478) );
  XOR U52371 ( .A(n52479), .B(n52480), .Z(n45198) );
  AND U52372 ( .A(n1043), .B(n52481), .Z(n52480) );
  XOR U52373 ( .A(n52482), .B(n52479), .Z(n52481) );
  XNOR U52374 ( .A(n45195), .B(n52475), .Z(n52477) );
  XOR U52375 ( .A(n52483), .B(n52484), .Z(n45195) );
  AND U52376 ( .A(n1040), .B(n52485), .Z(n52484) );
  XOR U52377 ( .A(n52486), .B(n52483), .Z(n52485) );
  XOR U52378 ( .A(n52487), .B(n52488), .Z(n52475) );
  AND U52379 ( .A(n52489), .B(n52490), .Z(n52488) );
  XOR U52380 ( .A(n52487), .B(n45210), .Z(n52490) );
  XOR U52381 ( .A(n52491), .B(n52492), .Z(n45210) );
  AND U52382 ( .A(n1043), .B(n52493), .Z(n52492) );
  XOR U52383 ( .A(n52494), .B(n52491), .Z(n52493) );
  XNOR U52384 ( .A(n45207), .B(n52487), .Z(n52489) );
  XOR U52385 ( .A(n52495), .B(n52496), .Z(n45207) );
  AND U52386 ( .A(n1040), .B(n52497), .Z(n52496) );
  XOR U52387 ( .A(n52498), .B(n52495), .Z(n52497) );
  XOR U52388 ( .A(n52499), .B(n52500), .Z(n52487) );
  AND U52389 ( .A(n52501), .B(n52502), .Z(n52500) );
  XOR U52390 ( .A(n52499), .B(n45222), .Z(n52502) );
  XOR U52391 ( .A(n52503), .B(n52504), .Z(n45222) );
  AND U52392 ( .A(n1043), .B(n52505), .Z(n52504) );
  XOR U52393 ( .A(n52506), .B(n52503), .Z(n52505) );
  XNOR U52394 ( .A(n45219), .B(n52499), .Z(n52501) );
  XOR U52395 ( .A(n52507), .B(n52508), .Z(n45219) );
  AND U52396 ( .A(n1040), .B(n52509), .Z(n52508) );
  XOR U52397 ( .A(n52510), .B(n52507), .Z(n52509) );
  XOR U52398 ( .A(n52511), .B(n52512), .Z(n52499) );
  AND U52399 ( .A(n52513), .B(n52514), .Z(n52512) );
  XOR U52400 ( .A(n52511), .B(n45234), .Z(n52514) );
  XOR U52401 ( .A(n52515), .B(n52516), .Z(n45234) );
  AND U52402 ( .A(n1043), .B(n52517), .Z(n52516) );
  XOR U52403 ( .A(n52518), .B(n52515), .Z(n52517) );
  XNOR U52404 ( .A(n45231), .B(n52511), .Z(n52513) );
  XOR U52405 ( .A(n52519), .B(n52520), .Z(n45231) );
  AND U52406 ( .A(n1040), .B(n52521), .Z(n52520) );
  XOR U52407 ( .A(n52522), .B(n52519), .Z(n52521) );
  XOR U52408 ( .A(n52523), .B(n52524), .Z(n52511) );
  AND U52409 ( .A(n52525), .B(n52526), .Z(n52524) );
  XNOR U52410 ( .A(n52527), .B(n45247), .Z(n52526) );
  XOR U52411 ( .A(n52528), .B(n52529), .Z(n45247) );
  AND U52412 ( .A(n1043), .B(n52530), .Z(n52529) );
  XOR U52413 ( .A(n52528), .B(n52531), .Z(n52530) );
  XNOR U52414 ( .A(n45244), .B(n52523), .Z(n52525) );
  XOR U52415 ( .A(n52532), .B(n52533), .Z(n45244) );
  AND U52416 ( .A(n1040), .B(n52534), .Z(n52533) );
  XOR U52417 ( .A(n52532), .B(n52535), .Z(n52534) );
  IV U52418 ( .A(n52527), .Z(n52523) );
  AND U52419 ( .A(n52159), .B(n52162), .Z(n52527) );
  XNOR U52420 ( .A(n52536), .B(n52537), .Z(n52162) );
  AND U52421 ( .A(n1043), .B(n52538), .Z(n52537) );
  XNOR U52422 ( .A(n52539), .B(n52536), .Z(n52538) );
  XOR U52423 ( .A(n52540), .B(n52541), .Z(n1043) );
  AND U52424 ( .A(n52542), .B(n52543), .Z(n52541) );
  XOR U52425 ( .A(n52540), .B(n52170), .Z(n52543) );
  XOR U52426 ( .A(n52544), .B(n52545), .Z(n52170) );
  AND U52427 ( .A(n915), .B(n52546), .Z(n52545) );
  XOR U52428 ( .A(n52547), .B(n52544), .Z(n52546) );
  XNOR U52429 ( .A(n52167), .B(n52540), .Z(n52542) );
  XOR U52430 ( .A(n52548), .B(n52549), .Z(n52167) );
  AND U52431 ( .A(n913), .B(n52550), .Z(n52549) );
  XOR U52432 ( .A(n52551), .B(n52548), .Z(n52550) );
  XOR U52433 ( .A(n52552), .B(n52553), .Z(n52540) );
  AND U52434 ( .A(n52554), .B(n52555), .Z(n52553) );
  XOR U52435 ( .A(n52552), .B(n52182), .Z(n52555) );
  XOR U52436 ( .A(n52556), .B(n52557), .Z(n52182) );
  AND U52437 ( .A(n915), .B(n52558), .Z(n52557) );
  XOR U52438 ( .A(n52559), .B(n52556), .Z(n52558) );
  XNOR U52439 ( .A(n52179), .B(n52552), .Z(n52554) );
  XOR U52440 ( .A(n52560), .B(n52561), .Z(n52179) );
  AND U52441 ( .A(n913), .B(n52562), .Z(n52561) );
  XOR U52442 ( .A(n52563), .B(n52560), .Z(n52562) );
  XOR U52443 ( .A(n52564), .B(n52565), .Z(n52552) );
  AND U52444 ( .A(n52566), .B(n52567), .Z(n52565) );
  XOR U52445 ( .A(n52564), .B(n52194), .Z(n52567) );
  XOR U52446 ( .A(n52568), .B(n52569), .Z(n52194) );
  AND U52447 ( .A(n915), .B(n52570), .Z(n52569) );
  XOR U52448 ( .A(n52571), .B(n52568), .Z(n52570) );
  XNOR U52449 ( .A(n52191), .B(n52564), .Z(n52566) );
  XOR U52450 ( .A(n52572), .B(n52573), .Z(n52191) );
  AND U52451 ( .A(n913), .B(n52574), .Z(n52573) );
  XOR U52452 ( .A(n52575), .B(n52572), .Z(n52574) );
  XOR U52453 ( .A(n52576), .B(n52577), .Z(n52564) );
  AND U52454 ( .A(n52578), .B(n52579), .Z(n52577) );
  XOR U52455 ( .A(n52576), .B(n52206), .Z(n52579) );
  XOR U52456 ( .A(n52580), .B(n52581), .Z(n52206) );
  AND U52457 ( .A(n915), .B(n52582), .Z(n52581) );
  XOR U52458 ( .A(n52583), .B(n52580), .Z(n52582) );
  XNOR U52459 ( .A(n52203), .B(n52576), .Z(n52578) );
  XOR U52460 ( .A(n52584), .B(n52585), .Z(n52203) );
  AND U52461 ( .A(n913), .B(n52586), .Z(n52585) );
  XOR U52462 ( .A(n52587), .B(n52584), .Z(n52586) );
  XOR U52463 ( .A(n52588), .B(n52589), .Z(n52576) );
  AND U52464 ( .A(n52590), .B(n52591), .Z(n52589) );
  XOR U52465 ( .A(n52588), .B(n52218), .Z(n52591) );
  XOR U52466 ( .A(n52592), .B(n52593), .Z(n52218) );
  AND U52467 ( .A(n915), .B(n52594), .Z(n52593) );
  XOR U52468 ( .A(n52595), .B(n52592), .Z(n52594) );
  XNOR U52469 ( .A(n52215), .B(n52588), .Z(n52590) );
  XOR U52470 ( .A(n52596), .B(n52597), .Z(n52215) );
  AND U52471 ( .A(n913), .B(n52598), .Z(n52597) );
  XOR U52472 ( .A(n52599), .B(n52596), .Z(n52598) );
  XOR U52473 ( .A(n52600), .B(n52601), .Z(n52588) );
  AND U52474 ( .A(n52602), .B(n52603), .Z(n52601) );
  XOR U52475 ( .A(n52600), .B(n52230), .Z(n52603) );
  XOR U52476 ( .A(n52604), .B(n52605), .Z(n52230) );
  AND U52477 ( .A(n915), .B(n52606), .Z(n52605) );
  XOR U52478 ( .A(n52607), .B(n52604), .Z(n52606) );
  XNOR U52479 ( .A(n52227), .B(n52600), .Z(n52602) );
  XOR U52480 ( .A(n52608), .B(n52609), .Z(n52227) );
  AND U52481 ( .A(n913), .B(n52610), .Z(n52609) );
  XOR U52482 ( .A(n52611), .B(n52608), .Z(n52610) );
  XOR U52483 ( .A(n52612), .B(n52613), .Z(n52600) );
  AND U52484 ( .A(n52614), .B(n52615), .Z(n52613) );
  XOR U52485 ( .A(n52612), .B(n52242), .Z(n52615) );
  XOR U52486 ( .A(n52616), .B(n52617), .Z(n52242) );
  AND U52487 ( .A(n915), .B(n52618), .Z(n52617) );
  XOR U52488 ( .A(n52619), .B(n52616), .Z(n52618) );
  XNOR U52489 ( .A(n52239), .B(n52612), .Z(n52614) );
  XOR U52490 ( .A(n52620), .B(n52621), .Z(n52239) );
  AND U52491 ( .A(n913), .B(n52622), .Z(n52621) );
  XOR U52492 ( .A(n52623), .B(n52620), .Z(n52622) );
  XOR U52493 ( .A(n52624), .B(n52625), .Z(n52612) );
  AND U52494 ( .A(n52626), .B(n52627), .Z(n52625) );
  XOR U52495 ( .A(n52624), .B(n52254), .Z(n52627) );
  XOR U52496 ( .A(n52628), .B(n52629), .Z(n52254) );
  AND U52497 ( .A(n915), .B(n52630), .Z(n52629) );
  XOR U52498 ( .A(n52631), .B(n52628), .Z(n52630) );
  XNOR U52499 ( .A(n52251), .B(n52624), .Z(n52626) );
  XOR U52500 ( .A(n52632), .B(n52633), .Z(n52251) );
  AND U52501 ( .A(n913), .B(n52634), .Z(n52633) );
  XOR U52502 ( .A(n52635), .B(n52632), .Z(n52634) );
  XOR U52503 ( .A(n52636), .B(n52637), .Z(n52624) );
  AND U52504 ( .A(n52638), .B(n52639), .Z(n52637) );
  XOR U52505 ( .A(n52636), .B(n52266), .Z(n52639) );
  XOR U52506 ( .A(n52640), .B(n52641), .Z(n52266) );
  AND U52507 ( .A(n915), .B(n52642), .Z(n52641) );
  XOR U52508 ( .A(n52643), .B(n52640), .Z(n52642) );
  XNOR U52509 ( .A(n52263), .B(n52636), .Z(n52638) );
  XOR U52510 ( .A(n52644), .B(n52645), .Z(n52263) );
  AND U52511 ( .A(n913), .B(n52646), .Z(n52645) );
  XOR U52512 ( .A(n52647), .B(n52644), .Z(n52646) );
  XOR U52513 ( .A(n52648), .B(n52649), .Z(n52636) );
  AND U52514 ( .A(n52650), .B(n52651), .Z(n52649) );
  XOR U52515 ( .A(n52648), .B(n52278), .Z(n52651) );
  XOR U52516 ( .A(n52652), .B(n52653), .Z(n52278) );
  AND U52517 ( .A(n915), .B(n52654), .Z(n52653) );
  XOR U52518 ( .A(n52655), .B(n52652), .Z(n52654) );
  XNOR U52519 ( .A(n52275), .B(n52648), .Z(n52650) );
  XOR U52520 ( .A(n52656), .B(n52657), .Z(n52275) );
  AND U52521 ( .A(n913), .B(n52658), .Z(n52657) );
  XOR U52522 ( .A(n52659), .B(n52656), .Z(n52658) );
  XOR U52523 ( .A(n52660), .B(n52661), .Z(n52648) );
  AND U52524 ( .A(n52662), .B(n52663), .Z(n52661) );
  XOR U52525 ( .A(n52660), .B(n52290), .Z(n52663) );
  XOR U52526 ( .A(n52664), .B(n52665), .Z(n52290) );
  AND U52527 ( .A(n915), .B(n52666), .Z(n52665) );
  XOR U52528 ( .A(n52667), .B(n52664), .Z(n52666) );
  XNOR U52529 ( .A(n52287), .B(n52660), .Z(n52662) );
  XOR U52530 ( .A(n52668), .B(n52669), .Z(n52287) );
  AND U52531 ( .A(n913), .B(n52670), .Z(n52669) );
  XOR U52532 ( .A(n52671), .B(n52668), .Z(n52670) );
  XOR U52533 ( .A(n52672), .B(n52673), .Z(n52660) );
  AND U52534 ( .A(n52674), .B(n52675), .Z(n52673) );
  XOR U52535 ( .A(n52672), .B(n52302), .Z(n52675) );
  XOR U52536 ( .A(n52676), .B(n52677), .Z(n52302) );
  AND U52537 ( .A(n915), .B(n52678), .Z(n52677) );
  XOR U52538 ( .A(n52679), .B(n52676), .Z(n52678) );
  XNOR U52539 ( .A(n52299), .B(n52672), .Z(n52674) );
  XOR U52540 ( .A(n52680), .B(n52681), .Z(n52299) );
  AND U52541 ( .A(n913), .B(n52682), .Z(n52681) );
  XOR U52542 ( .A(n52683), .B(n52680), .Z(n52682) );
  XOR U52543 ( .A(n52684), .B(n52685), .Z(n52672) );
  AND U52544 ( .A(n52686), .B(n52687), .Z(n52685) );
  XOR U52545 ( .A(n52684), .B(n52314), .Z(n52687) );
  XOR U52546 ( .A(n52688), .B(n52689), .Z(n52314) );
  AND U52547 ( .A(n915), .B(n52690), .Z(n52689) );
  XOR U52548 ( .A(n52691), .B(n52688), .Z(n52690) );
  XNOR U52549 ( .A(n52311), .B(n52684), .Z(n52686) );
  XOR U52550 ( .A(n52692), .B(n52693), .Z(n52311) );
  AND U52551 ( .A(n913), .B(n52694), .Z(n52693) );
  XOR U52552 ( .A(n52695), .B(n52692), .Z(n52694) );
  XOR U52553 ( .A(n52696), .B(n52697), .Z(n52684) );
  AND U52554 ( .A(n52698), .B(n52699), .Z(n52697) );
  XOR U52555 ( .A(n52696), .B(n52326), .Z(n52699) );
  XOR U52556 ( .A(n52700), .B(n52701), .Z(n52326) );
  AND U52557 ( .A(n915), .B(n52702), .Z(n52701) );
  XOR U52558 ( .A(n52703), .B(n52700), .Z(n52702) );
  XNOR U52559 ( .A(n52323), .B(n52696), .Z(n52698) );
  XOR U52560 ( .A(n52704), .B(n52705), .Z(n52323) );
  AND U52561 ( .A(n913), .B(n52706), .Z(n52705) );
  XOR U52562 ( .A(n52707), .B(n52704), .Z(n52706) );
  XOR U52563 ( .A(n52708), .B(n52709), .Z(n52696) );
  AND U52564 ( .A(n52710), .B(n52711), .Z(n52709) );
  XOR U52565 ( .A(n52708), .B(n52338), .Z(n52711) );
  XOR U52566 ( .A(n52712), .B(n52713), .Z(n52338) );
  AND U52567 ( .A(n915), .B(n52714), .Z(n52713) );
  XOR U52568 ( .A(n52715), .B(n52712), .Z(n52714) );
  XNOR U52569 ( .A(n52335), .B(n52708), .Z(n52710) );
  XOR U52570 ( .A(n52716), .B(n52717), .Z(n52335) );
  AND U52571 ( .A(n913), .B(n52718), .Z(n52717) );
  XOR U52572 ( .A(n52719), .B(n52716), .Z(n52718) );
  XOR U52573 ( .A(n52720), .B(n52721), .Z(n52708) );
  AND U52574 ( .A(n52722), .B(n52723), .Z(n52721) );
  XOR U52575 ( .A(n52720), .B(n52350), .Z(n52723) );
  XOR U52576 ( .A(n52724), .B(n52725), .Z(n52350) );
  AND U52577 ( .A(n915), .B(n52726), .Z(n52725) );
  XOR U52578 ( .A(n52727), .B(n52724), .Z(n52726) );
  XNOR U52579 ( .A(n52347), .B(n52720), .Z(n52722) );
  XOR U52580 ( .A(n52728), .B(n52729), .Z(n52347) );
  AND U52581 ( .A(n913), .B(n52730), .Z(n52729) );
  XOR U52582 ( .A(n52731), .B(n52728), .Z(n52730) );
  XOR U52583 ( .A(n52732), .B(n52733), .Z(n52720) );
  AND U52584 ( .A(n52734), .B(n52735), .Z(n52733) );
  XOR U52585 ( .A(n52732), .B(n52362), .Z(n52735) );
  XOR U52586 ( .A(n52736), .B(n52737), .Z(n52362) );
  AND U52587 ( .A(n915), .B(n52738), .Z(n52737) );
  XOR U52588 ( .A(n52739), .B(n52736), .Z(n52738) );
  XNOR U52589 ( .A(n52359), .B(n52732), .Z(n52734) );
  XOR U52590 ( .A(n52740), .B(n52741), .Z(n52359) );
  AND U52591 ( .A(n913), .B(n52742), .Z(n52741) );
  XOR U52592 ( .A(n52743), .B(n52740), .Z(n52742) );
  XOR U52593 ( .A(n52744), .B(n52745), .Z(n52732) );
  AND U52594 ( .A(n52746), .B(n52747), .Z(n52745) );
  XOR U52595 ( .A(n52744), .B(n52374), .Z(n52747) );
  XOR U52596 ( .A(n52748), .B(n52749), .Z(n52374) );
  AND U52597 ( .A(n915), .B(n52750), .Z(n52749) );
  XOR U52598 ( .A(n52751), .B(n52748), .Z(n52750) );
  XNOR U52599 ( .A(n52371), .B(n52744), .Z(n52746) );
  XOR U52600 ( .A(n52752), .B(n52753), .Z(n52371) );
  AND U52601 ( .A(n913), .B(n52754), .Z(n52753) );
  XOR U52602 ( .A(n52755), .B(n52752), .Z(n52754) );
  XOR U52603 ( .A(n52756), .B(n52757), .Z(n52744) );
  AND U52604 ( .A(n52758), .B(n52759), .Z(n52757) );
  XOR U52605 ( .A(n52756), .B(n52386), .Z(n52759) );
  XOR U52606 ( .A(n52760), .B(n52761), .Z(n52386) );
  AND U52607 ( .A(n915), .B(n52762), .Z(n52761) );
  XOR U52608 ( .A(n52763), .B(n52760), .Z(n52762) );
  XNOR U52609 ( .A(n52383), .B(n52756), .Z(n52758) );
  XOR U52610 ( .A(n52764), .B(n52765), .Z(n52383) );
  AND U52611 ( .A(n913), .B(n52766), .Z(n52765) );
  XOR U52612 ( .A(n52767), .B(n52764), .Z(n52766) );
  XOR U52613 ( .A(n52768), .B(n52769), .Z(n52756) );
  AND U52614 ( .A(n52770), .B(n52771), .Z(n52769) );
  XOR U52615 ( .A(n52768), .B(n52398), .Z(n52771) );
  XOR U52616 ( .A(n52772), .B(n52773), .Z(n52398) );
  AND U52617 ( .A(n915), .B(n52774), .Z(n52773) );
  XOR U52618 ( .A(n52775), .B(n52772), .Z(n52774) );
  XNOR U52619 ( .A(n52395), .B(n52768), .Z(n52770) );
  XOR U52620 ( .A(n52776), .B(n52777), .Z(n52395) );
  AND U52621 ( .A(n913), .B(n52778), .Z(n52777) );
  XOR U52622 ( .A(n52779), .B(n52776), .Z(n52778) );
  XOR U52623 ( .A(n52780), .B(n52781), .Z(n52768) );
  AND U52624 ( .A(n52782), .B(n52783), .Z(n52781) );
  XOR U52625 ( .A(n52780), .B(n52410), .Z(n52783) );
  XOR U52626 ( .A(n52784), .B(n52785), .Z(n52410) );
  AND U52627 ( .A(n915), .B(n52786), .Z(n52785) );
  XOR U52628 ( .A(n52787), .B(n52784), .Z(n52786) );
  XNOR U52629 ( .A(n52407), .B(n52780), .Z(n52782) );
  XOR U52630 ( .A(n52788), .B(n52789), .Z(n52407) );
  AND U52631 ( .A(n913), .B(n52790), .Z(n52789) );
  XOR U52632 ( .A(n52791), .B(n52788), .Z(n52790) );
  XOR U52633 ( .A(n52792), .B(n52793), .Z(n52780) );
  AND U52634 ( .A(n52794), .B(n52795), .Z(n52793) );
  XOR U52635 ( .A(n52792), .B(n52422), .Z(n52795) );
  XOR U52636 ( .A(n52796), .B(n52797), .Z(n52422) );
  AND U52637 ( .A(n915), .B(n52798), .Z(n52797) );
  XOR U52638 ( .A(n52799), .B(n52796), .Z(n52798) );
  XNOR U52639 ( .A(n52419), .B(n52792), .Z(n52794) );
  XOR U52640 ( .A(n52800), .B(n52801), .Z(n52419) );
  AND U52641 ( .A(n913), .B(n52802), .Z(n52801) );
  XOR U52642 ( .A(n52803), .B(n52800), .Z(n52802) );
  XOR U52643 ( .A(n52804), .B(n52805), .Z(n52792) );
  AND U52644 ( .A(n52806), .B(n52807), .Z(n52805) );
  XOR U52645 ( .A(n52804), .B(n52434), .Z(n52807) );
  XOR U52646 ( .A(n52808), .B(n52809), .Z(n52434) );
  AND U52647 ( .A(n915), .B(n52810), .Z(n52809) );
  XOR U52648 ( .A(n52811), .B(n52808), .Z(n52810) );
  XNOR U52649 ( .A(n52431), .B(n52804), .Z(n52806) );
  XOR U52650 ( .A(n52812), .B(n52813), .Z(n52431) );
  AND U52651 ( .A(n913), .B(n52814), .Z(n52813) );
  XOR U52652 ( .A(n52815), .B(n52812), .Z(n52814) );
  XOR U52653 ( .A(n52816), .B(n52817), .Z(n52804) );
  AND U52654 ( .A(n52818), .B(n52819), .Z(n52817) );
  XOR U52655 ( .A(n52816), .B(n52446), .Z(n52819) );
  XOR U52656 ( .A(n52820), .B(n52821), .Z(n52446) );
  AND U52657 ( .A(n915), .B(n52822), .Z(n52821) );
  XOR U52658 ( .A(n52823), .B(n52820), .Z(n52822) );
  XNOR U52659 ( .A(n52443), .B(n52816), .Z(n52818) );
  XOR U52660 ( .A(n52824), .B(n52825), .Z(n52443) );
  AND U52661 ( .A(n913), .B(n52826), .Z(n52825) );
  XOR U52662 ( .A(n52827), .B(n52824), .Z(n52826) );
  XOR U52663 ( .A(n52828), .B(n52829), .Z(n52816) );
  AND U52664 ( .A(n52830), .B(n52831), .Z(n52829) );
  XOR U52665 ( .A(n52828), .B(n52458), .Z(n52831) );
  XOR U52666 ( .A(n52832), .B(n52833), .Z(n52458) );
  AND U52667 ( .A(n915), .B(n52834), .Z(n52833) );
  XOR U52668 ( .A(n52835), .B(n52832), .Z(n52834) );
  XNOR U52669 ( .A(n52455), .B(n52828), .Z(n52830) );
  XOR U52670 ( .A(n52836), .B(n52837), .Z(n52455) );
  AND U52671 ( .A(n913), .B(n52838), .Z(n52837) );
  XOR U52672 ( .A(n52839), .B(n52836), .Z(n52838) );
  XOR U52673 ( .A(n52840), .B(n52841), .Z(n52828) );
  AND U52674 ( .A(n52842), .B(n52843), .Z(n52841) );
  XOR U52675 ( .A(n52840), .B(n52470), .Z(n52843) );
  XOR U52676 ( .A(n52844), .B(n52845), .Z(n52470) );
  AND U52677 ( .A(n915), .B(n52846), .Z(n52845) );
  XOR U52678 ( .A(n52847), .B(n52844), .Z(n52846) );
  XNOR U52679 ( .A(n52467), .B(n52840), .Z(n52842) );
  XOR U52680 ( .A(n52848), .B(n52849), .Z(n52467) );
  AND U52681 ( .A(n913), .B(n52850), .Z(n52849) );
  XOR U52682 ( .A(n52851), .B(n52848), .Z(n52850) );
  XOR U52683 ( .A(n52852), .B(n52853), .Z(n52840) );
  AND U52684 ( .A(n52854), .B(n52855), .Z(n52853) );
  XOR U52685 ( .A(n52852), .B(n52482), .Z(n52855) );
  XOR U52686 ( .A(n52856), .B(n52857), .Z(n52482) );
  AND U52687 ( .A(n915), .B(n52858), .Z(n52857) );
  XOR U52688 ( .A(n52859), .B(n52856), .Z(n52858) );
  XNOR U52689 ( .A(n52479), .B(n52852), .Z(n52854) );
  XOR U52690 ( .A(n52860), .B(n52861), .Z(n52479) );
  AND U52691 ( .A(n913), .B(n52862), .Z(n52861) );
  XOR U52692 ( .A(n52863), .B(n52860), .Z(n52862) );
  XOR U52693 ( .A(n52864), .B(n52865), .Z(n52852) );
  AND U52694 ( .A(n52866), .B(n52867), .Z(n52865) );
  XOR U52695 ( .A(n52864), .B(n52494), .Z(n52867) );
  XOR U52696 ( .A(n52868), .B(n52869), .Z(n52494) );
  AND U52697 ( .A(n915), .B(n52870), .Z(n52869) );
  XOR U52698 ( .A(n52871), .B(n52868), .Z(n52870) );
  XNOR U52699 ( .A(n52491), .B(n52864), .Z(n52866) );
  XOR U52700 ( .A(n52872), .B(n52873), .Z(n52491) );
  AND U52701 ( .A(n913), .B(n52874), .Z(n52873) );
  XOR U52702 ( .A(n52875), .B(n52872), .Z(n52874) );
  XOR U52703 ( .A(n52876), .B(n52877), .Z(n52864) );
  AND U52704 ( .A(n52878), .B(n52879), .Z(n52877) );
  XOR U52705 ( .A(n52876), .B(n52506), .Z(n52879) );
  XOR U52706 ( .A(n52880), .B(n52881), .Z(n52506) );
  AND U52707 ( .A(n915), .B(n52882), .Z(n52881) );
  XOR U52708 ( .A(n52883), .B(n52880), .Z(n52882) );
  XNOR U52709 ( .A(n52503), .B(n52876), .Z(n52878) );
  XOR U52710 ( .A(n52884), .B(n52885), .Z(n52503) );
  AND U52711 ( .A(n913), .B(n52886), .Z(n52885) );
  XOR U52712 ( .A(n52887), .B(n52884), .Z(n52886) );
  XOR U52713 ( .A(n52888), .B(n52889), .Z(n52876) );
  AND U52714 ( .A(n52890), .B(n52891), .Z(n52889) );
  XOR U52715 ( .A(n52888), .B(n52518), .Z(n52891) );
  XOR U52716 ( .A(n52892), .B(n52893), .Z(n52518) );
  AND U52717 ( .A(n915), .B(n52894), .Z(n52893) );
  XOR U52718 ( .A(n52895), .B(n52892), .Z(n52894) );
  XNOR U52719 ( .A(n52515), .B(n52888), .Z(n52890) );
  XOR U52720 ( .A(n52896), .B(n52897), .Z(n52515) );
  AND U52721 ( .A(n913), .B(n52898), .Z(n52897) );
  XOR U52722 ( .A(n52899), .B(n52896), .Z(n52898) );
  XOR U52723 ( .A(n52900), .B(n52901), .Z(n52888) );
  AND U52724 ( .A(n52902), .B(n52903), .Z(n52901) );
  XNOR U52725 ( .A(n52904), .B(n52531), .Z(n52903) );
  XOR U52726 ( .A(n52905), .B(n52906), .Z(n52531) );
  AND U52727 ( .A(n915), .B(n52907), .Z(n52906) );
  XOR U52728 ( .A(n52905), .B(n52908), .Z(n52907) );
  XNOR U52729 ( .A(n52528), .B(n52900), .Z(n52902) );
  XOR U52730 ( .A(n52909), .B(n52910), .Z(n52528) );
  AND U52731 ( .A(n913), .B(n52911), .Z(n52910) );
  XOR U52732 ( .A(n52909), .B(n52912), .Z(n52911) );
  IV U52733 ( .A(n52904), .Z(n52900) );
  AND U52734 ( .A(n52536), .B(n52539), .Z(n52904) );
  XNOR U52735 ( .A(n52913), .B(n52914), .Z(n52539) );
  AND U52736 ( .A(n915), .B(n52915), .Z(n52914) );
  XNOR U52737 ( .A(n52916), .B(n52913), .Z(n52915) );
  XOR U52738 ( .A(n52917), .B(n52918), .Z(n915) );
  AND U52739 ( .A(n52919), .B(n52920), .Z(n52918) );
  XOR U52740 ( .A(n52917), .B(n52547), .Z(n52920) );
  XNOR U52741 ( .A(n52921), .B(n52922), .Z(n52547) );
  AND U52742 ( .A(n52923), .B(n651), .Z(n52922) );
  AND U52743 ( .A(n52921), .B(n52924), .Z(n52923) );
  XNOR U52744 ( .A(n52544), .B(n52917), .Z(n52919) );
  XOR U52745 ( .A(n52925), .B(n52926), .Z(n52544) );
  AND U52746 ( .A(n52927), .B(n649), .Z(n52926) );
  NOR U52747 ( .A(n52925), .B(n52928), .Z(n52927) );
  XOR U52748 ( .A(n52929), .B(n52930), .Z(n52917) );
  AND U52749 ( .A(n52931), .B(n52932), .Z(n52930) );
  XOR U52750 ( .A(n52929), .B(n52559), .Z(n52932) );
  XOR U52751 ( .A(n52933), .B(n52934), .Z(n52559) );
  AND U52752 ( .A(n651), .B(n52935), .Z(n52934) );
  XOR U52753 ( .A(n52936), .B(n52933), .Z(n52935) );
  XNOR U52754 ( .A(n52556), .B(n52929), .Z(n52931) );
  XOR U52755 ( .A(n52937), .B(n52938), .Z(n52556) );
  AND U52756 ( .A(n649), .B(n52939), .Z(n52938) );
  XOR U52757 ( .A(n52940), .B(n52937), .Z(n52939) );
  XOR U52758 ( .A(n52941), .B(n52942), .Z(n52929) );
  AND U52759 ( .A(n52943), .B(n52944), .Z(n52942) );
  XOR U52760 ( .A(n52941), .B(n52571), .Z(n52944) );
  XOR U52761 ( .A(n52945), .B(n52946), .Z(n52571) );
  AND U52762 ( .A(n651), .B(n52947), .Z(n52946) );
  XOR U52763 ( .A(n52948), .B(n52945), .Z(n52947) );
  XNOR U52764 ( .A(n52568), .B(n52941), .Z(n52943) );
  XOR U52765 ( .A(n52949), .B(n52950), .Z(n52568) );
  AND U52766 ( .A(n649), .B(n52951), .Z(n52950) );
  XOR U52767 ( .A(n52952), .B(n52949), .Z(n52951) );
  XOR U52768 ( .A(n52953), .B(n52954), .Z(n52941) );
  AND U52769 ( .A(n52955), .B(n52956), .Z(n52954) );
  XOR U52770 ( .A(n52953), .B(n52583), .Z(n52956) );
  XOR U52771 ( .A(n52957), .B(n52958), .Z(n52583) );
  AND U52772 ( .A(n651), .B(n52959), .Z(n52958) );
  XOR U52773 ( .A(n52960), .B(n52957), .Z(n52959) );
  XNOR U52774 ( .A(n52580), .B(n52953), .Z(n52955) );
  XOR U52775 ( .A(n52961), .B(n52962), .Z(n52580) );
  AND U52776 ( .A(n649), .B(n52963), .Z(n52962) );
  XOR U52777 ( .A(n52964), .B(n52961), .Z(n52963) );
  XOR U52778 ( .A(n52965), .B(n52966), .Z(n52953) );
  AND U52779 ( .A(n52967), .B(n52968), .Z(n52966) );
  XOR U52780 ( .A(n52965), .B(n52595), .Z(n52968) );
  XOR U52781 ( .A(n52969), .B(n52970), .Z(n52595) );
  AND U52782 ( .A(n651), .B(n52971), .Z(n52970) );
  XOR U52783 ( .A(n52972), .B(n52969), .Z(n52971) );
  XNOR U52784 ( .A(n52592), .B(n52965), .Z(n52967) );
  XOR U52785 ( .A(n52973), .B(n52974), .Z(n52592) );
  AND U52786 ( .A(n649), .B(n52975), .Z(n52974) );
  XOR U52787 ( .A(n52976), .B(n52973), .Z(n52975) );
  XOR U52788 ( .A(n52977), .B(n52978), .Z(n52965) );
  AND U52789 ( .A(n52979), .B(n52980), .Z(n52978) );
  XOR U52790 ( .A(n52977), .B(n52607), .Z(n52980) );
  XOR U52791 ( .A(n52981), .B(n52982), .Z(n52607) );
  AND U52792 ( .A(n651), .B(n52983), .Z(n52982) );
  XOR U52793 ( .A(n52984), .B(n52981), .Z(n52983) );
  XNOR U52794 ( .A(n52604), .B(n52977), .Z(n52979) );
  XOR U52795 ( .A(n52985), .B(n52986), .Z(n52604) );
  AND U52796 ( .A(n649), .B(n52987), .Z(n52986) );
  XOR U52797 ( .A(n52988), .B(n52985), .Z(n52987) );
  XOR U52798 ( .A(n52989), .B(n52990), .Z(n52977) );
  AND U52799 ( .A(n52991), .B(n52992), .Z(n52990) );
  XOR U52800 ( .A(n52989), .B(n52619), .Z(n52992) );
  XOR U52801 ( .A(n52993), .B(n52994), .Z(n52619) );
  AND U52802 ( .A(n651), .B(n52995), .Z(n52994) );
  XOR U52803 ( .A(n52996), .B(n52993), .Z(n52995) );
  XNOR U52804 ( .A(n52616), .B(n52989), .Z(n52991) );
  XOR U52805 ( .A(n52997), .B(n52998), .Z(n52616) );
  AND U52806 ( .A(n649), .B(n52999), .Z(n52998) );
  XOR U52807 ( .A(n53000), .B(n52997), .Z(n52999) );
  XOR U52808 ( .A(n53001), .B(n53002), .Z(n52989) );
  AND U52809 ( .A(n53003), .B(n53004), .Z(n53002) );
  XOR U52810 ( .A(n53001), .B(n52631), .Z(n53004) );
  XOR U52811 ( .A(n53005), .B(n53006), .Z(n52631) );
  AND U52812 ( .A(n651), .B(n53007), .Z(n53006) );
  XOR U52813 ( .A(n53008), .B(n53005), .Z(n53007) );
  XNOR U52814 ( .A(n52628), .B(n53001), .Z(n53003) );
  XOR U52815 ( .A(n53009), .B(n53010), .Z(n52628) );
  AND U52816 ( .A(n649), .B(n53011), .Z(n53010) );
  XOR U52817 ( .A(n53012), .B(n53009), .Z(n53011) );
  XOR U52818 ( .A(n53013), .B(n53014), .Z(n53001) );
  AND U52819 ( .A(n53015), .B(n53016), .Z(n53014) );
  XOR U52820 ( .A(n53013), .B(n52643), .Z(n53016) );
  XOR U52821 ( .A(n53017), .B(n53018), .Z(n52643) );
  AND U52822 ( .A(n651), .B(n53019), .Z(n53018) );
  XOR U52823 ( .A(n53020), .B(n53017), .Z(n53019) );
  XNOR U52824 ( .A(n52640), .B(n53013), .Z(n53015) );
  XOR U52825 ( .A(n53021), .B(n53022), .Z(n52640) );
  AND U52826 ( .A(n649), .B(n53023), .Z(n53022) );
  XOR U52827 ( .A(n53024), .B(n53021), .Z(n53023) );
  XOR U52828 ( .A(n53025), .B(n53026), .Z(n53013) );
  AND U52829 ( .A(n53027), .B(n53028), .Z(n53026) );
  XOR U52830 ( .A(n53025), .B(n52655), .Z(n53028) );
  XOR U52831 ( .A(n53029), .B(n53030), .Z(n52655) );
  AND U52832 ( .A(n651), .B(n53031), .Z(n53030) );
  XOR U52833 ( .A(n53032), .B(n53029), .Z(n53031) );
  XNOR U52834 ( .A(n52652), .B(n53025), .Z(n53027) );
  XOR U52835 ( .A(n53033), .B(n53034), .Z(n52652) );
  AND U52836 ( .A(n649), .B(n53035), .Z(n53034) );
  XOR U52837 ( .A(n53036), .B(n53033), .Z(n53035) );
  XOR U52838 ( .A(n53037), .B(n53038), .Z(n53025) );
  AND U52839 ( .A(n53039), .B(n53040), .Z(n53038) );
  XOR U52840 ( .A(n53037), .B(n52667), .Z(n53040) );
  XOR U52841 ( .A(n53041), .B(n53042), .Z(n52667) );
  AND U52842 ( .A(n651), .B(n53043), .Z(n53042) );
  XOR U52843 ( .A(n53044), .B(n53041), .Z(n53043) );
  XNOR U52844 ( .A(n52664), .B(n53037), .Z(n53039) );
  XOR U52845 ( .A(n53045), .B(n53046), .Z(n52664) );
  AND U52846 ( .A(n649), .B(n53047), .Z(n53046) );
  XOR U52847 ( .A(n53048), .B(n53045), .Z(n53047) );
  XOR U52848 ( .A(n53049), .B(n53050), .Z(n53037) );
  AND U52849 ( .A(n53051), .B(n53052), .Z(n53050) );
  XOR U52850 ( .A(n53049), .B(n52679), .Z(n53052) );
  XOR U52851 ( .A(n53053), .B(n53054), .Z(n52679) );
  AND U52852 ( .A(n651), .B(n53055), .Z(n53054) );
  XOR U52853 ( .A(n53056), .B(n53053), .Z(n53055) );
  XNOR U52854 ( .A(n52676), .B(n53049), .Z(n53051) );
  XOR U52855 ( .A(n53057), .B(n53058), .Z(n52676) );
  AND U52856 ( .A(n649), .B(n53059), .Z(n53058) );
  XOR U52857 ( .A(n53060), .B(n53057), .Z(n53059) );
  XOR U52858 ( .A(n53061), .B(n53062), .Z(n53049) );
  AND U52859 ( .A(n53063), .B(n53064), .Z(n53062) );
  XOR U52860 ( .A(n53061), .B(n52691), .Z(n53064) );
  XOR U52861 ( .A(n53065), .B(n53066), .Z(n52691) );
  AND U52862 ( .A(n651), .B(n53067), .Z(n53066) );
  XOR U52863 ( .A(n53068), .B(n53065), .Z(n53067) );
  XNOR U52864 ( .A(n52688), .B(n53061), .Z(n53063) );
  XOR U52865 ( .A(n53069), .B(n53070), .Z(n52688) );
  AND U52866 ( .A(n649), .B(n53071), .Z(n53070) );
  XOR U52867 ( .A(n53072), .B(n53069), .Z(n53071) );
  XOR U52868 ( .A(n53073), .B(n53074), .Z(n53061) );
  AND U52869 ( .A(n53075), .B(n53076), .Z(n53074) );
  XOR U52870 ( .A(n53073), .B(n52703), .Z(n53076) );
  XOR U52871 ( .A(n53077), .B(n53078), .Z(n52703) );
  AND U52872 ( .A(n651), .B(n53079), .Z(n53078) );
  XOR U52873 ( .A(n53080), .B(n53077), .Z(n53079) );
  XNOR U52874 ( .A(n52700), .B(n53073), .Z(n53075) );
  XOR U52875 ( .A(n53081), .B(n53082), .Z(n52700) );
  AND U52876 ( .A(n649), .B(n53083), .Z(n53082) );
  XOR U52877 ( .A(n53084), .B(n53081), .Z(n53083) );
  XOR U52878 ( .A(n53085), .B(n53086), .Z(n53073) );
  AND U52879 ( .A(n53087), .B(n53088), .Z(n53086) );
  XOR U52880 ( .A(n53085), .B(n52715), .Z(n53088) );
  XOR U52881 ( .A(n53089), .B(n53090), .Z(n52715) );
  AND U52882 ( .A(n651), .B(n53091), .Z(n53090) );
  XOR U52883 ( .A(n53092), .B(n53089), .Z(n53091) );
  XNOR U52884 ( .A(n52712), .B(n53085), .Z(n53087) );
  XOR U52885 ( .A(n53093), .B(n53094), .Z(n52712) );
  AND U52886 ( .A(n649), .B(n53095), .Z(n53094) );
  XOR U52887 ( .A(n53096), .B(n53093), .Z(n53095) );
  XOR U52888 ( .A(n53097), .B(n53098), .Z(n53085) );
  AND U52889 ( .A(n53099), .B(n53100), .Z(n53098) );
  XOR U52890 ( .A(n53097), .B(n52727), .Z(n53100) );
  XOR U52891 ( .A(n53101), .B(n53102), .Z(n52727) );
  AND U52892 ( .A(n651), .B(n53103), .Z(n53102) );
  XOR U52893 ( .A(n53104), .B(n53101), .Z(n53103) );
  XNOR U52894 ( .A(n52724), .B(n53097), .Z(n53099) );
  XOR U52895 ( .A(n53105), .B(n53106), .Z(n52724) );
  AND U52896 ( .A(n649), .B(n53107), .Z(n53106) );
  XOR U52897 ( .A(n53108), .B(n53105), .Z(n53107) );
  XOR U52898 ( .A(n53109), .B(n53110), .Z(n53097) );
  AND U52899 ( .A(n53111), .B(n53112), .Z(n53110) );
  XOR U52900 ( .A(n53109), .B(n52739), .Z(n53112) );
  XOR U52901 ( .A(n53113), .B(n53114), .Z(n52739) );
  AND U52902 ( .A(n651), .B(n53115), .Z(n53114) );
  XOR U52903 ( .A(n53116), .B(n53113), .Z(n53115) );
  XNOR U52904 ( .A(n52736), .B(n53109), .Z(n53111) );
  XOR U52905 ( .A(n53117), .B(n53118), .Z(n52736) );
  AND U52906 ( .A(n649), .B(n53119), .Z(n53118) );
  XOR U52907 ( .A(n53120), .B(n53117), .Z(n53119) );
  XOR U52908 ( .A(n53121), .B(n53122), .Z(n53109) );
  AND U52909 ( .A(n53123), .B(n53124), .Z(n53122) );
  XOR U52910 ( .A(n53121), .B(n52751), .Z(n53124) );
  XOR U52911 ( .A(n53125), .B(n53126), .Z(n52751) );
  AND U52912 ( .A(n651), .B(n53127), .Z(n53126) );
  XOR U52913 ( .A(n53128), .B(n53125), .Z(n53127) );
  XNOR U52914 ( .A(n52748), .B(n53121), .Z(n53123) );
  XOR U52915 ( .A(n53129), .B(n53130), .Z(n52748) );
  AND U52916 ( .A(n649), .B(n53131), .Z(n53130) );
  XOR U52917 ( .A(n53132), .B(n53129), .Z(n53131) );
  XOR U52918 ( .A(n53133), .B(n53134), .Z(n53121) );
  AND U52919 ( .A(n53135), .B(n53136), .Z(n53134) );
  XOR U52920 ( .A(n53133), .B(n52763), .Z(n53136) );
  XOR U52921 ( .A(n53137), .B(n53138), .Z(n52763) );
  AND U52922 ( .A(n651), .B(n53139), .Z(n53138) );
  XOR U52923 ( .A(n53140), .B(n53137), .Z(n53139) );
  XNOR U52924 ( .A(n52760), .B(n53133), .Z(n53135) );
  XOR U52925 ( .A(n53141), .B(n53142), .Z(n52760) );
  AND U52926 ( .A(n649), .B(n53143), .Z(n53142) );
  XOR U52927 ( .A(n53144), .B(n53141), .Z(n53143) );
  XOR U52928 ( .A(n53145), .B(n53146), .Z(n53133) );
  AND U52929 ( .A(n53147), .B(n53148), .Z(n53146) );
  XOR U52930 ( .A(n53145), .B(n52775), .Z(n53148) );
  XOR U52931 ( .A(n53149), .B(n53150), .Z(n52775) );
  AND U52932 ( .A(n651), .B(n53151), .Z(n53150) );
  XOR U52933 ( .A(n53152), .B(n53149), .Z(n53151) );
  XNOR U52934 ( .A(n52772), .B(n53145), .Z(n53147) );
  XOR U52935 ( .A(n53153), .B(n53154), .Z(n52772) );
  AND U52936 ( .A(n649), .B(n53155), .Z(n53154) );
  XOR U52937 ( .A(n53156), .B(n53153), .Z(n53155) );
  XOR U52938 ( .A(n53157), .B(n53158), .Z(n53145) );
  AND U52939 ( .A(n53159), .B(n53160), .Z(n53158) );
  XOR U52940 ( .A(n53157), .B(n52787), .Z(n53160) );
  XOR U52941 ( .A(n53161), .B(n53162), .Z(n52787) );
  AND U52942 ( .A(n651), .B(n53163), .Z(n53162) );
  XOR U52943 ( .A(n53164), .B(n53161), .Z(n53163) );
  XNOR U52944 ( .A(n52784), .B(n53157), .Z(n53159) );
  XOR U52945 ( .A(n53165), .B(n53166), .Z(n52784) );
  AND U52946 ( .A(n649), .B(n53167), .Z(n53166) );
  XOR U52947 ( .A(n53168), .B(n53165), .Z(n53167) );
  XOR U52948 ( .A(n53169), .B(n53170), .Z(n53157) );
  AND U52949 ( .A(n53171), .B(n53172), .Z(n53170) );
  XOR U52950 ( .A(n53169), .B(n52799), .Z(n53172) );
  XOR U52951 ( .A(n53173), .B(n53174), .Z(n52799) );
  AND U52952 ( .A(n651), .B(n53175), .Z(n53174) );
  XOR U52953 ( .A(n53176), .B(n53173), .Z(n53175) );
  XNOR U52954 ( .A(n52796), .B(n53169), .Z(n53171) );
  XOR U52955 ( .A(n53177), .B(n53178), .Z(n52796) );
  AND U52956 ( .A(n649), .B(n53179), .Z(n53178) );
  XOR U52957 ( .A(n53180), .B(n53177), .Z(n53179) );
  XOR U52958 ( .A(n53181), .B(n53182), .Z(n53169) );
  AND U52959 ( .A(n53183), .B(n53184), .Z(n53182) );
  XOR U52960 ( .A(n53181), .B(n52811), .Z(n53184) );
  XOR U52961 ( .A(n53185), .B(n53186), .Z(n52811) );
  AND U52962 ( .A(n651), .B(n53187), .Z(n53186) );
  XOR U52963 ( .A(n53188), .B(n53185), .Z(n53187) );
  XNOR U52964 ( .A(n52808), .B(n53181), .Z(n53183) );
  XOR U52965 ( .A(n53189), .B(n53190), .Z(n52808) );
  AND U52966 ( .A(n649), .B(n53191), .Z(n53190) );
  XOR U52967 ( .A(n53192), .B(n53189), .Z(n53191) );
  XOR U52968 ( .A(n53193), .B(n53194), .Z(n53181) );
  AND U52969 ( .A(n53195), .B(n53196), .Z(n53194) );
  XOR U52970 ( .A(n53193), .B(n52823), .Z(n53196) );
  XOR U52971 ( .A(n53197), .B(n53198), .Z(n52823) );
  AND U52972 ( .A(n651), .B(n53199), .Z(n53198) );
  XOR U52973 ( .A(n53200), .B(n53197), .Z(n53199) );
  XNOR U52974 ( .A(n52820), .B(n53193), .Z(n53195) );
  XOR U52975 ( .A(n53201), .B(n53202), .Z(n52820) );
  AND U52976 ( .A(n649), .B(n53203), .Z(n53202) );
  XOR U52977 ( .A(n53204), .B(n53201), .Z(n53203) );
  XOR U52978 ( .A(n53205), .B(n53206), .Z(n53193) );
  AND U52979 ( .A(n53207), .B(n53208), .Z(n53206) );
  XOR U52980 ( .A(n53205), .B(n52835), .Z(n53208) );
  XOR U52981 ( .A(n53209), .B(n53210), .Z(n52835) );
  AND U52982 ( .A(n651), .B(n53211), .Z(n53210) );
  XOR U52983 ( .A(n53212), .B(n53209), .Z(n53211) );
  XNOR U52984 ( .A(n52832), .B(n53205), .Z(n53207) );
  XOR U52985 ( .A(n53213), .B(n53214), .Z(n52832) );
  AND U52986 ( .A(n649), .B(n53215), .Z(n53214) );
  XOR U52987 ( .A(n53216), .B(n53213), .Z(n53215) );
  XOR U52988 ( .A(n53217), .B(n53218), .Z(n53205) );
  AND U52989 ( .A(n53219), .B(n53220), .Z(n53218) );
  XOR U52990 ( .A(n53217), .B(n52847), .Z(n53220) );
  XOR U52991 ( .A(n53221), .B(n53222), .Z(n52847) );
  AND U52992 ( .A(n651), .B(n53223), .Z(n53222) );
  XOR U52993 ( .A(n53224), .B(n53221), .Z(n53223) );
  XNOR U52994 ( .A(n52844), .B(n53217), .Z(n53219) );
  XOR U52995 ( .A(n53225), .B(n53226), .Z(n52844) );
  AND U52996 ( .A(n649), .B(n53227), .Z(n53226) );
  XOR U52997 ( .A(n53228), .B(n53225), .Z(n53227) );
  XOR U52998 ( .A(n53229), .B(n53230), .Z(n53217) );
  AND U52999 ( .A(n53231), .B(n53232), .Z(n53230) );
  XOR U53000 ( .A(n53229), .B(n52859), .Z(n53232) );
  XOR U53001 ( .A(n53233), .B(n53234), .Z(n52859) );
  AND U53002 ( .A(n651), .B(n53235), .Z(n53234) );
  XOR U53003 ( .A(n53236), .B(n53233), .Z(n53235) );
  XNOR U53004 ( .A(n52856), .B(n53229), .Z(n53231) );
  XOR U53005 ( .A(n53237), .B(n53238), .Z(n52856) );
  AND U53006 ( .A(n649), .B(n53239), .Z(n53238) );
  XOR U53007 ( .A(n53240), .B(n53237), .Z(n53239) );
  XOR U53008 ( .A(n53241), .B(n53242), .Z(n53229) );
  AND U53009 ( .A(n53243), .B(n53244), .Z(n53242) );
  XOR U53010 ( .A(n53241), .B(n52871), .Z(n53244) );
  XOR U53011 ( .A(n53245), .B(n53246), .Z(n52871) );
  AND U53012 ( .A(n651), .B(n53247), .Z(n53246) );
  XOR U53013 ( .A(n53248), .B(n53245), .Z(n53247) );
  XNOR U53014 ( .A(n52868), .B(n53241), .Z(n53243) );
  XOR U53015 ( .A(n53249), .B(n53250), .Z(n52868) );
  AND U53016 ( .A(n649), .B(n53251), .Z(n53250) );
  XOR U53017 ( .A(n53252), .B(n53249), .Z(n53251) );
  XOR U53018 ( .A(n53253), .B(n53254), .Z(n53241) );
  AND U53019 ( .A(n53255), .B(n53256), .Z(n53254) );
  XOR U53020 ( .A(n53253), .B(n52883), .Z(n53256) );
  XOR U53021 ( .A(n53257), .B(n53258), .Z(n52883) );
  AND U53022 ( .A(n651), .B(n53259), .Z(n53258) );
  XOR U53023 ( .A(n53260), .B(n53257), .Z(n53259) );
  XNOR U53024 ( .A(n52880), .B(n53253), .Z(n53255) );
  XOR U53025 ( .A(n53261), .B(n53262), .Z(n52880) );
  AND U53026 ( .A(n649), .B(n53263), .Z(n53262) );
  XOR U53027 ( .A(n53264), .B(n53261), .Z(n53263) );
  XOR U53028 ( .A(n53265), .B(n53266), .Z(n53253) );
  AND U53029 ( .A(n53267), .B(n53268), .Z(n53266) );
  XOR U53030 ( .A(n53265), .B(n52895), .Z(n53268) );
  XOR U53031 ( .A(n53269), .B(n53270), .Z(n52895) );
  AND U53032 ( .A(n651), .B(n53271), .Z(n53270) );
  XOR U53033 ( .A(n53272), .B(n53269), .Z(n53271) );
  XNOR U53034 ( .A(n52892), .B(n53265), .Z(n53267) );
  XOR U53035 ( .A(n53273), .B(n53274), .Z(n52892) );
  AND U53036 ( .A(n649), .B(n53275), .Z(n53274) );
  XOR U53037 ( .A(n53276), .B(n53273), .Z(n53275) );
  XOR U53038 ( .A(n53277), .B(n53278), .Z(n53265) );
  AND U53039 ( .A(n53279), .B(n53280), .Z(n53278) );
  XNOR U53040 ( .A(n53281), .B(n52908), .Z(n53280) );
  XOR U53041 ( .A(n53282), .B(n53283), .Z(n52908) );
  AND U53042 ( .A(n651), .B(n53284), .Z(n53283) );
  XOR U53043 ( .A(n53282), .B(n53285), .Z(n53284) );
  XNOR U53044 ( .A(n52905), .B(n53277), .Z(n53279) );
  XOR U53045 ( .A(n53286), .B(n53287), .Z(n52905) );
  AND U53046 ( .A(n649), .B(n53288), .Z(n53287) );
  XOR U53047 ( .A(n53286), .B(n53289), .Z(n53288) );
  IV U53048 ( .A(n53281), .Z(n53277) );
  AND U53049 ( .A(n52913), .B(n52916), .Z(n53281) );
  XNOR U53050 ( .A(n53290), .B(n53291), .Z(n52916) );
  AND U53051 ( .A(n651), .B(n53292), .Z(n53291) );
  XNOR U53052 ( .A(n53293), .B(n53290), .Z(n53292) );
  XOR U53053 ( .A(n53294), .B(n53295), .Z(n651) );
  AND U53054 ( .A(n53296), .B(n53297), .Z(n53295) );
  XOR U53055 ( .A(n52924), .B(n53294), .Z(n53297) );
  IV U53056 ( .A(n53298), .Z(n52924) );
  AND U53057 ( .A(p_input[991]), .B(p_input[1023]), .Z(n53298) );
  XOR U53058 ( .A(n53294), .B(n52921), .Z(n53296) );
  AND U53059 ( .A(p_input[927]), .B(p_input[959]), .Z(n52921) );
  XOR U53060 ( .A(n53299), .B(n53300), .Z(n53294) );
  AND U53061 ( .A(n53301), .B(n53302), .Z(n53300) );
  XOR U53062 ( .A(n53299), .B(n52936), .Z(n53302) );
  XNOR U53063 ( .A(p_input[990]), .B(n53303), .Z(n52936) );
  AND U53064 ( .A(n1059), .B(n53304), .Z(n53303) );
  XOR U53065 ( .A(p_input[990]), .B(p_input[1022]), .Z(n53304) );
  XNOR U53066 ( .A(n52933), .B(n53299), .Z(n53301) );
  XOR U53067 ( .A(n53305), .B(n53306), .Z(n52933) );
  AND U53068 ( .A(n1057), .B(n53307), .Z(n53306) );
  XOR U53069 ( .A(p_input[958]), .B(p_input[926]), .Z(n53307) );
  XOR U53070 ( .A(n53308), .B(n53309), .Z(n53299) );
  AND U53071 ( .A(n53310), .B(n53311), .Z(n53309) );
  XOR U53072 ( .A(n53308), .B(n52948), .Z(n53311) );
  XNOR U53073 ( .A(p_input[989]), .B(n53312), .Z(n52948) );
  AND U53074 ( .A(n1059), .B(n53313), .Z(n53312) );
  XOR U53075 ( .A(p_input[989]), .B(p_input[1021]), .Z(n53313) );
  XNOR U53076 ( .A(n52945), .B(n53308), .Z(n53310) );
  XOR U53077 ( .A(n53314), .B(n53315), .Z(n52945) );
  AND U53078 ( .A(n1057), .B(n53316), .Z(n53315) );
  XOR U53079 ( .A(p_input[957]), .B(p_input[925]), .Z(n53316) );
  XOR U53080 ( .A(n53317), .B(n53318), .Z(n53308) );
  AND U53081 ( .A(n53319), .B(n53320), .Z(n53318) );
  XOR U53082 ( .A(n53317), .B(n52960), .Z(n53320) );
  XNOR U53083 ( .A(p_input[988]), .B(n53321), .Z(n52960) );
  AND U53084 ( .A(n1059), .B(n53322), .Z(n53321) );
  XOR U53085 ( .A(p_input[988]), .B(p_input[1020]), .Z(n53322) );
  XNOR U53086 ( .A(n52957), .B(n53317), .Z(n53319) );
  XOR U53087 ( .A(n53323), .B(n53324), .Z(n52957) );
  AND U53088 ( .A(n1057), .B(n53325), .Z(n53324) );
  XOR U53089 ( .A(p_input[956]), .B(p_input[924]), .Z(n53325) );
  XOR U53090 ( .A(n53326), .B(n53327), .Z(n53317) );
  AND U53091 ( .A(n53328), .B(n53329), .Z(n53327) );
  XOR U53092 ( .A(n53326), .B(n52972), .Z(n53329) );
  XNOR U53093 ( .A(p_input[987]), .B(n53330), .Z(n52972) );
  AND U53094 ( .A(n1059), .B(n53331), .Z(n53330) );
  XOR U53095 ( .A(p_input[987]), .B(p_input[1019]), .Z(n53331) );
  XNOR U53096 ( .A(n52969), .B(n53326), .Z(n53328) );
  XOR U53097 ( .A(n53332), .B(n53333), .Z(n52969) );
  AND U53098 ( .A(n1057), .B(n53334), .Z(n53333) );
  XOR U53099 ( .A(p_input[955]), .B(p_input[923]), .Z(n53334) );
  XOR U53100 ( .A(n53335), .B(n53336), .Z(n53326) );
  AND U53101 ( .A(n53337), .B(n53338), .Z(n53336) );
  XOR U53102 ( .A(n53335), .B(n52984), .Z(n53338) );
  XNOR U53103 ( .A(p_input[986]), .B(n53339), .Z(n52984) );
  AND U53104 ( .A(n1059), .B(n53340), .Z(n53339) );
  XOR U53105 ( .A(p_input[986]), .B(p_input[1018]), .Z(n53340) );
  XNOR U53106 ( .A(n52981), .B(n53335), .Z(n53337) );
  XOR U53107 ( .A(n53341), .B(n53342), .Z(n52981) );
  AND U53108 ( .A(n1057), .B(n53343), .Z(n53342) );
  XOR U53109 ( .A(p_input[954]), .B(p_input[922]), .Z(n53343) );
  XOR U53110 ( .A(n53344), .B(n53345), .Z(n53335) );
  AND U53111 ( .A(n53346), .B(n53347), .Z(n53345) );
  XOR U53112 ( .A(n53344), .B(n52996), .Z(n53347) );
  XNOR U53113 ( .A(p_input[985]), .B(n53348), .Z(n52996) );
  AND U53114 ( .A(n1059), .B(n53349), .Z(n53348) );
  XOR U53115 ( .A(p_input[985]), .B(p_input[1017]), .Z(n53349) );
  XNOR U53116 ( .A(n52993), .B(n53344), .Z(n53346) );
  XOR U53117 ( .A(n53350), .B(n53351), .Z(n52993) );
  AND U53118 ( .A(n1057), .B(n53352), .Z(n53351) );
  XOR U53119 ( .A(p_input[953]), .B(p_input[921]), .Z(n53352) );
  XOR U53120 ( .A(n53353), .B(n53354), .Z(n53344) );
  AND U53121 ( .A(n53355), .B(n53356), .Z(n53354) );
  XOR U53122 ( .A(n53353), .B(n53008), .Z(n53356) );
  XNOR U53123 ( .A(p_input[984]), .B(n53357), .Z(n53008) );
  AND U53124 ( .A(n1059), .B(n53358), .Z(n53357) );
  XOR U53125 ( .A(p_input[984]), .B(p_input[1016]), .Z(n53358) );
  XNOR U53126 ( .A(n53005), .B(n53353), .Z(n53355) );
  XOR U53127 ( .A(n53359), .B(n53360), .Z(n53005) );
  AND U53128 ( .A(n1057), .B(n53361), .Z(n53360) );
  XOR U53129 ( .A(p_input[952]), .B(p_input[920]), .Z(n53361) );
  XOR U53130 ( .A(n53362), .B(n53363), .Z(n53353) );
  AND U53131 ( .A(n53364), .B(n53365), .Z(n53363) );
  XOR U53132 ( .A(n53362), .B(n53020), .Z(n53365) );
  XNOR U53133 ( .A(p_input[983]), .B(n53366), .Z(n53020) );
  AND U53134 ( .A(n1059), .B(n53367), .Z(n53366) );
  XOR U53135 ( .A(p_input[983]), .B(p_input[1015]), .Z(n53367) );
  XNOR U53136 ( .A(n53017), .B(n53362), .Z(n53364) );
  XOR U53137 ( .A(n53368), .B(n53369), .Z(n53017) );
  AND U53138 ( .A(n1057), .B(n53370), .Z(n53369) );
  XOR U53139 ( .A(p_input[951]), .B(p_input[919]), .Z(n53370) );
  XOR U53140 ( .A(n53371), .B(n53372), .Z(n53362) );
  AND U53141 ( .A(n53373), .B(n53374), .Z(n53372) );
  XOR U53142 ( .A(n53371), .B(n53032), .Z(n53374) );
  XNOR U53143 ( .A(p_input[982]), .B(n53375), .Z(n53032) );
  AND U53144 ( .A(n1059), .B(n53376), .Z(n53375) );
  XOR U53145 ( .A(p_input[982]), .B(p_input[1014]), .Z(n53376) );
  XNOR U53146 ( .A(n53029), .B(n53371), .Z(n53373) );
  XOR U53147 ( .A(n53377), .B(n53378), .Z(n53029) );
  AND U53148 ( .A(n1057), .B(n53379), .Z(n53378) );
  XOR U53149 ( .A(p_input[950]), .B(p_input[918]), .Z(n53379) );
  XOR U53150 ( .A(n53380), .B(n53381), .Z(n53371) );
  AND U53151 ( .A(n53382), .B(n53383), .Z(n53381) );
  XOR U53152 ( .A(n53380), .B(n53044), .Z(n53383) );
  XNOR U53153 ( .A(p_input[981]), .B(n53384), .Z(n53044) );
  AND U53154 ( .A(n1059), .B(n53385), .Z(n53384) );
  XOR U53155 ( .A(p_input[981]), .B(p_input[1013]), .Z(n53385) );
  XNOR U53156 ( .A(n53041), .B(n53380), .Z(n53382) );
  XOR U53157 ( .A(n53386), .B(n53387), .Z(n53041) );
  AND U53158 ( .A(n1057), .B(n53388), .Z(n53387) );
  XOR U53159 ( .A(p_input[949]), .B(p_input[917]), .Z(n53388) );
  XOR U53160 ( .A(n53389), .B(n53390), .Z(n53380) );
  AND U53161 ( .A(n53391), .B(n53392), .Z(n53390) );
  XOR U53162 ( .A(n53389), .B(n53056), .Z(n53392) );
  XNOR U53163 ( .A(p_input[980]), .B(n53393), .Z(n53056) );
  AND U53164 ( .A(n1059), .B(n53394), .Z(n53393) );
  XOR U53165 ( .A(p_input[980]), .B(p_input[1012]), .Z(n53394) );
  XNOR U53166 ( .A(n53053), .B(n53389), .Z(n53391) );
  XOR U53167 ( .A(n53395), .B(n53396), .Z(n53053) );
  AND U53168 ( .A(n1057), .B(n53397), .Z(n53396) );
  XOR U53169 ( .A(p_input[948]), .B(p_input[916]), .Z(n53397) );
  XOR U53170 ( .A(n53398), .B(n53399), .Z(n53389) );
  AND U53171 ( .A(n53400), .B(n53401), .Z(n53399) );
  XOR U53172 ( .A(n53398), .B(n53068), .Z(n53401) );
  XNOR U53173 ( .A(p_input[979]), .B(n53402), .Z(n53068) );
  AND U53174 ( .A(n1059), .B(n53403), .Z(n53402) );
  XOR U53175 ( .A(p_input[979]), .B(p_input[1011]), .Z(n53403) );
  XNOR U53176 ( .A(n53065), .B(n53398), .Z(n53400) );
  XOR U53177 ( .A(n53404), .B(n53405), .Z(n53065) );
  AND U53178 ( .A(n1057), .B(n53406), .Z(n53405) );
  XOR U53179 ( .A(p_input[947]), .B(p_input[915]), .Z(n53406) );
  XOR U53180 ( .A(n53407), .B(n53408), .Z(n53398) );
  AND U53181 ( .A(n53409), .B(n53410), .Z(n53408) );
  XOR U53182 ( .A(n53407), .B(n53080), .Z(n53410) );
  XNOR U53183 ( .A(p_input[978]), .B(n53411), .Z(n53080) );
  AND U53184 ( .A(n1059), .B(n53412), .Z(n53411) );
  XOR U53185 ( .A(p_input[978]), .B(p_input[1010]), .Z(n53412) );
  XNOR U53186 ( .A(n53077), .B(n53407), .Z(n53409) );
  XOR U53187 ( .A(n53413), .B(n53414), .Z(n53077) );
  AND U53188 ( .A(n1057), .B(n53415), .Z(n53414) );
  XOR U53189 ( .A(p_input[946]), .B(p_input[914]), .Z(n53415) );
  XOR U53190 ( .A(n53416), .B(n53417), .Z(n53407) );
  AND U53191 ( .A(n53418), .B(n53419), .Z(n53417) );
  XOR U53192 ( .A(n53416), .B(n53092), .Z(n53419) );
  XNOR U53193 ( .A(p_input[977]), .B(n53420), .Z(n53092) );
  AND U53194 ( .A(n1059), .B(n53421), .Z(n53420) );
  XOR U53195 ( .A(p_input[977]), .B(p_input[1009]), .Z(n53421) );
  XNOR U53196 ( .A(n53089), .B(n53416), .Z(n53418) );
  XOR U53197 ( .A(n53422), .B(n53423), .Z(n53089) );
  AND U53198 ( .A(n1057), .B(n53424), .Z(n53423) );
  XOR U53199 ( .A(p_input[945]), .B(p_input[913]), .Z(n53424) );
  XOR U53200 ( .A(n53425), .B(n53426), .Z(n53416) );
  AND U53201 ( .A(n53427), .B(n53428), .Z(n53426) );
  XOR U53202 ( .A(n53425), .B(n53104), .Z(n53428) );
  XNOR U53203 ( .A(p_input[976]), .B(n53429), .Z(n53104) );
  AND U53204 ( .A(n1059), .B(n53430), .Z(n53429) );
  XOR U53205 ( .A(p_input[976]), .B(p_input[1008]), .Z(n53430) );
  XNOR U53206 ( .A(n53101), .B(n53425), .Z(n53427) );
  XOR U53207 ( .A(n53431), .B(n53432), .Z(n53101) );
  AND U53208 ( .A(n1057), .B(n53433), .Z(n53432) );
  XOR U53209 ( .A(p_input[944]), .B(p_input[912]), .Z(n53433) );
  XOR U53210 ( .A(n53434), .B(n53435), .Z(n53425) );
  AND U53211 ( .A(n53436), .B(n53437), .Z(n53435) );
  XOR U53212 ( .A(n53434), .B(n53116), .Z(n53437) );
  XNOR U53213 ( .A(p_input[975]), .B(n53438), .Z(n53116) );
  AND U53214 ( .A(n1059), .B(n53439), .Z(n53438) );
  XOR U53215 ( .A(p_input[975]), .B(p_input[1007]), .Z(n53439) );
  XNOR U53216 ( .A(n53113), .B(n53434), .Z(n53436) );
  XOR U53217 ( .A(n53440), .B(n53441), .Z(n53113) );
  AND U53218 ( .A(n1057), .B(n53442), .Z(n53441) );
  XOR U53219 ( .A(p_input[943]), .B(p_input[911]), .Z(n53442) );
  XOR U53220 ( .A(n53443), .B(n53444), .Z(n53434) );
  AND U53221 ( .A(n53445), .B(n53446), .Z(n53444) );
  XOR U53222 ( .A(n53443), .B(n53128), .Z(n53446) );
  XNOR U53223 ( .A(p_input[974]), .B(n53447), .Z(n53128) );
  AND U53224 ( .A(n1059), .B(n53448), .Z(n53447) );
  XOR U53225 ( .A(p_input[974]), .B(p_input[1006]), .Z(n53448) );
  XNOR U53226 ( .A(n53125), .B(n53443), .Z(n53445) );
  XOR U53227 ( .A(n53449), .B(n53450), .Z(n53125) );
  AND U53228 ( .A(n1057), .B(n53451), .Z(n53450) );
  XOR U53229 ( .A(p_input[942]), .B(p_input[910]), .Z(n53451) );
  XOR U53230 ( .A(n53452), .B(n53453), .Z(n53443) );
  AND U53231 ( .A(n53454), .B(n53455), .Z(n53453) );
  XOR U53232 ( .A(n53452), .B(n53140), .Z(n53455) );
  XNOR U53233 ( .A(p_input[973]), .B(n53456), .Z(n53140) );
  AND U53234 ( .A(n1059), .B(n53457), .Z(n53456) );
  XOR U53235 ( .A(p_input[973]), .B(p_input[1005]), .Z(n53457) );
  XNOR U53236 ( .A(n53137), .B(n53452), .Z(n53454) );
  XOR U53237 ( .A(n53458), .B(n53459), .Z(n53137) );
  AND U53238 ( .A(n1057), .B(n53460), .Z(n53459) );
  XOR U53239 ( .A(p_input[941]), .B(p_input[909]), .Z(n53460) );
  XOR U53240 ( .A(n53461), .B(n53462), .Z(n53452) );
  AND U53241 ( .A(n53463), .B(n53464), .Z(n53462) );
  XOR U53242 ( .A(n53461), .B(n53152), .Z(n53464) );
  XNOR U53243 ( .A(p_input[972]), .B(n53465), .Z(n53152) );
  AND U53244 ( .A(n1059), .B(n53466), .Z(n53465) );
  XOR U53245 ( .A(p_input[972]), .B(p_input[1004]), .Z(n53466) );
  XNOR U53246 ( .A(n53149), .B(n53461), .Z(n53463) );
  XOR U53247 ( .A(n53467), .B(n53468), .Z(n53149) );
  AND U53248 ( .A(n1057), .B(n53469), .Z(n53468) );
  XOR U53249 ( .A(p_input[940]), .B(p_input[908]), .Z(n53469) );
  XOR U53250 ( .A(n53470), .B(n53471), .Z(n53461) );
  AND U53251 ( .A(n53472), .B(n53473), .Z(n53471) );
  XOR U53252 ( .A(n53470), .B(n53164), .Z(n53473) );
  XNOR U53253 ( .A(p_input[971]), .B(n53474), .Z(n53164) );
  AND U53254 ( .A(n1059), .B(n53475), .Z(n53474) );
  XOR U53255 ( .A(p_input[971]), .B(p_input[1003]), .Z(n53475) );
  XNOR U53256 ( .A(n53161), .B(n53470), .Z(n53472) );
  XOR U53257 ( .A(n53476), .B(n53477), .Z(n53161) );
  AND U53258 ( .A(n1057), .B(n53478), .Z(n53477) );
  XOR U53259 ( .A(p_input[939]), .B(p_input[907]), .Z(n53478) );
  XOR U53260 ( .A(n53479), .B(n53480), .Z(n53470) );
  AND U53261 ( .A(n53481), .B(n53482), .Z(n53480) );
  XOR U53262 ( .A(n53479), .B(n53176), .Z(n53482) );
  XNOR U53263 ( .A(p_input[970]), .B(n53483), .Z(n53176) );
  AND U53264 ( .A(n1059), .B(n53484), .Z(n53483) );
  XOR U53265 ( .A(p_input[970]), .B(p_input[1002]), .Z(n53484) );
  XNOR U53266 ( .A(n53173), .B(n53479), .Z(n53481) );
  XOR U53267 ( .A(n53485), .B(n53486), .Z(n53173) );
  AND U53268 ( .A(n1057), .B(n53487), .Z(n53486) );
  XOR U53269 ( .A(p_input[938]), .B(p_input[906]), .Z(n53487) );
  XOR U53270 ( .A(n53488), .B(n53489), .Z(n53479) );
  AND U53271 ( .A(n53490), .B(n53491), .Z(n53489) );
  XOR U53272 ( .A(n53488), .B(n53188), .Z(n53491) );
  XNOR U53273 ( .A(p_input[969]), .B(n53492), .Z(n53188) );
  AND U53274 ( .A(n1059), .B(n53493), .Z(n53492) );
  XOR U53275 ( .A(p_input[969]), .B(p_input[1001]), .Z(n53493) );
  XNOR U53276 ( .A(n53185), .B(n53488), .Z(n53490) );
  XOR U53277 ( .A(n53494), .B(n53495), .Z(n53185) );
  AND U53278 ( .A(n1057), .B(n53496), .Z(n53495) );
  XOR U53279 ( .A(p_input[937]), .B(p_input[905]), .Z(n53496) );
  XOR U53280 ( .A(n53497), .B(n53498), .Z(n53488) );
  AND U53281 ( .A(n53499), .B(n53500), .Z(n53498) );
  XOR U53282 ( .A(n53497), .B(n53200), .Z(n53500) );
  XNOR U53283 ( .A(p_input[968]), .B(n53501), .Z(n53200) );
  AND U53284 ( .A(n1059), .B(n53502), .Z(n53501) );
  XOR U53285 ( .A(p_input[968]), .B(p_input[1000]), .Z(n53502) );
  XNOR U53286 ( .A(n53197), .B(n53497), .Z(n53499) );
  XOR U53287 ( .A(n53503), .B(n53504), .Z(n53197) );
  AND U53288 ( .A(n1057), .B(n53505), .Z(n53504) );
  XOR U53289 ( .A(p_input[936]), .B(p_input[904]), .Z(n53505) );
  XOR U53290 ( .A(n53506), .B(n53507), .Z(n53497) );
  AND U53291 ( .A(n53508), .B(n53509), .Z(n53507) );
  XOR U53292 ( .A(n53506), .B(n53212), .Z(n53509) );
  XNOR U53293 ( .A(p_input[967]), .B(n53510), .Z(n53212) );
  AND U53294 ( .A(n1059), .B(n53511), .Z(n53510) );
  XOR U53295 ( .A(p_input[999]), .B(p_input[967]), .Z(n53511) );
  XNOR U53296 ( .A(n53209), .B(n53506), .Z(n53508) );
  XOR U53297 ( .A(n53512), .B(n53513), .Z(n53209) );
  AND U53298 ( .A(n1057), .B(n53514), .Z(n53513) );
  XOR U53299 ( .A(p_input[935]), .B(p_input[903]), .Z(n53514) );
  XOR U53300 ( .A(n53515), .B(n53516), .Z(n53506) );
  AND U53301 ( .A(n53517), .B(n53518), .Z(n53516) );
  XOR U53302 ( .A(n53515), .B(n53224), .Z(n53518) );
  XNOR U53303 ( .A(p_input[966]), .B(n53519), .Z(n53224) );
  AND U53304 ( .A(n1059), .B(n53520), .Z(n53519) );
  XOR U53305 ( .A(p_input[998]), .B(p_input[966]), .Z(n53520) );
  XNOR U53306 ( .A(n53221), .B(n53515), .Z(n53517) );
  XOR U53307 ( .A(n53521), .B(n53522), .Z(n53221) );
  AND U53308 ( .A(n1057), .B(n53523), .Z(n53522) );
  XOR U53309 ( .A(p_input[934]), .B(p_input[902]), .Z(n53523) );
  XOR U53310 ( .A(n53524), .B(n53525), .Z(n53515) );
  AND U53311 ( .A(n53526), .B(n53527), .Z(n53525) );
  XOR U53312 ( .A(n53524), .B(n53236), .Z(n53527) );
  XNOR U53313 ( .A(p_input[965]), .B(n53528), .Z(n53236) );
  AND U53314 ( .A(n1059), .B(n53529), .Z(n53528) );
  XOR U53315 ( .A(p_input[997]), .B(p_input[965]), .Z(n53529) );
  XNOR U53316 ( .A(n53233), .B(n53524), .Z(n53526) );
  XOR U53317 ( .A(n53530), .B(n53531), .Z(n53233) );
  AND U53318 ( .A(n1057), .B(n53532), .Z(n53531) );
  XOR U53319 ( .A(p_input[933]), .B(p_input[901]), .Z(n53532) );
  XOR U53320 ( .A(n53533), .B(n53534), .Z(n53524) );
  AND U53321 ( .A(n53535), .B(n53536), .Z(n53534) );
  XOR U53322 ( .A(n53533), .B(n53248), .Z(n53536) );
  XNOR U53323 ( .A(p_input[964]), .B(n53537), .Z(n53248) );
  AND U53324 ( .A(n1059), .B(n53538), .Z(n53537) );
  XOR U53325 ( .A(p_input[996]), .B(p_input[964]), .Z(n53538) );
  XNOR U53326 ( .A(n53245), .B(n53533), .Z(n53535) );
  XOR U53327 ( .A(n53539), .B(n53540), .Z(n53245) );
  AND U53328 ( .A(n1057), .B(n53541), .Z(n53540) );
  XOR U53329 ( .A(p_input[932]), .B(p_input[900]), .Z(n53541) );
  XOR U53330 ( .A(n53542), .B(n53543), .Z(n53533) );
  AND U53331 ( .A(n53544), .B(n53545), .Z(n53543) );
  XOR U53332 ( .A(n53542), .B(n53260), .Z(n53545) );
  XNOR U53333 ( .A(p_input[963]), .B(n53546), .Z(n53260) );
  AND U53334 ( .A(n1059), .B(n53547), .Z(n53546) );
  XOR U53335 ( .A(p_input[995]), .B(p_input[963]), .Z(n53547) );
  XNOR U53336 ( .A(n53257), .B(n53542), .Z(n53544) );
  XOR U53337 ( .A(n53548), .B(n53549), .Z(n53257) );
  AND U53338 ( .A(n1057), .B(n53550), .Z(n53549) );
  XOR U53339 ( .A(p_input[931]), .B(p_input[899]), .Z(n53550) );
  XOR U53340 ( .A(n53551), .B(n53552), .Z(n53542) );
  AND U53341 ( .A(n53553), .B(n53554), .Z(n53552) );
  XOR U53342 ( .A(n53551), .B(n53272), .Z(n53554) );
  XNOR U53343 ( .A(p_input[962]), .B(n53555), .Z(n53272) );
  AND U53344 ( .A(n1059), .B(n53556), .Z(n53555) );
  XOR U53345 ( .A(p_input[994]), .B(p_input[962]), .Z(n53556) );
  XNOR U53346 ( .A(n53269), .B(n53551), .Z(n53553) );
  XOR U53347 ( .A(n53557), .B(n53558), .Z(n53269) );
  AND U53348 ( .A(n1057), .B(n53559), .Z(n53558) );
  XOR U53349 ( .A(p_input[930]), .B(p_input[898]), .Z(n53559) );
  XOR U53350 ( .A(n53560), .B(n53561), .Z(n53551) );
  AND U53351 ( .A(n53562), .B(n53563), .Z(n53561) );
  XNOR U53352 ( .A(n53564), .B(n53285), .Z(n53563) );
  XNOR U53353 ( .A(p_input[961]), .B(n53565), .Z(n53285) );
  AND U53354 ( .A(n1059), .B(n53566), .Z(n53565) );
  XNOR U53355 ( .A(p_input[993]), .B(n53567), .Z(n53566) );
  IV U53356 ( .A(p_input[961]), .Z(n53567) );
  XNOR U53357 ( .A(n53282), .B(n53560), .Z(n53562) );
  XNOR U53358 ( .A(p_input[897]), .B(n53568), .Z(n53282) );
  AND U53359 ( .A(n1057), .B(n53569), .Z(n53568) );
  XOR U53360 ( .A(p_input[929]), .B(p_input[897]), .Z(n53569) );
  IV U53361 ( .A(n53564), .Z(n53560) );
  AND U53362 ( .A(n53290), .B(n53293), .Z(n53564) );
  XOR U53363 ( .A(p_input[960]), .B(n53570), .Z(n53293) );
  AND U53364 ( .A(n1059), .B(n53571), .Z(n53570) );
  XOR U53365 ( .A(p_input[992]), .B(p_input[960]), .Z(n53571) );
  XOR U53366 ( .A(n53572), .B(n53573), .Z(n1059) );
  AND U53367 ( .A(n53574), .B(n53575), .Z(n53573) );
  XNOR U53368 ( .A(p_input[1023]), .B(n53572), .Z(n53575) );
  XOR U53369 ( .A(n53572), .B(p_input[991]), .Z(n53574) );
  XOR U53370 ( .A(n53576), .B(n53577), .Z(n53572) );
  AND U53371 ( .A(n53578), .B(n53579), .Z(n53577) );
  XNOR U53372 ( .A(p_input[1022]), .B(n53576), .Z(n53579) );
  XOR U53373 ( .A(n53576), .B(p_input[990]), .Z(n53578) );
  XOR U53374 ( .A(n53580), .B(n53581), .Z(n53576) );
  AND U53375 ( .A(n53582), .B(n53583), .Z(n53581) );
  XNOR U53376 ( .A(p_input[1021]), .B(n53580), .Z(n53583) );
  XOR U53377 ( .A(n53580), .B(p_input[989]), .Z(n53582) );
  XOR U53378 ( .A(n53584), .B(n53585), .Z(n53580) );
  AND U53379 ( .A(n53586), .B(n53587), .Z(n53585) );
  XNOR U53380 ( .A(p_input[1020]), .B(n53584), .Z(n53587) );
  XOR U53381 ( .A(n53584), .B(p_input[988]), .Z(n53586) );
  XOR U53382 ( .A(n53588), .B(n53589), .Z(n53584) );
  AND U53383 ( .A(n53590), .B(n53591), .Z(n53589) );
  XNOR U53384 ( .A(p_input[1019]), .B(n53588), .Z(n53591) );
  XOR U53385 ( .A(n53588), .B(p_input[987]), .Z(n53590) );
  XOR U53386 ( .A(n53592), .B(n53593), .Z(n53588) );
  AND U53387 ( .A(n53594), .B(n53595), .Z(n53593) );
  XNOR U53388 ( .A(p_input[1018]), .B(n53592), .Z(n53595) );
  XOR U53389 ( .A(n53592), .B(p_input[986]), .Z(n53594) );
  XOR U53390 ( .A(n53596), .B(n53597), .Z(n53592) );
  AND U53391 ( .A(n53598), .B(n53599), .Z(n53597) );
  XNOR U53392 ( .A(p_input[1017]), .B(n53596), .Z(n53599) );
  XOR U53393 ( .A(n53596), .B(p_input[985]), .Z(n53598) );
  XOR U53394 ( .A(n53600), .B(n53601), .Z(n53596) );
  AND U53395 ( .A(n53602), .B(n53603), .Z(n53601) );
  XNOR U53396 ( .A(p_input[1016]), .B(n53600), .Z(n53603) );
  XOR U53397 ( .A(n53600), .B(p_input[984]), .Z(n53602) );
  XOR U53398 ( .A(n53604), .B(n53605), .Z(n53600) );
  AND U53399 ( .A(n53606), .B(n53607), .Z(n53605) );
  XNOR U53400 ( .A(p_input[1015]), .B(n53604), .Z(n53607) );
  XOR U53401 ( .A(n53604), .B(p_input[983]), .Z(n53606) );
  XOR U53402 ( .A(n53608), .B(n53609), .Z(n53604) );
  AND U53403 ( .A(n53610), .B(n53611), .Z(n53609) );
  XNOR U53404 ( .A(p_input[1014]), .B(n53608), .Z(n53611) );
  XOR U53405 ( .A(n53608), .B(p_input[982]), .Z(n53610) );
  XOR U53406 ( .A(n53612), .B(n53613), .Z(n53608) );
  AND U53407 ( .A(n53614), .B(n53615), .Z(n53613) );
  XNOR U53408 ( .A(p_input[1013]), .B(n53612), .Z(n53615) );
  XOR U53409 ( .A(n53612), .B(p_input[981]), .Z(n53614) );
  XOR U53410 ( .A(n53616), .B(n53617), .Z(n53612) );
  AND U53411 ( .A(n53618), .B(n53619), .Z(n53617) );
  XNOR U53412 ( .A(p_input[1012]), .B(n53616), .Z(n53619) );
  XOR U53413 ( .A(n53616), .B(p_input[980]), .Z(n53618) );
  XOR U53414 ( .A(n53620), .B(n53621), .Z(n53616) );
  AND U53415 ( .A(n53622), .B(n53623), .Z(n53621) );
  XNOR U53416 ( .A(p_input[1011]), .B(n53620), .Z(n53623) );
  XOR U53417 ( .A(n53620), .B(p_input[979]), .Z(n53622) );
  XOR U53418 ( .A(n53624), .B(n53625), .Z(n53620) );
  AND U53419 ( .A(n53626), .B(n53627), .Z(n53625) );
  XNOR U53420 ( .A(p_input[1010]), .B(n53624), .Z(n53627) );
  XOR U53421 ( .A(n53624), .B(p_input[978]), .Z(n53626) );
  XOR U53422 ( .A(n53628), .B(n53629), .Z(n53624) );
  AND U53423 ( .A(n53630), .B(n53631), .Z(n53629) );
  XNOR U53424 ( .A(p_input[1009]), .B(n53628), .Z(n53631) );
  XOR U53425 ( .A(n53628), .B(p_input[977]), .Z(n53630) );
  XOR U53426 ( .A(n53632), .B(n53633), .Z(n53628) );
  AND U53427 ( .A(n53634), .B(n53635), .Z(n53633) );
  XNOR U53428 ( .A(p_input[1008]), .B(n53632), .Z(n53635) );
  XOR U53429 ( .A(n53632), .B(p_input[976]), .Z(n53634) );
  XOR U53430 ( .A(n53636), .B(n53637), .Z(n53632) );
  AND U53431 ( .A(n53638), .B(n53639), .Z(n53637) );
  XNOR U53432 ( .A(p_input[1007]), .B(n53636), .Z(n53639) );
  XOR U53433 ( .A(n53636), .B(p_input[975]), .Z(n53638) );
  XOR U53434 ( .A(n53640), .B(n53641), .Z(n53636) );
  AND U53435 ( .A(n53642), .B(n53643), .Z(n53641) );
  XNOR U53436 ( .A(p_input[1006]), .B(n53640), .Z(n53643) );
  XOR U53437 ( .A(n53640), .B(p_input[974]), .Z(n53642) );
  XOR U53438 ( .A(n53644), .B(n53645), .Z(n53640) );
  AND U53439 ( .A(n53646), .B(n53647), .Z(n53645) );
  XNOR U53440 ( .A(p_input[1005]), .B(n53644), .Z(n53647) );
  XOR U53441 ( .A(n53644), .B(p_input[973]), .Z(n53646) );
  XOR U53442 ( .A(n53648), .B(n53649), .Z(n53644) );
  AND U53443 ( .A(n53650), .B(n53651), .Z(n53649) );
  XNOR U53444 ( .A(p_input[1004]), .B(n53648), .Z(n53651) );
  XOR U53445 ( .A(n53648), .B(p_input[972]), .Z(n53650) );
  XOR U53446 ( .A(n53652), .B(n53653), .Z(n53648) );
  AND U53447 ( .A(n53654), .B(n53655), .Z(n53653) );
  XNOR U53448 ( .A(p_input[1003]), .B(n53652), .Z(n53655) );
  XOR U53449 ( .A(n53652), .B(p_input[971]), .Z(n53654) );
  XOR U53450 ( .A(n53656), .B(n53657), .Z(n53652) );
  AND U53451 ( .A(n53658), .B(n53659), .Z(n53657) );
  XNOR U53452 ( .A(p_input[1002]), .B(n53656), .Z(n53659) );
  XOR U53453 ( .A(n53656), .B(p_input[970]), .Z(n53658) );
  XOR U53454 ( .A(n53660), .B(n53661), .Z(n53656) );
  AND U53455 ( .A(n53662), .B(n53663), .Z(n53661) );
  XNOR U53456 ( .A(p_input[1001]), .B(n53660), .Z(n53663) );
  XOR U53457 ( .A(n53660), .B(p_input[969]), .Z(n53662) );
  XOR U53458 ( .A(n53664), .B(n53665), .Z(n53660) );
  AND U53459 ( .A(n53666), .B(n53667), .Z(n53665) );
  XNOR U53460 ( .A(p_input[1000]), .B(n53664), .Z(n53667) );
  XOR U53461 ( .A(n53664), .B(p_input[968]), .Z(n53666) );
  XOR U53462 ( .A(n53668), .B(n53669), .Z(n53664) );
  AND U53463 ( .A(n53670), .B(n53671), .Z(n53669) );
  XNOR U53464 ( .A(p_input[999]), .B(n53668), .Z(n53671) );
  XOR U53465 ( .A(n53668), .B(p_input[967]), .Z(n53670) );
  XOR U53466 ( .A(n53672), .B(n53673), .Z(n53668) );
  AND U53467 ( .A(n53674), .B(n53675), .Z(n53673) );
  XNOR U53468 ( .A(p_input[998]), .B(n53672), .Z(n53675) );
  XOR U53469 ( .A(n53672), .B(p_input[966]), .Z(n53674) );
  XOR U53470 ( .A(n53676), .B(n53677), .Z(n53672) );
  AND U53471 ( .A(n53678), .B(n53679), .Z(n53677) );
  XNOR U53472 ( .A(p_input[997]), .B(n53676), .Z(n53679) );
  XOR U53473 ( .A(n53676), .B(p_input[965]), .Z(n53678) );
  XOR U53474 ( .A(n53680), .B(n53681), .Z(n53676) );
  AND U53475 ( .A(n53682), .B(n53683), .Z(n53681) );
  XNOR U53476 ( .A(p_input[996]), .B(n53680), .Z(n53683) );
  XOR U53477 ( .A(n53680), .B(p_input[964]), .Z(n53682) );
  XOR U53478 ( .A(n53684), .B(n53685), .Z(n53680) );
  AND U53479 ( .A(n53686), .B(n53687), .Z(n53685) );
  XNOR U53480 ( .A(p_input[995]), .B(n53684), .Z(n53687) );
  XOR U53481 ( .A(n53684), .B(p_input[963]), .Z(n53686) );
  XOR U53482 ( .A(n53688), .B(n53689), .Z(n53684) );
  AND U53483 ( .A(n53690), .B(n53691), .Z(n53689) );
  XNOR U53484 ( .A(p_input[994]), .B(n53688), .Z(n53691) );
  XOR U53485 ( .A(n53688), .B(p_input[962]), .Z(n53690) );
  XNOR U53486 ( .A(n53692), .B(n53693), .Z(n53688) );
  AND U53487 ( .A(n53694), .B(n53695), .Z(n53693) );
  XOR U53488 ( .A(p_input[993]), .B(n53692), .Z(n53695) );
  XNOR U53489 ( .A(p_input[961]), .B(n53692), .Z(n53694) );
  AND U53490 ( .A(p_input[992]), .B(n53696), .Z(n53692) );
  IV U53491 ( .A(p_input[960]), .Z(n53696) );
  XNOR U53492 ( .A(p_input[896]), .B(n53697), .Z(n53290) );
  AND U53493 ( .A(n1057), .B(n53698), .Z(n53697) );
  XOR U53494 ( .A(p_input[928]), .B(p_input[896]), .Z(n53698) );
  XOR U53495 ( .A(n53699), .B(n53700), .Z(n1057) );
  AND U53496 ( .A(n53701), .B(n53702), .Z(n53700) );
  XNOR U53497 ( .A(p_input[959]), .B(n53699), .Z(n53702) );
  XOR U53498 ( .A(n53699), .B(p_input[927]), .Z(n53701) );
  XOR U53499 ( .A(n53703), .B(n53704), .Z(n53699) );
  AND U53500 ( .A(n53705), .B(n53706), .Z(n53704) );
  XNOR U53501 ( .A(p_input[958]), .B(n53703), .Z(n53706) );
  XNOR U53502 ( .A(n53703), .B(n53305), .Z(n53705) );
  IV U53503 ( .A(p_input[926]), .Z(n53305) );
  XOR U53504 ( .A(n53707), .B(n53708), .Z(n53703) );
  AND U53505 ( .A(n53709), .B(n53710), .Z(n53708) );
  XNOR U53506 ( .A(p_input[957]), .B(n53707), .Z(n53710) );
  XNOR U53507 ( .A(n53707), .B(n53314), .Z(n53709) );
  IV U53508 ( .A(p_input[925]), .Z(n53314) );
  XOR U53509 ( .A(n53711), .B(n53712), .Z(n53707) );
  AND U53510 ( .A(n53713), .B(n53714), .Z(n53712) );
  XNOR U53511 ( .A(p_input[956]), .B(n53711), .Z(n53714) );
  XNOR U53512 ( .A(n53711), .B(n53323), .Z(n53713) );
  IV U53513 ( .A(p_input[924]), .Z(n53323) );
  XOR U53514 ( .A(n53715), .B(n53716), .Z(n53711) );
  AND U53515 ( .A(n53717), .B(n53718), .Z(n53716) );
  XNOR U53516 ( .A(p_input[955]), .B(n53715), .Z(n53718) );
  XNOR U53517 ( .A(n53715), .B(n53332), .Z(n53717) );
  IV U53518 ( .A(p_input[923]), .Z(n53332) );
  XOR U53519 ( .A(n53719), .B(n53720), .Z(n53715) );
  AND U53520 ( .A(n53721), .B(n53722), .Z(n53720) );
  XNOR U53521 ( .A(p_input[954]), .B(n53719), .Z(n53722) );
  XNOR U53522 ( .A(n53719), .B(n53341), .Z(n53721) );
  IV U53523 ( .A(p_input[922]), .Z(n53341) );
  XOR U53524 ( .A(n53723), .B(n53724), .Z(n53719) );
  AND U53525 ( .A(n53725), .B(n53726), .Z(n53724) );
  XNOR U53526 ( .A(p_input[953]), .B(n53723), .Z(n53726) );
  XNOR U53527 ( .A(n53723), .B(n53350), .Z(n53725) );
  IV U53528 ( .A(p_input[921]), .Z(n53350) );
  XOR U53529 ( .A(n53727), .B(n53728), .Z(n53723) );
  AND U53530 ( .A(n53729), .B(n53730), .Z(n53728) );
  XNOR U53531 ( .A(p_input[952]), .B(n53727), .Z(n53730) );
  XNOR U53532 ( .A(n53727), .B(n53359), .Z(n53729) );
  IV U53533 ( .A(p_input[920]), .Z(n53359) );
  XOR U53534 ( .A(n53731), .B(n53732), .Z(n53727) );
  AND U53535 ( .A(n53733), .B(n53734), .Z(n53732) );
  XNOR U53536 ( .A(p_input[951]), .B(n53731), .Z(n53734) );
  XNOR U53537 ( .A(n53731), .B(n53368), .Z(n53733) );
  IV U53538 ( .A(p_input[919]), .Z(n53368) );
  XOR U53539 ( .A(n53735), .B(n53736), .Z(n53731) );
  AND U53540 ( .A(n53737), .B(n53738), .Z(n53736) );
  XNOR U53541 ( .A(p_input[950]), .B(n53735), .Z(n53738) );
  XNOR U53542 ( .A(n53735), .B(n53377), .Z(n53737) );
  IV U53543 ( .A(p_input[918]), .Z(n53377) );
  XOR U53544 ( .A(n53739), .B(n53740), .Z(n53735) );
  AND U53545 ( .A(n53741), .B(n53742), .Z(n53740) );
  XNOR U53546 ( .A(p_input[949]), .B(n53739), .Z(n53742) );
  XNOR U53547 ( .A(n53739), .B(n53386), .Z(n53741) );
  IV U53548 ( .A(p_input[917]), .Z(n53386) );
  XOR U53549 ( .A(n53743), .B(n53744), .Z(n53739) );
  AND U53550 ( .A(n53745), .B(n53746), .Z(n53744) );
  XNOR U53551 ( .A(p_input[948]), .B(n53743), .Z(n53746) );
  XNOR U53552 ( .A(n53743), .B(n53395), .Z(n53745) );
  IV U53553 ( .A(p_input[916]), .Z(n53395) );
  XOR U53554 ( .A(n53747), .B(n53748), .Z(n53743) );
  AND U53555 ( .A(n53749), .B(n53750), .Z(n53748) );
  XNOR U53556 ( .A(p_input[947]), .B(n53747), .Z(n53750) );
  XNOR U53557 ( .A(n53747), .B(n53404), .Z(n53749) );
  IV U53558 ( .A(p_input[915]), .Z(n53404) );
  XOR U53559 ( .A(n53751), .B(n53752), .Z(n53747) );
  AND U53560 ( .A(n53753), .B(n53754), .Z(n53752) );
  XNOR U53561 ( .A(p_input[946]), .B(n53751), .Z(n53754) );
  XNOR U53562 ( .A(n53751), .B(n53413), .Z(n53753) );
  IV U53563 ( .A(p_input[914]), .Z(n53413) );
  XOR U53564 ( .A(n53755), .B(n53756), .Z(n53751) );
  AND U53565 ( .A(n53757), .B(n53758), .Z(n53756) );
  XNOR U53566 ( .A(p_input[945]), .B(n53755), .Z(n53758) );
  XNOR U53567 ( .A(n53755), .B(n53422), .Z(n53757) );
  IV U53568 ( .A(p_input[913]), .Z(n53422) );
  XOR U53569 ( .A(n53759), .B(n53760), .Z(n53755) );
  AND U53570 ( .A(n53761), .B(n53762), .Z(n53760) );
  XNOR U53571 ( .A(p_input[944]), .B(n53759), .Z(n53762) );
  XNOR U53572 ( .A(n53759), .B(n53431), .Z(n53761) );
  IV U53573 ( .A(p_input[912]), .Z(n53431) );
  XOR U53574 ( .A(n53763), .B(n53764), .Z(n53759) );
  AND U53575 ( .A(n53765), .B(n53766), .Z(n53764) );
  XNOR U53576 ( .A(p_input[943]), .B(n53763), .Z(n53766) );
  XNOR U53577 ( .A(n53763), .B(n53440), .Z(n53765) );
  IV U53578 ( .A(p_input[911]), .Z(n53440) );
  XOR U53579 ( .A(n53767), .B(n53768), .Z(n53763) );
  AND U53580 ( .A(n53769), .B(n53770), .Z(n53768) );
  XNOR U53581 ( .A(p_input[942]), .B(n53767), .Z(n53770) );
  XNOR U53582 ( .A(n53767), .B(n53449), .Z(n53769) );
  IV U53583 ( .A(p_input[910]), .Z(n53449) );
  XOR U53584 ( .A(n53771), .B(n53772), .Z(n53767) );
  AND U53585 ( .A(n53773), .B(n53774), .Z(n53772) );
  XNOR U53586 ( .A(p_input[941]), .B(n53771), .Z(n53774) );
  XNOR U53587 ( .A(n53771), .B(n53458), .Z(n53773) );
  IV U53588 ( .A(p_input[909]), .Z(n53458) );
  XOR U53589 ( .A(n53775), .B(n53776), .Z(n53771) );
  AND U53590 ( .A(n53777), .B(n53778), .Z(n53776) );
  XNOR U53591 ( .A(p_input[940]), .B(n53775), .Z(n53778) );
  XNOR U53592 ( .A(n53775), .B(n53467), .Z(n53777) );
  IV U53593 ( .A(p_input[908]), .Z(n53467) );
  XOR U53594 ( .A(n53779), .B(n53780), .Z(n53775) );
  AND U53595 ( .A(n53781), .B(n53782), .Z(n53780) );
  XNOR U53596 ( .A(p_input[939]), .B(n53779), .Z(n53782) );
  XNOR U53597 ( .A(n53779), .B(n53476), .Z(n53781) );
  IV U53598 ( .A(p_input[907]), .Z(n53476) );
  XOR U53599 ( .A(n53783), .B(n53784), .Z(n53779) );
  AND U53600 ( .A(n53785), .B(n53786), .Z(n53784) );
  XNOR U53601 ( .A(p_input[938]), .B(n53783), .Z(n53786) );
  XNOR U53602 ( .A(n53783), .B(n53485), .Z(n53785) );
  IV U53603 ( .A(p_input[906]), .Z(n53485) );
  XOR U53604 ( .A(n53787), .B(n53788), .Z(n53783) );
  AND U53605 ( .A(n53789), .B(n53790), .Z(n53788) );
  XNOR U53606 ( .A(p_input[937]), .B(n53787), .Z(n53790) );
  XNOR U53607 ( .A(n53787), .B(n53494), .Z(n53789) );
  IV U53608 ( .A(p_input[905]), .Z(n53494) );
  XOR U53609 ( .A(n53791), .B(n53792), .Z(n53787) );
  AND U53610 ( .A(n53793), .B(n53794), .Z(n53792) );
  XNOR U53611 ( .A(p_input[936]), .B(n53791), .Z(n53794) );
  XNOR U53612 ( .A(n53791), .B(n53503), .Z(n53793) );
  IV U53613 ( .A(p_input[904]), .Z(n53503) );
  XOR U53614 ( .A(n53795), .B(n53796), .Z(n53791) );
  AND U53615 ( .A(n53797), .B(n53798), .Z(n53796) );
  XNOR U53616 ( .A(p_input[935]), .B(n53795), .Z(n53798) );
  XNOR U53617 ( .A(n53795), .B(n53512), .Z(n53797) );
  IV U53618 ( .A(p_input[903]), .Z(n53512) );
  XOR U53619 ( .A(n53799), .B(n53800), .Z(n53795) );
  AND U53620 ( .A(n53801), .B(n53802), .Z(n53800) );
  XNOR U53621 ( .A(p_input[934]), .B(n53799), .Z(n53802) );
  XNOR U53622 ( .A(n53799), .B(n53521), .Z(n53801) );
  IV U53623 ( .A(p_input[902]), .Z(n53521) );
  XOR U53624 ( .A(n53803), .B(n53804), .Z(n53799) );
  AND U53625 ( .A(n53805), .B(n53806), .Z(n53804) );
  XNOR U53626 ( .A(p_input[933]), .B(n53803), .Z(n53806) );
  XNOR U53627 ( .A(n53803), .B(n53530), .Z(n53805) );
  IV U53628 ( .A(p_input[901]), .Z(n53530) );
  XOR U53629 ( .A(n53807), .B(n53808), .Z(n53803) );
  AND U53630 ( .A(n53809), .B(n53810), .Z(n53808) );
  XNOR U53631 ( .A(p_input[932]), .B(n53807), .Z(n53810) );
  XNOR U53632 ( .A(n53807), .B(n53539), .Z(n53809) );
  IV U53633 ( .A(p_input[900]), .Z(n53539) );
  XOR U53634 ( .A(n53811), .B(n53812), .Z(n53807) );
  AND U53635 ( .A(n53813), .B(n53814), .Z(n53812) );
  XNOR U53636 ( .A(p_input[931]), .B(n53811), .Z(n53814) );
  XNOR U53637 ( .A(n53811), .B(n53548), .Z(n53813) );
  IV U53638 ( .A(p_input[899]), .Z(n53548) );
  XOR U53639 ( .A(n53815), .B(n53816), .Z(n53811) );
  AND U53640 ( .A(n53817), .B(n53818), .Z(n53816) );
  XNOR U53641 ( .A(p_input[930]), .B(n53815), .Z(n53818) );
  XNOR U53642 ( .A(n53815), .B(n53557), .Z(n53817) );
  IV U53643 ( .A(p_input[898]), .Z(n53557) );
  XNOR U53644 ( .A(n53819), .B(n53820), .Z(n53815) );
  AND U53645 ( .A(n53821), .B(n53822), .Z(n53820) );
  XOR U53646 ( .A(p_input[929]), .B(n53819), .Z(n53822) );
  XNOR U53647 ( .A(p_input[897]), .B(n53819), .Z(n53821) );
  AND U53648 ( .A(p_input[928]), .B(n53823), .Z(n53819) );
  IV U53649 ( .A(p_input[896]), .Z(n53823) );
  XOR U53650 ( .A(n53824), .B(n53825), .Z(n52913) );
  AND U53651 ( .A(n649), .B(n53826), .Z(n53825) );
  XNOR U53652 ( .A(n53827), .B(n53824), .Z(n53826) );
  XOR U53653 ( .A(n53828), .B(n53829), .Z(n649) );
  AND U53654 ( .A(n53830), .B(n53831), .Z(n53829) );
  XNOR U53655 ( .A(n52928), .B(n53828), .Z(n53831) );
  AND U53656 ( .A(p_input[895]), .B(p_input[863]), .Z(n52928) );
  XNOR U53657 ( .A(n53828), .B(n52925), .Z(n53830) );
  IV U53658 ( .A(n53832), .Z(n52925) );
  AND U53659 ( .A(p_input[799]), .B(p_input[831]), .Z(n53832) );
  XOR U53660 ( .A(n53833), .B(n53834), .Z(n53828) );
  AND U53661 ( .A(n53835), .B(n53836), .Z(n53834) );
  XOR U53662 ( .A(n53833), .B(n52940), .Z(n53836) );
  XNOR U53663 ( .A(p_input[862]), .B(n53837), .Z(n52940) );
  AND U53664 ( .A(n1063), .B(n53838), .Z(n53837) );
  XOR U53665 ( .A(p_input[894]), .B(p_input[862]), .Z(n53838) );
  XNOR U53666 ( .A(n52937), .B(n53833), .Z(n53835) );
  XOR U53667 ( .A(n53839), .B(n53840), .Z(n52937) );
  AND U53668 ( .A(n1060), .B(n53841), .Z(n53840) );
  XOR U53669 ( .A(p_input[830]), .B(p_input[798]), .Z(n53841) );
  XOR U53670 ( .A(n53842), .B(n53843), .Z(n53833) );
  AND U53671 ( .A(n53844), .B(n53845), .Z(n53843) );
  XOR U53672 ( .A(n53842), .B(n52952), .Z(n53845) );
  XNOR U53673 ( .A(p_input[861]), .B(n53846), .Z(n52952) );
  AND U53674 ( .A(n1063), .B(n53847), .Z(n53846) );
  XOR U53675 ( .A(p_input[893]), .B(p_input[861]), .Z(n53847) );
  XNOR U53676 ( .A(n52949), .B(n53842), .Z(n53844) );
  XOR U53677 ( .A(n53848), .B(n53849), .Z(n52949) );
  AND U53678 ( .A(n1060), .B(n53850), .Z(n53849) );
  XOR U53679 ( .A(p_input[829]), .B(p_input[797]), .Z(n53850) );
  XOR U53680 ( .A(n53851), .B(n53852), .Z(n53842) );
  AND U53681 ( .A(n53853), .B(n53854), .Z(n53852) );
  XOR U53682 ( .A(n53851), .B(n52964), .Z(n53854) );
  XNOR U53683 ( .A(p_input[860]), .B(n53855), .Z(n52964) );
  AND U53684 ( .A(n1063), .B(n53856), .Z(n53855) );
  XOR U53685 ( .A(p_input[892]), .B(p_input[860]), .Z(n53856) );
  XNOR U53686 ( .A(n52961), .B(n53851), .Z(n53853) );
  XOR U53687 ( .A(n53857), .B(n53858), .Z(n52961) );
  AND U53688 ( .A(n1060), .B(n53859), .Z(n53858) );
  XOR U53689 ( .A(p_input[828]), .B(p_input[796]), .Z(n53859) );
  XOR U53690 ( .A(n53860), .B(n53861), .Z(n53851) );
  AND U53691 ( .A(n53862), .B(n53863), .Z(n53861) );
  XOR U53692 ( .A(n53860), .B(n52976), .Z(n53863) );
  XNOR U53693 ( .A(p_input[859]), .B(n53864), .Z(n52976) );
  AND U53694 ( .A(n1063), .B(n53865), .Z(n53864) );
  XOR U53695 ( .A(p_input[891]), .B(p_input[859]), .Z(n53865) );
  XNOR U53696 ( .A(n52973), .B(n53860), .Z(n53862) );
  XOR U53697 ( .A(n53866), .B(n53867), .Z(n52973) );
  AND U53698 ( .A(n1060), .B(n53868), .Z(n53867) );
  XOR U53699 ( .A(p_input[827]), .B(p_input[795]), .Z(n53868) );
  XOR U53700 ( .A(n53869), .B(n53870), .Z(n53860) );
  AND U53701 ( .A(n53871), .B(n53872), .Z(n53870) );
  XOR U53702 ( .A(n53869), .B(n52988), .Z(n53872) );
  XNOR U53703 ( .A(p_input[858]), .B(n53873), .Z(n52988) );
  AND U53704 ( .A(n1063), .B(n53874), .Z(n53873) );
  XOR U53705 ( .A(p_input[890]), .B(p_input[858]), .Z(n53874) );
  XNOR U53706 ( .A(n52985), .B(n53869), .Z(n53871) );
  XOR U53707 ( .A(n53875), .B(n53876), .Z(n52985) );
  AND U53708 ( .A(n1060), .B(n53877), .Z(n53876) );
  XOR U53709 ( .A(p_input[826]), .B(p_input[794]), .Z(n53877) );
  XOR U53710 ( .A(n53878), .B(n53879), .Z(n53869) );
  AND U53711 ( .A(n53880), .B(n53881), .Z(n53879) );
  XOR U53712 ( .A(n53878), .B(n53000), .Z(n53881) );
  XNOR U53713 ( .A(p_input[857]), .B(n53882), .Z(n53000) );
  AND U53714 ( .A(n1063), .B(n53883), .Z(n53882) );
  XOR U53715 ( .A(p_input[889]), .B(p_input[857]), .Z(n53883) );
  XNOR U53716 ( .A(n52997), .B(n53878), .Z(n53880) );
  XOR U53717 ( .A(n53884), .B(n53885), .Z(n52997) );
  AND U53718 ( .A(n1060), .B(n53886), .Z(n53885) );
  XOR U53719 ( .A(p_input[825]), .B(p_input[793]), .Z(n53886) );
  XOR U53720 ( .A(n53887), .B(n53888), .Z(n53878) );
  AND U53721 ( .A(n53889), .B(n53890), .Z(n53888) );
  XOR U53722 ( .A(n53887), .B(n53012), .Z(n53890) );
  XNOR U53723 ( .A(p_input[856]), .B(n53891), .Z(n53012) );
  AND U53724 ( .A(n1063), .B(n53892), .Z(n53891) );
  XOR U53725 ( .A(p_input[888]), .B(p_input[856]), .Z(n53892) );
  XNOR U53726 ( .A(n53009), .B(n53887), .Z(n53889) );
  XOR U53727 ( .A(n53893), .B(n53894), .Z(n53009) );
  AND U53728 ( .A(n1060), .B(n53895), .Z(n53894) );
  XOR U53729 ( .A(p_input[824]), .B(p_input[792]), .Z(n53895) );
  XOR U53730 ( .A(n53896), .B(n53897), .Z(n53887) );
  AND U53731 ( .A(n53898), .B(n53899), .Z(n53897) );
  XOR U53732 ( .A(n53896), .B(n53024), .Z(n53899) );
  XNOR U53733 ( .A(p_input[855]), .B(n53900), .Z(n53024) );
  AND U53734 ( .A(n1063), .B(n53901), .Z(n53900) );
  XOR U53735 ( .A(p_input[887]), .B(p_input[855]), .Z(n53901) );
  XNOR U53736 ( .A(n53021), .B(n53896), .Z(n53898) );
  XOR U53737 ( .A(n53902), .B(n53903), .Z(n53021) );
  AND U53738 ( .A(n1060), .B(n53904), .Z(n53903) );
  XOR U53739 ( .A(p_input[823]), .B(p_input[791]), .Z(n53904) );
  XOR U53740 ( .A(n53905), .B(n53906), .Z(n53896) );
  AND U53741 ( .A(n53907), .B(n53908), .Z(n53906) );
  XOR U53742 ( .A(n53905), .B(n53036), .Z(n53908) );
  XNOR U53743 ( .A(p_input[854]), .B(n53909), .Z(n53036) );
  AND U53744 ( .A(n1063), .B(n53910), .Z(n53909) );
  XOR U53745 ( .A(p_input[886]), .B(p_input[854]), .Z(n53910) );
  XNOR U53746 ( .A(n53033), .B(n53905), .Z(n53907) );
  XOR U53747 ( .A(n53911), .B(n53912), .Z(n53033) );
  AND U53748 ( .A(n1060), .B(n53913), .Z(n53912) );
  XOR U53749 ( .A(p_input[822]), .B(p_input[790]), .Z(n53913) );
  XOR U53750 ( .A(n53914), .B(n53915), .Z(n53905) );
  AND U53751 ( .A(n53916), .B(n53917), .Z(n53915) );
  XOR U53752 ( .A(n53914), .B(n53048), .Z(n53917) );
  XNOR U53753 ( .A(p_input[853]), .B(n53918), .Z(n53048) );
  AND U53754 ( .A(n1063), .B(n53919), .Z(n53918) );
  XOR U53755 ( .A(p_input[885]), .B(p_input[853]), .Z(n53919) );
  XNOR U53756 ( .A(n53045), .B(n53914), .Z(n53916) );
  XOR U53757 ( .A(n53920), .B(n53921), .Z(n53045) );
  AND U53758 ( .A(n1060), .B(n53922), .Z(n53921) );
  XOR U53759 ( .A(p_input[821]), .B(p_input[789]), .Z(n53922) );
  XOR U53760 ( .A(n53923), .B(n53924), .Z(n53914) );
  AND U53761 ( .A(n53925), .B(n53926), .Z(n53924) );
  XOR U53762 ( .A(n53923), .B(n53060), .Z(n53926) );
  XNOR U53763 ( .A(p_input[852]), .B(n53927), .Z(n53060) );
  AND U53764 ( .A(n1063), .B(n53928), .Z(n53927) );
  XOR U53765 ( .A(p_input[884]), .B(p_input[852]), .Z(n53928) );
  XNOR U53766 ( .A(n53057), .B(n53923), .Z(n53925) );
  XOR U53767 ( .A(n53929), .B(n53930), .Z(n53057) );
  AND U53768 ( .A(n1060), .B(n53931), .Z(n53930) );
  XOR U53769 ( .A(p_input[820]), .B(p_input[788]), .Z(n53931) );
  XOR U53770 ( .A(n53932), .B(n53933), .Z(n53923) );
  AND U53771 ( .A(n53934), .B(n53935), .Z(n53933) );
  XOR U53772 ( .A(n53932), .B(n53072), .Z(n53935) );
  XNOR U53773 ( .A(p_input[851]), .B(n53936), .Z(n53072) );
  AND U53774 ( .A(n1063), .B(n53937), .Z(n53936) );
  XOR U53775 ( .A(p_input[883]), .B(p_input[851]), .Z(n53937) );
  XNOR U53776 ( .A(n53069), .B(n53932), .Z(n53934) );
  XOR U53777 ( .A(n53938), .B(n53939), .Z(n53069) );
  AND U53778 ( .A(n1060), .B(n53940), .Z(n53939) );
  XOR U53779 ( .A(p_input[819]), .B(p_input[787]), .Z(n53940) );
  XOR U53780 ( .A(n53941), .B(n53942), .Z(n53932) );
  AND U53781 ( .A(n53943), .B(n53944), .Z(n53942) );
  XOR U53782 ( .A(n53941), .B(n53084), .Z(n53944) );
  XNOR U53783 ( .A(p_input[850]), .B(n53945), .Z(n53084) );
  AND U53784 ( .A(n1063), .B(n53946), .Z(n53945) );
  XOR U53785 ( .A(p_input[882]), .B(p_input[850]), .Z(n53946) );
  XNOR U53786 ( .A(n53081), .B(n53941), .Z(n53943) );
  XOR U53787 ( .A(n53947), .B(n53948), .Z(n53081) );
  AND U53788 ( .A(n1060), .B(n53949), .Z(n53948) );
  XOR U53789 ( .A(p_input[818]), .B(p_input[786]), .Z(n53949) );
  XOR U53790 ( .A(n53950), .B(n53951), .Z(n53941) );
  AND U53791 ( .A(n53952), .B(n53953), .Z(n53951) );
  XOR U53792 ( .A(n53950), .B(n53096), .Z(n53953) );
  XNOR U53793 ( .A(p_input[849]), .B(n53954), .Z(n53096) );
  AND U53794 ( .A(n1063), .B(n53955), .Z(n53954) );
  XOR U53795 ( .A(p_input[881]), .B(p_input[849]), .Z(n53955) );
  XNOR U53796 ( .A(n53093), .B(n53950), .Z(n53952) );
  XOR U53797 ( .A(n53956), .B(n53957), .Z(n53093) );
  AND U53798 ( .A(n1060), .B(n53958), .Z(n53957) );
  XOR U53799 ( .A(p_input[817]), .B(p_input[785]), .Z(n53958) );
  XOR U53800 ( .A(n53959), .B(n53960), .Z(n53950) );
  AND U53801 ( .A(n53961), .B(n53962), .Z(n53960) );
  XOR U53802 ( .A(n53959), .B(n53108), .Z(n53962) );
  XNOR U53803 ( .A(p_input[848]), .B(n53963), .Z(n53108) );
  AND U53804 ( .A(n1063), .B(n53964), .Z(n53963) );
  XOR U53805 ( .A(p_input[880]), .B(p_input[848]), .Z(n53964) );
  XNOR U53806 ( .A(n53105), .B(n53959), .Z(n53961) );
  XOR U53807 ( .A(n53965), .B(n53966), .Z(n53105) );
  AND U53808 ( .A(n1060), .B(n53967), .Z(n53966) );
  XOR U53809 ( .A(p_input[816]), .B(p_input[784]), .Z(n53967) );
  XOR U53810 ( .A(n53968), .B(n53969), .Z(n53959) );
  AND U53811 ( .A(n53970), .B(n53971), .Z(n53969) );
  XOR U53812 ( .A(n53968), .B(n53120), .Z(n53971) );
  XNOR U53813 ( .A(p_input[847]), .B(n53972), .Z(n53120) );
  AND U53814 ( .A(n1063), .B(n53973), .Z(n53972) );
  XOR U53815 ( .A(p_input[879]), .B(p_input[847]), .Z(n53973) );
  XNOR U53816 ( .A(n53117), .B(n53968), .Z(n53970) );
  XOR U53817 ( .A(n53974), .B(n53975), .Z(n53117) );
  AND U53818 ( .A(n1060), .B(n53976), .Z(n53975) );
  XOR U53819 ( .A(p_input[815]), .B(p_input[783]), .Z(n53976) );
  XOR U53820 ( .A(n53977), .B(n53978), .Z(n53968) );
  AND U53821 ( .A(n53979), .B(n53980), .Z(n53978) );
  XOR U53822 ( .A(n53977), .B(n53132), .Z(n53980) );
  XNOR U53823 ( .A(p_input[846]), .B(n53981), .Z(n53132) );
  AND U53824 ( .A(n1063), .B(n53982), .Z(n53981) );
  XOR U53825 ( .A(p_input[878]), .B(p_input[846]), .Z(n53982) );
  XNOR U53826 ( .A(n53129), .B(n53977), .Z(n53979) );
  XOR U53827 ( .A(n53983), .B(n53984), .Z(n53129) );
  AND U53828 ( .A(n1060), .B(n53985), .Z(n53984) );
  XOR U53829 ( .A(p_input[814]), .B(p_input[782]), .Z(n53985) );
  XOR U53830 ( .A(n53986), .B(n53987), .Z(n53977) );
  AND U53831 ( .A(n53988), .B(n53989), .Z(n53987) );
  XOR U53832 ( .A(n53986), .B(n53144), .Z(n53989) );
  XNOR U53833 ( .A(p_input[845]), .B(n53990), .Z(n53144) );
  AND U53834 ( .A(n1063), .B(n53991), .Z(n53990) );
  XOR U53835 ( .A(p_input[877]), .B(p_input[845]), .Z(n53991) );
  XNOR U53836 ( .A(n53141), .B(n53986), .Z(n53988) );
  XOR U53837 ( .A(n53992), .B(n53993), .Z(n53141) );
  AND U53838 ( .A(n1060), .B(n53994), .Z(n53993) );
  XOR U53839 ( .A(p_input[813]), .B(p_input[781]), .Z(n53994) );
  XOR U53840 ( .A(n53995), .B(n53996), .Z(n53986) );
  AND U53841 ( .A(n53997), .B(n53998), .Z(n53996) );
  XOR U53842 ( .A(n53995), .B(n53156), .Z(n53998) );
  XNOR U53843 ( .A(p_input[844]), .B(n53999), .Z(n53156) );
  AND U53844 ( .A(n1063), .B(n54000), .Z(n53999) );
  XOR U53845 ( .A(p_input[876]), .B(p_input[844]), .Z(n54000) );
  XNOR U53846 ( .A(n53153), .B(n53995), .Z(n53997) );
  XOR U53847 ( .A(n54001), .B(n54002), .Z(n53153) );
  AND U53848 ( .A(n1060), .B(n54003), .Z(n54002) );
  XOR U53849 ( .A(p_input[812]), .B(p_input[780]), .Z(n54003) );
  XOR U53850 ( .A(n54004), .B(n54005), .Z(n53995) );
  AND U53851 ( .A(n54006), .B(n54007), .Z(n54005) );
  XOR U53852 ( .A(n54004), .B(n53168), .Z(n54007) );
  XNOR U53853 ( .A(p_input[843]), .B(n54008), .Z(n53168) );
  AND U53854 ( .A(n1063), .B(n54009), .Z(n54008) );
  XOR U53855 ( .A(p_input[875]), .B(p_input[843]), .Z(n54009) );
  XNOR U53856 ( .A(n53165), .B(n54004), .Z(n54006) );
  XOR U53857 ( .A(n54010), .B(n54011), .Z(n53165) );
  AND U53858 ( .A(n1060), .B(n54012), .Z(n54011) );
  XOR U53859 ( .A(p_input[811]), .B(p_input[779]), .Z(n54012) );
  XOR U53860 ( .A(n54013), .B(n54014), .Z(n54004) );
  AND U53861 ( .A(n54015), .B(n54016), .Z(n54014) );
  XOR U53862 ( .A(n54013), .B(n53180), .Z(n54016) );
  XNOR U53863 ( .A(p_input[842]), .B(n54017), .Z(n53180) );
  AND U53864 ( .A(n1063), .B(n54018), .Z(n54017) );
  XOR U53865 ( .A(p_input[874]), .B(p_input[842]), .Z(n54018) );
  XNOR U53866 ( .A(n53177), .B(n54013), .Z(n54015) );
  XOR U53867 ( .A(n54019), .B(n54020), .Z(n53177) );
  AND U53868 ( .A(n1060), .B(n54021), .Z(n54020) );
  XOR U53869 ( .A(p_input[810]), .B(p_input[778]), .Z(n54021) );
  XOR U53870 ( .A(n54022), .B(n54023), .Z(n54013) );
  AND U53871 ( .A(n54024), .B(n54025), .Z(n54023) );
  XOR U53872 ( .A(n54022), .B(n53192), .Z(n54025) );
  XNOR U53873 ( .A(p_input[841]), .B(n54026), .Z(n53192) );
  AND U53874 ( .A(n1063), .B(n54027), .Z(n54026) );
  XOR U53875 ( .A(p_input[873]), .B(p_input[841]), .Z(n54027) );
  XNOR U53876 ( .A(n53189), .B(n54022), .Z(n54024) );
  XOR U53877 ( .A(n54028), .B(n54029), .Z(n53189) );
  AND U53878 ( .A(n1060), .B(n54030), .Z(n54029) );
  XOR U53879 ( .A(p_input[809]), .B(p_input[777]), .Z(n54030) );
  XOR U53880 ( .A(n54031), .B(n54032), .Z(n54022) );
  AND U53881 ( .A(n54033), .B(n54034), .Z(n54032) );
  XOR U53882 ( .A(n54031), .B(n53204), .Z(n54034) );
  XNOR U53883 ( .A(p_input[840]), .B(n54035), .Z(n53204) );
  AND U53884 ( .A(n1063), .B(n54036), .Z(n54035) );
  XOR U53885 ( .A(p_input[872]), .B(p_input[840]), .Z(n54036) );
  XNOR U53886 ( .A(n53201), .B(n54031), .Z(n54033) );
  XOR U53887 ( .A(n54037), .B(n54038), .Z(n53201) );
  AND U53888 ( .A(n1060), .B(n54039), .Z(n54038) );
  XOR U53889 ( .A(p_input[808]), .B(p_input[776]), .Z(n54039) );
  XOR U53890 ( .A(n54040), .B(n54041), .Z(n54031) );
  AND U53891 ( .A(n54042), .B(n54043), .Z(n54041) );
  XOR U53892 ( .A(n54040), .B(n53216), .Z(n54043) );
  XNOR U53893 ( .A(p_input[839]), .B(n54044), .Z(n53216) );
  AND U53894 ( .A(n1063), .B(n54045), .Z(n54044) );
  XOR U53895 ( .A(p_input[871]), .B(p_input[839]), .Z(n54045) );
  XNOR U53896 ( .A(n53213), .B(n54040), .Z(n54042) );
  XOR U53897 ( .A(n54046), .B(n54047), .Z(n53213) );
  AND U53898 ( .A(n1060), .B(n54048), .Z(n54047) );
  XOR U53899 ( .A(p_input[807]), .B(p_input[775]), .Z(n54048) );
  XOR U53900 ( .A(n54049), .B(n54050), .Z(n54040) );
  AND U53901 ( .A(n54051), .B(n54052), .Z(n54050) );
  XOR U53902 ( .A(n54049), .B(n53228), .Z(n54052) );
  XNOR U53903 ( .A(p_input[838]), .B(n54053), .Z(n53228) );
  AND U53904 ( .A(n1063), .B(n54054), .Z(n54053) );
  XOR U53905 ( .A(p_input[870]), .B(p_input[838]), .Z(n54054) );
  XNOR U53906 ( .A(n53225), .B(n54049), .Z(n54051) );
  XOR U53907 ( .A(n54055), .B(n54056), .Z(n53225) );
  AND U53908 ( .A(n1060), .B(n54057), .Z(n54056) );
  XOR U53909 ( .A(p_input[806]), .B(p_input[774]), .Z(n54057) );
  XOR U53910 ( .A(n54058), .B(n54059), .Z(n54049) );
  AND U53911 ( .A(n54060), .B(n54061), .Z(n54059) );
  XOR U53912 ( .A(n54058), .B(n53240), .Z(n54061) );
  XNOR U53913 ( .A(p_input[837]), .B(n54062), .Z(n53240) );
  AND U53914 ( .A(n1063), .B(n54063), .Z(n54062) );
  XOR U53915 ( .A(p_input[869]), .B(p_input[837]), .Z(n54063) );
  XNOR U53916 ( .A(n53237), .B(n54058), .Z(n54060) );
  XOR U53917 ( .A(n54064), .B(n54065), .Z(n53237) );
  AND U53918 ( .A(n1060), .B(n54066), .Z(n54065) );
  XOR U53919 ( .A(p_input[805]), .B(p_input[773]), .Z(n54066) );
  XOR U53920 ( .A(n54067), .B(n54068), .Z(n54058) );
  AND U53921 ( .A(n54069), .B(n54070), .Z(n54068) );
  XOR U53922 ( .A(n54067), .B(n53252), .Z(n54070) );
  XNOR U53923 ( .A(p_input[836]), .B(n54071), .Z(n53252) );
  AND U53924 ( .A(n1063), .B(n54072), .Z(n54071) );
  XOR U53925 ( .A(p_input[868]), .B(p_input[836]), .Z(n54072) );
  XNOR U53926 ( .A(n53249), .B(n54067), .Z(n54069) );
  XOR U53927 ( .A(n54073), .B(n54074), .Z(n53249) );
  AND U53928 ( .A(n1060), .B(n54075), .Z(n54074) );
  XOR U53929 ( .A(p_input[804]), .B(p_input[772]), .Z(n54075) );
  XOR U53930 ( .A(n54076), .B(n54077), .Z(n54067) );
  AND U53931 ( .A(n54078), .B(n54079), .Z(n54077) );
  XOR U53932 ( .A(n54076), .B(n53264), .Z(n54079) );
  XNOR U53933 ( .A(p_input[835]), .B(n54080), .Z(n53264) );
  AND U53934 ( .A(n1063), .B(n54081), .Z(n54080) );
  XOR U53935 ( .A(p_input[867]), .B(p_input[835]), .Z(n54081) );
  XNOR U53936 ( .A(n53261), .B(n54076), .Z(n54078) );
  XOR U53937 ( .A(n54082), .B(n54083), .Z(n53261) );
  AND U53938 ( .A(n1060), .B(n54084), .Z(n54083) );
  XOR U53939 ( .A(p_input[803]), .B(p_input[771]), .Z(n54084) );
  XOR U53940 ( .A(n54085), .B(n54086), .Z(n54076) );
  AND U53941 ( .A(n54087), .B(n54088), .Z(n54086) );
  XOR U53942 ( .A(n54085), .B(n53276), .Z(n54088) );
  XNOR U53943 ( .A(p_input[834]), .B(n54089), .Z(n53276) );
  AND U53944 ( .A(n1063), .B(n54090), .Z(n54089) );
  XOR U53945 ( .A(p_input[866]), .B(p_input[834]), .Z(n54090) );
  XNOR U53946 ( .A(n53273), .B(n54085), .Z(n54087) );
  XOR U53947 ( .A(n54091), .B(n54092), .Z(n53273) );
  AND U53948 ( .A(n1060), .B(n54093), .Z(n54092) );
  XOR U53949 ( .A(p_input[802]), .B(p_input[770]), .Z(n54093) );
  XOR U53950 ( .A(n54094), .B(n54095), .Z(n54085) );
  AND U53951 ( .A(n54096), .B(n54097), .Z(n54095) );
  XNOR U53952 ( .A(n54098), .B(n53289), .Z(n54097) );
  XNOR U53953 ( .A(p_input[833]), .B(n54099), .Z(n53289) );
  AND U53954 ( .A(n1063), .B(n54100), .Z(n54099) );
  XNOR U53955 ( .A(p_input[865]), .B(n54101), .Z(n54100) );
  IV U53956 ( .A(p_input[833]), .Z(n54101) );
  XNOR U53957 ( .A(n53286), .B(n54094), .Z(n54096) );
  XNOR U53958 ( .A(p_input[769]), .B(n54102), .Z(n53286) );
  AND U53959 ( .A(n1060), .B(n54103), .Z(n54102) );
  XOR U53960 ( .A(p_input[801]), .B(p_input[769]), .Z(n54103) );
  IV U53961 ( .A(n54098), .Z(n54094) );
  AND U53962 ( .A(n53824), .B(n53827), .Z(n54098) );
  XOR U53963 ( .A(p_input[832]), .B(n54104), .Z(n53827) );
  AND U53964 ( .A(n1063), .B(n54105), .Z(n54104) );
  XOR U53965 ( .A(p_input[864]), .B(p_input[832]), .Z(n54105) );
  XOR U53966 ( .A(n54106), .B(n54107), .Z(n1063) );
  AND U53967 ( .A(n54108), .B(n54109), .Z(n54107) );
  XNOR U53968 ( .A(p_input[895]), .B(n54106), .Z(n54109) );
  XOR U53969 ( .A(n54106), .B(p_input[863]), .Z(n54108) );
  XOR U53970 ( .A(n54110), .B(n54111), .Z(n54106) );
  AND U53971 ( .A(n54112), .B(n54113), .Z(n54111) );
  XNOR U53972 ( .A(p_input[894]), .B(n54110), .Z(n54113) );
  XOR U53973 ( .A(n54110), .B(p_input[862]), .Z(n54112) );
  XOR U53974 ( .A(n54114), .B(n54115), .Z(n54110) );
  AND U53975 ( .A(n54116), .B(n54117), .Z(n54115) );
  XNOR U53976 ( .A(p_input[893]), .B(n54114), .Z(n54117) );
  XOR U53977 ( .A(n54114), .B(p_input[861]), .Z(n54116) );
  XOR U53978 ( .A(n54118), .B(n54119), .Z(n54114) );
  AND U53979 ( .A(n54120), .B(n54121), .Z(n54119) );
  XNOR U53980 ( .A(p_input[892]), .B(n54118), .Z(n54121) );
  XOR U53981 ( .A(n54118), .B(p_input[860]), .Z(n54120) );
  XOR U53982 ( .A(n54122), .B(n54123), .Z(n54118) );
  AND U53983 ( .A(n54124), .B(n54125), .Z(n54123) );
  XNOR U53984 ( .A(p_input[891]), .B(n54122), .Z(n54125) );
  XOR U53985 ( .A(n54122), .B(p_input[859]), .Z(n54124) );
  XOR U53986 ( .A(n54126), .B(n54127), .Z(n54122) );
  AND U53987 ( .A(n54128), .B(n54129), .Z(n54127) );
  XNOR U53988 ( .A(p_input[890]), .B(n54126), .Z(n54129) );
  XOR U53989 ( .A(n54126), .B(p_input[858]), .Z(n54128) );
  XOR U53990 ( .A(n54130), .B(n54131), .Z(n54126) );
  AND U53991 ( .A(n54132), .B(n54133), .Z(n54131) );
  XNOR U53992 ( .A(p_input[889]), .B(n54130), .Z(n54133) );
  XOR U53993 ( .A(n54130), .B(p_input[857]), .Z(n54132) );
  XOR U53994 ( .A(n54134), .B(n54135), .Z(n54130) );
  AND U53995 ( .A(n54136), .B(n54137), .Z(n54135) );
  XNOR U53996 ( .A(p_input[888]), .B(n54134), .Z(n54137) );
  XOR U53997 ( .A(n54134), .B(p_input[856]), .Z(n54136) );
  XOR U53998 ( .A(n54138), .B(n54139), .Z(n54134) );
  AND U53999 ( .A(n54140), .B(n54141), .Z(n54139) );
  XNOR U54000 ( .A(p_input[887]), .B(n54138), .Z(n54141) );
  XOR U54001 ( .A(n54138), .B(p_input[855]), .Z(n54140) );
  XOR U54002 ( .A(n54142), .B(n54143), .Z(n54138) );
  AND U54003 ( .A(n54144), .B(n54145), .Z(n54143) );
  XNOR U54004 ( .A(p_input[886]), .B(n54142), .Z(n54145) );
  XOR U54005 ( .A(n54142), .B(p_input[854]), .Z(n54144) );
  XOR U54006 ( .A(n54146), .B(n54147), .Z(n54142) );
  AND U54007 ( .A(n54148), .B(n54149), .Z(n54147) );
  XNOR U54008 ( .A(p_input[885]), .B(n54146), .Z(n54149) );
  XOR U54009 ( .A(n54146), .B(p_input[853]), .Z(n54148) );
  XOR U54010 ( .A(n54150), .B(n54151), .Z(n54146) );
  AND U54011 ( .A(n54152), .B(n54153), .Z(n54151) );
  XNOR U54012 ( .A(p_input[884]), .B(n54150), .Z(n54153) );
  XOR U54013 ( .A(n54150), .B(p_input[852]), .Z(n54152) );
  XOR U54014 ( .A(n54154), .B(n54155), .Z(n54150) );
  AND U54015 ( .A(n54156), .B(n54157), .Z(n54155) );
  XNOR U54016 ( .A(p_input[883]), .B(n54154), .Z(n54157) );
  XOR U54017 ( .A(n54154), .B(p_input[851]), .Z(n54156) );
  XOR U54018 ( .A(n54158), .B(n54159), .Z(n54154) );
  AND U54019 ( .A(n54160), .B(n54161), .Z(n54159) );
  XNOR U54020 ( .A(p_input[882]), .B(n54158), .Z(n54161) );
  XOR U54021 ( .A(n54158), .B(p_input[850]), .Z(n54160) );
  XOR U54022 ( .A(n54162), .B(n54163), .Z(n54158) );
  AND U54023 ( .A(n54164), .B(n54165), .Z(n54163) );
  XNOR U54024 ( .A(p_input[881]), .B(n54162), .Z(n54165) );
  XOR U54025 ( .A(n54162), .B(p_input[849]), .Z(n54164) );
  XOR U54026 ( .A(n54166), .B(n54167), .Z(n54162) );
  AND U54027 ( .A(n54168), .B(n54169), .Z(n54167) );
  XNOR U54028 ( .A(p_input[880]), .B(n54166), .Z(n54169) );
  XOR U54029 ( .A(n54166), .B(p_input[848]), .Z(n54168) );
  XOR U54030 ( .A(n54170), .B(n54171), .Z(n54166) );
  AND U54031 ( .A(n54172), .B(n54173), .Z(n54171) );
  XNOR U54032 ( .A(p_input[879]), .B(n54170), .Z(n54173) );
  XOR U54033 ( .A(n54170), .B(p_input[847]), .Z(n54172) );
  XOR U54034 ( .A(n54174), .B(n54175), .Z(n54170) );
  AND U54035 ( .A(n54176), .B(n54177), .Z(n54175) );
  XNOR U54036 ( .A(p_input[878]), .B(n54174), .Z(n54177) );
  XOR U54037 ( .A(n54174), .B(p_input[846]), .Z(n54176) );
  XOR U54038 ( .A(n54178), .B(n54179), .Z(n54174) );
  AND U54039 ( .A(n54180), .B(n54181), .Z(n54179) );
  XNOR U54040 ( .A(p_input[877]), .B(n54178), .Z(n54181) );
  XOR U54041 ( .A(n54178), .B(p_input[845]), .Z(n54180) );
  XOR U54042 ( .A(n54182), .B(n54183), .Z(n54178) );
  AND U54043 ( .A(n54184), .B(n54185), .Z(n54183) );
  XNOR U54044 ( .A(p_input[876]), .B(n54182), .Z(n54185) );
  XOR U54045 ( .A(n54182), .B(p_input[844]), .Z(n54184) );
  XOR U54046 ( .A(n54186), .B(n54187), .Z(n54182) );
  AND U54047 ( .A(n54188), .B(n54189), .Z(n54187) );
  XNOR U54048 ( .A(p_input[875]), .B(n54186), .Z(n54189) );
  XOR U54049 ( .A(n54186), .B(p_input[843]), .Z(n54188) );
  XOR U54050 ( .A(n54190), .B(n54191), .Z(n54186) );
  AND U54051 ( .A(n54192), .B(n54193), .Z(n54191) );
  XNOR U54052 ( .A(p_input[874]), .B(n54190), .Z(n54193) );
  XOR U54053 ( .A(n54190), .B(p_input[842]), .Z(n54192) );
  XOR U54054 ( .A(n54194), .B(n54195), .Z(n54190) );
  AND U54055 ( .A(n54196), .B(n54197), .Z(n54195) );
  XNOR U54056 ( .A(p_input[873]), .B(n54194), .Z(n54197) );
  XOR U54057 ( .A(n54194), .B(p_input[841]), .Z(n54196) );
  XOR U54058 ( .A(n54198), .B(n54199), .Z(n54194) );
  AND U54059 ( .A(n54200), .B(n54201), .Z(n54199) );
  XNOR U54060 ( .A(p_input[872]), .B(n54198), .Z(n54201) );
  XOR U54061 ( .A(n54198), .B(p_input[840]), .Z(n54200) );
  XOR U54062 ( .A(n54202), .B(n54203), .Z(n54198) );
  AND U54063 ( .A(n54204), .B(n54205), .Z(n54203) );
  XNOR U54064 ( .A(p_input[871]), .B(n54202), .Z(n54205) );
  XOR U54065 ( .A(n54202), .B(p_input[839]), .Z(n54204) );
  XOR U54066 ( .A(n54206), .B(n54207), .Z(n54202) );
  AND U54067 ( .A(n54208), .B(n54209), .Z(n54207) );
  XNOR U54068 ( .A(p_input[870]), .B(n54206), .Z(n54209) );
  XOR U54069 ( .A(n54206), .B(p_input[838]), .Z(n54208) );
  XOR U54070 ( .A(n54210), .B(n54211), .Z(n54206) );
  AND U54071 ( .A(n54212), .B(n54213), .Z(n54211) );
  XNOR U54072 ( .A(p_input[869]), .B(n54210), .Z(n54213) );
  XOR U54073 ( .A(n54210), .B(p_input[837]), .Z(n54212) );
  XOR U54074 ( .A(n54214), .B(n54215), .Z(n54210) );
  AND U54075 ( .A(n54216), .B(n54217), .Z(n54215) );
  XNOR U54076 ( .A(p_input[868]), .B(n54214), .Z(n54217) );
  XOR U54077 ( .A(n54214), .B(p_input[836]), .Z(n54216) );
  XOR U54078 ( .A(n54218), .B(n54219), .Z(n54214) );
  AND U54079 ( .A(n54220), .B(n54221), .Z(n54219) );
  XNOR U54080 ( .A(p_input[867]), .B(n54218), .Z(n54221) );
  XOR U54081 ( .A(n54218), .B(p_input[835]), .Z(n54220) );
  XOR U54082 ( .A(n54222), .B(n54223), .Z(n54218) );
  AND U54083 ( .A(n54224), .B(n54225), .Z(n54223) );
  XNOR U54084 ( .A(p_input[866]), .B(n54222), .Z(n54225) );
  XOR U54085 ( .A(n54222), .B(p_input[834]), .Z(n54224) );
  XNOR U54086 ( .A(n54226), .B(n54227), .Z(n54222) );
  AND U54087 ( .A(n54228), .B(n54229), .Z(n54227) );
  XOR U54088 ( .A(p_input[865]), .B(n54226), .Z(n54229) );
  XNOR U54089 ( .A(p_input[833]), .B(n54226), .Z(n54228) );
  AND U54090 ( .A(p_input[864]), .B(n54230), .Z(n54226) );
  IV U54091 ( .A(p_input[832]), .Z(n54230) );
  XNOR U54092 ( .A(p_input[768]), .B(n54231), .Z(n53824) );
  AND U54093 ( .A(n1060), .B(n54232), .Z(n54231) );
  XOR U54094 ( .A(p_input[800]), .B(p_input[768]), .Z(n54232) );
  XOR U54095 ( .A(n54233), .B(n54234), .Z(n1060) );
  AND U54096 ( .A(n54235), .B(n54236), .Z(n54234) );
  XNOR U54097 ( .A(p_input[831]), .B(n54233), .Z(n54236) );
  XOR U54098 ( .A(n54233), .B(p_input[799]), .Z(n54235) );
  XOR U54099 ( .A(n54237), .B(n54238), .Z(n54233) );
  AND U54100 ( .A(n54239), .B(n54240), .Z(n54238) );
  XNOR U54101 ( .A(p_input[830]), .B(n54237), .Z(n54240) );
  XNOR U54102 ( .A(n54237), .B(n53839), .Z(n54239) );
  IV U54103 ( .A(p_input[798]), .Z(n53839) );
  XOR U54104 ( .A(n54241), .B(n54242), .Z(n54237) );
  AND U54105 ( .A(n54243), .B(n54244), .Z(n54242) );
  XNOR U54106 ( .A(p_input[829]), .B(n54241), .Z(n54244) );
  XNOR U54107 ( .A(n54241), .B(n53848), .Z(n54243) );
  IV U54108 ( .A(p_input[797]), .Z(n53848) );
  XOR U54109 ( .A(n54245), .B(n54246), .Z(n54241) );
  AND U54110 ( .A(n54247), .B(n54248), .Z(n54246) );
  XNOR U54111 ( .A(p_input[828]), .B(n54245), .Z(n54248) );
  XNOR U54112 ( .A(n54245), .B(n53857), .Z(n54247) );
  IV U54113 ( .A(p_input[796]), .Z(n53857) );
  XOR U54114 ( .A(n54249), .B(n54250), .Z(n54245) );
  AND U54115 ( .A(n54251), .B(n54252), .Z(n54250) );
  XNOR U54116 ( .A(p_input[827]), .B(n54249), .Z(n54252) );
  XNOR U54117 ( .A(n54249), .B(n53866), .Z(n54251) );
  IV U54118 ( .A(p_input[795]), .Z(n53866) );
  XOR U54119 ( .A(n54253), .B(n54254), .Z(n54249) );
  AND U54120 ( .A(n54255), .B(n54256), .Z(n54254) );
  XNOR U54121 ( .A(p_input[826]), .B(n54253), .Z(n54256) );
  XNOR U54122 ( .A(n54253), .B(n53875), .Z(n54255) );
  IV U54123 ( .A(p_input[794]), .Z(n53875) );
  XOR U54124 ( .A(n54257), .B(n54258), .Z(n54253) );
  AND U54125 ( .A(n54259), .B(n54260), .Z(n54258) );
  XNOR U54126 ( .A(p_input[825]), .B(n54257), .Z(n54260) );
  XNOR U54127 ( .A(n54257), .B(n53884), .Z(n54259) );
  IV U54128 ( .A(p_input[793]), .Z(n53884) );
  XOR U54129 ( .A(n54261), .B(n54262), .Z(n54257) );
  AND U54130 ( .A(n54263), .B(n54264), .Z(n54262) );
  XNOR U54131 ( .A(p_input[824]), .B(n54261), .Z(n54264) );
  XNOR U54132 ( .A(n54261), .B(n53893), .Z(n54263) );
  IV U54133 ( .A(p_input[792]), .Z(n53893) );
  XOR U54134 ( .A(n54265), .B(n54266), .Z(n54261) );
  AND U54135 ( .A(n54267), .B(n54268), .Z(n54266) );
  XNOR U54136 ( .A(p_input[823]), .B(n54265), .Z(n54268) );
  XNOR U54137 ( .A(n54265), .B(n53902), .Z(n54267) );
  IV U54138 ( .A(p_input[791]), .Z(n53902) );
  XOR U54139 ( .A(n54269), .B(n54270), .Z(n54265) );
  AND U54140 ( .A(n54271), .B(n54272), .Z(n54270) );
  XNOR U54141 ( .A(p_input[822]), .B(n54269), .Z(n54272) );
  XNOR U54142 ( .A(n54269), .B(n53911), .Z(n54271) );
  IV U54143 ( .A(p_input[790]), .Z(n53911) );
  XOR U54144 ( .A(n54273), .B(n54274), .Z(n54269) );
  AND U54145 ( .A(n54275), .B(n54276), .Z(n54274) );
  XNOR U54146 ( .A(p_input[821]), .B(n54273), .Z(n54276) );
  XNOR U54147 ( .A(n54273), .B(n53920), .Z(n54275) );
  IV U54148 ( .A(p_input[789]), .Z(n53920) );
  XOR U54149 ( .A(n54277), .B(n54278), .Z(n54273) );
  AND U54150 ( .A(n54279), .B(n54280), .Z(n54278) );
  XNOR U54151 ( .A(p_input[820]), .B(n54277), .Z(n54280) );
  XNOR U54152 ( .A(n54277), .B(n53929), .Z(n54279) );
  IV U54153 ( .A(p_input[788]), .Z(n53929) );
  XOR U54154 ( .A(n54281), .B(n54282), .Z(n54277) );
  AND U54155 ( .A(n54283), .B(n54284), .Z(n54282) );
  XNOR U54156 ( .A(p_input[819]), .B(n54281), .Z(n54284) );
  XNOR U54157 ( .A(n54281), .B(n53938), .Z(n54283) );
  IV U54158 ( .A(p_input[787]), .Z(n53938) );
  XOR U54159 ( .A(n54285), .B(n54286), .Z(n54281) );
  AND U54160 ( .A(n54287), .B(n54288), .Z(n54286) );
  XNOR U54161 ( .A(p_input[818]), .B(n54285), .Z(n54288) );
  XNOR U54162 ( .A(n54285), .B(n53947), .Z(n54287) );
  IV U54163 ( .A(p_input[786]), .Z(n53947) );
  XOR U54164 ( .A(n54289), .B(n54290), .Z(n54285) );
  AND U54165 ( .A(n54291), .B(n54292), .Z(n54290) );
  XNOR U54166 ( .A(p_input[817]), .B(n54289), .Z(n54292) );
  XNOR U54167 ( .A(n54289), .B(n53956), .Z(n54291) );
  IV U54168 ( .A(p_input[785]), .Z(n53956) );
  XOR U54169 ( .A(n54293), .B(n54294), .Z(n54289) );
  AND U54170 ( .A(n54295), .B(n54296), .Z(n54294) );
  XNOR U54171 ( .A(p_input[816]), .B(n54293), .Z(n54296) );
  XNOR U54172 ( .A(n54293), .B(n53965), .Z(n54295) );
  IV U54173 ( .A(p_input[784]), .Z(n53965) );
  XOR U54174 ( .A(n54297), .B(n54298), .Z(n54293) );
  AND U54175 ( .A(n54299), .B(n54300), .Z(n54298) );
  XNOR U54176 ( .A(p_input[815]), .B(n54297), .Z(n54300) );
  XNOR U54177 ( .A(n54297), .B(n53974), .Z(n54299) );
  IV U54178 ( .A(p_input[783]), .Z(n53974) );
  XOR U54179 ( .A(n54301), .B(n54302), .Z(n54297) );
  AND U54180 ( .A(n54303), .B(n54304), .Z(n54302) );
  XNOR U54181 ( .A(p_input[814]), .B(n54301), .Z(n54304) );
  XNOR U54182 ( .A(n54301), .B(n53983), .Z(n54303) );
  IV U54183 ( .A(p_input[782]), .Z(n53983) );
  XOR U54184 ( .A(n54305), .B(n54306), .Z(n54301) );
  AND U54185 ( .A(n54307), .B(n54308), .Z(n54306) );
  XNOR U54186 ( .A(p_input[813]), .B(n54305), .Z(n54308) );
  XNOR U54187 ( .A(n54305), .B(n53992), .Z(n54307) );
  IV U54188 ( .A(p_input[781]), .Z(n53992) );
  XOR U54189 ( .A(n54309), .B(n54310), .Z(n54305) );
  AND U54190 ( .A(n54311), .B(n54312), .Z(n54310) );
  XNOR U54191 ( .A(p_input[812]), .B(n54309), .Z(n54312) );
  XNOR U54192 ( .A(n54309), .B(n54001), .Z(n54311) );
  IV U54193 ( .A(p_input[780]), .Z(n54001) );
  XOR U54194 ( .A(n54313), .B(n54314), .Z(n54309) );
  AND U54195 ( .A(n54315), .B(n54316), .Z(n54314) );
  XNOR U54196 ( .A(p_input[811]), .B(n54313), .Z(n54316) );
  XNOR U54197 ( .A(n54313), .B(n54010), .Z(n54315) );
  IV U54198 ( .A(p_input[779]), .Z(n54010) );
  XOR U54199 ( .A(n54317), .B(n54318), .Z(n54313) );
  AND U54200 ( .A(n54319), .B(n54320), .Z(n54318) );
  XNOR U54201 ( .A(p_input[810]), .B(n54317), .Z(n54320) );
  XNOR U54202 ( .A(n54317), .B(n54019), .Z(n54319) );
  IV U54203 ( .A(p_input[778]), .Z(n54019) );
  XOR U54204 ( .A(n54321), .B(n54322), .Z(n54317) );
  AND U54205 ( .A(n54323), .B(n54324), .Z(n54322) );
  XNOR U54206 ( .A(p_input[809]), .B(n54321), .Z(n54324) );
  XNOR U54207 ( .A(n54321), .B(n54028), .Z(n54323) );
  IV U54208 ( .A(p_input[777]), .Z(n54028) );
  XOR U54209 ( .A(n54325), .B(n54326), .Z(n54321) );
  AND U54210 ( .A(n54327), .B(n54328), .Z(n54326) );
  XNOR U54211 ( .A(p_input[808]), .B(n54325), .Z(n54328) );
  XNOR U54212 ( .A(n54325), .B(n54037), .Z(n54327) );
  IV U54213 ( .A(p_input[776]), .Z(n54037) );
  XOR U54214 ( .A(n54329), .B(n54330), .Z(n54325) );
  AND U54215 ( .A(n54331), .B(n54332), .Z(n54330) );
  XNOR U54216 ( .A(p_input[807]), .B(n54329), .Z(n54332) );
  XNOR U54217 ( .A(n54329), .B(n54046), .Z(n54331) );
  IV U54218 ( .A(p_input[775]), .Z(n54046) );
  XOR U54219 ( .A(n54333), .B(n54334), .Z(n54329) );
  AND U54220 ( .A(n54335), .B(n54336), .Z(n54334) );
  XNOR U54221 ( .A(p_input[806]), .B(n54333), .Z(n54336) );
  XNOR U54222 ( .A(n54333), .B(n54055), .Z(n54335) );
  IV U54223 ( .A(p_input[774]), .Z(n54055) );
  XOR U54224 ( .A(n54337), .B(n54338), .Z(n54333) );
  AND U54225 ( .A(n54339), .B(n54340), .Z(n54338) );
  XNOR U54226 ( .A(p_input[805]), .B(n54337), .Z(n54340) );
  XNOR U54227 ( .A(n54337), .B(n54064), .Z(n54339) );
  IV U54228 ( .A(p_input[773]), .Z(n54064) );
  XOR U54229 ( .A(n54341), .B(n54342), .Z(n54337) );
  AND U54230 ( .A(n54343), .B(n54344), .Z(n54342) );
  XNOR U54231 ( .A(p_input[804]), .B(n54341), .Z(n54344) );
  XNOR U54232 ( .A(n54341), .B(n54073), .Z(n54343) );
  IV U54233 ( .A(p_input[772]), .Z(n54073) );
  XOR U54234 ( .A(n54345), .B(n54346), .Z(n54341) );
  AND U54235 ( .A(n54347), .B(n54348), .Z(n54346) );
  XNOR U54236 ( .A(p_input[803]), .B(n54345), .Z(n54348) );
  XNOR U54237 ( .A(n54345), .B(n54082), .Z(n54347) );
  IV U54238 ( .A(p_input[771]), .Z(n54082) );
  XOR U54239 ( .A(n54349), .B(n54350), .Z(n54345) );
  AND U54240 ( .A(n54351), .B(n54352), .Z(n54350) );
  XNOR U54241 ( .A(p_input[802]), .B(n54349), .Z(n54352) );
  XNOR U54242 ( .A(n54349), .B(n54091), .Z(n54351) );
  IV U54243 ( .A(p_input[770]), .Z(n54091) );
  XNOR U54244 ( .A(n54353), .B(n54354), .Z(n54349) );
  AND U54245 ( .A(n54355), .B(n54356), .Z(n54354) );
  XOR U54246 ( .A(p_input[801]), .B(n54353), .Z(n54356) );
  XNOR U54247 ( .A(p_input[769]), .B(n54353), .Z(n54355) );
  AND U54248 ( .A(p_input[800]), .B(n54357), .Z(n54353) );
  IV U54249 ( .A(p_input[768]), .Z(n54357) );
  XOR U54250 ( .A(n54358), .B(n54359), .Z(n52536) );
  AND U54251 ( .A(n913), .B(n54360), .Z(n54359) );
  XNOR U54252 ( .A(n54361), .B(n54358), .Z(n54360) );
  XOR U54253 ( .A(n54362), .B(n54363), .Z(n913) );
  AND U54254 ( .A(n54364), .B(n54365), .Z(n54363) );
  XOR U54255 ( .A(n54362), .B(n52551), .Z(n54365) );
  XNOR U54256 ( .A(n54366), .B(n54367), .Z(n52551) );
  AND U54257 ( .A(n54368), .B(n655), .Z(n54367) );
  AND U54258 ( .A(n54366), .B(n54369), .Z(n54368) );
  XNOR U54259 ( .A(n52548), .B(n54362), .Z(n54364) );
  XOR U54260 ( .A(n54370), .B(n54371), .Z(n52548) );
  AND U54261 ( .A(n54372), .B(n652), .Z(n54371) );
  NOR U54262 ( .A(n54370), .B(n54373), .Z(n54372) );
  XOR U54263 ( .A(n54374), .B(n54375), .Z(n54362) );
  AND U54264 ( .A(n54376), .B(n54377), .Z(n54375) );
  XOR U54265 ( .A(n54374), .B(n52563), .Z(n54377) );
  XOR U54266 ( .A(n54378), .B(n54379), .Z(n52563) );
  AND U54267 ( .A(n655), .B(n54380), .Z(n54379) );
  XOR U54268 ( .A(n54381), .B(n54378), .Z(n54380) );
  XNOR U54269 ( .A(n52560), .B(n54374), .Z(n54376) );
  XOR U54270 ( .A(n54382), .B(n54383), .Z(n52560) );
  AND U54271 ( .A(n652), .B(n54384), .Z(n54383) );
  XOR U54272 ( .A(n54385), .B(n54382), .Z(n54384) );
  XOR U54273 ( .A(n54386), .B(n54387), .Z(n54374) );
  AND U54274 ( .A(n54388), .B(n54389), .Z(n54387) );
  XOR U54275 ( .A(n54386), .B(n52575), .Z(n54389) );
  XOR U54276 ( .A(n54390), .B(n54391), .Z(n52575) );
  AND U54277 ( .A(n655), .B(n54392), .Z(n54391) );
  XOR U54278 ( .A(n54393), .B(n54390), .Z(n54392) );
  XNOR U54279 ( .A(n52572), .B(n54386), .Z(n54388) );
  XOR U54280 ( .A(n54394), .B(n54395), .Z(n52572) );
  AND U54281 ( .A(n652), .B(n54396), .Z(n54395) );
  XOR U54282 ( .A(n54397), .B(n54394), .Z(n54396) );
  XOR U54283 ( .A(n54398), .B(n54399), .Z(n54386) );
  AND U54284 ( .A(n54400), .B(n54401), .Z(n54399) );
  XOR U54285 ( .A(n54398), .B(n52587), .Z(n54401) );
  XOR U54286 ( .A(n54402), .B(n54403), .Z(n52587) );
  AND U54287 ( .A(n655), .B(n54404), .Z(n54403) );
  XOR U54288 ( .A(n54405), .B(n54402), .Z(n54404) );
  XNOR U54289 ( .A(n52584), .B(n54398), .Z(n54400) );
  XOR U54290 ( .A(n54406), .B(n54407), .Z(n52584) );
  AND U54291 ( .A(n652), .B(n54408), .Z(n54407) );
  XOR U54292 ( .A(n54409), .B(n54406), .Z(n54408) );
  XOR U54293 ( .A(n54410), .B(n54411), .Z(n54398) );
  AND U54294 ( .A(n54412), .B(n54413), .Z(n54411) );
  XOR U54295 ( .A(n54410), .B(n52599), .Z(n54413) );
  XOR U54296 ( .A(n54414), .B(n54415), .Z(n52599) );
  AND U54297 ( .A(n655), .B(n54416), .Z(n54415) );
  XOR U54298 ( .A(n54417), .B(n54414), .Z(n54416) );
  XNOR U54299 ( .A(n52596), .B(n54410), .Z(n54412) );
  XOR U54300 ( .A(n54418), .B(n54419), .Z(n52596) );
  AND U54301 ( .A(n652), .B(n54420), .Z(n54419) );
  XOR U54302 ( .A(n54421), .B(n54418), .Z(n54420) );
  XOR U54303 ( .A(n54422), .B(n54423), .Z(n54410) );
  AND U54304 ( .A(n54424), .B(n54425), .Z(n54423) );
  XOR U54305 ( .A(n54422), .B(n52611), .Z(n54425) );
  XOR U54306 ( .A(n54426), .B(n54427), .Z(n52611) );
  AND U54307 ( .A(n655), .B(n54428), .Z(n54427) );
  XOR U54308 ( .A(n54429), .B(n54426), .Z(n54428) );
  XNOR U54309 ( .A(n52608), .B(n54422), .Z(n54424) );
  XOR U54310 ( .A(n54430), .B(n54431), .Z(n52608) );
  AND U54311 ( .A(n652), .B(n54432), .Z(n54431) );
  XOR U54312 ( .A(n54433), .B(n54430), .Z(n54432) );
  XOR U54313 ( .A(n54434), .B(n54435), .Z(n54422) );
  AND U54314 ( .A(n54436), .B(n54437), .Z(n54435) );
  XOR U54315 ( .A(n54434), .B(n52623), .Z(n54437) );
  XOR U54316 ( .A(n54438), .B(n54439), .Z(n52623) );
  AND U54317 ( .A(n655), .B(n54440), .Z(n54439) );
  XOR U54318 ( .A(n54441), .B(n54438), .Z(n54440) );
  XNOR U54319 ( .A(n52620), .B(n54434), .Z(n54436) );
  XOR U54320 ( .A(n54442), .B(n54443), .Z(n52620) );
  AND U54321 ( .A(n652), .B(n54444), .Z(n54443) );
  XOR U54322 ( .A(n54445), .B(n54442), .Z(n54444) );
  XOR U54323 ( .A(n54446), .B(n54447), .Z(n54434) );
  AND U54324 ( .A(n54448), .B(n54449), .Z(n54447) );
  XOR U54325 ( .A(n54446), .B(n52635), .Z(n54449) );
  XOR U54326 ( .A(n54450), .B(n54451), .Z(n52635) );
  AND U54327 ( .A(n655), .B(n54452), .Z(n54451) );
  XOR U54328 ( .A(n54453), .B(n54450), .Z(n54452) );
  XNOR U54329 ( .A(n52632), .B(n54446), .Z(n54448) );
  XOR U54330 ( .A(n54454), .B(n54455), .Z(n52632) );
  AND U54331 ( .A(n652), .B(n54456), .Z(n54455) );
  XOR U54332 ( .A(n54457), .B(n54454), .Z(n54456) );
  XOR U54333 ( .A(n54458), .B(n54459), .Z(n54446) );
  AND U54334 ( .A(n54460), .B(n54461), .Z(n54459) );
  XOR U54335 ( .A(n54458), .B(n52647), .Z(n54461) );
  XOR U54336 ( .A(n54462), .B(n54463), .Z(n52647) );
  AND U54337 ( .A(n655), .B(n54464), .Z(n54463) );
  XOR U54338 ( .A(n54465), .B(n54462), .Z(n54464) );
  XNOR U54339 ( .A(n52644), .B(n54458), .Z(n54460) );
  XOR U54340 ( .A(n54466), .B(n54467), .Z(n52644) );
  AND U54341 ( .A(n652), .B(n54468), .Z(n54467) );
  XOR U54342 ( .A(n54469), .B(n54466), .Z(n54468) );
  XOR U54343 ( .A(n54470), .B(n54471), .Z(n54458) );
  AND U54344 ( .A(n54472), .B(n54473), .Z(n54471) );
  XOR U54345 ( .A(n54470), .B(n52659), .Z(n54473) );
  XOR U54346 ( .A(n54474), .B(n54475), .Z(n52659) );
  AND U54347 ( .A(n655), .B(n54476), .Z(n54475) );
  XOR U54348 ( .A(n54477), .B(n54474), .Z(n54476) );
  XNOR U54349 ( .A(n52656), .B(n54470), .Z(n54472) );
  XOR U54350 ( .A(n54478), .B(n54479), .Z(n52656) );
  AND U54351 ( .A(n652), .B(n54480), .Z(n54479) );
  XOR U54352 ( .A(n54481), .B(n54478), .Z(n54480) );
  XOR U54353 ( .A(n54482), .B(n54483), .Z(n54470) );
  AND U54354 ( .A(n54484), .B(n54485), .Z(n54483) );
  XOR U54355 ( .A(n54482), .B(n52671), .Z(n54485) );
  XOR U54356 ( .A(n54486), .B(n54487), .Z(n52671) );
  AND U54357 ( .A(n655), .B(n54488), .Z(n54487) );
  XOR U54358 ( .A(n54489), .B(n54486), .Z(n54488) );
  XNOR U54359 ( .A(n52668), .B(n54482), .Z(n54484) );
  XOR U54360 ( .A(n54490), .B(n54491), .Z(n52668) );
  AND U54361 ( .A(n652), .B(n54492), .Z(n54491) );
  XOR U54362 ( .A(n54493), .B(n54490), .Z(n54492) );
  XOR U54363 ( .A(n54494), .B(n54495), .Z(n54482) );
  AND U54364 ( .A(n54496), .B(n54497), .Z(n54495) );
  XOR U54365 ( .A(n54494), .B(n52683), .Z(n54497) );
  XOR U54366 ( .A(n54498), .B(n54499), .Z(n52683) );
  AND U54367 ( .A(n655), .B(n54500), .Z(n54499) );
  XOR U54368 ( .A(n54501), .B(n54498), .Z(n54500) );
  XNOR U54369 ( .A(n52680), .B(n54494), .Z(n54496) );
  XOR U54370 ( .A(n54502), .B(n54503), .Z(n52680) );
  AND U54371 ( .A(n652), .B(n54504), .Z(n54503) );
  XOR U54372 ( .A(n54505), .B(n54502), .Z(n54504) );
  XOR U54373 ( .A(n54506), .B(n54507), .Z(n54494) );
  AND U54374 ( .A(n54508), .B(n54509), .Z(n54507) );
  XOR U54375 ( .A(n54506), .B(n52695), .Z(n54509) );
  XOR U54376 ( .A(n54510), .B(n54511), .Z(n52695) );
  AND U54377 ( .A(n655), .B(n54512), .Z(n54511) );
  XOR U54378 ( .A(n54513), .B(n54510), .Z(n54512) );
  XNOR U54379 ( .A(n52692), .B(n54506), .Z(n54508) );
  XOR U54380 ( .A(n54514), .B(n54515), .Z(n52692) );
  AND U54381 ( .A(n652), .B(n54516), .Z(n54515) );
  XOR U54382 ( .A(n54517), .B(n54514), .Z(n54516) );
  XOR U54383 ( .A(n54518), .B(n54519), .Z(n54506) );
  AND U54384 ( .A(n54520), .B(n54521), .Z(n54519) );
  XOR U54385 ( .A(n54518), .B(n52707), .Z(n54521) );
  XOR U54386 ( .A(n54522), .B(n54523), .Z(n52707) );
  AND U54387 ( .A(n655), .B(n54524), .Z(n54523) );
  XOR U54388 ( .A(n54525), .B(n54522), .Z(n54524) );
  XNOR U54389 ( .A(n52704), .B(n54518), .Z(n54520) );
  XOR U54390 ( .A(n54526), .B(n54527), .Z(n52704) );
  AND U54391 ( .A(n652), .B(n54528), .Z(n54527) );
  XOR U54392 ( .A(n54529), .B(n54526), .Z(n54528) );
  XOR U54393 ( .A(n54530), .B(n54531), .Z(n54518) );
  AND U54394 ( .A(n54532), .B(n54533), .Z(n54531) );
  XOR U54395 ( .A(n54530), .B(n52719), .Z(n54533) );
  XOR U54396 ( .A(n54534), .B(n54535), .Z(n52719) );
  AND U54397 ( .A(n655), .B(n54536), .Z(n54535) );
  XOR U54398 ( .A(n54537), .B(n54534), .Z(n54536) );
  XNOR U54399 ( .A(n52716), .B(n54530), .Z(n54532) );
  XOR U54400 ( .A(n54538), .B(n54539), .Z(n52716) );
  AND U54401 ( .A(n652), .B(n54540), .Z(n54539) );
  XOR U54402 ( .A(n54541), .B(n54538), .Z(n54540) );
  XOR U54403 ( .A(n54542), .B(n54543), .Z(n54530) );
  AND U54404 ( .A(n54544), .B(n54545), .Z(n54543) );
  XOR U54405 ( .A(n54542), .B(n52731), .Z(n54545) );
  XOR U54406 ( .A(n54546), .B(n54547), .Z(n52731) );
  AND U54407 ( .A(n655), .B(n54548), .Z(n54547) );
  XOR U54408 ( .A(n54549), .B(n54546), .Z(n54548) );
  XNOR U54409 ( .A(n52728), .B(n54542), .Z(n54544) );
  XOR U54410 ( .A(n54550), .B(n54551), .Z(n52728) );
  AND U54411 ( .A(n652), .B(n54552), .Z(n54551) );
  XOR U54412 ( .A(n54553), .B(n54550), .Z(n54552) );
  XOR U54413 ( .A(n54554), .B(n54555), .Z(n54542) );
  AND U54414 ( .A(n54556), .B(n54557), .Z(n54555) );
  XOR U54415 ( .A(n54554), .B(n52743), .Z(n54557) );
  XOR U54416 ( .A(n54558), .B(n54559), .Z(n52743) );
  AND U54417 ( .A(n655), .B(n54560), .Z(n54559) );
  XOR U54418 ( .A(n54561), .B(n54558), .Z(n54560) );
  XNOR U54419 ( .A(n52740), .B(n54554), .Z(n54556) );
  XOR U54420 ( .A(n54562), .B(n54563), .Z(n52740) );
  AND U54421 ( .A(n652), .B(n54564), .Z(n54563) );
  XOR U54422 ( .A(n54565), .B(n54562), .Z(n54564) );
  XOR U54423 ( .A(n54566), .B(n54567), .Z(n54554) );
  AND U54424 ( .A(n54568), .B(n54569), .Z(n54567) );
  XOR U54425 ( .A(n54566), .B(n52755), .Z(n54569) );
  XOR U54426 ( .A(n54570), .B(n54571), .Z(n52755) );
  AND U54427 ( .A(n655), .B(n54572), .Z(n54571) );
  XOR U54428 ( .A(n54573), .B(n54570), .Z(n54572) );
  XNOR U54429 ( .A(n52752), .B(n54566), .Z(n54568) );
  XOR U54430 ( .A(n54574), .B(n54575), .Z(n52752) );
  AND U54431 ( .A(n652), .B(n54576), .Z(n54575) );
  XOR U54432 ( .A(n54577), .B(n54574), .Z(n54576) );
  XOR U54433 ( .A(n54578), .B(n54579), .Z(n54566) );
  AND U54434 ( .A(n54580), .B(n54581), .Z(n54579) );
  XOR U54435 ( .A(n54578), .B(n52767), .Z(n54581) );
  XOR U54436 ( .A(n54582), .B(n54583), .Z(n52767) );
  AND U54437 ( .A(n655), .B(n54584), .Z(n54583) );
  XOR U54438 ( .A(n54585), .B(n54582), .Z(n54584) );
  XNOR U54439 ( .A(n52764), .B(n54578), .Z(n54580) );
  XOR U54440 ( .A(n54586), .B(n54587), .Z(n52764) );
  AND U54441 ( .A(n652), .B(n54588), .Z(n54587) );
  XOR U54442 ( .A(n54589), .B(n54586), .Z(n54588) );
  XOR U54443 ( .A(n54590), .B(n54591), .Z(n54578) );
  AND U54444 ( .A(n54592), .B(n54593), .Z(n54591) );
  XOR U54445 ( .A(n54590), .B(n52779), .Z(n54593) );
  XOR U54446 ( .A(n54594), .B(n54595), .Z(n52779) );
  AND U54447 ( .A(n655), .B(n54596), .Z(n54595) );
  XOR U54448 ( .A(n54597), .B(n54594), .Z(n54596) );
  XNOR U54449 ( .A(n52776), .B(n54590), .Z(n54592) );
  XOR U54450 ( .A(n54598), .B(n54599), .Z(n52776) );
  AND U54451 ( .A(n652), .B(n54600), .Z(n54599) );
  XOR U54452 ( .A(n54601), .B(n54598), .Z(n54600) );
  XOR U54453 ( .A(n54602), .B(n54603), .Z(n54590) );
  AND U54454 ( .A(n54604), .B(n54605), .Z(n54603) );
  XOR U54455 ( .A(n54602), .B(n52791), .Z(n54605) );
  XOR U54456 ( .A(n54606), .B(n54607), .Z(n52791) );
  AND U54457 ( .A(n655), .B(n54608), .Z(n54607) );
  XOR U54458 ( .A(n54609), .B(n54606), .Z(n54608) );
  XNOR U54459 ( .A(n52788), .B(n54602), .Z(n54604) );
  XOR U54460 ( .A(n54610), .B(n54611), .Z(n52788) );
  AND U54461 ( .A(n652), .B(n54612), .Z(n54611) );
  XOR U54462 ( .A(n54613), .B(n54610), .Z(n54612) );
  XOR U54463 ( .A(n54614), .B(n54615), .Z(n54602) );
  AND U54464 ( .A(n54616), .B(n54617), .Z(n54615) );
  XOR U54465 ( .A(n54614), .B(n52803), .Z(n54617) );
  XOR U54466 ( .A(n54618), .B(n54619), .Z(n52803) );
  AND U54467 ( .A(n655), .B(n54620), .Z(n54619) );
  XOR U54468 ( .A(n54621), .B(n54618), .Z(n54620) );
  XNOR U54469 ( .A(n52800), .B(n54614), .Z(n54616) );
  XOR U54470 ( .A(n54622), .B(n54623), .Z(n52800) );
  AND U54471 ( .A(n652), .B(n54624), .Z(n54623) );
  XOR U54472 ( .A(n54625), .B(n54622), .Z(n54624) );
  XOR U54473 ( .A(n54626), .B(n54627), .Z(n54614) );
  AND U54474 ( .A(n54628), .B(n54629), .Z(n54627) );
  XOR U54475 ( .A(n54626), .B(n52815), .Z(n54629) );
  XOR U54476 ( .A(n54630), .B(n54631), .Z(n52815) );
  AND U54477 ( .A(n655), .B(n54632), .Z(n54631) );
  XOR U54478 ( .A(n54633), .B(n54630), .Z(n54632) );
  XNOR U54479 ( .A(n52812), .B(n54626), .Z(n54628) );
  XOR U54480 ( .A(n54634), .B(n54635), .Z(n52812) );
  AND U54481 ( .A(n652), .B(n54636), .Z(n54635) );
  XOR U54482 ( .A(n54637), .B(n54634), .Z(n54636) );
  XOR U54483 ( .A(n54638), .B(n54639), .Z(n54626) );
  AND U54484 ( .A(n54640), .B(n54641), .Z(n54639) );
  XOR U54485 ( .A(n54638), .B(n52827), .Z(n54641) );
  XOR U54486 ( .A(n54642), .B(n54643), .Z(n52827) );
  AND U54487 ( .A(n655), .B(n54644), .Z(n54643) );
  XOR U54488 ( .A(n54645), .B(n54642), .Z(n54644) );
  XNOR U54489 ( .A(n52824), .B(n54638), .Z(n54640) );
  XOR U54490 ( .A(n54646), .B(n54647), .Z(n52824) );
  AND U54491 ( .A(n652), .B(n54648), .Z(n54647) );
  XOR U54492 ( .A(n54649), .B(n54646), .Z(n54648) );
  XOR U54493 ( .A(n54650), .B(n54651), .Z(n54638) );
  AND U54494 ( .A(n54652), .B(n54653), .Z(n54651) );
  XOR U54495 ( .A(n54650), .B(n52839), .Z(n54653) );
  XOR U54496 ( .A(n54654), .B(n54655), .Z(n52839) );
  AND U54497 ( .A(n655), .B(n54656), .Z(n54655) );
  XOR U54498 ( .A(n54657), .B(n54654), .Z(n54656) );
  XNOR U54499 ( .A(n52836), .B(n54650), .Z(n54652) );
  XOR U54500 ( .A(n54658), .B(n54659), .Z(n52836) );
  AND U54501 ( .A(n652), .B(n54660), .Z(n54659) );
  XOR U54502 ( .A(n54661), .B(n54658), .Z(n54660) );
  XOR U54503 ( .A(n54662), .B(n54663), .Z(n54650) );
  AND U54504 ( .A(n54664), .B(n54665), .Z(n54663) );
  XOR U54505 ( .A(n54662), .B(n52851), .Z(n54665) );
  XOR U54506 ( .A(n54666), .B(n54667), .Z(n52851) );
  AND U54507 ( .A(n655), .B(n54668), .Z(n54667) );
  XOR U54508 ( .A(n54669), .B(n54666), .Z(n54668) );
  XNOR U54509 ( .A(n52848), .B(n54662), .Z(n54664) );
  XOR U54510 ( .A(n54670), .B(n54671), .Z(n52848) );
  AND U54511 ( .A(n652), .B(n54672), .Z(n54671) );
  XOR U54512 ( .A(n54673), .B(n54670), .Z(n54672) );
  XOR U54513 ( .A(n54674), .B(n54675), .Z(n54662) );
  AND U54514 ( .A(n54676), .B(n54677), .Z(n54675) );
  XOR U54515 ( .A(n54674), .B(n52863), .Z(n54677) );
  XOR U54516 ( .A(n54678), .B(n54679), .Z(n52863) );
  AND U54517 ( .A(n655), .B(n54680), .Z(n54679) );
  XOR U54518 ( .A(n54681), .B(n54678), .Z(n54680) );
  XNOR U54519 ( .A(n52860), .B(n54674), .Z(n54676) );
  XOR U54520 ( .A(n54682), .B(n54683), .Z(n52860) );
  AND U54521 ( .A(n652), .B(n54684), .Z(n54683) );
  XOR U54522 ( .A(n54685), .B(n54682), .Z(n54684) );
  XOR U54523 ( .A(n54686), .B(n54687), .Z(n54674) );
  AND U54524 ( .A(n54688), .B(n54689), .Z(n54687) );
  XOR U54525 ( .A(n54686), .B(n52875), .Z(n54689) );
  XOR U54526 ( .A(n54690), .B(n54691), .Z(n52875) );
  AND U54527 ( .A(n655), .B(n54692), .Z(n54691) );
  XOR U54528 ( .A(n54693), .B(n54690), .Z(n54692) );
  XNOR U54529 ( .A(n52872), .B(n54686), .Z(n54688) );
  XOR U54530 ( .A(n54694), .B(n54695), .Z(n52872) );
  AND U54531 ( .A(n652), .B(n54696), .Z(n54695) );
  XOR U54532 ( .A(n54697), .B(n54694), .Z(n54696) );
  XOR U54533 ( .A(n54698), .B(n54699), .Z(n54686) );
  AND U54534 ( .A(n54700), .B(n54701), .Z(n54699) );
  XOR U54535 ( .A(n54698), .B(n52887), .Z(n54701) );
  XOR U54536 ( .A(n54702), .B(n54703), .Z(n52887) );
  AND U54537 ( .A(n655), .B(n54704), .Z(n54703) );
  XOR U54538 ( .A(n54705), .B(n54702), .Z(n54704) );
  XNOR U54539 ( .A(n52884), .B(n54698), .Z(n54700) );
  XOR U54540 ( .A(n54706), .B(n54707), .Z(n52884) );
  AND U54541 ( .A(n652), .B(n54708), .Z(n54707) );
  XOR U54542 ( .A(n54709), .B(n54706), .Z(n54708) );
  XOR U54543 ( .A(n54710), .B(n54711), .Z(n54698) );
  AND U54544 ( .A(n54712), .B(n54713), .Z(n54711) );
  XOR U54545 ( .A(n54710), .B(n52899), .Z(n54713) );
  XOR U54546 ( .A(n54714), .B(n54715), .Z(n52899) );
  AND U54547 ( .A(n655), .B(n54716), .Z(n54715) );
  XOR U54548 ( .A(n54717), .B(n54714), .Z(n54716) );
  XNOR U54549 ( .A(n52896), .B(n54710), .Z(n54712) );
  XOR U54550 ( .A(n54718), .B(n54719), .Z(n52896) );
  AND U54551 ( .A(n652), .B(n54720), .Z(n54719) );
  XOR U54552 ( .A(n54721), .B(n54718), .Z(n54720) );
  XOR U54553 ( .A(n54722), .B(n54723), .Z(n54710) );
  AND U54554 ( .A(n54724), .B(n54725), .Z(n54723) );
  XNOR U54555 ( .A(n54726), .B(n52912), .Z(n54725) );
  XOR U54556 ( .A(n54727), .B(n54728), .Z(n52912) );
  AND U54557 ( .A(n655), .B(n54729), .Z(n54728) );
  XOR U54558 ( .A(n54727), .B(n54730), .Z(n54729) );
  XNOR U54559 ( .A(n52909), .B(n54722), .Z(n54724) );
  XOR U54560 ( .A(n54731), .B(n54732), .Z(n52909) );
  AND U54561 ( .A(n652), .B(n54733), .Z(n54732) );
  XOR U54562 ( .A(n54731), .B(n54734), .Z(n54733) );
  IV U54563 ( .A(n54726), .Z(n54722) );
  AND U54564 ( .A(n54358), .B(n54361), .Z(n54726) );
  XNOR U54565 ( .A(n54735), .B(n54736), .Z(n54361) );
  AND U54566 ( .A(n655), .B(n54737), .Z(n54736) );
  XNOR U54567 ( .A(n54738), .B(n54735), .Z(n54737) );
  XOR U54568 ( .A(n54739), .B(n54740), .Z(n655) );
  AND U54569 ( .A(n54741), .B(n54742), .Z(n54740) );
  XOR U54570 ( .A(n54369), .B(n54739), .Z(n54742) );
  IV U54571 ( .A(n54743), .Z(n54369) );
  AND U54572 ( .A(p_input[767]), .B(p_input[735]), .Z(n54743) );
  XOR U54573 ( .A(n54739), .B(n54366), .Z(n54741) );
  AND U54574 ( .A(p_input[671]), .B(p_input[703]), .Z(n54366) );
  XOR U54575 ( .A(n54744), .B(n54745), .Z(n54739) );
  AND U54576 ( .A(n54746), .B(n54747), .Z(n54745) );
  XOR U54577 ( .A(n54744), .B(n54381), .Z(n54747) );
  XNOR U54578 ( .A(p_input[734]), .B(n54748), .Z(n54381) );
  AND U54579 ( .A(n1071), .B(n54749), .Z(n54748) );
  XOR U54580 ( .A(p_input[766]), .B(p_input[734]), .Z(n54749) );
  XNOR U54581 ( .A(n54378), .B(n54744), .Z(n54746) );
  XOR U54582 ( .A(n54750), .B(n54751), .Z(n54378) );
  AND U54583 ( .A(n1069), .B(n54752), .Z(n54751) );
  XOR U54584 ( .A(p_input[702]), .B(p_input[670]), .Z(n54752) );
  XOR U54585 ( .A(n54753), .B(n54754), .Z(n54744) );
  AND U54586 ( .A(n54755), .B(n54756), .Z(n54754) );
  XOR U54587 ( .A(n54753), .B(n54393), .Z(n54756) );
  XNOR U54588 ( .A(p_input[733]), .B(n54757), .Z(n54393) );
  AND U54589 ( .A(n1071), .B(n54758), .Z(n54757) );
  XOR U54590 ( .A(p_input[765]), .B(p_input[733]), .Z(n54758) );
  XNOR U54591 ( .A(n54390), .B(n54753), .Z(n54755) );
  XOR U54592 ( .A(n54759), .B(n54760), .Z(n54390) );
  AND U54593 ( .A(n1069), .B(n54761), .Z(n54760) );
  XOR U54594 ( .A(p_input[701]), .B(p_input[669]), .Z(n54761) );
  XOR U54595 ( .A(n54762), .B(n54763), .Z(n54753) );
  AND U54596 ( .A(n54764), .B(n54765), .Z(n54763) );
  XOR U54597 ( .A(n54762), .B(n54405), .Z(n54765) );
  XNOR U54598 ( .A(p_input[732]), .B(n54766), .Z(n54405) );
  AND U54599 ( .A(n1071), .B(n54767), .Z(n54766) );
  XOR U54600 ( .A(p_input[764]), .B(p_input[732]), .Z(n54767) );
  XNOR U54601 ( .A(n54402), .B(n54762), .Z(n54764) );
  XOR U54602 ( .A(n54768), .B(n54769), .Z(n54402) );
  AND U54603 ( .A(n1069), .B(n54770), .Z(n54769) );
  XOR U54604 ( .A(p_input[700]), .B(p_input[668]), .Z(n54770) );
  XOR U54605 ( .A(n54771), .B(n54772), .Z(n54762) );
  AND U54606 ( .A(n54773), .B(n54774), .Z(n54772) );
  XOR U54607 ( .A(n54771), .B(n54417), .Z(n54774) );
  XNOR U54608 ( .A(p_input[731]), .B(n54775), .Z(n54417) );
  AND U54609 ( .A(n1071), .B(n54776), .Z(n54775) );
  XOR U54610 ( .A(p_input[763]), .B(p_input[731]), .Z(n54776) );
  XNOR U54611 ( .A(n54414), .B(n54771), .Z(n54773) );
  XOR U54612 ( .A(n54777), .B(n54778), .Z(n54414) );
  AND U54613 ( .A(n1069), .B(n54779), .Z(n54778) );
  XOR U54614 ( .A(p_input[699]), .B(p_input[667]), .Z(n54779) );
  XOR U54615 ( .A(n54780), .B(n54781), .Z(n54771) );
  AND U54616 ( .A(n54782), .B(n54783), .Z(n54781) );
  XOR U54617 ( .A(n54780), .B(n54429), .Z(n54783) );
  XNOR U54618 ( .A(p_input[730]), .B(n54784), .Z(n54429) );
  AND U54619 ( .A(n1071), .B(n54785), .Z(n54784) );
  XOR U54620 ( .A(p_input[762]), .B(p_input[730]), .Z(n54785) );
  XNOR U54621 ( .A(n54426), .B(n54780), .Z(n54782) );
  XOR U54622 ( .A(n54786), .B(n54787), .Z(n54426) );
  AND U54623 ( .A(n1069), .B(n54788), .Z(n54787) );
  XOR U54624 ( .A(p_input[698]), .B(p_input[666]), .Z(n54788) );
  XOR U54625 ( .A(n54789), .B(n54790), .Z(n54780) );
  AND U54626 ( .A(n54791), .B(n54792), .Z(n54790) );
  XOR U54627 ( .A(n54789), .B(n54441), .Z(n54792) );
  XNOR U54628 ( .A(p_input[729]), .B(n54793), .Z(n54441) );
  AND U54629 ( .A(n1071), .B(n54794), .Z(n54793) );
  XOR U54630 ( .A(p_input[761]), .B(p_input[729]), .Z(n54794) );
  XNOR U54631 ( .A(n54438), .B(n54789), .Z(n54791) );
  XOR U54632 ( .A(n54795), .B(n54796), .Z(n54438) );
  AND U54633 ( .A(n1069), .B(n54797), .Z(n54796) );
  XOR U54634 ( .A(p_input[697]), .B(p_input[665]), .Z(n54797) );
  XOR U54635 ( .A(n54798), .B(n54799), .Z(n54789) );
  AND U54636 ( .A(n54800), .B(n54801), .Z(n54799) );
  XOR U54637 ( .A(n54798), .B(n54453), .Z(n54801) );
  XNOR U54638 ( .A(p_input[728]), .B(n54802), .Z(n54453) );
  AND U54639 ( .A(n1071), .B(n54803), .Z(n54802) );
  XOR U54640 ( .A(p_input[760]), .B(p_input[728]), .Z(n54803) );
  XNOR U54641 ( .A(n54450), .B(n54798), .Z(n54800) );
  XOR U54642 ( .A(n54804), .B(n54805), .Z(n54450) );
  AND U54643 ( .A(n1069), .B(n54806), .Z(n54805) );
  XOR U54644 ( .A(p_input[696]), .B(p_input[664]), .Z(n54806) );
  XOR U54645 ( .A(n54807), .B(n54808), .Z(n54798) );
  AND U54646 ( .A(n54809), .B(n54810), .Z(n54808) );
  XOR U54647 ( .A(n54807), .B(n54465), .Z(n54810) );
  XNOR U54648 ( .A(p_input[727]), .B(n54811), .Z(n54465) );
  AND U54649 ( .A(n1071), .B(n54812), .Z(n54811) );
  XOR U54650 ( .A(p_input[759]), .B(p_input[727]), .Z(n54812) );
  XNOR U54651 ( .A(n54462), .B(n54807), .Z(n54809) );
  XOR U54652 ( .A(n54813), .B(n54814), .Z(n54462) );
  AND U54653 ( .A(n1069), .B(n54815), .Z(n54814) );
  XOR U54654 ( .A(p_input[695]), .B(p_input[663]), .Z(n54815) );
  XOR U54655 ( .A(n54816), .B(n54817), .Z(n54807) );
  AND U54656 ( .A(n54818), .B(n54819), .Z(n54817) );
  XOR U54657 ( .A(n54816), .B(n54477), .Z(n54819) );
  XNOR U54658 ( .A(p_input[726]), .B(n54820), .Z(n54477) );
  AND U54659 ( .A(n1071), .B(n54821), .Z(n54820) );
  XOR U54660 ( .A(p_input[758]), .B(p_input[726]), .Z(n54821) );
  XNOR U54661 ( .A(n54474), .B(n54816), .Z(n54818) );
  XOR U54662 ( .A(n54822), .B(n54823), .Z(n54474) );
  AND U54663 ( .A(n1069), .B(n54824), .Z(n54823) );
  XOR U54664 ( .A(p_input[694]), .B(p_input[662]), .Z(n54824) );
  XOR U54665 ( .A(n54825), .B(n54826), .Z(n54816) );
  AND U54666 ( .A(n54827), .B(n54828), .Z(n54826) );
  XOR U54667 ( .A(n54825), .B(n54489), .Z(n54828) );
  XNOR U54668 ( .A(p_input[725]), .B(n54829), .Z(n54489) );
  AND U54669 ( .A(n1071), .B(n54830), .Z(n54829) );
  XOR U54670 ( .A(p_input[757]), .B(p_input[725]), .Z(n54830) );
  XNOR U54671 ( .A(n54486), .B(n54825), .Z(n54827) );
  XOR U54672 ( .A(n54831), .B(n54832), .Z(n54486) );
  AND U54673 ( .A(n1069), .B(n54833), .Z(n54832) );
  XOR U54674 ( .A(p_input[693]), .B(p_input[661]), .Z(n54833) );
  XOR U54675 ( .A(n54834), .B(n54835), .Z(n54825) );
  AND U54676 ( .A(n54836), .B(n54837), .Z(n54835) );
  XOR U54677 ( .A(n54834), .B(n54501), .Z(n54837) );
  XNOR U54678 ( .A(p_input[724]), .B(n54838), .Z(n54501) );
  AND U54679 ( .A(n1071), .B(n54839), .Z(n54838) );
  XOR U54680 ( .A(p_input[756]), .B(p_input[724]), .Z(n54839) );
  XNOR U54681 ( .A(n54498), .B(n54834), .Z(n54836) );
  XOR U54682 ( .A(n54840), .B(n54841), .Z(n54498) );
  AND U54683 ( .A(n1069), .B(n54842), .Z(n54841) );
  XOR U54684 ( .A(p_input[692]), .B(p_input[660]), .Z(n54842) );
  XOR U54685 ( .A(n54843), .B(n54844), .Z(n54834) );
  AND U54686 ( .A(n54845), .B(n54846), .Z(n54844) );
  XOR U54687 ( .A(n54843), .B(n54513), .Z(n54846) );
  XNOR U54688 ( .A(p_input[723]), .B(n54847), .Z(n54513) );
  AND U54689 ( .A(n1071), .B(n54848), .Z(n54847) );
  XOR U54690 ( .A(p_input[755]), .B(p_input[723]), .Z(n54848) );
  XNOR U54691 ( .A(n54510), .B(n54843), .Z(n54845) );
  XOR U54692 ( .A(n54849), .B(n54850), .Z(n54510) );
  AND U54693 ( .A(n1069), .B(n54851), .Z(n54850) );
  XOR U54694 ( .A(p_input[691]), .B(p_input[659]), .Z(n54851) );
  XOR U54695 ( .A(n54852), .B(n54853), .Z(n54843) );
  AND U54696 ( .A(n54854), .B(n54855), .Z(n54853) );
  XOR U54697 ( .A(n54852), .B(n54525), .Z(n54855) );
  XNOR U54698 ( .A(p_input[722]), .B(n54856), .Z(n54525) );
  AND U54699 ( .A(n1071), .B(n54857), .Z(n54856) );
  XOR U54700 ( .A(p_input[754]), .B(p_input[722]), .Z(n54857) );
  XNOR U54701 ( .A(n54522), .B(n54852), .Z(n54854) );
  XOR U54702 ( .A(n54858), .B(n54859), .Z(n54522) );
  AND U54703 ( .A(n1069), .B(n54860), .Z(n54859) );
  XOR U54704 ( .A(p_input[690]), .B(p_input[658]), .Z(n54860) );
  XOR U54705 ( .A(n54861), .B(n54862), .Z(n54852) );
  AND U54706 ( .A(n54863), .B(n54864), .Z(n54862) );
  XOR U54707 ( .A(n54861), .B(n54537), .Z(n54864) );
  XNOR U54708 ( .A(p_input[721]), .B(n54865), .Z(n54537) );
  AND U54709 ( .A(n1071), .B(n54866), .Z(n54865) );
  XOR U54710 ( .A(p_input[753]), .B(p_input[721]), .Z(n54866) );
  XNOR U54711 ( .A(n54534), .B(n54861), .Z(n54863) );
  XOR U54712 ( .A(n54867), .B(n54868), .Z(n54534) );
  AND U54713 ( .A(n1069), .B(n54869), .Z(n54868) );
  XOR U54714 ( .A(p_input[689]), .B(p_input[657]), .Z(n54869) );
  XOR U54715 ( .A(n54870), .B(n54871), .Z(n54861) );
  AND U54716 ( .A(n54872), .B(n54873), .Z(n54871) );
  XOR U54717 ( .A(n54870), .B(n54549), .Z(n54873) );
  XNOR U54718 ( .A(p_input[720]), .B(n54874), .Z(n54549) );
  AND U54719 ( .A(n1071), .B(n54875), .Z(n54874) );
  XOR U54720 ( .A(p_input[752]), .B(p_input[720]), .Z(n54875) );
  XNOR U54721 ( .A(n54546), .B(n54870), .Z(n54872) );
  XOR U54722 ( .A(n54876), .B(n54877), .Z(n54546) );
  AND U54723 ( .A(n1069), .B(n54878), .Z(n54877) );
  XOR U54724 ( .A(p_input[688]), .B(p_input[656]), .Z(n54878) );
  XOR U54725 ( .A(n54879), .B(n54880), .Z(n54870) );
  AND U54726 ( .A(n54881), .B(n54882), .Z(n54880) );
  XOR U54727 ( .A(n54879), .B(n54561), .Z(n54882) );
  XNOR U54728 ( .A(p_input[719]), .B(n54883), .Z(n54561) );
  AND U54729 ( .A(n1071), .B(n54884), .Z(n54883) );
  XOR U54730 ( .A(p_input[751]), .B(p_input[719]), .Z(n54884) );
  XNOR U54731 ( .A(n54558), .B(n54879), .Z(n54881) );
  XOR U54732 ( .A(n54885), .B(n54886), .Z(n54558) );
  AND U54733 ( .A(n1069), .B(n54887), .Z(n54886) );
  XOR U54734 ( .A(p_input[687]), .B(p_input[655]), .Z(n54887) );
  XOR U54735 ( .A(n54888), .B(n54889), .Z(n54879) );
  AND U54736 ( .A(n54890), .B(n54891), .Z(n54889) );
  XOR U54737 ( .A(n54888), .B(n54573), .Z(n54891) );
  XNOR U54738 ( .A(p_input[718]), .B(n54892), .Z(n54573) );
  AND U54739 ( .A(n1071), .B(n54893), .Z(n54892) );
  XOR U54740 ( .A(p_input[750]), .B(p_input[718]), .Z(n54893) );
  XNOR U54741 ( .A(n54570), .B(n54888), .Z(n54890) );
  XOR U54742 ( .A(n54894), .B(n54895), .Z(n54570) );
  AND U54743 ( .A(n1069), .B(n54896), .Z(n54895) );
  XOR U54744 ( .A(p_input[686]), .B(p_input[654]), .Z(n54896) );
  XOR U54745 ( .A(n54897), .B(n54898), .Z(n54888) );
  AND U54746 ( .A(n54899), .B(n54900), .Z(n54898) );
  XOR U54747 ( .A(n54897), .B(n54585), .Z(n54900) );
  XNOR U54748 ( .A(p_input[717]), .B(n54901), .Z(n54585) );
  AND U54749 ( .A(n1071), .B(n54902), .Z(n54901) );
  XOR U54750 ( .A(p_input[749]), .B(p_input[717]), .Z(n54902) );
  XNOR U54751 ( .A(n54582), .B(n54897), .Z(n54899) );
  XOR U54752 ( .A(n54903), .B(n54904), .Z(n54582) );
  AND U54753 ( .A(n1069), .B(n54905), .Z(n54904) );
  XOR U54754 ( .A(p_input[685]), .B(p_input[653]), .Z(n54905) );
  XOR U54755 ( .A(n54906), .B(n54907), .Z(n54897) );
  AND U54756 ( .A(n54908), .B(n54909), .Z(n54907) );
  XOR U54757 ( .A(n54906), .B(n54597), .Z(n54909) );
  XNOR U54758 ( .A(p_input[716]), .B(n54910), .Z(n54597) );
  AND U54759 ( .A(n1071), .B(n54911), .Z(n54910) );
  XOR U54760 ( .A(p_input[748]), .B(p_input[716]), .Z(n54911) );
  XNOR U54761 ( .A(n54594), .B(n54906), .Z(n54908) );
  XOR U54762 ( .A(n54912), .B(n54913), .Z(n54594) );
  AND U54763 ( .A(n1069), .B(n54914), .Z(n54913) );
  XOR U54764 ( .A(p_input[684]), .B(p_input[652]), .Z(n54914) );
  XOR U54765 ( .A(n54915), .B(n54916), .Z(n54906) );
  AND U54766 ( .A(n54917), .B(n54918), .Z(n54916) );
  XOR U54767 ( .A(n54915), .B(n54609), .Z(n54918) );
  XNOR U54768 ( .A(p_input[715]), .B(n54919), .Z(n54609) );
  AND U54769 ( .A(n1071), .B(n54920), .Z(n54919) );
  XOR U54770 ( .A(p_input[747]), .B(p_input[715]), .Z(n54920) );
  XNOR U54771 ( .A(n54606), .B(n54915), .Z(n54917) );
  XOR U54772 ( .A(n54921), .B(n54922), .Z(n54606) );
  AND U54773 ( .A(n1069), .B(n54923), .Z(n54922) );
  XOR U54774 ( .A(p_input[683]), .B(p_input[651]), .Z(n54923) );
  XOR U54775 ( .A(n54924), .B(n54925), .Z(n54915) );
  AND U54776 ( .A(n54926), .B(n54927), .Z(n54925) );
  XOR U54777 ( .A(n54924), .B(n54621), .Z(n54927) );
  XNOR U54778 ( .A(p_input[714]), .B(n54928), .Z(n54621) );
  AND U54779 ( .A(n1071), .B(n54929), .Z(n54928) );
  XOR U54780 ( .A(p_input[746]), .B(p_input[714]), .Z(n54929) );
  XNOR U54781 ( .A(n54618), .B(n54924), .Z(n54926) );
  XOR U54782 ( .A(n54930), .B(n54931), .Z(n54618) );
  AND U54783 ( .A(n1069), .B(n54932), .Z(n54931) );
  XOR U54784 ( .A(p_input[682]), .B(p_input[650]), .Z(n54932) );
  XOR U54785 ( .A(n54933), .B(n54934), .Z(n54924) );
  AND U54786 ( .A(n54935), .B(n54936), .Z(n54934) );
  XOR U54787 ( .A(n54933), .B(n54633), .Z(n54936) );
  XNOR U54788 ( .A(p_input[713]), .B(n54937), .Z(n54633) );
  AND U54789 ( .A(n1071), .B(n54938), .Z(n54937) );
  XOR U54790 ( .A(p_input[745]), .B(p_input[713]), .Z(n54938) );
  XNOR U54791 ( .A(n54630), .B(n54933), .Z(n54935) );
  XOR U54792 ( .A(n54939), .B(n54940), .Z(n54630) );
  AND U54793 ( .A(n1069), .B(n54941), .Z(n54940) );
  XOR U54794 ( .A(p_input[681]), .B(p_input[649]), .Z(n54941) );
  XOR U54795 ( .A(n54942), .B(n54943), .Z(n54933) );
  AND U54796 ( .A(n54944), .B(n54945), .Z(n54943) );
  XOR U54797 ( .A(n54942), .B(n54645), .Z(n54945) );
  XNOR U54798 ( .A(p_input[712]), .B(n54946), .Z(n54645) );
  AND U54799 ( .A(n1071), .B(n54947), .Z(n54946) );
  XOR U54800 ( .A(p_input[744]), .B(p_input[712]), .Z(n54947) );
  XNOR U54801 ( .A(n54642), .B(n54942), .Z(n54944) );
  XOR U54802 ( .A(n54948), .B(n54949), .Z(n54642) );
  AND U54803 ( .A(n1069), .B(n54950), .Z(n54949) );
  XOR U54804 ( .A(p_input[680]), .B(p_input[648]), .Z(n54950) );
  XOR U54805 ( .A(n54951), .B(n54952), .Z(n54942) );
  AND U54806 ( .A(n54953), .B(n54954), .Z(n54952) );
  XOR U54807 ( .A(n54951), .B(n54657), .Z(n54954) );
  XNOR U54808 ( .A(p_input[711]), .B(n54955), .Z(n54657) );
  AND U54809 ( .A(n1071), .B(n54956), .Z(n54955) );
  XOR U54810 ( .A(p_input[743]), .B(p_input[711]), .Z(n54956) );
  XNOR U54811 ( .A(n54654), .B(n54951), .Z(n54953) );
  XOR U54812 ( .A(n54957), .B(n54958), .Z(n54654) );
  AND U54813 ( .A(n1069), .B(n54959), .Z(n54958) );
  XOR U54814 ( .A(p_input[679]), .B(p_input[647]), .Z(n54959) );
  XOR U54815 ( .A(n54960), .B(n54961), .Z(n54951) );
  AND U54816 ( .A(n54962), .B(n54963), .Z(n54961) );
  XOR U54817 ( .A(n54960), .B(n54669), .Z(n54963) );
  XNOR U54818 ( .A(p_input[710]), .B(n54964), .Z(n54669) );
  AND U54819 ( .A(n1071), .B(n54965), .Z(n54964) );
  XOR U54820 ( .A(p_input[742]), .B(p_input[710]), .Z(n54965) );
  XNOR U54821 ( .A(n54666), .B(n54960), .Z(n54962) );
  XOR U54822 ( .A(n54966), .B(n54967), .Z(n54666) );
  AND U54823 ( .A(n1069), .B(n54968), .Z(n54967) );
  XOR U54824 ( .A(p_input[678]), .B(p_input[646]), .Z(n54968) );
  XOR U54825 ( .A(n54969), .B(n54970), .Z(n54960) );
  AND U54826 ( .A(n54971), .B(n54972), .Z(n54970) );
  XOR U54827 ( .A(n54969), .B(n54681), .Z(n54972) );
  XNOR U54828 ( .A(p_input[709]), .B(n54973), .Z(n54681) );
  AND U54829 ( .A(n1071), .B(n54974), .Z(n54973) );
  XOR U54830 ( .A(p_input[741]), .B(p_input[709]), .Z(n54974) );
  XNOR U54831 ( .A(n54678), .B(n54969), .Z(n54971) );
  XOR U54832 ( .A(n54975), .B(n54976), .Z(n54678) );
  AND U54833 ( .A(n1069), .B(n54977), .Z(n54976) );
  XOR U54834 ( .A(p_input[677]), .B(p_input[645]), .Z(n54977) );
  XOR U54835 ( .A(n54978), .B(n54979), .Z(n54969) );
  AND U54836 ( .A(n54980), .B(n54981), .Z(n54979) );
  XOR U54837 ( .A(n54978), .B(n54693), .Z(n54981) );
  XNOR U54838 ( .A(p_input[708]), .B(n54982), .Z(n54693) );
  AND U54839 ( .A(n1071), .B(n54983), .Z(n54982) );
  XOR U54840 ( .A(p_input[740]), .B(p_input[708]), .Z(n54983) );
  XNOR U54841 ( .A(n54690), .B(n54978), .Z(n54980) );
  XOR U54842 ( .A(n54984), .B(n54985), .Z(n54690) );
  AND U54843 ( .A(n1069), .B(n54986), .Z(n54985) );
  XOR U54844 ( .A(p_input[676]), .B(p_input[644]), .Z(n54986) );
  XOR U54845 ( .A(n54987), .B(n54988), .Z(n54978) );
  AND U54846 ( .A(n54989), .B(n54990), .Z(n54988) );
  XOR U54847 ( .A(n54987), .B(n54705), .Z(n54990) );
  XNOR U54848 ( .A(p_input[707]), .B(n54991), .Z(n54705) );
  AND U54849 ( .A(n1071), .B(n54992), .Z(n54991) );
  XOR U54850 ( .A(p_input[739]), .B(p_input[707]), .Z(n54992) );
  XNOR U54851 ( .A(n54702), .B(n54987), .Z(n54989) );
  XOR U54852 ( .A(n54993), .B(n54994), .Z(n54702) );
  AND U54853 ( .A(n1069), .B(n54995), .Z(n54994) );
  XOR U54854 ( .A(p_input[675]), .B(p_input[643]), .Z(n54995) );
  XOR U54855 ( .A(n54996), .B(n54997), .Z(n54987) );
  AND U54856 ( .A(n54998), .B(n54999), .Z(n54997) );
  XOR U54857 ( .A(n54996), .B(n54717), .Z(n54999) );
  XNOR U54858 ( .A(p_input[706]), .B(n55000), .Z(n54717) );
  AND U54859 ( .A(n1071), .B(n55001), .Z(n55000) );
  XOR U54860 ( .A(p_input[738]), .B(p_input[706]), .Z(n55001) );
  XNOR U54861 ( .A(n54714), .B(n54996), .Z(n54998) );
  XOR U54862 ( .A(n55002), .B(n55003), .Z(n54714) );
  AND U54863 ( .A(n1069), .B(n55004), .Z(n55003) );
  XOR U54864 ( .A(p_input[674]), .B(p_input[642]), .Z(n55004) );
  XOR U54865 ( .A(n55005), .B(n55006), .Z(n54996) );
  AND U54866 ( .A(n55007), .B(n55008), .Z(n55006) );
  XNOR U54867 ( .A(n55009), .B(n54730), .Z(n55008) );
  XNOR U54868 ( .A(p_input[705]), .B(n55010), .Z(n54730) );
  AND U54869 ( .A(n1071), .B(n55011), .Z(n55010) );
  XNOR U54870 ( .A(p_input[737]), .B(n55012), .Z(n55011) );
  IV U54871 ( .A(p_input[705]), .Z(n55012) );
  XNOR U54872 ( .A(n54727), .B(n55005), .Z(n55007) );
  XNOR U54873 ( .A(p_input[641]), .B(n55013), .Z(n54727) );
  AND U54874 ( .A(n1069), .B(n55014), .Z(n55013) );
  XOR U54875 ( .A(p_input[673]), .B(p_input[641]), .Z(n55014) );
  IV U54876 ( .A(n55009), .Z(n55005) );
  AND U54877 ( .A(n54735), .B(n54738), .Z(n55009) );
  XOR U54878 ( .A(p_input[704]), .B(n55015), .Z(n54738) );
  AND U54879 ( .A(n1071), .B(n55016), .Z(n55015) );
  XOR U54880 ( .A(p_input[736]), .B(p_input[704]), .Z(n55016) );
  XOR U54881 ( .A(n55017), .B(n55018), .Z(n1071) );
  AND U54882 ( .A(n55019), .B(n55020), .Z(n55018) );
  XNOR U54883 ( .A(p_input[767]), .B(n55017), .Z(n55020) );
  XOR U54884 ( .A(n55017), .B(p_input[735]), .Z(n55019) );
  XOR U54885 ( .A(n55021), .B(n55022), .Z(n55017) );
  AND U54886 ( .A(n55023), .B(n55024), .Z(n55022) );
  XNOR U54887 ( .A(p_input[766]), .B(n55021), .Z(n55024) );
  XOR U54888 ( .A(n55021), .B(p_input[734]), .Z(n55023) );
  XOR U54889 ( .A(n55025), .B(n55026), .Z(n55021) );
  AND U54890 ( .A(n55027), .B(n55028), .Z(n55026) );
  XNOR U54891 ( .A(p_input[765]), .B(n55025), .Z(n55028) );
  XOR U54892 ( .A(n55025), .B(p_input[733]), .Z(n55027) );
  XOR U54893 ( .A(n55029), .B(n55030), .Z(n55025) );
  AND U54894 ( .A(n55031), .B(n55032), .Z(n55030) );
  XNOR U54895 ( .A(p_input[764]), .B(n55029), .Z(n55032) );
  XOR U54896 ( .A(n55029), .B(p_input[732]), .Z(n55031) );
  XOR U54897 ( .A(n55033), .B(n55034), .Z(n55029) );
  AND U54898 ( .A(n55035), .B(n55036), .Z(n55034) );
  XNOR U54899 ( .A(p_input[763]), .B(n55033), .Z(n55036) );
  XOR U54900 ( .A(n55033), .B(p_input[731]), .Z(n55035) );
  XOR U54901 ( .A(n55037), .B(n55038), .Z(n55033) );
  AND U54902 ( .A(n55039), .B(n55040), .Z(n55038) );
  XNOR U54903 ( .A(p_input[762]), .B(n55037), .Z(n55040) );
  XOR U54904 ( .A(n55037), .B(p_input[730]), .Z(n55039) );
  XOR U54905 ( .A(n55041), .B(n55042), .Z(n55037) );
  AND U54906 ( .A(n55043), .B(n55044), .Z(n55042) );
  XNOR U54907 ( .A(p_input[761]), .B(n55041), .Z(n55044) );
  XOR U54908 ( .A(n55041), .B(p_input[729]), .Z(n55043) );
  XOR U54909 ( .A(n55045), .B(n55046), .Z(n55041) );
  AND U54910 ( .A(n55047), .B(n55048), .Z(n55046) );
  XNOR U54911 ( .A(p_input[760]), .B(n55045), .Z(n55048) );
  XOR U54912 ( .A(n55045), .B(p_input[728]), .Z(n55047) );
  XOR U54913 ( .A(n55049), .B(n55050), .Z(n55045) );
  AND U54914 ( .A(n55051), .B(n55052), .Z(n55050) );
  XNOR U54915 ( .A(p_input[759]), .B(n55049), .Z(n55052) );
  XOR U54916 ( .A(n55049), .B(p_input[727]), .Z(n55051) );
  XOR U54917 ( .A(n55053), .B(n55054), .Z(n55049) );
  AND U54918 ( .A(n55055), .B(n55056), .Z(n55054) );
  XNOR U54919 ( .A(p_input[758]), .B(n55053), .Z(n55056) );
  XOR U54920 ( .A(n55053), .B(p_input[726]), .Z(n55055) );
  XOR U54921 ( .A(n55057), .B(n55058), .Z(n55053) );
  AND U54922 ( .A(n55059), .B(n55060), .Z(n55058) );
  XNOR U54923 ( .A(p_input[757]), .B(n55057), .Z(n55060) );
  XOR U54924 ( .A(n55057), .B(p_input[725]), .Z(n55059) );
  XOR U54925 ( .A(n55061), .B(n55062), .Z(n55057) );
  AND U54926 ( .A(n55063), .B(n55064), .Z(n55062) );
  XNOR U54927 ( .A(p_input[756]), .B(n55061), .Z(n55064) );
  XOR U54928 ( .A(n55061), .B(p_input[724]), .Z(n55063) );
  XOR U54929 ( .A(n55065), .B(n55066), .Z(n55061) );
  AND U54930 ( .A(n55067), .B(n55068), .Z(n55066) );
  XNOR U54931 ( .A(p_input[755]), .B(n55065), .Z(n55068) );
  XOR U54932 ( .A(n55065), .B(p_input[723]), .Z(n55067) );
  XOR U54933 ( .A(n55069), .B(n55070), .Z(n55065) );
  AND U54934 ( .A(n55071), .B(n55072), .Z(n55070) );
  XNOR U54935 ( .A(p_input[754]), .B(n55069), .Z(n55072) );
  XOR U54936 ( .A(n55069), .B(p_input[722]), .Z(n55071) );
  XOR U54937 ( .A(n55073), .B(n55074), .Z(n55069) );
  AND U54938 ( .A(n55075), .B(n55076), .Z(n55074) );
  XNOR U54939 ( .A(p_input[753]), .B(n55073), .Z(n55076) );
  XOR U54940 ( .A(n55073), .B(p_input[721]), .Z(n55075) );
  XOR U54941 ( .A(n55077), .B(n55078), .Z(n55073) );
  AND U54942 ( .A(n55079), .B(n55080), .Z(n55078) );
  XNOR U54943 ( .A(p_input[752]), .B(n55077), .Z(n55080) );
  XOR U54944 ( .A(n55077), .B(p_input[720]), .Z(n55079) );
  XOR U54945 ( .A(n55081), .B(n55082), .Z(n55077) );
  AND U54946 ( .A(n55083), .B(n55084), .Z(n55082) );
  XNOR U54947 ( .A(p_input[751]), .B(n55081), .Z(n55084) );
  XOR U54948 ( .A(n55081), .B(p_input[719]), .Z(n55083) );
  XOR U54949 ( .A(n55085), .B(n55086), .Z(n55081) );
  AND U54950 ( .A(n55087), .B(n55088), .Z(n55086) );
  XNOR U54951 ( .A(p_input[750]), .B(n55085), .Z(n55088) );
  XOR U54952 ( .A(n55085), .B(p_input[718]), .Z(n55087) );
  XOR U54953 ( .A(n55089), .B(n55090), .Z(n55085) );
  AND U54954 ( .A(n55091), .B(n55092), .Z(n55090) );
  XNOR U54955 ( .A(p_input[749]), .B(n55089), .Z(n55092) );
  XOR U54956 ( .A(n55089), .B(p_input[717]), .Z(n55091) );
  XOR U54957 ( .A(n55093), .B(n55094), .Z(n55089) );
  AND U54958 ( .A(n55095), .B(n55096), .Z(n55094) );
  XNOR U54959 ( .A(p_input[748]), .B(n55093), .Z(n55096) );
  XOR U54960 ( .A(n55093), .B(p_input[716]), .Z(n55095) );
  XOR U54961 ( .A(n55097), .B(n55098), .Z(n55093) );
  AND U54962 ( .A(n55099), .B(n55100), .Z(n55098) );
  XNOR U54963 ( .A(p_input[747]), .B(n55097), .Z(n55100) );
  XOR U54964 ( .A(n55097), .B(p_input[715]), .Z(n55099) );
  XOR U54965 ( .A(n55101), .B(n55102), .Z(n55097) );
  AND U54966 ( .A(n55103), .B(n55104), .Z(n55102) );
  XNOR U54967 ( .A(p_input[746]), .B(n55101), .Z(n55104) );
  XOR U54968 ( .A(n55101), .B(p_input[714]), .Z(n55103) );
  XOR U54969 ( .A(n55105), .B(n55106), .Z(n55101) );
  AND U54970 ( .A(n55107), .B(n55108), .Z(n55106) );
  XNOR U54971 ( .A(p_input[745]), .B(n55105), .Z(n55108) );
  XOR U54972 ( .A(n55105), .B(p_input[713]), .Z(n55107) );
  XOR U54973 ( .A(n55109), .B(n55110), .Z(n55105) );
  AND U54974 ( .A(n55111), .B(n55112), .Z(n55110) );
  XNOR U54975 ( .A(p_input[744]), .B(n55109), .Z(n55112) );
  XOR U54976 ( .A(n55109), .B(p_input[712]), .Z(n55111) );
  XOR U54977 ( .A(n55113), .B(n55114), .Z(n55109) );
  AND U54978 ( .A(n55115), .B(n55116), .Z(n55114) );
  XNOR U54979 ( .A(p_input[743]), .B(n55113), .Z(n55116) );
  XOR U54980 ( .A(n55113), .B(p_input[711]), .Z(n55115) );
  XOR U54981 ( .A(n55117), .B(n55118), .Z(n55113) );
  AND U54982 ( .A(n55119), .B(n55120), .Z(n55118) );
  XNOR U54983 ( .A(p_input[742]), .B(n55117), .Z(n55120) );
  XOR U54984 ( .A(n55117), .B(p_input[710]), .Z(n55119) );
  XOR U54985 ( .A(n55121), .B(n55122), .Z(n55117) );
  AND U54986 ( .A(n55123), .B(n55124), .Z(n55122) );
  XNOR U54987 ( .A(p_input[741]), .B(n55121), .Z(n55124) );
  XOR U54988 ( .A(n55121), .B(p_input[709]), .Z(n55123) );
  XOR U54989 ( .A(n55125), .B(n55126), .Z(n55121) );
  AND U54990 ( .A(n55127), .B(n55128), .Z(n55126) );
  XNOR U54991 ( .A(p_input[740]), .B(n55125), .Z(n55128) );
  XOR U54992 ( .A(n55125), .B(p_input[708]), .Z(n55127) );
  XOR U54993 ( .A(n55129), .B(n55130), .Z(n55125) );
  AND U54994 ( .A(n55131), .B(n55132), .Z(n55130) );
  XNOR U54995 ( .A(p_input[739]), .B(n55129), .Z(n55132) );
  XOR U54996 ( .A(n55129), .B(p_input[707]), .Z(n55131) );
  XOR U54997 ( .A(n55133), .B(n55134), .Z(n55129) );
  AND U54998 ( .A(n55135), .B(n55136), .Z(n55134) );
  XNOR U54999 ( .A(p_input[738]), .B(n55133), .Z(n55136) );
  XOR U55000 ( .A(n55133), .B(p_input[706]), .Z(n55135) );
  XNOR U55001 ( .A(n55137), .B(n55138), .Z(n55133) );
  AND U55002 ( .A(n55139), .B(n55140), .Z(n55138) );
  XOR U55003 ( .A(p_input[737]), .B(n55137), .Z(n55140) );
  XNOR U55004 ( .A(p_input[705]), .B(n55137), .Z(n55139) );
  AND U55005 ( .A(p_input[736]), .B(n55141), .Z(n55137) );
  IV U55006 ( .A(p_input[704]), .Z(n55141) );
  XNOR U55007 ( .A(p_input[640]), .B(n55142), .Z(n54735) );
  AND U55008 ( .A(n1069), .B(n55143), .Z(n55142) );
  XOR U55009 ( .A(p_input[672]), .B(p_input[640]), .Z(n55143) );
  XOR U55010 ( .A(n55144), .B(n55145), .Z(n1069) );
  AND U55011 ( .A(n55146), .B(n55147), .Z(n55145) );
  XNOR U55012 ( .A(p_input[703]), .B(n55144), .Z(n55147) );
  XOR U55013 ( .A(n55144), .B(p_input[671]), .Z(n55146) );
  XOR U55014 ( .A(n55148), .B(n55149), .Z(n55144) );
  AND U55015 ( .A(n55150), .B(n55151), .Z(n55149) );
  XNOR U55016 ( .A(p_input[702]), .B(n55148), .Z(n55151) );
  XNOR U55017 ( .A(n55148), .B(n54750), .Z(n55150) );
  IV U55018 ( .A(p_input[670]), .Z(n54750) );
  XOR U55019 ( .A(n55152), .B(n55153), .Z(n55148) );
  AND U55020 ( .A(n55154), .B(n55155), .Z(n55153) );
  XNOR U55021 ( .A(p_input[701]), .B(n55152), .Z(n55155) );
  XNOR U55022 ( .A(n55152), .B(n54759), .Z(n55154) );
  IV U55023 ( .A(p_input[669]), .Z(n54759) );
  XOR U55024 ( .A(n55156), .B(n55157), .Z(n55152) );
  AND U55025 ( .A(n55158), .B(n55159), .Z(n55157) );
  XNOR U55026 ( .A(p_input[700]), .B(n55156), .Z(n55159) );
  XNOR U55027 ( .A(n55156), .B(n54768), .Z(n55158) );
  IV U55028 ( .A(p_input[668]), .Z(n54768) );
  XOR U55029 ( .A(n55160), .B(n55161), .Z(n55156) );
  AND U55030 ( .A(n55162), .B(n55163), .Z(n55161) );
  XNOR U55031 ( .A(p_input[699]), .B(n55160), .Z(n55163) );
  XNOR U55032 ( .A(n55160), .B(n54777), .Z(n55162) );
  IV U55033 ( .A(p_input[667]), .Z(n54777) );
  XOR U55034 ( .A(n55164), .B(n55165), .Z(n55160) );
  AND U55035 ( .A(n55166), .B(n55167), .Z(n55165) );
  XNOR U55036 ( .A(p_input[698]), .B(n55164), .Z(n55167) );
  XNOR U55037 ( .A(n55164), .B(n54786), .Z(n55166) );
  IV U55038 ( .A(p_input[666]), .Z(n54786) );
  XOR U55039 ( .A(n55168), .B(n55169), .Z(n55164) );
  AND U55040 ( .A(n55170), .B(n55171), .Z(n55169) );
  XNOR U55041 ( .A(p_input[697]), .B(n55168), .Z(n55171) );
  XNOR U55042 ( .A(n55168), .B(n54795), .Z(n55170) );
  IV U55043 ( .A(p_input[665]), .Z(n54795) );
  XOR U55044 ( .A(n55172), .B(n55173), .Z(n55168) );
  AND U55045 ( .A(n55174), .B(n55175), .Z(n55173) );
  XNOR U55046 ( .A(p_input[696]), .B(n55172), .Z(n55175) );
  XNOR U55047 ( .A(n55172), .B(n54804), .Z(n55174) );
  IV U55048 ( .A(p_input[664]), .Z(n54804) );
  XOR U55049 ( .A(n55176), .B(n55177), .Z(n55172) );
  AND U55050 ( .A(n55178), .B(n55179), .Z(n55177) );
  XNOR U55051 ( .A(p_input[695]), .B(n55176), .Z(n55179) );
  XNOR U55052 ( .A(n55176), .B(n54813), .Z(n55178) );
  IV U55053 ( .A(p_input[663]), .Z(n54813) );
  XOR U55054 ( .A(n55180), .B(n55181), .Z(n55176) );
  AND U55055 ( .A(n55182), .B(n55183), .Z(n55181) );
  XNOR U55056 ( .A(p_input[694]), .B(n55180), .Z(n55183) );
  XNOR U55057 ( .A(n55180), .B(n54822), .Z(n55182) );
  IV U55058 ( .A(p_input[662]), .Z(n54822) );
  XOR U55059 ( .A(n55184), .B(n55185), .Z(n55180) );
  AND U55060 ( .A(n55186), .B(n55187), .Z(n55185) );
  XNOR U55061 ( .A(p_input[693]), .B(n55184), .Z(n55187) );
  XNOR U55062 ( .A(n55184), .B(n54831), .Z(n55186) );
  IV U55063 ( .A(p_input[661]), .Z(n54831) );
  XOR U55064 ( .A(n55188), .B(n55189), .Z(n55184) );
  AND U55065 ( .A(n55190), .B(n55191), .Z(n55189) );
  XNOR U55066 ( .A(p_input[692]), .B(n55188), .Z(n55191) );
  XNOR U55067 ( .A(n55188), .B(n54840), .Z(n55190) );
  IV U55068 ( .A(p_input[660]), .Z(n54840) );
  XOR U55069 ( .A(n55192), .B(n55193), .Z(n55188) );
  AND U55070 ( .A(n55194), .B(n55195), .Z(n55193) );
  XNOR U55071 ( .A(p_input[691]), .B(n55192), .Z(n55195) );
  XNOR U55072 ( .A(n55192), .B(n54849), .Z(n55194) );
  IV U55073 ( .A(p_input[659]), .Z(n54849) );
  XOR U55074 ( .A(n55196), .B(n55197), .Z(n55192) );
  AND U55075 ( .A(n55198), .B(n55199), .Z(n55197) );
  XNOR U55076 ( .A(p_input[690]), .B(n55196), .Z(n55199) );
  XNOR U55077 ( .A(n55196), .B(n54858), .Z(n55198) );
  IV U55078 ( .A(p_input[658]), .Z(n54858) );
  XOR U55079 ( .A(n55200), .B(n55201), .Z(n55196) );
  AND U55080 ( .A(n55202), .B(n55203), .Z(n55201) );
  XNOR U55081 ( .A(p_input[689]), .B(n55200), .Z(n55203) );
  XNOR U55082 ( .A(n55200), .B(n54867), .Z(n55202) );
  IV U55083 ( .A(p_input[657]), .Z(n54867) );
  XOR U55084 ( .A(n55204), .B(n55205), .Z(n55200) );
  AND U55085 ( .A(n55206), .B(n55207), .Z(n55205) );
  XNOR U55086 ( .A(p_input[688]), .B(n55204), .Z(n55207) );
  XNOR U55087 ( .A(n55204), .B(n54876), .Z(n55206) );
  IV U55088 ( .A(p_input[656]), .Z(n54876) );
  XOR U55089 ( .A(n55208), .B(n55209), .Z(n55204) );
  AND U55090 ( .A(n55210), .B(n55211), .Z(n55209) );
  XNOR U55091 ( .A(p_input[687]), .B(n55208), .Z(n55211) );
  XNOR U55092 ( .A(n55208), .B(n54885), .Z(n55210) );
  IV U55093 ( .A(p_input[655]), .Z(n54885) );
  XOR U55094 ( .A(n55212), .B(n55213), .Z(n55208) );
  AND U55095 ( .A(n55214), .B(n55215), .Z(n55213) );
  XNOR U55096 ( .A(p_input[686]), .B(n55212), .Z(n55215) );
  XNOR U55097 ( .A(n55212), .B(n54894), .Z(n55214) );
  IV U55098 ( .A(p_input[654]), .Z(n54894) );
  XOR U55099 ( .A(n55216), .B(n55217), .Z(n55212) );
  AND U55100 ( .A(n55218), .B(n55219), .Z(n55217) );
  XNOR U55101 ( .A(p_input[685]), .B(n55216), .Z(n55219) );
  XNOR U55102 ( .A(n55216), .B(n54903), .Z(n55218) );
  IV U55103 ( .A(p_input[653]), .Z(n54903) );
  XOR U55104 ( .A(n55220), .B(n55221), .Z(n55216) );
  AND U55105 ( .A(n55222), .B(n55223), .Z(n55221) );
  XNOR U55106 ( .A(p_input[684]), .B(n55220), .Z(n55223) );
  XNOR U55107 ( .A(n55220), .B(n54912), .Z(n55222) );
  IV U55108 ( .A(p_input[652]), .Z(n54912) );
  XOR U55109 ( .A(n55224), .B(n55225), .Z(n55220) );
  AND U55110 ( .A(n55226), .B(n55227), .Z(n55225) );
  XNOR U55111 ( .A(p_input[683]), .B(n55224), .Z(n55227) );
  XNOR U55112 ( .A(n55224), .B(n54921), .Z(n55226) );
  IV U55113 ( .A(p_input[651]), .Z(n54921) );
  XOR U55114 ( .A(n55228), .B(n55229), .Z(n55224) );
  AND U55115 ( .A(n55230), .B(n55231), .Z(n55229) );
  XNOR U55116 ( .A(p_input[682]), .B(n55228), .Z(n55231) );
  XNOR U55117 ( .A(n55228), .B(n54930), .Z(n55230) );
  IV U55118 ( .A(p_input[650]), .Z(n54930) );
  XOR U55119 ( .A(n55232), .B(n55233), .Z(n55228) );
  AND U55120 ( .A(n55234), .B(n55235), .Z(n55233) );
  XNOR U55121 ( .A(p_input[681]), .B(n55232), .Z(n55235) );
  XNOR U55122 ( .A(n55232), .B(n54939), .Z(n55234) );
  IV U55123 ( .A(p_input[649]), .Z(n54939) );
  XOR U55124 ( .A(n55236), .B(n55237), .Z(n55232) );
  AND U55125 ( .A(n55238), .B(n55239), .Z(n55237) );
  XNOR U55126 ( .A(p_input[680]), .B(n55236), .Z(n55239) );
  XNOR U55127 ( .A(n55236), .B(n54948), .Z(n55238) );
  IV U55128 ( .A(p_input[648]), .Z(n54948) );
  XOR U55129 ( .A(n55240), .B(n55241), .Z(n55236) );
  AND U55130 ( .A(n55242), .B(n55243), .Z(n55241) );
  XNOR U55131 ( .A(p_input[679]), .B(n55240), .Z(n55243) );
  XNOR U55132 ( .A(n55240), .B(n54957), .Z(n55242) );
  IV U55133 ( .A(p_input[647]), .Z(n54957) );
  XOR U55134 ( .A(n55244), .B(n55245), .Z(n55240) );
  AND U55135 ( .A(n55246), .B(n55247), .Z(n55245) );
  XNOR U55136 ( .A(p_input[678]), .B(n55244), .Z(n55247) );
  XNOR U55137 ( .A(n55244), .B(n54966), .Z(n55246) );
  IV U55138 ( .A(p_input[646]), .Z(n54966) );
  XOR U55139 ( .A(n55248), .B(n55249), .Z(n55244) );
  AND U55140 ( .A(n55250), .B(n55251), .Z(n55249) );
  XNOR U55141 ( .A(p_input[677]), .B(n55248), .Z(n55251) );
  XNOR U55142 ( .A(n55248), .B(n54975), .Z(n55250) );
  IV U55143 ( .A(p_input[645]), .Z(n54975) );
  XOR U55144 ( .A(n55252), .B(n55253), .Z(n55248) );
  AND U55145 ( .A(n55254), .B(n55255), .Z(n55253) );
  XNOR U55146 ( .A(p_input[676]), .B(n55252), .Z(n55255) );
  XNOR U55147 ( .A(n55252), .B(n54984), .Z(n55254) );
  IV U55148 ( .A(p_input[644]), .Z(n54984) );
  XOR U55149 ( .A(n55256), .B(n55257), .Z(n55252) );
  AND U55150 ( .A(n55258), .B(n55259), .Z(n55257) );
  XNOR U55151 ( .A(p_input[675]), .B(n55256), .Z(n55259) );
  XNOR U55152 ( .A(n55256), .B(n54993), .Z(n55258) );
  IV U55153 ( .A(p_input[643]), .Z(n54993) );
  XOR U55154 ( .A(n55260), .B(n55261), .Z(n55256) );
  AND U55155 ( .A(n55262), .B(n55263), .Z(n55261) );
  XNOR U55156 ( .A(p_input[674]), .B(n55260), .Z(n55263) );
  XNOR U55157 ( .A(n55260), .B(n55002), .Z(n55262) );
  IV U55158 ( .A(p_input[642]), .Z(n55002) );
  XNOR U55159 ( .A(n55264), .B(n55265), .Z(n55260) );
  AND U55160 ( .A(n55266), .B(n55267), .Z(n55265) );
  XOR U55161 ( .A(p_input[673]), .B(n55264), .Z(n55267) );
  XNOR U55162 ( .A(p_input[641]), .B(n55264), .Z(n55266) );
  AND U55163 ( .A(p_input[672]), .B(n55268), .Z(n55264) );
  IV U55164 ( .A(p_input[640]), .Z(n55268) );
  XOR U55165 ( .A(n55269), .B(n55270), .Z(n54358) );
  AND U55166 ( .A(n652), .B(n55271), .Z(n55270) );
  XNOR U55167 ( .A(n55272), .B(n55269), .Z(n55271) );
  XOR U55168 ( .A(n55273), .B(n55274), .Z(n652) );
  AND U55169 ( .A(n55275), .B(n55276), .Z(n55274) );
  XNOR U55170 ( .A(n54373), .B(n55273), .Z(n55276) );
  AND U55171 ( .A(p_input[639]), .B(p_input[607]), .Z(n54373) );
  XNOR U55172 ( .A(n55273), .B(n54370), .Z(n55275) );
  IV U55173 ( .A(n55277), .Z(n54370) );
  AND U55174 ( .A(p_input[543]), .B(p_input[575]), .Z(n55277) );
  XOR U55175 ( .A(n55278), .B(n55279), .Z(n55273) );
  AND U55176 ( .A(n55280), .B(n55281), .Z(n55279) );
  XOR U55177 ( .A(n55278), .B(n54385), .Z(n55281) );
  XNOR U55178 ( .A(p_input[606]), .B(n55282), .Z(n54385) );
  AND U55179 ( .A(n1075), .B(n55283), .Z(n55282) );
  XOR U55180 ( .A(p_input[638]), .B(p_input[606]), .Z(n55283) );
  XNOR U55181 ( .A(n54382), .B(n55278), .Z(n55280) );
  XOR U55182 ( .A(n55284), .B(n55285), .Z(n54382) );
  AND U55183 ( .A(n1072), .B(n55286), .Z(n55285) );
  XOR U55184 ( .A(p_input[574]), .B(p_input[542]), .Z(n55286) );
  XOR U55185 ( .A(n55287), .B(n55288), .Z(n55278) );
  AND U55186 ( .A(n55289), .B(n55290), .Z(n55288) );
  XOR U55187 ( .A(n55287), .B(n54397), .Z(n55290) );
  XNOR U55188 ( .A(p_input[605]), .B(n55291), .Z(n54397) );
  AND U55189 ( .A(n1075), .B(n55292), .Z(n55291) );
  XOR U55190 ( .A(p_input[637]), .B(p_input[605]), .Z(n55292) );
  XNOR U55191 ( .A(n54394), .B(n55287), .Z(n55289) );
  XOR U55192 ( .A(n55293), .B(n55294), .Z(n54394) );
  AND U55193 ( .A(n1072), .B(n55295), .Z(n55294) );
  XOR U55194 ( .A(p_input[573]), .B(p_input[541]), .Z(n55295) );
  XOR U55195 ( .A(n55296), .B(n55297), .Z(n55287) );
  AND U55196 ( .A(n55298), .B(n55299), .Z(n55297) );
  XOR U55197 ( .A(n55296), .B(n54409), .Z(n55299) );
  XNOR U55198 ( .A(p_input[604]), .B(n55300), .Z(n54409) );
  AND U55199 ( .A(n1075), .B(n55301), .Z(n55300) );
  XOR U55200 ( .A(p_input[636]), .B(p_input[604]), .Z(n55301) );
  XNOR U55201 ( .A(n54406), .B(n55296), .Z(n55298) );
  XOR U55202 ( .A(n55302), .B(n55303), .Z(n54406) );
  AND U55203 ( .A(n1072), .B(n55304), .Z(n55303) );
  XOR U55204 ( .A(p_input[572]), .B(p_input[540]), .Z(n55304) );
  XOR U55205 ( .A(n55305), .B(n55306), .Z(n55296) );
  AND U55206 ( .A(n55307), .B(n55308), .Z(n55306) );
  XOR U55207 ( .A(n55305), .B(n54421), .Z(n55308) );
  XNOR U55208 ( .A(p_input[603]), .B(n55309), .Z(n54421) );
  AND U55209 ( .A(n1075), .B(n55310), .Z(n55309) );
  XOR U55210 ( .A(p_input[635]), .B(p_input[603]), .Z(n55310) );
  XNOR U55211 ( .A(n54418), .B(n55305), .Z(n55307) );
  XOR U55212 ( .A(n55311), .B(n55312), .Z(n54418) );
  AND U55213 ( .A(n1072), .B(n55313), .Z(n55312) );
  XOR U55214 ( .A(p_input[571]), .B(p_input[539]), .Z(n55313) );
  XOR U55215 ( .A(n55314), .B(n55315), .Z(n55305) );
  AND U55216 ( .A(n55316), .B(n55317), .Z(n55315) );
  XOR U55217 ( .A(n55314), .B(n54433), .Z(n55317) );
  XNOR U55218 ( .A(p_input[602]), .B(n55318), .Z(n54433) );
  AND U55219 ( .A(n1075), .B(n55319), .Z(n55318) );
  XOR U55220 ( .A(p_input[634]), .B(p_input[602]), .Z(n55319) );
  XNOR U55221 ( .A(n54430), .B(n55314), .Z(n55316) );
  XOR U55222 ( .A(n55320), .B(n55321), .Z(n54430) );
  AND U55223 ( .A(n1072), .B(n55322), .Z(n55321) );
  XOR U55224 ( .A(p_input[570]), .B(p_input[538]), .Z(n55322) );
  XOR U55225 ( .A(n55323), .B(n55324), .Z(n55314) );
  AND U55226 ( .A(n55325), .B(n55326), .Z(n55324) );
  XOR U55227 ( .A(n55323), .B(n54445), .Z(n55326) );
  XNOR U55228 ( .A(p_input[601]), .B(n55327), .Z(n54445) );
  AND U55229 ( .A(n1075), .B(n55328), .Z(n55327) );
  XOR U55230 ( .A(p_input[633]), .B(p_input[601]), .Z(n55328) );
  XNOR U55231 ( .A(n54442), .B(n55323), .Z(n55325) );
  XOR U55232 ( .A(n55329), .B(n55330), .Z(n54442) );
  AND U55233 ( .A(n1072), .B(n55331), .Z(n55330) );
  XOR U55234 ( .A(p_input[569]), .B(p_input[537]), .Z(n55331) );
  XOR U55235 ( .A(n55332), .B(n55333), .Z(n55323) );
  AND U55236 ( .A(n55334), .B(n55335), .Z(n55333) );
  XOR U55237 ( .A(n55332), .B(n54457), .Z(n55335) );
  XNOR U55238 ( .A(p_input[600]), .B(n55336), .Z(n54457) );
  AND U55239 ( .A(n1075), .B(n55337), .Z(n55336) );
  XOR U55240 ( .A(p_input[632]), .B(p_input[600]), .Z(n55337) );
  XNOR U55241 ( .A(n54454), .B(n55332), .Z(n55334) );
  XOR U55242 ( .A(n55338), .B(n55339), .Z(n54454) );
  AND U55243 ( .A(n1072), .B(n55340), .Z(n55339) );
  XOR U55244 ( .A(p_input[568]), .B(p_input[536]), .Z(n55340) );
  XOR U55245 ( .A(n55341), .B(n55342), .Z(n55332) );
  AND U55246 ( .A(n55343), .B(n55344), .Z(n55342) );
  XOR U55247 ( .A(n55341), .B(n54469), .Z(n55344) );
  XNOR U55248 ( .A(p_input[599]), .B(n55345), .Z(n54469) );
  AND U55249 ( .A(n1075), .B(n55346), .Z(n55345) );
  XOR U55250 ( .A(p_input[631]), .B(p_input[599]), .Z(n55346) );
  XNOR U55251 ( .A(n54466), .B(n55341), .Z(n55343) );
  XOR U55252 ( .A(n55347), .B(n55348), .Z(n54466) );
  AND U55253 ( .A(n1072), .B(n55349), .Z(n55348) );
  XOR U55254 ( .A(p_input[567]), .B(p_input[535]), .Z(n55349) );
  XOR U55255 ( .A(n55350), .B(n55351), .Z(n55341) );
  AND U55256 ( .A(n55352), .B(n55353), .Z(n55351) );
  XOR U55257 ( .A(n55350), .B(n54481), .Z(n55353) );
  XNOR U55258 ( .A(p_input[598]), .B(n55354), .Z(n54481) );
  AND U55259 ( .A(n1075), .B(n55355), .Z(n55354) );
  XOR U55260 ( .A(p_input[630]), .B(p_input[598]), .Z(n55355) );
  XNOR U55261 ( .A(n54478), .B(n55350), .Z(n55352) );
  XOR U55262 ( .A(n55356), .B(n55357), .Z(n54478) );
  AND U55263 ( .A(n1072), .B(n55358), .Z(n55357) );
  XOR U55264 ( .A(p_input[566]), .B(p_input[534]), .Z(n55358) );
  XOR U55265 ( .A(n55359), .B(n55360), .Z(n55350) );
  AND U55266 ( .A(n55361), .B(n55362), .Z(n55360) );
  XOR U55267 ( .A(n55359), .B(n54493), .Z(n55362) );
  XNOR U55268 ( .A(p_input[597]), .B(n55363), .Z(n54493) );
  AND U55269 ( .A(n1075), .B(n55364), .Z(n55363) );
  XOR U55270 ( .A(p_input[629]), .B(p_input[597]), .Z(n55364) );
  XNOR U55271 ( .A(n54490), .B(n55359), .Z(n55361) );
  XOR U55272 ( .A(n55365), .B(n55366), .Z(n54490) );
  AND U55273 ( .A(n1072), .B(n55367), .Z(n55366) );
  XOR U55274 ( .A(p_input[565]), .B(p_input[533]), .Z(n55367) );
  XOR U55275 ( .A(n55368), .B(n55369), .Z(n55359) );
  AND U55276 ( .A(n55370), .B(n55371), .Z(n55369) );
  XOR U55277 ( .A(n55368), .B(n54505), .Z(n55371) );
  XNOR U55278 ( .A(p_input[596]), .B(n55372), .Z(n54505) );
  AND U55279 ( .A(n1075), .B(n55373), .Z(n55372) );
  XOR U55280 ( .A(p_input[628]), .B(p_input[596]), .Z(n55373) );
  XNOR U55281 ( .A(n54502), .B(n55368), .Z(n55370) );
  XOR U55282 ( .A(n55374), .B(n55375), .Z(n54502) );
  AND U55283 ( .A(n1072), .B(n55376), .Z(n55375) );
  XOR U55284 ( .A(p_input[564]), .B(p_input[532]), .Z(n55376) );
  XOR U55285 ( .A(n55377), .B(n55378), .Z(n55368) );
  AND U55286 ( .A(n55379), .B(n55380), .Z(n55378) );
  XOR U55287 ( .A(n55377), .B(n54517), .Z(n55380) );
  XNOR U55288 ( .A(p_input[595]), .B(n55381), .Z(n54517) );
  AND U55289 ( .A(n1075), .B(n55382), .Z(n55381) );
  XOR U55290 ( .A(p_input[627]), .B(p_input[595]), .Z(n55382) );
  XNOR U55291 ( .A(n54514), .B(n55377), .Z(n55379) );
  XOR U55292 ( .A(n55383), .B(n55384), .Z(n54514) );
  AND U55293 ( .A(n1072), .B(n55385), .Z(n55384) );
  XOR U55294 ( .A(p_input[563]), .B(p_input[531]), .Z(n55385) );
  XOR U55295 ( .A(n55386), .B(n55387), .Z(n55377) );
  AND U55296 ( .A(n55388), .B(n55389), .Z(n55387) );
  XOR U55297 ( .A(n55386), .B(n54529), .Z(n55389) );
  XNOR U55298 ( .A(p_input[594]), .B(n55390), .Z(n54529) );
  AND U55299 ( .A(n1075), .B(n55391), .Z(n55390) );
  XOR U55300 ( .A(p_input[626]), .B(p_input[594]), .Z(n55391) );
  XNOR U55301 ( .A(n54526), .B(n55386), .Z(n55388) );
  XOR U55302 ( .A(n55392), .B(n55393), .Z(n54526) );
  AND U55303 ( .A(n1072), .B(n55394), .Z(n55393) );
  XOR U55304 ( .A(p_input[562]), .B(p_input[530]), .Z(n55394) );
  XOR U55305 ( .A(n55395), .B(n55396), .Z(n55386) );
  AND U55306 ( .A(n55397), .B(n55398), .Z(n55396) );
  XOR U55307 ( .A(n55395), .B(n54541), .Z(n55398) );
  XNOR U55308 ( .A(p_input[593]), .B(n55399), .Z(n54541) );
  AND U55309 ( .A(n1075), .B(n55400), .Z(n55399) );
  XOR U55310 ( .A(p_input[625]), .B(p_input[593]), .Z(n55400) );
  XNOR U55311 ( .A(n54538), .B(n55395), .Z(n55397) );
  XOR U55312 ( .A(n55401), .B(n55402), .Z(n54538) );
  AND U55313 ( .A(n1072), .B(n55403), .Z(n55402) );
  XOR U55314 ( .A(p_input[561]), .B(p_input[529]), .Z(n55403) );
  XOR U55315 ( .A(n55404), .B(n55405), .Z(n55395) );
  AND U55316 ( .A(n55406), .B(n55407), .Z(n55405) );
  XOR U55317 ( .A(n55404), .B(n54553), .Z(n55407) );
  XNOR U55318 ( .A(p_input[592]), .B(n55408), .Z(n54553) );
  AND U55319 ( .A(n1075), .B(n55409), .Z(n55408) );
  XOR U55320 ( .A(p_input[624]), .B(p_input[592]), .Z(n55409) );
  XNOR U55321 ( .A(n54550), .B(n55404), .Z(n55406) );
  XOR U55322 ( .A(n55410), .B(n55411), .Z(n54550) );
  AND U55323 ( .A(n1072), .B(n55412), .Z(n55411) );
  XOR U55324 ( .A(p_input[560]), .B(p_input[528]), .Z(n55412) );
  XOR U55325 ( .A(n55413), .B(n55414), .Z(n55404) );
  AND U55326 ( .A(n55415), .B(n55416), .Z(n55414) );
  XOR U55327 ( .A(n55413), .B(n54565), .Z(n55416) );
  XNOR U55328 ( .A(p_input[591]), .B(n55417), .Z(n54565) );
  AND U55329 ( .A(n1075), .B(n55418), .Z(n55417) );
  XOR U55330 ( .A(p_input[623]), .B(p_input[591]), .Z(n55418) );
  XNOR U55331 ( .A(n54562), .B(n55413), .Z(n55415) );
  XOR U55332 ( .A(n55419), .B(n55420), .Z(n54562) );
  AND U55333 ( .A(n1072), .B(n55421), .Z(n55420) );
  XOR U55334 ( .A(p_input[559]), .B(p_input[527]), .Z(n55421) );
  XOR U55335 ( .A(n55422), .B(n55423), .Z(n55413) );
  AND U55336 ( .A(n55424), .B(n55425), .Z(n55423) );
  XOR U55337 ( .A(n55422), .B(n54577), .Z(n55425) );
  XNOR U55338 ( .A(p_input[590]), .B(n55426), .Z(n54577) );
  AND U55339 ( .A(n1075), .B(n55427), .Z(n55426) );
  XOR U55340 ( .A(p_input[622]), .B(p_input[590]), .Z(n55427) );
  XNOR U55341 ( .A(n54574), .B(n55422), .Z(n55424) );
  XOR U55342 ( .A(n55428), .B(n55429), .Z(n54574) );
  AND U55343 ( .A(n1072), .B(n55430), .Z(n55429) );
  XOR U55344 ( .A(p_input[558]), .B(p_input[526]), .Z(n55430) );
  XOR U55345 ( .A(n55431), .B(n55432), .Z(n55422) );
  AND U55346 ( .A(n55433), .B(n55434), .Z(n55432) );
  XOR U55347 ( .A(n55431), .B(n54589), .Z(n55434) );
  XNOR U55348 ( .A(p_input[589]), .B(n55435), .Z(n54589) );
  AND U55349 ( .A(n1075), .B(n55436), .Z(n55435) );
  XOR U55350 ( .A(p_input[621]), .B(p_input[589]), .Z(n55436) );
  XNOR U55351 ( .A(n54586), .B(n55431), .Z(n55433) );
  XOR U55352 ( .A(n55437), .B(n55438), .Z(n54586) );
  AND U55353 ( .A(n1072), .B(n55439), .Z(n55438) );
  XOR U55354 ( .A(p_input[557]), .B(p_input[525]), .Z(n55439) );
  XOR U55355 ( .A(n55440), .B(n55441), .Z(n55431) );
  AND U55356 ( .A(n55442), .B(n55443), .Z(n55441) );
  XOR U55357 ( .A(n55440), .B(n54601), .Z(n55443) );
  XNOR U55358 ( .A(p_input[588]), .B(n55444), .Z(n54601) );
  AND U55359 ( .A(n1075), .B(n55445), .Z(n55444) );
  XOR U55360 ( .A(p_input[620]), .B(p_input[588]), .Z(n55445) );
  XNOR U55361 ( .A(n54598), .B(n55440), .Z(n55442) );
  XOR U55362 ( .A(n55446), .B(n55447), .Z(n54598) );
  AND U55363 ( .A(n1072), .B(n55448), .Z(n55447) );
  XOR U55364 ( .A(p_input[556]), .B(p_input[524]), .Z(n55448) );
  XOR U55365 ( .A(n55449), .B(n55450), .Z(n55440) );
  AND U55366 ( .A(n55451), .B(n55452), .Z(n55450) );
  XOR U55367 ( .A(n55449), .B(n54613), .Z(n55452) );
  XNOR U55368 ( .A(p_input[587]), .B(n55453), .Z(n54613) );
  AND U55369 ( .A(n1075), .B(n55454), .Z(n55453) );
  XOR U55370 ( .A(p_input[619]), .B(p_input[587]), .Z(n55454) );
  XNOR U55371 ( .A(n54610), .B(n55449), .Z(n55451) );
  XOR U55372 ( .A(n55455), .B(n55456), .Z(n54610) );
  AND U55373 ( .A(n1072), .B(n55457), .Z(n55456) );
  XOR U55374 ( .A(p_input[555]), .B(p_input[523]), .Z(n55457) );
  XOR U55375 ( .A(n55458), .B(n55459), .Z(n55449) );
  AND U55376 ( .A(n55460), .B(n55461), .Z(n55459) );
  XOR U55377 ( .A(n55458), .B(n54625), .Z(n55461) );
  XNOR U55378 ( .A(p_input[586]), .B(n55462), .Z(n54625) );
  AND U55379 ( .A(n1075), .B(n55463), .Z(n55462) );
  XOR U55380 ( .A(p_input[618]), .B(p_input[586]), .Z(n55463) );
  XNOR U55381 ( .A(n54622), .B(n55458), .Z(n55460) );
  XOR U55382 ( .A(n55464), .B(n55465), .Z(n54622) );
  AND U55383 ( .A(n1072), .B(n55466), .Z(n55465) );
  XOR U55384 ( .A(p_input[554]), .B(p_input[522]), .Z(n55466) );
  XOR U55385 ( .A(n55467), .B(n55468), .Z(n55458) );
  AND U55386 ( .A(n55469), .B(n55470), .Z(n55468) );
  XOR U55387 ( .A(n55467), .B(n54637), .Z(n55470) );
  XNOR U55388 ( .A(p_input[585]), .B(n55471), .Z(n54637) );
  AND U55389 ( .A(n1075), .B(n55472), .Z(n55471) );
  XOR U55390 ( .A(p_input[617]), .B(p_input[585]), .Z(n55472) );
  XNOR U55391 ( .A(n54634), .B(n55467), .Z(n55469) );
  XOR U55392 ( .A(n55473), .B(n55474), .Z(n54634) );
  AND U55393 ( .A(n1072), .B(n55475), .Z(n55474) );
  XOR U55394 ( .A(p_input[553]), .B(p_input[521]), .Z(n55475) );
  XOR U55395 ( .A(n55476), .B(n55477), .Z(n55467) );
  AND U55396 ( .A(n55478), .B(n55479), .Z(n55477) );
  XOR U55397 ( .A(n55476), .B(n54649), .Z(n55479) );
  XNOR U55398 ( .A(p_input[584]), .B(n55480), .Z(n54649) );
  AND U55399 ( .A(n1075), .B(n55481), .Z(n55480) );
  XOR U55400 ( .A(p_input[616]), .B(p_input[584]), .Z(n55481) );
  XNOR U55401 ( .A(n54646), .B(n55476), .Z(n55478) );
  XOR U55402 ( .A(n55482), .B(n55483), .Z(n54646) );
  AND U55403 ( .A(n1072), .B(n55484), .Z(n55483) );
  XOR U55404 ( .A(p_input[552]), .B(p_input[520]), .Z(n55484) );
  XOR U55405 ( .A(n55485), .B(n55486), .Z(n55476) );
  AND U55406 ( .A(n55487), .B(n55488), .Z(n55486) );
  XOR U55407 ( .A(n55485), .B(n54661), .Z(n55488) );
  XNOR U55408 ( .A(p_input[583]), .B(n55489), .Z(n54661) );
  AND U55409 ( .A(n1075), .B(n55490), .Z(n55489) );
  XOR U55410 ( .A(p_input[615]), .B(p_input[583]), .Z(n55490) );
  XNOR U55411 ( .A(n54658), .B(n55485), .Z(n55487) );
  XOR U55412 ( .A(n55491), .B(n55492), .Z(n54658) );
  AND U55413 ( .A(n1072), .B(n55493), .Z(n55492) );
  XOR U55414 ( .A(p_input[551]), .B(p_input[519]), .Z(n55493) );
  XOR U55415 ( .A(n55494), .B(n55495), .Z(n55485) );
  AND U55416 ( .A(n55496), .B(n55497), .Z(n55495) );
  XOR U55417 ( .A(n55494), .B(n54673), .Z(n55497) );
  XNOR U55418 ( .A(p_input[582]), .B(n55498), .Z(n54673) );
  AND U55419 ( .A(n1075), .B(n55499), .Z(n55498) );
  XOR U55420 ( .A(p_input[614]), .B(p_input[582]), .Z(n55499) );
  XNOR U55421 ( .A(n54670), .B(n55494), .Z(n55496) );
  XOR U55422 ( .A(n55500), .B(n55501), .Z(n54670) );
  AND U55423 ( .A(n1072), .B(n55502), .Z(n55501) );
  XOR U55424 ( .A(p_input[550]), .B(p_input[518]), .Z(n55502) );
  XOR U55425 ( .A(n55503), .B(n55504), .Z(n55494) );
  AND U55426 ( .A(n55505), .B(n55506), .Z(n55504) );
  XOR U55427 ( .A(n55503), .B(n54685), .Z(n55506) );
  XNOR U55428 ( .A(p_input[581]), .B(n55507), .Z(n54685) );
  AND U55429 ( .A(n1075), .B(n55508), .Z(n55507) );
  XOR U55430 ( .A(p_input[613]), .B(p_input[581]), .Z(n55508) );
  XNOR U55431 ( .A(n54682), .B(n55503), .Z(n55505) );
  XOR U55432 ( .A(n55509), .B(n55510), .Z(n54682) );
  AND U55433 ( .A(n1072), .B(n55511), .Z(n55510) );
  XOR U55434 ( .A(p_input[549]), .B(p_input[517]), .Z(n55511) );
  XOR U55435 ( .A(n55512), .B(n55513), .Z(n55503) );
  AND U55436 ( .A(n55514), .B(n55515), .Z(n55513) );
  XOR U55437 ( .A(n55512), .B(n54697), .Z(n55515) );
  XNOR U55438 ( .A(p_input[580]), .B(n55516), .Z(n54697) );
  AND U55439 ( .A(n1075), .B(n55517), .Z(n55516) );
  XOR U55440 ( .A(p_input[612]), .B(p_input[580]), .Z(n55517) );
  XNOR U55441 ( .A(n54694), .B(n55512), .Z(n55514) );
  XOR U55442 ( .A(n55518), .B(n55519), .Z(n54694) );
  AND U55443 ( .A(n1072), .B(n55520), .Z(n55519) );
  XOR U55444 ( .A(p_input[548]), .B(p_input[516]), .Z(n55520) );
  XOR U55445 ( .A(n55521), .B(n55522), .Z(n55512) );
  AND U55446 ( .A(n55523), .B(n55524), .Z(n55522) );
  XOR U55447 ( .A(n55521), .B(n54709), .Z(n55524) );
  XNOR U55448 ( .A(p_input[579]), .B(n55525), .Z(n54709) );
  AND U55449 ( .A(n1075), .B(n55526), .Z(n55525) );
  XOR U55450 ( .A(p_input[611]), .B(p_input[579]), .Z(n55526) );
  XNOR U55451 ( .A(n54706), .B(n55521), .Z(n55523) );
  XOR U55452 ( .A(n55527), .B(n55528), .Z(n54706) );
  AND U55453 ( .A(n1072), .B(n55529), .Z(n55528) );
  XOR U55454 ( .A(p_input[547]), .B(p_input[515]), .Z(n55529) );
  XOR U55455 ( .A(n55530), .B(n55531), .Z(n55521) );
  AND U55456 ( .A(n55532), .B(n55533), .Z(n55531) );
  XOR U55457 ( .A(n55530), .B(n54721), .Z(n55533) );
  XNOR U55458 ( .A(p_input[578]), .B(n55534), .Z(n54721) );
  AND U55459 ( .A(n1075), .B(n55535), .Z(n55534) );
  XOR U55460 ( .A(p_input[610]), .B(p_input[578]), .Z(n55535) );
  XNOR U55461 ( .A(n54718), .B(n55530), .Z(n55532) );
  XOR U55462 ( .A(n55536), .B(n55537), .Z(n54718) );
  AND U55463 ( .A(n1072), .B(n55538), .Z(n55537) );
  XOR U55464 ( .A(p_input[546]), .B(p_input[514]), .Z(n55538) );
  XOR U55465 ( .A(n55539), .B(n55540), .Z(n55530) );
  AND U55466 ( .A(n55541), .B(n55542), .Z(n55540) );
  XNOR U55467 ( .A(n55543), .B(n54734), .Z(n55542) );
  XNOR U55468 ( .A(p_input[577]), .B(n55544), .Z(n54734) );
  AND U55469 ( .A(n1075), .B(n55545), .Z(n55544) );
  XNOR U55470 ( .A(p_input[609]), .B(n55546), .Z(n55545) );
  IV U55471 ( .A(p_input[577]), .Z(n55546) );
  XNOR U55472 ( .A(n54731), .B(n55539), .Z(n55541) );
  XNOR U55473 ( .A(p_input[513]), .B(n55547), .Z(n54731) );
  AND U55474 ( .A(n1072), .B(n55548), .Z(n55547) );
  XOR U55475 ( .A(p_input[545]), .B(p_input[513]), .Z(n55548) );
  IV U55476 ( .A(n55543), .Z(n55539) );
  AND U55477 ( .A(n55269), .B(n55272), .Z(n55543) );
  XOR U55478 ( .A(p_input[576]), .B(n55549), .Z(n55272) );
  AND U55479 ( .A(n1075), .B(n55550), .Z(n55549) );
  XOR U55480 ( .A(p_input[608]), .B(p_input[576]), .Z(n55550) );
  XOR U55481 ( .A(n55551), .B(n55552), .Z(n1075) );
  AND U55482 ( .A(n55553), .B(n55554), .Z(n55552) );
  XNOR U55483 ( .A(p_input[639]), .B(n55551), .Z(n55554) );
  XOR U55484 ( .A(n55551), .B(p_input[607]), .Z(n55553) );
  XOR U55485 ( .A(n55555), .B(n55556), .Z(n55551) );
  AND U55486 ( .A(n55557), .B(n55558), .Z(n55556) );
  XNOR U55487 ( .A(p_input[638]), .B(n55555), .Z(n55558) );
  XOR U55488 ( .A(n55555), .B(p_input[606]), .Z(n55557) );
  XOR U55489 ( .A(n55559), .B(n55560), .Z(n55555) );
  AND U55490 ( .A(n55561), .B(n55562), .Z(n55560) );
  XNOR U55491 ( .A(p_input[637]), .B(n55559), .Z(n55562) );
  XOR U55492 ( .A(n55559), .B(p_input[605]), .Z(n55561) );
  XOR U55493 ( .A(n55563), .B(n55564), .Z(n55559) );
  AND U55494 ( .A(n55565), .B(n55566), .Z(n55564) );
  XNOR U55495 ( .A(p_input[636]), .B(n55563), .Z(n55566) );
  XOR U55496 ( .A(n55563), .B(p_input[604]), .Z(n55565) );
  XOR U55497 ( .A(n55567), .B(n55568), .Z(n55563) );
  AND U55498 ( .A(n55569), .B(n55570), .Z(n55568) );
  XNOR U55499 ( .A(p_input[635]), .B(n55567), .Z(n55570) );
  XOR U55500 ( .A(n55567), .B(p_input[603]), .Z(n55569) );
  XOR U55501 ( .A(n55571), .B(n55572), .Z(n55567) );
  AND U55502 ( .A(n55573), .B(n55574), .Z(n55572) );
  XNOR U55503 ( .A(p_input[634]), .B(n55571), .Z(n55574) );
  XOR U55504 ( .A(n55571), .B(p_input[602]), .Z(n55573) );
  XOR U55505 ( .A(n55575), .B(n55576), .Z(n55571) );
  AND U55506 ( .A(n55577), .B(n55578), .Z(n55576) );
  XNOR U55507 ( .A(p_input[633]), .B(n55575), .Z(n55578) );
  XOR U55508 ( .A(n55575), .B(p_input[601]), .Z(n55577) );
  XOR U55509 ( .A(n55579), .B(n55580), .Z(n55575) );
  AND U55510 ( .A(n55581), .B(n55582), .Z(n55580) );
  XNOR U55511 ( .A(p_input[632]), .B(n55579), .Z(n55582) );
  XOR U55512 ( .A(n55579), .B(p_input[600]), .Z(n55581) );
  XOR U55513 ( .A(n55583), .B(n55584), .Z(n55579) );
  AND U55514 ( .A(n55585), .B(n55586), .Z(n55584) );
  XNOR U55515 ( .A(p_input[631]), .B(n55583), .Z(n55586) );
  XOR U55516 ( .A(n55583), .B(p_input[599]), .Z(n55585) );
  XOR U55517 ( .A(n55587), .B(n55588), .Z(n55583) );
  AND U55518 ( .A(n55589), .B(n55590), .Z(n55588) );
  XNOR U55519 ( .A(p_input[630]), .B(n55587), .Z(n55590) );
  XOR U55520 ( .A(n55587), .B(p_input[598]), .Z(n55589) );
  XOR U55521 ( .A(n55591), .B(n55592), .Z(n55587) );
  AND U55522 ( .A(n55593), .B(n55594), .Z(n55592) );
  XNOR U55523 ( .A(p_input[629]), .B(n55591), .Z(n55594) );
  XOR U55524 ( .A(n55591), .B(p_input[597]), .Z(n55593) );
  XOR U55525 ( .A(n55595), .B(n55596), .Z(n55591) );
  AND U55526 ( .A(n55597), .B(n55598), .Z(n55596) );
  XNOR U55527 ( .A(p_input[628]), .B(n55595), .Z(n55598) );
  XOR U55528 ( .A(n55595), .B(p_input[596]), .Z(n55597) );
  XOR U55529 ( .A(n55599), .B(n55600), .Z(n55595) );
  AND U55530 ( .A(n55601), .B(n55602), .Z(n55600) );
  XNOR U55531 ( .A(p_input[627]), .B(n55599), .Z(n55602) );
  XOR U55532 ( .A(n55599), .B(p_input[595]), .Z(n55601) );
  XOR U55533 ( .A(n55603), .B(n55604), .Z(n55599) );
  AND U55534 ( .A(n55605), .B(n55606), .Z(n55604) );
  XNOR U55535 ( .A(p_input[626]), .B(n55603), .Z(n55606) );
  XOR U55536 ( .A(n55603), .B(p_input[594]), .Z(n55605) );
  XOR U55537 ( .A(n55607), .B(n55608), .Z(n55603) );
  AND U55538 ( .A(n55609), .B(n55610), .Z(n55608) );
  XNOR U55539 ( .A(p_input[625]), .B(n55607), .Z(n55610) );
  XOR U55540 ( .A(n55607), .B(p_input[593]), .Z(n55609) );
  XOR U55541 ( .A(n55611), .B(n55612), .Z(n55607) );
  AND U55542 ( .A(n55613), .B(n55614), .Z(n55612) );
  XNOR U55543 ( .A(p_input[624]), .B(n55611), .Z(n55614) );
  XOR U55544 ( .A(n55611), .B(p_input[592]), .Z(n55613) );
  XOR U55545 ( .A(n55615), .B(n55616), .Z(n55611) );
  AND U55546 ( .A(n55617), .B(n55618), .Z(n55616) );
  XNOR U55547 ( .A(p_input[623]), .B(n55615), .Z(n55618) );
  XOR U55548 ( .A(n55615), .B(p_input[591]), .Z(n55617) );
  XOR U55549 ( .A(n55619), .B(n55620), .Z(n55615) );
  AND U55550 ( .A(n55621), .B(n55622), .Z(n55620) );
  XNOR U55551 ( .A(p_input[622]), .B(n55619), .Z(n55622) );
  XOR U55552 ( .A(n55619), .B(p_input[590]), .Z(n55621) );
  XOR U55553 ( .A(n55623), .B(n55624), .Z(n55619) );
  AND U55554 ( .A(n55625), .B(n55626), .Z(n55624) );
  XNOR U55555 ( .A(p_input[621]), .B(n55623), .Z(n55626) );
  XOR U55556 ( .A(n55623), .B(p_input[589]), .Z(n55625) );
  XOR U55557 ( .A(n55627), .B(n55628), .Z(n55623) );
  AND U55558 ( .A(n55629), .B(n55630), .Z(n55628) );
  XNOR U55559 ( .A(p_input[620]), .B(n55627), .Z(n55630) );
  XOR U55560 ( .A(n55627), .B(p_input[588]), .Z(n55629) );
  XOR U55561 ( .A(n55631), .B(n55632), .Z(n55627) );
  AND U55562 ( .A(n55633), .B(n55634), .Z(n55632) );
  XNOR U55563 ( .A(p_input[619]), .B(n55631), .Z(n55634) );
  XOR U55564 ( .A(n55631), .B(p_input[587]), .Z(n55633) );
  XOR U55565 ( .A(n55635), .B(n55636), .Z(n55631) );
  AND U55566 ( .A(n55637), .B(n55638), .Z(n55636) );
  XNOR U55567 ( .A(p_input[618]), .B(n55635), .Z(n55638) );
  XOR U55568 ( .A(n55635), .B(p_input[586]), .Z(n55637) );
  XOR U55569 ( .A(n55639), .B(n55640), .Z(n55635) );
  AND U55570 ( .A(n55641), .B(n55642), .Z(n55640) );
  XNOR U55571 ( .A(p_input[617]), .B(n55639), .Z(n55642) );
  XOR U55572 ( .A(n55639), .B(p_input[585]), .Z(n55641) );
  XOR U55573 ( .A(n55643), .B(n55644), .Z(n55639) );
  AND U55574 ( .A(n55645), .B(n55646), .Z(n55644) );
  XNOR U55575 ( .A(p_input[616]), .B(n55643), .Z(n55646) );
  XOR U55576 ( .A(n55643), .B(p_input[584]), .Z(n55645) );
  XOR U55577 ( .A(n55647), .B(n55648), .Z(n55643) );
  AND U55578 ( .A(n55649), .B(n55650), .Z(n55648) );
  XNOR U55579 ( .A(p_input[615]), .B(n55647), .Z(n55650) );
  XOR U55580 ( .A(n55647), .B(p_input[583]), .Z(n55649) );
  XOR U55581 ( .A(n55651), .B(n55652), .Z(n55647) );
  AND U55582 ( .A(n55653), .B(n55654), .Z(n55652) );
  XNOR U55583 ( .A(p_input[614]), .B(n55651), .Z(n55654) );
  XOR U55584 ( .A(n55651), .B(p_input[582]), .Z(n55653) );
  XOR U55585 ( .A(n55655), .B(n55656), .Z(n55651) );
  AND U55586 ( .A(n55657), .B(n55658), .Z(n55656) );
  XNOR U55587 ( .A(p_input[613]), .B(n55655), .Z(n55658) );
  XOR U55588 ( .A(n55655), .B(p_input[581]), .Z(n55657) );
  XOR U55589 ( .A(n55659), .B(n55660), .Z(n55655) );
  AND U55590 ( .A(n55661), .B(n55662), .Z(n55660) );
  XNOR U55591 ( .A(p_input[612]), .B(n55659), .Z(n55662) );
  XOR U55592 ( .A(n55659), .B(p_input[580]), .Z(n55661) );
  XOR U55593 ( .A(n55663), .B(n55664), .Z(n55659) );
  AND U55594 ( .A(n55665), .B(n55666), .Z(n55664) );
  XNOR U55595 ( .A(p_input[611]), .B(n55663), .Z(n55666) );
  XOR U55596 ( .A(n55663), .B(p_input[579]), .Z(n55665) );
  XOR U55597 ( .A(n55667), .B(n55668), .Z(n55663) );
  AND U55598 ( .A(n55669), .B(n55670), .Z(n55668) );
  XNOR U55599 ( .A(p_input[610]), .B(n55667), .Z(n55670) );
  XOR U55600 ( .A(n55667), .B(p_input[578]), .Z(n55669) );
  XNOR U55601 ( .A(n55671), .B(n55672), .Z(n55667) );
  AND U55602 ( .A(n55673), .B(n55674), .Z(n55672) );
  XOR U55603 ( .A(p_input[609]), .B(n55671), .Z(n55674) );
  XNOR U55604 ( .A(p_input[577]), .B(n55671), .Z(n55673) );
  AND U55605 ( .A(p_input[608]), .B(n55675), .Z(n55671) );
  IV U55606 ( .A(p_input[576]), .Z(n55675) );
  XNOR U55607 ( .A(p_input[512]), .B(n55676), .Z(n55269) );
  AND U55608 ( .A(n1072), .B(n55677), .Z(n55676) );
  XOR U55609 ( .A(p_input[544]), .B(p_input[512]), .Z(n55677) );
  XOR U55610 ( .A(n55678), .B(n55679), .Z(n1072) );
  AND U55611 ( .A(n55680), .B(n55681), .Z(n55679) );
  XNOR U55612 ( .A(p_input[575]), .B(n55678), .Z(n55681) );
  XOR U55613 ( .A(n55678), .B(p_input[543]), .Z(n55680) );
  XOR U55614 ( .A(n55682), .B(n55683), .Z(n55678) );
  AND U55615 ( .A(n55684), .B(n55685), .Z(n55683) );
  XNOR U55616 ( .A(p_input[574]), .B(n55682), .Z(n55685) );
  XNOR U55617 ( .A(n55682), .B(n55284), .Z(n55684) );
  IV U55618 ( .A(p_input[542]), .Z(n55284) );
  XOR U55619 ( .A(n55686), .B(n55687), .Z(n55682) );
  AND U55620 ( .A(n55688), .B(n55689), .Z(n55687) );
  XNOR U55621 ( .A(p_input[573]), .B(n55686), .Z(n55689) );
  XNOR U55622 ( .A(n55686), .B(n55293), .Z(n55688) );
  IV U55623 ( .A(p_input[541]), .Z(n55293) );
  XOR U55624 ( .A(n55690), .B(n55691), .Z(n55686) );
  AND U55625 ( .A(n55692), .B(n55693), .Z(n55691) );
  XNOR U55626 ( .A(p_input[572]), .B(n55690), .Z(n55693) );
  XNOR U55627 ( .A(n55690), .B(n55302), .Z(n55692) );
  IV U55628 ( .A(p_input[540]), .Z(n55302) );
  XOR U55629 ( .A(n55694), .B(n55695), .Z(n55690) );
  AND U55630 ( .A(n55696), .B(n55697), .Z(n55695) );
  XNOR U55631 ( .A(p_input[571]), .B(n55694), .Z(n55697) );
  XNOR U55632 ( .A(n55694), .B(n55311), .Z(n55696) );
  IV U55633 ( .A(p_input[539]), .Z(n55311) );
  XOR U55634 ( .A(n55698), .B(n55699), .Z(n55694) );
  AND U55635 ( .A(n55700), .B(n55701), .Z(n55699) );
  XNOR U55636 ( .A(p_input[570]), .B(n55698), .Z(n55701) );
  XNOR U55637 ( .A(n55698), .B(n55320), .Z(n55700) );
  IV U55638 ( .A(p_input[538]), .Z(n55320) );
  XOR U55639 ( .A(n55702), .B(n55703), .Z(n55698) );
  AND U55640 ( .A(n55704), .B(n55705), .Z(n55703) );
  XNOR U55641 ( .A(p_input[569]), .B(n55702), .Z(n55705) );
  XNOR U55642 ( .A(n55702), .B(n55329), .Z(n55704) );
  IV U55643 ( .A(p_input[537]), .Z(n55329) );
  XOR U55644 ( .A(n55706), .B(n55707), .Z(n55702) );
  AND U55645 ( .A(n55708), .B(n55709), .Z(n55707) );
  XNOR U55646 ( .A(p_input[568]), .B(n55706), .Z(n55709) );
  XNOR U55647 ( .A(n55706), .B(n55338), .Z(n55708) );
  IV U55648 ( .A(p_input[536]), .Z(n55338) );
  XOR U55649 ( .A(n55710), .B(n55711), .Z(n55706) );
  AND U55650 ( .A(n55712), .B(n55713), .Z(n55711) );
  XNOR U55651 ( .A(p_input[567]), .B(n55710), .Z(n55713) );
  XNOR U55652 ( .A(n55710), .B(n55347), .Z(n55712) );
  IV U55653 ( .A(p_input[535]), .Z(n55347) );
  XOR U55654 ( .A(n55714), .B(n55715), .Z(n55710) );
  AND U55655 ( .A(n55716), .B(n55717), .Z(n55715) );
  XNOR U55656 ( .A(p_input[566]), .B(n55714), .Z(n55717) );
  XNOR U55657 ( .A(n55714), .B(n55356), .Z(n55716) );
  IV U55658 ( .A(p_input[534]), .Z(n55356) );
  XOR U55659 ( .A(n55718), .B(n55719), .Z(n55714) );
  AND U55660 ( .A(n55720), .B(n55721), .Z(n55719) );
  XNOR U55661 ( .A(p_input[565]), .B(n55718), .Z(n55721) );
  XNOR U55662 ( .A(n55718), .B(n55365), .Z(n55720) );
  IV U55663 ( .A(p_input[533]), .Z(n55365) );
  XOR U55664 ( .A(n55722), .B(n55723), .Z(n55718) );
  AND U55665 ( .A(n55724), .B(n55725), .Z(n55723) );
  XNOR U55666 ( .A(p_input[564]), .B(n55722), .Z(n55725) );
  XNOR U55667 ( .A(n55722), .B(n55374), .Z(n55724) );
  IV U55668 ( .A(p_input[532]), .Z(n55374) );
  XOR U55669 ( .A(n55726), .B(n55727), .Z(n55722) );
  AND U55670 ( .A(n55728), .B(n55729), .Z(n55727) );
  XNOR U55671 ( .A(p_input[563]), .B(n55726), .Z(n55729) );
  XNOR U55672 ( .A(n55726), .B(n55383), .Z(n55728) );
  IV U55673 ( .A(p_input[531]), .Z(n55383) );
  XOR U55674 ( .A(n55730), .B(n55731), .Z(n55726) );
  AND U55675 ( .A(n55732), .B(n55733), .Z(n55731) );
  XNOR U55676 ( .A(p_input[562]), .B(n55730), .Z(n55733) );
  XNOR U55677 ( .A(n55730), .B(n55392), .Z(n55732) );
  IV U55678 ( .A(p_input[530]), .Z(n55392) );
  XOR U55679 ( .A(n55734), .B(n55735), .Z(n55730) );
  AND U55680 ( .A(n55736), .B(n55737), .Z(n55735) );
  XNOR U55681 ( .A(p_input[561]), .B(n55734), .Z(n55737) );
  XNOR U55682 ( .A(n55734), .B(n55401), .Z(n55736) );
  IV U55683 ( .A(p_input[529]), .Z(n55401) );
  XOR U55684 ( .A(n55738), .B(n55739), .Z(n55734) );
  AND U55685 ( .A(n55740), .B(n55741), .Z(n55739) );
  XNOR U55686 ( .A(p_input[560]), .B(n55738), .Z(n55741) );
  XNOR U55687 ( .A(n55738), .B(n55410), .Z(n55740) );
  IV U55688 ( .A(p_input[528]), .Z(n55410) );
  XOR U55689 ( .A(n55742), .B(n55743), .Z(n55738) );
  AND U55690 ( .A(n55744), .B(n55745), .Z(n55743) );
  XNOR U55691 ( .A(p_input[559]), .B(n55742), .Z(n55745) );
  XNOR U55692 ( .A(n55742), .B(n55419), .Z(n55744) );
  IV U55693 ( .A(p_input[527]), .Z(n55419) );
  XOR U55694 ( .A(n55746), .B(n55747), .Z(n55742) );
  AND U55695 ( .A(n55748), .B(n55749), .Z(n55747) );
  XNOR U55696 ( .A(p_input[558]), .B(n55746), .Z(n55749) );
  XNOR U55697 ( .A(n55746), .B(n55428), .Z(n55748) );
  IV U55698 ( .A(p_input[526]), .Z(n55428) );
  XOR U55699 ( .A(n55750), .B(n55751), .Z(n55746) );
  AND U55700 ( .A(n55752), .B(n55753), .Z(n55751) );
  XNOR U55701 ( .A(p_input[557]), .B(n55750), .Z(n55753) );
  XNOR U55702 ( .A(n55750), .B(n55437), .Z(n55752) );
  IV U55703 ( .A(p_input[525]), .Z(n55437) );
  XOR U55704 ( .A(n55754), .B(n55755), .Z(n55750) );
  AND U55705 ( .A(n55756), .B(n55757), .Z(n55755) );
  XNOR U55706 ( .A(p_input[556]), .B(n55754), .Z(n55757) );
  XNOR U55707 ( .A(n55754), .B(n55446), .Z(n55756) );
  IV U55708 ( .A(p_input[524]), .Z(n55446) );
  XOR U55709 ( .A(n55758), .B(n55759), .Z(n55754) );
  AND U55710 ( .A(n55760), .B(n55761), .Z(n55759) );
  XNOR U55711 ( .A(p_input[555]), .B(n55758), .Z(n55761) );
  XNOR U55712 ( .A(n55758), .B(n55455), .Z(n55760) );
  IV U55713 ( .A(p_input[523]), .Z(n55455) );
  XOR U55714 ( .A(n55762), .B(n55763), .Z(n55758) );
  AND U55715 ( .A(n55764), .B(n55765), .Z(n55763) );
  XNOR U55716 ( .A(p_input[554]), .B(n55762), .Z(n55765) );
  XNOR U55717 ( .A(n55762), .B(n55464), .Z(n55764) );
  IV U55718 ( .A(p_input[522]), .Z(n55464) );
  XOR U55719 ( .A(n55766), .B(n55767), .Z(n55762) );
  AND U55720 ( .A(n55768), .B(n55769), .Z(n55767) );
  XNOR U55721 ( .A(p_input[553]), .B(n55766), .Z(n55769) );
  XNOR U55722 ( .A(n55766), .B(n55473), .Z(n55768) );
  IV U55723 ( .A(p_input[521]), .Z(n55473) );
  XOR U55724 ( .A(n55770), .B(n55771), .Z(n55766) );
  AND U55725 ( .A(n55772), .B(n55773), .Z(n55771) );
  XNOR U55726 ( .A(p_input[552]), .B(n55770), .Z(n55773) );
  XNOR U55727 ( .A(n55770), .B(n55482), .Z(n55772) );
  IV U55728 ( .A(p_input[520]), .Z(n55482) );
  XOR U55729 ( .A(n55774), .B(n55775), .Z(n55770) );
  AND U55730 ( .A(n55776), .B(n55777), .Z(n55775) );
  XNOR U55731 ( .A(p_input[551]), .B(n55774), .Z(n55777) );
  XNOR U55732 ( .A(n55774), .B(n55491), .Z(n55776) );
  IV U55733 ( .A(p_input[519]), .Z(n55491) );
  XOR U55734 ( .A(n55778), .B(n55779), .Z(n55774) );
  AND U55735 ( .A(n55780), .B(n55781), .Z(n55779) );
  XNOR U55736 ( .A(p_input[550]), .B(n55778), .Z(n55781) );
  XNOR U55737 ( .A(n55778), .B(n55500), .Z(n55780) );
  IV U55738 ( .A(p_input[518]), .Z(n55500) );
  XOR U55739 ( .A(n55782), .B(n55783), .Z(n55778) );
  AND U55740 ( .A(n55784), .B(n55785), .Z(n55783) );
  XNOR U55741 ( .A(p_input[549]), .B(n55782), .Z(n55785) );
  XNOR U55742 ( .A(n55782), .B(n55509), .Z(n55784) );
  IV U55743 ( .A(p_input[517]), .Z(n55509) );
  XOR U55744 ( .A(n55786), .B(n55787), .Z(n55782) );
  AND U55745 ( .A(n55788), .B(n55789), .Z(n55787) );
  XNOR U55746 ( .A(p_input[548]), .B(n55786), .Z(n55789) );
  XNOR U55747 ( .A(n55786), .B(n55518), .Z(n55788) );
  IV U55748 ( .A(p_input[516]), .Z(n55518) );
  XOR U55749 ( .A(n55790), .B(n55791), .Z(n55786) );
  AND U55750 ( .A(n55792), .B(n55793), .Z(n55791) );
  XNOR U55751 ( .A(p_input[547]), .B(n55790), .Z(n55793) );
  XNOR U55752 ( .A(n55790), .B(n55527), .Z(n55792) );
  IV U55753 ( .A(p_input[515]), .Z(n55527) );
  XOR U55754 ( .A(n55794), .B(n55795), .Z(n55790) );
  AND U55755 ( .A(n55796), .B(n55797), .Z(n55795) );
  XNOR U55756 ( .A(p_input[546]), .B(n55794), .Z(n55797) );
  XNOR U55757 ( .A(n55794), .B(n55536), .Z(n55796) );
  IV U55758 ( .A(p_input[514]), .Z(n55536) );
  XNOR U55759 ( .A(n55798), .B(n55799), .Z(n55794) );
  AND U55760 ( .A(n55800), .B(n55801), .Z(n55799) );
  XOR U55761 ( .A(p_input[545]), .B(n55798), .Z(n55801) );
  XNOR U55762 ( .A(p_input[513]), .B(n55798), .Z(n55800) );
  AND U55763 ( .A(p_input[544]), .B(n55802), .Z(n55798) );
  IV U55764 ( .A(p_input[512]), .Z(n55802) );
  XOR U55765 ( .A(n55803), .B(n55804), .Z(n52159) );
  AND U55766 ( .A(n1040), .B(n55805), .Z(n55804) );
  XNOR U55767 ( .A(n55806), .B(n55803), .Z(n55805) );
  XOR U55768 ( .A(n55807), .B(n55808), .Z(n1040) );
  AND U55769 ( .A(n55809), .B(n55810), .Z(n55808) );
  XOR U55770 ( .A(n55807), .B(n52174), .Z(n55810) );
  XOR U55771 ( .A(n55811), .B(n55812), .Z(n52174) );
  AND U55772 ( .A(n919), .B(n55813), .Z(n55812) );
  XOR U55773 ( .A(n55814), .B(n55811), .Z(n55813) );
  XNOR U55774 ( .A(n52171), .B(n55807), .Z(n55809) );
  XOR U55775 ( .A(n55815), .B(n55816), .Z(n52171) );
  AND U55776 ( .A(n916), .B(n55817), .Z(n55816) );
  XOR U55777 ( .A(n55818), .B(n55815), .Z(n55817) );
  XOR U55778 ( .A(n55819), .B(n55820), .Z(n55807) );
  AND U55779 ( .A(n55821), .B(n55822), .Z(n55820) );
  XOR U55780 ( .A(n55819), .B(n52186), .Z(n55822) );
  XOR U55781 ( .A(n55823), .B(n55824), .Z(n52186) );
  AND U55782 ( .A(n919), .B(n55825), .Z(n55824) );
  XOR U55783 ( .A(n55826), .B(n55823), .Z(n55825) );
  XNOR U55784 ( .A(n52183), .B(n55819), .Z(n55821) );
  XOR U55785 ( .A(n55827), .B(n55828), .Z(n52183) );
  AND U55786 ( .A(n916), .B(n55829), .Z(n55828) );
  XOR U55787 ( .A(n55830), .B(n55827), .Z(n55829) );
  XOR U55788 ( .A(n55831), .B(n55832), .Z(n55819) );
  AND U55789 ( .A(n55833), .B(n55834), .Z(n55832) );
  XOR U55790 ( .A(n55831), .B(n52198), .Z(n55834) );
  XOR U55791 ( .A(n55835), .B(n55836), .Z(n52198) );
  AND U55792 ( .A(n919), .B(n55837), .Z(n55836) );
  XOR U55793 ( .A(n55838), .B(n55835), .Z(n55837) );
  XNOR U55794 ( .A(n52195), .B(n55831), .Z(n55833) );
  XOR U55795 ( .A(n55839), .B(n55840), .Z(n52195) );
  AND U55796 ( .A(n916), .B(n55841), .Z(n55840) );
  XOR U55797 ( .A(n55842), .B(n55839), .Z(n55841) );
  XOR U55798 ( .A(n55843), .B(n55844), .Z(n55831) );
  AND U55799 ( .A(n55845), .B(n55846), .Z(n55844) );
  XOR U55800 ( .A(n55843), .B(n52210), .Z(n55846) );
  XOR U55801 ( .A(n55847), .B(n55848), .Z(n52210) );
  AND U55802 ( .A(n919), .B(n55849), .Z(n55848) );
  XOR U55803 ( .A(n55850), .B(n55847), .Z(n55849) );
  XNOR U55804 ( .A(n52207), .B(n55843), .Z(n55845) );
  XOR U55805 ( .A(n55851), .B(n55852), .Z(n52207) );
  AND U55806 ( .A(n916), .B(n55853), .Z(n55852) );
  XOR U55807 ( .A(n55854), .B(n55851), .Z(n55853) );
  XOR U55808 ( .A(n55855), .B(n55856), .Z(n55843) );
  AND U55809 ( .A(n55857), .B(n55858), .Z(n55856) );
  XOR U55810 ( .A(n55855), .B(n52222), .Z(n55858) );
  XOR U55811 ( .A(n55859), .B(n55860), .Z(n52222) );
  AND U55812 ( .A(n919), .B(n55861), .Z(n55860) );
  XOR U55813 ( .A(n55862), .B(n55859), .Z(n55861) );
  XNOR U55814 ( .A(n52219), .B(n55855), .Z(n55857) );
  XOR U55815 ( .A(n55863), .B(n55864), .Z(n52219) );
  AND U55816 ( .A(n916), .B(n55865), .Z(n55864) );
  XOR U55817 ( .A(n55866), .B(n55863), .Z(n55865) );
  XOR U55818 ( .A(n55867), .B(n55868), .Z(n55855) );
  AND U55819 ( .A(n55869), .B(n55870), .Z(n55868) );
  XOR U55820 ( .A(n55867), .B(n52234), .Z(n55870) );
  XOR U55821 ( .A(n55871), .B(n55872), .Z(n52234) );
  AND U55822 ( .A(n919), .B(n55873), .Z(n55872) );
  XOR U55823 ( .A(n55874), .B(n55871), .Z(n55873) );
  XNOR U55824 ( .A(n52231), .B(n55867), .Z(n55869) );
  XOR U55825 ( .A(n55875), .B(n55876), .Z(n52231) );
  AND U55826 ( .A(n916), .B(n55877), .Z(n55876) );
  XOR U55827 ( .A(n55878), .B(n55875), .Z(n55877) );
  XOR U55828 ( .A(n55879), .B(n55880), .Z(n55867) );
  AND U55829 ( .A(n55881), .B(n55882), .Z(n55880) );
  XOR U55830 ( .A(n55879), .B(n52246), .Z(n55882) );
  XOR U55831 ( .A(n55883), .B(n55884), .Z(n52246) );
  AND U55832 ( .A(n919), .B(n55885), .Z(n55884) );
  XOR U55833 ( .A(n55886), .B(n55883), .Z(n55885) );
  XNOR U55834 ( .A(n52243), .B(n55879), .Z(n55881) );
  XOR U55835 ( .A(n55887), .B(n55888), .Z(n52243) );
  AND U55836 ( .A(n916), .B(n55889), .Z(n55888) );
  XOR U55837 ( .A(n55890), .B(n55887), .Z(n55889) );
  XOR U55838 ( .A(n55891), .B(n55892), .Z(n55879) );
  AND U55839 ( .A(n55893), .B(n55894), .Z(n55892) );
  XOR U55840 ( .A(n55891), .B(n52258), .Z(n55894) );
  XOR U55841 ( .A(n55895), .B(n55896), .Z(n52258) );
  AND U55842 ( .A(n919), .B(n55897), .Z(n55896) );
  XOR U55843 ( .A(n55898), .B(n55895), .Z(n55897) );
  XNOR U55844 ( .A(n52255), .B(n55891), .Z(n55893) );
  XOR U55845 ( .A(n55899), .B(n55900), .Z(n52255) );
  AND U55846 ( .A(n916), .B(n55901), .Z(n55900) );
  XOR U55847 ( .A(n55902), .B(n55899), .Z(n55901) );
  XOR U55848 ( .A(n55903), .B(n55904), .Z(n55891) );
  AND U55849 ( .A(n55905), .B(n55906), .Z(n55904) );
  XOR U55850 ( .A(n55903), .B(n52270), .Z(n55906) );
  XOR U55851 ( .A(n55907), .B(n55908), .Z(n52270) );
  AND U55852 ( .A(n919), .B(n55909), .Z(n55908) );
  XOR U55853 ( .A(n55910), .B(n55907), .Z(n55909) );
  XNOR U55854 ( .A(n52267), .B(n55903), .Z(n55905) );
  XOR U55855 ( .A(n55911), .B(n55912), .Z(n52267) );
  AND U55856 ( .A(n916), .B(n55913), .Z(n55912) );
  XOR U55857 ( .A(n55914), .B(n55911), .Z(n55913) );
  XOR U55858 ( .A(n55915), .B(n55916), .Z(n55903) );
  AND U55859 ( .A(n55917), .B(n55918), .Z(n55916) );
  XOR U55860 ( .A(n55915), .B(n52282), .Z(n55918) );
  XOR U55861 ( .A(n55919), .B(n55920), .Z(n52282) );
  AND U55862 ( .A(n919), .B(n55921), .Z(n55920) );
  XOR U55863 ( .A(n55922), .B(n55919), .Z(n55921) );
  XNOR U55864 ( .A(n52279), .B(n55915), .Z(n55917) );
  XOR U55865 ( .A(n55923), .B(n55924), .Z(n52279) );
  AND U55866 ( .A(n916), .B(n55925), .Z(n55924) );
  XOR U55867 ( .A(n55926), .B(n55923), .Z(n55925) );
  XOR U55868 ( .A(n55927), .B(n55928), .Z(n55915) );
  AND U55869 ( .A(n55929), .B(n55930), .Z(n55928) );
  XOR U55870 ( .A(n55927), .B(n52294), .Z(n55930) );
  XOR U55871 ( .A(n55931), .B(n55932), .Z(n52294) );
  AND U55872 ( .A(n919), .B(n55933), .Z(n55932) );
  XOR U55873 ( .A(n55934), .B(n55931), .Z(n55933) );
  XNOR U55874 ( .A(n52291), .B(n55927), .Z(n55929) );
  XOR U55875 ( .A(n55935), .B(n55936), .Z(n52291) );
  AND U55876 ( .A(n916), .B(n55937), .Z(n55936) );
  XOR U55877 ( .A(n55938), .B(n55935), .Z(n55937) );
  XOR U55878 ( .A(n55939), .B(n55940), .Z(n55927) );
  AND U55879 ( .A(n55941), .B(n55942), .Z(n55940) );
  XOR U55880 ( .A(n55939), .B(n52306), .Z(n55942) );
  XOR U55881 ( .A(n55943), .B(n55944), .Z(n52306) );
  AND U55882 ( .A(n919), .B(n55945), .Z(n55944) );
  XOR U55883 ( .A(n55946), .B(n55943), .Z(n55945) );
  XNOR U55884 ( .A(n52303), .B(n55939), .Z(n55941) );
  XOR U55885 ( .A(n55947), .B(n55948), .Z(n52303) );
  AND U55886 ( .A(n916), .B(n55949), .Z(n55948) );
  XOR U55887 ( .A(n55950), .B(n55947), .Z(n55949) );
  XOR U55888 ( .A(n55951), .B(n55952), .Z(n55939) );
  AND U55889 ( .A(n55953), .B(n55954), .Z(n55952) );
  XOR U55890 ( .A(n55951), .B(n52318), .Z(n55954) );
  XOR U55891 ( .A(n55955), .B(n55956), .Z(n52318) );
  AND U55892 ( .A(n919), .B(n55957), .Z(n55956) );
  XOR U55893 ( .A(n55958), .B(n55955), .Z(n55957) );
  XNOR U55894 ( .A(n52315), .B(n55951), .Z(n55953) );
  XOR U55895 ( .A(n55959), .B(n55960), .Z(n52315) );
  AND U55896 ( .A(n916), .B(n55961), .Z(n55960) );
  XOR U55897 ( .A(n55962), .B(n55959), .Z(n55961) );
  XOR U55898 ( .A(n55963), .B(n55964), .Z(n55951) );
  AND U55899 ( .A(n55965), .B(n55966), .Z(n55964) );
  XOR U55900 ( .A(n55963), .B(n52330), .Z(n55966) );
  XOR U55901 ( .A(n55967), .B(n55968), .Z(n52330) );
  AND U55902 ( .A(n919), .B(n55969), .Z(n55968) );
  XOR U55903 ( .A(n55970), .B(n55967), .Z(n55969) );
  XNOR U55904 ( .A(n52327), .B(n55963), .Z(n55965) );
  XOR U55905 ( .A(n55971), .B(n55972), .Z(n52327) );
  AND U55906 ( .A(n916), .B(n55973), .Z(n55972) );
  XOR U55907 ( .A(n55974), .B(n55971), .Z(n55973) );
  XOR U55908 ( .A(n55975), .B(n55976), .Z(n55963) );
  AND U55909 ( .A(n55977), .B(n55978), .Z(n55976) );
  XOR U55910 ( .A(n55975), .B(n52342), .Z(n55978) );
  XOR U55911 ( .A(n55979), .B(n55980), .Z(n52342) );
  AND U55912 ( .A(n919), .B(n55981), .Z(n55980) );
  XOR U55913 ( .A(n55982), .B(n55979), .Z(n55981) );
  XNOR U55914 ( .A(n52339), .B(n55975), .Z(n55977) );
  XOR U55915 ( .A(n55983), .B(n55984), .Z(n52339) );
  AND U55916 ( .A(n916), .B(n55985), .Z(n55984) );
  XOR U55917 ( .A(n55986), .B(n55983), .Z(n55985) );
  XOR U55918 ( .A(n55987), .B(n55988), .Z(n55975) );
  AND U55919 ( .A(n55989), .B(n55990), .Z(n55988) );
  XOR U55920 ( .A(n55987), .B(n52354), .Z(n55990) );
  XOR U55921 ( .A(n55991), .B(n55992), .Z(n52354) );
  AND U55922 ( .A(n919), .B(n55993), .Z(n55992) );
  XOR U55923 ( .A(n55994), .B(n55991), .Z(n55993) );
  XNOR U55924 ( .A(n52351), .B(n55987), .Z(n55989) );
  XOR U55925 ( .A(n55995), .B(n55996), .Z(n52351) );
  AND U55926 ( .A(n916), .B(n55997), .Z(n55996) );
  XOR U55927 ( .A(n55998), .B(n55995), .Z(n55997) );
  XOR U55928 ( .A(n55999), .B(n56000), .Z(n55987) );
  AND U55929 ( .A(n56001), .B(n56002), .Z(n56000) );
  XOR U55930 ( .A(n55999), .B(n52366), .Z(n56002) );
  XOR U55931 ( .A(n56003), .B(n56004), .Z(n52366) );
  AND U55932 ( .A(n919), .B(n56005), .Z(n56004) );
  XOR U55933 ( .A(n56006), .B(n56003), .Z(n56005) );
  XNOR U55934 ( .A(n52363), .B(n55999), .Z(n56001) );
  XOR U55935 ( .A(n56007), .B(n56008), .Z(n52363) );
  AND U55936 ( .A(n916), .B(n56009), .Z(n56008) );
  XOR U55937 ( .A(n56010), .B(n56007), .Z(n56009) );
  XOR U55938 ( .A(n56011), .B(n56012), .Z(n55999) );
  AND U55939 ( .A(n56013), .B(n56014), .Z(n56012) );
  XOR U55940 ( .A(n56011), .B(n52378), .Z(n56014) );
  XOR U55941 ( .A(n56015), .B(n56016), .Z(n52378) );
  AND U55942 ( .A(n919), .B(n56017), .Z(n56016) );
  XOR U55943 ( .A(n56018), .B(n56015), .Z(n56017) );
  XNOR U55944 ( .A(n52375), .B(n56011), .Z(n56013) );
  XOR U55945 ( .A(n56019), .B(n56020), .Z(n52375) );
  AND U55946 ( .A(n916), .B(n56021), .Z(n56020) );
  XOR U55947 ( .A(n56022), .B(n56019), .Z(n56021) );
  XOR U55948 ( .A(n56023), .B(n56024), .Z(n56011) );
  AND U55949 ( .A(n56025), .B(n56026), .Z(n56024) );
  XOR U55950 ( .A(n56023), .B(n52390), .Z(n56026) );
  XOR U55951 ( .A(n56027), .B(n56028), .Z(n52390) );
  AND U55952 ( .A(n919), .B(n56029), .Z(n56028) );
  XOR U55953 ( .A(n56030), .B(n56027), .Z(n56029) );
  XNOR U55954 ( .A(n52387), .B(n56023), .Z(n56025) );
  XOR U55955 ( .A(n56031), .B(n56032), .Z(n52387) );
  AND U55956 ( .A(n916), .B(n56033), .Z(n56032) );
  XOR U55957 ( .A(n56034), .B(n56031), .Z(n56033) );
  XOR U55958 ( .A(n56035), .B(n56036), .Z(n56023) );
  AND U55959 ( .A(n56037), .B(n56038), .Z(n56036) );
  XOR U55960 ( .A(n56035), .B(n52402), .Z(n56038) );
  XOR U55961 ( .A(n56039), .B(n56040), .Z(n52402) );
  AND U55962 ( .A(n919), .B(n56041), .Z(n56040) );
  XOR U55963 ( .A(n56042), .B(n56039), .Z(n56041) );
  XNOR U55964 ( .A(n52399), .B(n56035), .Z(n56037) );
  XOR U55965 ( .A(n56043), .B(n56044), .Z(n52399) );
  AND U55966 ( .A(n916), .B(n56045), .Z(n56044) );
  XOR U55967 ( .A(n56046), .B(n56043), .Z(n56045) );
  XOR U55968 ( .A(n56047), .B(n56048), .Z(n56035) );
  AND U55969 ( .A(n56049), .B(n56050), .Z(n56048) );
  XOR U55970 ( .A(n56047), .B(n52414), .Z(n56050) );
  XOR U55971 ( .A(n56051), .B(n56052), .Z(n52414) );
  AND U55972 ( .A(n919), .B(n56053), .Z(n56052) );
  XOR U55973 ( .A(n56054), .B(n56051), .Z(n56053) );
  XNOR U55974 ( .A(n52411), .B(n56047), .Z(n56049) );
  XOR U55975 ( .A(n56055), .B(n56056), .Z(n52411) );
  AND U55976 ( .A(n916), .B(n56057), .Z(n56056) );
  XOR U55977 ( .A(n56058), .B(n56055), .Z(n56057) );
  XOR U55978 ( .A(n56059), .B(n56060), .Z(n56047) );
  AND U55979 ( .A(n56061), .B(n56062), .Z(n56060) );
  XOR U55980 ( .A(n56059), .B(n52426), .Z(n56062) );
  XOR U55981 ( .A(n56063), .B(n56064), .Z(n52426) );
  AND U55982 ( .A(n919), .B(n56065), .Z(n56064) );
  XOR U55983 ( .A(n56066), .B(n56063), .Z(n56065) );
  XNOR U55984 ( .A(n52423), .B(n56059), .Z(n56061) );
  XOR U55985 ( .A(n56067), .B(n56068), .Z(n52423) );
  AND U55986 ( .A(n916), .B(n56069), .Z(n56068) );
  XOR U55987 ( .A(n56070), .B(n56067), .Z(n56069) );
  XOR U55988 ( .A(n56071), .B(n56072), .Z(n56059) );
  AND U55989 ( .A(n56073), .B(n56074), .Z(n56072) );
  XOR U55990 ( .A(n56071), .B(n52438), .Z(n56074) );
  XOR U55991 ( .A(n56075), .B(n56076), .Z(n52438) );
  AND U55992 ( .A(n919), .B(n56077), .Z(n56076) );
  XOR U55993 ( .A(n56078), .B(n56075), .Z(n56077) );
  XNOR U55994 ( .A(n52435), .B(n56071), .Z(n56073) );
  XOR U55995 ( .A(n56079), .B(n56080), .Z(n52435) );
  AND U55996 ( .A(n916), .B(n56081), .Z(n56080) );
  XOR U55997 ( .A(n56082), .B(n56079), .Z(n56081) );
  XOR U55998 ( .A(n56083), .B(n56084), .Z(n56071) );
  AND U55999 ( .A(n56085), .B(n56086), .Z(n56084) );
  XOR U56000 ( .A(n56083), .B(n52450), .Z(n56086) );
  XOR U56001 ( .A(n56087), .B(n56088), .Z(n52450) );
  AND U56002 ( .A(n919), .B(n56089), .Z(n56088) );
  XOR U56003 ( .A(n56090), .B(n56087), .Z(n56089) );
  XNOR U56004 ( .A(n52447), .B(n56083), .Z(n56085) );
  XOR U56005 ( .A(n56091), .B(n56092), .Z(n52447) );
  AND U56006 ( .A(n916), .B(n56093), .Z(n56092) );
  XOR U56007 ( .A(n56094), .B(n56091), .Z(n56093) );
  XOR U56008 ( .A(n56095), .B(n56096), .Z(n56083) );
  AND U56009 ( .A(n56097), .B(n56098), .Z(n56096) );
  XOR U56010 ( .A(n56095), .B(n52462), .Z(n56098) );
  XOR U56011 ( .A(n56099), .B(n56100), .Z(n52462) );
  AND U56012 ( .A(n919), .B(n56101), .Z(n56100) );
  XOR U56013 ( .A(n56102), .B(n56099), .Z(n56101) );
  XNOR U56014 ( .A(n52459), .B(n56095), .Z(n56097) );
  XOR U56015 ( .A(n56103), .B(n56104), .Z(n52459) );
  AND U56016 ( .A(n916), .B(n56105), .Z(n56104) );
  XOR U56017 ( .A(n56106), .B(n56103), .Z(n56105) );
  XOR U56018 ( .A(n56107), .B(n56108), .Z(n56095) );
  AND U56019 ( .A(n56109), .B(n56110), .Z(n56108) );
  XOR U56020 ( .A(n56107), .B(n52474), .Z(n56110) );
  XOR U56021 ( .A(n56111), .B(n56112), .Z(n52474) );
  AND U56022 ( .A(n919), .B(n56113), .Z(n56112) );
  XOR U56023 ( .A(n56114), .B(n56111), .Z(n56113) );
  XNOR U56024 ( .A(n52471), .B(n56107), .Z(n56109) );
  XOR U56025 ( .A(n56115), .B(n56116), .Z(n52471) );
  AND U56026 ( .A(n916), .B(n56117), .Z(n56116) );
  XOR U56027 ( .A(n56118), .B(n56115), .Z(n56117) );
  XOR U56028 ( .A(n56119), .B(n56120), .Z(n56107) );
  AND U56029 ( .A(n56121), .B(n56122), .Z(n56120) );
  XOR U56030 ( .A(n56119), .B(n52486), .Z(n56122) );
  XOR U56031 ( .A(n56123), .B(n56124), .Z(n52486) );
  AND U56032 ( .A(n919), .B(n56125), .Z(n56124) );
  XOR U56033 ( .A(n56126), .B(n56123), .Z(n56125) );
  XNOR U56034 ( .A(n52483), .B(n56119), .Z(n56121) );
  XOR U56035 ( .A(n56127), .B(n56128), .Z(n52483) );
  AND U56036 ( .A(n916), .B(n56129), .Z(n56128) );
  XOR U56037 ( .A(n56130), .B(n56127), .Z(n56129) );
  XOR U56038 ( .A(n56131), .B(n56132), .Z(n56119) );
  AND U56039 ( .A(n56133), .B(n56134), .Z(n56132) );
  XOR U56040 ( .A(n56131), .B(n52498), .Z(n56134) );
  XOR U56041 ( .A(n56135), .B(n56136), .Z(n52498) );
  AND U56042 ( .A(n919), .B(n56137), .Z(n56136) );
  XOR U56043 ( .A(n56138), .B(n56135), .Z(n56137) );
  XNOR U56044 ( .A(n52495), .B(n56131), .Z(n56133) );
  XOR U56045 ( .A(n56139), .B(n56140), .Z(n52495) );
  AND U56046 ( .A(n916), .B(n56141), .Z(n56140) );
  XOR U56047 ( .A(n56142), .B(n56139), .Z(n56141) );
  XOR U56048 ( .A(n56143), .B(n56144), .Z(n56131) );
  AND U56049 ( .A(n56145), .B(n56146), .Z(n56144) );
  XOR U56050 ( .A(n56143), .B(n52510), .Z(n56146) );
  XOR U56051 ( .A(n56147), .B(n56148), .Z(n52510) );
  AND U56052 ( .A(n919), .B(n56149), .Z(n56148) );
  XOR U56053 ( .A(n56150), .B(n56147), .Z(n56149) );
  XNOR U56054 ( .A(n52507), .B(n56143), .Z(n56145) );
  XOR U56055 ( .A(n56151), .B(n56152), .Z(n52507) );
  AND U56056 ( .A(n916), .B(n56153), .Z(n56152) );
  XOR U56057 ( .A(n56154), .B(n56151), .Z(n56153) );
  XOR U56058 ( .A(n56155), .B(n56156), .Z(n56143) );
  AND U56059 ( .A(n56157), .B(n56158), .Z(n56156) );
  XOR U56060 ( .A(n56155), .B(n52522), .Z(n56158) );
  XOR U56061 ( .A(n56159), .B(n56160), .Z(n52522) );
  AND U56062 ( .A(n919), .B(n56161), .Z(n56160) );
  XOR U56063 ( .A(n56162), .B(n56159), .Z(n56161) );
  XNOR U56064 ( .A(n52519), .B(n56155), .Z(n56157) );
  XOR U56065 ( .A(n56163), .B(n56164), .Z(n52519) );
  AND U56066 ( .A(n916), .B(n56165), .Z(n56164) );
  XOR U56067 ( .A(n56166), .B(n56163), .Z(n56165) );
  XOR U56068 ( .A(n56167), .B(n56168), .Z(n56155) );
  AND U56069 ( .A(n56169), .B(n56170), .Z(n56168) );
  XNOR U56070 ( .A(n56171), .B(n52535), .Z(n56170) );
  XOR U56071 ( .A(n56172), .B(n56173), .Z(n52535) );
  AND U56072 ( .A(n919), .B(n56174), .Z(n56173) );
  XOR U56073 ( .A(n56172), .B(n56175), .Z(n56174) );
  XNOR U56074 ( .A(n52532), .B(n56167), .Z(n56169) );
  XOR U56075 ( .A(n56176), .B(n56177), .Z(n52532) );
  AND U56076 ( .A(n916), .B(n56178), .Z(n56177) );
  XOR U56077 ( .A(n56176), .B(n56179), .Z(n56178) );
  IV U56078 ( .A(n56171), .Z(n56167) );
  AND U56079 ( .A(n55803), .B(n55806), .Z(n56171) );
  XNOR U56080 ( .A(n56180), .B(n56181), .Z(n55806) );
  AND U56081 ( .A(n919), .B(n56182), .Z(n56181) );
  XNOR U56082 ( .A(n56183), .B(n56180), .Z(n56182) );
  XOR U56083 ( .A(n56184), .B(n56185), .Z(n919) );
  AND U56084 ( .A(n56186), .B(n56187), .Z(n56185) );
  XOR U56085 ( .A(n56184), .B(n55814), .Z(n56187) );
  XNOR U56086 ( .A(n56188), .B(n56189), .Z(n55814) );
  AND U56087 ( .A(n56190), .B(n663), .Z(n56189) );
  AND U56088 ( .A(n56188), .B(n56191), .Z(n56190) );
  XNOR U56089 ( .A(n55811), .B(n56184), .Z(n56186) );
  XOR U56090 ( .A(n56192), .B(n56193), .Z(n55811) );
  AND U56091 ( .A(n56194), .B(n661), .Z(n56193) );
  NOR U56092 ( .A(n56192), .B(n56195), .Z(n56194) );
  XOR U56093 ( .A(n56196), .B(n56197), .Z(n56184) );
  AND U56094 ( .A(n56198), .B(n56199), .Z(n56197) );
  XOR U56095 ( .A(n56196), .B(n55826), .Z(n56199) );
  XOR U56096 ( .A(n56200), .B(n56201), .Z(n55826) );
  AND U56097 ( .A(n663), .B(n56202), .Z(n56201) );
  XOR U56098 ( .A(n56203), .B(n56200), .Z(n56202) );
  XNOR U56099 ( .A(n55823), .B(n56196), .Z(n56198) );
  XOR U56100 ( .A(n56204), .B(n56205), .Z(n55823) );
  AND U56101 ( .A(n661), .B(n56206), .Z(n56205) );
  XOR U56102 ( .A(n56207), .B(n56204), .Z(n56206) );
  XOR U56103 ( .A(n56208), .B(n56209), .Z(n56196) );
  AND U56104 ( .A(n56210), .B(n56211), .Z(n56209) );
  XOR U56105 ( .A(n56208), .B(n55838), .Z(n56211) );
  XOR U56106 ( .A(n56212), .B(n56213), .Z(n55838) );
  AND U56107 ( .A(n663), .B(n56214), .Z(n56213) );
  XOR U56108 ( .A(n56215), .B(n56212), .Z(n56214) );
  XNOR U56109 ( .A(n55835), .B(n56208), .Z(n56210) );
  XOR U56110 ( .A(n56216), .B(n56217), .Z(n55835) );
  AND U56111 ( .A(n661), .B(n56218), .Z(n56217) );
  XOR U56112 ( .A(n56219), .B(n56216), .Z(n56218) );
  XOR U56113 ( .A(n56220), .B(n56221), .Z(n56208) );
  AND U56114 ( .A(n56222), .B(n56223), .Z(n56221) );
  XOR U56115 ( .A(n56220), .B(n55850), .Z(n56223) );
  XOR U56116 ( .A(n56224), .B(n56225), .Z(n55850) );
  AND U56117 ( .A(n663), .B(n56226), .Z(n56225) );
  XOR U56118 ( .A(n56227), .B(n56224), .Z(n56226) );
  XNOR U56119 ( .A(n55847), .B(n56220), .Z(n56222) );
  XOR U56120 ( .A(n56228), .B(n56229), .Z(n55847) );
  AND U56121 ( .A(n661), .B(n56230), .Z(n56229) );
  XOR U56122 ( .A(n56231), .B(n56228), .Z(n56230) );
  XOR U56123 ( .A(n56232), .B(n56233), .Z(n56220) );
  AND U56124 ( .A(n56234), .B(n56235), .Z(n56233) );
  XOR U56125 ( .A(n56232), .B(n55862), .Z(n56235) );
  XOR U56126 ( .A(n56236), .B(n56237), .Z(n55862) );
  AND U56127 ( .A(n663), .B(n56238), .Z(n56237) );
  XOR U56128 ( .A(n56239), .B(n56236), .Z(n56238) );
  XNOR U56129 ( .A(n55859), .B(n56232), .Z(n56234) );
  XOR U56130 ( .A(n56240), .B(n56241), .Z(n55859) );
  AND U56131 ( .A(n661), .B(n56242), .Z(n56241) );
  XOR U56132 ( .A(n56243), .B(n56240), .Z(n56242) );
  XOR U56133 ( .A(n56244), .B(n56245), .Z(n56232) );
  AND U56134 ( .A(n56246), .B(n56247), .Z(n56245) );
  XOR U56135 ( .A(n56244), .B(n55874), .Z(n56247) );
  XOR U56136 ( .A(n56248), .B(n56249), .Z(n55874) );
  AND U56137 ( .A(n663), .B(n56250), .Z(n56249) );
  XOR U56138 ( .A(n56251), .B(n56248), .Z(n56250) );
  XNOR U56139 ( .A(n55871), .B(n56244), .Z(n56246) );
  XOR U56140 ( .A(n56252), .B(n56253), .Z(n55871) );
  AND U56141 ( .A(n661), .B(n56254), .Z(n56253) );
  XOR U56142 ( .A(n56255), .B(n56252), .Z(n56254) );
  XOR U56143 ( .A(n56256), .B(n56257), .Z(n56244) );
  AND U56144 ( .A(n56258), .B(n56259), .Z(n56257) );
  XOR U56145 ( .A(n56256), .B(n55886), .Z(n56259) );
  XOR U56146 ( .A(n56260), .B(n56261), .Z(n55886) );
  AND U56147 ( .A(n663), .B(n56262), .Z(n56261) );
  XOR U56148 ( .A(n56263), .B(n56260), .Z(n56262) );
  XNOR U56149 ( .A(n55883), .B(n56256), .Z(n56258) );
  XOR U56150 ( .A(n56264), .B(n56265), .Z(n55883) );
  AND U56151 ( .A(n661), .B(n56266), .Z(n56265) );
  XOR U56152 ( .A(n56267), .B(n56264), .Z(n56266) );
  XOR U56153 ( .A(n56268), .B(n56269), .Z(n56256) );
  AND U56154 ( .A(n56270), .B(n56271), .Z(n56269) );
  XOR U56155 ( .A(n56268), .B(n55898), .Z(n56271) );
  XOR U56156 ( .A(n56272), .B(n56273), .Z(n55898) );
  AND U56157 ( .A(n663), .B(n56274), .Z(n56273) );
  XOR U56158 ( .A(n56275), .B(n56272), .Z(n56274) );
  XNOR U56159 ( .A(n55895), .B(n56268), .Z(n56270) );
  XOR U56160 ( .A(n56276), .B(n56277), .Z(n55895) );
  AND U56161 ( .A(n661), .B(n56278), .Z(n56277) );
  XOR U56162 ( .A(n56279), .B(n56276), .Z(n56278) );
  XOR U56163 ( .A(n56280), .B(n56281), .Z(n56268) );
  AND U56164 ( .A(n56282), .B(n56283), .Z(n56281) );
  XOR U56165 ( .A(n56280), .B(n55910), .Z(n56283) );
  XOR U56166 ( .A(n56284), .B(n56285), .Z(n55910) );
  AND U56167 ( .A(n663), .B(n56286), .Z(n56285) );
  XOR U56168 ( .A(n56287), .B(n56284), .Z(n56286) );
  XNOR U56169 ( .A(n55907), .B(n56280), .Z(n56282) );
  XOR U56170 ( .A(n56288), .B(n56289), .Z(n55907) );
  AND U56171 ( .A(n661), .B(n56290), .Z(n56289) );
  XOR U56172 ( .A(n56291), .B(n56288), .Z(n56290) );
  XOR U56173 ( .A(n56292), .B(n56293), .Z(n56280) );
  AND U56174 ( .A(n56294), .B(n56295), .Z(n56293) );
  XOR U56175 ( .A(n56292), .B(n55922), .Z(n56295) );
  XOR U56176 ( .A(n56296), .B(n56297), .Z(n55922) );
  AND U56177 ( .A(n663), .B(n56298), .Z(n56297) );
  XOR U56178 ( .A(n56299), .B(n56296), .Z(n56298) );
  XNOR U56179 ( .A(n55919), .B(n56292), .Z(n56294) );
  XOR U56180 ( .A(n56300), .B(n56301), .Z(n55919) );
  AND U56181 ( .A(n661), .B(n56302), .Z(n56301) );
  XOR U56182 ( .A(n56303), .B(n56300), .Z(n56302) );
  XOR U56183 ( .A(n56304), .B(n56305), .Z(n56292) );
  AND U56184 ( .A(n56306), .B(n56307), .Z(n56305) );
  XOR U56185 ( .A(n56304), .B(n55934), .Z(n56307) );
  XOR U56186 ( .A(n56308), .B(n56309), .Z(n55934) );
  AND U56187 ( .A(n663), .B(n56310), .Z(n56309) );
  XOR U56188 ( .A(n56311), .B(n56308), .Z(n56310) );
  XNOR U56189 ( .A(n55931), .B(n56304), .Z(n56306) );
  XOR U56190 ( .A(n56312), .B(n56313), .Z(n55931) );
  AND U56191 ( .A(n661), .B(n56314), .Z(n56313) );
  XOR U56192 ( .A(n56315), .B(n56312), .Z(n56314) );
  XOR U56193 ( .A(n56316), .B(n56317), .Z(n56304) );
  AND U56194 ( .A(n56318), .B(n56319), .Z(n56317) );
  XOR U56195 ( .A(n56316), .B(n55946), .Z(n56319) );
  XOR U56196 ( .A(n56320), .B(n56321), .Z(n55946) );
  AND U56197 ( .A(n663), .B(n56322), .Z(n56321) );
  XOR U56198 ( .A(n56323), .B(n56320), .Z(n56322) );
  XNOR U56199 ( .A(n55943), .B(n56316), .Z(n56318) );
  XOR U56200 ( .A(n56324), .B(n56325), .Z(n55943) );
  AND U56201 ( .A(n661), .B(n56326), .Z(n56325) );
  XOR U56202 ( .A(n56327), .B(n56324), .Z(n56326) );
  XOR U56203 ( .A(n56328), .B(n56329), .Z(n56316) );
  AND U56204 ( .A(n56330), .B(n56331), .Z(n56329) );
  XOR U56205 ( .A(n56328), .B(n55958), .Z(n56331) );
  XOR U56206 ( .A(n56332), .B(n56333), .Z(n55958) );
  AND U56207 ( .A(n663), .B(n56334), .Z(n56333) );
  XOR U56208 ( .A(n56335), .B(n56332), .Z(n56334) );
  XNOR U56209 ( .A(n55955), .B(n56328), .Z(n56330) );
  XOR U56210 ( .A(n56336), .B(n56337), .Z(n55955) );
  AND U56211 ( .A(n661), .B(n56338), .Z(n56337) );
  XOR U56212 ( .A(n56339), .B(n56336), .Z(n56338) );
  XOR U56213 ( .A(n56340), .B(n56341), .Z(n56328) );
  AND U56214 ( .A(n56342), .B(n56343), .Z(n56341) );
  XOR U56215 ( .A(n56340), .B(n55970), .Z(n56343) );
  XOR U56216 ( .A(n56344), .B(n56345), .Z(n55970) );
  AND U56217 ( .A(n663), .B(n56346), .Z(n56345) );
  XOR U56218 ( .A(n56347), .B(n56344), .Z(n56346) );
  XNOR U56219 ( .A(n55967), .B(n56340), .Z(n56342) );
  XOR U56220 ( .A(n56348), .B(n56349), .Z(n55967) );
  AND U56221 ( .A(n661), .B(n56350), .Z(n56349) );
  XOR U56222 ( .A(n56351), .B(n56348), .Z(n56350) );
  XOR U56223 ( .A(n56352), .B(n56353), .Z(n56340) );
  AND U56224 ( .A(n56354), .B(n56355), .Z(n56353) );
  XOR U56225 ( .A(n56352), .B(n55982), .Z(n56355) );
  XOR U56226 ( .A(n56356), .B(n56357), .Z(n55982) );
  AND U56227 ( .A(n663), .B(n56358), .Z(n56357) );
  XOR U56228 ( .A(n56359), .B(n56356), .Z(n56358) );
  XNOR U56229 ( .A(n55979), .B(n56352), .Z(n56354) );
  XOR U56230 ( .A(n56360), .B(n56361), .Z(n55979) );
  AND U56231 ( .A(n661), .B(n56362), .Z(n56361) );
  XOR U56232 ( .A(n56363), .B(n56360), .Z(n56362) );
  XOR U56233 ( .A(n56364), .B(n56365), .Z(n56352) );
  AND U56234 ( .A(n56366), .B(n56367), .Z(n56365) );
  XOR U56235 ( .A(n56364), .B(n55994), .Z(n56367) );
  XOR U56236 ( .A(n56368), .B(n56369), .Z(n55994) );
  AND U56237 ( .A(n663), .B(n56370), .Z(n56369) );
  XOR U56238 ( .A(n56371), .B(n56368), .Z(n56370) );
  XNOR U56239 ( .A(n55991), .B(n56364), .Z(n56366) );
  XOR U56240 ( .A(n56372), .B(n56373), .Z(n55991) );
  AND U56241 ( .A(n661), .B(n56374), .Z(n56373) );
  XOR U56242 ( .A(n56375), .B(n56372), .Z(n56374) );
  XOR U56243 ( .A(n56376), .B(n56377), .Z(n56364) );
  AND U56244 ( .A(n56378), .B(n56379), .Z(n56377) );
  XOR U56245 ( .A(n56376), .B(n56006), .Z(n56379) );
  XOR U56246 ( .A(n56380), .B(n56381), .Z(n56006) );
  AND U56247 ( .A(n663), .B(n56382), .Z(n56381) );
  XOR U56248 ( .A(n56383), .B(n56380), .Z(n56382) );
  XNOR U56249 ( .A(n56003), .B(n56376), .Z(n56378) );
  XOR U56250 ( .A(n56384), .B(n56385), .Z(n56003) );
  AND U56251 ( .A(n661), .B(n56386), .Z(n56385) );
  XOR U56252 ( .A(n56387), .B(n56384), .Z(n56386) );
  XOR U56253 ( .A(n56388), .B(n56389), .Z(n56376) );
  AND U56254 ( .A(n56390), .B(n56391), .Z(n56389) );
  XOR U56255 ( .A(n56388), .B(n56018), .Z(n56391) );
  XOR U56256 ( .A(n56392), .B(n56393), .Z(n56018) );
  AND U56257 ( .A(n663), .B(n56394), .Z(n56393) );
  XOR U56258 ( .A(n56395), .B(n56392), .Z(n56394) );
  XNOR U56259 ( .A(n56015), .B(n56388), .Z(n56390) );
  XOR U56260 ( .A(n56396), .B(n56397), .Z(n56015) );
  AND U56261 ( .A(n661), .B(n56398), .Z(n56397) );
  XOR U56262 ( .A(n56399), .B(n56396), .Z(n56398) );
  XOR U56263 ( .A(n56400), .B(n56401), .Z(n56388) );
  AND U56264 ( .A(n56402), .B(n56403), .Z(n56401) );
  XOR U56265 ( .A(n56400), .B(n56030), .Z(n56403) );
  XOR U56266 ( .A(n56404), .B(n56405), .Z(n56030) );
  AND U56267 ( .A(n663), .B(n56406), .Z(n56405) );
  XOR U56268 ( .A(n56407), .B(n56404), .Z(n56406) );
  XNOR U56269 ( .A(n56027), .B(n56400), .Z(n56402) );
  XOR U56270 ( .A(n56408), .B(n56409), .Z(n56027) );
  AND U56271 ( .A(n661), .B(n56410), .Z(n56409) );
  XOR U56272 ( .A(n56411), .B(n56408), .Z(n56410) );
  XOR U56273 ( .A(n56412), .B(n56413), .Z(n56400) );
  AND U56274 ( .A(n56414), .B(n56415), .Z(n56413) );
  XOR U56275 ( .A(n56412), .B(n56042), .Z(n56415) );
  XOR U56276 ( .A(n56416), .B(n56417), .Z(n56042) );
  AND U56277 ( .A(n663), .B(n56418), .Z(n56417) );
  XOR U56278 ( .A(n56419), .B(n56416), .Z(n56418) );
  XNOR U56279 ( .A(n56039), .B(n56412), .Z(n56414) );
  XOR U56280 ( .A(n56420), .B(n56421), .Z(n56039) );
  AND U56281 ( .A(n661), .B(n56422), .Z(n56421) );
  XOR U56282 ( .A(n56423), .B(n56420), .Z(n56422) );
  XOR U56283 ( .A(n56424), .B(n56425), .Z(n56412) );
  AND U56284 ( .A(n56426), .B(n56427), .Z(n56425) );
  XOR U56285 ( .A(n56424), .B(n56054), .Z(n56427) );
  XOR U56286 ( .A(n56428), .B(n56429), .Z(n56054) );
  AND U56287 ( .A(n663), .B(n56430), .Z(n56429) );
  XOR U56288 ( .A(n56431), .B(n56428), .Z(n56430) );
  XNOR U56289 ( .A(n56051), .B(n56424), .Z(n56426) );
  XOR U56290 ( .A(n56432), .B(n56433), .Z(n56051) );
  AND U56291 ( .A(n661), .B(n56434), .Z(n56433) );
  XOR U56292 ( .A(n56435), .B(n56432), .Z(n56434) );
  XOR U56293 ( .A(n56436), .B(n56437), .Z(n56424) );
  AND U56294 ( .A(n56438), .B(n56439), .Z(n56437) );
  XOR U56295 ( .A(n56436), .B(n56066), .Z(n56439) );
  XOR U56296 ( .A(n56440), .B(n56441), .Z(n56066) );
  AND U56297 ( .A(n663), .B(n56442), .Z(n56441) );
  XOR U56298 ( .A(n56443), .B(n56440), .Z(n56442) );
  XNOR U56299 ( .A(n56063), .B(n56436), .Z(n56438) );
  XOR U56300 ( .A(n56444), .B(n56445), .Z(n56063) );
  AND U56301 ( .A(n661), .B(n56446), .Z(n56445) );
  XOR U56302 ( .A(n56447), .B(n56444), .Z(n56446) );
  XOR U56303 ( .A(n56448), .B(n56449), .Z(n56436) );
  AND U56304 ( .A(n56450), .B(n56451), .Z(n56449) );
  XOR U56305 ( .A(n56448), .B(n56078), .Z(n56451) );
  XOR U56306 ( .A(n56452), .B(n56453), .Z(n56078) );
  AND U56307 ( .A(n663), .B(n56454), .Z(n56453) );
  XOR U56308 ( .A(n56455), .B(n56452), .Z(n56454) );
  XNOR U56309 ( .A(n56075), .B(n56448), .Z(n56450) );
  XOR U56310 ( .A(n56456), .B(n56457), .Z(n56075) );
  AND U56311 ( .A(n661), .B(n56458), .Z(n56457) );
  XOR U56312 ( .A(n56459), .B(n56456), .Z(n56458) );
  XOR U56313 ( .A(n56460), .B(n56461), .Z(n56448) );
  AND U56314 ( .A(n56462), .B(n56463), .Z(n56461) );
  XOR U56315 ( .A(n56460), .B(n56090), .Z(n56463) );
  XOR U56316 ( .A(n56464), .B(n56465), .Z(n56090) );
  AND U56317 ( .A(n663), .B(n56466), .Z(n56465) );
  XOR U56318 ( .A(n56467), .B(n56464), .Z(n56466) );
  XNOR U56319 ( .A(n56087), .B(n56460), .Z(n56462) );
  XOR U56320 ( .A(n56468), .B(n56469), .Z(n56087) );
  AND U56321 ( .A(n661), .B(n56470), .Z(n56469) );
  XOR U56322 ( .A(n56471), .B(n56468), .Z(n56470) );
  XOR U56323 ( .A(n56472), .B(n56473), .Z(n56460) );
  AND U56324 ( .A(n56474), .B(n56475), .Z(n56473) );
  XOR U56325 ( .A(n56472), .B(n56102), .Z(n56475) );
  XOR U56326 ( .A(n56476), .B(n56477), .Z(n56102) );
  AND U56327 ( .A(n663), .B(n56478), .Z(n56477) );
  XOR U56328 ( .A(n56479), .B(n56476), .Z(n56478) );
  XNOR U56329 ( .A(n56099), .B(n56472), .Z(n56474) );
  XOR U56330 ( .A(n56480), .B(n56481), .Z(n56099) );
  AND U56331 ( .A(n661), .B(n56482), .Z(n56481) );
  XOR U56332 ( .A(n56483), .B(n56480), .Z(n56482) );
  XOR U56333 ( .A(n56484), .B(n56485), .Z(n56472) );
  AND U56334 ( .A(n56486), .B(n56487), .Z(n56485) );
  XOR U56335 ( .A(n56484), .B(n56114), .Z(n56487) );
  XOR U56336 ( .A(n56488), .B(n56489), .Z(n56114) );
  AND U56337 ( .A(n663), .B(n56490), .Z(n56489) );
  XOR U56338 ( .A(n56491), .B(n56488), .Z(n56490) );
  XNOR U56339 ( .A(n56111), .B(n56484), .Z(n56486) );
  XOR U56340 ( .A(n56492), .B(n56493), .Z(n56111) );
  AND U56341 ( .A(n661), .B(n56494), .Z(n56493) );
  XOR U56342 ( .A(n56495), .B(n56492), .Z(n56494) );
  XOR U56343 ( .A(n56496), .B(n56497), .Z(n56484) );
  AND U56344 ( .A(n56498), .B(n56499), .Z(n56497) );
  XOR U56345 ( .A(n56496), .B(n56126), .Z(n56499) );
  XOR U56346 ( .A(n56500), .B(n56501), .Z(n56126) );
  AND U56347 ( .A(n663), .B(n56502), .Z(n56501) );
  XOR U56348 ( .A(n56503), .B(n56500), .Z(n56502) );
  XNOR U56349 ( .A(n56123), .B(n56496), .Z(n56498) );
  XOR U56350 ( .A(n56504), .B(n56505), .Z(n56123) );
  AND U56351 ( .A(n661), .B(n56506), .Z(n56505) );
  XOR U56352 ( .A(n56507), .B(n56504), .Z(n56506) );
  XOR U56353 ( .A(n56508), .B(n56509), .Z(n56496) );
  AND U56354 ( .A(n56510), .B(n56511), .Z(n56509) );
  XOR U56355 ( .A(n56508), .B(n56138), .Z(n56511) );
  XOR U56356 ( .A(n56512), .B(n56513), .Z(n56138) );
  AND U56357 ( .A(n663), .B(n56514), .Z(n56513) );
  XOR U56358 ( .A(n56515), .B(n56512), .Z(n56514) );
  XNOR U56359 ( .A(n56135), .B(n56508), .Z(n56510) );
  XOR U56360 ( .A(n56516), .B(n56517), .Z(n56135) );
  AND U56361 ( .A(n661), .B(n56518), .Z(n56517) );
  XOR U56362 ( .A(n56519), .B(n56516), .Z(n56518) );
  XOR U56363 ( .A(n56520), .B(n56521), .Z(n56508) );
  AND U56364 ( .A(n56522), .B(n56523), .Z(n56521) );
  XOR U56365 ( .A(n56520), .B(n56150), .Z(n56523) );
  XOR U56366 ( .A(n56524), .B(n56525), .Z(n56150) );
  AND U56367 ( .A(n663), .B(n56526), .Z(n56525) );
  XOR U56368 ( .A(n56527), .B(n56524), .Z(n56526) );
  XNOR U56369 ( .A(n56147), .B(n56520), .Z(n56522) );
  XOR U56370 ( .A(n56528), .B(n56529), .Z(n56147) );
  AND U56371 ( .A(n661), .B(n56530), .Z(n56529) );
  XOR U56372 ( .A(n56531), .B(n56528), .Z(n56530) );
  XOR U56373 ( .A(n56532), .B(n56533), .Z(n56520) );
  AND U56374 ( .A(n56534), .B(n56535), .Z(n56533) );
  XOR U56375 ( .A(n56532), .B(n56162), .Z(n56535) );
  XOR U56376 ( .A(n56536), .B(n56537), .Z(n56162) );
  AND U56377 ( .A(n663), .B(n56538), .Z(n56537) );
  XOR U56378 ( .A(n56539), .B(n56536), .Z(n56538) );
  XNOR U56379 ( .A(n56159), .B(n56532), .Z(n56534) );
  XOR U56380 ( .A(n56540), .B(n56541), .Z(n56159) );
  AND U56381 ( .A(n661), .B(n56542), .Z(n56541) );
  XOR U56382 ( .A(n56543), .B(n56540), .Z(n56542) );
  XOR U56383 ( .A(n56544), .B(n56545), .Z(n56532) );
  AND U56384 ( .A(n56546), .B(n56547), .Z(n56545) );
  XNOR U56385 ( .A(n56548), .B(n56175), .Z(n56547) );
  XOR U56386 ( .A(n56549), .B(n56550), .Z(n56175) );
  AND U56387 ( .A(n663), .B(n56551), .Z(n56550) );
  XOR U56388 ( .A(n56549), .B(n56552), .Z(n56551) );
  XNOR U56389 ( .A(n56172), .B(n56544), .Z(n56546) );
  XOR U56390 ( .A(n56553), .B(n56554), .Z(n56172) );
  AND U56391 ( .A(n661), .B(n56555), .Z(n56554) );
  XOR U56392 ( .A(n56553), .B(n56556), .Z(n56555) );
  IV U56393 ( .A(n56548), .Z(n56544) );
  AND U56394 ( .A(n56180), .B(n56183), .Z(n56548) );
  XNOR U56395 ( .A(n56557), .B(n56558), .Z(n56183) );
  AND U56396 ( .A(n663), .B(n56559), .Z(n56558) );
  XNOR U56397 ( .A(n56560), .B(n56557), .Z(n56559) );
  XOR U56398 ( .A(n56561), .B(n56562), .Z(n663) );
  AND U56399 ( .A(n56563), .B(n56564), .Z(n56562) );
  XOR U56400 ( .A(n56191), .B(n56561), .Z(n56564) );
  IV U56401 ( .A(n56565), .Z(n56191) );
  AND U56402 ( .A(p_input[511]), .B(p_input[479]), .Z(n56565) );
  XOR U56403 ( .A(n56561), .B(n56188), .Z(n56563) );
  AND U56404 ( .A(p_input[415]), .B(p_input[447]), .Z(n56188) );
  XOR U56405 ( .A(n56566), .B(n56567), .Z(n56561) );
  AND U56406 ( .A(n56568), .B(n56569), .Z(n56567) );
  XOR U56407 ( .A(n56566), .B(n56203), .Z(n56569) );
  XNOR U56408 ( .A(p_input[478]), .B(n56570), .Z(n56203) );
  AND U56409 ( .A(n1115), .B(n56571), .Z(n56570) );
  XOR U56410 ( .A(p_input[510]), .B(p_input[478]), .Z(n56571) );
  XNOR U56411 ( .A(n56200), .B(n56566), .Z(n56568) );
  XOR U56412 ( .A(n56572), .B(n56573), .Z(n56200) );
  AND U56413 ( .A(n1113), .B(n56574), .Z(n56573) );
  XOR U56414 ( .A(p_input[446]), .B(p_input[414]), .Z(n56574) );
  XOR U56415 ( .A(n56575), .B(n56576), .Z(n56566) );
  AND U56416 ( .A(n56577), .B(n56578), .Z(n56576) );
  XOR U56417 ( .A(n56575), .B(n56215), .Z(n56578) );
  XNOR U56418 ( .A(p_input[477]), .B(n56579), .Z(n56215) );
  AND U56419 ( .A(n1115), .B(n56580), .Z(n56579) );
  XOR U56420 ( .A(p_input[509]), .B(p_input[477]), .Z(n56580) );
  XNOR U56421 ( .A(n56212), .B(n56575), .Z(n56577) );
  XOR U56422 ( .A(n56581), .B(n56582), .Z(n56212) );
  AND U56423 ( .A(n1113), .B(n56583), .Z(n56582) );
  XOR U56424 ( .A(p_input[445]), .B(p_input[413]), .Z(n56583) );
  XOR U56425 ( .A(n56584), .B(n56585), .Z(n56575) );
  AND U56426 ( .A(n56586), .B(n56587), .Z(n56585) );
  XOR U56427 ( .A(n56584), .B(n56227), .Z(n56587) );
  XNOR U56428 ( .A(p_input[476]), .B(n56588), .Z(n56227) );
  AND U56429 ( .A(n1115), .B(n56589), .Z(n56588) );
  XOR U56430 ( .A(p_input[508]), .B(p_input[476]), .Z(n56589) );
  XNOR U56431 ( .A(n56224), .B(n56584), .Z(n56586) );
  XOR U56432 ( .A(n56590), .B(n56591), .Z(n56224) );
  AND U56433 ( .A(n1113), .B(n56592), .Z(n56591) );
  XOR U56434 ( .A(p_input[444]), .B(p_input[412]), .Z(n56592) );
  XOR U56435 ( .A(n56593), .B(n56594), .Z(n56584) );
  AND U56436 ( .A(n56595), .B(n56596), .Z(n56594) );
  XOR U56437 ( .A(n56593), .B(n56239), .Z(n56596) );
  XNOR U56438 ( .A(p_input[475]), .B(n56597), .Z(n56239) );
  AND U56439 ( .A(n1115), .B(n56598), .Z(n56597) );
  XOR U56440 ( .A(p_input[507]), .B(p_input[475]), .Z(n56598) );
  XNOR U56441 ( .A(n56236), .B(n56593), .Z(n56595) );
  XOR U56442 ( .A(n56599), .B(n56600), .Z(n56236) );
  AND U56443 ( .A(n1113), .B(n56601), .Z(n56600) );
  XOR U56444 ( .A(p_input[443]), .B(p_input[411]), .Z(n56601) );
  XOR U56445 ( .A(n56602), .B(n56603), .Z(n56593) );
  AND U56446 ( .A(n56604), .B(n56605), .Z(n56603) );
  XOR U56447 ( .A(n56602), .B(n56251), .Z(n56605) );
  XNOR U56448 ( .A(p_input[474]), .B(n56606), .Z(n56251) );
  AND U56449 ( .A(n1115), .B(n56607), .Z(n56606) );
  XOR U56450 ( .A(p_input[506]), .B(p_input[474]), .Z(n56607) );
  XNOR U56451 ( .A(n56248), .B(n56602), .Z(n56604) );
  XOR U56452 ( .A(n56608), .B(n56609), .Z(n56248) );
  AND U56453 ( .A(n1113), .B(n56610), .Z(n56609) );
  XOR U56454 ( .A(p_input[442]), .B(p_input[410]), .Z(n56610) );
  XOR U56455 ( .A(n56611), .B(n56612), .Z(n56602) );
  AND U56456 ( .A(n56613), .B(n56614), .Z(n56612) );
  XOR U56457 ( .A(n56611), .B(n56263), .Z(n56614) );
  XNOR U56458 ( .A(p_input[473]), .B(n56615), .Z(n56263) );
  AND U56459 ( .A(n1115), .B(n56616), .Z(n56615) );
  XOR U56460 ( .A(p_input[505]), .B(p_input[473]), .Z(n56616) );
  XNOR U56461 ( .A(n56260), .B(n56611), .Z(n56613) );
  XOR U56462 ( .A(n56617), .B(n56618), .Z(n56260) );
  AND U56463 ( .A(n1113), .B(n56619), .Z(n56618) );
  XOR U56464 ( .A(p_input[441]), .B(p_input[409]), .Z(n56619) );
  XOR U56465 ( .A(n56620), .B(n56621), .Z(n56611) );
  AND U56466 ( .A(n56622), .B(n56623), .Z(n56621) );
  XOR U56467 ( .A(n56620), .B(n56275), .Z(n56623) );
  XNOR U56468 ( .A(p_input[472]), .B(n56624), .Z(n56275) );
  AND U56469 ( .A(n1115), .B(n56625), .Z(n56624) );
  XOR U56470 ( .A(p_input[504]), .B(p_input[472]), .Z(n56625) );
  XNOR U56471 ( .A(n56272), .B(n56620), .Z(n56622) );
  XOR U56472 ( .A(n56626), .B(n56627), .Z(n56272) );
  AND U56473 ( .A(n1113), .B(n56628), .Z(n56627) );
  XOR U56474 ( .A(p_input[440]), .B(p_input[408]), .Z(n56628) );
  XOR U56475 ( .A(n56629), .B(n56630), .Z(n56620) );
  AND U56476 ( .A(n56631), .B(n56632), .Z(n56630) );
  XOR U56477 ( .A(n56629), .B(n56287), .Z(n56632) );
  XNOR U56478 ( .A(p_input[471]), .B(n56633), .Z(n56287) );
  AND U56479 ( .A(n1115), .B(n56634), .Z(n56633) );
  XOR U56480 ( .A(p_input[503]), .B(p_input[471]), .Z(n56634) );
  XNOR U56481 ( .A(n56284), .B(n56629), .Z(n56631) );
  XOR U56482 ( .A(n56635), .B(n56636), .Z(n56284) );
  AND U56483 ( .A(n1113), .B(n56637), .Z(n56636) );
  XOR U56484 ( .A(p_input[439]), .B(p_input[407]), .Z(n56637) );
  XOR U56485 ( .A(n56638), .B(n56639), .Z(n56629) );
  AND U56486 ( .A(n56640), .B(n56641), .Z(n56639) );
  XOR U56487 ( .A(n56638), .B(n56299), .Z(n56641) );
  XNOR U56488 ( .A(p_input[470]), .B(n56642), .Z(n56299) );
  AND U56489 ( .A(n1115), .B(n56643), .Z(n56642) );
  XOR U56490 ( .A(p_input[502]), .B(p_input[470]), .Z(n56643) );
  XNOR U56491 ( .A(n56296), .B(n56638), .Z(n56640) );
  XOR U56492 ( .A(n56644), .B(n56645), .Z(n56296) );
  AND U56493 ( .A(n1113), .B(n56646), .Z(n56645) );
  XOR U56494 ( .A(p_input[438]), .B(p_input[406]), .Z(n56646) );
  XOR U56495 ( .A(n56647), .B(n56648), .Z(n56638) );
  AND U56496 ( .A(n56649), .B(n56650), .Z(n56648) );
  XOR U56497 ( .A(n56647), .B(n56311), .Z(n56650) );
  XNOR U56498 ( .A(p_input[469]), .B(n56651), .Z(n56311) );
  AND U56499 ( .A(n1115), .B(n56652), .Z(n56651) );
  XOR U56500 ( .A(p_input[501]), .B(p_input[469]), .Z(n56652) );
  XNOR U56501 ( .A(n56308), .B(n56647), .Z(n56649) );
  XOR U56502 ( .A(n56653), .B(n56654), .Z(n56308) );
  AND U56503 ( .A(n1113), .B(n56655), .Z(n56654) );
  XOR U56504 ( .A(p_input[437]), .B(p_input[405]), .Z(n56655) );
  XOR U56505 ( .A(n56656), .B(n56657), .Z(n56647) );
  AND U56506 ( .A(n56658), .B(n56659), .Z(n56657) );
  XOR U56507 ( .A(n56656), .B(n56323), .Z(n56659) );
  XNOR U56508 ( .A(p_input[468]), .B(n56660), .Z(n56323) );
  AND U56509 ( .A(n1115), .B(n56661), .Z(n56660) );
  XOR U56510 ( .A(p_input[500]), .B(p_input[468]), .Z(n56661) );
  XNOR U56511 ( .A(n56320), .B(n56656), .Z(n56658) );
  XOR U56512 ( .A(n56662), .B(n56663), .Z(n56320) );
  AND U56513 ( .A(n1113), .B(n56664), .Z(n56663) );
  XOR U56514 ( .A(p_input[436]), .B(p_input[404]), .Z(n56664) );
  XOR U56515 ( .A(n56665), .B(n56666), .Z(n56656) );
  AND U56516 ( .A(n56667), .B(n56668), .Z(n56666) );
  XOR U56517 ( .A(n56665), .B(n56335), .Z(n56668) );
  XNOR U56518 ( .A(p_input[467]), .B(n56669), .Z(n56335) );
  AND U56519 ( .A(n1115), .B(n56670), .Z(n56669) );
  XOR U56520 ( .A(p_input[499]), .B(p_input[467]), .Z(n56670) );
  XNOR U56521 ( .A(n56332), .B(n56665), .Z(n56667) );
  XOR U56522 ( .A(n56671), .B(n56672), .Z(n56332) );
  AND U56523 ( .A(n1113), .B(n56673), .Z(n56672) );
  XOR U56524 ( .A(p_input[435]), .B(p_input[403]), .Z(n56673) );
  XOR U56525 ( .A(n56674), .B(n56675), .Z(n56665) );
  AND U56526 ( .A(n56676), .B(n56677), .Z(n56675) );
  XOR U56527 ( .A(n56674), .B(n56347), .Z(n56677) );
  XNOR U56528 ( .A(p_input[466]), .B(n56678), .Z(n56347) );
  AND U56529 ( .A(n1115), .B(n56679), .Z(n56678) );
  XOR U56530 ( .A(p_input[498]), .B(p_input[466]), .Z(n56679) );
  XNOR U56531 ( .A(n56344), .B(n56674), .Z(n56676) );
  XOR U56532 ( .A(n56680), .B(n56681), .Z(n56344) );
  AND U56533 ( .A(n1113), .B(n56682), .Z(n56681) );
  XOR U56534 ( .A(p_input[434]), .B(p_input[402]), .Z(n56682) );
  XOR U56535 ( .A(n56683), .B(n56684), .Z(n56674) );
  AND U56536 ( .A(n56685), .B(n56686), .Z(n56684) );
  XOR U56537 ( .A(n56683), .B(n56359), .Z(n56686) );
  XNOR U56538 ( .A(p_input[465]), .B(n56687), .Z(n56359) );
  AND U56539 ( .A(n1115), .B(n56688), .Z(n56687) );
  XOR U56540 ( .A(p_input[497]), .B(p_input[465]), .Z(n56688) );
  XNOR U56541 ( .A(n56356), .B(n56683), .Z(n56685) );
  XOR U56542 ( .A(n56689), .B(n56690), .Z(n56356) );
  AND U56543 ( .A(n1113), .B(n56691), .Z(n56690) );
  XOR U56544 ( .A(p_input[433]), .B(p_input[401]), .Z(n56691) );
  XOR U56545 ( .A(n56692), .B(n56693), .Z(n56683) );
  AND U56546 ( .A(n56694), .B(n56695), .Z(n56693) );
  XOR U56547 ( .A(n56692), .B(n56371), .Z(n56695) );
  XNOR U56548 ( .A(p_input[464]), .B(n56696), .Z(n56371) );
  AND U56549 ( .A(n1115), .B(n56697), .Z(n56696) );
  XOR U56550 ( .A(p_input[496]), .B(p_input[464]), .Z(n56697) );
  XNOR U56551 ( .A(n56368), .B(n56692), .Z(n56694) );
  XOR U56552 ( .A(n56698), .B(n56699), .Z(n56368) );
  AND U56553 ( .A(n1113), .B(n56700), .Z(n56699) );
  XOR U56554 ( .A(p_input[432]), .B(p_input[400]), .Z(n56700) );
  XOR U56555 ( .A(n56701), .B(n56702), .Z(n56692) );
  AND U56556 ( .A(n56703), .B(n56704), .Z(n56702) );
  XOR U56557 ( .A(n56701), .B(n56383), .Z(n56704) );
  XNOR U56558 ( .A(p_input[463]), .B(n56705), .Z(n56383) );
  AND U56559 ( .A(n1115), .B(n56706), .Z(n56705) );
  XOR U56560 ( .A(p_input[495]), .B(p_input[463]), .Z(n56706) );
  XNOR U56561 ( .A(n56380), .B(n56701), .Z(n56703) );
  XOR U56562 ( .A(n56707), .B(n56708), .Z(n56380) );
  AND U56563 ( .A(n1113), .B(n56709), .Z(n56708) );
  XOR U56564 ( .A(p_input[431]), .B(p_input[399]), .Z(n56709) );
  XOR U56565 ( .A(n56710), .B(n56711), .Z(n56701) );
  AND U56566 ( .A(n56712), .B(n56713), .Z(n56711) );
  XOR U56567 ( .A(n56710), .B(n56395), .Z(n56713) );
  XNOR U56568 ( .A(p_input[462]), .B(n56714), .Z(n56395) );
  AND U56569 ( .A(n1115), .B(n56715), .Z(n56714) );
  XOR U56570 ( .A(p_input[494]), .B(p_input[462]), .Z(n56715) );
  XNOR U56571 ( .A(n56392), .B(n56710), .Z(n56712) );
  XOR U56572 ( .A(n56716), .B(n56717), .Z(n56392) );
  AND U56573 ( .A(n1113), .B(n56718), .Z(n56717) );
  XOR U56574 ( .A(p_input[430]), .B(p_input[398]), .Z(n56718) );
  XOR U56575 ( .A(n56719), .B(n56720), .Z(n56710) );
  AND U56576 ( .A(n56721), .B(n56722), .Z(n56720) );
  XOR U56577 ( .A(n56719), .B(n56407), .Z(n56722) );
  XNOR U56578 ( .A(p_input[461]), .B(n56723), .Z(n56407) );
  AND U56579 ( .A(n1115), .B(n56724), .Z(n56723) );
  XOR U56580 ( .A(p_input[493]), .B(p_input[461]), .Z(n56724) );
  XNOR U56581 ( .A(n56404), .B(n56719), .Z(n56721) );
  XOR U56582 ( .A(n56725), .B(n56726), .Z(n56404) );
  AND U56583 ( .A(n1113), .B(n56727), .Z(n56726) );
  XOR U56584 ( .A(p_input[429]), .B(p_input[397]), .Z(n56727) );
  XOR U56585 ( .A(n56728), .B(n56729), .Z(n56719) );
  AND U56586 ( .A(n56730), .B(n56731), .Z(n56729) );
  XOR U56587 ( .A(n56728), .B(n56419), .Z(n56731) );
  XNOR U56588 ( .A(p_input[460]), .B(n56732), .Z(n56419) );
  AND U56589 ( .A(n1115), .B(n56733), .Z(n56732) );
  XOR U56590 ( .A(p_input[492]), .B(p_input[460]), .Z(n56733) );
  XNOR U56591 ( .A(n56416), .B(n56728), .Z(n56730) );
  XOR U56592 ( .A(n56734), .B(n56735), .Z(n56416) );
  AND U56593 ( .A(n1113), .B(n56736), .Z(n56735) );
  XOR U56594 ( .A(p_input[428]), .B(p_input[396]), .Z(n56736) );
  XOR U56595 ( .A(n56737), .B(n56738), .Z(n56728) );
  AND U56596 ( .A(n56739), .B(n56740), .Z(n56738) );
  XOR U56597 ( .A(n56737), .B(n56431), .Z(n56740) );
  XNOR U56598 ( .A(p_input[459]), .B(n56741), .Z(n56431) );
  AND U56599 ( .A(n1115), .B(n56742), .Z(n56741) );
  XOR U56600 ( .A(p_input[491]), .B(p_input[459]), .Z(n56742) );
  XNOR U56601 ( .A(n56428), .B(n56737), .Z(n56739) );
  XOR U56602 ( .A(n56743), .B(n56744), .Z(n56428) );
  AND U56603 ( .A(n1113), .B(n56745), .Z(n56744) );
  XOR U56604 ( .A(p_input[427]), .B(p_input[395]), .Z(n56745) );
  XOR U56605 ( .A(n56746), .B(n56747), .Z(n56737) );
  AND U56606 ( .A(n56748), .B(n56749), .Z(n56747) );
  XOR U56607 ( .A(n56746), .B(n56443), .Z(n56749) );
  XNOR U56608 ( .A(p_input[458]), .B(n56750), .Z(n56443) );
  AND U56609 ( .A(n1115), .B(n56751), .Z(n56750) );
  XOR U56610 ( .A(p_input[490]), .B(p_input[458]), .Z(n56751) );
  XNOR U56611 ( .A(n56440), .B(n56746), .Z(n56748) );
  XOR U56612 ( .A(n56752), .B(n56753), .Z(n56440) );
  AND U56613 ( .A(n1113), .B(n56754), .Z(n56753) );
  XOR U56614 ( .A(p_input[426]), .B(p_input[394]), .Z(n56754) );
  XOR U56615 ( .A(n56755), .B(n56756), .Z(n56746) );
  AND U56616 ( .A(n56757), .B(n56758), .Z(n56756) );
  XOR U56617 ( .A(n56755), .B(n56455), .Z(n56758) );
  XNOR U56618 ( .A(p_input[457]), .B(n56759), .Z(n56455) );
  AND U56619 ( .A(n1115), .B(n56760), .Z(n56759) );
  XOR U56620 ( .A(p_input[489]), .B(p_input[457]), .Z(n56760) );
  XNOR U56621 ( .A(n56452), .B(n56755), .Z(n56757) );
  XOR U56622 ( .A(n56761), .B(n56762), .Z(n56452) );
  AND U56623 ( .A(n1113), .B(n56763), .Z(n56762) );
  XOR U56624 ( .A(p_input[425]), .B(p_input[393]), .Z(n56763) );
  XOR U56625 ( .A(n56764), .B(n56765), .Z(n56755) );
  AND U56626 ( .A(n56766), .B(n56767), .Z(n56765) );
  XOR U56627 ( .A(n56764), .B(n56467), .Z(n56767) );
  XNOR U56628 ( .A(p_input[456]), .B(n56768), .Z(n56467) );
  AND U56629 ( .A(n1115), .B(n56769), .Z(n56768) );
  XOR U56630 ( .A(p_input[488]), .B(p_input[456]), .Z(n56769) );
  XNOR U56631 ( .A(n56464), .B(n56764), .Z(n56766) );
  XOR U56632 ( .A(n56770), .B(n56771), .Z(n56464) );
  AND U56633 ( .A(n1113), .B(n56772), .Z(n56771) );
  XOR U56634 ( .A(p_input[424]), .B(p_input[392]), .Z(n56772) );
  XOR U56635 ( .A(n56773), .B(n56774), .Z(n56764) );
  AND U56636 ( .A(n56775), .B(n56776), .Z(n56774) );
  XOR U56637 ( .A(n56773), .B(n56479), .Z(n56776) );
  XNOR U56638 ( .A(p_input[455]), .B(n56777), .Z(n56479) );
  AND U56639 ( .A(n1115), .B(n56778), .Z(n56777) );
  XOR U56640 ( .A(p_input[487]), .B(p_input[455]), .Z(n56778) );
  XNOR U56641 ( .A(n56476), .B(n56773), .Z(n56775) );
  XOR U56642 ( .A(n56779), .B(n56780), .Z(n56476) );
  AND U56643 ( .A(n1113), .B(n56781), .Z(n56780) );
  XOR U56644 ( .A(p_input[423]), .B(p_input[391]), .Z(n56781) );
  XOR U56645 ( .A(n56782), .B(n56783), .Z(n56773) );
  AND U56646 ( .A(n56784), .B(n56785), .Z(n56783) );
  XOR U56647 ( .A(n56782), .B(n56491), .Z(n56785) );
  XNOR U56648 ( .A(p_input[454]), .B(n56786), .Z(n56491) );
  AND U56649 ( .A(n1115), .B(n56787), .Z(n56786) );
  XOR U56650 ( .A(p_input[486]), .B(p_input[454]), .Z(n56787) );
  XNOR U56651 ( .A(n56488), .B(n56782), .Z(n56784) );
  XOR U56652 ( .A(n56788), .B(n56789), .Z(n56488) );
  AND U56653 ( .A(n1113), .B(n56790), .Z(n56789) );
  XOR U56654 ( .A(p_input[422]), .B(p_input[390]), .Z(n56790) );
  XOR U56655 ( .A(n56791), .B(n56792), .Z(n56782) );
  AND U56656 ( .A(n56793), .B(n56794), .Z(n56792) );
  XOR U56657 ( .A(n56791), .B(n56503), .Z(n56794) );
  XNOR U56658 ( .A(p_input[453]), .B(n56795), .Z(n56503) );
  AND U56659 ( .A(n1115), .B(n56796), .Z(n56795) );
  XOR U56660 ( .A(p_input[485]), .B(p_input[453]), .Z(n56796) );
  XNOR U56661 ( .A(n56500), .B(n56791), .Z(n56793) );
  XOR U56662 ( .A(n56797), .B(n56798), .Z(n56500) );
  AND U56663 ( .A(n1113), .B(n56799), .Z(n56798) );
  XOR U56664 ( .A(p_input[421]), .B(p_input[389]), .Z(n56799) );
  XOR U56665 ( .A(n56800), .B(n56801), .Z(n56791) );
  AND U56666 ( .A(n56802), .B(n56803), .Z(n56801) );
  XOR U56667 ( .A(n56800), .B(n56515), .Z(n56803) );
  XNOR U56668 ( .A(p_input[452]), .B(n56804), .Z(n56515) );
  AND U56669 ( .A(n1115), .B(n56805), .Z(n56804) );
  XOR U56670 ( .A(p_input[484]), .B(p_input[452]), .Z(n56805) );
  XNOR U56671 ( .A(n56512), .B(n56800), .Z(n56802) );
  XOR U56672 ( .A(n56806), .B(n56807), .Z(n56512) );
  AND U56673 ( .A(n1113), .B(n56808), .Z(n56807) );
  XOR U56674 ( .A(p_input[420]), .B(p_input[388]), .Z(n56808) );
  XOR U56675 ( .A(n56809), .B(n56810), .Z(n56800) );
  AND U56676 ( .A(n56811), .B(n56812), .Z(n56810) );
  XOR U56677 ( .A(n56809), .B(n56527), .Z(n56812) );
  XNOR U56678 ( .A(p_input[451]), .B(n56813), .Z(n56527) );
  AND U56679 ( .A(n1115), .B(n56814), .Z(n56813) );
  XOR U56680 ( .A(p_input[483]), .B(p_input[451]), .Z(n56814) );
  XNOR U56681 ( .A(n56524), .B(n56809), .Z(n56811) );
  XOR U56682 ( .A(n56815), .B(n56816), .Z(n56524) );
  AND U56683 ( .A(n1113), .B(n56817), .Z(n56816) );
  XOR U56684 ( .A(p_input[419]), .B(p_input[387]), .Z(n56817) );
  XOR U56685 ( .A(n56818), .B(n56819), .Z(n56809) );
  AND U56686 ( .A(n56820), .B(n56821), .Z(n56819) );
  XOR U56687 ( .A(n56818), .B(n56539), .Z(n56821) );
  XNOR U56688 ( .A(p_input[450]), .B(n56822), .Z(n56539) );
  AND U56689 ( .A(n1115), .B(n56823), .Z(n56822) );
  XOR U56690 ( .A(p_input[482]), .B(p_input[450]), .Z(n56823) );
  XNOR U56691 ( .A(n56536), .B(n56818), .Z(n56820) );
  XOR U56692 ( .A(n56824), .B(n56825), .Z(n56536) );
  AND U56693 ( .A(n1113), .B(n56826), .Z(n56825) );
  XOR U56694 ( .A(p_input[418]), .B(p_input[386]), .Z(n56826) );
  XOR U56695 ( .A(n56827), .B(n56828), .Z(n56818) );
  AND U56696 ( .A(n56829), .B(n56830), .Z(n56828) );
  XNOR U56697 ( .A(n56831), .B(n56552), .Z(n56830) );
  XNOR U56698 ( .A(p_input[449]), .B(n56832), .Z(n56552) );
  AND U56699 ( .A(n1115), .B(n56833), .Z(n56832) );
  XNOR U56700 ( .A(p_input[481]), .B(n56834), .Z(n56833) );
  IV U56701 ( .A(p_input[449]), .Z(n56834) );
  XNOR U56702 ( .A(n56549), .B(n56827), .Z(n56829) );
  XNOR U56703 ( .A(p_input[385]), .B(n56835), .Z(n56549) );
  AND U56704 ( .A(n1113), .B(n56836), .Z(n56835) );
  XOR U56705 ( .A(p_input[417]), .B(p_input[385]), .Z(n56836) );
  IV U56706 ( .A(n56831), .Z(n56827) );
  AND U56707 ( .A(n56557), .B(n56560), .Z(n56831) );
  XOR U56708 ( .A(p_input[448]), .B(n56837), .Z(n56560) );
  AND U56709 ( .A(n1115), .B(n56838), .Z(n56837) );
  XOR U56710 ( .A(p_input[480]), .B(p_input[448]), .Z(n56838) );
  XOR U56711 ( .A(n56839), .B(n56840), .Z(n1115) );
  AND U56712 ( .A(n56841), .B(n56842), .Z(n56840) );
  XNOR U56713 ( .A(p_input[511]), .B(n56839), .Z(n56842) );
  XOR U56714 ( .A(n56839), .B(p_input[479]), .Z(n56841) );
  XOR U56715 ( .A(n56843), .B(n56844), .Z(n56839) );
  AND U56716 ( .A(n56845), .B(n56846), .Z(n56844) );
  XNOR U56717 ( .A(p_input[510]), .B(n56843), .Z(n56846) );
  XOR U56718 ( .A(n56843), .B(p_input[478]), .Z(n56845) );
  XOR U56719 ( .A(n56847), .B(n56848), .Z(n56843) );
  AND U56720 ( .A(n56849), .B(n56850), .Z(n56848) );
  XNOR U56721 ( .A(p_input[509]), .B(n56847), .Z(n56850) );
  XOR U56722 ( .A(n56847), .B(p_input[477]), .Z(n56849) );
  XOR U56723 ( .A(n56851), .B(n56852), .Z(n56847) );
  AND U56724 ( .A(n56853), .B(n56854), .Z(n56852) );
  XNOR U56725 ( .A(p_input[508]), .B(n56851), .Z(n56854) );
  XOR U56726 ( .A(n56851), .B(p_input[476]), .Z(n56853) );
  XOR U56727 ( .A(n56855), .B(n56856), .Z(n56851) );
  AND U56728 ( .A(n56857), .B(n56858), .Z(n56856) );
  XNOR U56729 ( .A(p_input[507]), .B(n56855), .Z(n56858) );
  XOR U56730 ( .A(n56855), .B(p_input[475]), .Z(n56857) );
  XOR U56731 ( .A(n56859), .B(n56860), .Z(n56855) );
  AND U56732 ( .A(n56861), .B(n56862), .Z(n56860) );
  XNOR U56733 ( .A(p_input[506]), .B(n56859), .Z(n56862) );
  XOR U56734 ( .A(n56859), .B(p_input[474]), .Z(n56861) );
  XOR U56735 ( .A(n56863), .B(n56864), .Z(n56859) );
  AND U56736 ( .A(n56865), .B(n56866), .Z(n56864) );
  XNOR U56737 ( .A(p_input[505]), .B(n56863), .Z(n56866) );
  XOR U56738 ( .A(n56863), .B(p_input[473]), .Z(n56865) );
  XOR U56739 ( .A(n56867), .B(n56868), .Z(n56863) );
  AND U56740 ( .A(n56869), .B(n56870), .Z(n56868) );
  XNOR U56741 ( .A(p_input[504]), .B(n56867), .Z(n56870) );
  XOR U56742 ( .A(n56867), .B(p_input[472]), .Z(n56869) );
  XOR U56743 ( .A(n56871), .B(n56872), .Z(n56867) );
  AND U56744 ( .A(n56873), .B(n56874), .Z(n56872) );
  XNOR U56745 ( .A(p_input[503]), .B(n56871), .Z(n56874) );
  XOR U56746 ( .A(n56871), .B(p_input[471]), .Z(n56873) );
  XOR U56747 ( .A(n56875), .B(n56876), .Z(n56871) );
  AND U56748 ( .A(n56877), .B(n56878), .Z(n56876) );
  XNOR U56749 ( .A(p_input[502]), .B(n56875), .Z(n56878) );
  XOR U56750 ( .A(n56875), .B(p_input[470]), .Z(n56877) );
  XOR U56751 ( .A(n56879), .B(n56880), .Z(n56875) );
  AND U56752 ( .A(n56881), .B(n56882), .Z(n56880) );
  XNOR U56753 ( .A(p_input[501]), .B(n56879), .Z(n56882) );
  XOR U56754 ( .A(n56879), .B(p_input[469]), .Z(n56881) );
  XOR U56755 ( .A(n56883), .B(n56884), .Z(n56879) );
  AND U56756 ( .A(n56885), .B(n56886), .Z(n56884) );
  XNOR U56757 ( .A(p_input[500]), .B(n56883), .Z(n56886) );
  XOR U56758 ( .A(n56883), .B(p_input[468]), .Z(n56885) );
  XOR U56759 ( .A(n56887), .B(n56888), .Z(n56883) );
  AND U56760 ( .A(n56889), .B(n56890), .Z(n56888) );
  XNOR U56761 ( .A(p_input[499]), .B(n56887), .Z(n56890) );
  XOR U56762 ( .A(n56887), .B(p_input[467]), .Z(n56889) );
  XOR U56763 ( .A(n56891), .B(n56892), .Z(n56887) );
  AND U56764 ( .A(n56893), .B(n56894), .Z(n56892) );
  XNOR U56765 ( .A(p_input[498]), .B(n56891), .Z(n56894) );
  XOR U56766 ( .A(n56891), .B(p_input[466]), .Z(n56893) );
  XOR U56767 ( .A(n56895), .B(n56896), .Z(n56891) );
  AND U56768 ( .A(n56897), .B(n56898), .Z(n56896) );
  XNOR U56769 ( .A(p_input[497]), .B(n56895), .Z(n56898) );
  XOR U56770 ( .A(n56895), .B(p_input[465]), .Z(n56897) );
  XOR U56771 ( .A(n56899), .B(n56900), .Z(n56895) );
  AND U56772 ( .A(n56901), .B(n56902), .Z(n56900) );
  XNOR U56773 ( .A(p_input[496]), .B(n56899), .Z(n56902) );
  XOR U56774 ( .A(n56899), .B(p_input[464]), .Z(n56901) );
  XOR U56775 ( .A(n56903), .B(n56904), .Z(n56899) );
  AND U56776 ( .A(n56905), .B(n56906), .Z(n56904) );
  XNOR U56777 ( .A(p_input[495]), .B(n56903), .Z(n56906) );
  XOR U56778 ( .A(n56903), .B(p_input[463]), .Z(n56905) );
  XOR U56779 ( .A(n56907), .B(n56908), .Z(n56903) );
  AND U56780 ( .A(n56909), .B(n56910), .Z(n56908) );
  XNOR U56781 ( .A(p_input[494]), .B(n56907), .Z(n56910) );
  XOR U56782 ( .A(n56907), .B(p_input[462]), .Z(n56909) );
  XOR U56783 ( .A(n56911), .B(n56912), .Z(n56907) );
  AND U56784 ( .A(n56913), .B(n56914), .Z(n56912) );
  XNOR U56785 ( .A(p_input[493]), .B(n56911), .Z(n56914) );
  XOR U56786 ( .A(n56911), .B(p_input[461]), .Z(n56913) );
  XOR U56787 ( .A(n56915), .B(n56916), .Z(n56911) );
  AND U56788 ( .A(n56917), .B(n56918), .Z(n56916) );
  XNOR U56789 ( .A(p_input[492]), .B(n56915), .Z(n56918) );
  XOR U56790 ( .A(n56915), .B(p_input[460]), .Z(n56917) );
  XOR U56791 ( .A(n56919), .B(n56920), .Z(n56915) );
  AND U56792 ( .A(n56921), .B(n56922), .Z(n56920) );
  XNOR U56793 ( .A(p_input[491]), .B(n56919), .Z(n56922) );
  XOR U56794 ( .A(n56919), .B(p_input[459]), .Z(n56921) );
  XOR U56795 ( .A(n56923), .B(n56924), .Z(n56919) );
  AND U56796 ( .A(n56925), .B(n56926), .Z(n56924) );
  XNOR U56797 ( .A(p_input[490]), .B(n56923), .Z(n56926) );
  XOR U56798 ( .A(n56923), .B(p_input[458]), .Z(n56925) );
  XOR U56799 ( .A(n56927), .B(n56928), .Z(n56923) );
  AND U56800 ( .A(n56929), .B(n56930), .Z(n56928) );
  XNOR U56801 ( .A(p_input[489]), .B(n56927), .Z(n56930) );
  XOR U56802 ( .A(n56927), .B(p_input[457]), .Z(n56929) );
  XOR U56803 ( .A(n56931), .B(n56932), .Z(n56927) );
  AND U56804 ( .A(n56933), .B(n56934), .Z(n56932) );
  XNOR U56805 ( .A(p_input[488]), .B(n56931), .Z(n56934) );
  XOR U56806 ( .A(n56931), .B(p_input[456]), .Z(n56933) );
  XOR U56807 ( .A(n56935), .B(n56936), .Z(n56931) );
  AND U56808 ( .A(n56937), .B(n56938), .Z(n56936) );
  XNOR U56809 ( .A(p_input[487]), .B(n56935), .Z(n56938) );
  XOR U56810 ( .A(n56935), .B(p_input[455]), .Z(n56937) );
  XOR U56811 ( .A(n56939), .B(n56940), .Z(n56935) );
  AND U56812 ( .A(n56941), .B(n56942), .Z(n56940) );
  XNOR U56813 ( .A(p_input[486]), .B(n56939), .Z(n56942) );
  XOR U56814 ( .A(n56939), .B(p_input[454]), .Z(n56941) );
  XOR U56815 ( .A(n56943), .B(n56944), .Z(n56939) );
  AND U56816 ( .A(n56945), .B(n56946), .Z(n56944) );
  XNOR U56817 ( .A(p_input[485]), .B(n56943), .Z(n56946) );
  XOR U56818 ( .A(n56943), .B(p_input[453]), .Z(n56945) );
  XOR U56819 ( .A(n56947), .B(n56948), .Z(n56943) );
  AND U56820 ( .A(n56949), .B(n56950), .Z(n56948) );
  XNOR U56821 ( .A(p_input[484]), .B(n56947), .Z(n56950) );
  XOR U56822 ( .A(n56947), .B(p_input[452]), .Z(n56949) );
  XOR U56823 ( .A(n56951), .B(n56952), .Z(n56947) );
  AND U56824 ( .A(n56953), .B(n56954), .Z(n56952) );
  XNOR U56825 ( .A(p_input[483]), .B(n56951), .Z(n56954) );
  XOR U56826 ( .A(n56951), .B(p_input[451]), .Z(n56953) );
  XOR U56827 ( .A(n56955), .B(n56956), .Z(n56951) );
  AND U56828 ( .A(n56957), .B(n56958), .Z(n56956) );
  XNOR U56829 ( .A(p_input[482]), .B(n56955), .Z(n56958) );
  XOR U56830 ( .A(n56955), .B(p_input[450]), .Z(n56957) );
  XNOR U56831 ( .A(n56959), .B(n56960), .Z(n56955) );
  AND U56832 ( .A(n56961), .B(n56962), .Z(n56960) );
  XOR U56833 ( .A(p_input[481]), .B(n56959), .Z(n56962) );
  XNOR U56834 ( .A(p_input[449]), .B(n56959), .Z(n56961) );
  AND U56835 ( .A(p_input[480]), .B(n56963), .Z(n56959) );
  IV U56836 ( .A(p_input[448]), .Z(n56963) );
  XNOR U56837 ( .A(p_input[384]), .B(n56964), .Z(n56557) );
  AND U56838 ( .A(n1113), .B(n56965), .Z(n56964) );
  XOR U56839 ( .A(p_input[416]), .B(p_input[384]), .Z(n56965) );
  XOR U56840 ( .A(n56966), .B(n56967), .Z(n1113) );
  AND U56841 ( .A(n56968), .B(n56969), .Z(n56967) );
  XNOR U56842 ( .A(p_input[447]), .B(n56966), .Z(n56969) );
  XOR U56843 ( .A(n56966), .B(p_input[415]), .Z(n56968) );
  XOR U56844 ( .A(n56970), .B(n56971), .Z(n56966) );
  AND U56845 ( .A(n56972), .B(n56973), .Z(n56971) );
  XNOR U56846 ( .A(p_input[446]), .B(n56970), .Z(n56973) );
  XNOR U56847 ( .A(n56970), .B(n56572), .Z(n56972) );
  IV U56848 ( .A(p_input[414]), .Z(n56572) );
  XOR U56849 ( .A(n56974), .B(n56975), .Z(n56970) );
  AND U56850 ( .A(n56976), .B(n56977), .Z(n56975) );
  XNOR U56851 ( .A(p_input[445]), .B(n56974), .Z(n56977) );
  XNOR U56852 ( .A(n56974), .B(n56581), .Z(n56976) );
  IV U56853 ( .A(p_input[413]), .Z(n56581) );
  XOR U56854 ( .A(n56978), .B(n56979), .Z(n56974) );
  AND U56855 ( .A(n56980), .B(n56981), .Z(n56979) );
  XNOR U56856 ( .A(p_input[444]), .B(n56978), .Z(n56981) );
  XNOR U56857 ( .A(n56978), .B(n56590), .Z(n56980) );
  IV U56858 ( .A(p_input[412]), .Z(n56590) );
  XOR U56859 ( .A(n56982), .B(n56983), .Z(n56978) );
  AND U56860 ( .A(n56984), .B(n56985), .Z(n56983) );
  XNOR U56861 ( .A(p_input[443]), .B(n56982), .Z(n56985) );
  XNOR U56862 ( .A(n56982), .B(n56599), .Z(n56984) );
  IV U56863 ( .A(p_input[411]), .Z(n56599) );
  XOR U56864 ( .A(n56986), .B(n56987), .Z(n56982) );
  AND U56865 ( .A(n56988), .B(n56989), .Z(n56987) );
  XNOR U56866 ( .A(p_input[442]), .B(n56986), .Z(n56989) );
  XNOR U56867 ( .A(n56986), .B(n56608), .Z(n56988) );
  IV U56868 ( .A(p_input[410]), .Z(n56608) );
  XOR U56869 ( .A(n56990), .B(n56991), .Z(n56986) );
  AND U56870 ( .A(n56992), .B(n56993), .Z(n56991) );
  XNOR U56871 ( .A(p_input[441]), .B(n56990), .Z(n56993) );
  XNOR U56872 ( .A(n56990), .B(n56617), .Z(n56992) );
  IV U56873 ( .A(p_input[409]), .Z(n56617) );
  XOR U56874 ( .A(n56994), .B(n56995), .Z(n56990) );
  AND U56875 ( .A(n56996), .B(n56997), .Z(n56995) );
  XNOR U56876 ( .A(p_input[440]), .B(n56994), .Z(n56997) );
  XNOR U56877 ( .A(n56994), .B(n56626), .Z(n56996) );
  IV U56878 ( .A(p_input[408]), .Z(n56626) );
  XOR U56879 ( .A(n56998), .B(n56999), .Z(n56994) );
  AND U56880 ( .A(n57000), .B(n57001), .Z(n56999) );
  XNOR U56881 ( .A(p_input[439]), .B(n56998), .Z(n57001) );
  XNOR U56882 ( .A(n56998), .B(n56635), .Z(n57000) );
  IV U56883 ( .A(p_input[407]), .Z(n56635) );
  XOR U56884 ( .A(n57002), .B(n57003), .Z(n56998) );
  AND U56885 ( .A(n57004), .B(n57005), .Z(n57003) );
  XNOR U56886 ( .A(p_input[438]), .B(n57002), .Z(n57005) );
  XNOR U56887 ( .A(n57002), .B(n56644), .Z(n57004) );
  IV U56888 ( .A(p_input[406]), .Z(n56644) );
  XOR U56889 ( .A(n57006), .B(n57007), .Z(n57002) );
  AND U56890 ( .A(n57008), .B(n57009), .Z(n57007) );
  XNOR U56891 ( .A(p_input[437]), .B(n57006), .Z(n57009) );
  XNOR U56892 ( .A(n57006), .B(n56653), .Z(n57008) );
  IV U56893 ( .A(p_input[405]), .Z(n56653) );
  XOR U56894 ( .A(n57010), .B(n57011), .Z(n57006) );
  AND U56895 ( .A(n57012), .B(n57013), .Z(n57011) );
  XNOR U56896 ( .A(p_input[436]), .B(n57010), .Z(n57013) );
  XNOR U56897 ( .A(n57010), .B(n56662), .Z(n57012) );
  IV U56898 ( .A(p_input[404]), .Z(n56662) );
  XOR U56899 ( .A(n57014), .B(n57015), .Z(n57010) );
  AND U56900 ( .A(n57016), .B(n57017), .Z(n57015) );
  XNOR U56901 ( .A(p_input[435]), .B(n57014), .Z(n57017) );
  XNOR U56902 ( .A(n57014), .B(n56671), .Z(n57016) );
  IV U56903 ( .A(p_input[403]), .Z(n56671) );
  XOR U56904 ( .A(n57018), .B(n57019), .Z(n57014) );
  AND U56905 ( .A(n57020), .B(n57021), .Z(n57019) );
  XNOR U56906 ( .A(p_input[434]), .B(n57018), .Z(n57021) );
  XNOR U56907 ( .A(n57018), .B(n56680), .Z(n57020) );
  IV U56908 ( .A(p_input[402]), .Z(n56680) );
  XOR U56909 ( .A(n57022), .B(n57023), .Z(n57018) );
  AND U56910 ( .A(n57024), .B(n57025), .Z(n57023) );
  XNOR U56911 ( .A(p_input[433]), .B(n57022), .Z(n57025) );
  XNOR U56912 ( .A(n57022), .B(n56689), .Z(n57024) );
  IV U56913 ( .A(p_input[401]), .Z(n56689) );
  XOR U56914 ( .A(n57026), .B(n57027), .Z(n57022) );
  AND U56915 ( .A(n57028), .B(n57029), .Z(n57027) );
  XNOR U56916 ( .A(p_input[432]), .B(n57026), .Z(n57029) );
  XNOR U56917 ( .A(n57026), .B(n56698), .Z(n57028) );
  IV U56918 ( .A(p_input[400]), .Z(n56698) );
  XOR U56919 ( .A(n57030), .B(n57031), .Z(n57026) );
  AND U56920 ( .A(n57032), .B(n57033), .Z(n57031) );
  XNOR U56921 ( .A(p_input[431]), .B(n57030), .Z(n57033) );
  XNOR U56922 ( .A(n57030), .B(n56707), .Z(n57032) );
  IV U56923 ( .A(p_input[399]), .Z(n56707) );
  XOR U56924 ( .A(n57034), .B(n57035), .Z(n57030) );
  AND U56925 ( .A(n57036), .B(n57037), .Z(n57035) );
  XNOR U56926 ( .A(p_input[430]), .B(n57034), .Z(n57037) );
  XNOR U56927 ( .A(n57034), .B(n56716), .Z(n57036) );
  IV U56928 ( .A(p_input[398]), .Z(n56716) );
  XOR U56929 ( .A(n57038), .B(n57039), .Z(n57034) );
  AND U56930 ( .A(n57040), .B(n57041), .Z(n57039) );
  XNOR U56931 ( .A(p_input[429]), .B(n57038), .Z(n57041) );
  XNOR U56932 ( .A(n57038), .B(n56725), .Z(n57040) );
  IV U56933 ( .A(p_input[397]), .Z(n56725) );
  XOR U56934 ( .A(n57042), .B(n57043), .Z(n57038) );
  AND U56935 ( .A(n57044), .B(n57045), .Z(n57043) );
  XNOR U56936 ( .A(p_input[428]), .B(n57042), .Z(n57045) );
  XNOR U56937 ( .A(n57042), .B(n56734), .Z(n57044) );
  IV U56938 ( .A(p_input[396]), .Z(n56734) );
  XOR U56939 ( .A(n57046), .B(n57047), .Z(n57042) );
  AND U56940 ( .A(n57048), .B(n57049), .Z(n57047) );
  XNOR U56941 ( .A(p_input[427]), .B(n57046), .Z(n57049) );
  XNOR U56942 ( .A(n57046), .B(n56743), .Z(n57048) );
  IV U56943 ( .A(p_input[395]), .Z(n56743) );
  XOR U56944 ( .A(n57050), .B(n57051), .Z(n57046) );
  AND U56945 ( .A(n57052), .B(n57053), .Z(n57051) );
  XNOR U56946 ( .A(p_input[426]), .B(n57050), .Z(n57053) );
  XNOR U56947 ( .A(n57050), .B(n56752), .Z(n57052) );
  IV U56948 ( .A(p_input[394]), .Z(n56752) );
  XOR U56949 ( .A(n57054), .B(n57055), .Z(n57050) );
  AND U56950 ( .A(n57056), .B(n57057), .Z(n57055) );
  XNOR U56951 ( .A(p_input[425]), .B(n57054), .Z(n57057) );
  XNOR U56952 ( .A(n57054), .B(n56761), .Z(n57056) );
  IV U56953 ( .A(p_input[393]), .Z(n56761) );
  XOR U56954 ( .A(n57058), .B(n57059), .Z(n57054) );
  AND U56955 ( .A(n57060), .B(n57061), .Z(n57059) );
  XNOR U56956 ( .A(p_input[424]), .B(n57058), .Z(n57061) );
  XNOR U56957 ( .A(n57058), .B(n56770), .Z(n57060) );
  IV U56958 ( .A(p_input[392]), .Z(n56770) );
  XOR U56959 ( .A(n57062), .B(n57063), .Z(n57058) );
  AND U56960 ( .A(n57064), .B(n57065), .Z(n57063) );
  XNOR U56961 ( .A(p_input[423]), .B(n57062), .Z(n57065) );
  XNOR U56962 ( .A(n57062), .B(n56779), .Z(n57064) );
  IV U56963 ( .A(p_input[391]), .Z(n56779) );
  XOR U56964 ( .A(n57066), .B(n57067), .Z(n57062) );
  AND U56965 ( .A(n57068), .B(n57069), .Z(n57067) );
  XNOR U56966 ( .A(p_input[422]), .B(n57066), .Z(n57069) );
  XNOR U56967 ( .A(n57066), .B(n56788), .Z(n57068) );
  IV U56968 ( .A(p_input[390]), .Z(n56788) );
  XOR U56969 ( .A(n57070), .B(n57071), .Z(n57066) );
  AND U56970 ( .A(n57072), .B(n57073), .Z(n57071) );
  XNOR U56971 ( .A(p_input[421]), .B(n57070), .Z(n57073) );
  XNOR U56972 ( .A(n57070), .B(n56797), .Z(n57072) );
  IV U56973 ( .A(p_input[389]), .Z(n56797) );
  XOR U56974 ( .A(n57074), .B(n57075), .Z(n57070) );
  AND U56975 ( .A(n57076), .B(n57077), .Z(n57075) );
  XNOR U56976 ( .A(p_input[420]), .B(n57074), .Z(n57077) );
  XNOR U56977 ( .A(n57074), .B(n56806), .Z(n57076) );
  IV U56978 ( .A(p_input[388]), .Z(n56806) );
  XOR U56979 ( .A(n57078), .B(n57079), .Z(n57074) );
  AND U56980 ( .A(n57080), .B(n57081), .Z(n57079) );
  XNOR U56981 ( .A(p_input[419]), .B(n57078), .Z(n57081) );
  XNOR U56982 ( .A(n57078), .B(n56815), .Z(n57080) );
  IV U56983 ( .A(p_input[387]), .Z(n56815) );
  XOR U56984 ( .A(n57082), .B(n57083), .Z(n57078) );
  AND U56985 ( .A(n57084), .B(n57085), .Z(n57083) );
  XNOR U56986 ( .A(p_input[418]), .B(n57082), .Z(n57085) );
  XNOR U56987 ( .A(n57082), .B(n56824), .Z(n57084) );
  IV U56988 ( .A(p_input[386]), .Z(n56824) );
  XNOR U56989 ( .A(n57086), .B(n57087), .Z(n57082) );
  AND U56990 ( .A(n57088), .B(n57089), .Z(n57087) );
  XOR U56991 ( .A(p_input[417]), .B(n57086), .Z(n57089) );
  XNOR U56992 ( .A(p_input[385]), .B(n57086), .Z(n57088) );
  AND U56993 ( .A(p_input[416]), .B(n57090), .Z(n57086) );
  IV U56994 ( .A(p_input[384]), .Z(n57090) );
  XOR U56995 ( .A(n57091), .B(n57092), .Z(n56180) );
  AND U56996 ( .A(n661), .B(n57093), .Z(n57092) );
  XNOR U56997 ( .A(n57094), .B(n57091), .Z(n57093) );
  XOR U56998 ( .A(n57095), .B(n57096), .Z(n661) );
  AND U56999 ( .A(n57097), .B(n57098), .Z(n57096) );
  XNOR U57000 ( .A(n56195), .B(n57095), .Z(n57098) );
  AND U57001 ( .A(p_input[383]), .B(p_input[351]), .Z(n56195) );
  XNOR U57002 ( .A(n57095), .B(n56192), .Z(n57097) );
  IV U57003 ( .A(n57099), .Z(n56192) );
  AND U57004 ( .A(p_input[287]), .B(p_input[319]), .Z(n57099) );
  XOR U57005 ( .A(n57100), .B(n57101), .Z(n57095) );
  AND U57006 ( .A(n57102), .B(n57103), .Z(n57101) );
  XOR U57007 ( .A(n57100), .B(n56207), .Z(n57103) );
  XNOR U57008 ( .A(p_input[350]), .B(n57104), .Z(n56207) );
  AND U57009 ( .A(n1119), .B(n57105), .Z(n57104) );
  XOR U57010 ( .A(p_input[382]), .B(p_input[350]), .Z(n57105) );
  XNOR U57011 ( .A(n56204), .B(n57100), .Z(n57102) );
  XOR U57012 ( .A(n57106), .B(n57107), .Z(n56204) );
  AND U57013 ( .A(n1116), .B(n57108), .Z(n57107) );
  XOR U57014 ( .A(p_input[318]), .B(p_input[286]), .Z(n57108) );
  XOR U57015 ( .A(n57109), .B(n57110), .Z(n57100) );
  AND U57016 ( .A(n57111), .B(n57112), .Z(n57110) );
  XOR U57017 ( .A(n57109), .B(n56219), .Z(n57112) );
  XNOR U57018 ( .A(p_input[349]), .B(n57113), .Z(n56219) );
  AND U57019 ( .A(n1119), .B(n57114), .Z(n57113) );
  XOR U57020 ( .A(p_input[381]), .B(p_input[349]), .Z(n57114) );
  XNOR U57021 ( .A(n56216), .B(n57109), .Z(n57111) );
  XOR U57022 ( .A(n57115), .B(n57116), .Z(n56216) );
  AND U57023 ( .A(n1116), .B(n57117), .Z(n57116) );
  XOR U57024 ( .A(p_input[317]), .B(p_input[285]), .Z(n57117) );
  XOR U57025 ( .A(n57118), .B(n57119), .Z(n57109) );
  AND U57026 ( .A(n57120), .B(n57121), .Z(n57119) );
  XOR U57027 ( .A(n57118), .B(n56231), .Z(n57121) );
  XNOR U57028 ( .A(p_input[348]), .B(n57122), .Z(n56231) );
  AND U57029 ( .A(n1119), .B(n57123), .Z(n57122) );
  XOR U57030 ( .A(p_input[380]), .B(p_input[348]), .Z(n57123) );
  XNOR U57031 ( .A(n56228), .B(n57118), .Z(n57120) );
  XOR U57032 ( .A(n57124), .B(n57125), .Z(n56228) );
  AND U57033 ( .A(n1116), .B(n57126), .Z(n57125) );
  XOR U57034 ( .A(p_input[316]), .B(p_input[284]), .Z(n57126) );
  XOR U57035 ( .A(n57127), .B(n57128), .Z(n57118) );
  AND U57036 ( .A(n57129), .B(n57130), .Z(n57128) );
  XOR U57037 ( .A(n57127), .B(n56243), .Z(n57130) );
  XNOR U57038 ( .A(p_input[347]), .B(n57131), .Z(n56243) );
  AND U57039 ( .A(n1119), .B(n57132), .Z(n57131) );
  XOR U57040 ( .A(p_input[379]), .B(p_input[347]), .Z(n57132) );
  XNOR U57041 ( .A(n56240), .B(n57127), .Z(n57129) );
  XOR U57042 ( .A(n57133), .B(n57134), .Z(n56240) );
  AND U57043 ( .A(n1116), .B(n57135), .Z(n57134) );
  XOR U57044 ( .A(p_input[315]), .B(p_input[283]), .Z(n57135) );
  XOR U57045 ( .A(n57136), .B(n57137), .Z(n57127) );
  AND U57046 ( .A(n57138), .B(n57139), .Z(n57137) );
  XOR U57047 ( .A(n57136), .B(n56255), .Z(n57139) );
  XNOR U57048 ( .A(p_input[346]), .B(n57140), .Z(n56255) );
  AND U57049 ( .A(n1119), .B(n57141), .Z(n57140) );
  XOR U57050 ( .A(p_input[378]), .B(p_input[346]), .Z(n57141) );
  XNOR U57051 ( .A(n56252), .B(n57136), .Z(n57138) );
  XOR U57052 ( .A(n57142), .B(n57143), .Z(n56252) );
  AND U57053 ( .A(n1116), .B(n57144), .Z(n57143) );
  XOR U57054 ( .A(p_input[314]), .B(p_input[282]), .Z(n57144) );
  XOR U57055 ( .A(n57145), .B(n57146), .Z(n57136) );
  AND U57056 ( .A(n57147), .B(n57148), .Z(n57146) );
  XOR U57057 ( .A(n57145), .B(n56267), .Z(n57148) );
  XNOR U57058 ( .A(p_input[345]), .B(n57149), .Z(n56267) );
  AND U57059 ( .A(n1119), .B(n57150), .Z(n57149) );
  XOR U57060 ( .A(p_input[377]), .B(p_input[345]), .Z(n57150) );
  XNOR U57061 ( .A(n56264), .B(n57145), .Z(n57147) );
  XOR U57062 ( .A(n57151), .B(n57152), .Z(n56264) );
  AND U57063 ( .A(n1116), .B(n57153), .Z(n57152) );
  XOR U57064 ( .A(p_input[313]), .B(p_input[281]), .Z(n57153) );
  XOR U57065 ( .A(n57154), .B(n57155), .Z(n57145) );
  AND U57066 ( .A(n57156), .B(n57157), .Z(n57155) );
  XOR U57067 ( .A(n57154), .B(n56279), .Z(n57157) );
  XNOR U57068 ( .A(p_input[344]), .B(n57158), .Z(n56279) );
  AND U57069 ( .A(n1119), .B(n57159), .Z(n57158) );
  XOR U57070 ( .A(p_input[376]), .B(p_input[344]), .Z(n57159) );
  XNOR U57071 ( .A(n56276), .B(n57154), .Z(n57156) );
  XOR U57072 ( .A(n57160), .B(n57161), .Z(n56276) );
  AND U57073 ( .A(n1116), .B(n57162), .Z(n57161) );
  XOR U57074 ( .A(p_input[312]), .B(p_input[280]), .Z(n57162) );
  XOR U57075 ( .A(n57163), .B(n57164), .Z(n57154) );
  AND U57076 ( .A(n57165), .B(n57166), .Z(n57164) );
  XOR U57077 ( .A(n57163), .B(n56291), .Z(n57166) );
  XNOR U57078 ( .A(p_input[343]), .B(n57167), .Z(n56291) );
  AND U57079 ( .A(n1119), .B(n57168), .Z(n57167) );
  XOR U57080 ( .A(p_input[375]), .B(p_input[343]), .Z(n57168) );
  XNOR U57081 ( .A(n56288), .B(n57163), .Z(n57165) );
  XOR U57082 ( .A(n57169), .B(n57170), .Z(n56288) );
  AND U57083 ( .A(n1116), .B(n57171), .Z(n57170) );
  XOR U57084 ( .A(p_input[311]), .B(p_input[279]), .Z(n57171) );
  XOR U57085 ( .A(n57172), .B(n57173), .Z(n57163) );
  AND U57086 ( .A(n57174), .B(n57175), .Z(n57173) );
  XOR U57087 ( .A(n57172), .B(n56303), .Z(n57175) );
  XNOR U57088 ( .A(p_input[342]), .B(n57176), .Z(n56303) );
  AND U57089 ( .A(n1119), .B(n57177), .Z(n57176) );
  XOR U57090 ( .A(p_input[374]), .B(p_input[342]), .Z(n57177) );
  XNOR U57091 ( .A(n56300), .B(n57172), .Z(n57174) );
  XOR U57092 ( .A(n57178), .B(n57179), .Z(n56300) );
  AND U57093 ( .A(n1116), .B(n57180), .Z(n57179) );
  XOR U57094 ( .A(p_input[310]), .B(p_input[278]), .Z(n57180) );
  XOR U57095 ( .A(n57181), .B(n57182), .Z(n57172) );
  AND U57096 ( .A(n57183), .B(n57184), .Z(n57182) );
  XOR U57097 ( .A(n57181), .B(n56315), .Z(n57184) );
  XNOR U57098 ( .A(p_input[341]), .B(n57185), .Z(n56315) );
  AND U57099 ( .A(n1119), .B(n57186), .Z(n57185) );
  XOR U57100 ( .A(p_input[373]), .B(p_input[341]), .Z(n57186) );
  XNOR U57101 ( .A(n56312), .B(n57181), .Z(n57183) );
  XOR U57102 ( .A(n57187), .B(n57188), .Z(n56312) );
  AND U57103 ( .A(n1116), .B(n57189), .Z(n57188) );
  XOR U57104 ( .A(p_input[309]), .B(p_input[277]), .Z(n57189) );
  XOR U57105 ( .A(n57190), .B(n57191), .Z(n57181) );
  AND U57106 ( .A(n57192), .B(n57193), .Z(n57191) );
  XOR U57107 ( .A(n57190), .B(n56327), .Z(n57193) );
  XNOR U57108 ( .A(p_input[340]), .B(n57194), .Z(n56327) );
  AND U57109 ( .A(n1119), .B(n57195), .Z(n57194) );
  XOR U57110 ( .A(p_input[372]), .B(p_input[340]), .Z(n57195) );
  XNOR U57111 ( .A(n56324), .B(n57190), .Z(n57192) );
  XOR U57112 ( .A(n57196), .B(n57197), .Z(n56324) );
  AND U57113 ( .A(n1116), .B(n57198), .Z(n57197) );
  XOR U57114 ( .A(p_input[308]), .B(p_input[276]), .Z(n57198) );
  XOR U57115 ( .A(n57199), .B(n57200), .Z(n57190) );
  AND U57116 ( .A(n57201), .B(n57202), .Z(n57200) );
  XOR U57117 ( .A(n57199), .B(n56339), .Z(n57202) );
  XNOR U57118 ( .A(p_input[339]), .B(n57203), .Z(n56339) );
  AND U57119 ( .A(n1119), .B(n57204), .Z(n57203) );
  XOR U57120 ( .A(p_input[371]), .B(p_input[339]), .Z(n57204) );
  XNOR U57121 ( .A(n56336), .B(n57199), .Z(n57201) );
  XOR U57122 ( .A(n57205), .B(n57206), .Z(n56336) );
  AND U57123 ( .A(n1116), .B(n57207), .Z(n57206) );
  XOR U57124 ( .A(p_input[307]), .B(p_input[275]), .Z(n57207) );
  XOR U57125 ( .A(n57208), .B(n57209), .Z(n57199) );
  AND U57126 ( .A(n57210), .B(n57211), .Z(n57209) );
  XOR U57127 ( .A(n57208), .B(n56351), .Z(n57211) );
  XNOR U57128 ( .A(p_input[338]), .B(n57212), .Z(n56351) );
  AND U57129 ( .A(n1119), .B(n57213), .Z(n57212) );
  XOR U57130 ( .A(p_input[370]), .B(p_input[338]), .Z(n57213) );
  XNOR U57131 ( .A(n56348), .B(n57208), .Z(n57210) );
  XOR U57132 ( .A(n57214), .B(n57215), .Z(n56348) );
  AND U57133 ( .A(n1116), .B(n57216), .Z(n57215) );
  XOR U57134 ( .A(p_input[306]), .B(p_input[274]), .Z(n57216) );
  XOR U57135 ( .A(n57217), .B(n57218), .Z(n57208) );
  AND U57136 ( .A(n57219), .B(n57220), .Z(n57218) );
  XOR U57137 ( .A(n57217), .B(n56363), .Z(n57220) );
  XNOR U57138 ( .A(p_input[337]), .B(n57221), .Z(n56363) );
  AND U57139 ( .A(n1119), .B(n57222), .Z(n57221) );
  XOR U57140 ( .A(p_input[369]), .B(p_input[337]), .Z(n57222) );
  XNOR U57141 ( .A(n56360), .B(n57217), .Z(n57219) );
  XOR U57142 ( .A(n57223), .B(n57224), .Z(n56360) );
  AND U57143 ( .A(n1116), .B(n57225), .Z(n57224) );
  XOR U57144 ( .A(p_input[305]), .B(p_input[273]), .Z(n57225) );
  XOR U57145 ( .A(n57226), .B(n57227), .Z(n57217) );
  AND U57146 ( .A(n57228), .B(n57229), .Z(n57227) );
  XOR U57147 ( .A(n57226), .B(n56375), .Z(n57229) );
  XNOR U57148 ( .A(p_input[336]), .B(n57230), .Z(n56375) );
  AND U57149 ( .A(n1119), .B(n57231), .Z(n57230) );
  XOR U57150 ( .A(p_input[368]), .B(p_input[336]), .Z(n57231) );
  XNOR U57151 ( .A(n56372), .B(n57226), .Z(n57228) );
  XOR U57152 ( .A(n57232), .B(n57233), .Z(n56372) );
  AND U57153 ( .A(n1116), .B(n57234), .Z(n57233) );
  XOR U57154 ( .A(p_input[304]), .B(p_input[272]), .Z(n57234) );
  XOR U57155 ( .A(n57235), .B(n57236), .Z(n57226) );
  AND U57156 ( .A(n57237), .B(n57238), .Z(n57236) );
  XOR U57157 ( .A(n57235), .B(n56387), .Z(n57238) );
  XNOR U57158 ( .A(p_input[335]), .B(n57239), .Z(n56387) );
  AND U57159 ( .A(n1119), .B(n57240), .Z(n57239) );
  XOR U57160 ( .A(p_input[367]), .B(p_input[335]), .Z(n57240) );
  XNOR U57161 ( .A(n56384), .B(n57235), .Z(n57237) );
  XOR U57162 ( .A(n57241), .B(n57242), .Z(n56384) );
  AND U57163 ( .A(n1116), .B(n57243), .Z(n57242) );
  XOR U57164 ( .A(p_input[303]), .B(p_input[271]), .Z(n57243) );
  XOR U57165 ( .A(n57244), .B(n57245), .Z(n57235) );
  AND U57166 ( .A(n57246), .B(n57247), .Z(n57245) );
  XOR U57167 ( .A(n57244), .B(n56399), .Z(n57247) );
  XNOR U57168 ( .A(p_input[334]), .B(n57248), .Z(n56399) );
  AND U57169 ( .A(n1119), .B(n57249), .Z(n57248) );
  XOR U57170 ( .A(p_input[366]), .B(p_input[334]), .Z(n57249) );
  XNOR U57171 ( .A(n56396), .B(n57244), .Z(n57246) );
  XOR U57172 ( .A(n57250), .B(n57251), .Z(n56396) );
  AND U57173 ( .A(n1116), .B(n57252), .Z(n57251) );
  XOR U57174 ( .A(p_input[302]), .B(p_input[270]), .Z(n57252) );
  XOR U57175 ( .A(n57253), .B(n57254), .Z(n57244) );
  AND U57176 ( .A(n57255), .B(n57256), .Z(n57254) );
  XOR U57177 ( .A(n57253), .B(n56411), .Z(n57256) );
  XNOR U57178 ( .A(p_input[333]), .B(n57257), .Z(n56411) );
  AND U57179 ( .A(n1119), .B(n57258), .Z(n57257) );
  XOR U57180 ( .A(p_input[365]), .B(p_input[333]), .Z(n57258) );
  XNOR U57181 ( .A(n56408), .B(n57253), .Z(n57255) );
  XOR U57182 ( .A(n57259), .B(n57260), .Z(n56408) );
  AND U57183 ( .A(n1116), .B(n57261), .Z(n57260) );
  XOR U57184 ( .A(p_input[301]), .B(p_input[269]), .Z(n57261) );
  XOR U57185 ( .A(n57262), .B(n57263), .Z(n57253) );
  AND U57186 ( .A(n57264), .B(n57265), .Z(n57263) );
  XOR U57187 ( .A(n57262), .B(n56423), .Z(n57265) );
  XNOR U57188 ( .A(p_input[332]), .B(n57266), .Z(n56423) );
  AND U57189 ( .A(n1119), .B(n57267), .Z(n57266) );
  XOR U57190 ( .A(p_input[364]), .B(p_input[332]), .Z(n57267) );
  XNOR U57191 ( .A(n56420), .B(n57262), .Z(n57264) );
  XOR U57192 ( .A(n57268), .B(n57269), .Z(n56420) );
  AND U57193 ( .A(n1116), .B(n57270), .Z(n57269) );
  XOR U57194 ( .A(p_input[300]), .B(p_input[268]), .Z(n57270) );
  XOR U57195 ( .A(n57271), .B(n57272), .Z(n57262) );
  AND U57196 ( .A(n57273), .B(n57274), .Z(n57272) );
  XOR U57197 ( .A(n57271), .B(n56435), .Z(n57274) );
  XNOR U57198 ( .A(p_input[331]), .B(n57275), .Z(n56435) );
  AND U57199 ( .A(n1119), .B(n57276), .Z(n57275) );
  XOR U57200 ( .A(p_input[363]), .B(p_input[331]), .Z(n57276) );
  XNOR U57201 ( .A(n56432), .B(n57271), .Z(n57273) );
  XOR U57202 ( .A(n57277), .B(n57278), .Z(n56432) );
  AND U57203 ( .A(n1116), .B(n57279), .Z(n57278) );
  XOR U57204 ( .A(p_input[299]), .B(p_input[267]), .Z(n57279) );
  XOR U57205 ( .A(n57280), .B(n57281), .Z(n57271) );
  AND U57206 ( .A(n57282), .B(n57283), .Z(n57281) );
  XOR U57207 ( .A(n57280), .B(n56447), .Z(n57283) );
  XNOR U57208 ( .A(p_input[330]), .B(n57284), .Z(n56447) );
  AND U57209 ( .A(n1119), .B(n57285), .Z(n57284) );
  XOR U57210 ( .A(p_input[362]), .B(p_input[330]), .Z(n57285) );
  XNOR U57211 ( .A(n56444), .B(n57280), .Z(n57282) );
  XOR U57212 ( .A(n57286), .B(n57287), .Z(n56444) );
  AND U57213 ( .A(n1116), .B(n57288), .Z(n57287) );
  XOR U57214 ( .A(p_input[298]), .B(p_input[266]), .Z(n57288) );
  XOR U57215 ( .A(n57289), .B(n57290), .Z(n57280) );
  AND U57216 ( .A(n57291), .B(n57292), .Z(n57290) );
  XOR U57217 ( .A(n57289), .B(n56459), .Z(n57292) );
  XNOR U57218 ( .A(p_input[329]), .B(n57293), .Z(n56459) );
  AND U57219 ( .A(n1119), .B(n57294), .Z(n57293) );
  XOR U57220 ( .A(p_input[361]), .B(p_input[329]), .Z(n57294) );
  XNOR U57221 ( .A(n56456), .B(n57289), .Z(n57291) );
  XOR U57222 ( .A(n57295), .B(n57296), .Z(n56456) );
  AND U57223 ( .A(n1116), .B(n57297), .Z(n57296) );
  XOR U57224 ( .A(p_input[297]), .B(p_input[265]), .Z(n57297) );
  XOR U57225 ( .A(n57298), .B(n57299), .Z(n57289) );
  AND U57226 ( .A(n57300), .B(n57301), .Z(n57299) );
  XOR U57227 ( .A(n57298), .B(n56471), .Z(n57301) );
  XNOR U57228 ( .A(p_input[328]), .B(n57302), .Z(n56471) );
  AND U57229 ( .A(n1119), .B(n57303), .Z(n57302) );
  XOR U57230 ( .A(p_input[360]), .B(p_input[328]), .Z(n57303) );
  XNOR U57231 ( .A(n56468), .B(n57298), .Z(n57300) );
  XOR U57232 ( .A(n57304), .B(n57305), .Z(n56468) );
  AND U57233 ( .A(n1116), .B(n57306), .Z(n57305) );
  XOR U57234 ( .A(p_input[296]), .B(p_input[264]), .Z(n57306) );
  XOR U57235 ( .A(n57307), .B(n57308), .Z(n57298) );
  AND U57236 ( .A(n57309), .B(n57310), .Z(n57308) );
  XOR U57237 ( .A(n57307), .B(n56483), .Z(n57310) );
  XNOR U57238 ( .A(p_input[327]), .B(n57311), .Z(n56483) );
  AND U57239 ( .A(n1119), .B(n57312), .Z(n57311) );
  XOR U57240 ( .A(p_input[359]), .B(p_input[327]), .Z(n57312) );
  XNOR U57241 ( .A(n56480), .B(n57307), .Z(n57309) );
  XOR U57242 ( .A(n57313), .B(n57314), .Z(n56480) );
  AND U57243 ( .A(n1116), .B(n57315), .Z(n57314) );
  XOR U57244 ( .A(p_input[295]), .B(p_input[263]), .Z(n57315) );
  XOR U57245 ( .A(n57316), .B(n57317), .Z(n57307) );
  AND U57246 ( .A(n57318), .B(n57319), .Z(n57317) );
  XOR U57247 ( .A(n57316), .B(n56495), .Z(n57319) );
  XNOR U57248 ( .A(p_input[326]), .B(n57320), .Z(n56495) );
  AND U57249 ( .A(n1119), .B(n57321), .Z(n57320) );
  XOR U57250 ( .A(p_input[358]), .B(p_input[326]), .Z(n57321) );
  XNOR U57251 ( .A(n56492), .B(n57316), .Z(n57318) );
  XOR U57252 ( .A(n57322), .B(n57323), .Z(n56492) );
  AND U57253 ( .A(n1116), .B(n57324), .Z(n57323) );
  XOR U57254 ( .A(p_input[294]), .B(p_input[262]), .Z(n57324) );
  XOR U57255 ( .A(n57325), .B(n57326), .Z(n57316) );
  AND U57256 ( .A(n57327), .B(n57328), .Z(n57326) );
  XOR U57257 ( .A(n57325), .B(n56507), .Z(n57328) );
  XNOR U57258 ( .A(p_input[325]), .B(n57329), .Z(n56507) );
  AND U57259 ( .A(n1119), .B(n57330), .Z(n57329) );
  XOR U57260 ( .A(p_input[357]), .B(p_input[325]), .Z(n57330) );
  XNOR U57261 ( .A(n56504), .B(n57325), .Z(n57327) );
  XOR U57262 ( .A(n57331), .B(n57332), .Z(n56504) );
  AND U57263 ( .A(n1116), .B(n57333), .Z(n57332) );
  XOR U57264 ( .A(p_input[293]), .B(p_input[261]), .Z(n57333) );
  XOR U57265 ( .A(n57334), .B(n57335), .Z(n57325) );
  AND U57266 ( .A(n57336), .B(n57337), .Z(n57335) );
  XOR U57267 ( .A(n57334), .B(n56519), .Z(n57337) );
  XNOR U57268 ( .A(p_input[324]), .B(n57338), .Z(n56519) );
  AND U57269 ( .A(n1119), .B(n57339), .Z(n57338) );
  XOR U57270 ( .A(p_input[356]), .B(p_input[324]), .Z(n57339) );
  XNOR U57271 ( .A(n56516), .B(n57334), .Z(n57336) );
  XOR U57272 ( .A(n57340), .B(n57341), .Z(n56516) );
  AND U57273 ( .A(n1116), .B(n57342), .Z(n57341) );
  XOR U57274 ( .A(p_input[292]), .B(p_input[260]), .Z(n57342) );
  XOR U57275 ( .A(n57343), .B(n57344), .Z(n57334) );
  AND U57276 ( .A(n57345), .B(n57346), .Z(n57344) );
  XOR U57277 ( .A(n57343), .B(n56531), .Z(n57346) );
  XNOR U57278 ( .A(p_input[323]), .B(n57347), .Z(n56531) );
  AND U57279 ( .A(n1119), .B(n57348), .Z(n57347) );
  XOR U57280 ( .A(p_input[355]), .B(p_input[323]), .Z(n57348) );
  XNOR U57281 ( .A(n56528), .B(n57343), .Z(n57345) );
  XOR U57282 ( .A(n57349), .B(n57350), .Z(n56528) );
  AND U57283 ( .A(n1116), .B(n57351), .Z(n57350) );
  XOR U57284 ( .A(p_input[291]), .B(p_input[259]), .Z(n57351) );
  XOR U57285 ( .A(n57352), .B(n57353), .Z(n57343) );
  AND U57286 ( .A(n57354), .B(n57355), .Z(n57353) );
  XOR U57287 ( .A(n57352), .B(n56543), .Z(n57355) );
  XNOR U57288 ( .A(p_input[322]), .B(n57356), .Z(n56543) );
  AND U57289 ( .A(n1119), .B(n57357), .Z(n57356) );
  XOR U57290 ( .A(p_input[354]), .B(p_input[322]), .Z(n57357) );
  XNOR U57291 ( .A(n56540), .B(n57352), .Z(n57354) );
  XOR U57292 ( .A(n57358), .B(n57359), .Z(n56540) );
  AND U57293 ( .A(n1116), .B(n57360), .Z(n57359) );
  XOR U57294 ( .A(p_input[290]), .B(p_input[258]), .Z(n57360) );
  XOR U57295 ( .A(n57361), .B(n57362), .Z(n57352) );
  AND U57296 ( .A(n57363), .B(n57364), .Z(n57362) );
  XNOR U57297 ( .A(n57365), .B(n56556), .Z(n57364) );
  XNOR U57298 ( .A(p_input[321]), .B(n57366), .Z(n56556) );
  AND U57299 ( .A(n1119), .B(n57367), .Z(n57366) );
  XNOR U57300 ( .A(p_input[353]), .B(n57368), .Z(n57367) );
  IV U57301 ( .A(p_input[321]), .Z(n57368) );
  XNOR U57302 ( .A(n56553), .B(n57361), .Z(n57363) );
  XNOR U57303 ( .A(p_input[257]), .B(n57369), .Z(n56553) );
  AND U57304 ( .A(n1116), .B(n57370), .Z(n57369) );
  XOR U57305 ( .A(p_input[289]), .B(p_input[257]), .Z(n57370) );
  IV U57306 ( .A(n57365), .Z(n57361) );
  AND U57307 ( .A(n57091), .B(n57094), .Z(n57365) );
  XOR U57308 ( .A(p_input[320]), .B(n57371), .Z(n57094) );
  AND U57309 ( .A(n1119), .B(n57372), .Z(n57371) );
  XOR U57310 ( .A(p_input[352]), .B(p_input[320]), .Z(n57372) );
  XOR U57311 ( .A(n57373), .B(n57374), .Z(n1119) );
  AND U57312 ( .A(n57375), .B(n57376), .Z(n57374) );
  XNOR U57313 ( .A(p_input[383]), .B(n57373), .Z(n57376) );
  XOR U57314 ( .A(n57373), .B(p_input[351]), .Z(n57375) );
  XOR U57315 ( .A(n57377), .B(n57378), .Z(n57373) );
  AND U57316 ( .A(n57379), .B(n57380), .Z(n57378) );
  XNOR U57317 ( .A(p_input[382]), .B(n57377), .Z(n57380) );
  XOR U57318 ( .A(n57377), .B(p_input[350]), .Z(n57379) );
  XOR U57319 ( .A(n57381), .B(n57382), .Z(n57377) );
  AND U57320 ( .A(n57383), .B(n57384), .Z(n57382) );
  XNOR U57321 ( .A(p_input[381]), .B(n57381), .Z(n57384) );
  XOR U57322 ( .A(n57381), .B(p_input[349]), .Z(n57383) );
  XOR U57323 ( .A(n57385), .B(n57386), .Z(n57381) );
  AND U57324 ( .A(n57387), .B(n57388), .Z(n57386) );
  XNOR U57325 ( .A(p_input[380]), .B(n57385), .Z(n57388) );
  XOR U57326 ( .A(n57385), .B(p_input[348]), .Z(n57387) );
  XOR U57327 ( .A(n57389), .B(n57390), .Z(n57385) );
  AND U57328 ( .A(n57391), .B(n57392), .Z(n57390) );
  XNOR U57329 ( .A(p_input[379]), .B(n57389), .Z(n57392) );
  XOR U57330 ( .A(n57389), .B(p_input[347]), .Z(n57391) );
  XOR U57331 ( .A(n57393), .B(n57394), .Z(n57389) );
  AND U57332 ( .A(n57395), .B(n57396), .Z(n57394) );
  XNOR U57333 ( .A(p_input[378]), .B(n57393), .Z(n57396) );
  XOR U57334 ( .A(n57393), .B(p_input[346]), .Z(n57395) );
  XOR U57335 ( .A(n57397), .B(n57398), .Z(n57393) );
  AND U57336 ( .A(n57399), .B(n57400), .Z(n57398) );
  XNOR U57337 ( .A(p_input[377]), .B(n57397), .Z(n57400) );
  XOR U57338 ( .A(n57397), .B(p_input[345]), .Z(n57399) );
  XOR U57339 ( .A(n57401), .B(n57402), .Z(n57397) );
  AND U57340 ( .A(n57403), .B(n57404), .Z(n57402) );
  XNOR U57341 ( .A(p_input[376]), .B(n57401), .Z(n57404) );
  XOR U57342 ( .A(n57401), .B(p_input[344]), .Z(n57403) );
  XOR U57343 ( .A(n57405), .B(n57406), .Z(n57401) );
  AND U57344 ( .A(n57407), .B(n57408), .Z(n57406) );
  XNOR U57345 ( .A(p_input[375]), .B(n57405), .Z(n57408) );
  XOR U57346 ( .A(n57405), .B(p_input[343]), .Z(n57407) );
  XOR U57347 ( .A(n57409), .B(n57410), .Z(n57405) );
  AND U57348 ( .A(n57411), .B(n57412), .Z(n57410) );
  XNOR U57349 ( .A(p_input[374]), .B(n57409), .Z(n57412) );
  XOR U57350 ( .A(n57409), .B(p_input[342]), .Z(n57411) );
  XOR U57351 ( .A(n57413), .B(n57414), .Z(n57409) );
  AND U57352 ( .A(n57415), .B(n57416), .Z(n57414) );
  XNOR U57353 ( .A(p_input[373]), .B(n57413), .Z(n57416) );
  XOR U57354 ( .A(n57413), .B(p_input[341]), .Z(n57415) );
  XOR U57355 ( .A(n57417), .B(n57418), .Z(n57413) );
  AND U57356 ( .A(n57419), .B(n57420), .Z(n57418) );
  XNOR U57357 ( .A(p_input[372]), .B(n57417), .Z(n57420) );
  XOR U57358 ( .A(n57417), .B(p_input[340]), .Z(n57419) );
  XOR U57359 ( .A(n57421), .B(n57422), .Z(n57417) );
  AND U57360 ( .A(n57423), .B(n57424), .Z(n57422) );
  XNOR U57361 ( .A(p_input[371]), .B(n57421), .Z(n57424) );
  XOR U57362 ( .A(n57421), .B(p_input[339]), .Z(n57423) );
  XOR U57363 ( .A(n57425), .B(n57426), .Z(n57421) );
  AND U57364 ( .A(n57427), .B(n57428), .Z(n57426) );
  XNOR U57365 ( .A(p_input[370]), .B(n57425), .Z(n57428) );
  XOR U57366 ( .A(n57425), .B(p_input[338]), .Z(n57427) );
  XOR U57367 ( .A(n57429), .B(n57430), .Z(n57425) );
  AND U57368 ( .A(n57431), .B(n57432), .Z(n57430) );
  XNOR U57369 ( .A(p_input[369]), .B(n57429), .Z(n57432) );
  XOR U57370 ( .A(n57429), .B(p_input[337]), .Z(n57431) );
  XOR U57371 ( .A(n57433), .B(n57434), .Z(n57429) );
  AND U57372 ( .A(n57435), .B(n57436), .Z(n57434) );
  XNOR U57373 ( .A(p_input[368]), .B(n57433), .Z(n57436) );
  XOR U57374 ( .A(n57433), .B(p_input[336]), .Z(n57435) );
  XOR U57375 ( .A(n57437), .B(n57438), .Z(n57433) );
  AND U57376 ( .A(n57439), .B(n57440), .Z(n57438) );
  XNOR U57377 ( .A(p_input[367]), .B(n57437), .Z(n57440) );
  XOR U57378 ( .A(n57437), .B(p_input[335]), .Z(n57439) );
  XOR U57379 ( .A(n57441), .B(n57442), .Z(n57437) );
  AND U57380 ( .A(n57443), .B(n57444), .Z(n57442) );
  XNOR U57381 ( .A(p_input[366]), .B(n57441), .Z(n57444) );
  XOR U57382 ( .A(n57441), .B(p_input[334]), .Z(n57443) );
  XOR U57383 ( .A(n57445), .B(n57446), .Z(n57441) );
  AND U57384 ( .A(n57447), .B(n57448), .Z(n57446) );
  XNOR U57385 ( .A(p_input[365]), .B(n57445), .Z(n57448) );
  XOR U57386 ( .A(n57445), .B(p_input[333]), .Z(n57447) );
  XOR U57387 ( .A(n57449), .B(n57450), .Z(n57445) );
  AND U57388 ( .A(n57451), .B(n57452), .Z(n57450) );
  XNOR U57389 ( .A(p_input[364]), .B(n57449), .Z(n57452) );
  XOR U57390 ( .A(n57449), .B(p_input[332]), .Z(n57451) );
  XOR U57391 ( .A(n57453), .B(n57454), .Z(n57449) );
  AND U57392 ( .A(n57455), .B(n57456), .Z(n57454) );
  XNOR U57393 ( .A(p_input[363]), .B(n57453), .Z(n57456) );
  XOR U57394 ( .A(n57453), .B(p_input[331]), .Z(n57455) );
  XOR U57395 ( .A(n57457), .B(n57458), .Z(n57453) );
  AND U57396 ( .A(n57459), .B(n57460), .Z(n57458) );
  XNOR U57397 ( .A(p_input[362]), .B(n57457), .Z(n57460) );
  XOR U57398 ( .A(n57457), .B(p_input[330]), .Z(n57459) );
  XOR U57399 ( .A(n57461), .B(n57462), .Z(n57457) );
  AND U57400 ( .A(n57463), .B(n57464), .Z(n57462) );
  XNOR U57401 ( .A(p_input[361]), .B(n57461), .Z(n57464) );
  XOR U57402 ( .A(n57461), .B(p_input[329]), .Z(n57463) );
  XOR U57403 ( .A(n57465), .B(n57466), .Z(n57461) );
  AND U57404 ( .A(n57467), .B(n57468), .Z(n57466) );
  XNOR U57405 ( .A(p_input[360]), .B(n57465), .Z(n57468) );
  XOR U57406 ( .A(n57465), .B(p_input[328]), .Z(n57467) );
  XOR U57407 ( .A(n57469), .B(n57470), .Z(n57465) );
  AND U57408 ( .A(n57471), .B(n57472), .Z(n57470) );
  XNOR U57409 ( .A(p_input[359]), .B(n57469), .Z(n57472) );
  XOR U57410 ( .A(n57469), .B(p_input[327]), .Z(n57471) );
  XOR U57411 ( .A(n57473), .B(n57474), .Z(n57469) );
  AND U57412 ( .A(n57475), .B(n57476), .Z(n57474) );
  XNOR U57413 ( .A(p_input[358]), .B(n57473), .Z(n57476) );
  XOR U57414 ( .A(n57473), .B(p_input[326]), .Z(n57475) );
  XOR U57415 ( .A(n57477), .B(n57478), .Z(n57473) );
  AND U57416 ( .A(n57479), .B(n57480), .Z(n57478) );
  XNOR U57417 ( .A(p_input[357]), .B(n57477), .Z(n57480) );
  XOR U57418 ( .A(n57477), .B(p_input[325]), .Z(n57479) );
  XOR U57419 ( .A(n57481), .B(n57482), .Z(n57477) );
  AND U57420 ( .A(n57483), .B(n57484), .Z(n57482) );
  XNOR U57421 ( .A(p_input[356]), .B(n57481), .Z(n57484) );
  XOR U57422 ( .A(n57481), .B(p_input[324]), .Z(n57483) );
  XOR U57423 ( .A(n57485), .B(n57486), .Z(n57481) );
  AND U57424 ( .A(n57487), .B(n57488), .Z(n57486) );
  XNOR U57425 ( .A(p_input[355]), .B(n57485), .Z(n57488) );
  XOR U57426 ( .A(n57485), .B(p_input[323]), .Z(n57487) );
  XOR U57427 ( .A(n57489), .B(n57490), .Z(n57485) );
  AND U57428 ( .A(n57491), .B(n57492), .Z(n57490) );
  XNOR U57429 ( .A(p_input[354]), .B(n57489), .Z(n57492) );
  XOR U57430 ( .A(n57489), .B(p_input[322]), .Z(n57491) );
  XNOR U57431 ( .A(n57493), .B(n57494), .Z(n57489) );
  AND U57432 ( .A(n57495), .B(n57496), .Z(n57494) );
  XOR U57433 ( .A(p_input[353]), .B(n57493), .Z(n57496) );
  XNOR U57434 ( .A(p_input[321]), .B(n57493), .Z(n57495) );
  AND U57435 ( .A(p_input[352]), .B(n57497), .Z(n57493) );
  IV U57436 ( .A(p_input[320]), .Z(n57497) );
  XNOR U57437 ( .A(p_input[256]), .B(n57498), .Z(n57091) );
  AND U57438 ( .A(n1116), .B(n57499), .Z(n57498) );
  XOR U57439 ( .A(p_input[288]), .B(p_input[256]), .Z(n57499) );
  XOR U57440 ( .A(n57500), .B(n57501), .Z(n1116) );
  AND U57441 ( .A(n57502), .B(n57503), .Z(n57501) );
  XNOR U57442 ( .A(p_input[319]), .B(n57500), .Z(n57503) );
  XOR U57443 ( .A(n57500), .B(p_input[287]), .Z(n57502) );
  XOR U57444 ( .A(n57504), .B(n57505), .Z(n57500) );
  AND U57445 ( .A(n57506), .B(n57507), .Z(n57505) );
  XNOR U57446 ( .A(p_input[318]), .B(n57504), .Z(n57507) );
  XNOR U57447 ( .A(n57504), .B(n57106), .Z(n57506) );
  IV U57448 ( .A(p_input[286]), .Z(n57106) );
  XOR U57449 ( .A(n57508), .B(n57509), .Z(n57504) );
  AND U57450 ( .A(n57510), .B(n57511), .Z(n57509) );
  XNOR U57451 ( .A(p_input[317]), .B(n57508), .Z(n57511) );
  XNOR U57452 ( .A(n57508), .B(n57115), .Z(n57510) );
  IV U57453 ( .A(p_input[285]), .Z(n57115) );
  XOR U57454 ( .A(n57512), .B(n57513), .Z(n57508) );
  AND U57455 ( .A(n57514), .B(n57515), .Z(n57513) );
  XNOR U57456 ( .A(p_input[316]), .B(n57512), .Z(n57515) );
  XNOR U57457 ( .A(n57512), .B(n57124), .Z(n57514) );
  IV U57458 ( .A(p_input[284]), .Z(n57124) );
  XOR U57459 ( .A(n57516), .B(n57517), .Z(n57512) );
  AND U57460 ( .A(n57518), .B(n57519), .Z(n57517) );
  XNOR U57461 ( .A(p_input[315]), .B(n57516), .Z(n57519) );
  XNOR U57462 ( .A(n57516), .B(n57133), .Z(n57518) );
  IV U57463 ( .A(p_input[283]), .Z(n57133) );
  XOR U57464 ( .A(n57520), .B(n57521), .Z(n57516) );
  AND U57465 ( .A(n57522), .B(n57523), .Z(n57521) );
  XNOR U57466 ( .A(p_input[314]), .B(n57520), .Z(n57523) );
  XNOR U57467 ( .A(n57520), .B(n57142), .Z(n57522) );
  IV U57468 ( .A(p_input[282]), .Z(n57142) );
  XOR U57469 ( .A(n57524), .B(n57525), .Z(n57520) );
  AND U57470 ( .A(n57526), .B(n57527), .Z(n57525) );
  XNOR U57471 ( .A(p_input[313]), .B(n57524), .Z(n57527) );
  XNOR U57472 ( .A(n57524), .B(n57151), .Z(n57526) );
  IV U57473 ( .A(p_input[281]), .Z(n57151) );
  XOR U57474 ( .A(n57528), .B(n57529), .Z(n57524) );
  AND U57475 ( .A(n57530), .B(n57531), .Z(n57529) );
  XNOR U57476 ( .A(p_input[312]), .B(n57528), .Z(n57531) );
  XNOR U57477 ( .A(n57528), .B(n57160), .Z(n57530) );
  IV U57478 ( .A(p_input[280]), .Z(n57160) );
  XOR U57479 ( .A(n57532), .B(n57533), .Z(n57528) );
  AND U57480 ( .A(n57534), .B(n57535), .Z(n57533) );
  XNOR U57481 ( .A(p_input[311]), .B(n57532), .Z(n57535) );
  XNOR U57482 ( .A(n57532), .B(n57169), .Z(n57534) );
  IV U57483 ( .A(p_input[279]), .Z(n57169) );
  XOR U57484 ( .A(n57536), .B(n57537), .Z(n57532) );
  AND U57485 ( .A(n57538), .B(n57539), .Z(n57537) );
  XNOR U57486 ( .A(p_input[310]), .B(n57536), .Z(n57539) );
  XNOR U57487 ( .A(n57536), .B(n57178), .Z(n57538) );
  IV U57488 ( .A(p_input[278]), .Z(n57178) );
  XOR U57489 ( .A(n57540), .B(n57541), .Z(n57536) );
  AND U57490 ( .A(n57542), .B(n57543), .Z(n57541) );
  XNOR U57491 ( .A(p_input[309]), .B(n57540), .Z(n57543) );
  XNOR U57492 ( .A(n57540), .B(n57187), .Z(n57542) );
  IV U57493 ( .A(p_input[277]), .Z(n57187) );
  XOR U57494 ( .A(n57544), .B(n57545), .Z(n57540) );
  AND U57495 ( .A(n57546), .B(n57547), .Z(n57545) );
  XNOR U57496 ( .A(p_input[308]), .B(n57544), .Z(n57547) );
  XNOR U57497 ( .A(n57544), .B(n57196), .Z(n57546) );
  IV U57498 ( .A(p_input[276]), .Z(n57196) );
  XOR U57499 ( .A(n57548), .B(n57549), .Z(n57544) );
  AND U57500 ( .A(n57550), .B(n57551), .Z(n57549) );
  XNOR U57501 ( .A(p_input[307]), .B(n57548), .Z(n57551) );
  XNOR U57502 ( .A(n57548), .B(n57205), .Z(n57550) );
  IV U57503 ( .A(p_input[275]), .Z(n57205) );
  XOR U57504 ( .A(n57552), .B(n57553), .Z(n57548) );
  AND U57505 ( .A(n57554), .B(n57555), .Z(n57553) );
  XNOR U57506 ( .A(p_input[306]), .B(n57552), .Z(n57555) );
  XNOR U57507 ( .A(n57552), .B(n57214), .Z(n57554) );
  IV U57508 ( .A(p_input[274]), .Z(n57214) );
  XOR U57509 ( .A(n57556), .B(n57557), .Z(n57552) );
  AND U57510 ( .A(n57558), .B(n57559), .Z(n57557) );
  XNOR U57511 ( .A(p_input[305]), .B(n57556), .Z(n57559) );
  XNOR U57512 ( .A(n57556), .B(n57223), .Z(n57558) );
  IV U57513 ( .A(p_input[273]), .Z(n57223) );
  XOR U57514 ( .A(n57560), .B(n57561), .Z(n57556) );
  AND U57515 ( .A(n57562), .B(n57563), .Z(n57561) );
  XNOR U57516 ( .A(p_input[304]), .B(n57560), .Z(n57563) );
  XNOR U57517 ( .A(n57560), .B(n57232), .Z(n57562) );
  IV U57518 ( .A(p_input[272]), .Z(n57232) );
  XOR U57519 ( .A(n57564), .B(n57565), .Z(n57560) );
  AND U57520 ( .A(n57566), .B(n57567), .Z(n57565) );
  XNOR U57521 ( .A(p_input[303]), .B(n57564), .Z(n57567) );
  XNOR U57522 ( .A(n57564), .B(n57241), .Z(n57566) );
  IV U57523 ( .A(p_input[271]), .Z(n57241) );
  XOR U57524 ( .A(n57568), .B(n57569), .Z(n57564) );
  AND U57525 ( .A(n57570), .B(n57571), .Z(n57569) );
  XNOR U57526 ( .A(p_input[302]), .B(n57568), .Z(n57571) );
  XNOR U57527 ( .A(n57568), .B(n57250), .Z(n57570) );
  IV U57528 ( .A(p_input[270]), .Z(n57250) );
  XOR U57529 ( .A(n57572), .B(n57573), .Z(n57568) );
  AND U57530 ( .A(n57574), .B(n57575), .Z(n57573) );
  XNOR U57531 ( .A(p_input[301]), .B(n57572), .Z(n57575) );
  XNOR U57532 ( .A(n57572), .B(n57259), .Z(n57574) );
  IV U57533 ( .A(p_input[269]), .Z(n57259) );
  XOR U57534 ( .A(n57576), .B(n57577), .Z(n57572) );
  AND U57535 ( .A(n57578), .B(n57579), .Z(n57577) );
  XNOR U57536 ( .A(p_input[300]), .B(n57576), .Z(n57579) );
  XNOR U57537 ( .A(n57576), .B(n57268), .Z(n57578) );
  IV U57538 ( .A(p_input[268]), .Z(n57268) );
  XOR U57539 ( .A(n57580), .B(n57581), .Z(n57576) );
  AND U57540 ( .A(n57582), .B(n57583), .Z(n57581) );
  XNOR U57541 ( .A(p_input[299]), .B(n57580), .Z(n57583) );
  XNOR U57542 ( .A(n57580), .B(n57277), .Z(n57582) );
  IV U57543 ( .A(p_input[267]), .Z(n57277) );
  XOR U57544 ( .A(n57584), .B(n57585), .Z(n57580) );
  AND U57545 ( .A(n57586), .B(n57587), .Z(n57585) );
  XNOR U57546 ( .A(p_input[298]), .B(n57584), .Z(n57587) );
  XNOR U57547 ( .A(n57584), .B(n57286), .Z(n57586) );
  IV U57548 ( .A(p_input[266]), .Z(n57286) );
  XOR U57549 ( .A(n57588), .B(n57589), .Z(n57584) );
  AND U57550 ( .A(n57590), .B(n57591), .Z(n57589) );
  XNOR U57551 ( .A(p_input[297]), .B(n57588), .Z(n57591) );
  XNOR U57552 ( .A(n57588), .B(n57295), .Z(n57590) );
  IV U57553 ( .A(p_input[265]), .Z(n57295) );
  XOR U57554 ( .A(n57592), .B(n57593), .Z(n57588) );
  AND U57555 ( .A(n57594), .B(n57595), .Z(n57593) );
  XNOR U57556 ( .A(p_input[296]), .B(n57592), .Z(n57595) );
  XNOR U57557 ( .A(n57592), .B(n57304), .Z(n57594) );
  IV U57558 ( .A(p_input[264]), .Z(n57304) );
  XOR U57559 ( .A(n57596), .B(n57597), .Z(n57592) );
  AND U57560 ( .A(n57598), .B(n57599), .Z(n57597) );
  XNOR U57561 ( .A(p_input[295]), .B(n57596), .Z(n57599) );
  XNOR U57562 ( .A(n57596), .B(n57313), .Z(n57598) );
  IV U57563 ( .A(p_input[263]), .Z(n57313) );
  XOR U57564 ( .A(n57600), .B(n57601), .Z(n57596) );
  AND U57565 ( .A(n57602), .B(n57603), .Z(n57601) );
  XNOR U57566 ( .A(p_input[294]), .B(n57600), .Z(n57603) );
  XNOR U57567 ( .A(n57600), .B(n57322), .Z(n57602) );
  IV U57568 ( .A(p_input[262]), .Z(n57322) );
  XOR U57569 ( .A(n57604), .B(n57605), .Z(n57600) );
  AND U57570 ( .A(n57606), .B(n57607), .Z(n57605) );
  XNOR U57571 ( .A(p_input[293]), .B(n57604), .Z(n57607) );
  XNOR U57572 ( .A(n57604), .B(n57331), .Z(n57606) );
  IV U57573 ( .A(p_input[261]), .Z(n57331) );
  XOR U57574 ( .A(n57608), .B(n57609), .Z(n57604) );
  AND U57575 ( .A(n57610), .B(n57611), .Z(n57609) );
  XNOR U57576 ( .A(p_input[292]), .B(n57608), .Z(n57611) );
  XNOR U57577 ( .A(n57608), .B(n57340), .Z(n57610) );
  IV U57578 ( .A(p_input[260]), .Z(n57340) );
  XOR U57579 ( .A(n57612), .B(n57613), .Z(n57608) );
  AND U57580 ( .A(n57614), .B(n57615), .Z(n57613) );
  XNOR U57581 ( .A(p_input[291]), .B(n57612), .Z(n57615) );
  XNOR U57582 ( .A(n57612), .B(n57349), .Z(n57614) );
  IV U57583 ( .A(p_input[259]), .Z(n57349) );
  XOR U57584 ( .A(n57616), .B(n57617), .Z(n57612) );
  AND U57585 ( .A(n57618), .B(n57619), .Z(n57617) );
  XNOR U57586 ( .A(p_input[290]), .B(n57616), .Z(n57619) );
  XNOR U57587 ( .A(n57616), .B(n57358), .Z(n57618) );
  IV U57588 ( .A(p_input[258]), .Z(n57358) );
  XNOR U57589 ( .A(n57620), .B(n57621), .Z(n57616) );
  AND U57590 ( .A(n57622), .B(n57623), .Z(n57621) );
  XOR U57591 ( .A(p_input[289]), .B(n57620), .Z(n57623) );
  XNOR U57592 ( .A(p_input[257]), .B(n57620), .Z(n57622) );
  AND U57593 ( .A(p_input[288]), .B(n57624), .Z(n57620) );
  IV U57594 ( .A(p_input[256]), .Z(n57624) );
  XOR U57595 ( .A(n57625), .B(n57626), .Z(n55803) );
  AND U57596 ( .A(n916), .B(n57627), .Z(n57626) );
  XNOR U57597 ( .A(n57628), .B(n57625), .Z(n57627) );
  XOR U57598 ( .A(n57629), .B(n57630), .Z(n916) );
  AND U57599 ( .A(n57631), .B(n57632), .Z(n57630) );
  XOR U57600 ( .A(n57629), .B(n55818), .Z(n57632) );
  XNOR U57601 ( .A(n57633), .B(n57634), .Z(n55818) );
  AND U57602 ( .A(n57635), .B(n667), .Z(n57634) );
  AND U57603 ( .A(n57633), .B(n57636), .Z(n57635) );
  XNOR U57604 ( .A(n55815), .B(n57629), .Z(n57631) );
  XOR U57605 ( .A(n57637), .B(n57638), .Z(n55815) );
  AND U57606 ( .A(n57639), .B(n664), .Z(n57638) );
  NOR U57607 ( .A(n57637), .B(n57640), .Z(n57639) );
  XOR U57608 ( .A(n57641), .B(n57642), .Z(n57629) );
  AND U57609 ( .A(n57643), .B(n57644), .Z(n57642) );
  XOR U57610 ( .A(n57641), .B(n55830), .Z(n57644) );
  XOR U57611 ( .A(n57645), .B(n57646), .Z(n55830) );
  AND U57612 ( .A(n667), .B(n57647), .Z(n57646) );
  XOR U57613 ( .A(n57648), .B(n57645), .Z(n57647) );
  XNOR U57614 ( .A(n55827), .B(n57641), .Z(n57643) );
  XOR U57615 ( .A(n57649), .B(n57650), .Z(n55827) );
  AND U57616 ( .A(n664), .B(n57651), .Z(n57650) );
  XOR U57617 ( .A(n57652), .B(n57649), .Z(n57651) );
  XOR U57618 ( .A(n57653), .B(n57654), .Z(n57641) );
  AND U57619 ( .A(n57655), .B(n57656), .Z(n57654) );
  XOR U57620 ( .A(n57653), .B(n55842), .Z(n57656) );
  XOR U57621 ( .A(n57657), .B(n57658), .Z(n55842) );
  AND U57622 ( .A(n667), .B(n57659), .Z(n57658) );
  XOR U57623 ( .A(n57660), .B(n57657), .Z(n57659) );
  XNOR U57624 ( .A(n55839), .B(n57653), .Z(n57655) );
  XOR U57625 ( .A(n57661), .B(n57662), .Z(n55839) );
  AND U57626 ( .A(n664), .B(n57663), .Z(n57662) );
  XOR U57627 ( .A(n57664), .B(n57661), .Z(n57663) );
  XOR U57628 ( .A(n57665), .B(n57666), .Z(n57653) );
  AND U57629 ( .A(n57667), .B(n57668), .Z(n57666) );
  XOR U57630 ( .A(n57665), .B(n55854), .Z(n57668) );
  XOR U57631 ( .A(n57669), .B(n57670), .Z(n55854) );
  AND U57632 ( .A(n667), .B(n57671), .Z(n57670) );
  XOR U57633 ( .A(n57672), .B(n57669), .Z(n57671) );
  XNOR U57634 ( .A(n55851), .B(n57665), .Z(n57667) );
  XOR U57635 ( .A(n57673), .B(n57674), .Z(n55851) );
  AND U57636 ( .A(n664), .B(n57675), .Z(n57674) );
  XOR U57637 ( .A(n57676), .B(n57673), .Z(n57675) );
  XOR U57638 ( .A(n57677), .B(n57678), .Z(n57665) );
  AND U57639 ( .A(n57679), .B(n57680), .Z(n57678) );
  XOR U57640 ( .A(n57677), .B(n55866), .Z(n57680) );
  XOR U57641 ( .A(n57681), .B(n57682), .Z(n55866) );
  AND U57642 ( .A(n667), .B(n57683), .Z(n57682) );
  XOR U57643 ( .A(n57684), .B(n57681), .Z(n57683) );
  XNOR U57644 ( .A(n55863), .B(n57677), .Z(n57679) );
  XOR U57645 ( .A(n57685), .B(n57686), .Z(n55863) );
  AND U57646 ( .A(n664), .B(n57687), .Z(n57686) );
  XOR U57647 ( .A(n57688), .B(n57685), .Z(n57687) );
  XOR U57648 ( .A(n57689), .B(n57690), .Z(n57677) );
  AND U57649 ( .A(n57691), .B(n57692), .Z(n57690) );
  XOR U57650 ( .A(n57689), .B(n55878), .Z(n57692) );
  XOR U57651 ( .A(n57693), .B(n57694), .Z(n55878) );
  AND U57652 ( .A(n667), .B(n57695), .Z(n57694) );
  XOR U57653 ( .A(n57696), .B(n57693), .Z(n57695) );
  XNOR U57654 ( .A(n55875), .B(n57689), .Z(n57691) );
  XOR U57655 ( .A(n57697), .B(n57698), .Z(n55875) );
  AND U57656 ( .A(n664), .B(n57699), .Z(n57698) );
  XOR U57657 ( .A(n57700), .B(n57697), .Z(n57699) );
  XOR U57658 ( .A(n57701), .B(n57702), .Z(n57689) );
  AND U57659 ( .A(n57703), .B(n57704), .Z(n57702) );
  XOR U57660 ( .A(n57701), .B(n55890), .Z(n57704) );
  XOR U57661 ( .A(n57705), .B(n57706), .Z(n55890) );
  AND U57662 ( .A(n667), .B(n57707), .Z(n57706) );
  XOR U57663 ( .A(n57708), .B(n57705), .Z(n57707) );
  XNOR U57664 ( .A(n55887), .B(n57701), .Z(n57703) );
  XOR U57665 ( .A(n57709), .B(n57710), .Z(n55887) );
  AND U57666 ( .A(n664), .B(n57711), .Z(n57710) );
  XOR U57667 ( .A(n57712), .B(n57709), .Z(n57711) );
  XOR U57668 ( .A(n57713), .B(n57714), .Z(n57701) );
  AND U57669 ( .A(n57715), .B(n57716), .Z(n57714) );
  XOR U57670 ( .A(n57713), .B(n55902), .Z(n57716) );
  XOR U57671 ( .A(n57717), .B(n57718), .Z(n55902) );
  AND U57672 ( .A(n667), .B(n57719), .Z(n57718) );
  XOR U57673 ( .A(n57720), .B(n57717), .Z(n57719) );
  XNOR U57674 ( .A(n55899), .B(n57713), .Z(n57715) );
  XOR U57675 ( .A(n57721), .B(n57722), .Z(n55899) );
  AND U57676 ( .A(n664), .B(n57723), .Z(n57722) );
  XOR U57677 ( .A(n57724), .B(n57721), .Z(n57723) );
  XOR U57678 ( .A(n57725), .B(n57726), .Z(n57713) );
  AND U57679 ( .A(n57727), .B(n57728), .Z(n57726) );
  XOR U57680 ( .A(n57725), .B(n55914), .Z(n57728) );
  XOR U57681 ( .A(n57729), .B(n57730), .Z(n55914) );
  AND U57682 ( .A(n667), .B(n57731), .Z(n57730) );
  XOR U57683 ( .A(n57732), .B(n57729), .Z(n57731) );
  XNOR U57684 ( .A(n55911), .B(n57725), .Z(n57727) );
  XOR U57685 ( .A(n57733), .B(n57734), .Z(n55911) );
  AND U57686 ( .A(n664), .B(n57735), .Z(n57734) );
  XOR U57687 ( .A(n57736), .B(n57733), .Z(n57735) );
  XOR U57688 ( .A(n57737), .B(n57738), .Z(n57725) );
  AND U57689 ( .A(n57739), .B(n57740), .Z(n57738) );
  XOR U57690 ( .A(n57737), .B(n55926), .Z(n57740) );
  XOR U57691 ( .A(n57741), .B(n57742), .Z(n55926) );
  AND U57692 ( .A(n667), .B(n57743), .Z(n57742) );
  XOR U57693 ( .A(n57744), .B(n57741), .Z(n57743) );
  XNOR U57694 ( .A(n55923), .B(n57737), .Z(n57739) );
  XOR U57695 ( .A(n57745), .B(n57746), .Z(n55923) );
  AND U57696 ( .A(n664), .B(n57747), .Z(n57746) );
  XOR U57697 ( .A(n57748), .B(n57745), .Z(n57747) );
  XOR U57698 ( .A(n57749), .B(n57750), .Z(n57737) );
  AND U57699 ( .A(n57751), .B(n57752), .Z(n57750) );
  XOR U57700 ( .A(n57749), .B(n55938), .Z(n57752) );
  XOR U57701 ( .A(n57753), .B(n57754), .Z(n55938) );
  AND U57702 ( .A(n667), .B(n57755), .Z(n57754) );
  XOR U57703 ( .A(n57756), .B(n57753), .Z(n57755) );
  XNOR U57704 ( .A(n55935), .B(n57749), .Z(n57751) );
  XOR U57705 ( .A(n57757), .B(n57758), .Z(n55935) );
  AND U57706 ( .A(n664), .B(n57759), .Z(n57758) );
  XOR U57707 ( .A(n57760), .B(n57757), .Z(n57759) );
  XOR U57708 ( .A(n57761), .B(n57762), .Z(n57749) );
  AND U57709 ( .A(n57763), .B(n57764), .Z(n57762) );
  XOR U57710 ( .A(n57761), .B(n55950), .Z(n57764) );
  XOR U57711 ( .A(n57765), .B(n57766), .Z(n55950) );
  AND U57712 ( .A(n667), .B(n57767), .Z(n57766) );
  XOR U57713 ( .A(n57768), .B(n57765), .Z(n57767) );
  XNOR U57714 ( .A(n55947), .B(n57761), .Z(n57763) );
  XOR U57715 ( .A(n57769), .B(n57770), .Z(n55947) );
  AND U57716 ( .A(n664), .B(n57771), .Z(n57770) );
  XOR U57717 ( .A(n57772), .B(n57769), .Z(n57771) );
  XOR U57718 ( .A(n57773), .B(n57774), .Z(n57761) );
  AND U57719 ( .A(n57775), .B(n57776), .Z(n57774) );
  XOR U57720 ( .A(n57773), .B(n55962), .Z(n57776) );
  XOR U57721 ( .A(n57777), .B(n57778), .Z(n55962) );
  AND U57722 ( .A(n667), .B(n57779), .Z(n57778) );
  XOR U57723 ( .A(n57780), .B(n57777), .Z(n57779) );
  XNOR U57724 ( .A(n55959), .B(n57773), .Z(n57775) );
  XOR U57725 ( .A(n57781), .B(n57782), .Z(n55959) );
  AND U57726 ( .A(n664), .B(n57783), .Z(n57782) );
  XOR U57727 ( .A(n57784), .B(n57781), .Z(n57783) );
  XOR U57728 ( .A(n57785), .B(n57786), .Z(n57773) );
  AND U57729 ( .A(n57787), .B(n57788), .Z(n57786) );
  XOR U57730 ( .A(n57785), .B(n55974), .Z(n57788) );
  XOR U57731 ( .A(n57789), .B(n57790), .Z(n55974) );
  AND U57732 ( .A(n667), .B(n57791), .Z(n57790) );
  XOR U57733 ( .A(n57792), .B(n57789), .Z(n57791) );
  XNOR U57734 ( .A(n55971), .B(n57785), .Z(n57787) );
  XOR U57735 ( .A(n57793), .B(n57794), .Z(n55971) );
  AND U57736 ( .A(n664), .B(n57795), .Z(n57794) );
  XOR U57737 ( .A(n57796), .B(n57793), .Z(n57795) );
  XOR U57738 ( .A(n57797), .B(n57798), .Z(n57785) );
  AND U57739 ( .A(n57799), .B(n57800), .Z(n57798) );
  XOR U57740 ( .A(n57797), .B(n55986), .Z(n57800) );
  XOR U57741 ( .A(n57801), .B(n57802), .Z(n55986) );
  AND U57742 ( .A(n667), .B(n57803), .Z(n57802) );
  XOR U57743 ( .A(n57804), .B(n57801), .Z(n57803) );
  XNOR U57744 ( .A(n55983), .B(n57797), .Z(n57799) );
  XOR U57745 ( .A(n57805), .B(n57806), .Z(n55983) );
  AND U57746 ( .A(n664), .B(n57807), .Z(n57806) );
  XOR U57747 ( .A(n57808), .B(n57805), .Z(n57807) );
  XOR U57748 ( .A(n57809), .B(n57810), .Z(n57797) );
  AND U57749 ( .A(n57811), .B(n57812), .Z(n57810) );
  XOR U57750 ( .A(n57809), .B(n55998), .Z(n57812) );
  XOR U57751 ( .A(n57813), .B(n57814), .Z(n55998) );
  AND U57752 ( .A(n667), .B(n57815), .Z(n57814) );
  XOR U57753 ( .A(n57816), .B(n57813), .Z(n57815) );
  XNOR U57754 ( .A(n55995), .B(n57809), .Z(n57811) );
  XOR U57755 ( .A(n57817), .B(n57818), .Z(n55995) );
  AND U57756 ( .A(n664), .B(n57819), .Z(n57818) );
  XOR U57757 ( .A(n57820), .B(n57817), .Z(n57819) );
  XOR U57758 ( .A(n57821), .B(n57822), .Z(n57809) );
  AND U57759 ( .A(n57823), .B(n57824), .Z(n57822) );
  XOR U57760 ( .A(n57821), .B(n56010), .Z(n57824) );
  XOR U57761 ( .A(n57825), .B(n57826), .Z(n56010) );
  AND U57762 ( .A(n667), .B(n57827), .Z(n57826) );
  XOR U57763 ( .A(n57828), .B(n57825), .Z(n57827) );
  XNOR U57764 ( .A(n56007), .B(n57821), .Z(n57823) );
  XOR U57765 ( .A(n57829), .B(n57830), .Z(n56007) );
  AND U57766 ( .A(n664), .B(n57831), .Z(n57830) );
  XOR U57767 ( .A(n57832), .B(n57829), .Z(n57831) );
  XOR U57768 ( .A(n57833), .B(n57834), .Z(n57821) );
  AND U57769 ( .A(n57835), .B(n57836), .Z(n57834) );
  XOR U57770 ( .A(n57833), .B(n56022), .Z(n57836) );
  XOR U57771 ( .A(n57837), .B(n57838), .Z(n56022) );
  AND U57772 ( .A(n667), .B(n57839), .Z(n57838) );
  XOR U57773 ( .A(n57840), .B(n57837), .Z(n57839) );
  XNOR U57774 ( .A(n56019), .B(n57833), .Z(n57835) );
  XOR U57775 ( .A(n57841), .B(n57842), .Z(n56019) );
  AND U57776 ( .A(n664), .B(n57843), .Z(n57842) );
  XOR U57777 ( .A(n57844), .B(n57841), .Z(n57843) );
  XOR U57778 ( .A(n57845), .B(n57846), .Z(n57833) );
  AND U57779 ( .A(n57847), .B(n57848), .Z(n57846) );
  XOR U57780 ( .A(n57845), .B(n56034), .Z(n57848) );
  XOR U57781 ( .A(n57849), .B(n57850), .Z(n56034) );
  AND U57782 ( .A(n667), .B(n57851), .Z(n57850) );
  XOR U57783 ( .A(n57852), .B(n57849), .Z(n57851) );
  XNOR U57784 ( .A(n56031), .B(n57845), .Z(n57847) );
  XOR U57785 ( .A(n57853), .B(n57854), .Z(n56031) );
  AND U57786 ( .A(n664), .B(n57855), .Z(n57854) );
  XOR U57787 ( .A(n57856), .B(n57853), .Z(n57855) );
  XOR U57788 ( .A(n57857), .B(n57858), .Z(n57845) );
  AND U57789 ( .A(n57859), .B(n57860), .Z(n57858) );
  XOR U57790 ( .A(n57857), .B(n56046), .Z(n57860) );
  XOR U57791 ( .A(n57861), .B(n57862), .Z(n56046) );
  AND U57792 ( .A(n667), .B(n57863), .Z(n57862) );
  XOR U57793 ( .A(n57864), .B(n57861), .Z(n57863) );
  XNOR U57794 ( .A(n56043), .B(n57857), .Z(n57859) );
  XOR U57795 ( .A(n57865), .B(n57866), .Z(n56043) );
  AND U57796 ( .A(n664), .B(n57867), .Z(n57866) );
  XOR U57797 ( .A(n57868), .B(n57865), .Z(n57867) );
  XOR U57798 ( .A(n57869), .B(n57870), .Z(n57857) );
  AND U57799 ( .A(n57871), .B(n57872), .Z(n57870) );
  XOR U57800 ( .A(n57869), .B(n56058), .Z(n57872) );
  XOR U57801 ( .A(n57873), .B(n57874), .Z(n56058) );
  AND U57802 ( .A(n667), .B(n57875), .Z(n57874) );
  XOR U57803 ( .A(n57876), .B(n57873), .Z(n57875) );
  XNOR U57804 ( .A(n56055), .B(n57869), .Z(n57871) );
  XOR U57805 ( .A(n57877), .B(n57878), .Z(n56055) );
  AND U57806 ( .A(n664), .B(n57879), .Z(n57878) );
  XOR U57807 ( .A(n57880), .B(n57877), .Z(n57879) );
  XOR U57808 ( .A(n57881), .B(n57882), .Z(n57869) );
  AND U57809 ( .A(n57883), .B(n57884), .Z(n57882) );
  XOR U57810 ( .A(n57881), .B(n56070), .Z(n57884) );
  XOR U57811 ( .A(n57885), .B(n57886), .Z(n56070) );
  AND U57812 ( .A(n667), .B(n57887), .Z(n57886) );
  XOR U57813 ( .A(n57888), .B(n57885), .Z(n57887) );
  XNOR U57814 ( .A(n56067), .B(n57881), .Z(n57883) );
  XOR U57815 ( .A(n57889), .B(n57890), .Z(n56067) );
  AND U57816 ( .A(n664), .B(n57891), .Z(n57890) );
  XOR U57817 ( .A(n57892), .B(n57889), .Z(n57891) );
  XOR U57818 ( .A(n57893), .B(n57894), .Z(n57881) );
  AND U57819 ( .A(n57895), .B(n57896), .Z(n57894) );
  XOR U57820 ( .A(n57893), .B(n56082), .Z(n57896) );
  XOR U57821 ( .A(n57897), .B(n57898), .Z(n56082) );
  AND U57822 ( .A(n667), .B(n57899), .Z(n57898) );
  XOR U57823 ( .A(n57900), .B(n57897), .Z(n57899) );
  XNOR U57824 ( .A(n56079), .B(n57893), .Z(n57895) );
  XOR U57825 ( .A(n57901), .B(n57902), .Z(n56079) );
  AND U57826 ( .A(n664), .B(n57903), .Z(n57902) );
  XOR U57827 ( .A(n57904), .B(n57901), .Z(n57903) );
  XOR U57828 ( .A(n57905), .B(n57906), .Z(n57893) );
  AND U57829 ( .A(n57907), .B(n57908), .Z(n57906) );
  XOR U57830 ( .A(n57905), .B(n56094), .Z(n57908) );
  XOR U57831 ( .A(n57909), .B(n57910), .Z(n56094) );
  AND U57832 ( .A(n667), .B(n57911), .Z(n57910) );
  XOR U57833 ( .A(n57912), .B(n57909), .Z(n57911) );
  XNOR U57834 ( .A(n56091), .B(n57905), .Z(n57907) );
  XOR U57835 ( .A(n57913), .B(n57914), .Z(n56091) );
  AND U57836 ( .A(n664), .B(n57915), .Z(n57914) );
  XOR U57837 ( .A(n57916), .B(n57913), .Z(n57915) );
  XOR U57838 ( .A(n57917), .B(n57918), .Z(n57905) );
  AND U57839 ( .A(n57919), .B(n57920), .Z(n57918) );
  XOR U57840 ( .A(n57917), .B(n56106), .Z(n57920) );
  XOR U57841 ( .A(n57921), .B(n57922), .Z(n56106) );
  AND U57842 ( .A(n667), .B(n57923), .Z(n57922) );
  XOR U57843 ( .A(n57924), .B(n57921), .Z(n57923) );
  XNOR U57844 ( .A(n56103), .B(n57917), .Z(n57919) );
  XOR U57845 ( .A(n57925), .B(n57926), .Z(n56103) );
  AND U57846 ( .A(n664), .B(n57927), .Z(n57926) );
  XOR U57847 ( .A(n57928), .B(n57925), .Z(n57927) );
  XOR U57848 ( .A(n57929), .B(n57930), .Z(n57917) );
  AND U57849 ( .A(n57931), .B(n57932), .Z(n57930) );
  XOR U57850 ( .A(n57929), .B(n56118), .Z(n57932) );
  XOR U57851 ( .A(n57933), .B(n57934), .Z(n56118) );
  AND U57852 ( .A(n667), .B(n57935), .Z(n57934) );
  XOR U57853 ( .A(n57936), .B(n57933), .Z(n57935) );
  XNOR U57854 ( .A(n56115), .B(n57929), .Z(n57931) );
  XOR U57855 ( .A(n57937), .B(n57938), .Z(n56115) );
  AND U57856 ( .A(n664), .B(n57939), .Z(n57938) );
  XOR U57857 ( .A(n57940), .B(n57937), .Z(n57939) );
  XOR U57858 ( .A(n57941), .B(n57942), .Z(n57929) );
  AND U57859 ( .A(n57943), .B(n57944), .Z(n57942) );
  XOR U57860 ( .A(n57941), .B(n56130), .Z(n57944) );
  XOR U57861 ( .A(n57945), .B(n57946), .Z(n56130) );
  AND U57862 ( .A(n667), .B(n57947), .Z(n57946) );
  XOR U57863 ( .A(n57948), .B(n57945), .Z(n57947) );
  XNOR U57864 ( .A(n56127), .B(n57941), .Z(n57943) );
  XOR U57865 ( .A(n57949), .B(n57950), .Z(n56127) );
  AND U57866 ( .A(n664), .B(n57951), .Z(n57950) );
  XOR U57867 ( .A(n57952), .B(n57949), .Z(n57951) );
  XOR U57868 ( .A(n57953), .B(n57954), .Z(n57941) );
  AND U57869 ( .A(n57955), .B(n57956), .Z(n57954) );
  XOR U57870 ( .A(n57953), .B(n56142), .Z(n57956) );
  XOR U57871 ( .A(n57957), .B(n57958), .Z(n56142) );
  AND U57872 ( .A(n667), .B(n57959), .Z(n57958) );
  XOR U57873 ( .A(n57960), .B(n57957), .Z(n57959) );
  XNOR U57874 ( .A(n56139), .B(n57953), .Z(n57955) );
  XOR U57875 ( .A(n57961), .B(n57962), .Z(n56139) );
  AND U57876 ( .A(n664), .B(n57963), .Z(n57962) );
  XOR U57877 ( .A(n57964), .B(n57961), .Z(n57963) );
  XOR U57878 ( .A(n57965), .B(n57966), .Z(n57953) );
  AND U57879 ( .A(n57967), .B(n57968), .Z(n57966) );
  XOR U57880 ( .A(n57965), .B(n56154), .Z(n57968) );
  XOR U57881 ( .A(n57969), .B(n57970), .Z(n56154) );
  AND U57882 ( .A(n667), .B(n57971), .Z(n57970) );
  XOR U57883 ( .A(n57972), .B(n57969), .Z(n57971) );
  XNOR U57884 ( .A(n56151), .B(n57965), .Z(n57967) );
  XOR U57885 ( .A(n57973), .B(n57974), .Z(n56151) );
  AND U57886 ( .A(n664), .B(n57975), .Z(n57974) );
  XOR U57887 ( .A(n57976), .B(n57973), .Z(n57975) );
  XOR U57888 ( .A(n57977), .B(n57978), .Z(n57965) );
  AND U57889 ( .A(n57979), .B(n57980), .Z(n57978) );
  XOR U57890 ( .A(n57977), .B(n56166), .Z(n57980) );
  XOR U57891 ( .A(n57981), .B(n57982), .Z(n56166) );
  AND U57892 ( .A(n667), .B(n57983), .Z(n57982) );
  XOR U57893 ( .A(n57984), .B(n57981), .Z(n57983) );
  XNOR U57894 ( .A(n56163), .B(n57977), .Z(n57979) );
  XOR U57895 ( .A(n57985), .B(n57986), .Z(n56163) );
  AND U57896 ( .A(n664), .B(n57987), .Z(n57986) );
  XOR U57897 ( .A(n57988), .B(n57985), .Z(n57987) );
  XOR U57898 ( .A(n57989), .B(n57990), .Z(n57977) );
  AND U57899 ( .A(n57991), .B(n57992), .Z(n57990) );
  XNOR U57900 ( .A(n57993), .B(n56179), .Z(n57992) );
  XOR U57901 ( .A(n57994), .B(n57995), .Z(n56179) );
  AND U57902 ( .A(n667), .B(n57996), .Z(n57995) );
  XOR U57903 ( .A(n57994), .B(n57997), .Z(n57996) );
  XNOR U57904 ( .A(n56176), .B(n57989), .Z(n57991) );
  XOR U57905 ( .A(n57998), .B(n57999), .Z(n56176) );
  AND U57906 ( .A(n664), .B(n58000), .Z(n57999) );
  XOR U57907 ( .A(n57998), .B(n58001), .Z(n58000) );
  IV U57908 ( .A(n57993), .Z(n57989) );
  AND U57909 ( .A(n57625), .B(n57628), .Z(n57993) );
  XNOR U57910 ( .A(n58002), .B(n58003), .Z(n57628) );
  AND U57911 ( .A(n667), .B(n58004), .Z(n58003) );
  XNOR U57912 ( .A(n58005), .B(n58002), .Z(n58004) );
  XOR U57913 ( .A(n58006), .B(n58007), .Z(n667) );
  AND U57914 ( .A(n58008), .B(n58009), .Z(n58007) );
  XOR U57915 ( .A(n57636), .B(n58006), .Z(n58009) );
  IV U57916 ( .A(n58010), .Z(n57636) );
  AND U57917 ( .A(p_input[255]), .B(p_input[223]), .Z(n58010) );
  XOR U57918 ( .A(n58006), .B(n57633), .Z(n58008) );
  AND U57919 ( .A(p_input[159]), .B(p_input[191]), .Z(n57633) );
  XOR U57920 ( .A(n58011), .B(n58012), .Z(n58006) );
  AND U57921 ( .A(n58013), .B(n58014), .Z(n58012) );
  XOR U57922 ( .A(n58011), .B(n57648), .Z(n58014) );
  XNOR U57923 ( .A(p_input[222]), .B(n58015), .Z(n57648) );
  AND U57924 ( .A(n1139), .B(n58016), .Z(n58015) );
  XOR U57925 ( .A(p_input[254]), .B(p_input[222]), .Z(n58016) );
  XNOR U57926 ( .A(n57645), .B(n58011), .Z(n58013) );
  XOR U57927 ( .A(n58017), .B(n58018), .Z(n57645) );
  AND U57928 ( .A(n1137), .B(n58019), .Z(n58018) );
  XOR U57929 ( .A(p_input[190]), .B(p_input[158]), .Z(n58019) );
  XOR U57930 ( .A(n58020), .B(n58021), .Z(n58011) );
  AND U57931 ( .A(n58022), .B(n58023), .Z(n58021) );
  XOR U57932 ( .A(n58020), .B(n57660), .Z(n58023) );
  XNOR U57933 ( .A(p_input[221]), .B(n58024), .Z(n57660) );
  AND U57934 ( .A(n1139), .B(n58025), .Z(n58024) );
  XOR U57935 ( .A(p_input[253]), .B(p_input[221]), .Z(n58025) );
  XNOR U57936 ( .A(n57657), .B(n58020), .Z(n58022) );
  XOR U57937 ( .A(n58026), .B(n58027), .Z(n57657) );
  AND U57938 ( .A(n1137), .B(n58028), .Z(n58027) );
  XOR U57939 ( .A(p_input[189]), .B(p_input[157]), .Z(n58028) );
  XOR U57940 ( .A(n58029), .B(n58030), .Z(n58020) );
  AND U57941 ( .A(n58031), .B(n58032), .Z(n58030) );
  XOR U57942 ( .A(n58029), .B(n57672), .Z(n58032) );
  XNOR U57943 ( .A(p_input[220]), .B(n58033), .Z(n57672) );
  AND U57944 ( .A(n1139), .B(n58034), .Z(n58033) );
  XOR U57945 ( .A(p_input[252]), .B(p_input[220]), .Z(n58034) );
  XNOR U57946 ( .A(n57669), .B(n58029), .Z(n58031) );
  XOR U57947 ( .A(n58035), .B(n58036), .Z(n57669) );
  AND U57948 ( .A(n1137), .B(n58037), .Z(n58036) );
  XOR U57949 ( .A(p_input[188]), .B(p_input[156]), .Z(n58037) );
  XOR U57950 ( .A(n58038), .B(n58039), .Z(n58029) );
  AND U57951 ( .A(n58040), .B(n58041), .Z(n58039) );
  XOR U57952 ( .A(n58038), .B(n57684), .Z(n58041) );
  XNOR U57953 ( .A(p_input[219]), .B(n58042), .Z(n57684) );
  AND U57954 ( .A(n1139), .B(n58043), .Z(n58042) );
  XOR U57955 ( .A(p_input[251]), .B(p_input[219]), .Z(n58043) );
  XNOR U57956 ( .A(n57681), .B(n58038), .Z(n58040) );
  XOR U57957 ( .A(n58044), .B(n58045), .Z(n57681) );
  AND U57958 ( .A(n1137), .B(n58046), .Z(n58045) );
  XOR U57959 ( .A(p_input[187]), .B(p_input[155]), .Z(n58046) );
  XOR U57960 ( .A(n58047), .B(n58048), .Z(n58038) );
  AND U57961 ( .A(n58049), .B(n58050), .Z(n58048) );
  XOR U57962 ( .A(n58047), .B(n57696), .Z(n58050) );
  XNOR U57963 ( .A(p_input[218]), .B(n58051), .Z(n57696) );
  AND U57964 ( .A(n1139), .B(n58052), .Z(n58051) );
  XOR U57965 ( .A(p_input[250]), .B(p_input[218]), .Z(n58052) );
  XNOR U57966 ( .A(n57693), .B(n58047), .Z(n58049) );
  XOR U57967 ( .A(n58053), .B(n58054), .Z(n57693) );
  AND U57968 ( .A(n1137), .B(n58055), .Z(n58054) );
  XOR U57969 ( .A(p_input[186]), .B(p_input[154]), .Z(n58055) );
  XOR U57970 ( .A(n58056), .B(n58057), .Z(n58047) );
  AND U57971 ( .A(n58058), .B(n58059), .Z(n58057) );
  XOR U57972 ( .A(n58056), .B(n57708), .Z(n58059) );
  XNOR U57973 ( .A(p_input[217]), .B(n58060), .Z(n57708) );
  AND U57974 ( .A(n1139), .B(n58061), .Z(n58060) );
  XOR U57975 ( .A(p_input[249]), .B(p_input[217]), .Z(n58061) );
  XNOR U57976 ( .A(n57705), .B(n58056), .Z(n58058) );
  XOR U57977 ( .A(n58062), .B(n58063), .Z(n57705) );
  AND U57978 ( .A(n1137), .B(n58064), .Z(n58063) );
  XOR U57979 ( .A(p_input[185]), .B(p_input[153]), .Z(n58064) );
  XOR U57980 ( .A(n58065), .B(n58066), .Z(n58056) );
  AND U57981 ( .A(n58067), .B(n58068), .Z(n58066) );
  XOR U57982 ( .A(n58065), .B(n57720), .Z(n58068) );
  XNOR U57983 ( .A(p_input[216]), .B(n58069), .Z(n57720) );
  AND U57984 ( .A(n1139), .B(n58070), .Z(n58069) );
  XOR U57985 ( .A(p_input[248]), .B(p_input[216]), .Z(n58070) );
  XNOR U57986 ( .A(n57717), .B(n58065), .Z(n58067) );
  XOR U57987 ( .A(n58071), .B(n58072), .Z(n57717) );
  AND U57988 ( .A(n1137), .B(n58073), .Z(n58072) );
  XOR U57989 ( .A(p_input[184]), .B(p_input[152]), .Z(n58073) );
  XOR U57990 ( .A(n58074), .B(n58075), .Z(n58065) );
  AND U57991 ( .A(n58076), .B(n58077), .Z(n58075) );
  XOR U57992 ( .A(n58074), .B(n57732), .Z(n58077) );
  XNOR U57993 ( .A(p_input[215]), .B(n58078), .Z(n57732) );
  AND U57994 ( .A(n1139), .B(n58079), .Z(n58078) );
  XOR U57995 ( .A(p_input[247]), .B(p_input[215]), .Z(n58079) );
  XNOR U57996 ( .A(n57729), .B(n58074), .Z(n58076) );
  XOR U57997 ( .A(n58080), .B(n58081), .Z(n57729) );
  AND U57998 ( .A(n1137), .B(n58082), .Z(n58081) );
  XOR U57999 ( .A(p_input[183]), .B(p_input[151]), .Z(n58082) );
  XOR U58000 ( .A(n58083), .B(n58084), .Z(n58074) );
  AND U58001 ( .A(n58085), .B(n58086), .Z(n58084) );
  XOR U58002 ( .A(n58083), .B(n57744), .Z(n58086) );
  XNOR U58003 ( .A(p_input[214]), .B(n58087), .Z(n57744) );
  AND U58004 ( .A(n1139), .B(n58088), .Z(n58087) );
  XOR U58005 ( .A(p_input[246]), .B(p_input[214]), .Z(n58088) );
  XNOR U58006 ( .A(n57741), .B(n58083), .Z(n58085) );
  XOR U58007 ( .A(n58089), .B(n58090), .Z(n57741) );
  AND U58008 ( .A(n1137), .B(n58091), .Z(n58090) );
  XOR U58009 ( .A(p_input[182]), .B(p_input[150]), .Z(n58091) );
  XOR U58010 ( .A(n58092), .B(n58093), .Z(n58083) );
  AND U58011 ( .A(n58094), .B(n58095), .Z(n58093) );
  XOR U58012 ( .A(n58092), .B(n57756), .Z(n58095) );
  XNOR U58013 ( .A(p_input[213]), .B(n58096), .Z(n57756) );
  AND U58014 ( .A(n1139), .B(n58097), .Z(n58096) );
  XOR U58015 ( .A(p_input[245]), .B(p_input[213]), .Z(n58097) );
  XNOR U58016 ( .A(n57753), .B(n58092), .Z(n58094) );
  XOR U58017 ( .A(n58098), .B(n58099), .Z(n57753) );
  AND U58018 ( .A(n1137), .B(n58100), .Z(n58099) );
  XOR U58019 ( .A(p_input[181]), .B(p_input[149]), .Z(n58100) );
  XOR U58020 ( .A(n58101), .B(n58102), .Z(n58092) );
  AND U58021 ( .A(n58103), .B(n58104), .Z(n58102) );
  XOR U58022 ( .A(n58101), .B(n57768), .Z(n58104) );
  XNOR U58023 ( .A(p_input[212]), .B(n58105), .Z(n57768) );
  AND U58024 ( .A(n1139), .B(n58106), .Z(n58105) );
  XOR U58025 ( .A(p_input[244]), .B(p_input[212]), .Z(n58106) );
  XNOR U58026 ( .A(n57765), .B(n58101), .Z(n58103) );
  XOR U58027 ( .A(n58107), .B(n58108), .Z(n57765) );
  AND U58028 ( .A(n1137), .B(n58109), .Z(n58108) );
  XOR U58029 ( .A(p_input[180]), .B(p_input[148]), .Z(n58109) );
  XOR U58030 ( .A(n58110), .B(n58111), .Z(n58101) );
  AND U58031 ( .A(n58112), .B(n58113), .Z(n58111) );
  XOR U58032 ( .A(n58110), .B(n57780), .Z(n58113) );
  XNOR U58033 ( .A(p_input[211]), .B(n58114), .Z(n57780) );
  AND U58034 ( .A(n1139), .B(n58115), .Z(n58114) );
  XOR U58035 ( .A(p_input[243]), .B(p_input[211]), .Z(n58115) );
  XNOR U58036 ( .A(n57777), .B(n58110), .Z(n58112) );
  XOR U58037 ( .A(n58116), .B(n58117), .Z(n57777) );
  AND U58038 ( .A(n1137), .B(n58118), .Z(n58117) );
  XOR U58039 ( .A(p_input[179]), .B(p_input[147]), .Z(n58118) );
  XOR U58040 ( .A(n58119), .B(n58120), .Z(n58110) );
  AND U58041 ( .A(n58121), .B(n58122), .Z(n58120) );
  XOR U58042 ( .A(n58119), .B(n57792), .Z(n58122) );
  XNOR U58043 ( .A(p_input[210]), .B(n58123), .Z(n57792) );
  AND U58044 ( .A(n1139), .B(n58124), .Z(n58123) );
  XOR U58045 ( .A(p_input[242]), .B(p_input[210]), .Z(n58124) );
  XNOR U58046 ( .A(n57789), .B(n58119), .Z(n58121) );
  XOR U58047 ( .A(n58125), .B(n58126), .Z(n57789) );
  AND U58048 ( .A(n1137), .B(n58127), .Z(n58126) );
  XOR U58049 ( .A(p_input[178]), .B(p_input[146]), .Z(n58127) );
  XOR U58050 ( .A(n58128), .B(n58129), .Z(n58119) );
  AND U58051 ( .A(n58130), .B(n58131), .Z(n58129) );
  XOR U58052 ( .A(n58128), .B(n57804), .Z(n58131) );
  XNOR U58053 ( .A(p_input[209]), .B(n58132), .Z(n57804) );
  AND U58054 ( .A(n1139), .B(n58133), .Z(n58132) );
  XOR U58055 ( .A(p_input[241]), .B(p_input[209]), .Z(n58133) );
  XNOR U58056 ( .A(n57801), .B(n58128), .Z(n58130) );
  XOR U58057 ( .A(n58134), .B(n58135), .Z(n57801) );
  AND U58058 ( .A(n1137), .B(n58136), .Z(n58135) );
  XOR U58059 ( .A(p_input[177]), .B(p_input[145]), .Z(n58136) );
  XOR U58060 ( .A(n58137), .B(n58138), .Z(n58128) );
  AND U58061 ( .A(n58139), .B(n58140), .Z(n58138) );
  XOR U58062 ( .A(n58137), .B(n57816), .Z(n58140) );
  XNOR U58063 ( .A(p_input[208]), .B(n58141), .Z(n57816) );
  AND U58064 ( .A(n1139), .B(n58142), .Z(n58141) );
  XOR U58065 ( .A(p_input[240]), .B(p_input[208]), .Z(n58142) );
  XNOR U58066 ( .A(n57813), .B(n58137), .Z(n58139) );
  XOR U58067 ( .A(n58143), .B(n58144), .Z(n57813) );
  AND U58068 ( .A(n1137), .B(n58145), .Z(n58144) );
  XOR U58069 ( .A(p_input[176]), .B(p_input[144]), .Z(n58145) );
  XOR U58070 ( .A(n58146), .B(n58147), .Z(n58137) );
  AND U58071 ( .A(n58148), .B(n58149), .Z(n58147) );
  XOR U58072 ( .A(n58146), .B(n57828), .Z(n58149) );
  XNOR U58073 ( .A(p_input[207]), .B(n58150), .Z(n57828) );
  AND U58074 ( .A(n1139), .B(n58151), .Z(n58150) );
  XOR U58075 ( .A(p_input[239]), .B(p_input[207]), .Z(n58151) );
  XNOR U58076 ( .A(n57825), .B(n58146), .Z(n58148) );
  XOR U58077 ( .A(n58152), .B(n58153), .Z(n57825) );
  AND U58078 ( .A(n1137), .B(n58154), .Z(n58153) );
  XOR U58079 ( .A(p_input[175]), .B(p_input[143]), .Z(n58154) );
  XOR U58080 ( .A(n58155), .B(n58156), .Z(n58146) );
  AND U58081 ( .A(n58157), .B(n58158), .Z(n58156) );
  XOR U58082 ( .A(n58155), .B(n57840), .Z(n58158) );
  XNOR U58083 ( .A(p_input[206]), .B(n58159), .Z(n57840) );
  AND U58084 ( .A(n1139), .B(n58160), .Z(n58159) );
  XOR U58085 ( .A(p_input[238]), .B(p_input[206]), .Z(n58160) );
  XNOR U58086 ( .A(n57837), .B(n58155), .Z(n58157) );
  XOR U58087 ( .A(n58161), .B(n58162), .Z(n57837) );
  AND U58088 ( .A(n1137), .B(n58163), .Z(n58162) );
  XOR U58089 ( .A(p_input[174]), .B(p_input[142]), .Z(n58163) );
  XOR U58090 ( .A(n58164), .B(n58165), .Z(n58155) );
  AND U58091 ( .A(n58166), .B(n58167), .Z(n58165) );
  XOR U58092 ( .A(n58164), .B(n57852), .Z(n58167) );
  XNOR U58093 ( .A(p_input[205]), .B(n58168), .Z(n57852) );
  AND U58094 ( .A(n1139), .B(n58169), .Z(n58168) );
  XOR U58095 ( .A(p_input[237]), .B(p_input[205]), .Z(n58169) );
  XNOR U58096 ( .A(n57849), .B(n58164), .Z(n58166) );
  XOR U58097 ( .A(n58170), .B(n58171), .Z(n57849) );
  AND U58098 ( .A(n1137), .B(n58172), .Z(n58171) );
  XOR U58099 ( .A(p_input[173]), .B(p_input[141]), .Z(n58172) );
  XOR U58100 ( .A(n58173), .B(n58174), .Z(n58164) );
  AND U58101 ( .A(n58175), .B(n58176), .Z(n58174) );
  XOR U58102 ( .A(n58173), .B(n57864), .Z(n58176) );
  XNOR U58103 ( .A(p_input[204]), .B(n58177), .Z(n57864) );
  AND U58104 ( .A(n1139), .B(n58178), .Z(n58177) );
  XOR U58105 ( .A(p_input[236]), .B(p_input[204]), .Z(n58178) );
  XNOR U58106 ( .A(n57861), .B(n58173), .Z(n58175) );
  XOR U58107 ( .A(n58179), .B(n58180), .Z(n57861) );
  AND U58108 ( .A(n1137), .B(n58181), .Z(n58180) );
  XOR U58109 ( .A(p_input[172]), .B(p_input[140]), .Z(n58181) );
  XOR U58110 ( .A(n58182), .B(n58183), .Z(n58173) );
  AND U58111 ( .A(n58184), .B(n58185), .Z(n58183) );
  XOR U58112 ( .A(n58182), .B(n57876), .Z(n58185) );
  XNOR U58113 ( .A(p_input[203]), .B(n58186), .Z(n57876) );
  AND U58114 ( .A(n1139), .B(n58187), .Z(n58186) );
  XOR U58115 ( .A(p_input[235]), .B(p_input[203]), .Z(n58187) );
  XNOR U58116 ( .A(n57873), .B(n58182), .Z(n58184) );
  XOR U58117 ( .A(n58188), .B(n58189), .Z(n57873) );
  AND U58118 ( .A(n1137), .B(n58190), .Z(n58189) );
  XOR U58119 ( .A(p_input[171]), .B(p_input[139]), .Z(n58190) );
  XOR U58120 ( .A(n58191), .B(n58192), .Z(n58182) );
  AND U58121 ( .A(n58193), .B(n58194), .Z(n58192) );
  XOR U58122 ( .A(n58191), .B(n57888), .Z(n58194) );
  XNOR U58123 ( .A(p_input[202]), .B(n58195), .Z(n57888) );
  AND U58124 ( .A(n1139), .B(n58196), .Z(n58195) );
  XOR U58125 ( .A(p_input[234]), .B(p_input[202]), .Z(n58196) );
  XNOR U58126 ( .A(n57885), .B(n58191), .Z(n58193) );
  XOR U58127 ( .A(n58197), .B(n58198), .Z(n57885) );
  AND U58128 ( .A(n1137), .B(n58199), .Z(n58198) );
  XOR U58129 ( .A(p_input[170]), .B(p_input[138]), .Z(n58199) );
  XOR U58130 ( .A(n58200), .B(n58201), .Z(n58191) );
  AND U58131 ( .A(n58202), .B(n58203), .Z(n58201) );
  XOR U58132 ( .A(n58200), .B(n57900), .Z(n58203) );
  XNOR U58133 ( .A(p_input[201]), .B(n58204), .Z(n57900) );
  AND U58134 ( .A(n1139), .B(n58205), .Z(n58204) );
  XOR U58135 ( .A(p_input[233]), .B(p_input[201]), .Z(n58205) );
  XNOR U58136 ( .A(n57897), .B(n58200), .Z(n58202) );
  XOR U58137 ( .A(n58206), .B(n58207), .Z(n57897) );
  AND U58138 ( .A(n1137), .B(n58208), .Z(n58207) );
  XOR U58139 ( .A(p_input[169]), .B(p_input[137]), .Z(n58208) );
  XOR U58140 ( .A(n58209), .B(n58210), .Z(n58200) );
  AND U58141 ( .A(n58211), .B(n58212), .Z(n58210) );
  XOR U58142 ( .A(n58209), .B(n57912), .Z(n58212) );
  XNOR U58143 ( .A(p_input[200]), .B(n58213), .Z(n57912) );
  AND U58144 ( .A(n1139), .B(n58214), .Z(n58213) );
  XOR U58145 ( .A(p_input[232]), .B(p_input[200]), .Z(n58214) );
  XNOR U58146 ( .A(n57909), .B(n58209), .Z(n58211) );
  XOR U58147 ( .A(n58215), .B(n58216), .Z(n57909) );
  AND U58148 ( .A(n1137), .B(n58217), .Z(n58216) );
  XOR U58149 ( .A(p_input[168]), .B(p_input[136]), .Z(n58217) );
  XOR U58150 ( .A(n58218), .B(n58219), .Z(n58209) );
  AND U58151 ( .A(n58220), .B(n58221), .Z(n58219) );
  XOR U58152 ( .A(n58218), .B(n57924), .Z(n58221) );
  XNOR U58153 ( .A(p_input[199]), .B(n58222), .Z(n57924) );
  AND U58154 ( .A(n1139), .B(n58223), .Z(n58222) );
  XOR U58155 ( .A(p_input[231]), .B(p_input[199]), .Z(n58223) );
  XNOR U58156 ( .A(n57921), .B(n58218), .Z(n58220) );
  XOR U58157 ( .A(n58224), .B(n58225), .Z(n57921) );
  AND U58158 ( .A(n1137), .B(n58226), .Z(n58225) );
  XOR U58159 ( .A(p_input[167]), .B(p_input[135]), .Z(n58226) );
  XOR U58160 ( .A(n58227), .B(n58228), .Z(n58218) );
  AND U58161 ( .A(n58229), .B(n58230), .Z(n58228) );
  XOR U58162 ( .A(n58227), .B(n57936), .Z(n58230) );
  XNOR U58163 ( .A(p_input[198]), .B(n58231), .Z(n57936) );
  AND U58164 ( .A(n1139), .B(n58232), .Z(n58231) );
  XOR U58165 ( .A(p_input[230]), .B(p_input[198]), .Z(n58232) );
  XNOR U58166 ( .A(n57933), .B(n58227), .Z(n58229) );
  XOR U58167 ( .A(n58233), .B(n58234), .Z(n57933) );
  AND U58168 ( .A(n1137), .B(n58235), .Z(n58234) );
  XOR U58169 ( .A(p_input[166]), .B(p_input[134]), .Z(n58235) );
  XOR U58170 ( .A(n58236), .B(n58237), .Z(n58227) );
  AND U58171 ( .A(n58238), .B(n58239), .Z(n58237) );
  XOR U58172 ( .A(n58236), .B(n57948), .Z(n58239) );
  XNOR U58173 ( .A(p_input[197]), .B(n58240), .Z(n57948) );
  AND U58174 ( .A(n1139), .B(n58241), .Z(n58240) );
  XOR U58175 ( .A(p_input[229]), .B(p_input[197]), .Z(n58241) );
  XNOR U58176 ( .A(n57945), .B(n58236), .Z(n58238) );
  XOR U58177 ( .A(n58242), .B(n58243), .Z(n57945) );
  AND U58178 ( .A(n1137), .B(n58244), .Z(n58243) );
  XOR U58179 ( .A(p_input[165]), .B(p_input[133]), .Z(n58244) );
  XOR U58180 ( .A(n58245), .B(n58246), .Z(n58236) );
  AND U58181 ( .A(n58247), .B(n58248), .Z(n58246) );
  XOR U58182 ( .A(n58245), .B(n57960), .Z(n58248) );
  XNOR U58183 ( .A(p_input[196]), .B(n58249), .Z(n57960) );
  AND U58184 ( .A(n1139), .B(n58250), .Z(n58249) );
  XOR U58185 ( .A(p_input[228]), .B(p_input[196]), .Z(n58250) );
  XNOR U58186 ( .A(n57957), .B(n58245), .Z(n58247) );
  XOR U58187 ( .A(n58251), .B(n58252), .Z(n57957) );
  AND U58188 ( .A(n1137), .B(n58253), .Z(n58252) );
  XOR U58189 ( .A(p_input[164]), .B(p_input[132]), .Z(n58253) );
  XOR U58190 ( .A(n58254), .B(n58255), .Z(n58245) );
  AND U58191 ( .A(n58256), .B(n58257), .Z(n58255) );
  XOR U58192 ( .A(n58254), .B(n57972), .Z(n58257) );
  XNOR U58193 ( .A(p_input[195]), .B(n58258), .Z(n57972) );
  AND U58194 ( .A(n1139), .B(n58259), .Z(n58258) );
  XOR U58195 ( .A(p_input[227]), .B(p_input[195]), .Z(n58259) );
  XNOR U58196 ( .A(n57969), .B(n58254), .Z(n58256) );
  XOR U58197 ( .A(n58260), .B(n58261), .Z(n57969) );
  AND U58198 ( .A(n1137), .B(n58262), .Z(n58261) );
  XOR U58199 ( .A(p_input[163]), .B(p_input[131]), .Z(n58262) );
  XOR U58200 ( .A(n58263), .B(n58264), .Z(n58254) );
  AND U58201 ( .A(n58265), .B(n58266), .Z(n58264) );
  XOR U58202 ( .A(n58263), .B(n57984), .Z(n58266) );
  XNOR U58203 ( .A(p_input[194]), .B(n58267), .Z(n57984) );
  AND U58204 ( .A(n1139), .B(n58268), .Z(n58267) );
  XOR U58205 ( .A(p_input[226]), .B(p_input[194]), .Z(n58268) );
  XNOR U58206 ( .A(n57981), .B(n58263), .Z(n58265) );
  XOR U58207 ( .A(n58269), .B(n58270), .Z(n57981) );
  AND U58208 ( .A(n1137), .B(n58271), .Z(n58270) );
  XOR U58209 ( .A(p_input[162]), .B(p_input[130]), .Z(n58271) );
  XOR U58210 ( .A(n58272), .B(n58273), .Z(n58263) );
  AND U58211 ( .A(n58274), .B(n58275), .Z(n58273) );
  XNOR U58212 ( .A(n58276), .B(n57997), .Z(n58275) );
  XNOR U58213 ( .A(p_input[193]), .B(n58277), .Z(n57997) );
  AND U58214 ( .A(n1139), .B(n58278), .Z(n58277) );
  XNOR U58215 ( .A(p_input[225]), .B(n58279), .Z(n58278) );
  IV U58216 ( .A(p_input[193]), .Z(n58279) );
  XNOR U58217 ( .A(n57994), .B(n58272), .Z(n58274) );
  XNOR U58218 ( .A(p_input[129]), .B(n58280), .Z(n57994) );
  AND U58219 ( .A(n1137), .B(n58281), .Z(n58280) );
  XOR U58220 ( .A(p_input[161]), .B(p_input[129]), .Z(n58281) );
  IV U58221 ( .A(n58276), .Z(n58272) );
  AND U58222 ( .A(n58002), .B(n58005), .Z(n58276) );
  XOR U58223 ( .A(p_input[192]), .B(n58282), .Z(n58005) );
  AND U58224 ( .A(n1139), .B(n58283), .Z(n58282) );
  XOR U58225 ( .A(p_input[224]), .B(p_input[192]), .Z(n58283) );
  XOR U58226 ( .A(n58284), .B(n58285), .Z(n1139) );
  AND U58227 ( .A(n58286), .B(n58287), .Z(n58285) );
  XNOR U58228 ( .A(p_input[255]), .B(n58284), .Z(n58287) );
  XOR U58229 ( .A(n58284), .B(p_input[223]), .Z(n58286) );
  XOR U58230 ( .A(n58288), .B(n58289), .Z(n58284) );
  AND U58231 ( .A(n58290), .B(n58291), .Z(n58289) );
  XNOR U58232 ( .A(p_input[254]), .B(n58288), .Z(n58291) );
  XOR U58233 ( .A(n58288), .B(p_input[222]), .Z(n58290) );
  XOR U58234 ( .A(n58292), .B(n58293), .Z(n58288) );
  AND U58235 ( .A(n58294), .B(n58295), .Z(n58293) );
  XNOR U58236 ( .A(p_input[253]), .B(n58292), .Z(n58295) );
  XOR U58237 ( .A(n58292), .B(p_input[221]), .Z(n58294) );
  XOR U58238 ( .A(n58296), .B(n58297), .Z(n58292) );
  AND U58239 ( .A(n58298), .B(n58299), .Z(n58297) );
  XNOR U58240 ( .A(p_input[252]), .B(n58296), .Z(n58299) );
  XOR U58241 ( .A(n58296), .B(p_input[220]), .Z(n58298) );
  XOR U58242 ( .A(n58300), .B(n58301), .Z(n58296) );
  AND U58243 ( .A(n58302), .B(n58303), .Z(n58301) );
  XNOR U58244 ( .A(p_input[251]), .B(n58300), .Z(n58303) );
  XOR U58245 ( .A(n58300), .B(p_input[219]), .Z(n58302) );
  XOR U58246 ( .A(n58304), .B(n58305), .Z(n58300) );
  AND U58247 ( .A(n58306), .B(n58307), .Z(n58305) );
  XNOR U58248 ( .A(p_input[250]), .B(n58304), .Z(n58307) );
  XOR U58249 ( .A(n58304), .B(p_input[218]), .Z(n58306) );
  XOR U58250 ( .A(n58308), .B(n58309), .Z(n58304) );
  AND U58251 ( .A(n58310), .B(n58311), .Z(n58309) );
  XNOR U58252 ( .A(p_input[249]), .B(n58308), .Z(n58311) );
  XOR U58253 ( .A(n58308), .B(p_input[217]), .Z(n58310) );
  XOR U58254 ( .A(n58312), .B(n58313), .Z(n58308) );
  AND U58255 ( .A(n58314), .B(n58315), .Z(n58313) );
  XNOR U58256 ( .A(p_input[248]), .B(n58312), .Z(n58315) );
  XOR U58257 ( .A(n58312), .B(p_input[216]), .Z(n58314) );
  XOR U58258 ( .A(n58316), .B(n58317), .Z(n58312) );
  AND U58259 ( .A(n58318), .B(n58319), .Z(n58317) );
  XNOR U58260 ( .A(p_input[247]), .B(n58316), .Z(n58319) );
  XOR U58261 ( .A(n58316), .B(p_input[215]), .Z(n58318) );
  XOR U58262 ( .A(n58320), .B(n58321), .Z(n58316) );
  AND U58263 ( .A(n58322), .B(n58323), .Z(n58321) );
  XNOR U58264 ( .A(p_input[246]), .B(n58320), .Z(n58323) );
  XOR U58265 ( .A(n58320), .B(p_input[214]), .Z(n58322) );
  XOR U58266 ( .A(n58324), .B(n58325), .Z(n58320) );
  AND U58267 ( .A(n58326), .B(n58327), .Z(n58325) );
  XNOR U58268 ( .A(p_input[245]), .B(n58324), .Z(n58327) );
  XOR U58269 ( .A(n58324), .B(p_input[213]), .Z(n58326) );
  XOR U58270 ( .A(n58328), .B(n58329), .Z(n58324) );
  AND U58271 ( .A(n58330), .B(n58331), .Z(n58329) );
  XNOR U58272 ( .A(p_input[244]), .B(n58328), .Z(n58331) );
  XOR U58273 ( .A(n58328), .B(p_input[212]), .Z(n58330) );
  XOR U58274 ( .A(n58332), .B(n58333), .Z(n58328) );
  AND U58275 ( .A(n58334), .B(n58335), .Z(n58333) );
  XNOR U58276 ( .A(p_input[243]), .B(n58332), .Z(n58335) );
  XOR U58277 ( .A(n58332), .B(p_input[211]), .Z(n58334) );
  XOR U58278 ( .A(n58336), .B(n58337), .Z(n58332) );
  AND U58279 ( .A(n58338), .B(n58339), .Z(n58337) );
  XNOR U58280 ( .A(p_input[242]), .B(n58336), .Z(n58339) );
  XOR U58281 ( .A(n58336), .B(p_input[210]), .Z(n58338) );
  XOR U58282 ( .A(n58340), .B(n58341), .Z(n58336) );
  AND U58283 ( .A(n58342), .B(n58343), .Z(n58341) );
  XNOR U58284 ( .A(p_input[241]), .B(n58340), .Z(n58343) );
  XOR U58285 ( .A(n58340), .B(p_input[209]), .Z(n58342) );
  XOR U58286 ( .A(n58344), .B(n58345), .Z(n58340) );
  AND U58287 ( .A(n58346), .B(n58347), .Z(n58345) );
  XNOR U58288 ( .A(p_input[240]), .B(n58344), .Z(n58347) );
  XOR U58289 ( .A(n58344), .B(p_input[208]), .Z(n58346) );
  XOR U58290 ( .A(n58348), .B(n58349), .Z(n58344) );
  AND U58291 ( .A(n58350), .B(n58351), .Z(n58349) );
  XNOR U58292 ( .A(p_input[239]), .B(n58348), .Z(n58351) );
  XOR U58293 ( .A(n58348), .B(p_input[207]), .Z(n58350) );
  XOR U58294 ( .A(n58352), .B(n58353), .Z(n58348) );
  AND U58295 ( .A(n58354), .B(n58355), .Z(n58353) );
  XNOR U58296 ( .A(p_input[238]), .B(n58352), .Z(n58355) );
  XOR U58297 ( .A(n58352), .B(p_input[206]), .Z(n58354) );
  XOR U58298 ( .A(n58356), .B(n58357), .Z(n58352) );
  AND U58299 ( .A(n58358), .B(n58359), .Z(n58357) );
  XNOR U58300 ( .A(p_input[237]), .B(n58356), .Z(n58359) );
  XOR U58301 ( .A(n58356), .B(p_input[205]), .Z(n58358) );
  XOR U58302 ( .A(n58360), .B(n58361), .Z(n58356) );
  AND U58303 ( .A(n58362), .B(n58363), .Z(n58361) );
  XNOR U58304 ( .A(p_input[236]), .B(n58360), .Z(n58363) );
  XOR U58305 ( .A(n58360), .B(p_input[204]), .Z(n58362) );
  XOR U58306 ( .A(n58364), .B(n58365), .Z(n58360) );
  AND U58307 ( .A(n58366), .B(n58367), .Z(n58365) );
  XNOR U58308 ( .A(p_input[235]), .B(n58364), .Z(n58367) );
  XOR U58309 ( .A(n58364), .B(p_input[203]), .Z(n58366) );
  XOR U58310 ( .A(n58368), .B(n58369), .Z(n58364) );
  AND U58311 ( .A(n58370), .B(n58371), .Z(n58369) );
  XNOR U58312 ( .A(p_input[234]), .B(n58368), .Z(n58371) );
  XOR U58313 ( .A(n58368), .B(p_input[202]), .Z(n58370) );
  XOR U58314 ( .A(n58372), .B(n58373), .Z(n58368) );
  AND U58315 ( .A(n58374), .B(n58375), .Z(n58373) );
  XNOR U58316 ( .A(p_input[233]), .B(n58372), .Z(n58375) );
  XOR U58317 ( .A(n58372), .B(p_input[201]), .Z(n58374) );
  XOR U58318 ( .A(n58376), .B(n58377), .Z(n58372) );
  AND U58319 ( .A(n58378), .B(n58379), .Z(n58377) );
  XNOR U58320 ( .A(p_input[232]), .B(n58376), .Z(n58379) );
  XOR U58321 ( .A(n58376), .B(p_input[200]), .Z(n58378) );
  XOR U58322 ( .A(n58380), .B(n58381), .Z(n58376) );
  AND U58323 ( .A(n58382), .B(n58383), .Z(n58381) );
  XNOR U58324 ( .A(p_input[231]), .B(n58380), .Z(n58383) );
  XOR U58325 ( .A(n58380), .B(p_input[199]), .Z(n58382) );
  XOR U58326 ( .A(n58384), .B(n58385), .Z(n58380) );
  AND U58327 ( .A(n58386), .B(n58387), .Z(n58385) );
  XNOR U58328 ( .A(p_input[230]), .B(n58384), .Z(n58387) );
  XOR U58329 ( .A(n58384), .B(p_input[198]), .Z(n58386) );
  XOR U58330 ( .A(n58388), .B(n58389), .Z(n58384) );
  AND U58331 ( .A(n58390), .B(n58391), .Z(n58389) );
  XNOR U58332 ( .A(p_input[229]), .B(n58388), .Z(n58391) );
  XOR U58333 ( .A(n58388), .B(p_input[197]), .Z(n58390) );
  XOR U58334 ( .A(n58392), .B(n58393), .Z(n58388) );
  AND U58335 ( .A(n58394), .B(n58395), .Z(n58393) );
  XNOR U58336 ( .A(p_input[228]), .B(n58392), .Z(n58395) );
  XOR U58337 ( .A(n58392), .B(p_input[196]), .Z(n58394) );
  XOR U58338 ( .A(n58396), .B(n58397), .Z(n58392) );
  AND U58339 ( .A(n58398), .B(n58399), .Z(n58397) );
  XNOR U58340 ( .A(p_input[227]), .B(n58396), .Z(n58399) );
  XOR U58341 ( .A(n58396), .B(p_input[195]), .Z(n58398) );
  XOR U58342 ( .A(n58400), .B(n58401), .Z(n58396) );
  AND U58343 ( .A(n58402), .B(n58403), .Z(n58401) );
  XNOR U58344 ( .A(p_input[226]), .B(n58400), .Z(n58403) );
  XOR U58345 ( .A(n58400), .B(p_input[194]), .Z(n58402) );
  XNOR U58346 ( .A(n58404), .B(n58405), .Z(n58400) );
  AND U58347 ( .A(n58406), .B(n58407), .Z(n58405) );
  XOR U58348 ( .A(p_input[225]), .B(n58404), .Z(n58407) );
  XNOR U58349 ( .A(p_input[193]), .B(n58404), .Z(n58406) );
  AND U58350 ( .A(p_input[224]), .B(n58408), .Z(n58404) );
  IV U58351 ( .A(p_input[192]), .Z(n58408) );
  XNOR U58352 ( .A(p_input[128]), .B(n58409), .Z(n58002) );
  AND U58353 ( .A(n1137), .B(n58410), .Z(n58409) );
  XOR U58354 ( .A(p_input[160]), .B(p_input[128]), .Z(n58410) );
  XOR U58355 ( .A(n58411), .B(n58412), .Z(n1137) );
  AND U58356 ( .A(n58413), .B(n58414), .Z(n58412) );
  XNOR U58357 ( .A(p_input[191]), .B(n58411), .Z(n58414) );
  XOR U58358 ( .A(n58411), .B(p_input[159]), .Z(n58413) );
  XOR U58359 ( .A(n58415), .B(n58416), .Z(n58411) );
  AND U58360 ( .A(n58417), .B(n58418), .Z(n58416) );
  XNOR U58361 ( .A(p_input[190]), .B(n58415), .Z(n58418) );
  XNOR U58362 ( .A(n58415), .B(n58017), .Z(n58417) );
  IV U58363 ( .A(p_input[158]), .Z(n58017) );
  XOR U58364 ( .A(n58419), .B(n58420), .Z(n58415) );
  AND U58365 ( .A(n58421), .B(n58422), .Z(n58420) );
  XNOR U58366 ( .A(p_input[189]), .B(n58419), .Z(n58422) );
  XNOR U58367 ( .A(n58419), .B(n58026), .Z(n58421) );
  IV U58368 ( .A(p_input[157]), .Z(n58026) );
  XOR U58369 ( .A(n58423), .B(n58424), .Z(n58419) );
  AND U58370 ( .A(n58425), .B(n58426), .Z(n58424) );
  XNOR U58371 ( .A(p_input[188]), .B(n58423), .Z(n58426) );
  XNOR U58372 ( .A(n58423), .B(n58035), .Z(n58425) );
  IV U58373 ( .A(p_input[156]), .Z(n58035) );
  XOR U58374 ( .A(n58427), .B(n58428), .Z(n58423) );
  AND U58375 ( .A(n58429), .B(n58430), .Z(n58428) );
  XNOR U58376 ( .A(p_input[187]), .B(n58427), .Z(n58430) );
  XNOR U58377 ( .A(n58427), .B(n58044), .Z(n58429) );
  IV U58378 ( .A(p_input[155]), .Z(n58044) );
  XOR U58379 ( .A(n58431), .B(n58432), .Z(n58427) );
  AND U58380 ( .A(n58433), .B(n58434), .Z(n58432) );
  XNOR U58381 ( .A(p_input[186]), .B(n58431), .Z(n58434) );
  XNOR U58382 ( .A(n58431), .B(n58053), .Z(n58433) );
  IV U58383 ( .A(p_input[154]), .Z(n58053) );
  XOR U58384 ( .A(n58435), .B(n58436), .Z(n58431) );
  AND U58385 ( .A(n58437), .B(n58438), .Z(n58436) );
  XNOR U58386 ( .A(p_input[185]), .B(n58435), .Z(n58438) );
  XNOR U58387 ( .A(n58435), .B(n58062), .Z(n58437) );
  IV U58388 ( .A(p_input[153]), .Z(n58062) );
  XOR U58389 ( .A(n58439), .B(n58440), .Z(n58435) );
  AND U58390 ( .A(n58441), .B(n58442), .Z(n58440) );
  XNOR U58391 ( .A(p_input[184]), .B(n58439), .Z(n58442) );
  XNOR U58392 ( .A(n58439), .B(n58071), .Z(n58441) );
  IV U58393 ( .A(p_input[152]), .Z(n58071) );
  XOR U58394 ( .A(n58443), .B(n58444), .Z(n58439) );
  AND U58395 ( .A(n58445), .B(n58446), .Z(n58444) );
  XNOR U58396 ( .A(p_input[183]), .B(n58443), .Z(n58446) );
  XNOR U58397 ( .A(n58443), .B(n58080), .Z(n58445) );
  IV U58398 ( .A(p_input[151]), .Z(n58080) );
  XOR U58399 ( .A(n58447), .B(n58448), .Z(n58443) );
  AND U58400 ( .A(n58449), .B(n58450), .Z(n58448) );
  XNOR U58401 ( .A(p_input[182]), .B(n58447), .Z(n58450) );
  XNOR U58402 ( .A(n58447), .B(n58089), .Z(n58449) );
  IV U58403 ( .A(p_input[150]), .Z(n58089) );
  XOR U58404 ( .A(n58451), .B(n58452), .Z(n58447) );
  AND U58405 ( .A(n58453), .B(n58454), .Z(n58452) );
  XNOR U58406 ( .A(p_input[181]), .B(n58451), .Z(n58454) );
  XNOR U58407 ( .A(n58451), .B(n58098), .Z(n58453) );
  IV U58408 ( .A(p_input[149]), .Z(n58098) );
  XOR U58409 ( .A(n58455), .B(n58456), .Z(n58451) );
  AND U58410 ( .A(n58457), .B(n58458), .Z(n58456) );
  XNOR U58411 ( .A(p_input[180]), .B(n58455), .Z(n58458) );
  XNOR U58412 ( .A(n58455), .B(n58107), .Z(n58457) );
  IV U58413 ( .A(p_input[148]), .Z(n58107) );
  XOR U58414 ( .A(n58459), .B(n58460), .Z(n58455) );
  AND U58415 ( .A(n58461), .B(n58462), .Z(n58460) );
  XNOR U58416 ( .A(p_input[179]), .B(n58459), .Z(n58462) );
  XNOR U58417 ( .A(n58459), .B(n58116), .Z(n58461) );
  IV U58418 ( .A(p_input[147]), .Z(n58116) );
  XOR U58419 ( .A(n58463), .B(n58464), .Z(n58459) );
  AND U58420 ( .A(n58465), .B(n58466), .Z(n58464) );
  XNOR U58421 ( .A(p_input[178]), .B(n58463), .Z(n58466) );
  XNOR U58422 ( .A(n58463), .B(n58125), .Z(n58465) );
  IV U58423 ( .A(p_input[146]), .Z(n58125) );
  XOR U58424 ( .A(n58467), .B(n58468), .Z(n58463) );
  AND U58425 ( .A(n58469), .B(n58470), .Z(n58468) );
  XNOR U58426 ( .A(p_input[177]), .B(n58467), .Z(n58470) );
  XNOR U58427 ( .A(n58467), .B(n58134), .Z(n58469) );
  IV U58428 ( .A(p_input[145]), .Z(n58134) );
  XOR U58429 ( .A(n58471), .B(n58472), .Z(n58467) );
  AND U58430 ( .A(n58473), .B(n58474), .Z(n58472) );
  XNOR U58431 ( .A(p_input[176]), .B(n58471), .Z(n58474) );
  XNOR U58432 ( .A(n58471), .B(n58143), .Z(n58473) );
  IV U58433 ( .A(p_input[144]), .Z(n58143) );
  XOR U58434 ( .A(n58475), .B(n58476), .Z(n58471) );
  AND U58435 ( .A(n58477), .B(n58478), .Z(n58476) );
  XNOR U58436 ( .A(p_input[175]), .B(n58475), .Z(n58478) );
  XNOR U58437 ( .A(n58475), .B(n58152), .Z(n58477) );
  IV U58438 ( .A(p_input[143]), .Z(n58152) );
  XOR U58439 ( .A(n58479), .B(n58480), .Z(n58475) );
  AND U58440 ( .A(n58481), .B(n58482), .Z(n58480) );
  XNOR U58441 ( .A(p_input[174]), .B(n58479), .Z(n58482) );
  XNOR U58442 ( .A(n58479), .B(n58161), .Z(n58481) );
  IV U58443 ( .A(p_input[142]), .Z(n58161) );
  XOR U58444 ( .A(n58483), .B(n58484), .Z(n58479) );
  AND U58445 ( .A(n58485), .B(n58486), .Z(n58484) );
  XNOR U58446 ( .A(p_input[173]), .B(n58483), .Z(n58486) );
  XNOR U58447 ( .A(n58483), .B(n58170), .Z(n58485) );
  IV U58448 ( .A(p_input[141]), .Z(n58170) );
  XOR U58449 ( .A(n58487), .B(n58488), .Z(n58483) );
  AND U58450 ( .A(n58489), .B(n58490), .Z(n58488) );
  XNOR U58451 ( .A(p_input[172]), .B(n58487), .Z(n58490) );
  XNOR U58452 ( .A(n58487), .B(n58179), .Z(n58489) );
  IV U58453 ( .A(p_input[140]), .Z(n58179) );
  XOR U58454 ( .A(n58491), .B(n58492), .Z(n58487) );
  AND U58455 ( .A(n58493), .B(n58494), .Z(n58492) );
  XNOR U58456 ( .A(p_input[171]), .B(n58491), .Z(n58494) );
  XNOR U58457 ( .A(n58491), .B(n58188), .Z(n58493) );
  IV U58458 ( .A(p_input[139]), .Z(n58188) );
  XOR U58459 ( .A(n58495), .B(n58496), .Z(n58491) );
  AND U58460 ( .A(n58497), .B(n58498), .Z(n58496) );
  XNOR U58461 ( .A(p_input[170]), .B(n58495), .Z(n58498) );
  XNOR U58462 ( .A(n58495), .B(n58197), .Z(n58497) );
  IV U58463 ( .A(p_input[138]), .Z(n58197) );
  XOR U58464 ( .A(n58499), .B(n58500), .Z(n58495) );
  AND U58465 ( .A(n58501), .B(n58502), .Z(n58500) );
  XNOR U58466 ( .A(p_input[169]), .B(n58499), .Z(n58502) );
  XNOR U58467 ( .A(n58499), .B(n58206), .Z(n58501) );
  IV U58468 ( .A(p_input[137]), .Z(n58206) );
  XOR U58469 ( .A(n58503), .B(n58504), .Z(n58499) );
  AND U58470 ( .A(n58505), .B(n58506), .Z(n58504) );
  XNOR U58471 ( .A(p_input[168]), .B(n58503), .Z(n58506) );
  XNOR U58472 ( .A(n58503), .B(n58215), .Z(n58505) );
  IV U58473 ( .A(p_input[136]), .Z(n58215) );
  XOR U58474 ( .A(n58507), .B(n58508), .Z(n58503) );
  AND U58475 ( .A(n58509), .B(n58510), .Z(n58508) );
  XNOR U58476 ( .A(p_input[167]), .B(n58507), .Z(n58510) );
  XNOR U58477 ( .A(n58507), .B(n58224), .Z(n58509) );
  IV U58478 ( .A(p_input[135]), .Z(n58224) );
  XOR U58479 ( .A(n58511), .B(n58512), .Z(n58507) );
  AND U58480 ( .A(n58513), .B(n58514), .Z(n58512) );
  XNOR U58481 ( .A(p_input[166]), .B(n58511), .Z(n58514) );
  XNOR U58482 ( .A(n58511), .B(n58233), .Z(n58513) );
  IV U58483 ( .A(p_input[134]), .Z(n58233) );
  XOR U58484 ( .A(n58515), .B(n58516), .Z(n58511) );
  AND U58485 ( .A(n58517), .B(n58518), .Z(n58516) );
  XNOR U58486 ( .A(p_input[165]), .B(n58515), .Z(n58518) );
  XNOR U58487 ( .A(n58515), .B(n58242), .Z(n58517) );
  IV U58488 ( .A(p_input[133]), .Z(n58242) );
  XOR U58489 ( .A(n58519), .B(n58520), .Z(n58515) );
  AND U58490 ( .A(n58521), .B(n58522), .Z(n58520) );
  XNOR U58491 ( .A(p_input[164]), .B(n58519), .Z(n58522) );
  XNOR U58492 ( .A(n58519), .B(n58251), .Z(n58521) );
  IV U58493 ( .A(p_input[132]), .Z(n58251) );
  XOR U58494 ( .A(n58523), .B(n58524), .Z(n58519) );
  AND U58495 ( .A(n58525), .B(n58526), .Z(n58524) );
  XNOR U58496 ( .A(p_input[163]), .B(n58523), .Z(n58526) );
  XNOR U58497 ( .A(n58523), .B(n58260), .Z(n58525) );
  IV U58498 ( .A(p_input[131]), .Z(n58260) );
  XOR U58499 ( .A(n58527), .B(n58528), .Z(n58523) );
  AND U58500 ( .A(n58529), .B(n58530), .Z(n58528) );
  XNOR U58501 ( .A(p_input[162]), .B(n58527), .Z(n58530) );
  XNOR U58502 ( .A(n58527), .B(n58269), .Z(n58529) );
  IV U58503 ( .A(p_input[130]), .Z(n58269) );
  XNOR U58504 ( .A(n58531), .B(n58532), .Z(n58527) );
  AND U58505 ( .A(n58533), .B(n58534), .Z(n58532) );
  XOR U58506 ( .A(p_input[161]), .B(n58531), .Z(n58534) );
  XNOR U58507 ( .A(p_input[129]), .B(n58531), .Z(n58533) );
  AND U58508 ( .A(p_input[160]), .B(n58535), .Z(n58531) );
  IV U58509 ( .A(p_input[128]), .Z(n58535) );
  XOR U58510 ( .A(n58536), .B(n58537), .Z(n57625) );
  AND U58511 ( .A(n664), .B(n58538), .Z(n58537) );
  XNOR U58512 ( .A(n58539), .B(n58536), .Z(n58538) );
  XOR U58513 ( .A(n58540), .B(n58541), .Z(n664) );
  AND U58514 ( .A(n58542), .B(n58543), .Z(n58541) );
  XNOR U58515 ( .A(n57640), .B(n58540), .Z(n58543) );
  AND U58516 ( .A(p_input[95]), .B(p_input[127]), .Z(n57640) );
  XNOR U58517 ( .A(n58540), .B(n57637), .Z(n58542) );
  IV U58518 ( .A(n58544), .Z(n57637) );
  AND U58519 ( .A(p_input[31]), .B(p_input[63]), .Z(n58544) );
  XOR U58520 ( .A(n58545), .B(n58546), .Z(n58540) );
  AND U58521 ( .A(n58547), .B(n58548), .Z(n58546) );
  XOR U58522 ( .A(n58545), .B(n57652), .Z(n58548) );
  XNOR U58523 ( .A(p_input[94]), .B(n58549), .Z(n57652) );
  AND U58524 ( .A(n1147), .B(n58550), .Z(n58549) );
  XOR U58525 ( .A(p_input[94]), .B(p_input[126]), .Z(n58550) );
  XNOR U58526 ( .A(n57649), .B(n58545), .Z(n58547) );
  XOR U58527 ( .A(n58551), .B(n58552), .Z(n57649) );
  AND U58528 ( .A(n1144), .B(n58553), .Z(n58552) );
  XOR U58529 ( .A(p_input[62]), .B(p_input[30]), .Z(n58553) );
  XOR U58530 ( .A(n58554), .B(n58555), .Z(n58545) );
  AND U58531 ( .A(n58556), .B(n58557), .Z(n58555) );
  XOR U58532 ( .A(n58554), .B(n57664), .Z(n58557) );
  XNOR U58533 ( .A(p_input[93]), .B(n58558), .Z(n57664) );
  AND U58534 ( .A(n1147), .B(n58559), .Z(n58558) );
  XOR U58535 ( .A(p_input[93]), .B(p_input[125]), .Z(n58559) );
  XNOR U58536 ( .A(n57661), .B(n58554), .Z(n58556) );
  XOR U58537 ( .A(n58560), .B(n58561), .Z(n57661) );
  AND U58538 ( .A(n1144), .B(n58562), .Z(n58561) );
  XOR U58539 ( .A(p_input[61]), .B(p_input[29]), .Z(n58562) );
  XOR U58540 ( .A(n58563), .B(n58564), .Z(n58554) );
  AND U58541 ( .A(n58565), .B(n58566), .Z(n58564) );
  XOR U58542 ( .A(n58563), .B(n57676), .Z(n58566) );
  XNOR U58543 ( .A(p_input[92]), .B(n58567), .Z(n57676) );
  AND U58544 ( .A(n1147), .B(n58568), .Z(n58567) );
  XOR U58545 ( .A(p_input[92]), .B(p_input[124]), .Z(n58568) );
  XNOR U58546 ( .A(n57673), .B(n58563), .Z(n58565) );
  XOR U58547 ( .A(n58569), .B(n58570), .Z(n57673) );
  AND U58548 ( .A(n1144), .B(n58571), .Z(n58570) );
  XOR U58549 ( .A(p_input[60]), .B(p_input[28]), .Z(n58571) );
  XOR U58550 ( .A(n58572), .B(n58573), .Z(n58563) );
  AND U58551 ( .A(n58574), .B(n58575), .Z(n58573) );
  XOR U58552 ( .A(n58572), .B(n57688), .Z(n58575) );
  XNOR U58553 ( .A(p_input[91]), .B(n58576), .Z(n57688) );
  AND U58554 ( .A(n1147), .B(n58577), .Z(n58576) );
  XOR U58555 ( .A(p_input[91]), .B(p_input[123]), .Z(n58577) );
  XNOR U58556 ( .A(n57685), .B(n58572), .Z(n58574) );
  XOR U58557 ( .A(n58578), .B(n58579), .Z(n57685) );
  AND U58558 ( .A(n1144), .B(n58580), .Z(n58579) );
  XOR U58559 ( .A(p_input[59]), .B(p_input[27]), .Z(n58580) );
  XOR U58560 ( .A(n58581), .B(n58582), .Z(n58572) );
  AND U58561 ( .A(n58583), .B(n58584), .Z(n58582) );
  XOR U58562 ( .A(n58581), .B(n57700), .Z(n58584) );
  XNOR U58563 ( .A(p_input[90]), .B(n58585), .Z(n57700) );
  AND U58564 ( .A(n1147), .B(n58586), .Z(n58585) );
  XOR U58565 ( .A(p_input[90]), .B(p_input[122]), .Z(n58586) );
  XNOR U58566 ( .A(n57697), .B(n58581), .Z(n58583) );
  XOR U58567 ( .A(n58587), .B(n58588), .Z(n57697) );
  AND U58568 ( .A(n1144), .B(n58589), .Z(n58588) );
  XOR U58569 ( .A(p_input[58]), .B(p_input[26]), .Z(n58589) );
  XOR U58570 ( .A(n58590), .B(n58591), .Z(n58581) );
  AND U58571 ( .A(n58592), .B(n58593), .Z(n58591) );
  XOR U58572 ( .A(n58590), .B(n57712), .Z(n58593) );
  XNOR U58573 ( .A(p_input[89]), .B(n58594), .Z(n57712) );
  AND U58574 ( .A(n1147), .B(n58595), .Z(n58594) );
  XOR U58575 ( .A(p_input[89]), .B(p_input[121]), .Z(n58595) );
  XNOR U58576 ( .A(n57709), .B(n58590), .Z(n58592) );
  XOR U58577 ( .A(n58596), .B(n58597), .Z(n57709) );
  AND U58578 ( .A(n1144), .B(n58598), .Z(n58597) );
  XOR U58579 ( .A(p_input[57]), .B(p_input[25]), .Z(n58598) );
  XOR U58580 ( .A(n58599), .B(n58600), .Z(n58590) );
  AND U58581 ( .A(n58601), .B(n58602), .Z(n58600) );
  XOR U58582 ( .A(n58599), .B(n57724), .Z(n58602) );
  XNOR U58583 ( .A(p_input[88]), .B(n58603), .Z(n57724) );
  AND U58584 ( .A(n1147), .B(n58604), .Z(n58603) );
  XOR U58585 ( .A(p_input[88]), .B(p_input[120]), .Z(n58604) );
  XNOR U58586 ( .A(n57721), .B(n58599), .Z(n58601) );
  XOR U58587 ( .A(n58605), .B(n58606), .Z(n57721) );
  AND U58588 ( .A(n1144), .B(n58607), .Z(n58606) );
  XOR U58589 ( .A(p_input[56]), .B(p_input[24]), .Z(n58607) );
  XOR U58590 ( .A(n58608), .B(n58609), .Z(n58599) );
  AND U58591 ( .A(n58610), .B(n58611), .Z(n58609) );
  XOR U58592 ( .A(n58608), .B(n57736), .Z(n58611) );
  XNOR U58593 ( .A(p_input[87]), .B(n58612), .Z(n57736) );
  AND U58594 ( .A(n1147), .B(n58613), .Z(n58612) );
  XOR U58595 ( .A(p_input[87]), .B(p_input[119]), .Z(n58613) );
  XNOR U58596 ( .A(n57733), .B(n58608), .Z(n58610) );
  XOR U58597 ( .A(n58614), .B(n58615), .Z(n57733) );
  AND U58598 ( .A(n1144), .B(n58616), .Z(n58615) );
  XOR U58599 ( .A(p_input[55]), .B(p_input[23]), .Z(n58616) );
  XOR U58600 ( .A(n58617), .B(n58618), .Z(n58608) );
  AND U58601 ( .A(n58619), .B(n58620), .Z(n58618) );
  XOR U58602 ( .A(n58617), .B(n57748), .Z(n58620) );
  XNOR U58603 ( .A(p_input[86]), .B(n58621), .Z(n57748) );
  AND U58604 ( .A(n1147), .B(n58622), .Z(n58621) );
  XOR U58605 ( .A(p_input[86]), .B(p_input[118]), .Z(n58622) );
  XNOR U58606 ( .A(n57745), .B(n58617), .Z(n58619) );
  XOR U58607 ( .A(n58623), .B(n58624), .Z(n57745) );
  AND U58608 ( .A(n1144), .B(n58625), .Z(n58624) );
  XOR U58609 ( .A(p_input[54]), .B(p_input[22]), .Z(n58625) );
  XOR U58610 ( .A(n58626), .B(n58627), .Z(n58617) );
  AND U58611 ( .A(n58628), .B(n58629), .Z(n58627) );
  XOR U58612 ( .A(n58626), .B(n57760), .Z(n58629) );
  XNOR U58613 ( .A(p_input[85]), .B(n58630), .Z(n57760) );
  AND U58614 ( .A(n1147), .B(n58631), .Z(n58630) );
  XOR U58615 ( .A(p_input[85]), .B(p_input[117]), .Z(n58631) );
  XNOR U58616 ( .A(n57757), .B(n58626), .Z(n58628) );
  XOR U58617 ( .A(n58632), .B(n58633), .Z(n57757) );
  AND U58618 ( .A(n1144), .B(n58634), .Z(n58633) );
  XOR U58619 ( .A(p_input[53]), .B(p_input[21]), .Z(n58634) );
  XOR U58620 ( .A(n58635), .B(n58636), .Z(n58626) );
  AND U58621 ( .A(n58637), .B(n58638), .Z(n58636) );
  XOR U58622 ( .A(n58635), .B(n57772), .Z(n58638) );
  XNOR U58623 ( .A(p_input[84]), .B(n58639), .Z(n57772) );
  AND U58624 ( .A(n1147), .B(n58640), .Z(n58639) );
  XOR U58625 ( .A(p_input[84]), .B(p_input[116]), .Z(n58640) );
  XNOR U58626 ( .A(n57769), .B(n58635), .Z(n58637) );
  XOR U58627 ( .A(n58641), .B(n58642), .Z(n57769) );
  AND U58628 ( .A(n1144), .B(n58643), .Z(n58642) );
  XOR U58629 ( .A(p_input[52]), .B(p_input[20]), .Z(n58643) );
  XOR U58630 ( .A(n58644), .B(n58645), .Z(n58635) );
  AND U58631 ( .A(n58646), .B(n58647), .Z(n58645) );
  XOR U58632 ( .A(n58644), .B(n57784), .Z(n58647) );
  XNOR U58633 ( .A(p_input[83]), .B(n58648), .Z(n57784) );
  AND U58634 ( .A(n1147), .B(n58649), .Z(n58648) );
  XOR U58635 ( .A(p_input[83]), .B(p_input[115]), .Z(n58649) );
  XNOR U58636 ( .A(n57781), .B(n58644), .Z(n58646) );
  XOR U58637 ( .A(n58650), .B(n58651), .Z(n57781) );
  AND U58638 ( .A(n1144), .B(n58652), .Z(n58651) );
  XOR U58639 ( .A(p_input[51]), .B(p_input[19]), .Z(n58652) );
  XOR U58640 ( .A(n58653), .B(n58654), .Z(n58644) );
  AND U58641 ( .A(n58655), .B(n58656), .Z(n58654) );
  XOR U58642 ( .A(n58653), .B(n57796), .Z(n58656) );
  XNOR U58643 ( .A(p_input[82]), .B(n58657), .Z(n57796) );
  AND U58644 ( .A(n1147), .B(n58658), .Z(n58657) );
  XOR U58645 ( .A(p_input[82]), .B(p_input[114]), .Z(n58658) );
  XNOR U58646 ( .A(n57793), .B(n58653), .Z(n58655) );
  XOR U58647 ( .A(n58659), .B(n58660), .Z(n57793) );
  AND U58648 ( .A(n1144), .B(n58661), .Z(n58660) );
  XOR U58649 ( .A(p_input[50]), .B(p_input[18]), .Z(n58661) );
  XOR U58650 ( .A(n58662), .B(n58663), .Z(n58653) );
  AND U58651 ( .A(n58664), .B(n58665), .Z(n58663) );
  XOR U58652 ( .A(n58662), .B(n57808), .Z(n58665) );
  XNOR U58653 ( .A(p_input[81]), .B(n58666), .Z(n57808) );
  AND U58654 ( .A(n1147), .B(n58667), .Z(n58666) );
  XOR U58655 ( .A(p_input[81]), .B(p_input[113]), .Z(n58667) );
  XNOR U58656 ( .A(n57805), .B(n58662), .Z(n58664) );
  XOR U58657 ( .A(n58668), .B(n58669), .Z(n57805) );
  AND U58658 ( .A(n1144), .B(n58670), .Z(n58669) );
  XOR U58659 ( .A(p_input[49]), .B(p_input[17]), .Z(n58670) );
  XOR U58660 ( .A(n58671), .B(n58672), .Z(n58662) );
  AND U58661 ( .A(n58673), .B(n58674), .Z(n58672) );
  XOR U58662 ( .A(n58671), .B(n57820), .Z(n58674) );
  XNOR U58663 ( .A(p_input[80]), .B(n58675), .Z(n57820) );
  AND U58664 ( .A(n1147), .B(n58676), .Z(n58675) );
  XOR U58665 ( .A(p_input[80]), .B(p_input[112]), .Z(n58676) );
  XNOR U58666 ( .A(n57817), .B(n58671), .Z(n58673) );
  XOR U58667 ( .A(n58677), .B(n58678), .Z(n57817) );
  AND U58668 ( .A(n1144), .B(n58679), .Z(n58678) );
  XOR U58669 ( .A(p_input[48]), .B(p_input[16]), .Z(n58679) );
  XOR U58670 ( .A(n58680), .B(n58681), .Z(n58671) );
  AND U58671 ( .A(n58682), .B(n58683), .Z(n58681) );
  XOR U58672 ( .A(n58680), .B(n57832), .Z(n58683) );
  XNOR U58673 ( .A(p_input[79]), .B(n58684), .Z(n57832) );
  AND U58674 ( .A(n1147), .B(n58685), .Z(n58684) );
  XOR U58675 ( .A(p_input[79]), .B(p_input[111]), .Z(n58685) );
  XNOR U58676 ( .A(n57829), .B(n58680), .Z(n58682) );
  XOR U58677 ( .A(n58686), .B(n58687), .Z(n57829) );
  AND U58678 ( .A(n1144), .B(n58688), .Z(n58687) );
  XOR U58679 ( .A(p_input[47]), .B(p_input[15]), .Z(n58688) );
  XOR U58680 ( .A(n58689), .B(n58690), .Z(n58680) );
  AND U58681 ( .A(n58691), .B(n58692), .Z(n58690) );
  XOR U58682 ( .A(n58689), .B(n57844), .Z(n58692) );
  XNOR U58683 ( .A(p_input[78]), .B(n58693), .Z(n57844) );
  AND U58684 ( .A(n1147), .B(n58694), .Z(n58693) );
  XOR U58685 ( .A(p_input[78]), .B(p_input[110]), .Z(n58694) );
  XNOR U58686 ( .A(n57841), .B(n58689), .Z(n58691) );
  XOR U58687 ( .A(n58695), .B(n58696), .Z(n57841) );
  AND U58688 ( .A(n1144), .B(n58697), .Z(n58696) );
  XOR U58689 ( .A(p_input[46]), .B(p_input[14]), .Z(n58697) );
  XOR U58690 ( .A(n58698), .B(n58699), .Z(n58689) );
  AND U58691 ( .A(n58700), .B(n58701), .Z(n58699) );
  XOR U58692 ( .A(n58698), .B(n57856), .Z(n58701) );
  XNOR U58693 ( .A(p_input[77]), .B(n58702), .Z(n57856) );
  AND U58694 ( .A(n1147), .B(n58703), .Z(n58702) );
  XOR U58695 ( .A(p_input[77]), .B(p_input[109]), .Z(n58703) );
  XNOR U58696 ( .A(n57853), .B(n58698), .Z(n58700) );
  XOR U58697 ( .A(n58704), .B(n58705), .Z(n57853) );
  AND U58698 ( .A(n1144), .B(n58706), .Z(n58705) );
  XOR U58699 ( .A(p_input[45]), .B(p_input[13]), .Z(n58706) );
  XOR U58700 ( .A(n58707), .B(n58708), .Z(n58698) );
  AND U58701 ( .A(n58709), .B(n58710), .Z(n58708) );
  XOR U58702 ( .A(n58707), .B(n57868), .Z(n58710) );
  XNOR U58703 ( .A(p_input[76]), .B(n58711), .Z(n57868) );
  AND U58704 ( .A(n1147), .B(n58712), .Z(n58711) );
  XOR U58705 ( .A(p_input[76]), .B(p_input[108]), .Z(n58712) );
  XNOR U58706 ( .A(n57865), .B(n58707), .Z(n58709) );
  XOR U58707 ( .A(n58713), .B(n58714), .Z(n57865) );
  AND U58708 ( .A(n1144), .B(n58715), .Z(n58714) );
  XOR U58709 ( .A(p_input[44]), .B(p_input[12]), .Z(n58715) );
  XOR U58710 ( .A(n58716), .B(n58717), .Z(n58707) );
  AND U58711 ( .A(n58718), .B(n58719), .Z(n58717) );
  XOR U58712 ( .A(n58716), .B(n57880), .Z(n58719) );
  XNOR U58713 ( .A(p_input[75]), .B(n58720), .Z(n57880) );
  AND U58714 ( .A(n1147), .B(n58721), .Z(n58720) );
  XOR U58715 ( .A(p_input[75]), .B(p_input[107]), .Z(n58721) );
  XNOR U58716 ( .A(n57877), .B(n58716), .Z(n58718) );
  XOR U58717 ( .A(n58722), .B(n58723), .Z(n57877) );
  AND U58718 ( .A(n1144), .B(n58724), .Z(n58723) );
  XOR U58719 ( .A(p_input[43]), .B(p_input[11]), .Z(n58724) );
  XOR U58720 ( .A(n58725), .B(n58726), .Z(n58716) );
  AND U58721 ( .A(n58727), .B(n58728), .Z(n58726) );
  XOR U58722 ( .A(n58725), .B(n57892), .Z(n58728) );
  XNOR U58723 ( .A(p_input[74]), .B(n58729), .Z(n57892) );
  AND U58724 ( .A(n1147), .B(n58730), .Z(n58729) );
  XOR U58725 ( .A(p_input[74]), .B(p_input[106]), .Z(n58730) );
  XNOR U58726 ( .A(n57889), .B(n58725), .Z(n58727) );
  XOR U58727 ( .A(n58731), .B(n58732), .Z(n57889) );
  AND U58728 ( .A(n1144), .B(n58733), .Z(n58732) );
  XOR U58729 ( .A(p_input[42]), .B(p_input[10]), .Z(n58733) );
  XOR U58730 ( .A(n58734), .B(n58735), .Z(n58725) );
  AND U58731 ( .A(n58736), .B(n58737), .Z(n58735) );
  XOR U58732 ( .A(n58734), .B(n57904), .Z(n58737) );
  XNOR U58733 ( .A(p_input[73]), .B(n58738), .Z(n57904) );
  AND U58734 ( .A(n1147), .B(n58739), .Z(n58738) );
  XOR U58735 ( .A(p_input[73]), .B(p_input[105]), .Z(n58739) );
  XNOR U58736 ( .A(n57901), .B(n58734), .Z(n58736) );
  XOR U58737 ( .A(n58740), .B(n58741), .Z(n57901) );
  AND U58738 ( .A(n1144), .B(n58742), .Z(n58741) );
  XOR U58739 ( .A(p_input[9]), .B(p_input[41]), .Z(n58742) );
  XOR U58740 ( .A(n58743), .B(n58744), .Z(n58734) );
  AND U58741 ( .A(n58745), .B(n58746), .Z(n58744) );
  XOR U58742 ( .A(n58743), .B(n57916), .Z(n58746) );
  XNOR U58743 ( .A(p_input[72]), .B(n58747), .Z(n57916) );
  AND U58744 ( .A(n1147), .B(n58748), .Z(n58747) );
  XOR U58745 ( .A(p_input[72]), .B(p_input[104]), .Z(n58748) );
  XNOR U58746 ( .A(n57913), .B(n58743), .Z(n58745) );
  XOR U58747 ( .A(n58749), .B(n58750), .Z(n57913) );
  AND U58748 ( .A(n1144), .B(n58751), .Z(n58750) );
  XOR U58749 ( .A(p_input[8]), .B(p_input[40]), .Z(n58751) );
  XOR U58750 ( .A(n58752), .B(n58753), .Z(n58743) );
  AND U58751 ( .A(n58754), .B(n58755), .Z(n58753) );
  XOR U58752 ( .A(n58752), .B(n57928), .Z(n58755) );
  XNOR U58753 ( .A(p_input[71]), .B(n58756), .Z(n57928) );
  AND U58754 ( .A(n1147), .B(n58757), .Z(n58756) );
  XOR U58755 ( .A(p_input[71]), .B(p_input[103]), .Z(n58757) );
  XNOR U58756 ( .A(n57925), .B(n58752), .Z(n58754) );
  XOR U58757 ( .A(n58758), .B(n58759), .Z(n57925) );
  AND U58758 ( .A(n1144), .B(n58760), .Z(n58759) );
  XOR U58759 ( .A(p_input[7]), .B(p_input[39]), .Z(n58760) );
  XOR U58760 ( .A(n58761), .B(n58762), .Z(n58752) );
  AND U58761 ( .A(n58763), .B(n58764), .Z(n58762) );
  XOR U58762 ( .A(n58761), .B(n57940), .Z(n58764) );
  XNOR U58763 ( .A(p_input[70]), .B(n58765), .Z(n57940) );
  AND U58764 ( .A(n1147), .B(n58766), .Z(n58765) );
  XOR U58765 ( .A(p_input[70]), .B(p_input[102]), .Z(n58766) );
  XNOR U58766 ( .A(n57937), .B(n58761), .Z(n58763) );
  XOR U58767 ( .A(n58767), .B(n58768), .Z(n57937) );
  AND U58768 ( .A(n1144), .B(n58769), .Z(n58768) );
  XOR U58769 ( .A(p_input[6]), .B(p_input[38]), .Z(n58769) );
  XOR U58770 ( .A(n58770), .B(n58771), .Z(n58761) );
  AND U58771 ( .A(n58772), .B(n58773), .Z(n58771) );
  XOR U58772 ( .A(n58770), .B(n57952), .Z(n58773) );
  XNOR U58773 ( .A(p_input[69]), .B(n58774), .Z(n57952) );
  AND U58774 ( .A(n1147), .B(n58775), .Z(n58774) );
  XOR U58775 ( .A(p_input[69]), .B(p_input[101]), .Z(n58775) );
  XNOR U58776 ( .A(n57949), .B(n58770), .Z(n58772) );
  XOR U58777 ( .A(n58776), .B(n58777), .Z(n57949) );
  AND U58778 ( .A(n1144), .B(n58778), .Z(n58777) );
  XOR U58779 ( .A(p_input[5]), .B(p_input[37]), .Z(n58778) );
  XOR U58780 ( .A(n58779), .B(n58780), .Z(n58770) );
  AND U58781 ( .A(n58781), .B(n58782), .Z(n58780) );
  XOR U58782 ( .A(n58779), .B(n57964), .Z(n58782) );
  XNOR U58783 ( .A(p_input[68]), .B(n58783), .Z(n57964) );
  AND U58784 ( .A(n1147), .B(n58784), .Z(n58783) );
  XOR U58785 ( .A(p_input[68]), .B(p_input[100]), .Z(n58784) );
  XNOR U58786 ( .A(n57961), .B(n58779), .Z(n58781) );
  XOR U58787 ( .A(n58785), .B(n58786), .Z(n57961) );
  AND U58788 ( .A(n1144), .B(n58787), .Z(n58786) );
  XOR U58789 ( .A(p_input[4]), .B(p_input[36]), .Z(n58787) );
  XOR U58790 ( .A(n58788), .B(n58789), .Z(n58779) );
  AND U58791 ( .A(n58790), .B(n58791), .Z(n58789) );
  XOR U58792 ( .A(n58788), .B(n57976), .Z(n58791) );
  XNOR U58793 ( .A(p_input[67]), .B(n58792), .Z(n57976) );
  AND U58794 ( .A(n1147), .B(n58793), .Z(n58792) );
  XOR U58795 ( .A(p_input[99]), .B(p_input[67]), .Z(n58793) );
  XNOR U58796 ( .A(n57973), .B(n58788), .Z(n58790) );
  XOR U58797 ( .A(n58794), .B(n58795), .Z(n57973) );
  AND U58798 ( .A(n1144), .B(n58796), .Z(n58795) );
  XOR U58799 ( .A(p_input[3]), .B(p_input[35]), .Z(n58796) );
  XOR U58800 ( .A(n58797), .B(n58798), .Z(n58788) );
  AND U58801 ( .A(n58799), .B(n58800), .Z(n58798) );
  XOR U58802 ( .A(n58797), .B(n57988), .Z(n58800) );
  XNOR U58803 ( .A(p_input[66]), .B(n58801), .Z(n57988) );
  AND U58804 ( .A(n1147), .B(n58802), .Z(n58801) );
  XOR U58805 ( .A(p_input[98]), .B(p_input[66]), .Z(n58802) );
  XNOR U58806 ( .A(n57985), .B(n58797), .Z(n58799) );
  XOR U58807 ( .A(n58803), .B(n58804), .Z(n57985) );
  AND U58808 ( .A(n1144), .B(n58805), .Z(n58804) );
  XOR U58809 ( .A(p_input[34]), .B(p_input[2]), .Z(n58805) );
  XOR U58810 ( .A(n58806), .B(n58807), .Z(n58797) );
  AND U58811 ( .A(n58808), .B(n58809), .Z(n58807) );
  XNOR U58812 ( .A(n58810), .B(n58001), .Z(n58809) );
  XNOR U58813 ( .A(p_input[65]), .B(n58811), .Z(n58001) );
  AND U58814 ( .A(n1147), .B(n58812), .Z(n58811) );
  XNOR U58815 ( .A(p_input[97]), .B(n58813), .Z(n58812) );
  IV U58816 ( .A(p_input[65]), .Z(n58813) );
  XNOR U58817 ( .A(n57998), .B(n58806), .Z(n58808) );
  XNOR U58818 ( .A(p_input[1]), .B(n58814), .Z(n57998) );
  AND U58819 ( .A(n1144), .B(n58815), .Z(n58814) );
  XOR U58820 ( .A(p_input[33]), .B(p_input[1]), .Z(n58815) );
  IV U58821 ( .A(n58810), .Z(n58806) );
  AND U58822 ( .A(n58536), .B(n58539), .Z(n58810) );
  XOR U58823 ( .A(p_input[64]), .B(n58816), .Z(n58539) );
  AND U58824 ( .A(n1147), .B(n58817), .Z(n58816) );
  XOR U58825 ( .A(p_input[96]), .B(p_input[64]), .Z(n58817) );
  XOR U58826 ( .A(n58818), .B(n58819), .Z(n1147) );
  AND U58827 ( .A(n58820), .B(n58821), .Z(n58819) );
  XNOR U58828 ( .A(p_input[127]), .B(n58818), .Z(n58821) );
  XOR U58829 ( .A(n58818), .B(p_input[95]), .Z(n58820) );
  XOR U58830 ( .A(n58822), .B(n58823), .Z(n58818) );
  AND U58831 ( .A(n58824), .B(n58825), .Z(n58823) );
  XNOR U58832 ( .A(p_input[126]), .B(n58822), .Z(n58825) );
  XOR U58833 ( .A(n58822), .B(p_input[94]), .Z(n58824) );
  XOR U58834 ( .A(n58826), .B(n58827), .Z(n58822) );
  AND U58835 ( .A(n58828), .B(n58829), .Z(n58827) );
  XNOR U58836 ( .A(p_input[125]), .B(n58826), .Z(n58829) );
  XOR U58837 ( .A(n58826), .B(p_input[93]), .Z(n58828) );
  XOR U58838 ( .A(n58830), .B(n58831), .Z(n58826) );
  AND U58839 ( .A(n58832), .B(n58833), .Z(n58831) );
  XNOR U58840 ( .A(p_input[124]), .B(n58830), .Z(n58833) );
  XOR U58841 ( .A(n58830), .B(p_input[92]), .Z(n58832) );
  XOR U58842 ( .A(n58834), .B(n58835), .Z(n58830) );
  AND U58843 ( .A(n58836), .B(n58837), .Z(n58835) );
  XNOR U58844 ( .A(p_input[123]), .B(n58834), .Z(n58837) );
  XOR U58845 ( .A(n58834), .B(p_input[91]), .Z(n58836) );
  XOR U58846 ( .A(n58838), .B(n58839), .Z(n58834) );
  AND U58847 ( .A(n58840), .B(n58841), .Z(n58839) );
  XNOR U58848 ( .A(p_input[122]), .B(n58838), .Z(n58841) );
  XOR U58849 ( .A(n58838), .B(p_input[90]), .Z(n58840) );
  XOR U58850 ( .A(n58842), .B(n58843), .Z(n58838) );
  AND U58851 ( .A(n58844), .B(n58845), .Z(n58843) );
  XNOR U58852 ( .A(p_input[121]), .B(n58842), .Z(n58845) );
  XOR U58853 ( .A(n58842), .B(p_input[89]), .Z(n58844) );
  XOR U58854 ( .A(n58846), .B(n58847), .Z(n58842) );
  AND U58855 ( .A(n58848), .B(n58849), .Z(n58847) );
  XNOR U58856 ( .A(p_input[120]), .B(n58846), .Z(n58849) );
  XOR U58857 ( .A(n58846), .B(p_input[88]), .Z(n58848) );
  XOR U58858 ( .A(n58850), .B(n58851), .Z(n58846) );
  AND U58859 ( .A(n58852), .B(n58853), .Z(n58851) );
  XNOR U58860 ( .A(p_input[119]), .B(n58850), .Z(n58853) );
  XOR U58861 ( .A(n58850), .B(p_input[87]), .Z(n58852) );
  XOR U58862 ( .A(n58854), .B(n58855), .Z(n58850) );
  AND U58863 ( .A(n58856), .B(n58857), .Z(n58855) );
  XNOR U58864 ( .A(p_input[118]), .B(n58854), .Z(n58857) );
  XOR U58865 ( .A(n58854), .B(p_input[86]), .Z(n58856) );
  XOR U58866 ( .A(n58858), .B(n58859), .Z(n58854) );
  AND U58867 ( .A(n58860), .B(n58861), .Z(n58859) );
  XNOR U58868 ( .A(p_input[117]), .B(n58858), .Z(n58861) );
  XOR U58869 ( .A(n58858), .B(p_input[85]), .Z(n58860) );
  XOR U58870 ( .A(n58862), .B(n58863), .Z(n58858) );
  AND U58871 ( .A(n58864), .B(n58865), .Z(n58863) );
  XNOR U58872 ( .A(p_input[116]), .B(n58862), .Z(n58865) );
  XOR U58873 ( .A(n58862), .B(p_input[84]), .Z(n58864) );
  XOR U58874 ( .A(n58866), .B(n58867), .Z(n58862) );
  AND U58875 ( .A(n58868), .B(n58869), .Z(n58867) );
  XNOR U58876 ( .A(p_input[115]), .B(n58866), .Z(n58869) );
  XOR U58877 ( .A(n58866), .B(p_input[83]), .Z(n58868) );
  XOR U58878 ( .A(n58870), .B(n58871), .Z(n58866) );
  AND U58879 ( .A(n58872), .B(n58873), .Z(n58871) );
  XNOR U58880 ( .A(p_input[114]), .B(n58870), .Z(n58873) );
  XOR U58881 ( .A(n58870), .B(p_input[82]), .Z(n58872) );
  XOR U58882 ( .A(n58874), .B(n58875), .Z(n58870) );
  AND U58883 ( .A(n58876), .B(n58877), .Z(n58875) );
  XNOR U58884 ( .A(p_input[113]), .B(n58874), .Z(n58877) );
  XOR U58885 ( .A(n58874), .B(p_input[81]), .Z(n58876) );
  XOR U58886 ( .A(n58878), .B(n58879), .Z(n58874) );
  AND U58887 ( .A(n58880), .B(n58881), .Z(n58879) );
  XNOR U58888 ( .A(p_input[112]), .B(n58878), .Z(n58881) );
  XOR U58889 ( .A(n58878), .B(p_input[80]), .Z(n58880) );
  XOR U58890 ( .A(n58882), .B(n58883), .Z(n58878) );
  AND U58891 ( .A(n58884), .B(n58885), .Z(n58883) );
  XNOR U58892 ( .A(p_input[111]), .B(n58882), .Z(n58885) );
  XOR U58893 ( .A(n58882), .B(p_input[79]), .Z(n58884) );
  XOR U58894 ( .A(n58886), .B(n58887), .Z(n58882) );
  AND U58895 ( .A(n58888), .B(n58889), .Z(n58887) );
  XNOR U58896 ( .A(p_input[110]), .B(n58886), .Z(n58889) );
  XOR U58897 ( .A(n58886), .B(p_input[78]), .Z(n58888) );
  XOR U58898 ( .A(n58890), .B(n58891), .Z(n58886) );
  AND U58899 ( .A(n58892), .B(n58893), .Z(n58891) );
  XNOR U58900 ( .A(p_input[109]), .B(n58890), .Z(n58893) );
  XOR U58901 ( .A(n58890), .B(p_input[77]), .Z(n58892) );
  XOR U58902 ( .A(n58894), .B(n58895), .Z(n58890) );
  AND U58903 ( .A(n58896), .B(n58897), .Z(n58895) );
  XNOR U58904 ( .A(p_input[108]), .B(n58894), .Z(n58897) );
  XOR U58905 ( .A(n58894), .B(p_input[76]), .Z(n58896) );
  XOR U58906 ( .A(n58898), .B(n58899), .Z(n58894) );
  AND U58907 ( .A(n58900), .B(n58901), .Z(n58899) );
  XNOR U58908 ( .A(p_input[107]), .B(n58898), .Z(n58901) );
  XOR U58909 ( .A(n58898), .B(p_input[75]), .Z(n58900) );
  XOR U58910 ( .A(n58902), .B(n58903), .Z(n58898) );
  AND U58911 ( .A(n58904), .B(n58905), .Z(n58903) );
  XNOR U58912 ( .A(p_input[106]), .B(n58902), .Z(n58905) );
  XOR U58913 ( .A(n58902), .B(p_input[74]), .Z(n58904) );
  XOR U58914 ( .A(n58906), .B(n58907), .Z(n58902) );
  AND U58915 ( .A(n58908), .B(n58909), .Z(n58907) );
  XNOR U58916 ( .A(p_input[105]), .B(n58906), .Z(n58909) );
  XOR U58917 ( .A(n58906), .B(p_input[73]), .Z(n58908) );
  XOR U58918 ( .A(n58910), .B(n58911), .Z(n58906) );
  AND U58919 ( .A(n58912), .B(n58913), .Z(n58911) );
  XNOR U58920 ( .A(p_input[104]), .B(n58910), .Z(n58913) );
  XOR U58921 ( .A(n58910), .B(p_input[72]), .Z(n58912) );
  XOR U58922 ( .A(n58914), .B(n58915), .Z(n58910) );
  AND U58923 ( .A(n58916), .B(n58917), .Z(n58915) );
  XNOR U58924 ( .A(p_input[103]), .B(n58914), .Z(n58917) );
  XOR U58925 ( .A(n58914), .B(p_input[71]), .Z(n58916) );
  XOR U58926 ( .A(n58918), .B(n58919), .Z(n58914) );
  AND U58927 ( .A(n58920), .B(n58921), .Z(n58919) );
  XNOR U58928 ( .A(p_input[102]), .B(n58918), .Z(n58921) );
  XOR U58929 ( .A(n58918), .B(p_input[70]), .Z(n58920) );
  XOR U58930 ( .A(n58922), .B(n58923), .Z(n58918) );
  AND U58931 ( .A(n58924), .B(n58925), .Z(n58923) );
  XNOR U58932 ( .A(p_input[101]), .B(n58922), .Z(n58925) );
  XOR U58933 ( .A(n58922), .B(p_input[69]), .Z(n58924) );
  XOR U58934 ( .A(n58926), .B(n58927), .Z(n58922) );
  AND U58935 ( .A(n58928), .B(n58929), .Z(n58927) );
  XNOR U58936 ( .A(p_input[100]), .B(n58926), .Z(n58929) );
  XOR U58937 ( .A(n58926), .B(p_input[68]), .Z(n58928) );
  XOR U58938 ( .A(n58930), .B(n58931), .Z(n58926) );
  AND U58939 ( .A(n58932), .B(n58933), .Z(n58931) );
  XNOR U58940 ( .A(p_input[99]), .B(n58930), .Z(n58933) );
  XOR U58941 ( .A(n58930), .B(p_input[67]), .Z(n58932) );
  XOR U58942 ( .A(n58934), .B(n58935), .Z(n58930) );
  AND U58943 ( .A(n58936), .B(n58937), .Z(n58935) );
  XNOR U58944 ( .A(p_input[98]), .B(n58934), .Z(n58937) );
  XOR U58945 ( .A(n58934), .B(p_input[66]), .Z(n58936) );
  XNOR U58946 ( .A(n58938), .B(n58939), .Z(n58934) );
  AND U58947 ( .A(n58940), .B(n58941), .Z(n58939) );
  XOR U58948 ( .A(p_input[97]), .B(n58938), .Z(n58941) );
  XNOR U58949 ( .A(p_input[65]), .B(n58938), .Z(n58940) );
  AND U58950 ( .A(p_input[96]), .B(n58942), .Z(n58938) );
  IV U58951 ( .A(p_input[64]), .Z(n58942) );
  XNOR U58952 ( .A(p_input[0]), .B(n58943), .Z(n58536) );
  AND U58953 ( .A(n1144), .B(n58944), .Z(n58943) );
  XOR U58954 ( .A(p_input[32]), .B(p_input[0]), .Z(n58944) );
  XOR U58955 ( .A(n58945), .B(n58946), .Z(n1144) );
  AND U58956 ( .A(n58947), .B(n58948), .Z(n58946) );
  XNOR U58957 ( .A(p_input[63]), .B(n58945), .Z(n58948) );
  XOR U58958 ( .A(n58945), .B(p_input[31]), .Z(n58947) );
  XOR U58959 ( .A(n58949), .B(n58950), .Z(n58945) );
  AND U58960 ( .A(n58951), .B(n58952), .Z(n58950) );
  XNOR U58961 ( .A(p_input[62]), .B(n58949), .Z(n58952) );
  XNOR U58962 ( .A(n58949), .B(n58551), .Z(n58951) );
  IV U58963 ( .A(p_input[30]), .Z(n58551) );
  XOR U58964 ( .A(n58953), .B(n58954), .Z(n58949) );
  AND U58965 ( .A(n58955), .B(n58956), .Z(n58954) );
  XNOR U58966 ( .A(p_input[61]), .B(n58953), .Z(n58956) );
  XNOR U58967 ( .A(n58953), .B(n58560), .Z(n58955) );
  IV U58968 ( .A(p_input[29]), .Z(n58560) );
  XOR U58969 ( .A(n58957), .B(n58958), .Z(n58953) );
  AND U58970 ( .A(n58959), .B(n58960), .Z(n58958) );
  XNOR U58971 ( .A(p_input[60]), .B(n58957), .Z(n58960) );
  XNOR U58972 ( .A(n58957), .B(n58569), .Z(n58959) );
  IV U58973 ( .A(p_input[28]), .Z(n58569) );
  XOR U58974 ( .A(n58961), .B(n58962), .Z(n58957) );
  AND U58975 ( .A(n58963), .B(n58964), .Z(n58962) );
  XNOR U58976 ( .A(p_input[59]), .B(n58961), .Z(n58964) );
  XNOR U58977 ( .A(n58961), .B(n58578), .Z(n58963) );
  IV U58978 ( .A(p_input[27]), .Z(n58578) );
  XOR U58979 ( .A(n58965), .B(n58966), .Z(n58961) );
  AND U58980 ( .A(n58967), .B(n58968), .Z(n58966) );
  XNOR U58981 ( .A(p_input[58]), .B(n58965), .Z(n58968) );
  XNOR U58982 ( .A(n58965), .B(n58587), .Z(n58967) );
  IV U58983 ( .A(p_input[26]), .Z(n58587) );
  XOR U58984 ( .A(n58969), .B(n58970), .Z(n58965) );
  AND U58985 ( .A(n58971), .B(n58972), .Z(n58970) );
  XNOR U58986 ( .A(p_input[57]), .B(n58969), .Z(n58972) );
  XNOR U58987 ( .A(n58969), .B(n58596), .Z(n58971) );
  IV U58988 ( .A(p_input[25]), .Z(n58596) );
  XOR U58989 ( .A(n58973), .B(n58974), .Z(n58969) );
  AND U58990 ( .A(n58975), .B(n58976), .Z(n58974) );
  XNOR U58991 ( .A(p_input[56]), .B(n58973), .Z(n58976) );
  XNOR U58992 ( .A(n58973), .B(n58605), .Z(n58975) );
  IV U58993 ( .A(p_input[24]), .Z(n58605) );
  XOR U58994 ( .A(n58977), .B(n58978), .Z(n58973) );
  AND U58995 ( .A(n58979), .B(n58980), .Z(n58978) );
  XNOR U58996 ( .A(p_input[55]), .B(n58977), .Z(n58980) );
  XNOR U58997 ( .A(n58977), .B(n58614), .Z(n58979) );
  IV U58998 ( .A(p_input[23]), .Z(n58614) );
  XOR U58999 ( .A(n58981), .B(n58982), .Z(n58977) );
  AND U59000 ( .A(n58983), .B(n58984), .Z(n58982) );
  XNOR U59001 ( .A(p_input[54]), .B(n58981), .Z(n58984) );
  XNOR U59002 ( .A(n58981), .B(n58623), .Z(n58983) );
  IV U59003 ( .A(p_input[22]), .Z(n58623) );
  XOR U59004 ( .A(n58985), .B(n58986), .Z(n58981) );
  AND U59005 ( .A(n58987), .B(n58988), .Z(n58986) );
  XNOR U59006 ( .A(p_input[53]), .B(n58985), .Z(n58988) );
  XNOR U59007 ( .A(n58985), .B(n58632), .Z(n58987) );
  IV U59008 ( .A(p_input[21]), .Z(n58632) );
  XOR U59009 ( .A(n58989), .B(n58990), .Z(n58985) );
  AND U59010 ( .A(n58991), .B(n58992), .Z(n58990) );
  XNOR U59011 ( .A(p_input[52]), .B(n58989), .Z(n58992) );
  XNOR U59012 ( .A(n58989), .B(n58641), .Z(n58991) );
  IV U59013 ( .A(p_input[20]), .Z(n58641) );
  XOR U59014 ( .A(n58993), .B(n58994), .Z(n58989) );
  AND U59015 ( .A(n58995), .B(n58996), .Z(n58994) );
  XNOR U59016 ( .A(p_input[51]), .B(n58993), .Z(n58996) );
  XNOR U59017 ( .A(n58993), .B(n58650), .Z(n58995) );
  IV U59018 ( .A(p_input[19]), .Z(n58650) );
  XOR U59019 ( .A(n58997), .B(n58998), .Z(n58993) );
  AND U59020 ( .A(n58999), .B(n59000), .Z(n58998) );
  XNOR U59021 ( .A(p_input[50]), .B(n58997), .Z(n59000) );
  XNOR U59022 ( .A(n58997), .B(n58659), .Z(n58999) );
  IV U59023 ( .A(p_input[18]), .Z(n58659) );
  XOR U59024 ( .A(n59001), .B(n59002), .Z(n58997) );
  AND U59025 ( .A(n59003), .B(n59004), .Z(n59002) );
  XNOR U59026 ( .A(p_input[49]), .B(n59001), .Z(n59004) );
  XNOR U59027 ( .A(n59001), .B(n58668), .Z(n59003) );
  IV U59028 ( .A(p_input[17]), .Z(n58668) );
  XOR U59029 ( .A(n59005), .B(n59006), .Z(n59001) );
  AND U59030 ( .A(n59007), .B(n59008), .Z(n59006) );
  XNOR U59031 ( .A(p_input[48]), .B(n59005), .Z(n59008) );
  XNOR U59032 ( .A(n59005), .B(n58677), .Z(n59007) );
  IV U59033 ( .A(p_input[16]), .Z(n58677) );
  XOR U59034 ( .A(n59009), .B(n59010), .Z(n59005) );
  AND U59035 ( .A(n59011), .B(n59012), .Z(n59010) );
  XNOR U59036 ( .A(p_input[47]), .B(n59009), .Z(n59012) );
  XNOR U59037 ( .A(n59009), .B(n58686), .Z(n59011) );
  IV U59038 ( .A(p_input[15]), .Z(n58686) );
  XOR U59039 ( .A(n59013), .B(n59014), .Z(n59009) );
  AND U59040 ( .A(n59015), .B(n59016), .Z(n59014) );
  XNOR U59041 ( .A(p_input[46]), .B(n59013), .Z(n59016) );
  XNOR U59042 ( .A(n59013), .B(n58695), .Z(n59015) );
  IV U59043 ( .A(p_input[14]), .Z(n58695) );
  XOR U59044 ( .A(n59017), .B(n59018), .Z(n59013) );
  AND U59045 ( .A(n59019), .B(n59020), .Z(n59018) );
  XNOR U59046 ( .A(p_input[45]), .B(n59017), .Z(n59020) );
  XNOR U59047 ( .A(n59017), .B(n58704), .Z(n59019) );
  IV U59048 ( .A(p_input[13]), .Z(n58704) );
  XOR U59049 ( .A(n59021), .B(n59022), .Z(n59017) );
  AND U59050 ( .A(n59023), .B(n59024), .Z(n59022) );
  XNOR U59051 ( .A(p_input[44]), .B(n59021), .Z(n59024) );
  XNOR U59052 ( .A(n59021), .B(n58713), .Z(n59023) );
  IV U59053 ( .A(p_input[12]), .Z(n58713) );
  XOR U59054 ( .A(n59025), .B(n59026), .Z(n59021) );
  AND U59055 ( .A(n59027), .B(n59028), .Z(n59026) );
  XNOR U59056 ( .A(p_input[43]), .B(n59025), .Z(n59028) );
  XNOR U59057 ( .A(n59025), .B(n58722), .Z(n59027) );
  IV U59058 ( .A(p_input[11]), .Z(n58722) );
  XOR U59059 ( .A(n59029), .B(n59030), .Z(n59025) );
  AND U59060 ( .A(n59031), .B(n59032), .Z(n59030) );
  XNOR U59061 ( .A(p_input[42]), .B(n59029), .Z(n59032) );
  XNOR U59062 ( .A(n59029), .B(n58731), .Z(n59031) );
  IV U59063 ( .A(p_input[10]), .Z(n58731) );
  XOR U59064 ( .A(n59033), .B(n59034), .Z(n59029) );
  AND U59065 ( .A(n59035), .B(n59036), .Z(n59034) );
  XNOR U59066 ( .A(p_input[41]), .B(n59033), .Z(n59036) );
  XNOR U59067 ( .A(n59033), .B(n58740), .Z(n59035) );
  IV U59068 ( .A(p_input[9]), .Z(n58740) );
  XOR U59069 ( .A(n59037), .B(n59038), .Z(n59033) );
  AND U59070 ( .A(n59039), .B(n59040), .Z(n59038) );
  XNOR U59071 ( .A(p_input[40]), .B(n59037), .Z(n59040) );
  XNOR U59072 ( .A(n59037), .B(n58749), .Z(n59039) );
  IV U59073 ( .A(p_input[8]), .Z(n58749) );
  XOR U59074 ( .A(n59041), .B(n59042), .Z(n59037) );
  AND U59075 ( .A(n59043), .B(n59044), .Z(n59042) );
  XNOR U59076 ( .A(p_input[39]), .B(n59041), .Z(n59044) );
  XNOR U59077 ( .A(n59041), .B(n58758), .Z(n59043) );
  IV U59078 ( .A(p_input[7]), .Z(n58758) );
  XOR U59079 ( .A(n59045), .B(n59046), .Z(n59041) );
  AND U59080 ( .A(n59047), .B(n59048), .Z(n59046) );
  XNOR U59081 ( .A(p_input[38]), .B(n59045), .Z(n59048) );
  XNOR U59082 ( .A(n59045), .B(n58767), .Z(n59047) );
  IV U59083 ( .A(p_input[6]), .Z(n58767) );
  XOR U59084 ( .A(n59049), .B(n59050), .Z(n59045) );
  AND U59085 ( .A(n59051), .B(n59052), .Z(n59050) );
  XNOR U59086 ( .A(p_input[37]), .B(n59049), .Z(n59052) );
  XNOR U59087 ( .A(n59049), .B(n58776), .Z(n59051) );
  IV U59088 ( .A(p_input[5]), .Z(n58776) );
  XOR U59089 ( .A(n59053), .B(n59054), .Z(n59049) );
  AND U59090 ( .A(n59055), .B(n59056), .Z(n59054) );
  XNOR U59091 ( .A(p_input[36]), .B(n59053), .Z(n59056) );
  XNOR U59092 ( .A(n59053), .B(n58785), .Z(n59055) );
  IV U59093 ( .A(p_input[4]), .Z(n58785) );
  XOR U59094 ( .A(n59057), .B(n59058), .Z(n59053) );
  AND U59095 ( .A(n59059), .B(n59060), .Z(n59058) );
  XNOR U59096 ( .A(p_input[35]), .B(n59057), .Z(n59060) );
  XNOR U59097 ( .A(n59057), .B(n58794), .Z(n59059) );
  IV U59098 ( .A(p_input[3]), .Z(n58794) );
  XOR U59099 ( .A(n59061), .B(n59062), .Z(n59057) );
  AND U59100 ( .A(n59063), .B(n59064), .Z(n59062) );
  XNOR U59101 ( .A(p_input[34]), .B(n59061), .Z(n59064) );
  XNOR U59102 ( .A(n59061), .B(n58803), .Z(n59063) );
  IV U59103 ( .A(p_input[2]), .Z(n58803) );
  XNOR U59104 ( .A(n59065), .B(n59066), .Z(n59061) );
  AND U59105 ( .A(n59067), .B(n59068), .Z(n59066) );
  XOR U59106 ( .A(p_input[33]), .B(n59065), .Z(n59068) );
  XNOR U59107 ( .A(p_input[1]), .B(n59065), .Z(n59067) );
  AND U59108 ( .A(p_input[32]), .B(n59069), .Z(n59065) );
  IV U59109 ( .A(p_input[0]), .Z(n59069) );
endmodule

